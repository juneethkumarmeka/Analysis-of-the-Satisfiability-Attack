module basic_1000_10000_1500_10_levels_10xor_1(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999;
nand U0 (N_0,In_160,In_53);
or U1 (N_1,In_55,In_948);
xnor U2 (N_2,In_776,In_422);
nor U3 (N_3,In_850,In_741);
nor U4 (N_4,In_381,In_870);
xnor U5 (N_5,In_211,In_472);
nor U6 (N_6,In_426,In_378);
nand U7 (N_7,In_563,In_33);
nor U8 (N_8,In_181,In_201);
nor U9 (N_9,In_78,In_102);
and U10 (N_10,In_159,In_128);
nand U11 (N_11,In_855,In_879);
or U12 (N_12,In_600,In_659);
or U13 (N_13,In_954,In_215);
nand U14 (N_14,In_272,In_788);
nand U15 (N_15,In_35,In_235);
and U16 (N_16,In_108,In_152);
xnor U17 (N_17,In_232,In_736);
xnor U18 (N_18,In_701,In_813);
xnor U19 (N_19,In_22,In_1);
or U20 (N_20,In_4,In_284);
xnor U21 (N_21,In_570,In_256);
and U22 (N_22,In_196,In_264);
nand U23 (N_23,In_873,In_591);
nor U24 (N_24,In_923,In_492);
xnor U25 (N_25,In_573,In_519);
xor U26 (N_26,In_603,In_351);
and U27 (N_27,In_302,In_314);
or U28 (N_28,In_937,In_347);
nand U29 (N_29,In_468,In_966);
nand U30 (N_30,In_892,In_738);
nor U31 (N_31,In_987,In_764);
nand U32 (N_32,In_312,In_491);
nor U33 (N_33,In_864,In_599);
or U34 (N_34,In_276,In_438);
and U35 (N_35,In_993,In_151);
nand U36 (N_36,In_714,In_79);
nand U37 (N_37,In_625,In_619);
nor U38 (N_38,In_127,In_867);
or U39 (N_39,In_396,In_739);
nand U40 (N_40,In_118,In_546);
nor U41 (N_41,In_495,In_214);
nand U42 (N_42,In_432,In_157);
or U43 (N_43,In_985,In_901);
nand U44 (N_44,In_863,In_928);
nand U45 (N_45,In_847,In_47);
and U46 (N_46,In_56,In_656);
xor U47 (N_47,In_226,In_655);
nor U48 (N_48,In_222,In_877);
nand U49 (N_49,In_476,In_992);
or U50 (N_50,In_130,In_690);
nand U51 (N_51,In_524,In_915);
nand U52 (N_52,In_882,In_433);
nor U53 (N_53,In_355,In_558);
nand U54 (N_54,In_750,In_303);
xor U55 (N_55,In_149,In_729);
nand U56 (N_56,In_178,In_539);
xnor U57 (N_57,In_971,In_323);
nand U58 (N_58,In_114,In_747);
or U59 (N_59,In_192,In_38);
xor U60 (N_60,In_672,In_854);
nand U61 (N_61,In_846,In_2);
nor U62 (N_62,In_359,In_231);
or U63 (N_63,In_150,In_481);
nand U64 (N_64,In_28,In_541);
nand U65 (N_65,In_113,In_562);
nor U66 (N_66,In_278,In_91);
or U67 (N_67,In_169,In_477);
nor U68 (N_68,In_994,In_857);
and U69 (N_69,In_129,In_485);
or U70 (N_70,In_945,In_975);
or U71 (N_71,In_990,In_259);
and U72 (N_72,In_221,In_121);
xnor U73 (N_73,In_429,In_779);
nand U74 (N_74,In_550,In_699);
xnor U75 (N_75,In_875,In_759);
xnor U76 (N_76,In_988,In_430);
and U77 (N_77,In_934,In_380);
xnor U78 (N_78,In_164,In_397);
and U79 (N_79,In_82,In_122);
nand U80 (N_80,In_271,In_100);
or U81 (N_81,In_958,In_978);
nor U82 (N_82,In_838,In_266);
nand U83 (N_83,In_290,In_880);
nand U84 (N_84,In_329,In_564);
nand U85 (N_85,In_131,In_924);
nand U86 (N_86,In_249,In_810);
and U87 (N_87,In_860,In_876);
nor U88 (N_88,In_182,In_483);
nand U89 (N_89,In_703,In_856);
xor U90 (N_90,In_289,In_452);
nor U91 (N_91,In_6,In_50);
nor U92 (N_92,In_417,In_777);
xor U93 (N_93,In_908,In_252);
or U94 (N_94,In_306,In_427);
xor U95 (N_95,In_853,In_658);
xor U96 (N_96,In_205,In_488);
and U97 (N_97,In_138,In_5);
and U98 (N_98,In_409,In_280);
nand U99 (N_99,In_845,In_581);
or U100 (N_100,In_177,In_935);
nor U101 (N_101,In_700,In_733);
nor U102 (N_102,In_645,In_243);
nand U103 (N_103,In_447,In_115);
or U104 (N_104,In_315,In_957);
nor U105 (N_105,In_773,In_156);
and U106 (N_106,In_512,In_44);
or U107 (N_107,In_155,In_92);
nand U108 (N_108,In_808,In_520);
xor U109 (N_109,In_852,In_939);
nand U110 (N_110,In_745,In_633);
and U111 (N_111,In_202,In_394);
xor U112 (N_112,In_926,In_567);
nor U113 (N_113,In_571,In_916);
nor U114 (N_114,In_525,In_842);
nand U115 (N_115,In_18,In_363);
nor U116 (N_116,In_498,In_905);
nor U117 (N_117,In_677,In_542);
nand U118 (N_118,In_976,In_653);
and U119 (N_119,In_610,In_360);
nand U120 (N_120,In_757,In_999);
or U121 (N_121,In_95,In_722);
or U122 (N_122,In_348,In_187);
xnor U123 (N_123,In_240,In_829);
nand U124 (N_124,In_774,In_642);
or U125 (N_125,In_93,In_210);
or U126 (N_126,In_490,In_967);
and U127 (N_127,In_494,In_596);
xnor U128 (N_128,In_902,In_531);
nand U129 (N_129,In_503,In_42);
xnor U130 (N_130,In_101,In_732);
or U131 (N_131,In_449,In_273);
nor U132 (N_132,In_899,In_62);
xor U133 (N_133,In_995,In_41);
nand U134 (N_134,In_316,In_12);
or U135 (N_135,In_478,In_909);
or U136 (N_136,In_604,In_184);
and U137 (N_137,In_644,In_237);
or U138 (N_138,In_116,In_301);
xnor U139 (N_139,In_465,In_711);
nor U140 (N_140,In_505,In_811);
and U141 (N_141,In_960,In_756);
nor U142 (N_142,In_986,In_720);
nor U143 (N_143,In_444,In_285);
or U144 (N_144,In_803,In_96);
and U145 (N_145,In_245,In_470);
and U146 (N_146,In_34,In_442);
nand U147 (N_147,In_998,In_622);
nor U148 (N_148,In_357,In_896);
and U149 (N_149,In_223,In_330);
nand U150 (N_150,In_372,In_588);
xnor U151 (N_151,In_668,In_8);
nor U152 (N_152,In_766,In_453);
xnor U153 (N_153,In_724,In_293);
and U154 (N_154,In_545,In_540);
nor U155 (N_155,In_250,In_175);
xor U156 (N_156,In_612,In_61);
or U157 (N_157,In_806,In_383);
nand U158 (N_158,In_63,In_286);
xnor U159 (N_159,In_632,In_337);
and U160 (N_160,In_922,In_36);
nor U161 (N_161,In_415,In_959);
nor U162 (N_162,In_740,In_40);
xnor U163 (N_163,In_715,In_74);
or U164 (N_164,In_514,In_549);
xnor U165 (N_165,In_784,In_669);
nand U166 (N_166,In_207,In_173);
or U167 (N_167,In_972,In_809);
or U168 (N_168,In_464,In_39);
nand U169 (N_169,In_538,In_327);
and U170 (N_170,In_961,In_30);
or U171 (N_171,In_627,In_869);
and U172 (N_172,In_20,In_946);
nand U173 (N_173,In_137,In_933);
and U174 (N_174,In_601,In_718);
nand U175 (N_175,In_927,In_818);
and U176 (N_176,In_375,In_942);
and U177 (N_177,In_25,In_459);
and U178 (N_178,In_313,In_194);
nor U179 (N_179,In_537,In_70);
nor U180 (N_180,In_413,In_404);
or U181 (N_181,In_532,In_613);
or U182 (N_182,In_765,In_799);
and U183 (N_183,In_621,In_435);
and U184 (N_184,In_421,In_769);
or U185 (N_185,In_792,In_480);
nand U186 (N_186,In_457,In_172);
xor U187 (N_187,In_382,In_410);
nor U188 (N_188,In_517,In_296);
nor U189 (N_189,In_735,In_812);
and U190 (N_190,In_979,In_213);
and U191 (N_191,In_667,In_338);
nand U192 (N_192,In_257,In_258);
xor U193 (N_193,In_572,In_768);
and U194 (N_194,In_88,In_721);
nor U195 (N_195,In_815,In_665);
nand U196 (N_196,In_199,In_414);
nand U197 (N_197,In_52,In_328);
or U198 (N_198,In_636,In_681);
nand U199 (N_199,In_43,In_795);
nor U200 (N_200,In_191,In_955);
nor U201 (N_201,In_696,In_746);
nor U202 (N_202,In_179,In_661);
nor U203 (N_203,In_166,In_439);
or U204 (N_204,In_475,In_797);
nor U205 (N_205,In_220,In_448);
and U206 (N_206,In_962,In_597);
and U207 (N_207,In_111,In_650);
nor U208 (N_208,In_965,In_405);
xnor U209 (N_209,In_502,In_450);
xnor U210 (N_210,In_85,In_866);
nand U211 (N_211,In_474,In_910);
or U212 (N_212,In_268,In_657);
and U213 (N_213,In_731,In_224);
or U214 (N_214,In_824,In_865);
nand U215 (N_215,In_605,In_14);
or U216 (N_216,In_443,In_592);
nand U217 (N_217,In_639,In_99);
and U218 (N_218,In_200,In_489);
and U219 (N_219,In_791,In_473);
or U220 (N_220,In_743,In_536);
nor U221 (N_221,In_446,In_590);
or U222 (N_222,In_834,In_90);
or U223 (N_223,In_456,In_664);
nor U224 (N_224,In_107,In_814);
xor U225 (N_225,In_663,In_911);
and U226 (N_226,In_886,In_727);
and U227 (N_227,In_823,In_557);
nand U228 (N_228,In_325,In_526);
xnor U229 (N_229,In_789,In_707);
nand U230 (N_230,In_618,In_333);
nand U231 (N_231,In_120,In_75);
xnor U232 (N_232,In_734,In_726);
nand U233 (N_233,In_13,In_135);
nor U234 (N_234,In_343,In_335);
xor U235 (N_235,In_291,In_298);
and U236 (N_236,In_511,In_602);
nand U237 (N_237,In_80,In_785);
or U238 (N_238,In_826,In_407);
or U239 (N_239,In_804,In_830);
nor U240 (N_240,In_951,In_680);
nor U241 (N_241,In_180,In_903);
or U242 (N_242,In_940,In_686);
xnor U243 (N_243,In_676,In_145);
or U244 (N_244,In_796,In_518);
or U245 (N_245,In_529,In_970);
or U246 (N_246,In_165,In_522);
xor U247 (N_247,In_648,In_793);
nor U248 (N_248,In_68,In_820);
xnor U249 (N_249,In_460,In_932);
nor U250 (N_250,In_832,In_698);
nor U251 (N_251,In_533,In_119);
or U252 (N_252,In_772,In_168);
or U253 (N_253,In_914,In_471);
or U254 (N_254,In_624,In_246);
and U255 (N_255,In_654,In_72);
and U256 (N_256,In_188,In_705);
nand U257 (N_257,In_358,In_19);
nand U258 (N_258,In_637,In_949);
nand U259 (N_259,In_354,In_373);
and U260 (N_260,In_693,In_559);
nand U261 (N_261,In_279,In_390);
xor U262 (N_262,In_682,In_29);
nand U263 (N_263,In_629,In_305);
nand U264 (N_264,In_780,In_640);
or U265 (N_265,In_261,In_260);
nor U266 (N_266,In_831,In_649);
or U267 (N_267,In_283,In_606);
nor U268 (N_268,In_320,In_938);
and U269 (N_269,In_493,In_379);
xor U270 (N_270,In_952,In_614);
or U271 (N_271,In_46,In_479);
xor U272 (N_272,In_675,In_125);
or U273 (N_273,In_717,In_913);
nand U274 (N_274,In_974,In_781);
nor U275 (N_275,In_827,In_255);
and U276 (N_276,In_977,In_263);
and U277 (N_277,In_27,In_436);
nor U278 (N_278,In_311,In_595);
xor U279 (N_279,In_146,In_197);
and U280 (N_280,In_352,In_218);
xnor U281 (N_281,In_560,In_349);
or U282 (N_282,In_620,In_425);
nor U283 (N_283,In_837,In_84);
xnor U284 (N_284,In_535,In_611);
xor U285 (N_285,In_798,In_32);
and U286 (N_286,In_185,In_692);
nor U287 (N_287,In_944,In_434);
nor U288 (N_288,In_134,In_893);
nor U289 (N_289,In_907,In_49);
and U290 (N_290,In_345,In_384);
or U291 (N_291,In_919,In_616);
or U292 (N_292,In_819,In_513);
nor U293 (N_293,In_755,In_859);
nor U294 (N_294,In_651,In_751);
or U295 (N_295,In_767,In_984);
and U296 (N_296,In_275,In_297);
or U297 (N_297,In_497,In_728);
nand U298 (N_298,In_684,In_7);
or U299 (N_299,In_300,In_318);
nor U300 (N_300,In_506,In_891);
or U301 (N_301,In_76,In_890);
nand U302 (N_302,In_399,In_282);
nand U303 (N_303,In_760,In_515);
nor U304 (N_304,In_148,In_694);
nor U305 (N_305,In_752,In_11);
and U306 (N_306,In_17,In_816);
or U307 (N_307,In_411,In_917);
and U308 (N_308,In_981,In_635);
nand U309 (N_309,In_241,In_678);
and U310 (N_310,In_805,In_445);
nor U311 (N_311,In_801,In_10);
xnor U312 (N_312,In_615,In_208);
xor U313 (N_313,In_139,In_86);
xnor U314 (N_314,In_59,In_144);
nor U315 (N_315,In_212,In_983);
nor U316 (N_316,In_871,In_190);
and U317 (N_317,In_548,In_16);
xnor U318 (N_318,In_771,In_868);
or U319 (N_319,In_786,In_238);
xnor U320 (N_320,In_802,In_454);
nor U321 (N_321,In_523,In_841);
xnor U322 (N_322,In_183,In_60);
and U323 (N_323,In_964,In_527);
nand U324 (N_324,In_626,In_790);
and U325 (N_325,In_561,In_496);
nand U326 (N_326,In_69,In_265);
and U327 (N_327,In_424,In_216);
nor U328 (N_328,In_670,In_206);
xnor U329 (N_329,In_304,In_953);
and U330 (N_330,In_292,In_376);
and U331 (N_331,In_594,In_991);
or U332 (N_332,In_554,In_929);
or U333 (N_333,In_585,In_883);
xor U334 (N_334,In_671,In_825);
or U335 (N_335,In_881,In_507);
nor U336 (N_336,In_132,In_336);
nor U337 (N_337,In_725,In_377);
nor U338 (N_338,In_689,In_844);
and U339 (N_339,In_467,In_37);
nor U340 (N_340,In_341,In_849);
nor U341 (N_341,In_712,In_709);
and U342 (N_342,In_609,In_888);
and U343 (N_343,In_912,In_420);
nor U344 (N_344,In_71,In_24);
and U345 (N_345,In_904,In_307);
and U346 (N_346,In_242,In_136);
xnor U347 (N_347,In_925,In_23);
nor U348 (N_348,In_673,In_385);
nor U349 (N_349,In_73,In_294);
nor U350 (N_350,In_862,In_687);
or U351 (N_351,In_392,In_254);
xnor U352 (N_352,In_638,In_339);
and U353 (N_353,In_142,In_288);
or U354 (N_354,In_455,In_921);
or U355 (N_355,In_509,In_486);
or U356 (N_356,In_186,In_848);
or U357 (N_357,In_583,In_287);
xor U358 (N_358,In_487,In_94);
nand U359 (N_359,In_274,In_387);
or U360 (N_360,In_482,In_577);
nand U361 (N_361,In_817,In_451);
or U362 (N_362,In_501,In_401);
and U363 (N_363,In_646,In_106);
nor U364 (N_364,In_586,In_758);
xnor U365 (N_365,In_851,In_887);
or U366 (N_366,In_81,In_406);
xnor U367 (N_367,In_269,In_389);
and U368 (N_368,In_982,In_783);
xor U369 (N_369,In_299,In_141);
xnor U370 (N_370,In_956,In_950);
nor U371 (N_371,In_836,In_652);
nor U372 (N_372,In_872,In_0);
and U373 (N_373,In_229,In_326);
nand U374 (N_374,In_695,In_9);
and U375 (N_375,In_551,In_716);
xor U376 (N_376,In_174,In_204);
xnor U377 (N_377,In_463,In_861);
nor U378 (N_378,In_147,In_388);
xor U379 (N_379,In_688,In_217);
and U380 (N_380,In_97,In_930);
or U381 (N_381,In_57,In_143);
xnor U382 (N_382,In_331,In_441);
or U383 (N_383,In_484,In_508);
nor U384 (N_384,In_225,In_973);
nand U385 (N_385,In_770,In_947);
and U386 (N_386,In_516,In_374);
xnor U387 (N_387,In_170,In_126);
nand U388 (N_388,In_674,In_219);
and U389 (N_389,In_361,In_344);
xnor U390 (N_390,In_15,In_340);
nor U391 (N_391,In_666,In_628);
xor U392 (N_392,In_462,In_247);
or U393 (N_393,In_920,In_176);
nor U394 (N_394,In_353,In_569);
and U395 (N_395,In_500,In_158);
nor U396 (N_396,In_858,In_321);
xnor U397 (N_397,In_369,In_277);
xnor U398 (N_398,In_308,In_575);
xnor U399 (N_399,In_748,In_897);
nand U400 (N_400,In_54,In_310);
xnor U401 (N_401,In_706,In_763);
nor U402 (N_402,In_133,In_153);
nor U403 (N_403,In_440,In_742);
nor U404 (N_404,In_634,In_236);
and U405 (N_405,In_461,In_83);
nor U406 (N_406,In_104,In_840);
and U407 (N_407,In_356,In_45);
or U408 (N_408,In_775,In_889);
and U409 (N_409,In_87,In_77);
nand U410 (N_410,In_51,In_608);
xor U411 (N_411,In_895,In_364);
nand U412 (N_412,In_267,In_556);
or U413 (N_413,In_193,In_21);
and U414 (N_414,In_794,In_112);
and U415 (N_415,In_822,In_346);
or U416 (N_416,In_281,In_64);
or U417 (N_417,In_547,In_579);
nand U418 (N_418,In_617,In_140);
and U419 (N_419,In_968,In_552);
and U420 (N_420,In_408,In_350);
nand U421 (N_421,In_574,In_874);
nand U422 (N_422,In_737,In_26);
or U423 (N_423,In_839,In_761);
xnor U424 (N_424,In_253,In_702);
nand U425 (N_425,In_233,In_662);
or U426 (N_426,In_386,In_553);
and U427 (N_427,In_400,In_431);
or U428 (N_428,In_109,In_393);
xnor U429 (N_429,In_368,In_969);
or U430 (N_430,In_641,In_989);
and U431 (N_431,In_807,In_568);
nor U432 (N_432,In_898,In_458);
or U433 (N_433,In_931,In_117);
nor U434 (N_434,In_469,In_370);
xor U435 (N_435,In_593,In_821);
or U436 (N_436,In_48,In_203);
nor U437 (N_437,In_248,In_787);
xnor U438 (N_438,In_366,In_828);
or U439 (N_439,In_402,In_528);
nor U440 (N_440,In_322,In_744);
and U441 (N_441,In_623,In_521);
or U442 (N_442,In_660,In_607);
xnor U443 (N_443,In_209,In_227);
and U444 (N_444,In_884,In_3);
nor U445 (N_445,In_324,In_423);
nand U446 (N_446,In_710,In_365);
nor U447 (N_447,In_504,In_67);
nor U448 (N_448,In_943,In_403);
nor U449 (N_449,In_543,In_189);
or U450 (N_450,In_997,In_162);
xor U451 (N_451,In_510,In_171);
or U452 (N_452,In_123,In_412);
nand U453 (N_453,In_371,In_587);
or U454 (N_454,In_835,In_643);
and U455 (N_455,In_228,In_565);
and U456 (N_456,In_391,In_582);
and U457 (N_457,In_418,In_918);
and U458 (N_458,In_124,In_906);
and U459 (N_459,In_941,In_395);
xor U460 (N_460,In_154,In_198);
or U461 (N_461,In_270,In_367);
nand U462 (N_462,In_584,In_578);
and U463 (N_463,In_244,In_530);
or U464 (N_464,In_334,In_894);
and U465 (N_465,In_782,In_980);
nor U466 (N_466,In_58,In_566);
xnor U467 (N_467,In_239,In_723);
and U468 (N_468,In_885,In_309);
nand U469 (N_469,In_89,In_598);
and U470 (N_470,In_996,In_555);
nand U471 (N_471,In_534,In_936);
or U472 (N_472,In_833,In_362);
nand U473 (N_473,In_685,In_437);
nand U474 (N_474,In_589,In_631);
nor U475 (N_475,In_580,In_262);
or U476 (N_476,In_466,In_163);
nor U477 (N_477,In_98,In_753);
or U478 (N_478,In_499,In_105);
xnor U479 (N_479,In_230,In_167);
nor U480 (N_480,In_697,In_963);
or U481 (N_481,In_319,In_65);
nor U482 (N_482,In_398,In_762);
nand U483 (N_483,In_103,In_416);
and U484 (N_484,In_843,In_544);
and U485 (N_485,In_778,In_295);
nand U486 (N_486,In_251,In_708);
nor U487 (N_487,In_878,In_110);
nand U488 (N_488,In_749,In_713);
or U489 (N_489,In_332,In_428);
nor U490 (N_490,In_576,In_630);
and U491 (N_491,In_900,In_691);
or U492 (N_492,In_647,In_342);
or U493 (N_493,In_679,In_800);
nor U494 (N_494,In_754,In_31);
nor U495 (N_495,In_730,In_195);
nand U496 (N_496,In_683,In_234);
nor U497 (N_497,In_419,In_161);
xnor U498 (N_498,In_66,In_719);
xnor U499 (N_499,In_317,In_704);
xor U500 (N_500,In_713,In_821);
and U501 (N_501,In_493,In_840);
nand U502 (N_502,In_786,In_964);
and U503 (N_503,In_914,In_627);
nand U504 (N_504,In_128,In_183);
nor U505 (N_505,In_793,In_632);
xnor U506 (N_506,In_305,In_751);
xnor U507 (N_507,In_224,In_362);
and U508 (N_508,In_890,In_292);
and U509 (N_509,In_629,In_372);
xnor U510 (N_510,In_527,In_444);
xnor U511 (N_511,In_541,In_428);
and U512 (N_512,In_403,In_169);
or U513 (N_513,In_929,In_276);
and U514 (N_514,In_14,In_177);
nor U515 (N_515,In_16,In_806);
xnor U516 (N_516,In_348,In_222);
xnor U517 (N_517,In_285,In_700);
nand U518 (N_518,In_253,In_709);
nor U519 (N_519,In_223,In_712);
nand U520 (N_520,In_529,In_436);
and U521 (N_521,In_486,In_5);
or U522 (N_522,In_3,In_418);
nand U523 (N_523,In_538,In_273);
nor U524 (N_524,In_623,In_711);
nor U525 (N_525,In_810,In_191);
xnor U526 (N_526,In_435,In_553);
and U527 (N_527,In_56,In_410);
and U528 (N_528,In_827,In_872);
or U529 (N_529,In_361,In_978);
or U530 (N_530,In_121,In_909);
nor U531 (N_531,In_725,In_642);
nand U532 (N_532,In_733,In_949);
nor U533 (N_533,In_31,In_46);
nor U534 (N_534,In_664,In_413);
nor U535 (N_535,In_827,In_18);
xnor U536 (N_536,In_965,In_43);
xor U537 (N_537,In_755,In_813);
nor U538 (N_538,In_954,In_574);
or U539 (N_539,In_666,In_577);
xnor U540 (N_540,In_901,In_567);
or U541 (N_541,In_951,In_639);
xor U542 (N_542,In_254,In_810);
or U543 (N_543,In_309,In_823);
and U544 (N_544,In_480,In_360);
xor U545 (N_545,In_406,In_86);
and U546 (N_546,In_638,In_38);
xnor U547 (N_547,In_809,In_321);
nand U548 (N_548,In_303,In_178);
nor U549 (N_549,In_524,In_399);
nand U550 (N_550,In_570,In_216);
and U551 (N_551,In_575,In_57);
nor U552 (N_552,In_160,In_817);
nand U553 (N_553,In_518,In_650);
nand U554 (N_554,In_230,In_527);
and U555 (N_555,In_517,In_727);
or U556 (N_556,In_284,In_363);
xor U557 (N_557,In_129,In_65);
nand U558 (N_558,In_305,In_942);
or U559 (N_559,In_870,In_792);
xnor U560 (N_560,In_809,In_297);
xnor U561 (N_561,In_446,In_10);
nand U562 (N_562,In_530,In_871);
nand U563 (N_563,In_386,In_260);
nand U564 (N_564,In_553,In_793);
xnor U565 (N_565,In_151,In_373);
nor U566 (N_566,In_229,In_48);
and U567 (N_567,In_178,In_405);
nor U568 (N_568,In_802,In_925);
or U569 (N_569,In_486,In_411);
xnor U570 (N_570,In_612,In_185);
and U571 (N_571,In_256,In_182);
xnor U572 (N_572,In_870,In_658);
or U573 (N_573,In_815,In_436);
or U574 (N_574,In_391,In_923);
xnor U575 (N_575,In_610,In_554);
xor U576 (N_576,In_738,In_435);
xor U577 (N_577,In_626,In_43);
nor U578 (N_578,In_549,In_86);
nor U579 (N_579,In_447,In_227);
xor U580 (N_580,In_716,In_803);
and U581 (N_581,In_445,In_232);
or U582 (N_582,In_89,In_846);
or U583 (N_583,In_475,In_695);
xnor U584 (N_584,In_983,In_708);
nor U585 (N_585,In_484,In_523);
and U586 (N_586,In_201,In_486);
and U587 (N_587,In_209,In_585);
or U588 (N_588,In_641,In_555);
nor U589 (N_589,In_825,In_868);
nor U590 (N_590,In_981,In_849);
and U591 (N_591,In_136,In_542);
or U592 (N_592,In_23,In_147);
nand U593 (N_593,In_112,In_770);
and U594 (N_594,In_686,In_680);
nand U595 (N_595,In_324,In_422);
nand U596 (N_596,In_483,In_42);
or U597 (N_597,In_104,In_914);
nand U598 (N_598,In_208,In_618);
and U599 (N_599,In_845,In_301);
nor U600 (N_600,In_494,In_369);
or U601 (N_601,In_492,In_934);
nor U602 (N_602,In_401,In_170);
xnor U603 (N_603,In_252,In_293);
xnor U604 (N_604,In_724,In_350);
xnor U605 (N_605,In_994,In_498);
nor U606 (N_606,In_700,In_891);
nor U607 (N_607,In_903,In_820);
and U608 (N_608,In_495,In_18);
nand U609 (N_609,In_7,In_774);
or U610 (N_610,In_822,In_976);
nand U611 (N_611,In_272,In_546);
and U612 (N_612,In_664,In_622);
nor U613 (N_613,In_290,In_96);
xnor U614 (N_614,In_638,In_471);
nand U615 (N_615,In_279,In_437);
and U616 (N_616,In_977,In_280);
nor U617 (N_617,In_937,In_279);
nor U618 (N_618,In_5,In_306);
and U619 (N_619,In_45,In_501);
or U620 (N_620,In_494,In_566);
or U621 (N_621,In_578,In_357);
nor U622 (N_622,In_212,In_122);
and U623 (N_623,In_523,In_747);
or U624 (N_624,In_939,In_20);
xnor U625 (N_625,In_115,In_306);
or U626 (N_626,In_831,In_676);
nand U627 (N_627,In_574,In_857);
xnor U628 (N_628,In_364,In_315);
nor U629 (N_629,In_317,In_758);
nor U630 (N_630,In_843,In_292);
nor U631 (N_631,In_511,In_81);
or U632 (N_632,In_266,In_900);
and U633 (N_633,In_749,In_791);
nor U634 (N_634,In_611,In_168);
nand U635 (N_635,In_925,In_968);
nand U636 (N_636,In_728,In_240);
and U637 (N_637,In_438,In_131);
or U638 (N_638,In_700,In_737);
xnor U639 (N_639,In_970,In_917);
nor U640 (N_640,In_55,In_776);
xor U641 (N_641,In_829,In_801);
nand U642 (N_642,In_906,In_44);
nor U643 (N_643,In_194,In_705);
and U644 (N_644,In_184,In_185);
nand U645 (N_645,In_927,In_836);
nand U646 (N_646,In_212,In_796);
xnor U647 (N_647,In_412,In_541);
xor U648 (N_648,In_902,In_642);
and U649 (N_649,In_152,In_488);
or U650 (N_650,In_976,In_111);
nor U651 (N_651,In_514,In_773);
xor U652 (N_652,In_728,In_614);
nand U653 (N_653,In_0,In_348);
nor U654 (N_654,In_650,In_77);
and U655 (N_655,In_689,In_180);
or U656 (N_656,In_747,In_864);
nor U657 (N_657,In_16,In_790);
xnor U658 (N_658,In_836,In_305);
or U659 (N_659,In_724,In_563);
nand U660 (N_660,In_991,In_875);
nor U661 (N_661,In_250,In_405);
xor U662 (N_662,In_379,In_919);
and U663 (N_663,In_458,In_352);
and U664 (N_664,In_749,In_581);
or U665 (N_665,In_38,In_956);
nor U666 (N_666,In_822,In_818);
nor U667 (N_667,In_97,In_95);
nand U668 (N_668,In_449,In_595);
nor U669 (N_669,In_640,In_805);
and U670 (N_670,In_288,In_460);
nand U671 (N_671,In_917,In_271);
nor U672 (N_672,In_993,In_941);
xnor U673 (N_673,In_296,In_455);
nand U674 (N_674,In_615,In_93);
xor U675 (N_675,In_942,In_291);
nor U676 (N_676,In_763,In_504);
and U677 (N_677,In_384,In_42);
nor U678 (N_678,In_315,In_28);
or U679 (N_679,In_18,In_912);
nand U680 (N_680,In_48,In_78);
nor U681 (N_681,In_931,In_388);
nand U682 (N_682,In_281,In_101);
or U683 (N_683,In_503,In_665);
nand U684 (N_684,In_343,In_651);
nor U685 (N_685,In_960,In_959);
and U686 (N_686,In_314,In_353);
nor U687 (N_687,In_602,In_443);
nand U688 (N_688,In_875,In_778);
or U689 (N_689,In_26,In_563);
and U690 (N_690,In_999,In_901);
and U691 (N_691,In_155,In_786);
and U692 (N_692,In_943,In_831);
or U693 (N_693,In_983,In_603);
nor U694 (N_694,In_197,In_279);
xor U695 (N_695,In_874,In_383);
or U696 (N_696,In_641,In_239);
nor U697 (N_697,In_957,In_741);
xor U698 (N_698,In_845,In_785);
or U699 (N_699,In_418,In_895);
xor U700 (N_700,In_829,In_554);
or U701 (N_701,In_873,In_806);
and U702 (N_702,In_769,In_654);
xor U703 (N_703,In_700,In_839);
xnor U704 (N_704,In_267,In_433);
xor U705 (N_705,In_317,In_355);
nor U706 (N_706,In_535,In_628);
or U707 (N_707,In_512,In_569);
and U708 (N_708,In_752,In_805);
nand U709 (N_709,In_342,In_131);
nor U710 (N_710,In_300,In_140);
nor U711 (N_711,In_255,In_477);
or U712 (N_712,In_215,In_415);
nand U713 (N_713,In_703,In_834);
nand U714 (N_714,In_417,In_810);
nor U715 (N_715,In_927,In_41);
nor U716 (N_716,In_766,In_257);
or U717 (N_717,In_327,In_333);
nand U718 (N_718,In_684,In_682);
nand U719 (N_719,In_561,In_860);
nor U720 (N_720,In_585,In_861);
and U721 (N_721,In_485,In_559);
xor U722 (N_722,In_162,In_788);
and U723 (N_723,In_409,In_83);
and U724 (N_724,In_176,In_503);
nand U725 (N_725,In_457,In_999);
or U726 (N_726,In_461,In_19);
xor U727 (N_727,In_644,In_903);
nor U728 (N_728,In_812,In_132);
xnor U729 (N_729,In_488,In_622);
nand U730 (N_730,In_584,In_107);
xnor U731 (N_731,In_624,In_61);
nor U732 (N_732,In_909,In_772);
nand U733 (N_733,In_168,In_522);
xor U734 (N_734,In_973,In_486);
or U735 (N_735,In_421,In_706);
or U736 (N_736,In_744,In_484);
nor U737 (N_737,In_846,In_778);
or U738 (N_738,In_758,In_904);
xor U739 (N_739,In_427,In_940);
nand U740 (N_740,In_991,In_574);
nor U741 (N_741,In_268,In_167);
nor U742 (N_742,In_970,In_793);
or U743 (N_743,In_953,In_522);
nor U744 (N_744,In_702,In_550);
or U745 (N_745,In_608,In_517);
or U746 (N_746,In_404,In_575);
nand U747 (N_747,In_737,In_220);
nor U748 (N_748,In_607,In_643);
nor U749 (N_749,In_6,In_158);
nor U750 (N_750,In_451,In_526);
or U751 (N_751,In_423,In_801);
nor U752 (N_752,In_485,In_245);
or U753 (N_753,In_31,In_64);
nand U754 (N_754,In_412,In_608);
nand U755 (N_755,In_486,In_213);
nor U756 (N_756,In_785,In_842);
and U757 (N_757,In_240,In_180);
nand U758 (N_758,In_375,In_125);
nor U759 (N_759,In_659,In_511);
or U760 (N_760,In_300,In_389);
nor U761 (N_761,In_587,In_901);
or U762 (N_762,In_596,In_777);
xnor U763 (N_763,In_415,In_115);
and U764 (N_764,In_604,In_251);
nor U765 (N_765,In_728,In_637);
and U766 (N_766,In_148,In_872);
nand U767 (N_767,In_61,In_613);
and U768 (N_768,In_924,In_541);
xnor U769 (N_769,In_220,In_335);
and U770 (N_770,In_360,In_378);
xor U771 (N_771,In_674,In_323);
nand U772 (N_772,In_927,In_926);
xor U773 (N_773,In_420,In_943);
nand U774 (N_774,In_8,In_749);
nand U775 (N_775,In_846,In_828);
and U776 (N_776,In_113,In_553);
nor U777 (N_777,In_134,In_400);
or U778 (N_778,In_199,In_854);
nor U779 (N_779,In_807,In_394);
nand U780 (N_780,In_450,In_33);
nor U781 (N_781,In_204,In_680);
nor U782 (N_782,In_456,In_193);
xor U783 (N_783,In_385,In_386);
nand U784 (N_784,In_688,In_19);
xor U785 (N_785,In_807,In_314);
nand U786 (N_786,In_389,In_449);
nand U787 (N_787,In_116,In_752);
xor U788 (N_788,In_525,In_310);
nor U789 (N_789,In_401,In_699);
nor U790 (N_790,In_340,In_415);
nor U791 (N_791,In_971,In_211);
xor U792 (N_792,In_842,In_67);
and U793 (N_793,In_673,In_767);
nand U794 (N_794,In_356,In_182);
xor U795 (N_795,In_938,In_426);
nand U796 (N_796,In_681,In_198);
xnor U797 (N_797,In_489,In_169);
xnor U798 (N_798,In_821,In_191);
or U799 (N_799,In_887,In_101);
and U800 (N_800,In_825,In_459);
or U801 (N_801,In_182,In_247);
xor U802 (N_802,In_778,In_952);
xor U803 (N_803,In_913,In_342);
and U804 (N_804,In_839,In_104);
nand U805 (N_805,In_0,In_586);
nand U806 (N_806,In_434,In_452);
nand U807 (N_807,In_831,In_68);
or U808 (N_808,In_989,In_78);
nor U809 (N_809,In_362,In_226);
nand U810 (N_810,In_613,In_244);
and U811 (N_811,In_456,In_769);
xnor U812 (N_812,In_334,In_397);
and U813 (N_813,In_865,In_399);
and U814 (N_814,In_141,In_91);
or U815 (N_815,In_579,In_635);
nand U816 (N_816,In_608,In_301);
nor U817 (N_817,In_584,In_975);
xor U818 (N_818,In_907,In_679);
xnor U819 (N_819,In_126,In_515);
xor U820 (N_820,In_612,In_130);
nor U821 (N_821,In_963,In_66);
xnor U822 (N_822,In_113,In_811);
nor U823 (N_823,In_355,In_941);
xnor U824 (N_824,In_168,In_399);
or U825 (N_825,In_99,In_96);
xor U826 (N_826,In_803,In_134);
nand U827 (N_827,In_453,In_692);
and U828 (N_828,In_969,In_693);
and U829 (N_829,In_719,In_964);
or U830 (N_830,In_9,In_370);
and U831 (N_831,In_451,In_826);
or U832 (N_832,In_40,In_721);
nor U833 (N_833,In_858,In_922);
or U834 (N_834,In_473,In_658);
nor U835 (N_835,In_111,In_766);
and U836 (N_836,In_811,In_320);
and U837 (N_837,In_498,In_541);
or U838 (N_838,In_761,In_429);
nor U839 (N_839,In_790,In_615);
nor U840 (N_840,In_459,In_699);
or U841 (N_841,In_290,In_199);
and U842 (N_842,In_41,In_301);
and U843 (N_843,In_583,In_770);
or U844 (N_844,In_996,In_146);
or U845 (N_845,In_938,In_35);
nor U846 (N_846,In_96,In_171);
nand U847 (N_847,In_813,In_273);
or U848 (N_848,In_0,In_735);
and U849 (N_849,In_380,In_549);
or U850 (N_850,In_943,In_61);
or U851 (N_851,In_906,In_453);
or U852 (N_852,In_714,In_927);
nand U853 (N_853,In_551,In_633);
nand U854 (N_854,In_557,In_43);
or U855 (N_855,In_334,In_603);
xnor U856 (N_856,In_187,In_750);
xor U857 (N_857,In_952,In_328);
nand U858 (N_858,In_318,In_210);
and U859 (N_859,In_560,In_203);
or U860 (N_860,In_61,In_540);
nor U861 (N_861,In_779,In_943);
nor U862 (N_862,In_630,In_145);
nand U863 (N_863,In_267,In_986);
and U864 (N_864,In_514,In_9);
nor U865 (N_865,In_713,In_455);
nor U866 (N_866,In_622,In_537);
or U867 (N_867,In_582,In_863);
xnor U868 (N_868,In_766,In_700);
and U869 (N_869,In_564,In_662);
xnor U870 (N_870,In_166,In_423);
and U871 (N_871,In_714,In_113);
and U872 (N_872,In_226,In_266);
or U873 (N_873,In_813,In_581);
nor U874 (N_874,In_511,In_536);
nand U875 (N_875,In_758,In_520);
xor U876 (N_876,In_374,In_211);
xnor U877 (N_877,In_341,In_79);
nor U878 (N_878,In_724,In_597);
or U879 (N_879,In_825,In_281);
xnor U880 (N_880,In_18,In_65);
nand U881 (N_881,In_243,In_631);
or U882 (N_882,In_704,In_308);
and U883 (N_883,In_652,In_558);
nand U884 (N_884,In_171,In_612);
xor U885 (N_885,In_392,In_528);
and U886 (N_886,In_393,In_838);
or U887 (N_887,In_466,In_704);
nor U888 (N_888,In_162,In_30);
or U889 (N_889,In_497,In_308);
xnor U890 (N_890,In_779,In_260);
xnor U891 (N_891,In_711,In_368);
xor U892 (N_892,In_323,In_639);
or U893 (N_893,In_830,In_644);
nor U894 (N_894,In_828,In_16);
xnor U895 (N_895,In_204,In_414);
and U896 (N_896,In_85,In_685);
nand U897 (N_897,In_187,In_12);
nand U898 (N_898,In_968,In_609);
nand U899 (N_899,In_538,In_492);
nand U900 (N_900,In_691,In_541);
xor U901 (N_901,In_535,In_386);
nand U902 (N_902,In_749,In_99);
or U903 (N_903,In_164,In_954);
and U904 (N_904,In_98,In_222);
nor U905 (N_905,In_816,In_577);
xor U906 (N_906,In_270,In_106);
or U907 (N_907,In_663,In_386);
xor U908 (N_908,In_197,In_264);
and U909 (N_909,In_724,In_752);
nand U910 (N_910,In_977,In_803);
nor U911 (N_911,In_494,In_434);
and U912 (N_912,In_780,In_278);
nand U913 (N_913,In_840,In_34);
and U914 (N_914,In_289,In_637);
or U915 (N_915,In_902,In_759);
nand U916 (N_916,In_336,In_591);
or U917 (N_917,In_685,In_978);
xor U918 (N_918,In_951,In_580);
nand U919 (N_919,In_364,In_51);
and U920 (N_920,In_24,In_203);
nand U921 (N_921,In_881,In_662);
and U922 (N_922,In_123,In_43);
nand U923 (N_923,In_488,In_105);
or U924 (N_924,In_119,In_368);
and U925 (N_925,In_812,In_718);
nor U926 (N_926,In_486,In_494);
and U927 (N_927,In_631,In_132);
xnor U928 (N_928,In_262,In_965);
or U929 (N_929,In_835,In_481);
nor U930 (N_930,In_695,In_868);
xor U931 (N_931,In_607,In_622);
xnor U932 (N_932,In_853,In_927);
nor U933 (N_933,In_786,In_537);
xor U934 (N_934,In_245,In_999);
xnor U935 (N_935,In_762,In_598);
or U936 (N_936,In_627,In_434);
and U937 (N_937,In_186,In_833);
and U938 (N_938,In_131,In_404);
or U939 (N_939,In_229,In_788);
and U940 (N_940,In_738,In_873);
nor U941 (N_941,In_731,In_961);
and U942 (N_942,In_320,In_365);
nand U943 (N_943,In_39,In_855);
or U944 (N_944,In_795,In_193);
and U945 (N_945,In_539,In_59);
xnor U946 (N_946,In_975,In_74);
nand U947 (N_947,In_500,In_795);
and U948 (N_948,In_641,In_375);
nand U949 (N_949,In_268,In_7);
and U950 (N_950,In_56,In_169);
or U951 (N_951,In_15,In_479);
nor U952 (N_952,In_170,In_485);
nor U953 (N_953,In_388,In_357);
nor U954 (N_954,In_109,In_876);
nand U955 (N_955,In_489,In_607);
nand U956 (N_956,In_74,In_297);
or U957 (N_957,In_357,In_772);
nor U958 (N_958,In_412,In_984);
nor U959 (N_959,In_415,In_110);
nand U960 (N_960,In_341,In_991);
nand U961 (N_961,In_489,In_760);
nand U962 (N_962,In_625,In_775);
xor U963 (N_963,In_31,In_165);
or U964 (N_964,In_976,In_841);
nand U965 (N_965,In_45,In_975);
xnor U966 (N_966,In_811,In_553);
and U967 (N_967,In_599,In_70);
nand U968 (N_968,In_985,In_629);
xor U969 (N_969,In_399,In_514);
nor U970 (N_970,In_22,In_28);
and U971 (N_971,In_59,In_294);
xnor U972 (N_972,In_187,In_217);
or U973 (N_973,In_784,In_969);
and U974 (N_974,In_78,In_316);
nand U975 (N_975,In_296,In_705);
and U976 (N_976,In_987,In_58);
xnor U977 (N_977,In_88,In_291);
and U978 (N_978,In_127,In_642);
and U979 (N_979,In_215,In_532);
nand U980 (N_980,In_598,In_419);
nand U981 (N_981,In_359,In_129);
nand U982 (N_982,In_947,In_184);
xor U983 (N_983,In_444,In_299);
and U984 (N_984,In_306,In_889);
nor U985 (N_985,In_972,In_471);
nor U986 (N_986,In_977,In_766);
xor U987 (N_987,In_240,In_253);
nand U988 (N_988,In_186,In_933);
xor U989 (N_989,In_847,In_954);
nand U990 (N_990,In_837,In_925);
nor U991 (N_991,In_623,In_495);
xnor U992 (N_992,In_604,In_617);
nand U993 (N_993,In_998,In_106);
or U994 (N_994,In_939,In_984);
or U995 (N_995,In_160,In_888);
or U996 (N_996,In_917,In_865);
nor U997 (N_997,In_267,In_509);
nor U998 (N_998,In_854,In_544);
nand U999 (N_999,In_974,In_832);
nand U1000 (N_1000,N_526,N_527);
and U1001 (N_1001,N_814,N_324);
nor U1002 (N_1002,N_406,N_907);
or U1003 (N_1003,N_105,N_33);
or U1004 (N_1004,N_973,N_504);
nor U1005 (N_1005,N_201,N_939);
xor U1006 (N_1006,N_878,N_340);
nand U1007 (N_1007,N_350,N_432);
nand U1008 (N_1008,N_557,N_582);
nor U1009 (N_1009,N_363,N_47);
nor U1010 (N_1010,N_334,N_698);
nor U1011 (N_1011,N_172,N_49);
or U1012 (N_1012,N_393,N_822);
or U1013 (N_1013,N_162,N_695);
xor U1014 (N_1014,N_665,N_141);
or U1015 (N_1015,N_946,N_866);
and U1016 (N_1016,N_271,N_355);
and U1017 (N_1017,N_349,N_658);
or U1018 (N_1018,N_98,N_899);
nand U1019 (N_1019,N_78,N_837);
and U1020 (N_1020,N_293,N_482);
xnor U1021 (N_1021,N_303,N_756);
or U1022 (N_1022,N_358,N_203);
nand U1023 (N_1023,N_921,N_360);
nor U1024 (N_1024,N_93,N_429);
xor U1025 (N_1025,N_241,N_515);
xnor U1026 (N_1026,N_976,N_811);
nor U1027 (N_1027,N_932,N_23);
and U1028 (N_1028,N_993,N_356);
and U1029 (N_1029,N_65,N_151);
nand U1030 (N_1030,N_501,N_160);
or U1031 (N_1031,N_436,N_736);
or U1032 (N_1032,N_31,N_353);
nor U1033 (N_1033,N_717,N_280);
and U1034 (N_1034,N_536,N_73);
or U1035 (N_1035,N_640,N_895);
nand U1036 (N_1036,N_458,N_194);
or U1037 (N_1037,N_192,N_569);
nor U1038 (N_1038,N_588,N_125);
nor U1039 (N_1039,N_290,N_461);
or U1040 (N_1040,N_738,N_239);
nand U1041 (N_1041,N_322,N_116);
nor U1042 (N_1042,N_108,N_253);
xnor U1043 (N_1043,N_408,N_633);
and U1044 (N_1044,N_900,N_602);
and U1045 (N_1045,N_776,N_221);
nor U1046 (N_1046,N_10,N_88);
nor U1047 (N_1047,N_265,N_890);
nor U1048 (N_1048,N_594,N_209);
and U1049 (N_1049,N_53,N_860);
or U1050 (N_1050,N_3,N_785);
xnor U1051 (N_1051,N_445,N_631);
nand U1052 (N_1052,N_54,N_904);
nand U1053 (N_1053,N_998,N_875);
nand U1054 (N_1054,N_145,N_273);
nand U1055 (N_1055,N_779,N_962);
and U1056 (N_1056,N_924,N_628);
and U1057 (N_1057,N_743,N_252);
nor U1058 (N_1058,N_331,N_202);
nor U1059 (N_1059,N_827,N_975);
xnor U1060 (N_1060,N_958,N_772);
xor U1061 (N_1061,N_180,N_989);
xnor U1062 (N_1062,N_212,N_763);
or U1063 (N_1063,N_609,N_138);
nand U1064 (N_1064,N_573,N_128);
nor U1065 (N_1065,N_777,N_189);
or U1066 (N_1066,N_555,N_300);
nand U1067 (N_1067,N_951,N_641);
and U1068 (N_1068,N_456,N_991);
and U1069 (N_1069,N_694,N_560);
and U1070 (N_1070,N_457,N_635);
and U1071 (N_1071,N_943,N_682);
xnor U1072 (N_1072,N_846,N_918);
and U1073 (N_1073,N_441,N_134);
nand U1074 (N_1074,N_732,N_700);
or U1075 (N_1075,N_184,N_509);
or U1076 (N_1076,N_646,N_643);
or U1077 (N_1077,N_37,N_264);
xnor U1078 (N_1078,N_351,N_66);
nand U1079 (N_1079,N_314,N_323);
xor U1080 (N_1080,N_873,N_531);
nor U1081 (N_1081,N_181,N_967);
xor U1082 (N_1082,N_905,N_693);
nand U1083 (N_1083,N_940,N_106);
nand U1084 (N_1084,N_86,N_140);
and U1085 (N_1085,N_269,N_268);
xnor U1086 (N_1086,N_887,N_439);
nand U1087 (N_1087,N_608,N_295);
or U1088 (N_1088,N_90,N_662);
xor U1089 (N_1089,N_489,N_699);
nand U1090 (N_1090,N_27,N_716);
or U1091 (N_1091,N_882,N_492);
nor U1092 (N_1092,N_744,N_908);
nand U1093 (N_1093,N_460,N_751);
xor U1094 (N_1094,N_177,N_922);
nand U1095 (N_1095,N_583,N_22);
or U1096 (N_1096,N_824,N_650);
or U1097 (N_1097,N_412,N_316);
and U1098 (N_1098,N_839,N_183);
or U1099 (N_1099,N_20,N_934);
nor U1100 (N_1100,N_791,N_136);
nor U1101 (N_1101,N_486,N_844);
nand U1102 (N_1102,N_339,N_519);
nor U1103 (N_1103,N_668,N_186);
nand U1104 (N_1104,N_85,N_567);
nand U1105 (N_1105,N_233,N_413);
or U1106 (N_1106,N_649,N_352);
xnor U1107 (N_1107,N_75,N_701);
nor U1108 (N_1108,N_220,N_817);
nor U1109 (N_1109,N_16,N_69);
or U1110 (N_1110,N_821,N_771);
nor U1111 (N_1111,N_227,N_472);
or U1112 (N_1112,N_605,N_284);
and U1113 (N_1113,N_45,N_659);
or U1114 (N_1114,N_135,N_288);
and U1115 (N_1115,N_596,N_72);
xor U1116 (N_1116,N_56,N_29);
or U1117 (N_1117,N_276,N_706);
nor U1118 (N_1118,N_679,N_48);
nand U1119 (N_1119,N_789,N_784);
nand U1120 (N_1120,N_988,N_571);
nor U1121 (N_1121,N_496,N_217);
nand U1122 (N_1122,N_347,N_868);
or U1123 (N_1123,N_291,N_512);
nor U1124 (N_1124,N_144,N_684);
nor U1125 (N_1125,N_651,N_267);
nor U1126 (N_1126,N_657,N_911);
and U1127 (N_1127,N_714,N_286);
xnor U1128 (N_1128,N_21,N_500);
xor U1129 (N_1129,N_188,N_617);
nor U1130 (N_1130,N_179,N_497);
and U1131 (N_1131,N_977,N_213);
nor U1132 (N_1132,N_343,N_366);
nand U1133 (N_1133,N_468,N_38);
nor U1134 (N_1134,N_781,N_398);
or U1135 (N_1135,N_954,N_678);
nor U1136 (N_1136,N_431,N_402);
xnor U1137 (N_1137,N_113,N_426);
nor U1138 (N_1138,N_82,N_257);
xor U1139 (N_1139,N_287,N_546);
nor U1140 (N_1140,N_238,N_455);
xnor U1141 (N_1141,N_169,N_676);
nor U1142 (N_1142,N_454,N_537);
and U1143 (N_1143,N_542,N_522);
or U1144 (N_1144,N_99,N_381);
and U1145 (N_1145,N_463,N_312);
nand U1146 (N_1146,N_948,N_775);
xnor U1147 (N_1147,N_764,N_936);
and U1148 (N_1148,N_139,N_773);
or U1149 (N_1149,N_346,N_564);
nand U1150 (N_1150,N_880,N_229);
xor U1151 (N_1151,N_618,N_262);
or U1152 (N_1152,N_100,N_972);
and U1153 (N_1153,N_103,N_261);
and U1154 (N_1154,N_929,N_577);
xnor U1155 (N_1155,N_226,N_80);
or U1156 (N_1156,N_995,N_417);
xnor U1157 (N_1157,N_845,N_986);
nor U1158 (N_1158,N_345,N_656);
xnor U1159 (N_1159,N_94,N_167);
nor U1160 (N_1160,N_187,N_697);
xnor U1161 (N_1161,N_329,N_753);
nand U1162 (N_1162,N_881,N_807);
xnor U1163 (N_1163,N_163,N_947);
nand U1164 (N_1164,N_626,N_175);
xor U1165 (N_1165,N_11,N_132);
nand U1166 (N_1166,N_67,N_421);
nor U1167 (N_1167,N_600,N_142);
xnor U1168 (N_1168,N_690,N_199);
or U1169 (N_1169,N_525,N_185);
nand U1170 (N_1170,N_853,N_884);
nand U1171 (N_1171,N_996,N_502);
nor U1172 (N_1172,N_57,N_237);
or U1173 (N_1173,N_969,N_704);
nand U1174 (N_1174,N_126,N_475);
nor U1175 (N_1175,N_828,N_892);
nand U1176 (N_1176,N_916,N_244);
nor U1177 (N_1177,N_545,N_733);
nor U1178 (N_1178,N_757,N_487);
or U1179 (N_1179,N_231,N_89);
xor U1180 (N_1180,N_466,N_133);
nand U1181 (N_1181,N_832,N_485);
and U1182 (N_1182,N_556,N_34);
nand U1183 (N_1183,N_13,N_745);
nand U1184 (N_1184,N_77,N_585);
or U1185 (N_1185,N_4,N_159);
nor U1186 (N_1186,N_154,N_374);
nand U1187 (N_1187,N_917,N_114);
or U1188 (N_1188,N_834,N_430);
and U1189 (N_1189,N_120,N_869);
and U1190 (N_1190,N_831,N_801);
nand U1191 (N_1191,N_153,N_83);
or U1192 (N_1192,N_514,N_559);
xor U1193 (N_1193,N_388,N_891);
xor U1194 (N_1194,N_170,N_30);
or U1195 (N_1195,N_857,N_122);
and U1196 (N_1196,N_318,N_95);
nor U1197 (N_1197,N_914,N_576);
and U1198 (N_1198,N_942,N_893);
xnor U1199 (N_1199,N_214,N_127);
nand U1200 (N_1200,N_117,N_754);
nand U1201 (N_1201,N_40,N_630);
nor U1202 (N_1202,N_768,N_964);
and U1203 (N_1203,N_840,N_790);
xnor U1204 (N_1204,N_750,N_561);
xor U1205 (N_1205,N_637,N_889);
nor U1206 (N_1206,N_176,N_401);
or U1207 (N_1207,N_107,N_632);
or U1208 (N_1208,N_713,N_647);
or U1209 (N_1209,N_808,N_440);
and U1210 (N_1210,N_562,N_61);
and U1211 (N_1211,N_357,N_477);
nor U1212 (N_1212,N_666,N_616);
xor U1213 (N_1213,N_341,N_302);
or U1214 (N_1214,N_849,N_685);
nor U1215 (N_1215,N_191,N_143);
and U1216 (N_1216,N_830,N_944);
nor U1217 (N_1217,N_933,N_671);
nand U1218 (N_1218,N_478,N_660);
xnor U1219 (N_1219,N_782,N_405);
or U1220 (N_1220,N_173,N_242);
or U1221 (N_1221,N_369,N_119);
nand U1222 (N_1222,N_850,N_858);
nand U1223 (N_1223,N_864,N_935);
nor U1224 (N_1224,N_292,N_499);
or U1225 (N_1225,N_696,N_879);
or U1226 (N_1226,N_980,N_816);
nor U1227 (N_1227,N_952,N_9);
nor U1228 (N_1228,N_473,N_957);
nor U1229 (N_1229,N_810,N_897);
xor U1230 (N_1230,N_488,N_256);
or U1231 (N_1231,N_688,N_418);
or U1232 (N_1232,N_606,N_877);
nand U1233 (N_1233,N_419,N_551);
or U1234 (N_1234,N_307,N_298);
and U1235 (N_1235,N_396,N_788);
nand U1236 (N_1236,N_380,N_338);
and U1237 (N_1237,N_901,N_270);
and U1238 (N_1238,N_155,N_792);
xor U1239 (N_1239,N_841,N_87);
xor U1240 (N_1240,N_411,N_394);
xor U1241 (N_1241,N_912,N_211);
or U1242 (N_1242,N_580,N_547);
nand U1243 (N_1243,N_661,N_336);
or U1244 (N_1244,N_722,N_758);
nand U1245 (N_1245,N_655,N_513);
or U1246 (N_1246,N_102,N_390);
and U1247 (N_1247,N_335,N_855);
nand U1248 (N_1248,N_386,N_495);
xor U1249 (N_1249,N_702,N_131);
nand U1250 (N_1250,N_615,N_886);
and U1251 (N_1251,N_503,N_210);
or U1252 (N_1252,N_578,N_910);
and U1253 (N_1253,N_802,N_888);
or U1254 (N_1254,N_813,N_624);
nand U1255 (N_1255,N_692,N_876);
nor U1256 (N_1256,N_620,N_568);
or U1257 (N_1257,N_740,N_613);
and U1258 (N_1258,N_505,N_433);
or U1259 (N_1259,N_634,N_234);
xor U1260 (N_1260,N_370,N_611);
and U1261 (N_1261,N_196,N_344);
and U1262 (N_1262,N_803,N_109);
nand U1263 (N_1263,N_373,N_994);
nand U1264 (N_1264,N_843,N_248);
nand U1265 (N_1265,N_446,N_423);
and U1266 (N_1266,N_91,N_365);
and U1267 (N_1267,N_317,N_539);
and U1268 (N_1268,N_493,N_883);
nor U1269 (N_1269,N_200,N_552);
nand U1270 (N_1270,N_19,N_277);
nand U1271 (N_1271,N_62,N_726);
nand U1272 (N_1272,N_854,N_484);
xnor U1273 (N_1273,N_79,N_289);
nand U1274 (N_1274,N_36,N_558);
or U1275 (N_1275,N_310,N_171);
nand U1276 (N_1276,N_621,N_965);
nor U1277 (N_1277,N_639,N_377);
nor U1278 (N_1278,N_950,N_581);
nor U1279 (N_1279,N_451,N_689);
and U1280 (N_1280,N_819,N_586);
and U1281 (N_1281,N_861,N_115);
or U1282 (N_1282,N_607,N_833);
and U1283 (N_1283,N_326,N_245);
or U1284 (N_1284,N_464,N_297);
and U1285 (N_1285,N_315,N_938);
xnor U1286 (N_1286,N_206,N_870);
xnor U1287 (N_1287,N_541,N_760);
xnor U1288 (N_1288,N_70,N_663);
nand U1289 (N_1289,N_50,N_687);
nor U1290 (N_1290,N_710,N_24);
or U1291 (N_1291,N_762,N_707);
nand U1292 (N_1292,N_332,N_735);
nand U1293 (N_1293,N_305,N_376);
nand U1294 (N_1294,N_325,N_770);
or U1295 (N_1295,N_26,N_992);
nor U1296 (N_1296,N_761,N_966);
or U1297 (N_1297,N_285,N_711);
or U1298 (N_1298,N_529,N_595);
or U1299 (N_1299,N_592,N_272);
nand U1300 (N_1300,N_926,N_767);
nor U1301 (N_1301,N_250,N_806);
xor U1302 (N_1302,N_58,N_584);
and U1303 (N_1303,N_224,N_118);
nor U1304 (N_1304,N_982,N_450);
nand U1305 (N_1305,N_727,N_246);
xnor U1306 (N_1306,N_235,N_553);
nand U1307 (N_1307,N_826,N_511);
or U1308 (N_1308,N_368,N_533);
nand U1309 (N_1309,N_166,N_674);
xnor U1310 (N_1310,N_379,N_614);
or U1311 (N_1311,N_375,N_793);
and U1312 (N_1312,N_798,N_636);
and U1313 (N_1313,N_794,N_18);
nor U1314 (N_1314,N_404,N_981);
and U1315 (N_1315,N_540,N_372);
nand U1316 (N_1316,N_797,N_931);
nor U1317 (N_1317,N_730,N_769);
and U1318 (N_1318,N_232,N_104);
and U1319 (N_1319,N_84,N_279);
and U1320 (N_1320,N_945,N_572);
xnor U1321 (N_1321,N_111,N_480);
or U1322 (N_1322,N_178,N_601);
or U1323 (N_1323,N_847,N_101);
or U1324 (N_1324,N_920,N_60);
nand U1325 (N_1325,N_452,N_364);
and U1326 (N_1326,N_563,N_648);
nand U1327 (N_1327,N_25,N_174);
or U1328 (N_1328,N_459,N_925);
nor U1329 (N_1329,N_491,N_407);
nor U1330 (N_1330,N_76,N_215);
xor U1331 (N_1331,N_448,N_680);
xor U1332 (N_1332,N_971,N_731);
nand U1333 (N_1333,N_937,N_720);
and U1334 (N_1334,N_543,N_240);
nor U1335 (N_1335,N_677,N_409);
or U1336 (N_1336,N_725,N_422);
and U1337 (N_1337,N_208,N_321);
or U1338 (N_1338,N_534,N_746);
xnor U1339 (N_1339,N_742,N_361);
nand U1340 (N_1340,N_851,N_623);
xnor U1341 (N_1341,N_471,N_774);
nor U1342 (N_1342,N_523,N_367);
nand U1343 (N_1343,N_425,N_110);
xor U1344 (N_1344,N_909,N_255);
nor U1345 (N_1345,N_301,N_752);
nand U1346 (N_1346,N_81,N_427);
or U1347 (N_1347,N_2,N_462);
nor U1348 (N_1348,N_283,N_236);
xnor U1349 (N_1349,N_818,N_566);
and U1350 (N_1350,N_223,N_453);
nor U1351 (N_1351,N_872,N_734);
or U1352 (N_1352,N_469,N_867);
or U1353 (N_1353,N_391,N_309);
xnor U1354 (N_1354,N_7,N_260);
nand U1355 (N_1355,N_902,N_664);
or U1356 (N_1356,N_549,N_741);
or U1357 (N_1357,N_724,N_805);
nor U1358 (N_1358,N_795,N_579);
or U1359 (N_1359,N_359,N_517);
or U1360 (N_1360,N_149,N_984);
nand U1361 (N_1361,N_955,N_979);
and U1362 (N_1362,N_796,N_719);
nor U1363 (N_1363,N_447,N_894);
nor U1364 (N_1364,N_63,N_230);
or U1365 (N_1365,N_997,N_765);
or U1366 (N_1366,N_197,N_544);
or U1367 (N_1367,N_251,N_382);
and U1368 (N_1368,N_550,N_348);
or U1369 (N_1369,N_28,N_778);
or U1370 (N_1370,N_823,N_296);
xor U1371 (N_1371,N_333,N_403);
xnor U1372 (N_1372,N_434,N_538);
nand U1373 (N_1373,N_465,N_928);
xnor U1374 (N_1374,N_903,N_653);
xor U1375 (N_1375,N_723,N_121);
or U1376 (N_1376,N_686,N_780);
xor U1377 (N_1377,N_627,N_195);
nand U1378 (N_1378,N_198,N_168);
or U1379 (N_1379,N_718,N_494);
or U1380 (N_1380,N_51,N_825);
nor U1381 (N_1381,N_598,N_378);
nand U1382 (N_1382,N_961,N_281);
xnor U1383 (N_1383,N_507,N_629);
xor U1384 (N_1384,N_354,N_739);
nand U1385 (N_1385,N_518,N_150);
nor U1386 (N_1386,N_304,N_275);
and U1387 (N_1387,N_809,N_205);
or U1388 (N_1388,N_15,N_165);
or U1389 (N_1389,N_812,N_371);
nor U1390 (N_1390,N_673,N_152);
nor U1391 (N_1391,N_599,N_216);
and U1392 (N_1392,N_521,N_330);
nand U1393 (N_1393,N_68,N_766);
nor U1394 (N_1394,N_278,N_532);
nor U1395 (N_1395,N_565,N_164);
or U1396 (N_1396,N_476,N_604);
nand U1397 (N_1397,N_247,N_474);
or U1398 (N_1398,N_428,N_863);
nor U1399 (N_1399,N_587,N_672);
xor U1400 (N_1400,N_397,N_35);
xnor U1401 (N_1401,N_342,N_968);
nor U1402 (N_1402,N_148,N_498);
nand U1403 (N_1403,N_258,N_470);
xor U1404 (N_1404,N_786,N_392);
nand U1405 (N_1405,N_667,N_927);
and U1406 (N_1406,N_449,N_414);
xnor U1407 (N_1407,N_747,N_259);
xnor U1408 (N_1408,N_591,N_898);
nand U1409 (N_1409,N_835,N_437);
nor U1410 (N_1410,N_820,N_842);
xor U1411 (N_1411,N_1,N_737);
and U1412 (N_1412,N_856,N_622);
nand U1413 (N_1413,N_983,N_956);
xnor U1414 (N_1414,N_158,N_263);
nor U1415 (N_1415,N_570,N_438);
or U1416 (N_1416,N_970,N_865);
nor U1417 (N_1417,N_852,N_593);
nor U1418 (N_1418,N_416,N_721);
and U1419 (N_1419,N_590,N_311);
xnor U1420 (N_1420,N_222,N_74);
or U1421 (N_1421,N_654,N_64);
nand U1422 (N_1422,N_193,N_467);
nor U1423 (N_1423,N_389,N_574);
or U1424 (N_1424,N_32,N_508);
nand U1425 (N_1425,N_182,N_642);
and U1426 (N_1426,N_915,N_479);
nand U1427 (N_1427,N_97,N_400);
and U1428 (N_1428,N_528,N_759);
nor U1429 (N_1429,N_729,N_638);
nor U1430 (N_1430,N_225,N_249);
or U1431 (N_1431,N_218,N_254);
nor U1432 (N_1432,N_669,N_804);
nor U1433 (N_1433,N_683,N_39);
and U1434 (N_1434,N_597,N_589);
nand U1435 (N_1435,N_274,N_874);
and U1436 (N_1436,N_815,N_749);
and U1437 (N_1437,N_974,N_319);
nor U1438 (N_1438,N_55,N_999);
nand U1439 (N_1439,N_435,N_306);
xnor U1440 (N_1440,N_112,N_395);
nand U1441 (N_1441,N_930,N_207);
nor U1442 (N_1442,N_399,N_712);
nand U1443 (N_1443,N_941,N_219);
xnor U1444 (N_1444,N_548,N_266);
xnor U1445 (N_1445,N_510,N_953);
nor U1446 (N_1446,N_337,N_985);
or U1447 (N_1447,N_92,N_294);
xor U1448 (N_1448,N_123,N_146);
nor U1449 (N_1449,N_520,N_137);
nor U1450 (N_1450,N_282,N_243);
xor U1451 (N_1451,N_709,N_645);
nand U1452 (N_1452,N_885,N_385);
xor U1453 (N_1453,N_490,N_836);
xor U1454 (N_1454,N_859,N_524);
and U1455 (N_1455,N_862,N_681);
xnor U1456 (N_1456,N_299,N_228);
and U1457 (N_1457,N_147,N_44);
and U1458 (N_1458,N_670,N_161);
or U1459 (N_1459,N_619,N_506);
and U1460 (N_1460,N_575,N_0);
nor U1461 (N_1461,N_46,N_43);
xor U1462 (N_1462,N_424,N_799);
and U1463 (N_1463,N_313,N_481);
nor U1464 (N_1464,N_124,N_913);
and U1465 (N_1465,N_6,N_8);
nand U1466 (N_1466,N_415,N_443);
or U1467 (N_1467,N_554,N_848);
and U1468 (N_1468,N_204,N_17);
nor U1469 (N_1469,N_444,N_990);
nor U1470 (N_1470,N_5,N_320);
or U1471 (N_1471,N_59,N_328);
and U1472 (N_1472,N_705,N_71);
xor U1473 (N_1473,N_715,N_978);
nor U1474 (N_1474,N_420,N_703);
xor U1475 (N_1475,N_516,N_652);
and U1476 (N_1476,N_963,N_362);
xor U1477 (N_1477,N_42,N_327);
and U1478 (N_1478,N_41,N_829);
and U1479 (N_1479,N_383,N_535);
nor U1480 (N_1480,N_919,N_800);
nor U1481 (N_1481,N_783,N_384);
and U1482 (N_1482,N_308,N_675);
nor U1483 (N_1483,N_387,N_987);
nor U1484 (N_1484,N_923,N_442);
or U1485 (N_1485,N_96,N_483);
or U1486 (N_1486,N_755,N_906);
and U1487 (N_1487,N_130,N_871);
nand U1488 (N_1488,N_612,N_129);
nand U1489 (N_1489,N_748,N_12);
nor U1490 (N_1490,N_959,N_838);
or U1491 (N_1491,N_787,N_603);
xor U1492 (N_1492,N_728,N_52);
and U1493 (N_1493,N_14,N_625);
or U1494 (N_1494,N_949,N_691);
nor U1495 (N_1495,N_610,N_708);
nand U1496 (N_1496,N_156,N_530);
nand U1497 (N_1497,N_896,N_644);
or U1498 (N_1498,N_410,N_960);
and U1499 (N_1499,N_190,N_157);
xor U1500 (N_1500,N_891,N_39);
or U1501 (N_1501,N_867,N_543);
and U1502 (N_1502,N_908,N_980);
nand U1503 (N_1503,N_307,N_617);
nor U1504 (N_1504,N_297,N_184);
nand U1505 (N_1505,N_451,N_641);
nor U1506 (N_1506,N_380,N_476);
nand U1507 (N_1507,N_149,N_645);
xnor U1508 (N_1508,N_438,N_33);
nand U1509 (N_1509,N_542,N_734);
nor U1510 (N_1510,N_469,N_490);
nor U1511 (N_1511,N_41,N_359);
nor U1512 (N_1512,N_514,N_82);
nand U1513 (N_1513,N_788,N_466);
nand U1514 (N_1514,N_68,N_797);
nor U1515 (N_1515,N_891,N_136);
and U1516 (N_1516,N_995,N_117);
xnor U1517 (N_1517,N_769,N_867);
nand U1518 (N_1518,N_764,N_381);
and U1519 (N_1519,N_841,N_141);
nor U1520 (N_1520,N_350,N_493);
and U1521 (N_1521,N_576,N_743);
nand U1522 (N_1522,N_92,N_752);
or U1523 (N_1523,N_83,N_143);
nor U1524 (N_1524,N_804,N_994);
or U1525 (N_1525,N_848,N_394);
nand U1526 (N_1526,N_641,N_733);
and U1527 (N_1527,N_751,N_75);
nand U1528 (N_1528,N_776,N_361);
and U1529 (N_1529,N_420,N_812);
or U1530 (N_1530,N_299,N_974);
nor U1531 (N_1531,N_430,N_245);
or U1532 (N_1532,N_249,N_419);
nor U1533 (N_1533,N_284,N_863);
nor U1534 (N_1534,N_260,N_457);
nor U1535 (N_1535,N_514,N_524);
or U1536 (N_1536,N_513,N_924);
and U1537 (N_1537,N_302,N_956);
nand U1538 (N_1538,N_97,N_325);
xnor U1539 (N_1539,N_375,N_962);
xor U1540 (N_1540,N_553,N_236);
xnor U1541 (N_1541,N_1,N_346);
and U1542 (N_1542,N_624,N_795);
nand U1543 (N_1543,N_818,N_454);
nand U1544 (N_1544,N_254,N_322);
nand U1545 (N_1545,N_873,N_647);
nor U1546 (N_1546,N_745,N_153);
and U1547 (N_1547,N_394,N_966);
xor U1548 (N_1548,N_955,N_950);
xor U1549 (N_1549,N_808,N_386);
nand U1550 (N_1550,N_458,N_473);
nor U1551 (N_1551,N_631,N_124);
nand U1552 (N_1552,N_217,N_275);
or U1553 (N_1553,N_332,N_846);
nand U1554 (N_1554,N_178,N_467);
nand U1555 (N_1555,N_631,N_619);
or U1556 (N_1556,N_111,N_626);
nor U1557 (N_1557,N_866,N_87);
xor U1558 (N_1558,N_79,N_165);
nor U1559 (N_1559,N_281,N_938);
or U1560 (N_1560,N_684,N_298);
nand U1561 (N_1561,N_348,N_575);
nor U1562 (N_1562,N_338,N_896);
or U1563 (N_1563,N_335,N_851);
xnor U1564 (N_1564,N_811,N_773);
or U1565 (N_1565,N_201,N_570);
or U1566 (N_1566,N_710,N_190);
nand U1567 (N_1567,N_154,N_234);
nor U1568 (N_1568,N_113,N_173);
or U1569 (N_1569,N_894,N_707);
xnor U1570 (N_1570,N_732,N_811);
and U1571 (N_1571,N_293,N_201);
xnor U1572 (N_1572,N_881,N_711);
and U1573 (N_1573,N_386,N_957);
nand U1574 (N_1574,N_67,N_678);
nor U1575 (N_1575,N_983,N_230);
nand U1576 (N_1576,N_191,N_583);
nand U1577 (N_1577,N_773,N_763);
xor U1578 (N_1578,N_367,N_305);
nand U1579 (N_1579,N_459,N_621);
nand U1580 (N_1580,N_136,N_811);
nand U1581 (N_1581,N_922,N_930);
nand U1582 (N_1582,N_871,N_415);
xnor U1583 (N_1583,N_840,N_94);
xor U1584 (N_1584,N_158,N_865);
nor U1585 (N_1585,N_567,N_952);
nor U1586 (N_1586,N_765,N_249);
nor U1587 (N_1587,N_770,N_379);
nor U1588 (N_1588,N_954,N_788);
nor U1589 (N_1589,N_553,N_801);
and U1590 (N_1590,N_999,N_519);
nor U1591 (N_1591,N_980,N_496);
and U1592 (N_1592,N_487,N_674);
nand U1593 (N_1593,N_489,N_374);
nor U1594 (N_1594,N_168,N_788);
or U1595 (N_1595,N_374,N_25);
and U1596 (N_1596,N_959,N_17);
and U1597 (N_1597,N_463,N_147);
and U1598 (N_1598,N_781,N_568);
nand U1599 (N_1599,N_131,N_851);
nor U1600 (N_1600,N_871,N_756);
nor U1601 (N_1601,N_866,N_927);
nor U1602 (N_1602,N_495,N_787);
and U1603 (N_1603,N_266,N_193);
xor U1604 (N_1604,N_833,N_198);
xor U1605 (N_1605,N_89,N_234);
nor U1606 (N_1606,N_908,N_454);
xnor U1607 (N_1607,N_459,N_902);
or U1608 (N_1608,N_603,N_152);
nand U1609 (N_1609,N_589,N_221);
xor U1610 (N_1610,N_165,N_569);
and U1611 (N_1611,N_179,N_711);
and U1612 (N_1612,N_592,N_634);
or U1613 (N_1613,N_728,N_311);
and U1614 (N_1614,N_674,N_311);
xnor U1615 (N_1615,N_35,N_83);
nand U1616 (N_1616,N_945,N_732);
or U1617 (N_1617,N_793,N_526);
and U1618 (N_1618,N_553,N_743);
or U1619 (N_1619,N_159,N_188);
xnor U1620 (N_1620,N_93,N_407);
nor U1621 (N_1621,N_318,N_90);
or U1622 (N_1622,N_459,N_831);
xor U1623 (N_1623,N_944,N_574);
nor U1624 (N_1624,N_32,N_494);
and U1625 (N_1625,N_497,N_30);
and U1626 (N_1626,N_264,N_5);
nand U1627 (N_1627,N_900,N_685);
nand U1628 (N_1628,N_681,N_972);
nor U1629 (N_1629,N_607,N_807);
or U1630 (N_1630,N_116,N_74);
nand U1631 (N_1631,N_24,N_533);
and U1632 (N_1632,N_639,N_541);
or U1633 (N_1633,N_983,N_72);
xor U1634 (N_1634,N_937,N_282);
and U1635 (N_1635,N_147,N_439);
nor U1636 (N_1636,N_38,N_940);
and U1637 (N_1637,N_219,N_643);
nand U1638 (N_1638,N_420,N_987);
nor U1639 (N_1639,N_361,N_630);
nor U1640 (N_1640,N_826,N_47);
xnor U1641 (N_1641,N_556,N_53);
or U1642 (N_1642,N_15,N_317);
xnor U1643 (N_1643,N_577,N_154);
nand U1644 (N_1644,N_628,N_31);
or U1645 (N_1645,N_143,N_81);
nand U1646 (N_1646,N_844,N_415);
nand U1647 (N_1647,N_921,N_354);
nand U1648 (N_1648,N_896,N_141);
nor U1649 (N_1649,N_314,N_329);
xnor U1650 (N_1650,N_44,N_398);
nand U1651 (N_1651,N_473,N_596);
nand U1652 (N_1652,N_937,N_333);
nor U1653 (N_1653,N_55,N_433);
xnor U1654 (N_1654,N_145,N_287);
nor U1655 (N_1655,N_307,N_369);
nor U1656 (N_1656,N_332,N_788);
and U1657 (N_1657,N_514,N_504);
xnor U1658 (N_1658,N_420,N_82);
and U1659 (N_1659,N_861,N_998);
and U1660 (N_1660,N_908,N_898);
xnor U1661 (N_1661,N_807,N_400);
nor U1662 (N_1662,N_722,N_164);
and U1663 (N_1663,N_741,N_986);
and U1664 (N_1664,N_382,N_905);
and U1665 (N_1665,N_588,N_222);
or U1666 (N_1666,N_800,N_758);
nor U1667 (N_1667,N_113,N_436);
xnor U1668 (N_1668,N_245,N_449);
and U1669 (N_1669,N_598,N_958);
and U1670 (N_1670,N_219,N_112);
xor U1671 (N_1671,N_461,N_283);
nor U1672 (N_1672,N_892,N_442);
xnor U1673 (N_1673,N_704,N_185);
nor U1674 (N_1674,N_487,N_625);
or U1675 (N_1675,N_726,N_173);
nand U1676 (N_1676,N_180,N_236);
nand U1677 (N_1677,N_649,N_20);
nor U1678 (N_1678,N_167,N_89);
or U1679 (N_1679,N_226,N_64);
xnor U1680 (N_1680,N_807,N_216);
or U1681 (N_1681,N_368,N_56);
and U1682 (N_1682,N_445,N_257);
xnor U1683 (N_1683,N_602,N_494);
xor U1684 (N_1684,N_530,N_296);
nor U1685 (N_1685,N_851,N_774);
nor U1686 (N_1686,N_700,N_712);
nand U1687 (N_1687,N_326,N_404);
nor U1688 (N_1688,N_452,N_473);
or U1689 (N_1689,N_628,N_944);
nand U1690 (N_1690,N_121,N_394);
nor U1691 (N_1691,N_473,N_185);
nor U1692 (N_1692,N_491,N_848);
and U1693 (N_1693,N_319,N_814);
xor U1694 (N_1694,N_972,N_170);
nor U1695 (N_1695,N_2,N_675);
xor U1696 (N_1696,N_965,N_194);
and U1697 (N_1697,N_455,N_935);
nor U1698 (N_1698,N_536,N_550);
xor U1699 (N_1699,N_971,N_255);
xnor U1700 (N_1700,N_798,N_563);
nand U1701 (N_1701,N_724,N_599);
xor U1702 (N_1702,N_710,N_734);
nor U1703 (N_1703,N_968,N_138);
nor U1704 (N_1704,N_369,N_372);
and U1705 (N_1705,N_51,N_450);
nand U1706 (N_1706,N_856,N_935);
and U1707 (N_1707,N_23,N_178);
nor U1708 (N_1708,N_819,N_284);
nor U1709 (N_1709,N_931,N_749);
xnor U1710 (N_1710,N_109,N_100);
and U1711 (N_1711,N_381,N_104);
nor U1712 (N_1712,N_651,N_537);
xor U1713 (N_1713,N_34,N_152);
and U1714 (N_1714,N_673,N_510);
and U1715 (N_1715,N_854,N_602);
or U1716 (N_1716,N_757,N_732);
nor U1717 (N_1717,N_234,N_949);
and U1718 (N_1718,N_197,N_360);
or U1719 (N_1719,N_597,N_549);
nand U1720 (N_1720,N_220,N_777);
nor U1721 (N_1721,N_45,N_112);
or U1722 (N_1722,N_627,N_823);
or U1723 (N_1723,N_880,N_449);
or U1724 (N_1724,N_96,N_622);
nand U1725 (N_1725,N_459,N_115);
nor U1726 (N_1726,N_955,N_138);
nor U1727 (N_1727,N_791,N_908);
nand U1728 (N_1728,N_134,N_591);
or U1729 (N_1729,N_364,N_313);
nor U1730 (N_1730,N_671,N_759);
nand U1731 (N_1731,N_23,N_45);
nor U1732 (N_1732,N_835,N_937);
nor U1733 (N_1733,N_804,N_299);
and U1734 (N_1734,N_539,N_453);
and U1735 (N_1735,N_339,N_172);
and U1736 (N_1736,N_614,N_293);
nor U1737 (N_1737,N_175,N_903);
nor U1738 (N_1738,N_58,N_158);
and U1739 (N_1739,N_421,N_27);
nand U1740 (N_1740,N_97,N_694);
nor U1741 (N_1741,N_57,N_885);
nor U1742 (N_1742,N_578,N_966);
and U1743 (N_1743,N_636,N_933);
and U1744 (N_1744,N_546,N_88);
nand U1745 (N_1745,N_91,N_869);
nand U1746 (N_1746,N_197,N_699);
and U1747 (N_1747,N_926,N_952);
xnor U1748 (N_1748,N_795,N_915);
or U1749 (N_1749,N_753,N_121);
nand U1750 (N_1750,N_923,N_405);
and U1751 (N_1751,N_358,N_666);
nand U1752 (N_1752,N_725,N_614);
xnor U1753 (N_1753,N_218,N_156);
nor U1754 (N_1754,N_659,N_923);
or U1755 (N_1755,N_690,N_713);
xnor U1756 (N_1756,N_842,N_188);
nor U1757 (N_1757,N_676,N_357);
and U1758 (N_1758,N_140,N_277);
nand U1759 (N_1759,N_403,N_238);
nand U1760 (N_1760,N_966,N_76);
nor U1761 (N_1761,N_408,N_510);
or U1762 (N_1762,N_5,N_724);
and U1763 (N_1763,N_944,N_740);
nor U1764 (N_1764,N_273,N_695);
nand U1765 (N_1765,N_413,N_797);
xnor U1766 (N_1766,N_763,N_795);
and U1767 (N_1767,N_429,N_830);
nand U1768 (N_1768,N_196,N_655);
nand U1769 (N_1769,N_732,N_768);
or U1770 (N_1770,N_236,N_671);
nand U1771 (N_1771,N_626,N_814);
nand U1772 (N_1772,N_597,N_174);
nand U1773 (N_1773,N_169,N_957);
and U1774 (N_1774,N_551,N_379);
nand U1775 (N_1775,N_80,N_135);
and U1776 (N_1776,N_28,N_345);
xnor U1777 (N_1777,N_581,N_202);
xor U1778 (N_1778,N_679,N_322);
and U1779 (N_1779,N_772,N_427);
or U1780 (N_1780,N_819,N_661);
nor U1781 (N_1781,N_629,N_157);
and U1782 (N_1782,N_956,N_153);
nor U1783 (N_1783,N_244,N_248);
nor U1784 (N_1784,N_427,N_415);
or U1785 (N_1785,N_481,N_715);
nand U1786 (N_1786,N_365,N_876);
nor U1787 (N_1787,N_722,N_118);
nor U1788 (N_1788,N_501,N_585);
nor U1789 (N_1789,N_461,N_762);
or U1790 (N_1790,N_379,N_413);
or U1791 (N_1791,N_849,N_592);
and U1792 (N_1792,N_645,N_196);
and U1793 (N_1793,N_792,N_428);
and U1794 (N_1794,N_837,N_214);
nand U1795 (N_1795,N_370,N_423);
nand U1796 (N_1796,N_706,N_58);
and U1797 (N_1797,N_291,N_530);
and U1798 (N_1798,N_344,N_658);
or U1799 (N_1799,N_802,N_791);
xor U1800 (N_1800,N_569,N_986);
and U1801 (N_1801,N_663,N_354);
or U1802 (N_1802,N_906,N_332);
nor U1803 (N_1803,N_594,N_805);
and U1804 (N_1804,N_278,N_269);
or U1805 (N_1805,N_827,N_638);
nand U1806 (N_1806,N_46,N_141);
and U1807 (N_1807,N_270,N_25);
and U1808 (N_1808,N_69,N_64);
xnor U1809 (N_1809,N_204,N_99);
xor U1810 (N_1810,N_890,N_991);
and U1811 (N_1811,N_323,N_312);
or U1812 (N_1812,N_588,N_883);
nor U1813 (N_1813,N_735,N_365);
or U1814 (N_1814,N_257,N_745);
xnor U1815 (N_1815,N_193,N_959);
nor U1816 (N_1816,N_558,N_216);
nor U1817 (N_1817,N_133,N_991);
and U1818 (N_1818,N_825,N_365);
nor U1819 (N_1819,N_309,N_248);
nand U1820 (N_1820,N_280,N_608);
nand U1821 (N_1821,N_536,N_288);
xor U1822 (N_1822,N_919,N_261);
xor U1823 (N_1823,N_877,N_654);
and U1824 (N_1824,N_537,N_81);
nor U1825 (N_1825,N_3,N_568);
or U1826 (N_1826,N_552,N_942);
nor U1827 (N_1827,N_372,N_254);
nor U1828 (N_1828,N_744,N_585);
nor U1829 (N_1829,N_979,N_379);
nor U1830 (N_1830,N_691,N_302);
and U1831 (N_1831,N_536,N_389);
xor U1832 (N_1832,N_927,N_602);
nand U1833 (N_1833,N_924,N_153);
and U1834 (N_1834,N_477,N_744);
xnor U1835 (N_1835,N_366,N_894);
xnor U1836 (N_1836,N_598,N_404);
or U1837 (N_1837,N_547,N_841);
and U1838 (N_1838,N_519,N_229);
xnor U1839 (N_1839,N_59,N_997);
nor U1840 (N_1840,N_449,N_144);
or U1841 (N_1841,N_892,N_472);
xnor U1842 (N_1842,N_955,N_117);
and U1843 (N_1843,N_583,N_403);
or U1844 (N_1844,N_387,N_411);
nor U1845 (N_1845,N_535,N_953);
or U1846 (N_1846,N_988,N_981);
nor U1847 (N_1847,N_137,N_927);
and U1848 (N_1848,N_492,N_588);
or U1849 (N_1849,N_761,N_904);
xor U1850 (N_1850,N_320,N_323);
or U1851 (N_1851,N_21,N_419);
xnor U1852 (N_1852,N_171,N_678);
or U1853 (N_1853,N_238,N_669);
nand U1854 (N_1854,N_405,N_456);
nor U1855 (N_1855,N_491,N_437);
and U1856 (N_1856,N_613,N_504);
or U1857 (N_1857,N_999,N_425);
nor U1858 (N_1858,N_737,N_658);
and U1859 (N_1859,N_362,N_649);
nor U1860 (N_1860,N_263,N_968);
nand U1861 (N_1861,N_546,N_539);
and U1862 (N_1862,N_951,N_155);
nor U1863 (N_1863,N_659,N_182);
and U1864 (N_1864,N_314,N_702);
nor U1865 (N_1865,N_252,N_665);
nor U1866 (N_1866,N_395,N_509);
nand U1867 (N_1867,N_321,N_731);
xor U1868 (N_1868,N_959,N_556);
or U1869 (N_1869,N_255,N_534);
and U1870 (N_1870,N_637,N_560);
and U1871 (N_1871,N_158,N_768);
nand U1872 (N_1872,N_365,N_657);
or U1873 (N_1873,N_180,N_755);
nor U1874 (N_1874,N_990,N_146);
xor U1875 (N_1875,N_291,N_311);
or U1876 (N_1876,N_427,N_607);
and U1877 (N_1877,N_368,N_97);
nand U1878 (N_1878,N_703,N_548);
xor U1879 (N_1879,N_103,N_868);
xnor U1880 (N_1880,N_114,N_281);
and U1881 (N_1881,N_624,N_432);
nor U1882 (N_1882,N_143,N_357);
nor U1883 (N_1883,N_391,N_1);
nand U1884 (N_1884,N_813,N_332);
xnor U1885 (N_1885,N_531,N_399);
and U1886 (N_1886,N_297,N_201);
nor U1887 (N_1887,N_300,N_3);
or U1888 (N_1888,N_770,N_963);
xnor U1889 (N_1889,N_932,N_625);
nor U1890 (N_1890,N_240,N_772);
nand U1891 (N_1891,N_835,N_426);
xnor U1892 (N_1892,N_441,N_684);
nor U1893 (N_1893,N_936,N_896);
xnor U1894 (N_1894,N_956,N_303);
or U1895 (N_1895,N_449,N_364);
or U1896 (N_1896,N_151,N_142);
or U1897 (N_1897,N_839,N_622);
nor U1898 (N_1898,N_552,N_880);
and U1899 (N_1899,N_897,N_814);
xor U1900 (N_1900,N_386,N_320);
xor U1901 (N_1901,N_728,N_139);
xnor U1902 (N_1902,N_813,N_11);
xor U1903 (N_1903,N_61,N_850);
xor U1904 (N_1904,N_837,N_934);
and U1905 (N_1905,N_576,N_780);
or U1906 (N_1906,N_409,N_54);
nor U1907 (N_1907,N_809,N_745);
xnor U1908 (N_1908,N_359,N_880);
nand U1909 (N_1909,N_898,N_25);
xor U1910 (N_1910,N_411,N_422);
and U1911 (N_1911,N_301,N_556);
and U1912 (N_1912,N_626,N_902);
xor U1913 (N_1913,N_534,N_286);
nor U1914 (N_1914,N_342,N_911);
or U1915 (N_1915,N_388,N_15);
or U1916 (N_1916,N_992,N_658);
or U1917 (N_1917,N_14,N_407);
nand U1918 (N_1918,N_733,N_627);
nand U1919 (N_1919,N_415,N_515);
and U1920 (N_1920,N_453,N_521);
or U1921 (N_1921,N_406,N_846);
or U1922 (N_1922,N_873,N_944);
xnor U1923 (N_1923,N_729,N_213);
xnor U1924 (N_1924,N_449,N_999);
xnor U1925 (N_1925,N_293,N_51);
and U1926 (N_1926,N_226,N_152);
nand U1927 (N_1927,N_990,N_623);
or U1928 (N_1928,N_883,N_241);
nor U1929 (N_1929,N_134,N_115);
nor U1930 (N_1930,N_735,N_606);
and U1931 (N_1931,N_601,N_618);
xnor U1932 (N_1932,N_485,N_329);
and U1933 (N_1933,N_685,N_178);
nand U1934 (N_1934,N_210,N_570);
and U1935 (N_1935,N_50,N_77);
and U1936 (N_1936,N_467,N_533);
nor U1937 (N_1937,N_486,N_768);
nand U1938 (N_1938,N_835,N_923);
nand U1939 (N_1939,N_555,N_628);
or U1940 (N_1940,N_728,N_523);
nor U1941 (N_1941,N_573,N_862);
nor U1942 (N_1942,N_448,N_431);
xnor U1943 (N_1943,N_687,N_157);
nand U1944 (N_1944,N_581,N_855);
xor U1945 (N_1945,N_217,N_928);
nand U1946 (N_1946,N_779,N_411);
or U1947 (N_1947,N_208,N_85);
nor U1948 (N_1948,N_95,N_171);
nor U1949 (N_1949,N_233,N_5);
and U1950 (N_1950,N_597,N_350);
nor U1951 (N_1951,N_813,N_274);
nor U1952 (N_1952,N_771,N_585);
nand U1953 (N_1953,N_509,N_187);
nand U1954 (N_1954,N_761,N_312);
or U1955 (N_1955,N_89,N_226);
and U1956 (N_1956,N_339,N_164);
nor U1957 (N_1957,N_186,N_443);
or U1958 (N_1958,N_26,N_834);
nand U1959 (N_1959,N_408,N_194);
or U1960 (N_1960,N_457,N_187);
nor U1961 (N_1961,N_463,N_92);
or U1962 (N_1962,N_550,N_622);
nor U1963 (N_1963,N_741,N_819);
or U1964 (N_1964,N_301,N_46);
and U1965 (N_1965,N_750,N_641);
or U1966 (N_1966,N_408,N_562);
xnor U1967 (N_1967,N_15,N_865);
or U1968 (N_1968,N_782,N_584);
nor U1969 (N_1969,N_545,N_109);
nor U1970 (N_1970,N_386,N_549);
nor U1971 (N_1971,N_882,N_481);
nand U1972 (N_1972,N_441,N_888);
xor U1973 (N_1973,N_955,N_272);
xnor U1974 (N_1974,N_564,N_71);
and U1975 (N_1975,N_873,N_817);
xor U1976 (N_1976,N_485,N_188);
nand U1977 (N_1977,N_970,N_739);
nor U1978 (N_1978,N_882,N_377);
or U1979 (N_1979,N_847,N_925);
xor U1980 (N_1980,N_109,N_217);
or U1981 (N_1981,N_32,N_164);
or U1982 (N_1982,N_192,N_503);
and U1983 (N_1983,N_299,N_101);
or U1984 (N_1984,N_374,N_515);
and U1985 (N_1985,N_695,N_368);
or U1986 (N_1986,N_851,N_768);
or U1987 (N_1987,N_890,N_586);
and U1988 (N_1988,N_991,N_883);
and U1989 (N_1989,N_983,N_613);
nand U1990 (N_1990,N_219,N_72);
and U1991 (N_1991,N_832,N_719);
nor U1992 (N_1992,N_656,N_665);
or U1993 (N_1993,N_427,N_467);
nor U1994 (N_1994,N_508,N_168);
or U1995 (N_1995,N_40,N_203);
xor U1996 (N_1996,N_184,N_660);
or U1997 (N_1997,N_361,N_469);
or U1998 (N_1998,N_238,N_34);
or U1999 (N_1999,N_103,N_196);
xnor U2000 (N_2000,N_1738,N_1061);
nand U2001 (N_2001,N_1794,N_1627);
and U2002 (N_2002,N_1455,N_1765);
or U2003 (N_2003,N_1001,N_1870);
xor U2004 (N_2004,N_1380,N_1043);
and U2005 (N_2005,N_1178,N_1593);
xnor U2006 (N_2006,N_1493,N_1138);
xnor U2007 (N_2007,N_1237,N_1480);
and U2008 (N_2008,N_1093,N_1559);
nor U2009 (N_2009,N_1787,N_1377);
nor U2010 (N_2010,N_1321,N_1430);
or U2011 (N_2011,N_1920,N_1468);
nor U2012 (N_2012,N_1740,N_1501);
and U2013 (N_2013,N_1716,N_1616);
nor U2014 (N_2014,N_1766,N_1524);
or U2015 (N_2015,N_1102,N_1204);
or U2016 (N_2016,N_1585,N_1503);
nand U2017 (N_2017,N_1365,N_1550);
nor U2018 (N_2018,N_1723,N_1763);
and U2019 (N_2019,N_1890,N_1844);
nor U2020 (N_2020,N_1450,N_1908);
or U2021 (N_2021,N_1255,N_1996);
or U2022 (N_2022,N_1213,N_1872);
nor U2023 (N_2023,N_1999,N_1597);
nor U2024 (N_2024,N_1910,N_1047);
or U2025 (N_2025,N_1913,N_1124);
and U2026 (N_2026,N_1816,N_1303);
xnor U2027 (N_2027,N_1170,N_1697);
nor U2028 (N_2028,N_1532,N_1878);
xor U2029 (N_2029,N_1614,N_1301);
xnor U2030 (N_2030,N_1055,N_1647);
and U2031 (N_2031,N_1214,N_1580);
nand U2032 (N_2032,N_1531,N_1635);
nand U2033 (N_2033,N_1352,N_1820);
nand U2034 (N_2034,N_1744,N_1025);
or U2035 (N_2035,N_1200,N_1813);
and U2036 (N_2036,N_1322,N_1408);
nand U2037 (N_2037,N_1160,N_1489);
and U2038 (N_2038,N_1404,N_1161);
xor U2039 (N_2039,N_1021,N_1305);
xnor U2040 (N_2040,N_1695,N_1613);
xnor U2041 (N_2041,N_1173,N_1278);
xor U2042 (N_2042,N_1112,N_1109);
xor U2043 (N_2043,N_1714,N_1041);
nor U2044 (N_2044,N_1015,N_1054);
and U2045 (N_2045,N_1642,N_1163);
nand U2046 (N_2046,N_1414,N_1022);
nand U2047 (N_2047,N_1909,N_1181);
nor U2048 (N_2048,N_1098,N_1222);
nand U2049 (N_2049,N_1148,N_1106);
nand U2050 (N_2050,N_1590,N_1553);
xnor U2051 (N_2051,N_1520,N_1267);
nor U2052 (N_2052,N_1494,N_1554);
or U2053 (N_2053,N_1522,N_1737);
nand U2054 (N_2054,N_1973,N_1433);
nor U2055 (N_2055,N_1634,N_1065);
xnor U2056 (N_2056,N_1857,N_1435);
nand U2057 (N_2057,N_1626,N_1502);
and U2058 (N_2058,N_1917,N_1608);
or U2059 (N_2059,N_1272,N_1361);
xor U2060 (N_2060,N_1762,N_1534);
xnor U2061 (N_2061,N_1758,N_1883);
nand U2062 (N_2062,N_1957,N_1491);
nor U2063 (N_2063,N_1351,N_1072);
and U2064 (N_2064,N_1075,N_1335);
nand U2065 (N_2065,N_1464,N_1241);
nand U2066 (N_2066,N_1226,N_1159);
nor U2067 (N_2067,N_1423,N_1736);
or U2068 (N_2068,N_1829,N_1775);
xor U2069 (N_2069,N_1839,N_1067);
nand U2070 (N_2070,N_1177,N_1333);
xnor U2071 (N_2071,N_1753,N_1235);
or U2072 (N_2072,N_1541,N_1013);
or U2073 (N_2073,N_1094,N_1891);
xnor U2074 (N_2074,N_1183,N_1980);
xnor U2075 (N_2075,N_1718,N_1436);
or U2076 (N_2076,N_1115,N_1769);
nor U2077 (N_2077,N_1947,N_1584);
nor U2078 (N_2078,N_1289,N_1245);
or U2079 (N_2079,N_1664,N_1552);
and U2080 (N_2080,N_1147,N_1398);
nor U2081 (N_2081,N_1448,N_1258);
nor U2082 (N_2082,N_1686,N_1709);
xnor U2083 (N_2083,N_1533,N_1789);
nand U2084 (N_2084,N_1997,N_1964);
nand U2085 (N_2085,N_1291,N_1924);
xnor U2086 (N_2086,N_1332,N_1700);
xor U2087 (N_2087,N_1154,N_1195);
and U2088 (N_2088,N_1317,N_1757);
and U2089 (N_2089,N_1347,N_1282);
nor U2090 (N_2090,N_1251,N_1228);
nor U2091 (N_2091,N_1643,N_1132);
and U2092 (N_2092,N_1837,N_1174);
and U2093 (N_2093,N_1962,N_1044);
nor U2094 (N_2094,N_1928,N_1551);
xnor U2095 (N_2095,N_1394,N_1326);
and U2096 (N_2096,N_1268,N_1578);
xnor U2097 (N_2097,N_1529,N_1682);
nand U2098 (N_2098,N_1687,N_1633);
nor U2099 (N_2099,N_1199,N_1086);
xnor U2100 (N_2100,N_1095,N_1416);
or U2101 (N_2101,N_1986,N_1281);
nor U2102 (N_2102,N_1549,N_1063);
nand U2103 (N_2103,N_1208,N_1421);
nand U2104 (N_2104,N_1655,N_1712);
or U2105 (N_2105,N_1396,N_1573);
xnor U2106 (N_2106,N_1311,N_1219);
nand U2107 (N_2107,N_1806,N_1577);
or U2108 (N_2108,N_1447,N_1755);
nor U2109 (N_2109,N_1631,N_1561);
xor U2110 (N_2110,N_1851,N_1636);
and U2111 (N_2111,N_1020,N_1466);
and U2112 (N_2112,N_1772,N_1711);
nand U2113 (N_2113,N_1587,N_1370);
and U2114 (N_2114,N_1230,N_1900);
or U2115 (N_2115,N_1030,N_1749);
nand U2116 (N_2116,N_1952,N_1676);
or U2117 (N_2117,N_1732,N_1701);
nand U2118 (N_2118,N_1412,N_1345);
xor U2119 (N_2119,N_1855,N_1899);
or U2120 (N_2120,N_1420,N_1796);
xor U2121 (N_2121,N_1788,N_1343);
or U2122 (N_2122,N_1638,N_1456);
xnor U2123 (N_2123,N_1440,N_1988);
or U2124 (N_2124,N_1939,N_1336);
or U2125 (N_2125,N_1034,N_1128);
and U2126 (N_2126,N_1292,N_1624);
and U2127 (N_2127,N_1426,N_1401);
nand U2128 (N_2128,N_1100,N_1166);
nand U2129 (N_2129,N_1706,N_1575);
and U2130 (N_2130,N_1096,N_1266);
and U2131 (N_2131,N_1665,N_1340);
xnor U2132 (N_2132,N_1386,N_1497);
nand U2133 (N_2133,N_1231,N_1881);
nand U2134 (N_2134,N_1995,N_1607);
nand U2135 (N_2135,N_1410,N_1261);
nor U2136 (N_2136,N_1923,N_1894);
nand U2137 (N_2137,N_1803,N_1530);
xor U2138 (N_2138,N_1859,N_1216);
xnor U2139 (N_2139,N_1594,N_1259);
nor U2140 (N_2140,N_1821,N_1505);
nand U2141 (N_2141,N_1619,N_1157);
nand U2142 (N_2142,N_1233,N_1925);
nor U2143 (N_2143,N_1622,N_1754);
nor U2144 (N_2144,N_1595,N_1203);
and U2145 (N_2145,N_1084,N_1629);
and U2146 (N_2146,N_1387,N_1557);
nand U2147 (N_2147,N_1571,N_1419);
and U2148 (N_2148,N_1432,N_1521);
nor U2149 (N_2149,N_1373,N_1186);
nor U2150 (N_2150,N_1428,N_1846);
nor U2151 (N_2151,N_1271,N_1699);
and U2152 (N_2152,N_1562,N_1201);
xor U2153 (N_2153,N_1838,N_1091);
nor U2154 (N_2154,N_1669,N_1652);
xnor U2155 (N_2155,N_1623,N_1003);
or U2156 (N_2156,N_1116,N_1739);
or U2157 (N_2157,N_1232,N_1029);
xnor U2158 (N_2158,N_1300,N_1889);
or U2159 (N_2159,N_1689,N_1366);
nand U2160 (N_2160,N_1004,N_1472);
nand U2161 (N_2161,N_1684,N_1628);
nor U2162 (N_2162,N_1783,N_1114);
nor U2163 (N_2163,N_1514,N_1184);
or U2164 (N_2164,N_1108,N_1053);
xnor U2165 (N_2165,N_1008,N_1290);
nor U2166 (N_2166,N_1475,N_1621);
nor U2167 (N_2167,N_1018,N_1127);
nor U2168 (N_2168,N_1485,N_1062);
or U2169 (N_2169,N_1984,N_1904);
nor U2170 (N_2170,N_1598,N_1005);
xor U2171 (N_2171,N_1405,N_1297);
nand U2172 (N_2172,N_1617,N_1210);
and U2173 (N_2173,N_1499,N_1037);
nand U2174 (N_2174,N_1945,N_1651);
and U2175 (N_2175,N_1922,N_1158);
and U2176 (N_2176,N_1673,N_1819);
or U2177 (N_2177,N_1444,N_1759);
xor U2178 (N_2178,N_1971,N_1832);
nor U2179 (N_2179,N_1705,N_1197);
xor U2180 (N_2180,N_1659,N_1082);
and U2181 (N_2181,N_1645,N_1523);
xnor U2182 (N_2182,N_1660,N_1779);
nor U2183 (N_2183,N_1615,N_1318);
nand U2184 (N_2184,N_1936,N_1884);
nor U2185 (N_2185,N_1861,N_1639);
and U2186 (N_2186,N_1312,N_1830);
nand U2187 (N_2187,N_1747,N_1583);
nand U2188 (N_2188,N_1745,N_1896);
xnor U2189 (N_2189,N_1257,N_1556);
xor U2190 (N_2190,N_1911,N_1589);
nand U2191 (N_2191,N_1600,N_1512);
and U2192 (N_2192,N_1176,N_1653);
and U2193 (N_2193,N_1579,N_1049);
nor U2194 (N_2194,N_1058,N_1007);
nand U2195 (N_2195,N_1938,N_1515);
nor U2196 (N_2196,N_1536,N_1866);
or U2197 (N_2197,N_1721,N_1346);
or U2198 (N_2198,N_1814,N_1059);
or U2199 (N_2199,N_1375,N_1954);
or U2200 (N_2200,N_1169,N_1193);
or U2201 (N_2201,N_1354,N_1823);
or U2202 (N_2202,N_1833,N_1519);
xnor U2203 (N_2203,N_1471,N_1513);
and U2204 (N_2204,N_1798,N_1850);
and U2205 (N_2205,N_1319,N_1630);
nand U2206 (N_2206,N_1473,N_1175);
nor U2207 (N_2207,N_1249,N_1134);
nor U2208 (N_2208,N_1090,N_1875);
xnor U2209 (N_2209,N_1641,N_1189);
nor U2210 (N_2210,N_1761,N_1194);
and U2211 (N_2211,N_1567,N_1205);
nand U2212 (N_2212,N_1331,N_1726);
and U2213 (N_2213,N_1088,N_1618);
nor U2214 (N_2214,N_1596,N_1477);
xor U2215 (N_2215,N_1168,N_1284);
xnor U2216 (N_2216,N_1842,N_1767);
and U2217 (N_2217,N_1256,N_1707);
xor U2218 (N_2218,N_1588,N_1240);
nor U2219 (N_2219,N_1637,N_1264);
nand U2220 (N_2220,N_1155,N_1625);
nand U2221 (N_2221,N_1474,N_1402);
xor U2222 (N_2222,N_1974,N_1307);
and U2223 (N_2223,N_1068,N_1555);
or U2224 (N_2224,N_1934,N_1677);
or U2225 (N_2225,N_1895,N_1323);
or U2226 (N_2226,N_1042,N_1150);
xnor U2227 (N_2227,N_1191,N_1886);
or U2228 (N_2228,N_1118,N_1733);
nor U2229 (N_2229,N_1792,N_1446);
xor U2230 (N_2230,N_1805,N_1657);
and U2231 (N_2231,N_1632,N_1039);
nand U2232 (N_2232,N_1977,N_1591);
nor U2233 (N_2233,N_1927,N_1164);
nand U2234 (N_2234,N_1569,N_1675);
and U2235 (N_2235,N_1449,N_1247);
xnor U2236 (N_2236,N_1717,N_1965);
nand U2237 (N_2237,N_1431,N_1269);
nand U2238 (N_2238,N_1000,N_1339);
nor U2239 (N_2239,N_1295,N_1946);
nor U2240 (N_2240,N_1143,N_1836);
and U2241 (N_2241,N_1488,N_1198);
or U2242 (N_2242,N_1860,N_1125);
nor U2243 (N_2243,N_1688,N_1454);
nor U2244 (N_2244,N_1831,N_1678);
or U2245 (N_2245,N_1422,N_1356);
and U2246 (N_2246,N_1804,N_1451);
or U2247 (N_2247,N_1461,N_1847);
or U2248 (N_2248,N_1970,N_1683);
nand U2249 (N_2249,N_1320,N_1563);
nor U2250 (N_2250,N_1381,N_1242);
or U2251 (N_2251,N_1570,N_1288);
and U2252 (N_2252,N_1192,N_1076);
or U2253 (N_2253,N_1864,N_1824);
and U2254 (N_2254,N_1481,N_1774);
xnor U2255 (N_2255,N_1012,N_1385);
nor U2256 (N_2256,N_1901,N_1324);
nor U2257 (N_2257,N_1854,N_1685);
xor U2258 (N_2258,N_1538,N_1378);
or U2259 (N_2259,N_1452,N_1048);
or U2260 (N_2260,N_1863,N_1442);
xnor U2261 (N_2261,N_1834,N_1293);
xnor U2262 (N_2262,N_1907,N_1807);
or U2263 (N_2263,N_1565,N_1800);
xnor U2264 (N_2264,N_1897,N_1006);
or U2265 (N_2265,N_1942,N_1188);
and U2266 (N_2266,N_1145,N_1179);
nor U2267 (N_2267,N_1244,N_1119);
and U2268 (N_2268,N_1182,N_1713);
or U2269 (N_2269,N_1564,N_1526);
or U2270 (N_2270,N_1500,N_1342);
and U2271 (N_2271,N_1703,N_1056);
or U2272 (N_2272,N_1040,N_1328);
nor U2273 (N_2273,N_1142,N_1724);
nor U2274 (N_2274,N_1666,N_1202);
xnor U2275 (N_2275,N_1959,N_1975);
nor U2276 (N_2276,N_1028,N_1799);
or U2277 (N_2277,N_1443,N_1490);
xnor U2278 (N_2278,N_1882,N_1963);
xor U2279 (N_2279,N_1438,N_1960);
and U2280 (N_2280,N_1606,N_1137);
or U2281 (N_2281,N_1852,N_1495);
and U2282 (N_2282,N_1105,N_1372);
or U2283 (N_2283,N_1994,N_1131);
xnor U2284 (N_2284,N_1399,N_1967);
nand U2285 (N_2285,N_1395,N_1727);
and U2286 (N_2286,N_1704,N_1310);
or U2287 (N_2287,N_1640,N_1384);
or U2288 (N_2288,N_1141,N_1254);
xor U2289 (N_2289,N_1873,N_1708);
xnor U2290 (N_2290,N_1092,N_1341);
or U2291 (N_2291,N_1252,N_1113);
xnor U2292 (N_2292,N_1933,N_1123);
nand U2293 (N_2293,N_1802,N_1646);
nand U2294 (N_2294,N_1835,N_1045);
xnor U2295 (N_2295,N_1892,N_1729);
or U2296 (N_2296,N_1893,N_1064);
nor U2297 (N_2297,N_1698,N_1280);
or U2298 (N_2298,N_1620,N_1014);
and U2299 (N_2299,N_1809,N_1434);
or U2300 (N_2300,N_1770,N_1560);
or U2301 (N_2301,N_1248,N_1702);
or U2302 (N_2302,N_1275,N_1010);
or U2303 (N_2303,N_1601,N_1283);
and U2304 (N_2304,N_1528,N_1407);
nand U2305 (N_2305,N_1060,N_1476);
nand U2306 (N_2306,N_1050,N_1427);
nor U2307 (N_2307,N_1167,N_1424);
or U2308 (N_2308,N_1843,N_1773);
or U2309 (N_2309,N_1391,N_1825);
xnor U2310 (N_2310,N_1644,N_1187);
and U2311 (N_2311,N_1841,N_1019);
xor U2312 (N_2312,N_1360,N_1879);
or U2313 (N_2313,N_1912,N_1990);
or U2314 (N_2314,N_1741,N_1956);
nand U2315 (N_2315,N_1299,N_1720);
nor U2316 (N_2316,N_1916,N_1535);
nor U2317 (N_2317,N_1171,N_1822);
nand U2318 (N_2318,N_1991,N_1782);
xor U2319 (N_2319,N_1696,N_1129);
nand U2320 (N_2320,N_1218,N_1797);
and U2321 (N_2321,N_1415,N_1070);
nor U2322 (N_2322,N_1350,N_1462);
and U2323 (N_2323,N_1868,N_1856);
nand U2324 (N_2324,N_1888,N_1458);
and U2325 (N_2325,N_1215,N_1057);
xnor U2326 (N_2326,N_1826,N_1981);
or U2327 (N_2327,N_1220,N_1778);
xnor U2328 (N_2328,N_1517,N_1349);
nor U2329 (N_2329,N_1389,N_1496);
nor U2330 (N_2330,N_1487,N_1080);
nor U2331 (N_2331,N_1140,N_1110);
xnor U2332 (N_2332,N_1694,N_1966);
nor U2333 (N_2333,N_1603,N_1876);
nand U2334 (N_2334,N_1217,N_1316);
and U2335 (N_2335,N_1149,N_1101);
nor U2336 (N_2336,N_1085,N_1661);
xor U2337 (N_2337,N_1035,N_1576);
xor U2338 (N_2338,N_1547,N_1120);
nor U2339 (N_2339,N_1172,N_1367);
nor U2340 (N_2340,N_1469,N_1382);
nor U2341 (N_2341,N_1355,N_1815);
xnor U2342 (N_2342,N_1107,N_1812);
nor U2343 (N_2343,N_1568,N_1719);
nor U2344 (N_2344,N_1898,N_1304);
nor U2345 (N_2345,N_1944,N_1046);
nor U2346 (N_2346,N_1374,N_1031);
or U2347 (N_2347,N_1270,N_1441);
xnor U2348 (N_2348,N_1650,N_1506);
or U2349 (N_2349,N_1949,N_1081);
and U2350 (N_2350,N_1581,N_1152);
nand U2351 (N_2351,N_1992,N_1906);
nand U2352 (N_2352,N_1950,N_1406);
or U2353 (N_2353,N_1818,N_1781);
xor U2354 (N_2354,N_1544,N_1425);
or U2355 (N_2355,N_1302,N_1453);
nor U2356 (N_2356,N_1731,N_1691);
nor U2357 (N_2357,N_1027,N_1246);
or U2358 (N_2358,N_1486,N_1734);
and U2359 (N_2359,N_1122,N_1791);
xnor U2360 (N_2360,N_1546,N_1445);
xnor U2361 (N_2361,N_1961,N_1368);
and U2362 (N_2362,N_1253,N_1602);
and U2363 (N_2363,N_1089,N_1274);
nor U2364 (N_2364,N_1077,N_1146);
xnor U2365 (N_2365,N_1853,N_1483);
and U2366 (N_2366,N_1752,N_1038);
nor U2367 (N_2367,N_1470,N_1599);
nand U2368 (N_2368,N_1905,N_1674);
xor U2369 (N_2369,N_1941,N_1390);
xor U2370 (N_2370,N_1828,N_1180);
or U2371 (N_2371,N_1211,N_1511);
and U2372 (N_2372,N_1662,N_1279);
nand U2373 (N_2373,N_1358,N_1315);
xnor U2374 (N_2374,N_1403,N_1073);
xnor U2375 (N_2375,N_1069,N_1654);
or U2376 (N_2376,N_1545,N_1735);
nand U2377 (N_2377,N_1325,N_1418);
or U2378 (N_2378,N_1071,N_1457);
or U2379 (N_2379,N_1760,N_1238);
nand U2380 (N_2380,N_1880,N_1224);
nand U2381 (N_2381,N_1286,N_1926);
nand U2382 (N_2382,N_1586,N_1771);
and U2383 (N_2383,N_1784,N_1572);
xnor U2384 (N_2384,N_1276,N_1314);
nor U2385 (N_2385,N_1026,N_1681);
nor U2386 (N_2386,N_1392,N_1658);
or U2387 (N_2387,N_1097,N_1672);
nand U2388 (N_2388,N_1207,N_1337);
xnor U2389 (N_2389,N_1227,N_1103);
nor U2390 (N_2390,N_1052,N_1982);
nor U2391 (N_2391,N_1265,N_1348);
nor U2392 (N_2392,N_1225,N_1376);
nand U2393 (N_2393,N_1915,N_1362);
nor U2394 (N_2394,N_1811,N_1680);
or U2395 (N_2395,N_1751,N_1429);
and U2396 (N_2396,N_1958,N_1969);
xnor U2397 (N_2397,N_1871,N_1785);
and U2398 (N_2398,N_1397,N_1649);
or U2399 (N_2399,N_1463,N_1921);
and U2400 (N_2400,N_1036,N_1298);
nand U2401 (N_2401,N_1359,N_1692);
xnor U2402 (N_2402,N_1239,N_1801);
nand U2403 (N_2403,N_1083,N_1032);
or U2404 (N_2404,N_1605,N_1937);
or U2405 (N_2405,N_1542,N_1849);
or U2406 (N_2406,N_1260,N_1327);
nand U2407 (N_2407,N_1287,N_1306);
and U2408 (N_2408,N_1329,N_1940);
and U2409 (N_2409,N_1510,N_1409);
or U2410 (N_2410,N_1467,N_1002);
and U2411 (N_2411,N_1604,N_1989);
nor U2412 (N_2412,N_1948,N_1943);
nand U2413 (N_2413,N_1743,N_1411);
and U2414 (N_2414,N_1263,N_1111);
nor U2415 (N_2415,N_1117,N_1371);
xnor U2416 (N_2416,N_1011,N_1715);
xor U2417 (N_2417,N_1756,N_1236);
or U2418 (N_2418,N_1285,N_1492);
nor U2419 (N_2419,N_1887,N_1104);
or U2420 (N_2420,N_1874,N_1344);
nor U2421 (N_2421,N_1776,N_1417);
nor U2422 (N_2422,N_1221,N_1670);
and U2423 (N_2423,N_1478,N_1525);
xnor U2424 (N_2424,N_1139,N_1196);
xnor U2425 (N_2425,N_1592,N_1250);
and U2426 (N_2426,N_1330,N_1223);
nor U2427 (N_2427,N_1273,N_1983);
nand U2428 (N_2428,N_1612,N_1017);
xor U2429 (N_2429,N_1507,N_1338);
xor U2430 (N_2430,N_1185,N_1364);
nand U2431 (N_2431,N_1133,N_1079);
nor U2432 (N_2432,N_1935,N_1135);
or U2433 (N_2433,N_1931,N_1827);
xor U2434 (N_2434,N_1051,N_1725);
nand U2435 (N_2435,N_1817,N_1509);
and U2436 (N_2436,N_1610,N_1460);
nand U2437 (N_2437,N_1130,N_1126);
or U2438 (N_2438,N_1611,N_1978);
nor U2439 (N_2439,N_1439,N_1858);
and U2440 (N_2440,N_1566,N_1979);
nor U2441 (N_2441,N_1667,N_1777);
and U2442 (N_2442,N_1987,N_1877);
nand U2443 (N_2443,N_1209,N_1516);
nor U2444 (N_2444,N_1465,N_1537);
nand U2445 (N_2445,N_1919,N_1929);
nand U2446 (N_2446,N_1121,N_1388);
xor U2447 (N_2447,N_1722,N_1024);
or U2448 (N_2448,N_1527,N_1151);
xor U2449 (N_2449,N_1459,N_1206);
and U2450 (N_2450,N_1993,N_1998);
xnor U2451 (N_2451,N_1144,N_1930);
and U2452 (N_2452,N_1710,N_1504);
and U2453 (N_2453,N_1539,N_1479);
and U2454 (N_2454,N_1369,N_1790);
and U2455 (N_2455,N_1484,N_1296);
or U2456 (N_2456,N_1609,N_1951);
nand U2457 (N_2457,N_1243,N_1548);
xnor U2458 (N_2458,N_1742,N_1968);
xor U2459 (N_2459,N_1023,N_1136);
nor U2460 (N_2460,N_1190,N_1748);
nor U2461 (N_2461,N_1540,N_1648);
or U2462 (N_2462,N_1016,N_1400);
xor U2463 (N_2463,N_1543,N_1156);
nand U2464 (N_2464,N_1074,N_1165);
or U2465 (N_2465,N_1728,N_1867);
xnor U2466 (N_2466,N_1313,N_1099);
or U2467 (N_2467,N_1308,N_1914);
and U2468 (N_2468,N_1383,N_1558);
or U2469 (N_2469,N_1656,N_1972);
xor U2470 (N_2470,N_1848,N_1334);
xnor U2471 (N_2471,N_1212,N_1869);
nor U2472 (N_2472,N_1845,N_1730);
and U2473 (N_2473,N_1780,N_1363);
nor U2474 (N_2474,N_1768,N_1309);
and U2475 (N_2475,N_1574,N_1508);
and U2476 (N_2476,N_1087,N_1795);
xor U2477 (N_2477,N_1033,N_1668);
nor U2478 (N_2478,N_1750,N_1229);
or U2479 (N_2479,N_1393,N_1746);
nand U2480 (N_2480,N_1413,N_1066);
nor U2481 (N_2481,N_1865,N_1482);
nand U2482 (N_2482,N_1903,N_1353);
xor U2483 (N_2483,N_1277,N_1162);
and U2484 (N_2484,N_1840,N_1902);
or U2485 (N_2485,N_1498,N_1808);
or U2486 (N_2486,N_1985,N_1078);
xnor U2487 (N_2487,N_1437,N_1932);
xor U2488 (N_2488,N_1294,N_1693);
nor U2489 (N_2489,N_1764,N_1955);
nand U2490 (N_2490,N_1679,N_1671);
nand U2491 (N_2491,N_1379,N_1862);
xor U2492 (N_2492,N_1953,N_1518);
nor U2493 (N_2493,N_1262,N_1234);
or U2494 (N_2494,N_1793,N_1786);
and U2495 (N_2495,N_1009,N_1582);
and U2496 (N_2496,N_1357,N_1663);
nand U2497 (N_2497,N_1153,N_1690);
or U2498 (N_2498,N_1976,N_1810);
nand U2499 (N_2499,N_1885,N_1918);
or U2500 (N_2500,N_1331,N_1840);
or U2501 (N_2501,N_1079,N_1075);
or U2502 (N_2502,N_1173,N_1794);
and U2503 (N_2503,N_1323,N_1800);
nor U2504 (N_2504,N_1504,N_1037);
and U2505 (N_2505,N_1252,N_1652);
and U2506 (N_2506,N_1564,N_1140);
nor U2507 (N_2507,N_1925,N_1041);
nor U2508 (N_2508,N_1153,N_1875);
nor U2509 (N_2509,N_1787,N_1689);
or U2510 (N_2510,N_1613,N_1828);
and U2511 (N_2511,N_1940,N_1345);
or U2512 (N_2512,N_1770,N_1124);
xnor U2513 (N_2513,N_1498,N_1724);
nor U2514 (N_2514,N_1837,N_1288);
nand U2515 (N_2515,N_1724,N_1901);
xnor U2516 (N_2516,N_1013,N_1511);
xor U2517 (N_2517,N_1877,N_1772);
nor U2518 (N_2518,N_1826,N_1533);
xnor U2519 (N_2519,N_1269,N_1488);
or U2520 (N_2520,N_1340,N_1059);
nor U2521 (N_2521,N_1584,N_1076);
or U2522 (N_2522,N_1408,N_1371);
xnor U2523 (N_2523,N_1779,N_1535);
nor U2524 (N_2524,N_1053,N_1472);
or U2525 (N_2525,N_1692,N_1189);
nor U2526 (N_2526,N_1620,N_1848);
xnor U2527 (N_2527,N_1518,N_1309);
xor U2528 (N_2528,N_1525,N_1796);
xnor U2529 (N_2529,N_1491,N_1631);
or U2530 (N_2530,N_1977,N_1803);
and U2531 (N_2531,N_1793,N_1168);
nor U2532 (N_2532,N_1729,N_1992);
xor U2533 (N_2533,N_1760,N_1691);
or U2534 (N_2534,N_1321,N_1337);
nand U2535 (N_2535,N_1750,N_1970);
nand U2536 (N_2536,N_1310,N_1493);
nor U2537 (N_2537,N_1633,N_1438);
xnor U2538 (N_2538,N_1149,N_1301);
nor U2539 (N_2539,N_1623,N_1516);
xnor U2540 (N_2540,N_1010,N_1011);
or U2541 (N_2541,N_1487,N_1482);
xor U2542 (N_2542,N_1817,N_1671);
nor U2543 (N_2543,N_1875,N_1313);
xor U2544 (N_2544,N_1480,N_1238);
xnor U2545 (N_2545,N_1875,N_1179);
nand U2546 (N_2546,N_1545,N_1940);
nand U2547 (N_2547,N_1455,N_1975);
and U2548 (N_2548,N_1843,N_1805);
and U2549 (N_2549,N_1233,N_1391);
nor U2550 (N_2550,N_1274,N_1474);
xnor U2551 (N_2551,N_1641,N_1890);
xnor U2552 (N_2552,N_1924,N_1889);
and U2553 (N_2553,N_1179,N_1064);
and U2554 (N_2554,N_1674,N_1127);
or U2555 (N_2555,N_1366,N_1427);
xnor U2556 (N_2556,N_1152,N_1376);
and U2557 (N_2557,N_1592,N_1907);
nor U2558 (N_2558,N_1863,N_1342);
nand U2559 (N_2559,N_1010,N_1291);
nor U2560 (N_2560,N_1117,N_1867);
nand U2561 (N_2561,N_1005,N_1151);
and U2562 (N_2562,N_1278,N_1767);
or U2563 (N_2563,N_1241,N_1355);
nor U2564 (N_2564,N_1638,N_1708);
xor U2565 (N_2565,N_1600,N_1203);
or U2566 (N_2566,N_1466,N_1817);
or U2567 (N_2567,N_1335,N_1170);
xnor U2568 (N_2568,N_1796,N_1234);
nand U2569 (N_2569,N_1802,N_1408);
or U2570 (N_2570,N_1330,N_1160);
xor U2571 (N_2571,N_1002,N_1348);
nand U2572 (N_2572,N_1583,N_1690);
xnor U2573 (N_2573,N_1660,N_1372);
or U2574 (N_2574,N_1147,N_1745);
xor U2575 (N_2575,N_1099,N_1623);
nor U2576 (N_2576,N_1079,N_1361);
xor U2577 (N_2577,N_1959,N_1304);
xor U2578 (N_2578,N_1453,N_1077);
nor U2579 (N_2579,N_1317,N_1163);
nor U2580 (N_2580,N_1902,N_1857);
xnor U2581 (N_2581,N_1683,N_1700);
and U2582 (N_2582,N_1422,N_1934);
nand U2583 (N_2583,N_1935,N_1892);
and U2584 (N_2584,N_1617,N_1627);
nor U2585 (N_2585,N_1363,N_1807);
nor U2586 (N_2586,N_1446,N_1246);
nor U2587 (N_2587,N_1569,N_1695);
nor U2588 (N_2588,N_1498,N_1120);
or U2589 (N_2589,N_1623,N_1281);
nand U2590 (N_2590,N_1182,N_1307);
nor U2591 (N_2591,N_1821,N_1165);
nand U2592 (N_2592,N_1017,N_1990);
xnor U2593 (N_2593,N_1288,N_1072);
and U2594 (N_2594,N_1148,N_1323);
or U2595 (N_2595,N_1677,N_1957);
nand U2596 (N_2596,N_1659,N_1976);
or U2597 (N_2597,N_1117,N_1320);
and U2598 (N_2598,N_1384,N_1613);
xor U2599 (N_2599,N_1659,N_1484);
or U2600 (N_2600,N_1747,N_1955);
and U2601 (N_2601,N_1790,N_1031);
nor U2602 (N_2602,N_1100,N_1430);
nor U2603 (N_2603,N_1519,N_1787);
xor U2604 (N_2604,N_1512,N_1375);
nor U2605 (N_2605,N_1601,N_1649);
nor U2606 (N_2606,N_1628,N_1482);
and U2607 (N_2607,N_1087,N_1375);
nor U2608 (N_2608,N_1720,N_1149);
xor U2609 (N_2609,N_1868,N_1070);
and U2610 (N_2610,N_1206,N_1407);
nor U2611 (N_2611,N_1659,N_1415);
nor U2612 (N_2612,N_1700,N_1334);
and U2613 (N_2613,N_1728,N_1619);
nand U2614 (N_2614,N_1150,N_1068);
nor U2615 (N_2615,N_1322,N_1164);
nor U2616 (N_2616,N_1678,N_1199);
xnor U2617 (N_2617,N_1408,N_1032);
or U2618 (N_2618,N_1480,N_1455);
nor U2619 (N_2619,N_1041,N_1000);
nor U2620 (N_2620,N_1135,N_1042);
xor U2621 (N_2621,N_1729,N_1293);
nand U2622 (N_2622,N_1419,N_1099);
and U2623 (N_2623,N_1329,N_1693);
nor U2624 (N_2624,N_1350,N_1025);
xor U2625 (N_2625,N_1065,N_1063);
xnor U2626 (N_2626,N_1499,N_1311);
and U2627 (N_2627,N_1961,N_1069);
nor U2628 (N_2628,N_1657,N_1989);
or U2629 (N_2629,N_1255,N_1861);
nor U2630 (N_2630,N_1082,N_1362);
or U2631 (N_2631,N_1110,N_1541);
nand U2632 (N_2632,N_1769,N_1305);
xor U2633 (N_2633,N_1591,N_1785);
and U2634 (N_2634,N_1676,N_1420);
nand U2635 (N_2635,N_1853,N_1604);
or U2636 (N_2636,N_1572,N_1766);
and U2637 (N_2637,N_1624,N_1012);
nor U2638 (N_2638,N_1598,N_1324);
xor U2639 (N_2639,N_1368,N_1800);
xnor U2640 (N_2640,N_1241,N_1177);
or U2641 (N_2641,N_1472,N_1016);
or U2642 (N_2642,N_1194,N_1461);
xor U2643 (N_2643,N_1788,N_1048);
nand U2644 (N_2644,N_1250,N_1031);
nor U2645 (N_2645,N_1567,N_1101);
nand U2646 (N_2646,N_1967,N_1973);
and U2647 (N_2647,N_1424,N_1559);
nor U2648 (N_2648,N_1156,N_1571);
nand U2649 (N_2649,N_1608,N_1315);
or U2650 (N_2650,N_1091,N_1043);
and U2651 (N_2651,N_1126,N_1265);
and U2652 (N_2652,N_1266,N_1627);
and U2653 (N_2653,N_1370,N_1618);
nand U2654 (N_2654,N_1786,N_1911);
and U2655 (N_2655,N_1403,N_1412);
xnor U2656 (N_2656,N_1997,N_1600);
xor U2657 (N_2657,N_1756,N_1311);
nor U2658 (N_2658,N_1676,N_1759);
xor U2659 (N_2659,N_1088,N_1923);
xor U2660 (N_2660,N_1763,N_1686);
nor U2661 (N_2661,N_1830,N_1048);
and U2662 (N_2662,N_1672,N_1610);
xor U2663 (N_2663,N_1280,N_1233);
nor U2664 (N_2664,N_1893,N_1260);
xor U2665 (N_2665,N_1069,N_1975);
or U2666 (N_2666,N_1897,N_1186);
xnor U2667 (N_2667,N_1649,N_1715);
nor U2668 (N_2668,N_1912,N_1622);
nand U2669 (N_2669,N_1860,N_1550);
nand U2670 (N_2670,N_1845,N_1338);
and U2671 (N_2671,N_1727,N_1255);
nor U2672 (N_2672,N_1097,N_1990);
or U2673 (N_2673,N_1351,N_1575);
nand U2674 (N_2674,N_1769,N_1197);
nor U2675 (N_2675,N_1919,N_1150);
nand U2676 (N_2676,N_1272,N_1382);
nand U2677 (N_2677,N_1355,N_1690);
and U2678 (N_2678,N_1424,N_1213);
or U2679 (N_2679,N_1245,N_1565);
nand U2680 (N_2680,N_1779,N_1380);
xnor U2681 (N_2681,N_1369,N_1072);
nor U2682 (N_2682,N_1113,N_1295);
xor U2683 (N_2683,N_1155,N_1775);
nor U2684 (N_2684,N_1559,N_1378);
xnor U2685 (N_2685,N_1221,N_1808);
or U2686 (N_2686,N_1071,N_1901);
or U2687 (N_2687,N_1714,N_1966);
nand U2688 (N_2688,N_1974,N_1410);
and U2689 (N_2689,N_1948,N_1812);
xor U2690 (N_2690,N_1746,N_1674);
xnor U2691 (N_2691,N_1394,N_1956);
or U2692 (N_2692,N_1078,N_1617);
and U2693 (N_2693,N_1056,N_1961);
nand U2694 (N_2694,N_1927,N_1821);
and U2695 (N_2695,N_1069,N_1969);
nand U2696 (N_2696,N_1243,N_1026);
nor U2697 (N_2697,N_1441,N_1494);
xor U2698 (N_2698,N_1009,N_1848);
xor U2699 (N_2699,N_1102,N_1899);
and U2700 (N_2700,N_1718,N_1563);
nor U2701 (N_2701,N_1016,N_1721);
nand U2702 (N_2702,N_1983,N_1613);
nor U2703 (N_2703,N_1270,N_1070);
nor U2704 (N_2704,N_1901,N_1510);
xor U2705 (N_2705,N_1738,N_1603);
xnor U2706 (N_2706,N_1856,N_1050);
nand U2707 (N_2707,N_1442,N_1944);
xnor U2708 (N_2708,N_1542,N_1505);
xor U2709 (N_2709,N_1374,N_1912);
and U2710 (N_2710,N_1768,N_1851);
nand U2711 (N_2711,N_1967,N_1655);
and U2712 (N_2712,N_1331,N_1725);
xor U2713 (N_2713,N_1691,N_1476);
or U2714 (N_2714,N_1888,N_1445);
nand U2715 (N_2715,N_1418,N_1140);
xnor U2716 (N_2716,N_1174,N_1648);
and U2717 (N_2717,N_1209,N_1459);
xor U2718 (N_2718,N_1329,N_1873);
or U2719 (N_2719,N_1091,N_1205);
nor U2720 (N_2720,N_1713,N_1850);
xor U2721 (N_2721,N_1337,N_1424);
xor U2722 (N_2722,N_1866,N_1232);
and U2723 (N_2723,N_1068,N_1075);
nor U2724 (N_2724,N_1061,N_1680);
or U2725 (N_2725,N_1032,N_1981);
nor U2726 (N_2726,N_1313,N_1643);
or U2727 (N_2727,N_1908,N_1333);
nand U2728 (N_2728,N_1024,N_1482);
xor U2729 (N_2729,N_1406,N_1726);
and U2730 (N_2730,N_1858,N_1514);
nor U2731 (N_2731,N_1558,N_1437);
or U2732 (N_2732,N_1120,N_1677);
or U2733 (N_2733,N_1161,N_1542);
nand U2734 (N_2734,N_1206,N_1813);
or U2735 (N_2735,N_1941,N_1595);
xor U2736 (N_2736,N_1985,N_1211);
nand U2737 (N_2737,N_1925,N_1593);
xor U2738 (N_2738,N_1803,N_1952);
nor U2739 (N_2739,N_1621,N_1966);
and U2740 (N_2740,N_1012,N_1405);
or U2741 (N_2741,N_1654,N_1719);
and U2742 (N_2742,N_1704,N_1001);
and U2743 (N_2743,N_1027,N_1551);
and U2744 (N_2744,N_1625,N_1394);
nor U2745 (N_2745,N_1969,N_1570);
or U2746 (N_2746,N_1724,N_1515);
or U2747 (N_2747,N_1600,N_1162);
and U2748 (N_2748,N_1990,N_1895);
nand U2749 (N_2749,N_1223,N_1762);
xor U2750 (N_2750,N_1448,N_1101);
nand U2751 (N_2751,N_1651,N_1772);
xor U2752 (N_2752,N_1748,N_1664);
xor U2753 (N_2753,N_1420,N_1852);
or U2754 (N_2754,N_1637,N_1465);
or U2755 (N_2755,N_1124,N_1140);
xnor U2756 (N_2756,N_1753,N_1977);
xor U2757 (N_2757,N_1604,N_1584);
xnor U2758 (N_2758,N_1537,N_1877);
or U2759 (N_2759,N_1008,N_1132);
and U2760 (N_2760,N_1070,N_1605);
xor U2761 (N_2761,N_1428,N_1478);
nor U2762 (N_2762,N_1884,N_1060);
or U2763 (N_2763,N_1177,N_1842);
nor U2764 (N_2764,N_1075,N_1852);
and U2765 (N_2765,N_1758,N_1611);
xnor U2766 (N_2766,N_1825,N_1794);
nand U2767 (N_2767,N_1214,N_1911);
or U2768 (N_2768,N_1009,N_1660);
or U2769 (N_2769,N_1766,N_1731);
nand U2770 (N_2770,N_1667,N_1473);
and U2771 (N_2771,N_1701,N_1559);
and U2772 (N_2772,N_1566,N_1806);
nor U2773 (N_2773,N_1150,N_1501);
xor U2774 (N_2774,N_1555,N_1338);
or U2775 (N_2775,N_1338,N_1440);
nor U2776 (N_2776,N_1137,N_1861);
xor U2777 (N_2777,N_1643,N_1010);
and U2778 (N_2778,N_1878,N_1143);
xnor U2779 (N_2779,N_1003,N_1567);
nor U2780 (N_2780,N_1904,N_1951);
nand U2781 (N_2781,N_1322,N_1166);
xor U2782 (N_2782,N_1919,N_1720);
xnor U2783 (N_2783,N_1955,N_1719);
nor U2784 (N_2784,N_1679,N_1763);
nand U2785 (N_2785,N_1729,N_1421);
xnor U2786 (N_2786,N_1250,N_1216);
nor U2787 (N_2787,N_1038,N_1890);
nor U2788 (N_2788,N_1890,N_1152);
or U2789 (N_2789,N_1755,N_1214);
nor U2790 (N_2790,N_1530,N_1686);
nor U2791 (N_2791,N_1693,N_1903);
nor U2792 (N_2792,N_1405,N_1424);
xnor U2793 (N_2793,N_1525,N_1289);
nor U2794 (N_2794,N_1496,N_1783);
or U2795 (N_2795,N_1770,N_1754);
nand U2796 (N_2796,N_1452,N_1712);
or U2797 (N_2797,N_1146,N_1803);
xor U2798 (N_2798,N_1477,N_1888);
nor U2799 (N_2799,N_1759,N_1254);
and U2800 (N_2800,N_1537,N_1424);
nand U2801 (N_2801,N_1674,N_1508);
or U2802 (N_2802,N_1240,N_1404);
and U2803 (N_2803,N_1665,N_1713);
nor U2804 (N_2804,N_1768,N_1803);
and U2805 (N_2805,N_1204,N_1604);
or U2806 (N_2806,N_1530,N_1795);
nor U2807 (N_2807,N_1146,N_1008);
or U2808 (N_2808,N_1107,N_1568);
xor U2809 (N_2809,N_1144,N_1105);
nand U2810 (N_2810,N_1404,N_1313);
or U2811 (N_2811,N_1791,N_1337);
nor U2812 (N_2812,N_1229,N_1946);
and U2813 (N_2813,N_1322,N_1474);
xnor U2814 (N_2814,N_1280,N_1084);
xnor U2815 (N_2815,N_1326,N_1162);
xnor U2816 (N_2816,N_1213,N_1007);
or U2817 (N_2817,N_1790,N_1661);
nor U2818 (N_2818,N_1700,N_1035);
xnor U2819 (N_2819,N_1119,N_1197);
and U2820 (N_2820,N_1307,N_1253);
and U2821 (N_2821,N_1042,N_1488);
nor U2822 (N_2822,N_1265,N_1960);
nand U2823 (N_2823,N_1160,N_1587);
or U2824 (N_2824,N_1133,N_1173);
xor U2825 (N_2825,N_1619,N_1602);
nor U2826 (N_2826,N_1361,N_1664);
xor U2827 (N_2827,N_1311,N_1257);
xor U2828 (N_2828,N_1264,N_1306);
nand U2829 (N_2829,N_1015,N_1810);
nor U2830 (N_2830,N_1542,N_1407);
or U2831 (N_2831,N_1681,N_1171);
xnor U2832 (N_2832,N_1767,N_1743);
nand U2833 (N_2833,N_1852,N_1235);
xnor U2834 (N_2834,N_1132,N_1634);
and U2835 (N_2835,N_1006,N_1294);
xor U2836 (N_2836,N_1537,N_1003);
and U2837 (N_2837,N_1578,N_1274);
or U2838 (N_2838,N_1661,N_1769);
nand U2839 (N_2839,N_1672,N_1359);
xor U2840 (N_2840,N_1698,N_1181);
nand U2841 (N_2841,N_1439,N_1856);
nor U2842 (N_2842,N_1086,N_1421);
xnor U2843 (N_2843,N_1671,N_1636);
nor U2844 (N_2844,N_1378,N_1130);
nor U2845 (N_2845,N_1118,N_1799);
and U2846 (N_2846,N_1431,N_1543);
or U2847 (N_2847,N_1132,N_1130);
or U2848 (N_2848,N_1798,N_1608);
nor U2849 (N_2849,N_1462,N_1036);
nand U2850 (N_2850,N_1126,N_1206);
nor U2851 (N_2851,N_1153,N_1150);
and U2852 (N_2852,N_1579,N_1443);
or U2853 (N_2853,N_1925,N_1245);
or U2854 (N_2854,N_1226,N_1235);
nor U2855 (N_2855,N_1511,N_1992);
nand U2856 (N_2856,N_1826,N_1757);
and U2857 (N_2857,N_1578,N_1567);
nor U2858 (N_2858,N_1282,N_1899);
nand U2859 (N_2859,N_1816,N_1550);
nand U2860 (N_2860,N_1166,N_1973);
nor U2861 (N_2861,N_1251,N_1979);
xnor U2862 (N_2862,N_1635,N_1487);
nand U2863 (N_2863,N_1337,N_1959);
or U2864 (N_2864,N_1396,N_1308);
nand U2865 (N_2865,N_1125,N_1849);
xnor U2866 (N_2866,N_1722,N_1620);
xnor U2867 (N_2867,N_1074,N_1912);
nor U2868 (N_2868,N_1390,N_1460);
or U2869 (N_2869,N_1598,N_1594);
xnor U2870 (N_2870,N_1518,N_1047);
xnor U2871 (N_2871,N_1424,N_1705);
nand U2872 (N_2872,N_1158,N_1647);
nor U2873 (N_2873,N_1489,N_1132);
nor U2874 (N_2874,N_1969,N_1517);
and U2875 (N_2875,N_1905,N_1010);
xor U2876 (N_2876,N_1216,N_1493);
nand U2877 (N_2877,N_1129,N_1899);
and U2878 (N_2878,N_1025,N_1936);
nand U2879 (N_2879,N_1868,N_1226);
nor U2880 (N_2880,N_1257,N_1084);
or U2881 (N_2881,N_1751,N_1868);
nand U2882 (N_2882,N_1863,N_1808);
nor U2883 (N_2883,N_1015,N_1869);
xor U2884 (N_2884,N_1064,N_1198);
nor U2885 (N_2885,N_1635,N_1693);
nor U2886 (N_2886,N_1850,N_1031);
or U2887 (N_2887,N_1956,N_1734);
and U2888 (N_2888,N_1631,N_1346);
xnor U2889 (N_2889,N_1595,N_1421);
and U2890 (N_2890,N_1690,N_1403);
or U2891 (N_2891,N_1526,N_1907);
and U2892 (N_2892,N_1484,N_1782);
or U2893 (N_2893,N_1902,N_1788);
or U2894 (N_2894,N_1900,N_1612);
xnor U2895 (N_2895,N_1303,N_1985);
nand U2896 (N_2896,N_1888,N_1884);
nand U2897 (N_2897,N_1511,N_1163);
nor U2898 (N_2898,N_1499,N_1292);
xnor U2899 (N_2899,N_1026,N_1204);
nand U2900 (N_2900,N_1423,N_1394);
and U2901 (N_2901,N_1525,N_1687);
xor U2902 (N_2902,N_1521,N_1129);
nor U2903 (N_2903,N_1932,N_1258);
nand U2904 (N_2904,N_1352,N_1887);
nand U2905 (N_2905,N_1179,N_1900);
xor U2906 (N_2906,N_1151,N_1530);
nor U2907 (N_2907,N_1482,N_1249);
nor U2908 (N_2908,N_1099,N_1947);
xor U2909 (N_2909,N_1397,N_1247);
nand U2910 (N_2910,N_1033,N_1945);
xnor U2911 (N_2911,N_1741,N_1626);
nor U2912 (N_2912,N_1703,N_1261);
and U2913 (N_2913,N_1502,N_1004);
nor U2914 (N_2914,N_1257,N_1871);
nor U2915 (N_2915,N_1630,N_1957);
nor U2916 (N_2916,N_1638,N_1190);
and U2917 (N_2917,N_1733,N_1989);
nand U2918 (N_2918,N_1481,N_1524);
nand U2919 (N_2919,N_1968,N_1098);
and U2920 (N_2920,N_1337,N_1541);
and U2921 (N_2921,N_1383,N_1931);
xor U2922 (N_2922,N_1452,N_1180);
and U2923 (N_2923,N_1916,N_1761);
nand U2924 (N_2924,N_1898,N_1120);
or U2925 (N_2925,N_1213,N_1771);
xnor U2926 (N_2926,N_1101,N_1525);
or U2927 (N_2927,N_1810,N_1178);
nor U2928 (N_2928,N_1963,N_1019);
nor U2929 (N_2929,N_1494,N_1895);
nor U2930 (N_2930,N_1507,N_1904);
or U2931 (N_2931,N_1868,N_1355);
xnor U2932 (N_2932,N_1733,N_1553);
nand U2933 (N_2933,N_1546,N_1203);
nand U2934 (N_2934,N_1876,N_1815);
nand U2935 (N_2935,N_1960,N_1388);
nor U2936 (N_2936,N_1141,N_1715);
xor U2937 (N_2937,N_1302,N_1888);
nor U2938 (N_2938,N_1551,N_1538);
and U2939 (N_2939,N_1080,N_1202);
xor U2940 (N_2940,N_1487,N_1341);
nor U2941 (N_2941,N_1611,N_1502);
and U2942 (N_2942,N_1157,N_1651);
or U2943 (N_2943,N_1186,N_1708);
xor U2944 (N_2944,N_1132,N_1837);
or U2945 (N_2945,N_1987,N_1719);
nand U2946 (N_2946,N_1071,N_1042);
nand U2947 (N_2947,N_1205,N_1360);
and U2948 (N_2948,N_1458,N_1753);
and U2949 (N_2949,N_1727,N_1543);
and U2950 (N_2950,N_1374,N_1618);
xnor U2951 (N_2951,N_1525,N_1419);
and U2952 (N_2952,N_1105,N_1535);
xor U2953 (N_2953,N_1964,N_1633);
or U2954 (N_2954,N_1585,N_1875);
nand U2955 (N_2955,N_1655,N_1762);
nor U2956 (N_2956,N_1621,N_1201);
and U2957 (N_2957,N_1208,N_1899);
xnor U2958 (N_2958,N_1073,N_1789);
xnor U2959 (N_2959,N_1551,N_1387);
nor U2960 (N_2960,N_1412,N_1285);
and U2961 (N_2961,N_1677,N_1002);
nor U2962 (N_2962,N_1597,N_1249);
xnor U2963 (N_2963,N_1701,N_1299);
and U2964 (N_2964,N_1411,N_1877);
and U2965 (N_2965,N_1620,N_1823);
nand U2966 (N_2966,N_1349,N_1825);
nand U2967 (N_2967,N_1610,N_1002);
nand U2968 (N_2968,N_1404,N_1560);
xor U2969 (N_2969,N_1843,N_1424);
nor U2970 (N_2970,N_1767,N_1783);
xor U2971 (N_2971,N_1241,N_1084);
or U2972 (N_2972,N_1324,N_1305);
xnor U2973 (N_2973,N_1649,N_1029);
or U2974 (N_2974,N_1022,N_1211);
xor U2975 (N_2975,N_1091,N_1932);
xor U2976 (N_2976,N_1547,N_1151);
and U2977 (N_2977,N_1311,N_1046);
nand U2978 (N_2978,N_1588,N_1298);
or U2979 (N_2979,N_1138,N_1999);
nand U2980 (N_2980,N_1560,N_1593);
nor U2981 (N_2981,N_1348,N_1651);
or U2982 (N_2982,N_1741,N_1270);
and U2983 (N_2983,N_1558,N_1609);
nor U2984 (N_2984,N_1603,N_1359);
nand U2985 (N_2985,N_1056,N_1042);
or U2986 (N_2986,N_1598,N_1453);
nor U2987 (N_2987,N_1180,N_1466);
or U2988 (N_2988,N_1269,N_1421);
nor U2989 (N_2989,N_1707,N_1419);
xnor U2990 (N_2990,N_1344,N_1015);
and U2991 (N_2991,N_1394,N_1603);
nand U2992 (N_2992,N_1535,N_1610);
xor U2993 (N_2993,N_1673,N_1427);
and U2994 (N_2994,N_1137,N_1406);
nor U2995 (N_2995,N_1790,N_1276);
nand U2996 (N_2996,N_1808,N_1914);
nor U2997 (N_2997,N_1214,N_1793);
and U2998 (N_2998,N_1304,N_1121);
nand U2999 (N_2999,N_1220,N_1668);
or U3000 (N_3000,N_2132,N_2504);
nand U3001 (N_3001,N_2452,N_2774);
nand U3002 (N_3002,N_2742,N_2749);
and U3003 (N_3003,N_2770,N_2645);
xor U3004 (N_3004,N_2884,N_2978);
or U3005 (N_3005,N_2034,N_2004);
nand U3006 (N_3006,N_2793,N_2913);
and U3007 (N_3007,N_2574,N_2692);
xor U3008 (N_3008,N_2607,N_2276);
xor U3009 (N_3009,N_2135,N_2334);
nand U3010 (N_3010,N_2141,N_2703);
xor U3011 (N_3011,N_2191,N_2327);
nor U3012 (N_3012,N_2182,N_2260);
xnor U3013 (N_3013,N_2393,N_2031);
nor U3014 (N_3014,N_2454,N_2128);
or U3015 (N_3015,N_2652,N_2587);
xnor U3016 (N_3016,N_2596,N_2012);
nor U3017 (N_3017,N_2569,N_2251);
xor U3018 (N_3018,N_2522,N_2874);
xnor U3019 (N_3019,N_2972,N_2778);
or U3020 (N_3020,N_2529,N_2390);
or U3021 (N_3021,N_2910,N_2151);
xor U3022 (N_3022,N_2642,N_2268);
nor U3023 (N_3023,N_2581,N_2729);
nand U3024 (N_3024,N_2253,N_2954);
nand U3025 (N_3025,N_2612,N_2364);
nand U3026 (N_3026,N_2624,N_2289);
nand U3027 (N_3027,N_2506,N_2285);
and U3028 (N_3028,N_2055,N_2365);
nor U3029 (N_3029,N_2863,N_2834);
and U3030 (N_3030,N_2472,N_2675);
xor U3031 (N_3031,N_2678,N_2809);
or U3032 (N_3032,N_2585,N_2259);
xnor U3033 (N_3033,N_2228,N_2795);
nor U3034 (N_3034,N_2730,N_2707);
nand U3035 (N_3035,N_2881,N_2629);
and U3036 (N_3036,N_2027,N_2265);
nor U3037 (N_3037,N_2616,N_2889);
nor U3038 (N_3038,N_2469,N_2628);
nor U3039 (N_3039,N_2308,N_2747);
nand U3040 (N_3040,N_2048,N_2483);
nor U3041 (N_3041,N_2754,N_2174);
nor U3042 (N_3042,N_2420,N_2914);
nor U3043 (N_3043,N_2131,N_2006);
and U3044 (N_3044,N_2557,N_2467);
and U3045 (N_3045,N_2150,N_2275);
xnor U3046 (N_3046,N_2019,N_2744);
or U3047 (N_3047,N_2377,N_2400);
nor U3048 (N_3048,N_2800,N_2716);
nor U3049 (N_3049,N_2503,N_2891);
or U3050 (N_3050,N_2931,N_2790);
nand U3051 (N_3051,N_2297,N_2223);
nand U3052 (N_3052,N_2201,N_2161);
or U3053 (N_3053,N_2808,N_2571);
nand U3054 (N_3054,N_2429,N_2110);
nor U3055 (N_3055,N_2180,N_2382);
and U3056 (N_3056,N_2448,N_2944);
or U3057 (N_3057,N_2195,N_2908);
nor U3058 (N_3058,N_2833,N_2821);
or U3059 (N_3059,N_2030,N_2368);
or U3060 (N_3060,N_2967,N_2722);
and U3061 (N_3061,N_2178,N_2915);
or U3062 (N_3062,N_2058,N_2855);
xnor U3063 (N_3063,N_2322,N_2745);
nor U3064 (N_3064,N_2138,N_2667);
xnor U3065 (N_3065,N_2041,N_2426);
and U3066 (N_3066,N_2613,N_2005);
and U3067 (N_3067,N_2816,N_2782);
or U3068 (N_3068,N_2969,N_2530);
and U3069 (N_3069,N_2282,N_2639);
xor U3070 (N_3070,N_2611,N_2388);
and U3071 (N_3071,N_2872,N_2278);
xnor U3072 (N_3072,N_2220,N_2057);
and U3073 (N_3073,N_2591,N_2066);
xnor U3074 (N_3074,N_2568,N_2051);
or U3075 (N_3075,N_2542,N_2803);
nor U3076 (N_3076,N_2122,N_2828);
or U3077 (N_3077,N_2362,N_2428);
or U3078 (N_3078,N_2453,N_2636);
xnor U3079 (N_3079,N_2622,N_2398);
xnor U3080 (N_3080,N_2167,N_2498);
nand U3081 (N_3081,N_2290,N_2149);
xnor U3082 (N_3082,N_2423,N_2419);
and U3083 (N_3083,N_2996,N_2570);
xor U3084 (N_3084,N_2521,N_2080);
nor U3085 (N_3085,N_2214,N_2394);
nor U3086 (N_3086,N_2438,N_2170);
nand U3087 (N_3087,N_2105,N_2540);
xor U3088 (N_3088,N_2020,N_2450);
and U3089 (N_3089,N_2553,N_2734);
nor U3090 (N_3090,N_2205,N_2474);
nor U3091 (N_3091,N_2113,N_2852);
nand U3092 (N_3092,N_2162,N_2582);
and U3093 (N_3093,N_2086,N_2430);
or U3094 (N_3094,N_2077,N_2475);
nand U3095 (N_3095,N_2664,N_2039);
nand U3096 (N_3096,N_2177,N_2898);
nand U3097 (N_3097,N_2072,N_2208);
nor U3098 (N_3098,N_2378,N_2273);
xnor U3099 (N_3099,N_2641,N_2185);
or U3100 (N_3100,N_2106,N_2773);
xor U3101 (N_3101,N_2402,N_2488);
and U3102 (N_3102,N_2603,N_2391);
nand U3103 (N_3103,N_2695,N_2785);
nor U3104 (N_3104,N_2319,N_2901);
xor U3105 (N_3105,N_2239,N_2335);
xnor U3106 (N_3106,N_2490,N_2941);
nand U3107 (N_3107,N_2753,N_2231);
xor U3108 (N_3108,N_2776,N_2865);
and U3109 (N_3109,N_2791,N_2410);
nand U3110 (N_3110,N_2395,N_2010);
nand U3111 (N_3111,N_2731,N_2196);
or U3112 (N_3112,N_2594,N_2677);
and U3113 (N_3113,N_2092,N_2932);
or U3114 (N_3114,N_2071,N_2534);
and U3115 (N_3115,N_2123,N_2281);
or U3116 (N_3116,N_2623,N_2213);
or U3117 (N_3117,N_2366,N_2272);
xnor U3118 (N_3118,N_2054,N_2445);
or U3119 (N_3119,N_2826,N_2310);
nand U3120 (N_3120,N_2087,N_2741);
nand U3121 (N_3121,N_2997,N_2274);
nand U3122 (N_3122,N_2358,N_2599);
or U3123 (N_3123,N_2818,N_2606);
nand U3124 (N_3124,N_2447,N_2882);
nand U3125 (N_3125,N_2936,N_2985);
nand U3126 (N_3126,N_2783,N_2421);
nor U3127 (N_3127,N_2680,N_2073);
nand U3128 (N_3128,N_2644,N_2844);
or U3129 (N_3129,N_2805,N_2084);
and U3130 (N_3130,N_2346,N_2560);
xnor U3131 (N_3131,N_2902,N_2397);
or U3132 (N_3132,N_2219,N_2948);
and U3133 (N_3133,N_2441,N_2842);
nand U3134 (N_3134,N_2971,N_2524);
or U3135 (N_3135,N_2576,N_2189);
nor U3136 (N_3136,N_2924,N_2956);
and U3137 (N_3137,N_2942,N_2115);
or U3138 (N_3138,N_2008,N_2876);
nand U3139 (N_3139,N_2082,N_2089);
xor U3140 (N_3140,N_2526,N_2212);
and U3141 (N_3141,N_2171,N_2871);
nor U3142 (N_3142,N_2246,N_2563);
xor U3143 (N_3143,N_2837,N_2090);
and U3144 (N_3144,N_2007,N_2751);
nor U3145 (N_3145,N_2977,N_2512);
nor U3146 (N_3146,N_2919,N_2333);
nand U3147 (N_3147,N_2799,N_2342);
xnor U3148 (N_3148,N_2381,N_2687);
or U3149 (N_3149,N_2555,N_2721);
and U3150 (N_3150,N_2098,N_2849);
or U3151 (N_3151,N_2957,N_2864);
xnor U3152 (N_3152,N_2466,N_2166);
and U3153 (N_3153,N_2422,N_2187);
nor U3154 (N_3154,N_2806,N_2893);
xnor U3155 (N_3155,N_2029,N_2050);
or U3156 (N_3156,N_2096,N_2955);
xor U3157 (N_3157,N_2302,N_2037);
nor U3158 (N_3158,N_2094,N_2032);
or U3159 (N_3159,N_2065,N_2810);
nor U3160 (N_3160,N_2271,N_2341);
xor U3161 (N_3161,N_2789,N_2159);
nor U3162 (N_3162,N_2222,N_2655);
nor U3163 (N_3163,N_2857,N_2701);
nor U3164 (N_3164,N_2277,N_2895);
nand U3165 (N_3165,N_2356,N_2286);
xor U3166 (N_3166,N_2224,N_2234);
nand U3167 (N_3167,N_2750,N_2387);
and U3168 (N_3168,N_2817,N_2074);
nor U3169 (N_3169,N_2492,N_2173);
nor U3170 (N_3170,N_2543,N_2998);
xor U3171 (N_3171,N_2043,N_2210);
nor U3172 (N_3172,N_2939,N_2482);
or U3173 (N_3173,N_2497,N_2653);
or U3174 (N_3174,N_2347,N_2249);
or U3175 (N_3175,N_2349,N_2245);
nand U3176 (N_3176,N_2413,N_2651);
and U3177 (N_3177,N_2489,N_2772);
xor U3178 (N_3178,N_2904,N_2179);
or U3179 (N_3179,N_2888,N_2003);
nand U3180 (N_3180,N_2233,N_2781);
nor U3181 (N_3181,N_2705,N_2883);
xnor U3182 (N_3182,N_2737,N_2207);
or U3183 (N_3183,N_2539,N_2965);
nor U3184 (N_3184,N_2983,N_2614);
nand U3185 (N_3185,N_2892,N_2843);
nor U3186 (N_3186,N_2520,N_2432);
nand U3187 (N_3187,N_2476,N_2330);
or U3188 (N_3188,N_2313,N_2134);
nor U3189 (N_3189,N_2403,N_2236);
and U3190 (N_3190,N_2494,N_2684);
nor U3191 (N_3191,N_2221,N_2683);
nand U3192 (N_3192,N_2145,N_2647);
nor U3193 (N_3193,N_2460,N_2862);
xnor U3194 (N_3194,N_2363,N_2093);
xor U3195 (N_3195,N_2300,N_2414);
nor U3196 (N_3196,N_2181,N_2155);
or U3197 (N_3197,N_2981,N_2657);
or U3198 (N_3198,N_2905,N_2242);
nor U3199 (N_3199,N_2456,N_2798);
xor U3200 (N_3200,N_2124,N_2121);
xnor U3201 (N_3201,N_2449,N_2505);
and U3202 (N_3202,N_2694,N_2348);
and U3203 (N_3203,N_2112,N_2192);
and U3204 (N_3204,N_2411,N_2148);
nor U3205 (N_3205,N_2235,N_2127);
and U3206 (N_3206,N_2633,N_2225);
or U3207 (N_3207,N_2600,N_2825);
nor U3208 (N_3208,N_2867,N_2117);
nor U3209 (N_3209,N_2375,N_2940);
xor U3210 (N_3210,N_2909,N_2620);
nand U3211 (N_3211,N_2823,N_2764);
or U3212 (N_3212,N_2704,N_2357);
xnor U3213 (N_3213,N_2204,N_2696);
or U3214 (N_3214,N_2929,N_2401);
xor U3215 (N_3215,N_2514,N_2784);
or U3216 (N_3216,N_2672,N_2922);
xor U3217 (N_3217,N_2943,N_2464);
nand U3218 (N_3218,N_2194,N_2009);
xor U3219 (N_3219,N_2021,N_2994);
nand U3220 (N_3220,N_2176,N_2638);
nor U3221 (N_3221,N_2011,N_2339);
nor U3222 (N_3222,N_2495,N_2075);
nor U3223 (N_3223,N_2232,N_2602);
xor U3224 (N_3224,N_2693,N_2937);
nand U3225 (N_3225,N_2987,N_2318);
or U3226 (N_3226,N_2735,N_2136);
nor U3227 (N_3227,N_2711,N_2169);
nand U3228 (N_3228,N_2851,N_2934);
nor U3229 (N_3229,N_2928,N_2760);
or U3230 (N_3230,N_2739,N_2984);
xor U3231 (N_3231,N_2437,N_2714);
xor U3232 (N_3232,N_2118,N_2590);
nand U3233 (N_3233,N_2518,N_2355);
or U3234 (N_3234,N_2293,N_2650);
and U3235 (N_3235,N_2493,N_2689);
nor U3236 (N_3236,N_2660,N_2314);
xnor U3237 (N_3237,N_2218,N_2091);
nand U3238 (N_3238,N_2970,N_2921);
or U3239 (N_3239,N_2879,N_2758);
or U3240 (N_3240,N_2897,N_2042);
and U3241 (N_3241,N_2966,N_2140);
and U3242 (N_3242,N_2211,N_2299);
xnor U3243 (N_3243,N_2431,N_2632);
nor U3244 (N_3244,N_2510,N_2200);
xor U3245 (N_3245,N_2160,N_2325);
nor U3246 (N_3246,N_2605,N_2545);
nor U3247 (N_3247,N_2583,N_2918);
or U3248 (N_3248,N_2811,N_2724);
or U3249 (N_3249,N_2875,N_2107);
or U3250 (N_3250,N_2045,N_2307);
and U3251 (N_3251,N_2827,N_2700);
and U3252 (N_3252,N_2960,N_2238);
and U3253 (N_3253,N_2787,N_2685);
nand U3254 (N_3254,N_2499,N_2873);
and U3255 (N_3255,N_2777,N_2755);
nand U3256 (N_3256,N_2559,N_2748);
xor U3257 (N_3257,N_2911,N_2535);
and U3258 (N_3258,N_2095,N_2324);
and U3259 (N_3259,N_2573,N_2321);
and U3260 (N_3260,N_2417,N_2354);
nor U3261 (N_3261,N_2199,N_2163);
or U3262 (N_3262,N_2820,N_2968);
or U3263 (N_3263,N_2501,N_2567);
or U3264 (N_3264,N_2193,N_2989);
nand U3265 (N_3265,N_2933,N_2230);
xnor U3266 (N_3266,N_2668,N_2125);
nor U3267 (N_3267,N_2598,N_2103);
xor U3268 (N_3268,N_2725,N_2993);
nor U3269 (N_3269,N_2838,N_2627);
xnor U3270 (N_3270,N_2283,N_2457);
nand U3271 (N_3271,N_2593,N_2718);
or U3272 (N_3272,N_2076,N_2126);
or U3273 (N_3273,N_2771,N_2938);
nand U3274 (N_3274,N_2081,N_2059);
nor U3275 (N_3275,N_2443,N_2544);
and U3276 (N_3276,N_2070,N_2502);
nand U3277 (N_3277,N_2309,N_2509);
or U3278 (N_3278,N_2405,N_2579);
nand U3279 (N_3279,N_2369,N_2184);
or U3280 (N_3280,N_2002,N_2669);
or U3281 (N_3281,N_2486,N_2962);
or U3282 (N_3282,N_2990,N_2562);
and U3283 (N_3283,N_2247,N_2709);
or U3284 (N_3284,N_2830,N_2255);
or U3285 (N_3285,N_2374,N_2508);
nor U3286 (N_3286,N_2014,N_2604);
nand U3287 (N_3287,N_2847,N_2699);
nor U3288 (N_3288,N_2434,N_2815);
or U3289 (N_3289,N_2404,N_2547);
nand U3290 (N_3290,N_2767,N_2440);
or U3291 (N_3291,N_2532,N_2640);
xnor U3292 (N_3292,N_2757,N_2017);
or U3293 (N_3293,N_2515,N_2558);
nand U3294 (N_3294,N_2244,N_2676);
or U3295 (N_3295,N_2491,N_2780);
xor U3296 (N_3296,N_2878,N_2360);
or U3297 (N_3297,N_2198,N_2974);
or U3298 (N_3298,N_2999,N_2415);
and U3299 (N_3299,N_2992,N_2241);
or U3300 (N_3300,N_2619,N_2144);
and U3301 (N_3301,N_2101,N_2258);
nand U3302 (N_3302,N_2868,N_2018);
or U3303 (N_3303,N_2775,N_2370);
xor U3304 (N_3304,N_2083,N_2697);
or U3305 (N_3305,N_2100,N_2439);
nor U3306 (N_3306,N_2756,N_2950);
and U3307 (N_3307,N_2061,N_2485);
and U3308 (N_3308,N_2550,N_2295);
and U3309 (N_3309,N_2446,N_2848);
or U3310 (N_3310,N_2723,N_2040);
xor U3311 (N_3311,N_2383,N_2407);
or U3312 (N_3312,N_2761,N_2986);
and U3313 (N_3313,N_2461,N_2656);
nor U3314 (N_3314,N_2496,N_2713);
nor U3315 (N_3315,N_2001,N_2738);
nand U3316 (N_3316,N_2376,N_2399);
xor U3317 (N_3317,N_2870,N_2715);
nor U3318 (N_3318,N_2326,N_2609);
nor U3319 (N_3319,N_2779,N_2952);
xor U3320 (N_3320,N_2597,N_2462);
or U3321 (N_3321,N_2511,N_2786);
or U3322 (N_3322,N_2280,N_2353);
xor U3323 (N_3323,N_2287,N_2079);
or U3324 (N_3324,N_2643,N_2266);
nor U3325 (N_3325,N_2953,N_2133);
xor U3326 (N_3326,N_2886,N_2740);
xor U3327 (N_3327,N_2478,N_2566);
and U3328 (N_3328,N_2424,N_2256);
xnor U3329 (N_3329,N_2473,N_2154);
or U3330 (N_3330,N_2719,N_2139);
or U3331 (N_3331,N_2267,N_2637);
nor U3332 (N_3332,N_2618,N_2853);
xnor U3333 (N_3333,N_2792,N_2099);
and U3334 (N_3334,N_2682,N_2991);
or U3335 (N_3335,N_2537,N_2608);
and U3336 (N_3336,N_2046,N_2052);
xor U3337 (N_3337,N_2209,N_2869);
and U3338 (N_3338,N_2379,N_2964);
nand U3339 (N_3339,N_2935,N_2727);
and U3340 (N_3340,N_2726,N_2056);
or U3341 (N_3341,N_2328,N_2690);
nand U3342 (N_3342,N_2028,N_2038);
xor U3343 (N_3343,N_2890,N_2471);
nand U3344 (N_3344,N_2575,N_2912);
nor U3345 (N_3345,N_2016,N_2049);
xor U3346 (N_3346,N_2044,N_2930);
xor U3347 (N_3347,N_2634,N_2681);
xnor U3348 (N_3348,N_2958,N_2973);
nand U3349 (N_3349,N_2345,N_2728);
and U3350 (N_3350,N_2085,N_2708);
or U3351 (N_3351,N_2227,N_2367);
nor U3352 (N_3352,N_2769,N_2666);
or U3353 (N_3353,N_2114,N_2832);
xor U3354 (N_3354,N_2361,N_2250);
xor U3355 (N_3355,N_2329,N_2949);
xnor U3356 (N_3356,N_2311,N_2860);
and U3357 (N_3357,N_2617,N_2768);
nand U3358 (N_3358,N_2269,N_2903);
and U3359 (N_3359,N_2648,N_2317);
or U3360 (N_3360,N_2839,N_2679);
and U3361 (N_3361,N_2976,N_2854);
nor U3362 (N_3362,N_2262,N_2572);
nand U3363 (N_3363,N_2923,N_2487);
and U3364 (N_3364,N_2023,N_2392);
nand U3365 (N_3365,N_2752,N_2175);
nand U3366 (N_3366,N_2635,N_2665);
or U3367 (N_3367,N_2000,N_2925);
xor U3368 (N_3368,N_2945,N_2386);
nand U3369 (N_3369,N_2384,N_2845);
nand U3370 (N_3370,N_2859,N_2894);
or U3371 (N_3371,N_2344,N_2906);
xnor U3372 (N_3372,N_2822,N_2243);
nor U3373 (N_3373,N_2546,N_2097);
nand U3374 (N_3374,N_2146,N_2663);
nand U3375 (N_3375,N_2481,N_2433);
xor U3376 (N_3376,N_2470,N_2900);
xor U3377 (N_3377,N_2759,N_2961);
or U3378 (N_3378,N_2720,N_2920);
or U3379 (N_3379,N_2408,N_2406);
nand U3380 (N_3380,N_2197,N_2359);
xnor U3381 (N_3381,N_2766,N_2418);
and U3382 (N_3382,N_2584,N_2024);
and U3383 (N_3383,N_2458,N_2531);
nor U3384 (N_3384,N_2129,N_2158);
and U3385 (N_3385,N_2896,N_2371);
xnor U3386 (N_3386,N_2631,N_2240);
nor U3387 (N_3387,N_2698,N_2588);
xor U3388 (N_3388,N_2980,N_2975);
and U3389 (N_3389,N_2229,N_2202);
or U3390 (N_3390,N_2063,N_2168);
xor U3391 (N_3391,N_2257,N_2717);
nand U3392 (N_3392,N_2686,N_2802);
nor U3393 (N_3393,N_2765,N_2654);
or U3394 (N_3394,N_2601,N_2336);
nand U3395 (N_3395,N_2551,N_2533);
nor U3396 (N_3396,N_2813,N_2270);
and U3397 (N_3397,N_2047,N_2477);
or U3398 (N_3398,N_2812,N_2840);
nor U3399 (N_3399,N_2069,N_2068);
xnor U3400 (N_3400,N_2885,N_2248);
xnor U3401 (N_3401,N_2733,N_2111);
nand U3402 (N_3402,N_2856,N_2416);
and U3403 (N_3403,N_2465,N_2157);
xnor U3404 (N_3404,N_2804,N_2442);
or U3405 (N_3405,N_2331,N_2078);
nor U3406 (N_3406,N_2396,N_2525);
or U3407 (N_3407,N_2261,N_2165);
xor U3408 (N_3408,N_2507,N_2523);
or U3409 (N_3409,N_2385,N_2025);
nand U3410 (N_3410,N_2022,N_2142);
xor U3411 (N_3411,N_2702,N_2190);
xnor U3412 (N_3412,N_2062,N_2305);
or U3413 (N_3413,N_2425,N_2389);
or U3414 (N_3414,N_2484,N_2147);
xnor U3415 (N_3415,N_2254,N_2796);
nand U3416 (N_3416,N_2186,N_2116);
xor U3417 (N_3417,N_2807,N_2444);
and U3418 (N_3418,N_2982,N_2380);
and U3419 (N_3419,N_2671,N_2836);
nand U3420 (N_3420,N_2516,N_2252);
or U3421 (N_3421,N_2762,N_2829);
nand U3422 (N_3422,N_2203,N_2578);
or U3423 (N_3423,N_2794,N_2427);
xor U3424 (N_3424,N_2947,N_2564);
or U3425 (N_3425,N_2661,N_2053);
nor U3426 (N_3426,N_2372,N_2625);
and U3427 (N_3427,N_2797,N_2988);
or U3428 (N_3428,N_2130,N_2877);
nand U3429 (N_3429,N_2549,N_2188);
and U3430 (N_3430,N_2951,N_2670);
and U3431 (N_3431,N_2435,N_2412);
xnor U3432 (N_3432,N_2480,N_2340);
or U3433 (N_3433,N_2035,N_2292);
and U3434 (N_3434,N_2580,N_2338);
and U3435 (N_3435,N_2519,N_2887);
nand U3436 (N_3436,N_2291,N_2217);
nand U3437 (N_3437,N_2926,N_2284);
nand U3438 (N_3438,N_2527,N_2301);
nor U3439 (N_3439,N_2541,N_2710);
or U3440 (N_3440,N_2343,N_2835);
xnor U3441 (N_3441,N_2263,N_2577);
xnor U3442 (N_3442,N_2658,N_2064);
nand U3443 (N_3443,N_2468,N_2850);
xnor U3444 (N_3444,N_2436,N_2517);
and U3445 (N_3445,N_2528,N_2088);
and U3446 (N_3446,N_2621,N_2659);
or U3447 (N_3447,N_2538,N_2109);
nor U3448 (N_3448,N_2674,N_2595);
xnor U3449 (N_3449,N_2688,N_2556);
and U3450 (N_3450,N_2673,N_2033);
nand U3451 (N_3451,N_2552,N_2662);
and U3452 (N_3452,N_2409,N_2226);
xnor U3453 (N_3453,N_2959,N_2108);
nor U3454 (N_3454,N_2036,N_2646);
and U3455 (N_3455,N_2104,N_2626);
nor U3456 (N_3456,N_2801,N_2479);
and U3457 (N_3457,N_2963,N_2015);
nor U3458 (N_3458,N_2536,N_2592);
nor U3459 (N_3459,N_2630,N_2706);
nand U3460 (N_3460,N_2119,N_2164);
and U3461 (N_3461,N_2907,N_2548);
nand U3462 (N_3462,N_2067,N_2831);
and U3463 (N_3463,N_2819,N_2183);
nand U3464 (N_3464,N_2026,N_2060);
nor U3465 (N_3465,N_2712,N_2846);
xnor U3466 (N_3466,N_2264,N_2215);
and U3467 (N_3467,N_2102,N_2298);
xor U3468 (N_3468,N_2373,N_2861);
and U3469 (N_3469,N_2736,N_2615);
xor U3470 (N_3470,N_2320,N_2927);
xor U3471 (N_3471,N_2788,N_2206);
nand U3472 (N_3472,N_2610,N_2814);
nand U3473 (N_3473,N_2316,N_2216);
nor U3474 (N_3474,N_2120,N_2352);
xnor U3475 (N_3475,N_2153,N_2979);
xor U3476 (N_3476,N_2294,N_2137);
xor U3477 (N_3477,N_2451,N_2732);
and U3478 (N_3478,N_2312,N_2306);
nor U3479 (N_3479,N_2279,N_2500);
or U3480 (N_3480,N_2691,N_2143);
nand U3481 (N_3481,N_2995,N_2323);
and U3482 (N_3482,N_2296,N_2351);
or U3483 (N_3483,N_2237,N_2589);
xor U3484 (N_3484,N_2586,N_2916);
or U3485 (N_3485,N_2350,N_2332);
and U3486 (N_3486,N_2172,N_2866);
nand U3487 (N_3487,N_2763,N_2463);
xor U3488 (N_3488,N_2315,N_2152);
nor U3489 (N_3489,N_2858,N_2561);
xnor U3490 (N_3490,N_2565,N_2013);
nor U3491 (N_3491,N_2880,N_2917);
xnor U3492 (N_3492,N_2455,N_2899);
or U3493 (N_3493,N_2288,N_2459);
nor U3494 (N_3494,N_2946,N_2303);
or U3495 (N_3495,N_2513,N_2743);
nand U3496 (N_3496,N_2841,N_2337);
nor U3497 (N_3497,N_2746,N_2156);
or U3498 (N_3498,N_2304,N_2649);
and U3499 (N_3499,N_2824,N_2554);
or U3500 (N_3500,N_2773,N_2763);
xnor U3501 (N_3501,N_2467,N_2679);
nand U3502 (N_3502,N_2782,N_2705);
xnor U3503 (N_3503,N_2795,N_2403);
and U3504 (N_3504,N_2697,N_2196);
nand U3505 (N_3505,N_2940,N_2641);
and U3506 (N_3506,N_2011,N_2899);
or U3507 (N_3507,N_2966,N_2251);
or U3508 (N_3508,N_2333,N_2426);
nor U3509 (N_3509,N_2246,N_2904);
xnor U3510 (N_3510,N_2734,N_2995);
and U3511 (N_3511,N_2032,N_2492);
and U3512 (N_3512,N_2401,N_2264);
or U3513 (N_3513,N_2036,N_2517);
nor U3514 (N_3514,N_2350,N_2314);
nor U3515 (N_3515,N_2014,N_2934);
nor U3516 (N_3516,N_2711,N_2904);
xor U3517 (N_3517,N_2240,N_2148);
or U3518 (N_3518,N_2678,N_2252);
nor U3519 (N_3519,N_2051,N_2902);
nor U3520 (N_3520,N_2360,N_2106);
xnor U3521 (N_3521,N_2711,N_2887);
nor U3522 (N_3522,N_2507,N_2353);
xnor U3523 (N_3523,N_2040,N_2511);
xnor U3524 (N_3524,N_2344,N_2572);
nand U3525 (N_3525,N_2132,N_2821);
nand U3526 (N_3526,N_2005,N_2768);
nor U3527 (N_3527,N_2305,N_2399);
nand U3528 (N_3528,N_2353,N_2899);
or U3529 (N_3529,N_2680,N_2100);
xnor U3530 (N_3530,N_2031,N_2740);
nand U3531 (N_3531,N_2275,N_2544);
nand U3532 (N_3532,N_2797,N_2927);
nand U3533 (N_3533,N_2195,N_2565);
and U3534 (N_3534,N_2681,N_2353);
or U3535 (N_3535,N_2594,N_2457);
xnor U3536 (N_3536,N_2601,N_2054);
or U3537 (N_3537,N_2469,N_2093);
xnor U3538 (N_3538,N_2490,N_2225);
nand U3539 (N_3539,N_2072,N_2804);
xor U3540 (N_3540,N_2708,N_2842);
nor U3541 (N_3541,N_2761,N_2714);
xor U3542 (N_3542,N_2503,N_2210);
or U3543 (N_3543,N_2681,N_2770);
nor U3544 (N_3544,N_2847,N_2921);
nor U3545 (N_3545,N_2009,N_2827);
or U3546 (N_3546,N_2992,N_2972);
nand U3547 (N_3547,N_2704,N_2766);
and U3548 (N_3548,N_2700,N_2841);
xor U3549 (N_3549,N_2858,N_2376);
or U3550 (N_3550,N_2838,N_2292);
nor U3551 (N_3551,N_2281,N_2249);
and U3552 (N_3552,N_2639,N_2989);
nor U3553 (N_3553,N_2773,N_2313);
or U3554 (N_3554,N_2888,N_2593);
nand U3555 (N_3555,N_2235,N_2012);
and U3556 (N_3556,N_2609,N_2526);
and U3557 (N_3557,N_2217,N_2352);
nor U3558 (N_3558,N_2757,N_2177);
or U3559 (N_3559,N_2521,N_2005);
and U3560 (N_3560,N_2188,N_2520);
xor U3561 (N_3561,N_2022,N_2224);
nand U3562 (N_3562,N_2702,N_2544);
nand U3563 (N_3563,N_2737,N_2875);
or U3564 (N_3564,N_2680,N_2582);
and U3565 (N_3565,N_2430,N_2571);
or U3566 (N_3566,N_2695,N_2184);
nand U3567 (N_3567,N_2884,N_2223);
or U3568 (N_3568,N_2547,N_2417);
nand U3569 (N_3569,N_2655,N_2154);
and U3570 (N_3570,N_2208,N_2657);
and U3571 (N_3571,N_2466,N_2519);
nand U3572 (N_3572,N_2561,N_2390);
and U3573 (N_3573,N_2871,N_2860);
or U3574 (N_3574,N_2325,N_2354);
or U3575 (N_3575,N_2578,N_2112);
and U3576 (N_3576,N_2757,N_2403);
and U3577 (N_3577,N_2232,N_2247);
and U3578 (N_3578,N_2246,N_2244);
or U3579 (N_3579,N_2318,N_2288);
or U3580 (N_3580,N_2352,N_2750);
nand U3581 (N_3581,N_2910,N_2549);
and U3582 (N_3582,N_2927,N_2697);
and U3583 (N_3583,N_2533,N_2555);
nand U3584 (N_3584,N_2208,N_2904);
nand U3585 (N_3585,N_2261,N_2588);
nor U3586 (N_3586,N_2768,N_2557);
and U3587 (N_3587,N_2753,N_2466);
or U3588 (N_3588,N_2884,N_2101);
xor U3589 (N_3589,N_2654,N_2627);
and U3590 (N_3590,N_2123,N_2932);
nor U3591 (N_3591,N_2279,N_2528);
nor U3592 (N_3592,N_2744,N_2726);
or U3593 (N_3593,N_2702,N_2262);
nand U3594 (N_3594,N_2097,N_2685);
xnor U3595 (N_3595,N_2722,N_2112);
nand U3596 (N_3596,N_2129,N_2335);
nand U3597 (N_3597,N_2340,N_2538);
nor U3598 (N_3598,N_2020,N_2586);
nand U3599 (N_3599,N_2510,N_2747);
and U3600 (N_3600,N_2693,N_2811);
xnor U3601 (N_3601,N_2805,N_2610);
nor U3602 (N_3602,N_2430,N_2136);
xnor U3603 (N_3603,N_2547,N_2982);
nor U3604 (N_3604,N_2463,N_2483);
nand U3605 (N_3605,N_2757,N_2598);
nor U3606 (N_3606,N_2565,N_2158);
and U3607 (N_3607,N_2083,N_2361);
and U3608 (N_3608,N_2584,N_2820);
xnor U3609 (N_3609,N_2024,N_2462);
or U3610 (N_3610,N_2740,N_2624);
and U3611 (N_3611,N_2263,N_2372);
or U3612 (N_3612,N_2654,N_2220);
nand U3613 (N_3613,N_2859,N_2167);
or U3614 (N_3614,N_2961,N_2377);
nand U3615 (N_3615,N_2947,N_2474);
nand U3616 (N_3616,N_2089,N_2063);
and U3617 (N_3617,N_2828,N_2944);
nand U3618 (N_3618,N_2721,N_2107);
and U3619 (N_3619,N_2040,N_2667);
and U3620 (N_3620,N_2890,N_2048);
xnor U3621 (N_3621,N_2048,N_2362);
and U3622 (N_3622,N_2567,N_2806);
and U3623 (N_3623,N_2393,N_2867);
xor U3624 (N_3624,N_2215,N_2649);
nor U3625 (N_3625,N_2205,N_2118);
nand U3626 (N_3626,N_2713,N_2664);
or U3627 (N_3627,N_2009,N_2859);
or U3628 (N_3628,N_2227,N_2275);
and U3629 (N_3629,N_2355,N_2100);
and U3630 (N_3630,N_2983,N_2284);
nor U3631 (N_3631,N_2644,N_2036);
nand U3632 (N_3632,N_2453,N_2980);
nand U3633 (N_3633,N_2760,N_2510);
nand U3634 (N_3634,N_2551,N_2549);
nand U3635 (N_3635,N_2969,N_2874);
xnor U3636 (N_3636,N_2139,N_2198);
nand U3637 (N_3637,N_2658,N_2909);
nand U3638 (N_3638,N_2943,N_2685);
xor U3639 (N_3639,N_2378,N_2482);
nand U3640 (N_3640,N_2769,N_2002);
and U3641 (N_3641,N_2460,N_2350);
nand U3642 (N_3642,N_2988,N_2737);
nor U3643 (N_3643,N_2860,N_2613);
xor U3644 (N_3644,N_2295,N_2269);
nand U3645 (N_3645,N_2406,N_2754);
nand U3646 (N_3646,N_2114,N_2675);
nor U3647 (N_3647,N_2941,N_2768);
or U3648 (N_3648,N_2527,N_2403);
nand U3649 (N_3649,N_2808,N_2313);
or U3650 (N_3650,N_2651,N_2115);
nor U3651 (N_3651,N_2648,N_2882);
or U3652 (N_3652,N_2989,N_2767);
or U3653 (N_3653,N_2764,N_2745);
nor U3654 (N_3654,N_2436,N_2069);
xor U3655 (N_3655,N_2509,N_2304);
nor U3656 (N_3656,N_2726,N_2613);
or U3657 (N_3657,N_2766,N_2583);
or U3658 (N_3658,N_2376,N_2175);
xnor U3659 (N_3659,N_2722,N_2236);
and U3660 (N_3660,N_2846,N_2016);
nand U3661 (N_3661,N_2619,N_2206);
nor U3662 (N_3662,N_2982,N_2287);
or U3663 (N_3663,N_2008,N_2548);
or U3664 (N_3664,N_2090,N_2746);
or U3665 (N_3665,N_2884,N_2965);
xor U3666 (N_3666,N_2572,N_2376);
nor U3667 (N_3667,N_2669,N_2017);
nor U3668 (N_3668,N_2152,N_2326);
nor U3669 (N_3669,N_2317,N_2297);
and U3670 (N_3670,N_2861,N_2968);
and U3671 (N_3671,N_2471,N_2223);
nor U3672 (N_3672,N_2590,N_2615);
or U3673 (N_3673,N_2262,N_2479);
and U3674 (N_3674,N_2138,N_2063);
nor U3675 (N_3675,N_2477,N_2348);
nor U3676 (N_3676,N_2976,N_2290);
or U3677 (N_3677,N_2671,N_2637);
nor U3678 (N_3678,N_2095,N_2835);
nor U3679 (N_3679,N_2691,N_2510);
nor U3680 (N_3680,N_2636,N_2635);
and U3681 (N_3681,N_2527,N_2014);
and U3682 (N_3682,N_2399,N_2714);
and U3683 (N_3683,N_2847,N_2427);
nor U3684 (N_3684,N_2237,N_2198);
nand U3685 (N_3685,N_2984,N_2273);
or U3686 (N_3686,N_2600,N_2592);
nand U3687 (N_3687,N_2584,N_2290);
or U3688 (N_3688,N_2209,N_2563);
or U3689 (N_3689,N_2784,N_2001);
nor U3690 (N_3690,N_2533,N_2670);
or U3691 (N_3691,N_2703,N_2176);
nand U3692 (N_3692,N_2933,N_2344);
nand U3693 (N_3693,N_2172,N_2965);
or U3694 (N_3694,N_2202,N_2467);
xnor U3695 (N_3695,N_2783,N_2284);
or U3696 (N_3696,N_2979,N_2393);
nand U3697 (N_3697,N_2810,N_2241);
nor U3698 (N_3698,N_2384,N_2631);
nand U3699 (N_3699,N_2853,N_2985);
xor U3700 (N_3700,N_2225,N_2076);
and U3701 (N_3701,N_2022,N_2789);
or U3702 (N_3702,N_2690,N_2360);
nor U3703 (N_3703,N_2829,N_2708);
nand U3704 (N_3704,N_2075,N_2188);
or U3705 (N_3705,N_2340,N_2799);
nand U3706 (N_3706,N_2057,N_2148);
or U3707 (N_3707,N_2679,N_2874);
xor U3708 (N_3708,N_2476,N_2364);
or U3709 (N_3709,N_2456,N_2618);
and U3710 (N_3710,N_2489,N_2114);
or U3711 (N_3711,N_2006,N_2366);
or U3712 (N_3712,N_2836,N_2482);
nand U3713 (N_3713,N_2952,N_2043);
xnor U3714 (N_3714,N_2285,N_2784);
xor U3715 (N_3715,N_2103,N_2264);
nor U3716 (N_3716,N_2631,N_2265);
and U3717 (N_3717,N_2514,N_2228);
or U3718 (N_3718,N_2076,N_2925);
nand U3719 (N_3719,N_2545,N_2678);
or U3720 (N_3720,N_2630,N_2995);
nand U3721 (N_3721,N_2372,N_2700);
and U3722 (N_3722,N_2625,N_2232);
and U3723 (N_3723,N_2061,N_2256);
or U3724 (N_3724,N_2548,N_2656);
and U3725 (N_3725,N_2789,N_2432);
nor U3726 (N_3726,N_2216,N_2590);
and U3727 (N_3727,N_2466,N_2331);
nor U3728 (N_3728,N_2667,N_2812);
xnor U3729 (N_3729,N_2600,N_2402);
nor U3730 (N_3730,N_2918,N_2067);
xor U3731 (N_3731,N_2590,N_2962);
or U3732 (N_3732,N_2814,N_2710);
and U3733 (N_3733,N_2954,N_2354);
xnor U3734 (N_3734,N_2232,N_2162);
nand U3735 (N_3735,N_2276,N_2650);
xnor U3736 (N_3736,N_2950,N_2873);
or U3737 (N_3737,N_2993,N_2075);
and U3738 (N_3738,N_2413,N_2900);
nor U3739 (N_3739,N_2579,N_2304);
nor U3740 (N_3740,N_2674,N_2453);
or U3741 (N_3741,N_2777,N_2253);
nand U3742 (N_3742,N_2146,N_2422);
nand U3743 (N_3743,N_2152,N_2944);
xor U3744 (N_3744,N_2537,N_2492);
nand U3745 (N_3745,N_2878,N_2520);
nor U3746 (N_3746,N_2779,N_2224);
nand U3747 (N_3747,N_2057,N_2969);
nor U3748 (N_3748,N_2389,N_2627);
and U3749 (N_3749,N_2299,N_2057);
nor U3750 (N_3750,N_2414,N_2246);
or U3751 (N_3751,N_2545,N_2150);
and U3752 (N_3752,N_2467,N_2510);
xnor U3753 (N_3753,N_2512,N_2483);
xor U3754 (N_3754,N_2368,N_2502);
nand U3755 (N_3755,N_2840,N_2959);
or U3756 (N_3756,N_2865,N_2642);
nor U3757 (N_3757,N_2318,N_2597);
xnor U3758 (N_3758,N_2205,N_2259);
nand U3759 (N_3759,N_2212,N_2986);
and U3760 (N_3760,N_2187,N_2731);
nand U3761 (N_3761,N_2592,N_2732);
and U3762 (N_3762,N_2724,N_2744);
nand U3763 (N_3763,N_2562,N_2425);
and U3764 (N_3764,N_2541,N_2046);
xor U3765 (N_3765,N_2888,N_2935);
and U3766 (N_3766,N_2378,N_2704);
or U3767 (N_3767,N_2557,N_2035);
xor U3768 (N_3768,N_2812,N_2832);
nor U3769 (N_3769,N_2884,N_2143);
nor U3770 (N_3770,N_2332,N_2095);
or U3771 (N_3771,N_2174,N_2784);
nor U3772 (N_3772,N_2540,N_2068);
xnor U3773 (N_3773,N_2752,N_2038);
nor U3774 (N_3774,N_2298,N_2263);
nor U3775 (N_3775,N_2278,N_2468);
or U3776 (N_3776,N_2835,N_2256);
or U3777 (N_3777,N_2076,N_2746);
or U3778 (N_3778,N_2773,N_2585);
or U3779 (N_3779,N_2386,N_2882);
or U3780 (N_3780,N_2965,N_2599);
nor U3781 (N_3781,N_2611,N_2904);
or U3782 (N_3782,N_2115,N_2412);
xor U3783 (N_3783,N_2877,N_2947);
nor U3784 (N_3784,N_2121,N_2945);
or U3785 (N_3785,N_2614,N_2099);
xor U3786 (N_3786,N_2666,N_2746);
or U3787 (N_3787,N_2134,N_2527);
and U3788 (N_3788,N_2280,N_2701);
and U3789 (N_3789,N_2960,N_2909);
and U3790 (N_3790,N_2941,N_2672);
nor U3791 (N_3791,N_2624,N_2767);
or U3792 (N_3792,N_2789,N_2013);
nand U3793 (N_3793,N_2097,N_2480);
xnor U3794 (N_3794,N_2422,N_2467);
nand U3795 (N_3795,N_2851,N_2565);
xor U3796 (N_3796,N_2368,N_2771);
or U3797 (N_3797,N_2295,N_2739);
nor U3798 (N_3798,N_2010,N_2356);
xor U3799 (N_3799,N_2076,N_2468);
and U3800 (N_3800,N_2182,N_2285);
xnor U3801 (N_3801,N_2130,N_2668);
or U3802 (N_3802,N_2525,N_2330);
or U3803 (N_3803,N_2743,N_2617);
nand U3804 (N_3804,N_2038,N_2783);
xor U3805 (N_3805,N_2765,N_2637);
xnor U3806 (N_3806,N_2617,N_2870);
xnor U3807 (N_3807,N_2355,N_2362);
nand U3808 (N_3808,N_2264,N_2667);
nand U3809 (N_3809,N_2943,N_2555);
xnor U3810 (N_3810,N_2987,N_2256);
xnor U3811 (N_3811,N_2305,N_2232);
nand U3812 (N_3812,N_2270,N_2288);
nand U3813 (N_3813,N_2015,N_2597);
or U3814 (N_3814,N_2537,N_2434);
nor U3815 (N_3815,N_2810,N_2532);
nor U3816 (N_3816,N_2261,N_2939);
nor U3817 (N_3817,N_2455,N_2295);
or U3818 (N_3818,N_2330,N_2583);
xnor U3819 (N_3819,N_2404,N_2825);
and U3820 (N_3820,N_2178,N_2701);
or U3821 (N_3821,N_2726,N_2925);
xnor U3822 (N_3822,N_2358,N_2845);
xor U3823 (N_3823,N_2127,N_2154);
xor U3824 (N_3824,N_2947,N_2076);
and U3825 (N_3825,N_2656,N_2506);
xnor U3826 (N_3826,N_2080,N_2645);
and U3827 (N_3827,N_2441,N_2975);
and U3828 (N_3828,N_2703,N_2847);
nor U3829 (N_3829,N_2469,N_2358);
xor U3830 (N_3830,N_2000,N_2696);
xnor U3831 (N_3831,N_2354,N_2591);
nor U3832 (N_3832,N_2362,N_2519);
nor U3833 (N_3833,N_2601,N_2083);
or U3834 (N_3834,N_2098,N_2836);
and U3835 (N_3835,N_2200,N_2231);
nand U3836 (N_3836,N_2974,N_2950);
or U3837 (N_3837,N_2521,N_2095);
nand U3838 (N_3838,N_2500,N_2257);
and U3839 (N_3839,N_2336,N_2010);
nor U3840 (N_3840,N_2095,N_2269);
nor U3841 (N_3841,N_2975,N_2810);
xnor U3842 (N_3842,N_2768,N_2010);
xor U3843 (N_3843,N_2664,N_2659);
xor U3844 (N_3844,N_2357,N_2982);
nor U3845 (N_3845,N_2197,N_2331);
nor U3846 (N_3846,N_2405,N_2680);
nor U3847 (N_3847,N_2801,N_2790);
nand U3848 (N_3848,N_2263,N_2996);
nand U3849 (N_3849,N_2601,N_2067);
nor U3850 (N_3850,N_2437,N_2020);
and U3851 (N_3851,N_2044,N_2124);
xor U3852 (N_3852,N_2293,N_2155);
nor U3853 (N_3853,N_2555,N_2333);
or U3854 (N_3854,N_2732,N_2708);
nand U3855 (N_3855,N_2707,N_2591);
nor U3856 (N_3856,N_2391,N_2122);
xnor U3857 (N_3857,N_2580,N_2476);
and U3858 (N_3858,N_2553,N_2165);
or U3859 (N_3859,N_2571,N_2380);
and U3860 (N_3860,N_2857,N_2427);
xor U3861 (N_3861,N_2190,N_2825);
nand U3862 (N_3862,N_2639,N_2197);
xor U3863 (N_3863,N_2578,N_2595);
xor U3864 (N_3864,N_2395,N_2414);
and U3865 (N_3865,N_2359,N_2386);
nand U3866 (N_3866,N_2848,N_2811);
or U3867 (N_3867,N_2243,N_2364);
and U3868 (N_3868,N_2193,N_2470);
or U3869 (N_3869,N_2955,N_2323);
or U3870 (N_3870,N_2996,N_2300);
nor U3871 (N_3871,N_2518,N_2698);
and U3872 (N_3872,N_2869,N_2053);
nand U3873 (N_3873,N_2725,N_2502);
xor U3874 (N_3874,N_2987,N_2266);
or U3875 (N_3875,N_2870,N_2859);
nor U3876 (N_3876,N_2776,N_2367);
or U3877 (N_3877,N_2740,N_2224);
nor U3878 (N_3878,N_2262,N_2918);
and U3879 (N_3879,N_2513,N_2480);
nor U3880 (N_3880,N_2573,N_2711);
nand U3881 (N_3881,N_2053,N_2767);
nand U3882 (N_3882,N_2171,N_2372);
xnor U3883 (N_3883,N_2360,N_2983);
nand U3884 (N_3884,N_2529,N_2627);
nor U3885 (N_3885,N_2777,N_2472);
and U3886 (N_3886,N_2657,N_2621);
nand U3887 (N_3887,N_2124,N_2499);
or U3888 (N_3888,N_2634,N_2523);
xnor U3889 (N_3889,N_2225,N_2129);
or U3890 (N_3890,N_2774,N_2652);
nand U3891 (N_3891,N_2066,N_2162);
xor U3892 (N_3892,N_2695,N_2577);
nor U3893 (N_3893,N_2457,N_2498);
and U3894 (N_3894,N_2197,N_2375);
and U3895 (N_3895,N_2998,N_2172);
xor U3896 (N_3896,N_2808,N_2979);
or U3897 (N_3897,N_2815,N_2992);
xor U3898 (N_3898,N_2347,N_2058);
and U3899 (N_3899,N_2830,N_2534);
nand U3900 (N_3900,N_2073,N_2138);
nand U3901 (N_3901,N_2250,N_2682);
nor U3902 (N_3902,N_2614,N_2174);
and U3903 (N_3903,N_2643,N_2453);
and U3904 (N_3904,N_2798,N_2029);
nand U3905 (N_3905,N_2823,N_2605);
nand U3906 (N_3906,N_2925,N_2982);
nand U3907 (N_3907,N_2512,N_2152);
xor U3908 (N_3908,N_2230,N_2541);
xnor U3909 (N_3909,N_2370,N_2262);
xor U3910 (N_3910,N_2205,N_2003);
xnor U3911 (N_3911,N_2049,N_2026);
or U3912 (N_3912,N_2402,N_2268);
xnor U3913 (N_3913,N_2132,N_2031);
and U3914 (N_3914,N_2591,N_2246);
and U3915 (N_3915,N_2818,N_2021);
and U3916 (N_3916,N_2727,N_2678);
and U3917 (N_3917,N_2981,N_2008);
nor U3918 (N_3918,N_2525,N_2630);
nor U3919 (N_3919,N_2588,N_2454);
or U3920 (N_3920,N_2752,N_2593);
nor U3921 (N_3921,N_2295,N_2053);
xor U3922 (N_3922,N_2647,N_2114);
nand U3923 (N_3923,N_2376,N_2038);
xnor U3924 (N_3924,N_2950,N_2043);
xnor U3925 (N_3925,N_2154,N_2918);
and U3926 (N_3926,N_2312,N_2670);
or U3927 (N_3927,N_2940,N_2002);
nand U3928 (N_3928,N_2388,N_2689);
xor U3929 (N_3929,N_2580,N_2226);
xnor U3930 (N_3930,N_2511,N_2732);
nand U3931 (N_3931,N_2986,N_2345);
xnor U3932 (N_3932,N_2000,N_2179);
nor U3933 (N_3933,N_2793,N_2838);
xnor U3934 (N_3934,N_2251,N_2395);
xnor U3935 (N_3935,N_2537,N_2422);
xor U3936 (N_3936,N_2810,N_2168);
and U3937 (N_3937,N_2116,N_2129);
nand U3938 (N_3938,N_2934,N_2244);
nand U3939 (N_3939,N_2330,N_2591);
xnor U3940 (N_3940,N_2836,N_2767);
and U3941 (N_3941,N_2614,N_2618);
and U3942 (N_3942,N_2196,N_2455);
or U3943 (N_3943,N_2064,N_2008);
nand U3944 (N_3944,N_2741,N_2861);
nor U3945 (N_3945,N_2702,N_2396);
nand U3946 (N_3946,N_2681,N_2571);
and U3947 (N_3947,N_2213,N_2333);
nand U3948 (N_3948,N_2362,N_2792);
nor U3949 (N_3949,N_2037,N_2885);
and U3950 (N_3950,N_2355,N_2816);
and U3951 (N_3951,N_2052,N_2516);
nand U3952 (N_3952,N_2114,N_2781);
nor U3953 (N_3953,N_2848,N_2465);
nand U3954 (N_3954,N_2329,N_2762);
or U3955 (N_3955,N_2758,N_2443);
nand U3956 (N_3956,N_2348,N_2763);
nand U3957 (N_3957,N_2061,N_2676);
and U3958 (N_3958,N_2318,N_2763);
xor U3959 (N_3959,N_2851,N_2581);
or U3960 (N_3960,N_2981,N_2713);
or U3961 (N_3961,N_2664,N_2038);
xnor U3962 (N_3962,N_2296,N_2590);
or U3963 (N_3963,N_2472,N_2523);
nand U3964 (N_3964,N_2211,N_2736);
nor U3965 (N_3965,N_2695,N_2536);
nand U3966 (N_3966,N_2472,N_2201);
or U3967 (N_3967,N_2337,N_2844);
or U3968 (N_3968,N_2820,N_2799);
nand U3969 (N_3969,N_2998,N_2462);
and U3970 (N_3970,N_2488,N_2261);
nor U3971 (N_3971,N_2457,N_2133);
and U3972 (N_3972,N_2721,N_2222);
nor U3973 (N_3973,N_2073,N_2086);
and U3974 (N_3974,N_2616,N_2065);
xor U3975 (N_3975,N_2835,N_2755);
nand U3976 (N_3976,N_2318,N_2567);
or U3977 (N_3977,N_2956,N_2881);
nor U3978 (N_3978,N_2158,N_2786);
xor U3979 (N_3979,N_2579,N_2460);
or U3980 (N_3980,N_2668,N_2924);
nor U3981 (N_3981,N_2232,N_2815);
nand U3982 (N_3982,N_2023,N_2062);
and U3983 (N_3983,N_2720,N_2457);
and U3984 (N_3984,N_2492,N_2666);
and U3985 (N_3985,N_2011,N_2065);
nand U3986 (N_3986,N_2672,N_2174);
or U3987 (N_3987,N_2962,N_2474);
and U3988 (N_3988,N_2685,N_2883);
or U3989 (N_3989,N_2886,N_2688);
xnor U3990 (N_3990,N_2130,N_2713);
or U3991 (N_3991,N_2062,N_2625);
and U3992 (N_3992,N_2815,N_2656);
nand U3993 (N_3993,N_2297,N_2824);
and U3994 (N_3994,N_2563,N_2582);
nor U3995 (N_3995,N_2500,N_2187);
nor U3996 (N_3996,N_2593,N_2665);
and U3997 (N_3997,N_2272,N_2239);
and U3998 (N_3998,N_2642,N_2021);
xor U3999 (N_3999,N_2292,N_2185);
nand U4000 (N_4000,N_3987,N_3378);
or U4001 (N_4001,N_3808,N_3464);
nor U4002 (N_4002,N_3973,N_3603);
xor U4003 (N_4003,N_3752,N_3506);
nand U4004 (N_4004,N_3666,N_3228);
xor U4005 (N_4005,N_3685,N_3801);
and U4006 (N_4006,N_3495,N_3065);
or U4007 (N_4007,N_3853,N_3848);
nor U4008 (N_4008,N_3929,N_3935);
nor U4009 (N_4009,N_3241,N_3533);
nor U4010 (N_4010,N_3689,N_3042);
or U4011 (N_4011,N_3069,N_3424);
and U4012 (N_4012,N_3851,N_3707);
or U4013 (N_4013,N_3056,N_3868);
nand U4014 (N_4014,N_3679,N_3649);
nor U4015 (N_4015,N_3718,N_3030);
or U4016 (N_4016,N_3058,N_3341);
xnor U4017 (N_4017,N_3842,N_3107);
nand U4018 (N_4018,N_3849,N_3158);
and U4019 (N_4019,N_3912,N_3717);
nor U4020 (N_4020,N_3772,N_3338);
and U4021 (N_4021,N_3913,N_3402);
nand U4022 (N_4022,N_3963,N_3719);
nor U4023 (N_4023,N_3833,N_3596);
nor U4024 (N_4024,N_3996,N_3906);
xor U4025 (N_4025,N_3527,N_3617);
nor U4026 (N_4026,N_3359,N_3890);
nor U4027 (N_4027,N_3975,N_3312);
or U4028 (N_4028,N_3780,N_3151);
nand U4029 (N_4029,N_3447,N_3381);
nand U4030 (N_4030,N_3931,N_3462);
nor U4031 (N_4031,N_3737,N_3574);
nor U4032 (N_4032,N_3052,N_3310);
and U4033 (N_4033,N_3543,N_3037);
nor U4034 (N_4034,N_3704,N_3117);
xor U4035 (N_4035,N_3620,N_3003);
xor U4036 (N_4036,N_3271,N_3641);
nor U4037 (N_4037,N_3962,N_3988);
nand U4038 (N_4038,N_3916,N_3759);
and U4039 (N_4039,N_3284,N_3604);
xor U4040 (N_4040,N_3933,N_3440);
xor U4041 (N_4041,N_3882,N_3231);
nor U4042 (N_4042,N_3026,N_3124);
nor U4043 (N_4043,N_3136,N_3751);
nor U4044 (N_4044,N_3125,N_3781);
xor U4045 (N_4045,N_3484,N_3471);
and U4046 (N_4046,N_3370,N_3578);
nand U4047 (N_4047,N_3302,N_3485);
nor U4048 (N_4048,N_3678,N_3909);
and U4049 (N_4049,N_3840,N_3281);
xor U4050 (N_4050,N_3315,N_3092);
or U4051 (N_4051,N_3353,N_3735);
or U4052 (N_4052,N_3309,N_3754);
nand U4053 (N_4053,N_3984,N_3562);
xnor U4054 (N_4054,N_3321,N_3957);
and U4055 (N_4055,N_3000,N_3624);
or U4056 (N_4056,N_3896,N_3655);
nand U4057 (N_4057,N_3073,N_3016);
nor U4058 (N_4058,N_3263,N_3764);
or U4059 (N_4059,N_3580,N_3377);
and U4060 (N_4060,N_3834,N_3443);
or U4061 (N_4061,N_3932,N_3711);
xnor U4062 (N_4062,N_3811,N_3647);
or U4063 (N_4063,N_3285,N_3040);
xnor U4064 (N_4064,N_3223,N_3989);
nor U4065 (N_4065,N_3945,N_3725);
nand U4066 (N_4066,N_3750,N_3260);
nand U4067 (N_4067,N_3045,N_3998);
nor U4068 (N_4068,N_3164,N_3943);
xnor U4069 (N_4069,N_3809,N_3976);
or U4070 (N_4070,N_3209,N_3034);
nor U4071 (N_4071,N_3863,N_3036);
and U4072 (N_4072,N_3395,N_3902);
nand U4073 (N_4073,N_3010,N_3382);
or U4074 (N_4074,N_3047,N_3537);
or U4075 (N_4075,N_3978,N_3405);
or U4076 (N_4076,N_3161,N_3992);
or U4077 (N_4077,N_3272,N_3584);
and U4078 (N_4078,N_3638,N_3111);
nor U4079 (N_4079,N_3736,N_3261);
nand U4080 (N_4080,N_3441,N_3345);
and U4081 (N_4081,N_3545,N_3552);
nand U4082 (N_4082,N_3091,N_3756);
xor U4083 (N_4083,N_3313,N_3077);
nor U4084 (N_4084,N_3776,N_3292);
and U4085 (N_4085,N_3826,N_3248);
nand U4086 (N_4086,N_3726,N_3390);
nand U4087 (N_4087,N_3720,N_3773);
nand U4088 (N_4088,N_3525,N_3983);
and U4089 (N_4089,N_3924,N_3814);
xnor U4090 (N_4090,N_3761,N_3386);
xor U4091 (N_4091,N_3192,N_3547);
and U4092 (N_4092,N_3593,N_3577);
or U4093 (N_4093,N_3796,N_3822);
and U4094 (N_4094,N_3304,N_3152);
xor U4095 (N_4095,N_3234,N_3439);
or U4096 (N_4096,N_3371,N_3326);
nand U4097 (N_4097,N_3046,N_3160);
nand U4098 (N_4098,N_3749,N_3592);
or U4099 (N_4099,N_3004,N_3907);
and U4100 (N_4100,N_3311,N_3400);
nand U4101 (N_4101,N_3994,N_3430);
nor U4102 (N_4102,N_3431,N_3145);
and U4103 (N_4103,N_3274,N_3905);
and U4104 (N_4104,N_3232,N_3007);
or U4105 (N_4105,N_3089,N_3183);
and U4106 (N_4106,N_3275,N_3565);
nor U4107 (N_4107,N_3657,N_3013);
nor U4108 (N_4108,N_3434,N_3939);
and U4109 (N_4109,N_3143,N_3385);
and U4110 (N_4110,N_3952,N_3530);
and U4111 (N_4111,N_3605,N_3061);
nor U4112 (N_4112,N_3244,N_3934);
xor U4113 (N_4113,N_3612,N_3100);
nand U4114 (N_4114,N_3887,N_3406);
nand U4115 (N_4115,N_3366,N_3599);
nor U4116 (N_4116,N_3129,N_3270);
xnor U4117 (N_4117,N_3810,N_3384);
and U4118 (N_4118,N_3731,N_3419);
nand U4119 (N_4119,N_3873,N_3049);
and U4120 (N_4120,N_3150,N_3894);
xnor U4121 (N_4121,N_3408,N_3460);
xor U4122 (N_4122,N_3410,N_3482);
and U4123 (N_4123,N_3297,N_3096);
nand U4124 (N_4124,N_3173,N_3277);
and U4125 (N_4125,N_3211,N_3680);
nand U4126 (N_4126,N_3083,N_3288);
nand U4127 (N_4127,N_3551,N_3131);
nand U4128 (N_4128,N_3889,N_3835);
and U4129 (N_4129,N_3119,N_3216);
nor U4130 (N_4130,N_3937,N_3573);
nand U4131 (N_4131,N_3587,N_3757);
xnor U4132 (N_4132,N_3886,N_3306);
or U4133 (N_4133,N_3544,N_3861);
or U4134 (N_4134,N_3249,N_3301);
and U4135 (N_4135,N_3815,N_3467);
and U4136 (N_4136,N_3613,N_3895);
or U4137 (N_4137,N_3528,N_3546);
nand U4138 (N_4138,N_3182,N_3576);
xor U4139 (N_4139,N_3739,N_3661);
nor U4140 (N_4140,N_3558,N_3062);
nor U4141 (N_4141,N_3219,N_3702);
xnor U4142 (N_4142,N_3942,N_3884);
and U4143 (N_4143,N_3463,N_3137);
xnor U4144 (N_4144,N_3729,N_3695);
nand U4145 (N_4145,N_3893,N_3944);
and U4146 (N_4146,N_3844,N_3287);
and U4147 (N_4147,N_3608,N_3162);
xnor U4148 (N_4148,N_3171,N_3144);
nand U4149 (N_4149,N_3289,N_3930);
nand U4150 (N_4150,N_3841,N_3324);
nand U4151 (N_4151,N_3305,N_3455);
or U4152 (N_4152,N_3266,N_3224);
and U4153 (N_4153,N_3466,N_3489);
nand U4154 (N_4154,N_3519,N_3332);
nand U4155 (N_4155,N_3350,N_3559);
nand U4156 (N_4156,N_3213,N_3012);
nor U4157 (N_4157,N_3548,N_3361);
and U4158 (N_4158,N_3867,N_3128);
or U4159 (N_4159,N_3018,N_3958);
nand U4160 (N_4160,N_3947,N_3193);
nor U4161 (N_4161,N_3043,N_3391);
or U4162 (N_4162,N_3334,N_3102);
and U4163 (N_4163,N_3741,N_3055);
nand U4164 (N_4164,N_3793,N_3493);
nor U4165 (N_4165,N_3340,N_3885);
and U4166 (N_4166,N_3291,N_3174);
xnor U4167 (N_4167,N_3600,N_3870);
or U4168 (N_4168,N_3633,N_3966);
or U4169 (N_4169,N_3444,N_3675);
nand U4170 (N_4170,N_3714,N_3303);
xnor U4171 (N_4171,N_3256,N_3081);
or U4172 (N_4172,N_3433,N_3713);
or U4173 (N_4173,N_3412,N_3662);
nand U4174 (N_4174,N_3509,N_3101);
nand U4175 (N_4175,N_3368,N_3403);
nand U4176 (N_4176,N_3053,N_3316);
nor U4177 (N_4177,N_3293,N_3511);
nand U4178 (N_4178,N_3166,N_3106);
nand U4179 (N_4179,N_3372,N_3563);
nor U4180 (N_4180,N_3154,N_3995);
nand U4181 (N_4181,N_3398,N_3888);
xnor U4182 (N_4182,N_3926,N_3855);
xor U4183 (N_4183,N_3475,N_3588);
or U4184 (N_4184,N_3454,N_3199);
xnor U4185 (N_4185,N_3308,N_3407);
xnor U4186 (N_4186,N_3524,N_3487);
nor U4187 (N_4187,N_3254,N_3597);
and U4188 (N_4188,N_3832,N_3622);
nand U4189 (N_4189,N_3257,N_3207);
or U4190 (N_4190,N_3985,N_3428);
xor U4191 (N_4191,N_3222,N_3342);
or U4192 (N_4192,N_3255,N_3025);
and U4193 (N_4193,N_3331,N_3191);
or U4194 (N_4194,N_3696,N_3076);
nand U4195 (N_4195,N_3630,N_3730);
xnor U4196 (N_4196,N_3420,N_3079);
nor U4197 (N_4197,N_3669,N_3602);
or U4198 (N_4198,N_3869,N_3517);
nor U4199 (N_4199,N_3582,N_3024);
and U4200 (N_4200,N_3964,N_3903);
xor U4201 (N_4201,N_3456,N_3364);
nand U4202 (N_4202,N_3522,N_3508);
nand U4203 (N_4203,N_3017,N_3296);
and U4204 (N_4204,N_3705,N_3011);
or U4205 (N_4205,N_3362,N_3948);
and U4206 (N_4206,N_3616,N_3442);
nand U4207 (N_4207,N_3072,N_3694);
nand U4208 (N_4208,N_3572,N_3346);
nand U4209 (N_4209,N_3220,N_3828);
or U4210 (N_4210,N_3788,N_3418);
and U4211 (N_4211,N_3583,N_3795);
or U4212 (N_4212,N_3469,N_3784);
xnor U4213 (N_4213,N_3697,N_3643);
nand U4214 (N_4214,N_3591,N_3892);
nor U4215 (N_4215,N_3797,N_3733);
nand U4216 (N_4216,N_3259,N_3268);
xor U4217 (N_4217,N_3575,N_3184);
and U4218 (N_4218,N_3557,N_3067);
and U4219 (N_4219,N_3656,N_3491);
and U4220 (N_4220,N_3701,N_3437);
nand U4221 (N_4221,N_3860,N_3549);
xor U4222 (N_4222,N_3258,N_3969);
nor U4223 (N_4223,N_3170,N_3569);
xnor U4224 (N_4224,N_3060,N_3674);
xor U4225 (N_4225,N_3082,N_3827);
nor U4226 (N_4226,N_3854,N_3817);
xor U4227 (N_4227,N_3747,N_3415);
or U4228 (N_4228,N_3140,N_3483);
and U4229 (N_4229,N_3252,N_3824);
nand U4230 (N_4230,N_3659,N_3745);
and U4231 (N_4231,N_3721,N_3812);
xor U4232 (N_4232,N_3946,N_3997);
nand U4233 (N_4233,N_3635,N_3397);
or U4234 (N_4234,N_3080,N_3028);
and U4235 (N_4235,N_3423,N_3778);
xnor U4236 (N_4236,N_3194,N_3532);
nand U4237 (N_4237,N_3526,N_3123);
nor U4238 (N_4238,N_3634,N_3910);
and U4239 (N_4239,N_3542,N_3044);
nand U4240 (N_4240,N_3746,N_3093);
xor U4241 (N_4241,N_3130,N_3658);
nand U4242 (N_4242,N_3202,N_3319);
xor U4243 (N_4243,N_3878,N_3108);
and U4244 (N_4244,N_3027,N_3858);
or U4245 (N_4245,N_3829,N_3663);
xnor U4246 (N_4246,N_3497,N_3956);
nor U4247 (N_4247,N_3201,N_3413);
nor U4248 (N_4248,N_3198,N_3240);
or U4249 (N_4249,N_3369,N_3498);
and U4250 (N_4250,N_3251,N_3344);
nor U4251 (N_4251,N_3514,N_3059);
xnor U4252 (N_4252,N_3667,N_3054);
xor U4253 (N_4253,N_3438,N_3767);
or U4254 (N_4254,N_3609,N_3404);
nor U4255 (N_4255,N_3477,N_3769);
and U4256 (N_4256,N_3347,N_3226);
xor U4257 (N_4257,N_3928,N_3792);
xnor U4258 (N_4258,N_3621,N_3105);
nor U4259 (N_4259,N_3852,N_3126);
and U4260 (N_4260,N_3200,N_3090);
nand U4261 (N_4261,N_3692,N_3961);
xor U4262 (N_4262,N_3765,N_3560);
or U4263 (N_4263,N_3221,N_3023);
nor U4264 (N_4264,N_3639,N_3210);
or U4265 (N_4265,N_3640,N_3122);
or U4266 (N_4266,N_3180,N_3539);
and U4267 (N_4267,N_3771,N_3927);
xor U4268 (N_4268,N_3020,N_3941);
xor U4269 (N_4269,N_3472,N_3185);
xor U4270 (N_4270,N_3022,N_3499);
xor U4271 (N_4271,N_3611,N_3336);
nor U4272 (N_4272,N_3269,N_3755);
nor U4273 (N_4273,N_3116,N_3950);
nand U4274 (N_4274,N_3488,N_3607);
or U4275 (N_4275,N_3283,N_3389);
nor U4276 (N_4276,N_3553,N_3461);
xnor U4277 (N_4277,N_3529,N_3001);
nor U4278 (N_4278,N_3307,N_3416);
nor U4279 (N_4279,N_3479,N_3146);
and U4280 (N_4280,N_3156,N_3979);
xor U4281 (N_4281,N_3917,N_3169);
or U4282 (N_4282,N_3791,N_3465);
and U4283 (N_4283,N_3084,N_3758);
or U4284 (N_4284,N_3686,N_3352);
nor U4285 (N_4285,N_3951,N_3449);
or U4286 (N_4286,N_3682,N_3057);
xnor U4287 (N_4287,N_3967,N_3496);
xnor U4288 (N_4288,N_3866,N_3133);
nand U4289 (N_4289,N_3401,N_3790);
or U4290 (N_4290,N_3919,N_3448);
xnor U4291 (N_4291,N_3877,N_3214);
and U4292 (N_4292,N_3710,N_3328);
or U4293 (N_4293,N_3492,N_3881);
nor U4294 (N_4294,N_3006,N_3627);
nand U4295 (N_4295,N_3243,N_3282);
nor U4296 (N_4296,N_3699,N_3501);
xor U4297 (N_4297,N_3783,N_3922);
nor U4298 (N_4298,N_3333,N_3744);
nand U4299 (N_4299,N_3112,N_3982);
nor U4300 (N_4300,N_3348,N_3625);
xor U4301 (N_4301,N_3644,N_3891);
xnor U4302 (N_4302,N_3949,N_3993);
and U4303 (N_4303,N_3300,N_3915);
nor U4304 (N_4304,N_3740,N_3113);
nor U4305 (N_4305,N_3110,N_3299);
nor U4306 (N_4306,N_3276,N_3516);
and U4307 (N_4307,N_3706,N_3375);
and U4308 (N_4308,N_3864,N_3693);
nor U4309 (N_4309,N_3813,N_3615);
and U4310 (N_4310,N_3816,N_3339);
or U4311 (N_4311,N_3230,N_3148);
nor U4312 (N_4312,N_3770,N_3436);
nor U4313 (N_4313,N_3618,N_3388);
nand U4314 (N_4314,N_3322,N_3538);
xor U4315 (N_4315,N_3677,N_3581);
nand U4316 (N_4316,N_3651,N_3648);
and U4317 (N_4317,N_3349,N_3088);
or U4318 (N_4318,N_3005,N_3262);
xor U4319 (N_4319,N_3728,N_3103);
or U4320 (N_4320,N_3354,N_3186);
nor U4321 (N_4321,N_3986,N_3195);
nor U4322 (N_4322,N_3253,N_3033);
and U4323 (N_4323,N_3175,N_3245);
nand U4324 (N_4324,N_3280,N_3120);
nand U4325 (N_4325,N_3642,N_3564);
and U4326 (N_4326,N_3490,N_3954);
or U4327 (N_4327,N_3601,N_3804);
and U4328 (N_4328,N_3229,N_3874);
nor U4329 (N_4329,N_3021,N_3380);
xor U4330 (N_4330,N_3698,N_3898);
and U4331 (N_4331,N_3178,N_3504);
nor U4332 (N_4332,N_3862,N_3429);
or U4333 (N_4333,N_3879,N_3500);
or U4334 (N_4334,N_3654,N_3708);
nor U4335 (N_4335,N_3847,N_3723);
nor U4336 (N_4336,N_3665,N_3290);
and U4337 (N_4337,N_3494,N_3238);
nor U4338 (N_4338,N_3074,N_3265);
nor U4339 (N_4339,N_3645,N_3684);
or U4340 (N_4340,N_3821,N_3298);
or U4341 (N_4341,N_3660,N_3980);
nor U4342 (N_4342,N_3267,N_3035);
or U4343 (N_4343,N_3365,N_3203);
and U4344 (N_4344,N_3337,N_3176);
and U4345 (N_4345,N_3807,N_3716);
or U4346 (N_4346,N_3722,N_3872);
nand U4347 (N_4347,N_3513,N_3589);
nand U4348 (N_4348,N_3383,N_3078);
nor U4349 (N_4349,N_3512,N_3357);
and U4350 (N_4350,N_3628,N_3838);
or U4351 (N_4351,N_3570,N_3374);
and U4352 (N_4352,N_3970,N_3085);
or U4353 (N_4353,N_3250,N_3457);
nor U4354 (N_4354,N_3568,N_3155);
or U4355 (N_4355,N_3118,N_3846);
nor U4356 (N_4356,N_3075,N_3048);
or U4357 (N_4357,N_3911,N_3918);
nor U4358 (N_4358,N_3990,N_3836);
xor U4359 (N_4359,N_3865,N_3738);
or U4360 (N_4360,N_3327,N_3031);
nor U4361 (N_4361,N_3190,N_3206);
and U4362 (N_4362,N_3139,N_3953);
or U4363 (N_4363,N_3153,N_3217);
nor U4364 (N_4364,N_3550,N_3786);
nand U4365 (N_4365,N_3317,N_3325);
xnor U4366 (N_4366,N_3205,N_3278);
nand U4367 (N_4367,N_3646,N_3520);
and U4368 (N_4368,N_3938,N_3831);
nand U4369 (N_4369,N_3687,N_3051);
nor U4370 (N_4370,N_3802,N_3399);
nor U4371 (N_4371,N_3329,N_3104);
nand U4372 (N_4372,N_3664,N_3474);
nand U4373 (N_4373,N_3215,N_3800);
nor U4374 (N_4374,N_3163,N_3727);
or U4375 (N_4375,N_3411,N_3534);
nor U4376 (N_4376,N_3187,N_3619);
nor U4377 (N_4377,N_3273,N_3503);
and U4378 (N_4378,N_3114,N_3820);
nor U4379 (N_4379,N_3880,N_3452);
and U4380 (N_4380,N_3787,N_3782);
nor U4381 (N_4381,N_3435,N_3159);
or U4382 (N_4382,N_3335,N_3507);
nor U4383 (N_4383,N_3960,N_3505);
nand U4384 (N_4384,N_3502,N_3806);
nand U4385 (N_4385,N_3775,N_3768);
nand U4386 (N_4386,N_3459,N_3330);
or U4387 (N_4387,N_3208,N_3177);
or U4388 (N_4388,N_3715,N_3473);
nor U4389 (N_4389,N_3421,N_3856);
xor U4390 (N_4390,N_3556,N_3355);
or U4391 (N_4391,N_3540,N_3805);
nand U4392 (N_4392,N_3039,N_3753);
xnor U4393 (N_4393,N_3971,N_3585);
nand U4394 (N_4394,N_3900,N_3940);
nand U4395 (N_4395,N_3566,N_3636);
nor U4396 (N_4396,N_3819,N_3923);
or U4397 (N_4397,N_3393,N_3857);
nor U4398 (N_4398,N_3671,N_3426);
xnor U4399 (N_4399,N_3632,N_3172);
or U4400 (N_4400,N_3785,N_3087);
or U4401 (N_4401,N_3631,N_3571);
nor U4402 (N_4402,N_3458,N_3009);
or U4403 (N_4403,N_3233,N_3239);
nor U4404 (N_4404,N_3595,N_3068);
xor U4405 (N_4405,N_3681,N_3070);
or U4406 (N_4406,N_3237,N_3181);
or U4407 (N_4407,N_3127,N_3132);
or U4408 (N_4408,N_3323,N_3379);
nor U4409 (N_4409,N_3197,N_3314);
xnor U4410 (N_4410,N_3981,N_3871);
nor U4411 (N_4411,N_3883,N_3991);
and U4412 (N_4412,N_3904,N_3286);
nand U4413 (N_4413,N_3097,N_3225);
or U4414 (N_4414,N_3610,N_3486);
nand U4415 (N_4415,N_3959,N_3850);
nor U4416 (N_4416,N_3914,N_3320);
xor U4417 (N_4417,N_3394,N_3936);
or U4418 (N_4418,N_3859,N_3157);
or U4419 (N_4419,N_3015,N_3732);
and U4420 (N_4420,N_3515,N_3830);
nand U4421 (N_4421,N_3897,N_3598);
nand U4422 (N_4422,N_3766,N_3446);
nor U4423 (N_4423,N_3799,N_3196);
nand U4424 (N_4424,N_3063,N_3724);
xor U4425 (N_4425,N_3367,N_3818);
or U4426 (N_4426,N_3652,N_3843);
xnor U4427 (N_4427,N_3774,N_3521);
or U4428 (N_4428,N_3358,N_3242);
nand U4429 (N_4429,N_3373,N_3476);
nand U4430 (N_4430,N_3637,N_3921);
nor U4431 (N_4431,N_3279,N_3029);
nor U4432 (N_4432,N_3032,N_3204);
nand U4433 (N_4433,N_3839,N_3343);
nor U4434 (N_4434,N_3518,N_3363);
xor U4435 (N_4435,N_3541,N_3086);
xnor U4436 (N_4436,N_3825,N_3974);
or U4437 (N_4437,N_3920,N_3908);
nand U4438 (N_4438,N_3392,N_3899);
or U4439 (N_4439,N_3236,N_3734);
and U4440 (N_4440,N_3650,N_3246);
nor U4441 (N_4441,N_3167,N_3823);
or U4442 (N_4442,N_3700,N_3218);
xnor U4443 (N_4443,N_3064,N_3247);
or U4444 (N_4444,N_3789,N_3691);
nand U4445 (N_4445,N_3586,N_3555);
xnor U4446 (N_4446,N_3189,N_3427);
xnor U4447 (N_4447,N_3876,N_3703);
nand U4448 (N_4448,N_3968,N_3095);
and U4449 (N_4449,N_3676,N_3134);
nor U4450 (N_4450,N_3417,N_3121);
xor U4451 (N_4451,N_3478,N_3451);
or U4452 (N_4452,N_3606,N_3875);
xnor U4453 (N_4453,N_3779,N_3227);
xnor U4454 (N_4454,N_3977,N_3019);
nor U4455 (N_4455,N_3623,N_3798);
or U4456 (N_4456,N_3235,N_3688);
and U4457 (N_4457,N_3098,N_3748);
nand U4458 (N_4458,N_3387,N_3165);
xor U4459 (N_4459,N_3099,N_3425);
xor U4460 (N_4460,N_3535,N_3432);
nor U4461 (N_4461,N_3803,N_3683);
and U4462 (N_4462,N_3561,N_3837);
nand U4463 (N_4463,N_3450,N_3554);
and U4464 (N_4464,N_3742,N_3453);
and U4465 (N_4465,N_3149,N_3673);
xnor U4466 (N_4466,N_3445,N_3041);
xnor U4467 (N_4467,N_3179,N_3141);
and U4468 (N_4468,N_3138,N_3579);
nor U4469 (N_4469,N_3999,N_3972);
and U4470 (N_4470,N_3531,N_3294);
and U4471 (N_4471,N_3212,N_3360);
nor U4472 (N_4472,N_3925,N_3653);
xor U4473 (N_4473,N_3050,N_3008);
nand U4474 (N_4474,N_3762,N_3590);
xor U4475 (N_4475,N_3168,N_3743);
nor U4476 (N_4476,N_3955,N_3071);
and U4477 (N_4477,N_3147,N_3709);
nor U4478 (N_4478,N_3115,N_3794);
nand U4479 (N_4479,N_3094,N_3629);
and U4480 (N_4480,N_3760,N_3356);
nand U4481 (N_4481,N_3965,N_3712);
and U4482 (N_4482,N_3002,N_3066);
and U4483 (N_4483,N_3038,N_3422);
or U4484 (N_4484,N_3777,N_3376);
and U4485 (N_4485,N_3264,N_3351);
or U4486 (N_4486,N_3670,N_3594);
nand U4487 (N_4487,N_3481,N_3295);
nor U4488 (N_4488,N_3480,N_3672);
or U4489 (N_4489,N_3409,N_3845);
nand U4490 (N_4490,N_3135,N_3536);
nand U4491 (N_4491,N_3614,N_3510);
nand U4492 (N_4492,N_3690,N_3901);
and U4493 (N_4493,N_3142,N_3414);
nand U4494 (N_4494,N_3188,N_3523);
nor U4495 (N_4495,N_3763,N_3668);
xnor U4496 (N_4496,N_3014,N_3470);
xnor U4497 (N_4497,N_3567,N_3396);
nand U4498 (N_4498,N_3626,N_3109);
nor U4499 (N_4499,N_3318,N_3468);
or U4500 (N_4500,N_3595,N_3805);
or U4501 (N_4501,N_3592,N_3188);
xor U4502 (N_4502,N_3427,N_3895);
and U4503 (N_4503,N_3366,N_3334);
and U4504 (N_4504,N_3282,N_3995);
or U4505 (N_4505,N_3831,N_3125);
or U4506 (N_4506,N_3492,N_3038);
nor U4507 (N_4507,N_3258,N_3276);
and U4508 (N_4508,N_3712,N_3466);
and U4509 (N_4509,N_3469,N_3400);
nor U4510 (N_4510,N_3557,N_3693);
nand U4511 (N_4511,N_3094,N_3127);
nand U4512 (N_4512,N_3746,N_3463);
or U4513 (N_4513,N_3476,N_3473);
and U4514 (N_4514,N_3244,N_3667);
or U4515 (N_4515,N_3534,N_3607);
or U4516 (N_4516,N_3051,N_3981);
and U4517 (N_4517,N_3313,N_3588);
and U4518 (N_4518,N_3719,N_3863);
and U4519 (N_4519,N_3482,N_3670);
nor U4520 (N_4520,N_3217,N_3473);
xor U4521 (N_4521,N_3538,N_3936);
or U4522 (N_4522,N_3697,N_3605);
and U4523 (N_4523,N_3610,N_3411);
nor U4524 (N_4524,N_3208,N_3693);
nor U4525 (N_4525,N_3439,N_3656);
or U4526 (N_4526,N_3738,N_3764);
or U4527 (N_4527,N_3212,N_3452);
or U4528 (N_4528,N_3509,N_3048);
or U4529 (N_4529,N_3901,N_3100);
or U4530 (N_4530,N_3519,N_3856);
and U4531 (N_4531,N_3481,N_3732);
nor U4532 (N_4532,N_3552,N_3618);
xnor U4533 (N_4533,N_3595,N_3900);
nand U4534 (N_4534,N_3889,N_3907);
nand U4535 (N_4535,N_3211,N_3051);
nor U4536 (N_4536,N_3716,N_3068);
nand U4537 (N_4537,N_3890,N_3044);
and U4538 (N_4538,N_3129,N_3648);
and U4539 (N_4539,N_3826,N_3617);
nor U4540 (N_4540,N_3263,N_3521);
or U4541 (N_4541,N_3462,N_3340);
nand U4542 (N_4542,N_3195,N_3875);
xnor U4543 (N_4543,N_3432,N_3244);
or U4544 (N_4544,N_3584,N_3044);
and U4545 (N_4545,N_3157,N_3167);
or U4546 (N_4546,N_3840,N_3624);
nand U4547 (N_4547,N_3280,N_3668);
or U4548 (N_4548,N_3093,N_3099);
nand U4549 (N_4549,N_3958,N_3732);
xnor U4550 (N_4550,N_3667,N_3780);
nor U4551 (N_4551,N_3977,N_3909);
xor U4552 (N_4552,N_3169,N_3391);
and U4553 (N_4553,N_3870,N_3733);
and U4554 (N_4554,N_3824,N_3697);
or U4555 (N_4555,N_3637,N_3837);
nor U4556 (N_4556,N_3062,N_3184);
and U4557 (N_4557,N_3199,N_3273);
nand U4558 (N_4558,N_3165,N_3237);
xnor U4559 (N_4559,N_3583,N_3607);
nand U4560 (N_4560,N_3206,N_3291);
and U4561 (N_4561,N_3689,N_3193);
nor U4562 (N_4562,N_3735,N_3220);
nand U4563 (N_4563,N_3360,N_3146);
nand U4564 (N_4564,N_3093,N_3834);
nor U4565 (N_4565,N_3902,N_3530);
xnor U4566 (N_4566,N_3886,N_3919);
nor U4567 (N_4567,N_3397,N_3062);
xnor U4568 (N_4568,N_3947,N_3035);
xor U4569 (N_4569,N_3011,N_3561);
and U4570 (N_4570,N_3946,N_3210);
nor U4571 (N_4571,N_3049,N_3191);
or U4572 (N_4572,N_3726,N_3239);
and U4573 (N_4573,N_3841,N_3457);
and U4574 (N_4574,N_3292,N_3793);
nand U4575 (N_4575,N_3487,N_3372);
and U4576 (N_4576,N_3671,N_3973);
and U4577 (N_4577,N_3419,N_3771);
nor U4578 (N_4578,N_3041,N_3446);
or U4579 (N_4579,N_3878,N_3344);
and U4580 (N_4580,N_3939,N_3509);
nor U4581 (N_4581,N_3484,N_3075);
and U4582 (N_4582,N_3836,N_3989);
nor U4583 (N_4583,N_3047,N_3990);
or U4584 (N_4584,N_3064,N_3137);
xor U4585 (N_4585,N_3617,N_3697);
and U4586 (N_4586,N_3560,N_3627);
xor U4587 (N_4587,N_3891,N_3328);
nor U4588 (N_4588,N_3561,N_3781);
or U4589 (N_4589,N_3332,N_3174);
or U4590 (N_4590,N_3335,N_3038);
and U4591 (N_4591,N_3844,N_3624);
and U4592 (N_4592,N_3708,N_3962);
and U4593 (N_4593,N_3129,N_3237);
and U4594 (N_4594,N_3068,N_3263);
nor U4595 (N_4595,N_3826,N_3723);
nand U4596 (N_4596,N_3304,N_3833);
nand U4597 (N_4597,N_3901,N_3896);
and U4598 (N_4598,N_3094,N_3775);
nand U4599 (N_4599,N_3958,N_3482);
xnor U4600 (N_4600,N_3769,N_3232);
nor U4601 (N_4601,N_3780,N_3364);
or U4602 (N_4602,N_3701,N_3048);
nand U4603 (N_4603,N_3516,N_3605);
nor U4604 (N_4604,N_3503,N_3993);
nand U4605 (N_4605,N_3416,N_3546);
or U4606 (N_4606,N_3269,N_3858);
xor U4607 (N_4607,N_3681,N_3672);
or U4608 (N_4608,N_3376,N_3115);
nor U4609 (N_4609,N_3672,N_3529);
and U4610 (N_4610,N_3667,N_3074);
and U4611 (N_4611,N_3483,N_3536);
nand U4612 (N_4612,N_3714,N_3491);
or U4613 (N_4613,N_3515,N_3846);
nand U4614 (N_4614,N_3432,N_3958);
xnor U4615 (N_4615,N_3053,N_3622);
or U4616 (N_4616,N_3808,N_3175);
and U4617 (N_4617,N_3285,N_3337);
or U4618 (N_4618,N_3725,N_3156);
nor U4619 (N_4619,N_3183,N_3722);
and U4620 (N_4620,N_3794,N_3350);
or U4621 (N_4621,N_3771,N_3308);
and U4622 (N_4622,N_3279,N_3416);
xor U4623 (N_4623,N_3443,N_3108);
or U4624 (N_4624,N_3489,N_3949);
xor U4625 (N_4625,N_3567,N_3875);
or U4626 (N_4626,N_3701,N_3271);
and U4627 (N_4627,N_3859,N_3413);
nand U4628 (N_4628,N_3990,N_3206);
and U4629 (N_4629,N_3948,N_3729);
or U4630 (N_4630,N_3428,N_3458);
or U4631 (N_4631,N_3664,N_3482);
nor U4632 (N_4632,N_3646,N_3458);
nand U4633 (N_4633,N_3537,N_3669);
nand U4634 (N_4634,N_3478,N_3905);
nand U4635 (N_4635,N_3587,N_3021);
nand U4636 (N_4636,N_3913,N_3946);
nor U4637 (N_4637,N_3340,N_3235);
or U4638 (N_4638,N_3777,N_3308);
xnor U4639 (N_4639,N_3463,N_3550);
or U4640 (N_4640,N_3691,N_3964);
xnor U4641 (N_4641,N_3762,N_3060);
or U4642 (N_4642,N_3574,N_3567);
xor U4643 (N_4643,N_3665,N_3227);
or U4644 (N_4644,N_3434,N_3775);
nand U4645 (N_4645,N_3079,N_3491);
xor U4646 (N_4646,N_3267,N_3743);
and U4647 (N_4647,N_3481,N_3409);
nor U4648 (N_4648,N_3635,N_3882);
xnor U4649 (N_4649,N_3814,N_3305);
xor U4650 (N_4650,N_3670,N_3204);
and U4651 (N_4651,N_3682,N_3650);
nand U4652 (N_4652,N_3811,N_3498);
and U4653 (N_4653,N_3195,N_3039);
nor U4654 (N_4654,N_3716,N_3616);
and U4655 (N_4655,N_3318,N_3774);
and U4656 (N_4656,N_3215,N_3104);
and U4657 (N_4657,N_3390,N_3146);
nor U4658 (N_4658,N_3932,N_3887);
nor U4659 (N_4659,N_3913,N_3005);
nand U4660 (N_4660,N_3495,N_3071);
or U4661 (N_4661,N_3384,N_3914);
or U4662 (N_4662,N_3584,N_3428);
nand U4663 (N_4663,N_3448,N_3278);
nor U4664 (N_4664,N_3521,N_3566);
and U4665 (N_4665,N_3887,N_3300);
xor U4666 (N_4666,N_3039,N_3197);
xor U4667 (N_4667,N_3084,N_3557);
xor U4668 (N_4668,N_3757,N_3036);
or U4669 (N_4669,N_3202,N_3766);
nand U4670 (N_4670,N_3219,N_3968);
or U4671 (N_4671,N_3677,N_3578);
and U4672 (N_4672,N_3190,N_3032);
and U4673 (N_4673,N_3966,N_3836);
nand U4674 (N_4674,N_3206,N_3449);
and U4675 (N_4675,N_3937,N_3927);
nand U4676 (N_4676,N_3459,N_3149);
xnor U4677 (N_4677,N_3753,N_3096);
nor U4678 (N_4678,N_3139,N_3510);
nor U4679 (N_4679,N_3319,N_3973);
nand U4680 (N_4680,N_3618,N_3451);
nand U4681 (N_4681,N_3929,N_3415);
xnor U4682 (N_4682,N_3442,N_3863);
and U4683 (N_4683,N_3702,N_3320);
nand U4684 (N_4684,N_3834,N_3388);
or U4685 (N_4685,N_3619,N_3639);
nor U4686 (N_4686,N_3827,N_3960);
xor U4687 (N_4687,N_3689,N_3559);
nand U4688 (N_4688,N_3234,N_3272);
xnor U4689 (N_4689,N_3317,N_3451);
or U4690 (N_4690,N_3048,N_3161);
nand U4691 (N_4691,N_3460,N_3734);
or U4692 (N_4692,N_3369,N_3857);
xor U4693 (N_4693,N_3312,N_3688);
and U4694 (N_4694,N_3846,N_3211);
xor U4695 (N_4695,N_3054,N_3930);
and U4696 (N_4696,N_3609,N_3535);
nand U4697 (N_4697,N_3507,N_3981);
and U4698 (N_4698,N_3574,N_3419);
nor U4699 (N_4699,N_3413,N_3899);
nand U4700 (N_4700,N_3298,N_3775);
or U4701 (N_4701,N_3615,N_3105);
and U4702 (N_4702,N_3906,N_3535);
xor U4703 (N_4703,N_3424,N_3683);
nand U4704 (N_4704,N_3310,N_3044);
xor U4705 (N_4705,N_3523,N_3706);
nand U4706 (N_4706,N_3340,N_3218);
and U4707 (N_4707,N_3379,N_3405);
nor U4708 (N_4708,N_3597,N_3962);
nand U4709 (N_4709,N_3673,N_3724);
nand U4710 (N_4710,N_3296,N_3009);
and U4711 (N_4711,N_3663,N_3458);
or U4712 (N_4712,N_3107,N_3102);
nor U4713 (N_4713,N_3228,N_3574);
or U4714 (N_4714,N_3060,N_3588);
xnor U4715 (N_4715,N_3173,N_3539);
nor U4716 (N_4716,N_3274,N_3791);
nand U4717 (N_4717,N_3300,N_3155);
nor U4718 (N_4718,N_3087,N_3722);
xor U4719 (N_4719,N_3563,N_3385);
and U4720 (N_4720,N_3419,N_3805);
or U4721 (N_4721,N_3354,N_3834);
nor U4722 (N_4722,N_3381,N_3698);
nand U4723 (N_4723,N_3657,N_3850);
nand U4724 (N_4724,N_3092,N_3864);
nand U4725 (N_4725,N_3335,N_3433);
or U4726 (N_4726,N_3515,N_3591);
and U4727 (N_4727,N_3634,N_3670);
or U4728 (N_4728,N_3817,N_3474);
xnor U4729 (N_4729,N_3271,N_3029);
nand U4730 (N_4730,N_3046,N_3856);
nor U4731 (N_4731,N_3224,N_3371);
and U4732 (N_4732,N_3684,N_3788);
xor U4733 (N_4733,N_3204,N_3316);
nand U4734 (N_4734,N_3756,N_3035);
nor U4735 (N_4735,N_3519,N_3604);
xor U4736 (N_4736,N_3683,N_3467);
nand U4737 (N_4737,N_3406,N_3359);
nor U4738 (N_4738,N_3395,N_3817);
nand U4739 (N_4739,N_3014,N_3161);
and U4740 (N_4740,N_3735,N_3578);
nand U4741 (N_4741,N_3816,N_3078);
xnor U4742 (N_4742,N_3100,N_3647);
nor U4743 (N_4743,N_3293,N_3126);
and U4744 (N_4744,N_3573,N_3742);
and U4745 (N_4745,N_3248,N_3358);
or U4746 (N_4746,N_3448,N_3878);
and U4747 (N_4747,N_3038,N_3572);
nor U4748 (N_4748,N_3049,N_3651);
or U4749 (N_4749,N_3753,N_3136);
or U4750 (N_4750,N_3633,N_3100);
nor U4751 (N_4751,N_3842,N_3336);
and U4752 (N_4752,N_3549,N_3662);
nor U4753 (N_4753,N_3694,N_3286);
and U4754 (N_4754,N_3563,N_3642);
nand U4755 (N_4755,N_3161,N_3689);
nand U4756 (N_4756,N_3318,N_3033);
nor U4757 (N_4757,N_3551,N_3022);
and U4758 (N_4758,N_3960,N_3495);
nor U4759 (N_4759,N_3874,N_3984);
nor U4760 (N_4760,N_3090,N_3887);
nand U4761 (N_4761,N_3504,N_3776);
nor U4762 (N_4762,N_3629,N_3181);
xor U4763 (N_4763,N_3396,N_3388);
or U4764 (N_4764,N_3458,N_3032);
and U4765 (N_4765,N_3924,N_3067);
and U4766 (N_4766,N_3214,N_3682);
or U4767 (N_4767,N_3053,N_3571);
or U4768 (N_4768,N_3023,N_3268);
xor U4769 (N_4769,N_3557,N_3585);
xor U4770 (N_4770,N_3143,N_3745);
nand U4771 (N_4771,N_3506,N_3761);
nor U4772 (N_4772,N_3347,N_3437);
xor U4773 (N_4773,N_3042,N_3022);
nor U4774 (N_4774,N_3644,N_3706);
and U4775 (N_4775,N_3634,N_3544);
or U4776 (N_4776,N_3328,N_3702);
and U4777 (N_4777,N_3201,N_3049);
nor U4778 (N_4778,N_3766,N_3916);
xnor U4779 (N_4779,N_3152,N_3570);
or U4780 (N_4780,N_3817,N_3167);
and U4781 (N_4781,N_3171,N_3317);
nor U4782 (N_4782,N_3838,N_3123);
nor U4783 (N_4783,N_3580,N_3407);
nor U4784 (N_4784,N_3664,N_3307);
or U4785 (N_4785,N_3289,N_3836);
nor U4786 (N_4786,N_3682,N_3562);
or U4787 (N_4787,N_3237,N_3367);
and U4788 (N_4788,N_3268,N_3961);
or U4789 (N_4789,N_3233,N_3369);
nor U4790 (N_4790,N_3418,N_3544);
nor U4791 (N_4791,N_3680,N_3859);
nand U4792 (N_4792,N_3817,N_3460);
and U4793 (N_4793,N_3371,N_3907);
nand U4794 (N_4794,N_3550,N_3841);
nor U4795 (N_4795,N_3703,N_3013);
and U4796 (N_4796,N_3343,N_3210);
nand U4797 (N_4797,N_3639,N_3618);
nand U4798 (N_4798,N_3499,N_3183);
nor U4799 (N_4799,N_3137,N_3439);
xnor U4800 (N_4800,N_3034,N_3000);
or U4801 (N_4801,N_3700,N_3651);
xor U4802 (N_4802,N_3333,N_3633);
or U4803 (N_4803,N_3027,N_3917);
xnor U4804 (N_4804,N_3517,N_3340);
or U4805 (N_4805,N_3652,N_3658);
and U4806 (N_4806,N_3323,N_3004);
nand U4807 (N_4807,N_3627,N_3127);
xor U4808 (N_4808,N_3399,N_3805);
xor U4809 (N_4809,N_3291,N_3685);
or U4810 (N_4810,N_3604,N_3271);
and U4811 (N_4811,N_3920,N_3601);
xor U4812 (N_4812,N_3204,N_3805);
nor U4813 (N_4813,N_3652,N_3109);
nand U4814 (N_4814,N_3767,N_3815);
nand U4815 (N_4815,N_3058,N_3005);
xor U4816 (N_4816,N_3858,N_3262);
nand U4817 (N_4817,N_3479,N_3777);
or U4818 (N_4818,N_3524,N_3843);
nor U4819 (N_4819,N_3471,N_3518);
and U4820 (N_4820,N_3695,N_3674);
or U4821 (N_4821,N_3067,N_3179);
and U4822 (N_4822,N_3036,N_3461);
xnor U4823 (N_4823,N_3597,N_3928);
nor U4824 (N_4824,N_3651,N_3172);
and U4825 (N_4825,N_3378,N_3214);
nand U4826 (N_4826,N_3154,N_3069);
nor U4827 (N_4827,N_3453,N_3673);
xor U4828 (N_4828,N_3450,N_3335);
nor U4829 (N_4829,N_3027,N_3279);
or U4830 (N_4830,N_3580,N_3624);
and U4831 (N_4831,N_3143,N_3296);
or U4832 (N_4832,N_3393,N_3455);
nor U4833 (N_4833,N_3657,N_3731);
nand U4834 (N_4834,N_3656,N_3312);
or U4835 (N_4835,N_3310,N_3568);
xnor U4836 (N_4836,N_3803,N_3321);
xnor U4837 (N_4837,N_3571,N_3715);
nand U4838 (N_4838,N_3357,N_3940);
nor U4839 (N_4839,N_3920,N_3257);
nand U4840 (N_4840,N_3292,N_3270);
or U4841 (N_4841,N_3621,N_3825);
nand U4842 (N_4842,N_3325,N_3689);
nor U4843 (N_4843,N_3413,N_3597);
nor U4844 (N_4844,N_3838,N_3779);
xnor U4845 (N_4845,N_3099,N_3233);
and U4846 (N_4846,N_3361,N_3710);
and U4847 (N_4847,N_3364,N_3218);
and U4848 (N_4848,N_3347,N_3595);
or U4849 (N_4849,N_3207,N_3414);
xnor U4850 (N_4850,N_3109,N_3524);
or U4851 (N_4851,N_3262,N_3107);
or U4852 (N_4852,N_3010,N_3786);
and U4853 (N_4853,N_3634,N_3863);
xor U4854 (N_4854,N_3357,N_3328);
or U4855 (N_4855,N_3266,N_3564);
or U4856 (N_4856,N_3822,N_3957);
or U4857 (N_4857,N_3368,N_3747);
xnor U4858 (N_4858,N_3137,N_3464);
nand U4859 (N_4859,N_3157,N_3753);
or U4860 (N_4860,N_3277,N_3781);
xor U4861 (N_4861,N_3129,N_3686);
nor U4862 (N_4862,N_3971,N_3796);
nor U4863 (N_4863,N_3205,N_3273);
nand U4864 (N_4864,N_3477,N_3837);
nor U4865 (N_4865,N_3593,N_3282);
or U4866 (N_4866,N_3883,N_3933);
xnor U4867 (N_4867,N_3392,N_3426);
and U4868 (N_4868,N_3733,N_3584);
or U4869 (N_4869,N_3110,N_3291);
nor U4870 (N_4870,N_3138,N_3537);
nor U4871 (N_4871,N_3453,N_3106);
nor U4872 (N_4872,N_3885,N_3667);
or U4873 (N_4873,N_3966,N_3919);
xor U4874 (N_4874,N_3981,N_3759);
nand U4875 (N_4875,N_3198,N_3401);
nor U4876 (N_4876,N_3988,N_3046);
nor U4877 (N_4877,N_3674,N_3609);
nor U4878 (N_4878,N_3124,N_3793);
xnor U4879 (N_4879,N_3161,N_3820);
or U4880 (N_4880,N_3948,N_3249);
nor U4881 (N_4881,N_3650,N_3823);
and U4882 (N_4882,N_3480,N_3016);
or U4883 (N_4883,N_3132,N_3787);
and U4884 (N_4884,N_3403,N_3666);
nor U4885 (N_4885,N_3448,N_3494);
and U4886 (N_4886,N_3720,N_3393);
nand U4887 (N_4887,N_3629,N_3371);
nand U4888 (N_4888,N_3843,N_3850);
nor U4889 (N_4889,N_3153,N_3830);
xnor U4890 (N_4890,N_3895,N_3844);
nand U4891 (N_4891,N_3712,N_3629);
and U4892 (N_4892,N_3594,N_3000);
nand U4893 (N_4893,N_3999,N_3316);
nor U4894 (N_4894,N_3699,N_3847);
and U4895 (N_4895,N_3868,N_3842);
nand U4896 (N_4896,N_3427,N_3754);
nand U4897 (N_4897,N_3880,N_3172);
or U4898 (N_4898,N_3112,N_3254);
nor U4899 (N_4899,N_3754,N_3421);
and U4900 (N_4900,N_3559,N_3716);
and U4901 (N_4901,N_3189,N_3646);
nor U4902 (N_4902,N_3703,N_3697);
xnor U4903 (N_4903,N_3518,N_3743);
or U4904 (N_4904,N_3362,N_3860);
or U4905 (N_4905,N_3887,N_3994);
nor U4906 (N_4906,N_3816,N_3222);
or U4907 (N_4907,N_3234,N_3382);
or U4908 (N_4908,N_3083,N_3645);
xnor U4909 (N_4909,N_3178,N_3686);
and U4910 (N_4910,N_3248,N_3057);
or U4911 (N_4911,N_3720,N_3370);
and U4912 (N_4912,N_3236,N_3064);
and U4913 (N_4913,N_3405,N_3217);
xnor U4914 (N_4914,N_3145,N_3881);
and U4915 (N_4915,N_3382,N_3360);
nor U4916 (N_4916,N_3046,N_3521);
or U4917 (N_4917,N_3055,N_3239);
or U4918 (N_4918,N_3651,N_3236);
or U4919 (N_4919,N_3129,N_3369);
nor U4920 (N_4920,N_3282,N_3055);
or U4921 (N_4921,N_3927,N_3986);
nand U4922 (N_4922,N_3041,N_3897);
nor U4923 (N_4923,N_3610,N_3373);
and U4924 (N_4924,N_3571,N_3165);
nand U4925 (N_4925,N_3953,N_3044);
nor U4926 (N_4926,N_3067,N_3923);
xnor U4927 (N_4927,N_3028,N_3187);
nand U4928 (N_4928,N_3457,N_3111);
xnor U4929 (N_4929,N_3947,N_3504);
or U4930 (N_4930,N_3899,N_3328);
or U4931 (N_4931,N_3527,N_3284);
or U4932 (N_4932,N_3010,N_3974);
nor U4933 (N_4933,N_3830,N_3821);
or U4934 (N_4934,N_3110,N_3720);
nor U4935 (N_4935,N_3201,N_3979);
nand U4936 (N_4936,N_3243,N_3850);
nor U4937 (N_4937,N_3784,N_3123);
nand U4938 (N_4938,N_3967,N_3294);
xor U4939 (N_4939,N_3914,N_3827);
xor U4940 (N_4940,N_3592,N_3244);
nor U4941 (N_4941,N_3104,N_3490);
nor U4942 (N_4942,N_3270,N_3093);
nor U4943 (N_4943,N_3799,N_3193);
nand U4944 (N_4944,N_3080,N_3144);
xnor U4945 (N_4945,N_3118,N_3007);
nor U4946 (N_4946,N_3694,N_3760);
xnor U4947 (N_4947,N_3259,N_3975);
xor U4948 (N_4948,N_3607,N_3870);
and U4949 (N_4949,N_3101,N_3142);
or U4950 (N_4950,N_3360,N_3493);
or U4951 (N_4951,N_3352,N_3163);
or U4952 (N_4952,N_3960,N_3016);
xor U4953 (N_4953,N_3610,N_3710);
nand U4954 (N_4954,N_3677,N_3626);
and U4955 (N_4955,N_3523,N_3635);
or U4956 (N_4956,N_3350,N_3092);
or U4957 (N_4957,N_3250,N_3412);
nand U4958 (N_4958,N_3635,N_3160);
nand U4959 (N_4959,N_3404,N_3420);
xnor U4960 (N_4960,N_3097,N_3697);
or U4961 (N_4961,N_3214,N_3561);
nand U4962 (N_4962,N_3845,N_3114);
nand U4963 (N_4963,N_3343,N_3043);
and U4964 (N_4964,N_3081,N_3456);
nor U4965 (N_4965,N_3157,N_3243);
nand U4966 (N_4966,N_3090,N_3595);
or U4967 (N_4967,N_3557,N_3543);
xnor U4968 (N_4968,N_3166,N_3307);
xor U4969 (N_4969,N_3446,N_3323);
nor U4970 (N_4970,N_3599,N_3249);
or U4971 (N_4971,N_3790,N_3545);
nor U4972 (N_4972,N_3445,N_3437);
or U4973 (N_4973,N_3686,N_3883);
nor U4974 (N_4974,N_3110,N_3464);
and U4975 (N_4975,N_3345,N_3641);
xnor U4976 (N_4976,N_3657,N_3576);
nor U4977 (N_4977,N_3341,N_3561);
and U4978 (N_4978,N_3465,N_3821);
or U4979 (N_4979,N_3294,N_3947);
nand U4980 (N_4980,N_3171,N_3965);
and U4981 (N_4981,N_3976,N_3385);
and U4982 (N_4982,N_3448,N_3566);
xor U4983 (N_4983,N_3547,N_3565);
nand U4984 (N_4984,N_3915,N_3734);
nand U4985 (N_4985,N_3592,N_3435);
nor U4986 (N_4986,N_3983,N_3828);
or U4987 (N_4987,N_3561,N_3867);
nor U4988 (N_4988,N_3807,N_3978);
nand U4989 (N_4989,N_3060,N_3859);
nor U4990 (N_4990,N_3348,N_3633);
nand U4991 (N_4991,N_3109,N_3164);
nand U4992 (N_4992,N_3654,N_3018);
nor U4993 (N_4993,N_3942,N_3357);
and U4994 (N_4994,N_3291,N_3902);
nand U4995 (N_4995,N_3230,N_3040);
nor U4996 (N_4996,N_3370,N_3380);
and U4997 (N_4997,N_3586,N_3635);
or U4998 (N_4998,N_3678,N_3251);
or U4999 (N_4999,N_3631,N_3263);
or U5000 (N_5000,N_4627,N_4169);
nor U5001 (N_5001,N_4254,N_4320);
and U5002 (N_5002,N_4142,N_4565);
nand U5003 (N_5003,N_4676,N_4209);
nand U5004 (N_5004,N_4573,N_4753);
or U5005 (N_5005,N_4268,N_4233);
or U5006 (N_5006,N_4333,N_4099);
xnor U5007 (N_5007,N_4399,N_4134);
nor U5008 (N_5008,N_4110,N_4473);
nor U5009 (N_5009,N_4535,N_4723);
or U5010 (N_5010,N_4612,N_4450);
nand U5011 (N_5011,N_4445,N_4347);
nand U5012 (N_5012,N_4467,N_4179);
nor U5013 (N_5013,N_4167,N_4215);
or U5014 (N_5014,N_4860,N_4464);
nor U5015 (N_5015,N_4117,N_4139);
or U5016 (N_5016,N_4075,N_4512);
xnor U5017 (N_5017,N_4901,N_4204);
nor U5018 (N_5018,N_4218,N_4704);
or U5019 (N_5019,N_4242,N_4985);
or U5020 (N_5020,N_4505,N_4217);
nand U5021 (N_5021,N_4593,N_4590);
nand U5022 (N_5022,N_4664,N_4061);
and U5023 (N_5023,N_4706,N_4471);
nand U5024 (N_5024,N_4380,N_4720);
xnor U5025 (N_5025,N_4479,N_4662);
and U5026 (N_5026,N_4772,N_4929);
and U5027 (N_5027,N_4731,N_4172);
and U5028 (N_5028,N_4582,N_4097);
nor U5029 (N_5029,N_4787,N_4950);
nand U5030 (N_5030,N_4230,N_4231);
or U5031 (N_5031,N_4629,N_4086);
nor U5032 (N_5032,N_4425,N_4503);
and U5033 (N_5033,N_4406,N_4971);
or U5034 (N_5034,N_4456,N_4304);
or U5035 (N_5035,N_4875,N_4962);
xor U5036 (N_5036,N_4776,N_4454);
or U5037 (N_5037,N_4244,N_4779);
and U5038 (N_5038,N_4543,N_4128);
xor U5039 (N_5039,N_4190,N_4859);
nand U5040 (N_5040,N_4600,N_4730);
or U5041 (N_5041,N_4129,N_4090);
nor U5042 (N_5042,N_4837,N_4422);
nor U5043 (N_5043,N_4031,N_4791);
nor U5044 (N_5044,N_4712,N_4684);
nand U5045 (N_5045,N_4146,N_4625);
xor U5046 (N_5046,N_4006,N_4141);
xnor U5047 (N_5047,N_4558,N_4135);
nor U5048 (N_5048,N_4057,N_4289);
and U5049 (N_5049,N_4883,N_4449);
nor U5050 (N_5050,N_4891,N_4997);
xnor U5051 (N_5051,N_4123,N_4821);
nand U5052 (N_5052,N_4411,N_4307);
or U5053 (N_5053,N_4935,N_4184);
xnor U5054 (N_5054,N_4862,N_4197);
nand U5055 (N_5055,N_4822,N_4889);
or U5056 (N_5056,N_4896,N_4622);
or U5057 (N_5057,N_4469,N_4395);
nor U5058 (N_5058,N_4126,N_4548);
or U5059 (N_5059,N_4127,N_4601);
nand U5060 (N_5060,N_4626,N_4897);
xor U5061 (N_5061,N_4604,N_4843);
xor U5062 (N_5062,N_4178,N_4828);
nor U5063 (N_5063,N_4579,N_4793);
nor U5064 (N_5064,N_4430,N_4675);
or U5065 (N_5065,N_4107,N_4481);
nor U5066 (N_5066,N_4853,N_4749);
or U5067 (N_5067,N_4359,N_4506);
and U5068 (N_5068,N_4115,N_4522);
xor U5069 (N_5069,N_4465,N_4315);
or U5070 (N_5070,N_4887,N_4306);
and U5071 (N_5071,N_4510,N_4874);
nor U5072 (N_5072,N_4188,N_4265);
and U5073 (N_5073,N_4211,N_4034);
or U5074 (N_5074,N_4576,N_4092);
and U5075 (N_5075,N_4832,N_4458);
and U5076 (N_5076,N_4383,N_4526);
or U5077 (N_5077,N_4181,N_4861);
xor U5078 (N_5078,N_4421,N_4413);
nor U5079 (N_5079,N_4235,N_4195);
xor U5080 (N_5080,N_4741,N_4603);
nor U5081 (N_5081,N_4803,N_4963);
and U5082 (N_5082,N_4894,N_4282);
xnor U5083 (N_5083,N_4330,N_4416);
and U5084 (N_5084,N_4846,N_4670);
and U5085 (N_5085,N_4041,N_4327);
xor U5086 (N_5086,N_4507,N_4940);
xor U5087 (N_5087,N_4063,N_4970);
and U5088 (N_5088,N_4234,N_4702);
and U5089 (N_5089,N_4909,N_4984);
nand U5090 (N_5090,N_4767,N_4212);
xnor U5091 (N_5091,N_4453,N_4830);
nor U5092 (N_5092,N_4087,N_4933);
nand U5093 (N_5093,N_4278,N_4228);
nor U5094 (N_5094,N_4485,N_4199);
xor U5095 (N_5095,N_4324,N_4257);
and U5096 (N_5096,N_4343,N_4977);
nand U5097 (N_5097,N_4848,N_4969);
and U5098 (N_5098,N_4439,N_4983);
nor U5099 (N_5099,N_4353,N_4089);
nor U5100 (N_5100,N_4295,N_4067);
xor U5101 (N_5101,N_4293,N_4375);
and U5102 (N_5102,N_4085,N_4273);
nor U5103 (N_5103,N_4666,N_4116);
or U5104 (N_5104,N_4276,N_4559);
or U5105 (N_5105,N_4882,N_4423);
or U5106 (N_5106,N_4342,N_4237);
or U5107 (N_5107,N_4624,N_4154);
xor U5108 (N_5108,N_4007,N_4433);
nand U5109 (N_5109,N_4054,N_4227);
xor U5110 (N_5110,N_4491,N_4694);
nor U5111 (N_5111,N_4403,N_4372);
and U5112 (N_5112,N_4334,N_4355);
xor U5113 (N_5113,N_4957,N_4937);
nand U5114 (N_5114,N_4104,N_4518);
or U5115 (N_5115,N_4816,N_4895);
and U5116 (N_5116,N_4310,N_4258);
and U5117 (N_5117,N_4917,N_4575);
and U5118 (N_5118,N_4768,N_4497);
or U5119 (N_5119,N_4322,N_4932);
or U5120 (N_5120,N_4136,N_4055);
and U5121 (N_5121,N_4384,N_4047);
nor U5122 (N_5122,N_4189,N_4836);
xor U5123 (N_5123,N_4714,N_4763);
and U5124 (N_5124,N_4571,N_4408);
xor U5125 (N_5125,N_4761,N_4160);
or U5126 (N_5126,N_4132,N_4605);
xnor U5127 (N_5127,N_4206,N_4683);
or U5128 (N_5128,N_4918,N_4879);
or U5129 (N_5129,N_4125,N_4030);
or U5130 (N_5130,N_4377,N_4806);
xor U5131 (N_5131,N_4908,N_4020);
nor U5132 (N_5132,N_4826,N_4261);
and U5133 (N_5133,N_4297,N_4825);
or U5134 (N_5134,N_4781,N_4975);
nor U5135 (N_5135,N_4990,N_4474);
or U5136 (N_5136,N_4868,N_4775);
xor U5137 (N_5137,N_4805,N_4358);
or U5138 (N_5138,N_4101,N_4910);
nand U5139 (N_5139,N_4241,N_4298);
or U5140 (N_5140,N_4053,N_4019);
and U5141 (N_5141,N_4687,N_4336);
or U5142 (N_5142,N_4354,N_4619);
and U5143 (N_5143,N_4637,N_4038);
xnor U5144 (N_5144,N_4998,N_4771);
xor U5145 (N_5145,N_4546,N_4913);
nand U5146 (N_5146,N_4109,N_4356);
xnor U5147 (N_5147,N_4371,N_4597);
nor U5148 (N_5148,N_4568,N_4577);
xor U5149 (N_5149,N_4401,N_4900);
nor U5150 (N_5150,N_4810,N_4795);
or U5151 (N_5151,N_4530,N_4120);
or U5152 (N_5152,N_4193,N_4924);
or U5153 (N_5153,N_4713,N_4743);
or U5154 (N_5154,N_4751,N_4317);
or U5155 (N_5155,N_4851,N_4946);
and U5156 (N_5156,N_4740,N_4165);
nand U5157 (N_5157,N_4588,N_4486);
xnor U5158 (N_5158,N_4489,N_4820);
or U5159 (N_5159,N_4798,N_4326);
or U5160 (N_5160,N_4378,N_4688);
nand U5161 (N_5161,N_4583,N_4958);
nor U5162 (N_5162,N_4790,N_4774);
nor U5163 (N_5163,N_4052,N_4321);
nor U5164 (N_5164,N_4400,N_4312);
nand U5165 (N_5165,N_4980,N_4916);
nor U5166 (N_5166,N_4693,N_4208);
and U5167 (N_5167,N_4852,N_4196);
nand U5168 (N_5168,N_4682,N_4564);
nand U5169 (N_5169,N_4490,N_4251);
xnor U5170 (N_5170,N_4750,N_4191);
nor U5171 (N_5171,N_4815,N_4618);
or U5172 (N_5172,N_4655,N_4700);
nor U5173 (N_5173,N_4496,N_4978);
nor U5174 (N_5174,N_4414,N_4850);
and U5175 (N_5175,N_4262,N_4633);
or U5176 (N_5176,N_4721,N_4615);
and U5177 (N_5177,N_4009,N_4867);
and U5178 (N_5178,N_4589,N_4899);
or U5179 (N_5179,N_4029,N_4608);
or U5180 (N_5180,N_4287,N_4886);
xor U5181 (N_5181,N_4409,N_4448);
xnor U5182 (N_5182,N_4728,N_4492);
or U5183 (N_5183,N_4680,N_4532);
nor U5184 (N_5184,N_4701,N_4500);
xor U5185 (N_5185,N_4267,N_4171);
nand U5186 (N_5186,N_4288,N_4480);
nand U5187 (N_5187,N_4407,N_4082);
xnor U5188 (N_5188,N_4854,N_4569);
xnor U5189 (N_5189,N_4441,N_4804);
xnor U5190 (N_5190,N_4494,N_4229);
or U5191 (N_5191,N_4762,N_4391);
nand U5192 (N_5192,N_4769,N_4717);
nand U5193 (N_5193,N_4677,N_4996);
nand U5194 (N_5194,N_4736,N_4443);
xnor U5195 (N_5195,N_4782,N_4872);
nor U5196 (N_5196,N_4809,N_4557);
or U5197 (N_5197,N_4335,N_4551);
or U5198 (N_5198,N_4549,N_4379);
nor U5199 (N_5199,N_4185,N_4180);
xor U5200 (N_5200,N_4245,N_4368);
or U5201 (N_5201,N_4631,N_4387);
and U5202 (N_5202,N_4755,N_4111);
and U5203 (N_5203,N_4070,N_4361);
nor U5204 (N_5204,N_4722,N_4130);
and U5205 (N_5205,N_4028,N_4654);
nand U5206 (N_5206,N_4214,N_4538);
xor U5207 (N_5207,N_4813,N_4079);
nand U5208 (N_5208,N_4147,N_4898);
and U5209 (N_5209,N_4968,N_4133);
nor U5210 (N_5210,N_4071,N_4436);
nor U5211 (N_5211,N_4328,N_4166);
and U5212 (N_5212,N_4834,N_4398);
nor U5213 (N_5213,N_4643,N_4542);
nand U5214 (N_5214,N_4617,N_4058);
or U5215 (N_5215,N_4737,N_4502);
nand U5216 (N_5216,N_4396,N_4650);
xor U5217 (N_5217,N_4056,N_4594);
or U5218 (N_5218,N_4742,N_4153);
nor U5219 (N_5219,N_4942,N_4556);
nand U5220 (N_5220,N_4939,N_4709);
and U5221 (N_5221,N_4632,N_4536);
or U5222 (N_5222,N_4033,N_4673);
or U5223 (N_5223,N_4841,N_4840);
and U5224 (N_5224,N_4961,N_4255);
xor U5225 (N_5225,N_4784,N_4907);
and U5226 (N_5226,N_4048,N_4162);
or U5227 (N_5227,N_4220,N_4871);
nor U5228 (N_5228,N_4074,N_4902);
or U5229 (N_5229,N_4386,N_4691);
and U5230 (N_5230,N_4931,N_4149);
xnor U5231 (N_5231,N_4246,N_4508);
and U5232 (N_5232,N_4986,N_4999);
nand U5233 (N_5233,N_4202,N_4570);
nor U5234 (N_5234,N_4766,N_4599);
nor U5235 (N_5235,N_4281,N_4801);
xor U5236 (N_5236,N_4818,N_4194);
nor U5237 (N_5237,N_4174,N_4018);
nand U5238 (N_5238,N_4253,N_4435);
nand U5239 (N_5239,N_4004,N_4187);
nor U5240 (N_5240,N_4960,N_4303);
or U5241 (N_5241,N_4719,N_4598);
xnor U5242 (N_5242,N_4225,N_4865);
nor U5243 (N_5243,N_4844,N_4239);
nor U5244 (N_5244,N_4431,N_4905);
nand U5245 (N_5245,N_4145,N_4829);
nor U5246 (N_5246,N_4487,N_4752);
nand U5247 (N_5247,N_4892,N_4735);
nand U5248 (N_5248,N_4754,N_4498);
nor U5249 (N_5249,N_4934,N_4250);
and U5250 (N_5250,N_4385,N_4357);
and U5251 (N_5251,N_4098,N_4163);
nand U5252 (N_5252,N_4182,N_4533);
or U5253 (N_5253,N_4340,N_4159);
and U5254 (N_5254,N_4432,N_4168);
or U5255 (N_5255,N_4124,N_4362);
nor U5256 (N_5256,N_4524,N_4103);
and U5257 (N_5257,N_4842,N_4786);
xor U5258 (N_5258,N_4084,N_4747);
nand U5259 (N_5259,N_4122,N_4277);
nor U5260 (N_5260,N_4069,N_4773);
xnor U5261 (N_5261,N_4010,N_4881);
and U5262 (N_5262,N_4945,N_4925);
nand U5263 (N_5263,N_4025,N_4649);
or U5264 (N_5264,N_4402,N_4364);
or U5265 (N_5265,N_4140,N_4080);
and U5266 (N_5266,N_4560,N_4764);
xor U5267 (N_5267,N_4003,N_4628);
and U5268 (N_5268,N_4988,N_4219);
nand U5269 (N_5269,N_4390,N_4667);
xnor U5270 (N_5270,N_4726,N_4252);
xor U5271 (N_5271,N_4697,N_4725);
or U5272 (N_5272,N_4272,N_4156);
and U5273 (N_5273,N_4873,N_4311);
and U5274 (N_5274,N_4426,N_4921);
and U5275 (N_5275,N_4641,N_4094);
and U5276 (N_5276,N_4758,N_4724);
nand U5277 (N_5277,N_4483,N_4213);
or U5278 (N_5278,N_4991,N_4249);
xnor U5279 (N_5279,N_4926,N_4944);
or U5280 (N_5280,N_4349,N_4592);
and U5281 (N_5281,N_4528,N_4525);
nor U5282 (N_5282,N_4200,N_4746);
xnor U5283 (N_5283,N_4131,N_4201);
or U5284 (N_5284,N_4639,N_4482);
xor U5285 (N_5285,N_4039,N_4634);
or U5286 (N_5286,N_4472,N_4927);
or U5287 (N_5287,N_4337,N_4008);
and U5288 (N_5288,N_4351,N_4578);
nand U5289 (N_5289,N_4083,N_4964);
or U5290 (N_5290,N_4446,N_4797);
or U5291 (N_5291,N_4610,N_4369);
nor U5292 (N_5292,N_4022,N_4602);
nor U5293 (N_5293,N_4271,N_4611);
or U5294 (N_5294,N_4096,N_4877);
or U5295 (N_5295,N_4609,N_4965);
nor U5296 (N_5296,N_4065,N_4236);
and U5297 (N_5297,N_4711,N_4366);
and U5298 (N_5298,N_4049,N_4305);
xor U5299 (N_5299,N_4373,N_4027);
or U5300 (N_5300,N_4095,N_4014);
xor U5301 (N_5301,N_4114,N_4678);
or U5302 (N_5302,N_4948,N_4833);
and U5303 (N_5303,N_4459,N_4817);
xnor U5304 (N_5304,N_4428,N_4488);
nor U5305 (N_5305,N_4484,N_4911);
or U5306 (N_5306,N_4581,N_4827);
xor U5307 (N_5307,N_4299,N_4922);
nor U5308 (N_5308,N_4292,N_4596);
xor U5309 (N_5309,N_4947,N_4309);
or U5310 (N_5310,N_4238,N_4112);
or U5311 (N_5311,N_4091,N_4669);
nor U5312 (N_5312,N_4325,N_4595);
xnor U5313 (N_5313,N_4653,N_4170);
and U5314 (N_5314,N_4011,N_4656);
nor U5315 (N_5315,N_4718,N_4685);
and U5316 (N_5316,N_4405,N_4072);
nand U5317 (N_5317,N_4995,N_4585);
nand U5318 (N_5318,N_4759,N_4420);
xor U5319 (N_5319,N_4294,N_4616);
and U5320 (N_5320,N_4550,N_4823);
nor U5321 (N_5321,N_4527,N_4463);
xor U5322 (N_5322,N_4059,N_4920);
or U5323 (N_5323,N_4175,N_4308);
or U5324 (N_5324,N_4705,N_4376);
nor U5325 (N_5325,N_4350,N_4799);
xor U5326 (N_5326,N_4475,N_4105);
or U5327 (N_5327,N_4690,N_4462);
nand U5328 (N_5328,N_4260,N_4976);
and U5329 (N_5329,N_4332,N_4903);
nand U5330 (N_5330,N_4037,N_4437);
xor U5331 (N_5331,N_4040,N_4857);
nor U5332 (N_5332,N_4062,N_4523);
nor U5333 (N_5333,N_4606,N_4138);
nor U5334 (N_5334,N_4636,N_4973);
and U5335 (N_5335,N_4839,N_4064);
or U5336 (N_5336,N_4382,N_4994);
or U5337 (N_5337,N_4584,N_4447);
and U5338 (N_5338,N_4539,N_4158);
xor U5339 (N_5339,N_4613,N_4203);
nor U5340 (N_5340,N_4692,N_4470);
nand U5341 (N_5341,N_4076,N_4529);
xor U5342 (N_5342,N_4013,N_4001);
nand U5343 (N_5343,N_4733,N_4681);
and U5344 (N_5344,N_4424,N_4966);
nor U5345 (N_5345,N_4992,N_4652);
nor U5346 (N_5346,N_4679,N_4906);
or U5347 (N_5347,N_4161,N_4346);
nor U5348 (N_5348,N_4374,N_4869);
nor U5349 (N_5349,N_4476,N_4739);
and U5350 (N_5350,N_4716,N_4183);
xnor U5351 (N_5351,N_4151,N_4205);
xnor U5352 (N_5352,N_4732,N_4660);
nand U5353 (N_5353,N_4291,N_4164);
nand U5354 (N_5354,N_4864,N_4541);
and U5355 (N_5355,N_4259,N_4845);
or U5356 (N_5356,N_4017,N_4381);
or U5357 (N_5357,N_4285,N_4956);
and U5358 (N_5358,N_4300,N_4658);
nand U5359 (N_5359,N_4770,N_4699);
xnor U5360 (N_5360,N_4545,N_4955);
or U5361 (N_5361,N_4587,N_4444);
xor U5362 (N_5362,N_4243,N_4521);
or U5363 (N_5363,N_4301,N_4876);
and U5364 (N_5364,N_4941,N_4451);
nand U5365 (N_5365,N_4478,N_4689);
nor U5366 (N_5366,N_4284,N_4024);
and U5367 (N_5367,N_4914,N_4972);
nor U5368 (N_5368,N_4323,N_4365);
and U5369 (N_5369,N_4192,N_4951);
nor U5370 (N_5370,N_4068,N_4002);
nand U5371 (N_5371,N_4514,N_4102);
nand U5372 (N_5372,N_4638,N_4341);
xor U5373 (N_5373,N_4847,N_4930);
nand U5374 (N_5374,N_4989,N_4499);
nand U5375 (N_5375,N_4248,N_4835);
nand U5376 (N_5376,N_4223,N_4155);
and U5377 (N_5377,N_4412,N_4574);
or U5378 (N_5378,N_4783,N_4352);
nor U5379 (N_5379,N_4173,N_4734);
and U5380 (N_5380,N_4504,N_4296);
nor U5381 (N_5381,N_4036,N_4012);
and U5382 (N_5382,N_4893,N_4544);
nor U5383 (N_5383,N_4046,N_4313);
nand U5384 (N_5384,N_4657,N_4866);
and U5385 (N_5385,N_4547,N_4814);
xor U5386 (N_5386,N_4005,N_4645);
nor U5387 (N_5387,N_4552,N_4648);
nor U5388 (N_5388,N_4247,N_4954);
nand U5389 (N_5389,N_4035,N_4021);
xnor U5390 (N_5390,N_4216,N_4890);
or U5391 (N_5391,N_4952,N_4338);
nor U5392 (N_5392,N_4452,N_4415);
nand U5393 (N_5393,N_4222,N_4517);
or U5394 (N_5394,N_4477,N_4642);
nor U5395 (N_5395,N_4043,N_4286);
and U5396 (N_5396,N_4591,N_4417);
xor U5397 (N_5397,N_4392,N_4314);
and U5398 (N_5398,N_4858,N_4393);
nand U5399 (N_5399,N_4788,N_4904);
nand U5400 (N_5400,N_4959,N_4348);
xnor U5401 (N_5401,N_4993,N_4811);
and U5402 (N_5402,N_4949,N_4644);
nand U5403 (N_5403,N_4884,N_4695);
or U5404 (N_5404,N_4661,N_4427);
nand U5405 (N_5405,N_4290,N_4620);
and U5406 (N_5406,N_4461,N_4434);
and U5407 (N_5407,N_4531,N_4831);
nor U5408 (N_5408,N_4520,N_4455);
nand U5409 (N_5409,N_4912,N_4388);
and U5410 (N_5410,N_4800,N_4081);
nand U5411 (N_5411,N_4729,N_4672);
nor U5412 (N_5412,N_4256,N_4240);
xnor U5413 (N_5413,N_4855,N_4280);
or U5414 (N_5414,N_4563,N_4647);
nor U5415 (N_5415,N_4807,N_4275);
or U5416 (N_5416,N_4819,N_4878);
or U5417 (N_5417,N_4345,N_4440);
xor U5418 (N_5418,N_4051,N_4953);
xnor U5419 (N_5419,N_4106,N_4316);
nor U5420 (N_5420,N_4785,N_4418);
or U5421 (N_5421,N_4000,N_4319);
xor U5422 (N_5422,N_4015,N_4023);
or U5423 (N_5423,N_4756,N_4630);
nand U5424 (N_5424,N_4108,N_4410);
nor U5425 (N_5425,N_4457,N_4659);
or U5426 (N_5426,N_4938,N_4077);
nand U5427 (N_5427,N_4363,N_4495);
and U5428 (N_5428,N_4519,N_4580);
nor U5429 (N_5429,N_4042,N_4438);
xnor U5430 (N_5430,N_4137,N_4561);
nor U5431 (N_5431,N_4674,N_4148);
xnor U5432 (N_5432,N_4808,N_4232);
nand U5433 (N_5433,N_4651,N_4397);
xor U5434 (N_5434,N_4748,N_4572);
and U5435 (N_5435,N_4974,N_4936);
nand U5436 (N_5436,N_4671,N_4144);
xor U5437 (N_5437,N_4554,N_4515);
nand U5438 (N_5438,N_4744,N_4555);
or U5439 (N_5439,N_4943,N_4923);
or U5440 (N_5440,N_4640,N_4915);
nand U5441 (N_5441,N_4919,N_4266);
and U5442 (N_5442,N_4856,N_4665);
or U5443 (N_5443,N_4646,N_4981);
nor U5444 (N_5444,N_4329,N_4143);
or U5445 (N_5445,N_4442,N_4812);
or U5446 (N_5446,N_4460,N_4210);
nor U5447 (N_5447,N_4738,N_4849);
nor U5448 (N_5448,N_4698,N_4283);
nand U5449 (N_5449,N_4888,N_4429);
xor U5450 (N_5450,N_4982,N_4780);
nor U5451 (N_5451,N_4838,N_4073);
or U5452 (N_5452,N_4668,N_4635);
nor U5453 (N_5453,N_4745,N_4318);
xnor U5454 (N_5454,N_4663,N_4686);
nand U5455 (N_5455,N_4100,N_4778);
nor U5456 (N_5456,N_4331,N_4026);
xor U5457 (N_5457,N_4757,N_4198);
and U5458 (N_5458,N_4501,N_4870);
nor U5459 (N_5459,N_4789,N_4511);
nand U5460 (N_5460,N_4760,N_4207);
nor U5461 (N_5461,N_4157,N_4302);
and U5462 (N_5462,N_4270,N_4703);
nand U5463 (N_5463,N_4078,N_4880);
nor U5464 (N_5464,N_4045,N_4050);
and U5465 (N_5465,N_4516,N_4710);
nand U5466 (N_5466,N_4404,N_4562);
xor U5467 (N_5467,N_4623,N_4269);
and U5468 (N_5468,N_4513,N_4987);
nand U5469 (N_5469,N_4979,N_4032);
nor U5470 (N_5470,N_4567,N_4824);
and U5471 (N_5471,N_4044,N_4696);
or U5472 (N_5472,N_4152,N_4176);
and U5473 (N_5473,N_4367,N_4607);
and U5474 (N_5474,N_4279,N_4389);
nand U5475 (N_5475,N_4493,N_4863);
or U5476 (N_5476,N_4534,N_4088);
nor U5477 (N_5477,N_4707,N_4274);
nor U5478 (N_5478,N_4553,N_4468);
or U5479 (N_5479,N_4509,N_4466);
nand U5480 (N_5480,N_4419,N_4118);
and U5481 (N_5481,N_4708,N_4540);
xor U5482 (N_5482,N_4177,N_4794);
and U5483 (N_5483,N_4967,N_4715);
nor U5484 (N_5484,N_4765,N_4360);
xor U5485 (N_5485,N_4928,N_4537);
xor U5486 (N_5486,N_4113,N_4586);
xor U5487 (N_5487,N_4263,N_4221);
nor U5488 (N_5488,N_4119,N_4264);
xnor U5489 (N_5489,N_4796,N_4614);
nor U5490 (N_5490,N_4792,N_4224);
nand U5491 (N_5491,N_4121,N_4802);
nor U5492 (N_5492,N_4066,N_4150);
nor U5493 (N_5493,N_4727,N_4060);
nor U5494 (N_5494,N_4777,N_4621);
and U5495 (N_5495,N_4186,N_4344);
and U5496 (N_5496,N_4226,N_4339);
nand U5497 (N_5497,N_4885,N_4093);
xnor U5498 (N_5498,N_4370,N_4394);
and U5499 (N_5499,N_4016,N_4566);
xnor U5500 (N_5500,N_4826,N_4692);
and U5501 (N_5501,N_4747,N_4374);
and U5502 (N_5502,N_4670,N_4820);
xor U5503 (N_5503,N_4709,N_4920);
xor U5504 (N_5504,N_4090,N_4841);
xnor U5505 (N_5505,N_4917,N_4424);
and U5506 (N_5506,N_4957,N_4546);
nand U5507 (N_5507,N_4122,N_4017);
nand U5508 (N_5508,N_4025,N_4765);
xnor U5509 (N_5509,N_4680,N_4561);
and U5510 (N_5510,N_4820,N_4407);
nand U5511 (N_5511,N_4391,N_4884);
xnor U5512 (N_5512,N_4369,N_4124);
nor U5513 (N_5513,N_4517,N_4209);
nor U5514 (N_5514,N_4067,N_4576);
and U5515 (N_5515,N_4183,N_4351);
nor U5516 (N_5516,N_4511,N_4646);
nor U5517 (N_5517,N_4010,N_4614);
and U5518 (N_5518,N_4663,N_4146);
nor U5519 (N_5519,N_4680,N_4656);
xor U5520 (N_5520,N_4147,N_4826);
or U5521 (N_5521,N_4218,N_4914);
xor U5522 (N_5522,N_4216,N_4611);
xnor U5523 (N_5523,N_4251,N_4197);
and U5524 (N_5524,N_4883,N_4815);
and U5525 (N_5525,N_4014,N_4532);
nand U5526 (N_5526,N_4409,N_4942);
xnor U5527 (N_5527,N_4289,N_4445);
nand U5528 (N_5528,N_4031,N_4512);
nand U5529 (N_5529,N_4945,N_4412);
xor U5530 (N_5530,N_4309,N_4638);
nand U5531 (N_5531,N_4479,N_4116);
nor U5532 (N_5532,N_4210,N_4014);
nor U5533 (N_5533,N_4180,N_4676);
xnor U5534 (N_5534,N_4779,N_4088);
nand U5535 (N_5535,N_4490,N_4550);
nand U5536 (N_5536,N_4481,N_4583);
or U5537 (N_5537,N_4676,N_4962);
or U5538 (N_5538,N_4058,N_4606);
nor U5539 (N_5539,N_4266,N_4804);
and U5540 (N_5540,N_4196,N_4831);
nor U5541 (N_5541,N_4520,N_4563);
or U5542 (N_5542,N_4112,N_4473);
or U5543 (N_5543,N_4418,N_4331);
or U5544 (N_5544,N_4382,N_4085);
and U5545 (N_5545,N_4202,N_4614);
nor U5546 (N_5546,N_4516,N_4844);
or U5547 (N_5547,N_4946,N_4766);
or U5548 (N_5548,N_4499,N_4256);
or U5549 (N_5549,N_4188,N_4864);
xnor U5550 (N_5550,N_4388,N_4262);
nand U5551 (N_5551,N_4541,N_4983);
xnor U5552 (N_5552,N_4218,N_4286);
nor U5553 (N_5553,N_4184,N_4035);
xnor U5554 (N_5554,N_4329,N_4410);
and U5555 (N_5555,N_4289,N_4628);
nand U5556 (N_5556,N_4909,N_4765);
or U5557 (N_5557,N_4638,N_4843);
nand U5558 (N_5558,N_4409,N_4536);
and U5559 (N_5559,N_4229,N_4730);
nand U5560 (N_5560,N_4141,N_4529);
or U5561 (N_5561,N_4326,N_4725);
nor U5562 (N_5562,N_4969,N_4959);
nor U5563 (N_5563,N_4861,N_4102);
and U5564 (N_5564,N_4044,N_4522);
or U5565 (N_5565,N_4755,N_4734);
nand U5566 (N_5566,N_4568,N_4122);
nand U5567 (N_5567,N_4784,N_4645);
and U5568 (N_5568,N_4948,N_4318);
or U5569 (N_5569,N_4323,N_4389);
nand U5570 (N_5570,N_4460,N_4517);
and U5571 (N_5571,N_4960,N_4992);
nand U5572 (N_5572,N_4409,N_4143);
xnor U5573 (N_5573,N_4714,N_4895);
or U5574 (N_5574,N_4091,N_4413);
and U5575 (N_5575,N_4240,N_4281);
nor U5576 (N_5576,N_4655,N_4641);
and U5577 (N_5577,N_4074,N_4337);
and U5578 (N_5578,N_4248,N_4369);
xor U5579 (N_5579,N_4568,N_4600);
and U5580 (N_5580,N_4111,N_4827);
or U5581 (N_5581,N_4757,N_4329);
xnor U5582 (N_5582,N_4851,N_4588);
xor U5583 (N_5583,N_4129,N_4108);
xnor U5584 (N_5584,N_4423,N_4604);
and U5585 (N_5585,N_4988,N_4820);
nand U5586 (N_5586,N_4845,N_4880);
nor U5587 (N_5587,N_4183,N_4103);
nand U5588 (N_5588,N_4619,N_4188);
and U5589 (N_5589,N_4609,N_4996);
xor U5590 (N_5590,N_4287,N_4081);
and U5591 (N_5591,N_4541,N_4457);
or U5592 (N_5592,N_4535,N_4482);
and U5593 (N_5593,N_4133,N_4311);
or U5594 (N_5594,N_4946,N_4857);
and U5595 (N_5595,N_4531,N_4766);
nor U5596 (N_5596,N_4448,N_4887);
or U5597 (N_5597,N_4804,N_4506);
nand U5598 (N_5598,N_4412,N_4861);
nor U5599 (N_5599,N_4234,N_4797);
and U5600 (N_5600,N_4992,N_4203);
xnor U5601 (N_5601,N_4901,N_4115);
nand U5602 (N_5602,N_4075,N_4297);
and U5603 (N_5603,N_4208,N_4037);
or U5604 (N_5604,N_4141,N_4183);
xnor U5605 (N_5605,N_4750,N_4622);
xnor U5606 (N_5606,N_4812,N_4036);
nand U5607 (N_5607,N_4274,N_4420);
or U5608 (N_5608,N_4333,N_4839);
or U5609 (N_5609,N_4212,N_4173);
nand U5610 (N_5610,N_4987,N_4324);
or U5611 (N_5611,N_4905,N_4731);
xnor U5612 (N_5612,N_4365,N_4688);
nor U5613 (N_5613,N_4466,N_4675);
nand U5614 (N_5614,N_4644,N_4225);
nand U5615 (N_5615,N_4112,N_4128);
nand U5616 (N_5616,N_4450,N_4458);
nor U5617 (N_5617,N_4841,N_4344);
or U5618 (N_5618,N_4610,N_4453);
nand U5619 (N_5619,N_4741,N_4844);
xor U5620 (N_5620,N_4903,N_4301);
and U5621 (N_5621,N_4809,N_4960);
and U5622 (N_5622,N_4068,N_4851);
nor U5623 (N_5623,N_4659,N_4765);
nand U5624 (N_5624,N_4703,N_4637);
xor U5625 (N_5625,N_4451,N_4575);
nand U5626 (N_5626,N_4615,N_4384);
nor U5627 (N_5627,N_4308,N_4753);
xnor U5628 (N_5628,N_4555,N_4935);
xnor U5629 (N_5629,N_4344,N_4792);
or U5630 (N_5630,N_4803,N_4377);
nand U5631 (N_5631,N_4929,N_4473);
or U5632 (N_5632,N_4991,N_4458);
nor U5633 (N_5633,N_4030,N_4131);
and U5634 (N_5634,N_4724,N_4981);
nor U5635 (N_5635,N_4908,N_4673);
nand U5636 (N_5636,N_4123,N_4131);
nor U5637 (N_5637,N_4689,N_4591);
and U5638 (N_5638,N_4505,N_4741);
or U5639 (N_5639,N_4070,N_4191);
and U5640 (N_5640,N_4767,N_4303);
xnor U5641 (N_5641,N_4764,N_4719);
nand U5642 (N_5642,N_4347,N_4737);
and U5643 (N_5643,N_4777,N_4044);
nor U5644 (N_5644,N_4621,N_4390);
xor U5645 (N_5645,N_4187,N_4875);
xnor U5646 (N_5646,N_4427,N_4484);
nand U5647 (N_5647,N_4451,N_4025);
xnor U5648 (N_5648,N_4140,N_4790);
nand U5649 (N_5649,N_4709,N_4313);
nor U5650 (N_5650,N_4014,N_4430);
or U5651 (N_5651,N_4702,N_4230);
or U5652 (N_5652,N_4125,N_4138);
or U5653 (N_5653,N_4634,N_4189);
nor U5654 (N_5654,N_4098,N_4601);
nand U5655 (N_5655,N_4302,N_4295);
xnor U5656 (N_5656,N_4136,N_4158);
nand U5657 (N_5657,N_4123,N_4414);
nor U5658 (N_5658,N_4928,N_4121);
xnor U5659 (N_5659,N_4279,N_4719);
nand U5660 (N_5660,N_4894,N_4597);
or U5661 (N_5661,N_4408,N_4866);
xnor U5662 (N_5662,N_4904,N_4029);
xor U5663 (N_5663,N_4640,N_4426);
nor U5664 (N_5664,N_4843,N_4664);
xnor U5665 (N_5665,N_4041,N_4679);
nand U5666 (N_5666,N_4815,N_4192);
nand U5667 (N_5667,N_4054,N_4241);
and U5668 (N_5668,N_4233,N_4421);
xor U5669 (N_5669,N_4399,N_4660);
and U5670 (N_5670,N_4364,N_4470);
xor U5671 (N_5671,N_4410,N_4902);
and U5672 (N_5672,N_4590,N_4748);
and U5673 (N_5673,N_4398,N_4044);
nand U5674 (N_5674,N_4140,N_4380);
xor U5675 (N_5675,N_4010,N_4639);
nand U5676 (N_5676,N_4961,N_4212);
xor U5677 (N_5677,N_4921,N_4892);
xor U5678 (N_5678,N_4204,N_4019);
xor U5679 (N_5679,N_4646,N_4344);
nand U5680 (N_5680,N_4570,N_4069);
xnor U5681 (N_5681,N_4328,N_4747);
xor U5682 (N_5682,N_4477,N_4625);
nor U5683 (N_5683,N_4060,N_4689);
and U5684 (N_5684,N_4631,N_4573);
xnor U5685 (N_5685,N_4441,N_4647);
xor U5686 (N_5686,N_4048,N_4757);
nor U5687 (N_5687,N_4248,N_4298);
nor U5688 (N_5688,N_4046,N_4531);
nor U5689 (N_5689,N_4500,N_4493);
xor U5690 (N_5690,N_4196,N_4430);
or U5691 (N_5691,N_4957,N_4775);
or U5692 (N_5692,N_4389,N_4798);
xnor U5693 (N_5693,N_4538,N_4944);
xor U5694 (N_5694,N_4778,N_4114);
nor U5695 (N_5695,N_4473,N_4020);
and U5696 (N_5696,N_4834,N_4740);
nand U5697 (N_5697,N_4620,N_4988);
or U5698 (N_5698,N_4590,N_4170);
nor U5699 (N_5699,N_4080,N_4628);
nand U5700 (N_5700,N_4398,N_4417);
xnor U5701 (N_5701,N_4378,N_4177);
and U5702 (N_5702,N_4852,N_4604);
xor U5703 (N_5703,N_4675,N_4110);
nor U5704 (N_5704,N_4362,N_4911);
xnor U5705 (N_5705,N_4696,N_4950);
nand U5706 (N_5706,N_4878,N_4542);
nand U5707 (N_5707,N_4589,N_4059);
or U5708 (N_5708,N_4496,N_4825);
and U5709 (N_5709,N_4998,N_4774);
or U5710 (N_5710,N_4006,N_4612);
and U5711 (N_5711,N_4255,N_4680);
or U5712 (N_5712,N_4433,N_4649);
nand U5713 (N_5713,N_4267,N_4609);
or U5714 (N_5714,N_4722,N_4382);
and U5715 (N_5715,N_4297,N_4316);
nor U5716 (N_5716,N_4813,N_4108);
and U5717 (N_5717,N_4863,N_4149);
or U5718 (N_5718,N_4851,N_4050);
nor U5719 (N_5719,N_4862,N_4320);
nand U5720 (N_5720,N_4761,N_4208);
and U5721 (N_5721,N_4874,N_4357);
nand U5722 (N_5722,N_4710,N_4083);
nand U5723 (N_5723,N_4478,N_4650);
nand U5724 (N_5724,N_4401,N_4122);
nand U5725 (N_5725,N_4899,N_4475);
or U5726 (N_5726,N_4291,N_4306);
nand U5727 (N_5727,N_4042,N_4331);
nor U5728 (N_5728,N_4384,N_4935);
xor U5729 (N_5729,N_4896,N_4027);
xor U5730 (N_5730,N_4983,N_4158);
and U5731 (N_5731,N_4823,N_4322);
nor U5732 (N_5732,N_4847,N_4801);
xnor U5733 (N_5733,N_4690,N_4886);
or U5734 (N_5734,N_4600,N_4319);
or U5735 (N_5735,N_4531,N_4025);
or U5736 (N_5736,N_4222,N_4229);
nor U5737 (N_5737,N_4386,N_4445);
nor U5738 (N_5738,N_4928,N_4520);
nand U5739 (N_5739,N_4035,N_4878);
or U5740 (N_5740,N_4450,N_4611);
and U5741 (N_5741,N_4435,N_4138);
or U5742 (N_5742,N_4592,N_4322);
xor U5743 (N_5743,N_4857,N_4224);
and U5744 (N_5744,N_4479,N_4324);
nand U5745 (N_5745,N_4764,N_4566);
or U5746 (N_5746,N_4781,N_4527);
or U5747 (N_5747,N_4509,N_4473);
nand U5748 (N_5748,N_4544,N_4576);
or U5749 (N_5749,N_4685,N_4271);
nor U5750 (N_5750,N_4122,N_4618);
and U5751 (N_5751,N_4492,N_4864);
and U5752 (N_5752,N_4930,N_4413);
xor U5753 (N_5753,N_4057,N_4584);
or U5754 (N_5754,N_4531,N_4593);
nor U5755 (N_5755,N_4907,N_4545);
and U5756 (N_5756,N_4239,N_4553);
or U5757 (N_5757,N_4183,N_4615);
xnor U5758 (N_5758,N_4913,N_4942);
xnor U5759 (N_5759,N_4886,N_4314);
and U5760 (N_5760,N_4613,N_4864);
or U5761 (N_5761,N_4206,N_4541);
xnor U5762 (N_5762,N_4120,N_4655);
xor U5763 (N_5763,N_4854,N_4006);
nand U5764 (N_5764,N_4669,N_4507);
nand U5765 (N_5765,N_4782,N_4709);
xnor U5766 (N_5766,N_4769,N_4854);
nor U5767 (N_5767,N_4095,N_4265);
and U5768 (N_5768,N_4557,N_4529);
and U5769 (N_5769,N_4911,N_4935);
xnor U5770 (N_5770,N_4889,N_4870);
nand U5771 (N_5771,N_4552,N_4771);
or U5772 (N_5772,N_4638,N_4180);
and U5773 (N_5773,N_4811,N_4079);
xor U5774 (N_5774,N_4154,N_4880);
or U5775 (N_5775,N_4867,N_4008);
or U5776 (N_5776,N_4337,N_4228);
xor U5777 (N_5777,N_4254,N_4422);
nor U5778 (N_5778,N_4813,N_4982);
or U5779 (N_5779,N_4162,N_4673);
nor U5780 (N_5780,N_4816,N_4270);
nand U5781 (N_5781,N_4431,N_4536);
or U5782 (N_5782,N_4279,N_4451);
and U5783 (N_5783,N_4389,N_4124);
nor U5784 (N_5784,N_4600,N_4934);
nor U5785 (N_5785,N_4183,N_4500);
nor U5786 (N_5786,N_4520,N_4492);
and U5787 (N_5787,N_4400,N_4500);
nand U5788 (N_5788,N_4668,N_4491);
and U5789 (N_5789,N_4415,N_4311);
nand U5790 (N_5790,N_4305,N_4778);
nor U5791 (N_5791,N_4383,N_4483);
and U5792 (N_5792,N_4658,N_4901);
xnor U5793 (N_5793,N_4430,N_4071);
or U5794 (N_5794,N_4426,N_4441);
nor U5795 (N_5795,N_4843,N_4812);
nor U5796 (N_5796,N_4988,N_4874);
nor U5797 (N_5797,N_4810,N_4231);
xnor U5798 (N_5798,N_4238,N_4924);
nor U5799 (N_5799,N_4203,N_4600);
and U5800 (N_5800,N_4669,N_4836);
or U5801 (N_5801,N_4193,N_4039);
nor U5802 (N_5802,N_4370,N_4514);
nand U5803 (N_5803,N_4951,N_4598);
nor U5804 (N_5804,N_4506,N_4581);
xnor U5805 (N_5805,N_4715,N_4215);
nor U5806 (N_5806,N_4132,N_4055);
or U5807 (N_5807,N_4350,N_4555);
nand U5808 (N_5808,N_4913,N_4460);
and U5809 (N_5809,N_4791,N_4200);
nor U5810 (N_5810,N_4014,N_4146);
or U5811 (N_5811,N_4822,N_4432);
nand U5812 (N_5812,N_4137,N_4665);
nor U5813 (N_5813,N_4950,N_4794);
and U5814 (N_5814,N_4350,N_4032);
xnor U5815 (N_5815,N_4459,N_4171);
and U5816 (N_5816,N_4527,N_4889);
nand U5817 (N_5817,N_4650,N_4470);
or U5818 (N_5818,N_4173,N_4589);
xor U5819 (N_5819,N_4891,N_4191);
nor U5820 (N_5820,N_4972,N_4644);
and U5821 (N_5821,N_4315,N_4982);
and U5822 (N_5822,N_4605,N_4522);
xnor U5823 (N_5823,N_4173,N_4230);
or U5824 (N_5824,N_4352,N_4547);
nor U5825 (N_5825,N_4761,N_4518);
nand U5826 (N_5826,N_4758,N_4999);
nor U5827 (N_5827,N_4106,N_4202);
and U5828 (N_5828,N_4708,N_4546);
or U5829 (N_5829,N_4939,N_4262);
and U5830 (N_5830,N_4882,N_4369);
and U5831 (N_5831,N_4532,N_4397);
or U5832 (N_5832,N_4384,N_4195);
or U5833 (N_5833,N_4386,N_4969);
and U5834 (N_5834,N_4625,N_4041);
or U5835 (N_5835,N_4110,N_4800);
nor U5836 (N_5836,N_4149,N_4636);
or U5837 (N_5837,N_4994,N_4651);
or U5838 (N_5838,N_4423,N_4735);
nand U5839 (N_5839,N_4557,N_4561);
nor U5840 (N_5840,N_4227,N_4926);
and U5841 (N_5841,N_4415,N_4306);
nor U5842 (N_5842,N_4681,N_4650);
xnor U5843 (N_5843,N_4245,N_4295);
and U5844 (N_5844,N_4779,N_4354);
xnor U5845 (N_5845,N_4453,N_4011);
xnor U5846 (N_5846,N_4769,N_4459);
or U5847 (N_5847,N_4020,N_4762);
xnor U5848 (N_5848,N_4265,N_4304);
or U5849 (N_5849,N_4036,N_4554);
xnor U5850 (N_5850,N_4035,N_4564);
nand U5851 (N_5851,N_4007,N_4680);
nor U5852 (N_5852,N_4704,N_4360);
or U5853 (N_5853,N_4751,N_4602);
xnor U5854 (N_5854,N_4741,N_4827);
xor U5855 (N_5855,N_4519,N_4330);
nand U5856 (N_5856,N_4535,N_4464);
xor U5857 (N_5857,N_4480,N_4854);
nor U5858 (N_5858,N_4960,N_4891);
xnor U5859 (N_5859,N_4031,N_4884);
or U5860 (N_5860,N_4970,N_4746);
or U5861 (N_5861,N_4925,N_4303);
xnor U5862 (N_5862,N_4146,N_4608);
and U5863 (N_5863,N_4093,N_4979);
xor U5864 (N_5864,N_4641,N_4169);
xnor U5865 (N_5865,N_4370,N_4666);
or U5866 (N_5866,N_4839,N_4178);
xnor U5867 (N_5867,N_4314,N_4800);
nor U5868 (N_5868,N_4479,N_4034);
and U5869 (N_5869,N_4891,N_4920);
and U5870 (N_5870,N_4042,N_4395);
and U5871 (N_5871,N_4732,N_4625);
and U5872 (N_5872,N_4850,N_4433);
and U5873 (N_5873,N_4899,N_4648);
and U5874 (N_5874,N_4323,N_4192);
nand U5875 (N_5875,N_4700,N_4641);
and U5876 (N_5876,N_4205,N_4053);
nand U5877 (N_5877,N_4678,N_4914);
or U5878 (N_5878,N_4316,N_4709);
xnor U5879 (N_5879,N_4272,N_4394);
nor U5880 (N_5880,N_4755,N_4747);
nand U5881 (N_5881,N_4138,N_4932);
nand U5882 (N_5882,N_4268,N_4365);
xnor U5883 (N_5883,N_4307,N_4199);
and U5884 (N_5884,N_4043,N_4506);
xor U5885 (N_5885,N_4916,N_4519);
or U5886 (N_5886,N_4195,N_4340);
nor U5887 (N_5887,N_4734,N_4598);
nand U5888 (N_5888,N_4039,N_4767);
nor U5889 (N_5889,N_4617,N_4412);
nor U5890 (N_5890,N_4203,N_4777);
and U5891 (N_5891,N_4963,N_4473);
or U5892 (N_5892,N_4191,N_4557);
and U5893 (N_5893,N_4088,N_4998);
nand U5894 (N_5894,N_4089,N_4517);
nor U5895 (N_5895,N_4148,N_4522);
nor U5896 (N_5896,N_4690,N_4560);
nand U5897 (N_5897,N_4455,N_4238);
xnor U5898 (N_5898,N_4296,N_4559);
xnor U5899 (N_5899,N_4428,N_4480);
or U5900 (N_5900,N_4939,N_4657);
and U5901 (N_5901,N_4809,N_4703);
or U5902 (N_5902,N_4896,N_4768);
xnor U5903 (N_5903,N_4014,N_4273);
nand U5904 (N_5904,N_4801,N_4442);
or U5905 (N_5905,N_4671,N_4452);
or U5906 (N_5906,N_4010,N_4026);
xnor U5907 (N_5907,N_4808,N_4654);
or U5908 (N_5908,N_4982,N_4222);
nor U5909 (N_5909,N_4267,N_4132);
nand U5910 (N_5910,N_4152,N_4170);
nand U5911 (N_5911,N_4912,N_4140);
nand U5912 (N_5912,N_4094,N_4755);
xor U5913 (N_5913,N_4166,N_4894);
or U5914 (N_5914,N_4403,N_4896);
and U5915 (N_5915,N_4673,N_4625);
xnor U5916 (N_5916,N_4519,N_4507);
nor U5917 (N_5917,N_4427,N_4500);
xnor U5918 (N_5918,N_4767,N_4377);
or U5919 (N_5919,N_4618,N_4411);
and U5920 (N_5920,N_4474,N_4435);
and U5921 (N_5921,N_4112,N_4243);
xor U5922 (N_5922,N_4204,N_4316);
nand U5923 (N_5923,N_4839,N_4304);
xor U5924 (N_5924,N_4001,N_4122);
or U5925 (N_5925,N_4723,N_4124);
nand U5926 (N_5926,N_4632,N_4669);
or U5927 (N_5927,N_4792,N_4776);
nand U5928 (N_5928,N_4151,N_4032);
xnor U5929 (N_5929,N_4936,N_4344);
nand U5930 (N_5930,N_4855,N_4510);
and U5931 (N_5931,N_4573,N_4377);
nand U5932 (N_5932,N_4646,N_4140);
or U5933 (N_5933,N_4227,N_4388);
nand U5934 (N_5934,N_4782,N_4188);
xor U5935 (N_5935,N_4164,N_4148);
or U5936 (N_5936,N_4991,N_4319);
or U5937 (N_5937,N_4463,N_4899);
and U5938 (N_5938,N_4793,N_4080);
nor U5939 (N_5939,N_4288,N_4945);
xnor U5940 (N_5940,N_4483,N_4643);
nand U5941 (N_5941,N_4344,N_4734);
xnor U5942 (N_5942,N_4704,N_4679);
nor U5943 (N_5943,N_4578,N_4106);
nand U5944 (N_5944,N_4771,N_4600);
nand U5945 (N_5945,N_4250,N_4840);
nor U5946 (N_5946,N_4339,N_4622);
or U5947 (N_5947,N_4744,N_4661);
xnor U5948 (N_5948,N_4987,N_4873);
nand U5949 (N_5949,N_4549,N_4319);
nand U5950 (N_5950,N_4678,N_4977);
xor U5951 (N_5951,N_4286,N_4543);
or U5952 (N_5952,N_4184,N_4248);
or U5953 (N_5953,N_4347,N_4367);
xnor U5954 (N_5954,N_4172,N_4366);
or U5955 (N_5955,N_4959,N_4269);
and U5956 (N_5956,N_4110,N_4919);
and U5957 (N_5957,N_4496,N_4888);
nor U5958 (N_5958,N_4793,N_4382);
nand U5959 (N_5959,N_4504,N_4616);
xnor U5960 (N_5960,N_4675,N_4012);
or U5961 (N_5961,N_4004,N_4397);
and U5962 (N_5962,N_4836,N_4055);
xor U5963 (N_5963,N_4906,N_4597);
xor U5964 (N_5964,N_4500,N_4128);
nand U5965 (N_5965,N_4176,N_4683);
and U5966 (N_5966,N_4268,N_4726);
and U5967 (N_5967,N_4992,N_4914);
xnor U5968 (N_5968,N_4749,N_4672);
or U5969 (N_5969,N_4781,N_4102);
and U5970 (N_5970,N_4759,N_4969);
nand U5971 (N_5971,N_4880,N_4321);
xnor U5972 (N_5972,N_4769,N_4545);
xor U5973 (N_5973,N_4377,N_4116);
nand U5974 (N_5974,N_4101,N_4334);
nor U5975 (N_5975,N_4939,N_4852);
nor U5976 (N_5976,N_4148,N_4185);
and U5977 (N_5977,N_4532,N_4201);
nand U5978 (N_5978,N_4411,N_4912);
and U5979 (N_5979,N_4302,N_4627);
or U5980 (N_5980,N_4899,N_4412);
nand U5981 (N_5981,N_4780,N_4634);
or U5982 (N_5982,N_4457,N_4387);
nand U5983 (N_5983,N_4319,N_4398);
xor U5984 (N_5984,N_4669,N_4232);
nand U5985 (N_5985,N_4796,N_4164);
nand U5986 (N_5986,N_4949,N_4870);
or U5987 (N_5987,N_4397,N_4281);
nor U5988 (N_5988,N_4423,N_4331);
or U5989 (N_5989,N_4016,N_4246);
or U5990 (N_5990,N_4639,N_4067);
or U5991 (N_5991,N_4027,N_4399);
and U5992 (N_5992,N_4268,N_4098);
xor U5993 (N_5993,N_4448,N_4057);
or U5994 (N_5994,N_4650,N_4721);
and U5995 (N_5995,N_4602,N_4255);
nand U5996 (N_5996,N_4727,N_4640);
or U5997 (N_5997,N_4714,N_4174);
or U5998 (N_5998,N_4946,N_4328);
xnor U5999 (N_5999,N_4140,N_4546);
or U6000 (N_6000,N_5981,N_5234);
xnor U6001 (N_6001,N_5236,N_5156);
or U6002 (N_6002,N_5283,N_5772);
and U6003 (N_6003,N_5763,N_5690);
or U6004 (N_6004,N_5363,N_5972);
nor U6005 (N_6005,N_5113,N_5200);
nand U6006 (N_6006,N_5189,N_5872);
or U6007 (N_6007,N_5180,N_5678);
or U6008 (N_6008,N_5030,N_5616);
xnor U6009 (N_6009,N_5639,N_5734);
xnor U6010 (N_6010,N_5093,N_5530);
nand U6011 (N_6011,N_5099,N_5259);
nand U6012 (N_6012,N_5911,N_5759);
or U6013 (N_6013,N_5367,N_5455);
or U6014 (N_6014,N_5342,N_5277);
nor U6015 (N_6015,N_5798,N_5097);
and U6016 (N_6016,N_5661,N_5577);
or U6017 (N_6017,N_5288,N_5468);
and U6018 (N_6018,N_5773,N_5496);
or U6019 (N_6019,N_5660,N_5703);
nor U6020 (N_6020,N_5243,N_5725);
nor U6021 (N_6021,N_5306,N_5008);
xnor U6022 (N_6022,N_5434,N_5887);
xor U6023 (N_6023,N_5810,N_5522);
nand U6024 (N_6024,N_5818,N_5158);
xor U6025 (N_6025,N_5094,N_5088);
xnor U6026 (N_6026,N_5405,N_5428);
and U6027 (N_6027,N_5697,N_5276);
and U6028 (N_6028,N_5321,N_5744);
nand U6029 (N_6029,N_5217,N_5326);
nor U6030 (N_6030,N_5543,N_5664);
nor U6031 (N_6031,N_5412,N_5054);
nor U6032 (N_6032,N_5635,N_5935);
nand U6033 (N_6033,N_5868,N_5318);
or U6034 (N_6034,N_5401,N_5470);
nor U6035 (N_6035,N_5372,N_5481);
nor U6036 (N_6036,N_5732,N_5501);
nor U6037 (N_6037,N_5375,N_5369);
and U6038 (N_6038,N_5056,N_5513);
and U6039 (N_6039,N_5881,N_5139);
nor U6040 (N_6040,N_5124,N_5349);
or U6041 (N_6041,N_5615,N_5399);
xnor U6042 (N_6042,N_5076,N_5392);
nand U6043 (N_6043,N_5979,N_5644);
or U6044 (N_6044,N_5589,N_5676);
nor U6045 (N_6045,N_5581,N_5339);
nor U6046 (N_6046,N_5982,N_5044);
nand U6047 (N_6047,N_5737,N_5782);
nor U6048 (N_6048,N_5413,N_5694);
and U6049 (N_6049,N_5835,N_5880);
nand U6050 (N_6050,N_5939,N_5209);
and U6051 (N_6051,N_5319,N_5366);
or U6052 (N_6052,N_5724,N_5707);
nand U6053 (N_6053,N_5202,N_5147);
xnor U6054 (N_6054,N_5790,N_5927);
and U6055 (N_6055,N_5518,N_5580);
xor U6056 (N_6056,N_5842,N_5439);
or U6057 (N_6057,N_5805,N_5447);
xor U6058 (N_6058,N_5251,N_5996);
and U6059 (N_6059,N_5316,N_5203);
xor U6060 (N_6060,N_5086,N_5229);
nand U6061 (N_6061,N_5856,N_5018);
nand U6062 (N_6062,N_5774,N_5134);
nor U6063 (N_6063,N_5072,N_5095);
or U6064 (N_6064,N_5371,N_5081);
nand U6065 (N_6065,N_5809,N_5874);
or U6066 (N_6066,N_5264,N_5598);
or U6067 (N_6067,N_5652,N_5869);
and U6068 (N_6068,N_5188,N_5378);
nand U6069 (N_6069,N_5552,N_5531);
nand U6070 (N_6070,N_5228,N_5951);
nand U6071 (N_6071,N_5914,N_5353);
and U6072 (N_6072,N_5899,N_5999);
and U6073 (N_6073,N_5104,N_5721);
nor U6074 (N_6074,N_5106,N_5947);
nand U6075 (N_6075,N_5022,N_5706);
nor U6076 (N_6076,N_5799,N_5222);
or U6077 (N_6077,N_5923,N_5685);
and U6078 (N_6078,N_5421,N_5519);
nor U6079 (N_6079,N_5383,N_5298);
xor U6080 (N_6080,N_5900,N_5073);
nand U6081 (N_6081,N_5904,N_5829);
xor U6082 (N_6082,N_5016,N_5688);
nand U6083 (N_6083,N_5764,N_5704);
nor U6084 (N_6084,N_5400,N_5360);
xor U6085 (N_6085,N_5131,N_5994);
and U6086 (N_6086,N_5558,N_5140);
nand U6087 (N_6087,N_5407,N_5323);
xor U6088 (N_6088,N_5021,N_5064);
and U6089 (N_6089,N_5959,N_5731);
nor U6090 (N_6090,N_5687,N_5791);
xnor U6091 (N_6091,N_5517,N_5756);
xor U6092 (N_6092,N_5625,N_5789);
or U6093 (N_6093,N_5191,N_5520);
and U6094 (N_6094,N_5100,N_5491);
nand U6095 (N_6095,N_5172,N_5962);
nor U6096 (N_6096,N_5847,N_5309);
xor U6097 (N_6097,N_5343,N_5453);
xnor U6098 (N_6098,N_5740,N_5257);
nor U6099 (N_6099,N_5148,N_5406);
nor U6100 (N_6100,N_5898,N_5928);
and U6101 (N_6101,N_5057,N_5459);
and U6102 (N_6102,N_5844,N_5278);
and U6103 (N_6103,N_5307,N_5565);
nor U6104 (N_6104,N_5142,N_5219);
nand U6105 (N_6105,N_5152,N_5634);
nor U6106 (N_6106,N_5071,N_5215);
nand U6107 (N_6107,N_5049,N_5542);
nor U6108 (N_6108,N_5454,N_5702);
nor U6109 (N_6109,N_5235,N_5166);
or U6110 (N_6110,N_5467,N_5777);
or U6111 (N_6111,N_5848,N_5084);
and U6112 (N_6112,N_5608,N_5955);
nand U6113 (N_6113,N_5225,N_5752);
nor U6114 (N_6114,N_5083,N_5750);
or U6115 (N_6115,N_5233,N_5877);
and U6116 (N_6116,N_5793,N_5977);
nor U6117 (N_6117,N_5444,N_5862);
nand U6118 (N_6118,N_5282,N_5313);
nor U6119 (N_6119,N_5133,N_5260);
nand U6120 (N_6120,N_5328,N_5013);
and U6121 (N_6121,N_5286,N_5143);
nand U6122 (N_6122,N_5418,N_5490);
nor U6123 (N_6123,N_5419,N_5729);
or U6124 (N_6124,N_5301,N_5079);
or U6125 (N_6125,N_5843,N_5956);
nor U6126 (N_6126,N_5859,N_5250);
nand U6127 (N_6127,N_5595,N_5273);
and U6128 (N_6128,N_5157,N_5484);
nor U6129 (N_6129,N_5550,N_5146);
nand U6130 (N_6130,N_5443,N_5770);
and U6131 (N_6131,N_5866,N_5695);
or U6132 (N_6132,N_5429,N_5967);
nor U6133 (N_6133,N_5457,N_5508);
or U6134 (N_6134,N_5480,N_5244);
xnor U6135 (N_6135,N_5091,N_5776);
and U6136 (N_6136,N_5003,N_5575);
nor U6137 (N_6137,N_5514,N_5510);
or U6138 (N_6138,N_5918,N_5446);
nand U6139 (N_6139,N_5493,N_5155);
xor U6140 (N_6140,N_5034,N_5998);
and U6141 (N_6141,N_5512,N_5162);
nand U6142 (N_6142,N_5631,N_5934);
xor U6143 (N_6143,N_5677,N_5322);
or U6144 (N_6144,N_5980,N_5292);
and U6145 (N_6145,N_5875,N_5332);
or U6146 (N_6146,N_5930,N_5945);
nand U6147 (N_6147,N_5127,N_5701);
nor U6148 (N_6148,N_5983,N_5314);
nand U6149 (N_6149,N_5135,N_5674);
xor U6150 (N_6150,N_5495,N_5267);
or U6151 (N_6151,N_5386,N_5043);
nand U6152 (N_6152,N_5297,N_5252);
and U6153 (N_6153,N_5103,N_5573);
nor U6154 (N_6154,N_5402,N_5964);
or U6155 (N_6155,N_5111,N_5170);
or U6156 (N_6156,N_5730,N_5938);
nand U6157 (N_6157,N_5673,N_5836);
nand U6158 (N_6158,N_5272,N_5061);
xor U6159 (N_6159,N_5028,N_5940);
or U6160 (N_6160,N_5352,N_5985);
nand U6161 (N_6161,N_5715,N_5171);
nand U6162 (N_6162,N_5141,N_5201);
and U6163 (N_6163,N_5090,N_5990);
and U6164 (N_6164,N_5416,N_5845);
or U6165 (N_6165,N_5640,N_5775);
and U6166 (N_6166,N_5409,N_5485);
or U6167 (N_6167,N_5237,N_5831);
nand U6168 (N_6168,N_5821,N_5672);
nand U6169 (N_6169,N_5153,N_5144);
nor U6170 (N_6170,N_5867,N_5966);
xnor U6171 (N_6171,N_5190,N_5341);
xnor U6172 (N_6172,N_5958,N_5816);
nand U6173 (N_6173,N_5345,N_5394);
nand U6174 (N_6174,N_5193,N_5710);
or U6175 (N_6175,N_5840,N_5693);
or U6176 (N_6176,N_5922,N_5174);
and U6177 (N_6177,N_5108,N_5572);
and U6178 (N_6178,N_5539,N_5115);
and U6179 (N_6179,N_5813,N_5364);
and U6180 (N_6180,N_5596,N_5340);
and U6181 (N_6181,N_5834,N_5683);
nor U6182 (N_6182,N_5936,N_5850);
and U6183 (N_6183,N_5971,N_5526);
and U6184 (N_6184,N_5554,N_5746);
and U6185 (N_6185,N_5311,N_5507);
or U6186 (N_6186,N_5965,N_5077);
and U6187 (N_6187,N_5886,N_5211);
nor U6188 (N_6188,N_5380,N_5637);
nand U6189 (N_6189,N_5643,N_5449);
nor U6190 (N_6190,N_5164,N_5795);
nor U6191 (N_6191,N_5646,N_5827);
nand U6192 (N_6192,N_5524,N_5536);
or U6193 (N_6193,N_5270,N_5390);
or U6194 (N_6194,N_5240,N_5778);
xor U6195 (N_6195,N_5261,N_5611);
xor U6196 (N_6196,N_5080,N_5442);
nor U6197 (N_6197,N_5648,N_5258);
xor U6198 (N_6198,N_5659,N_5448);
nand U6199 (N_6199,N_5151,N_5293);
nor U6200 (N_6200,N_5186,N_5224);
nand U6201 (N_6201,N_5102,N_5503);
xor U6202 (N_6202,N_5395,N_5838);
nor U6203 (N_6203,N_5864,N_5205);
xnor U6204 (N_6204,N_5132,N_5888);
xnor U6205 (N_6205,N_5576,N_5279);
nand U6206 (N_6206,N_5599,N_5903);
xor U6207 (N_6207,N_5749,N_5296);
and U6208 (N_6208,N_5876,N_5336);
and U6209 (N_6209,N_5976,N_5338);
and U6210 (N_6210,N_5846,N_5492);
nand U6211 (N_6211,N_5780,N_5743);
nand U6212 (N_6212,N_5570,N_5535);
or U6213 (N_6213,N_5566,N_5074);
nand U6214 (N_6214,N_5559,N_5105);
or U6215 (N_6215,N_5063,N_5089);
nor U6216 (N_6216,N_5398,N_5689);
or U6217 (N_6217,N_5545,N_5471);
nor U6218 (N_6218,N_5437,N_5871);
nand U6219 (N_6219,N_5050,N_5195);
or U6220 (N_6220,N_5450,N_5046);
nand U6221 (N_6221,N_5065,N_5751);
and U6222 (N_6222,N_5878,N_5067);
nand U6223 (N_6223,N_5389,N_5001);
nor U6224 (N_6224,N_5256,N_5109);
xor U6225 (N_6225,N_5808,N_5404);
or U6226 (N_6226,N_5606,N_5494);
xnor U6227 (N_6227,N_5424,N_5933);
xor U6228 (N_6228,N_5671,N_5331);
or U6229 (N_6229,N_5642,N_5445);
nand U6230 (N_6230,N_5950,N_5879);
nand U6231 (N_6231,N_5187,N_5804);
nand U6232 (N_6232,N_5137,N_5223);
and U6233 (N_6233,N_5308,N_5946);
nand U6234 (N_6234,N_5691,N_5628);
and U6235 (N_6235,N_5742,N_5489);
nand U6236 (N_6236,N_5220,N_5912);
nand U6237 (N_6237,N_5285,N_5663);
nor U6238 (N_6238,N_5511,N_5477);
or U6239 (N_6239,N_5833,N_5609);
nor U6240 (N_6240,N_5023,N_5629);
nand U6241 (N_6241,N_5783,N_5905);
or U6242 (N_6242,N_5852,N_5801);
and U6243 (N_6243,N_5368,N_5408);
nor U6244 (N_6244,N_5052,N_5374);
nor U6245 (N_6245,N_5832,N_5909);
nand U6246 (N_6246,N_5692,N_5226);
nand U6247 (N_6247,N_5126,N_5465);
xor U6248 (N_6248,N_5433,N_5123);
nor U6249 (N_6249,N_5587,N_5654);
or U6250 (N_6250,N_5183,N_5529);
nand U6251 (N_6251,N_5410,N_5117);
xor U6252 (N_6252,N_5423,N_5622);
xor U6253 (N_6253,N_5555,N_5841);
or U6254 (N_6254,N_5921,N_5620);
nand U6255 (N_6255,N_5767,N_5107);
xor U6256 (N_6256,N_5662,N_5348);
or U6257 (N_6257,N_5942,N_5861);
nand U6258 (N_6258,N_5145,N_5865);
xnor U6259 (N_6259,N_5765,N_5361);
or U6260 (N_6260,N_5325,N_5883);
nand U6261 (N_6261,N_5451,N_5020);
or U6262 (N_6262,N_5739,N_5828);
xor U6263 (N_6263,N_5178,N_5379);
or U6264 (N_6264,N_5588,N_5993);
nand U6265 (N_6265,N_5525,N_5557);
nand U6266 (N_6266,N_5009,N_5357);
and U6267 (N_6267,N_5249,N_5087);
nor U6268 (N_6268,N_5870,N_5463);
nor U6269 (N_6269,N_5114,N_5185);
nand U6270 (N_6270,N_5456,N_5974);
nor U6271 (N_6271,N_5638,N_5562);
xnor U6272 (N_6272,N_5907,N_5438);
or U6273 (N_6273,N_5925,N_5128);
and U6274 (N_6274,N_5610,N_5591);
nand U6275 (N_6275,N_5995,N_5122);
or U6276 (N_6276,N_5024,N_5992);
or U6277 (N_6277,N_5414,N_5823);
and U6278 (N_6278,N_5027,N_5641);
nand U6279 (N_6279,N_5381,N_5159);
nor U6280 (N_6280,N_5239,N_5556);
or U6281 (N_6281,N_5953,N_5210);
nor U6282 (N_6282,N_5506,N_5800);
or U6283 (N_6283,N_5462,N_5890);
and U6284 (N_6284,N_5284,N_5594);
nor U6285 (N_6285,N_5294,N_5365);
and U6286 (N_6286,N_5165,N_5901);
xnor U6287 (N_6287,N_5602,N_5315);
nor U6288 (N_6288,N_5411,N_5991);
and U6289 (N_6289,N_5712,N_5769);
xor U6290 (N_6290,N_5475,N_5649);
xor U6291 (N_6291,N_5048,N_5658);
nand U6292 (N_6292,N_5384,N_5047);
nand U6293 (N_6293,N_5943,N_5670);
nor U6294 (N_6294,N_5177,N_5055);
or U6295 (N_6295,N_5247,N_5680);
or U6296 (N_6296,N_5902,N_5125);
or U6297 (N_6297,N_5548,N_5310);
nor U6298 (N_6298,N_5726,N_5426);
or U6299 (N_6299,N_5889,N_5120);
nand U6300 (N_6300,N_5632,N_5618);
and U6301 (N_6301,N_5483,N_5619);
nor U6302 (N_6302,N_5388,N_5207);
nand U6303 (N_6303,N_5216,N_5295);
xor U6304 (N_6304,N_5913,N_5385);
nand U6305 (N_6305,N_5154,N_5041);
and U6306 (N_6306,N_5425,N_5245);
and U6307 (N_6307,N_5929,N_5657);
nor U6308 (N_6308,N_5987,N_5698);
or U6309 (N_6309,N_5708,N_5858);
and U6310 (N_6310,N_5238,N_5350);
nor U6311 (N_6311,N_5906,N_5521);
and U6312 (N_6312,N_5837,N_5498);
or U6313 (N_6313,N_5544,N_5747);
nand U6314 (N_6314,N_5553,N_5184);
or U6315 (N_6315,N_5949,N_5705);
xnor U6316 (N_6316,N_5176,N_5377);
nor U6317 (N_6317,N_5299,N_5417);
xor U6318 (N_6318,N_5231,N_5317);
nor U6319 (N_6319,N_5329,N_5478);
nor U6320 (N_6320,N_5253,N_5578);
xnor U6321 (N_6321,N_5717,N_5568);
xor U6322 (N_6322,N_5075,N_5458);
nor U6323 (N_6323,N_5356,N_5957);
xor U6324 (N_6324,N_5007,N_5917);
nand U6325 (N_6325,N_5391,N_5716);
and U6326 (N_6326,N_5825,N_5011);
and U6327 (N_6327,N_5579,N_5476);
xor U6328 (N_6328,N_5300,N_5466);
or U6329 (N_6329,N_5666,N_5582);
nor U6330 (N_6330,N_5645,N_5452);
or U6331 (N_6331,N_5005,N_5713);
nor U6332 (N_6332,N_5714,N_5460);
and U6333 (N_6333,N_5312,N_5085);
xor U6334 (N_6334,N_5000,N_5359);
and U6335 (N_6335,N_5968,N_5647);
and U6336 (N_6336,N_5370,N_5474);
nor U6337 (N_6337,N_5305,N_5741);
xor U6338 (N_6338,N_5497,N_5214);
xnor U6339 (N_6339,N_5121,N_5811);
nor U6340 (N_6340,N_5802,N_5192);
nor U6341 (N_6341,N_5129,N_5334);
or U6342 (N_6342,N_5196,N_5160);
or U6343 (N_6343,N_5179,N_5118);
and U6344 (N_6344,N_5266,N_5910);
nor U6345 (N_6345,N_5788,N_5597);
nand U6346 (N_6346,N_5627,N_5042);
nor U6347 (N_6347,N_5039,N_5528);
and U6348 (N_6348,N_5605,N_5723);
nor U6349 (N_6349,N_5792,N_5150);
or U6350 (N_6350,N_5330,N_5019);
and U6351 (N_6351,N_5839,N_5337);
and U6352 (N_6352,N_5218,N_5797);
nand U6353 (N_6353,N_5516,N_5393);
or U6354 (N_6354,N_5614,N_5853);
nand U6355 (N_6355,N_5346,N_5537);
xnor U6356 (N_6356,N_5561,N_5116);
or U6357 (N_6357,N_5194,N_5601);
nor U6358 (N_6358,N_5623,N_5937);
or U6359 (N_6359,N_5822,N_5675);
nand U6360 (N_6360,N_5268,N_5563);
and U6361 (N_6361,N_5633,N_5699);
xnor U6362 (N_6362,N_5255,N_5718);
nor U6363 (N_6363,N_5978,N_5504);
xor U6364 (N_6364,N_5882,N_5803);
nor U6365 (N_6365,N_5590,N_5854);
xor U6366 (N_6366,N_5376,N_5230);
nor U6367 (N_6367,N_5096,N_5851);
nand U6368 (N_6368,N_5058,N_5895);
xor U6369 (N_6369,N_5213,N_5785);
nand U6370 (N_6370,N_5894,N_5029);
or U6371 (N_6371,N_5728,N_5893);
nand U6372 (N_6372,N_5500,N_5280);
and U6373 (N_6373,N_5373,N_5897);
xnor U6374 (N_6374,N_5422,N_5527);
xor U6375 (N_6375,N_5035,N_5208);
or U6376 (N_6376,N_5062,N_5168);
or U6377 (N_6377,N_5271,N_5066);
nor U6378 (N_6378,N_5650,N_5396);
xnor U6379 (N_6379,N_5138,N_5092);
or U6380 (N_6380,N_5430,N_5748);
nand U6381 (N_6381,N_5669,N_5733);
nand U6382 (N_6382,N_5397,N_5970);
nand U6383 (N_6383,N_5932,N_5204);
xor U6384 (N_6384,N_5040,N_5078);
and U6385 (N_6385,N_5681,N_5173);
and U6386 (N_6386,N_5855,N_5988);
or U6387 (N_6387,N_5546,N_5163);
xor U6388 (N_6388,N_5771,N_5857);
nor U6389 (N_6389,N_5781,N_5863);
nand U6390 (N_6390,N_5014,N_5119);
and U6391 (N_6391,N_5549,N_5161);
xnor U6392 (N_6392,N_5098,N_5358);
nand U6393 (N_6393,N_5432,N_5636);
xor U6394 (N_6394,N_5753,N_5651);
nand U6395 (N_6395,N_5344,N_5586);
nor U6396 (N_6396,N_5473,N_5761);
nor U6397 (N_6397,N_5564,N_5817);
or U6398 (N_6398,N_5320,N_5915);
and U6399 (N_6399,N_5482,N_5051);
nor U6400 (N_6400,N_5427,N_5354);
nand U6401 (N_6401,N_5025,N_5711);
and U6402 (N_6402,N_5656,N_5860);
nor U6403 (N_6403,N_5515,N_5626);
and U6404 (N_6404,N_5924,N_5045);
nand U6405 (N_6405,N_5505,N_5824);
nor U6406 (N_6406,N_5002,N_5262);
nand U6407 (N_6407,N_5873,N_5420);
and U6408 (N_6408,N_5963,N_5812);
nand U6409 (N_6409,N_5436,N_5274);
and U6410 (N_6410,N_5944,N_5952);
nand U6411 (N_6411,N_5585,N_5415);
or U6412 (N_6412,N_5206,N_5973);
and U6413 (N_6413,N_5440,N_5403);
or U6414 (N_6414,N_5607,N_5031);
xnor U6415 (N_6415,N_5149,N_5613);
nand U6416 (N_6416,N_5068,N_5069);
xnor U6417 (N_6417,N_5571,N_5441);
and U6418 (N_6418,N_5291,N_5032);
nand U6419 (N_6419,N_5461,N_5469);
nand U6420 (N_6420,N_5668,N_5181);
or U6421 (N_6421,N_5722,N_5700);
or U6422 (N_6422,N_5665,N_5303);
xor U6423 (N_6423,N_5603,N_5199);
xor U6424 (N_6424,N_5479,N_5324);
and U6425 (N_6425,N_5806,N_5975);
or U6426 (N_6426,N_5532,N_5534);
nor U6427 (N_6427,N_5584,N_5241);
nor U6428 (N_6428,N_5169,N_5221);
or U6429 (N_6429,N_5604,N_5538);
and U6430 (N_6430,N_5768,N_5621);
and U6431 (N_6431,N_5896,N_5017);
or U6432 (N_6432,N_5541,N_5814);
nand U6433 (N_6433,N_5026,N_5004);
nor U6434 (N_6434,N_5038,N_5060);
or U6435 (N_6435,N_5488,N_5254);
and U6436 (N_6436,N_5709,N_5754);
and U6437 (N_6437,N_5997,N_5112);
and U6438 (N_6438,N_5036,N_5757);
nor U6439 (N_6439,N_5919,N_5736);
or U6440 (N_6440,N_5612,N_5263);
or U6441 (N_6441,N_5807,N_5053);
nor U6442 (N_6442,N_5265,N_5684);
nand U6443 (N_6443,N_5275,N_5540);
nor U6444 (N_6444,N_5227,N_5015);
and U6445 (N_6445,N_5986,N_5486);
xnor U6446 (N_6446,N_5762,N_5755);
and U6447 (N_6447,N_5281,N_5033);
nor U6448 (N_6448,N_5667,N_5686);
or U6449 (N_6449,N_5600,N_5327);
nor U6450 (N_6450,N_5891,N_5787);
nand U6451 (N_6451,N_5735,N_5760);
nand U6452 (N_6452,N_5849,N_5198);
and U6453 (N_6453,N_5796,N_5786);
and U6454 (N_6454,N_5246,N_5130);
nand U6455 (N_6455,N_5961,N_5302);
xnor U6456 (N_6456,N_5569,N_5885);
and U6457 (N_6457,N_5779,N_5989);
nor U6458 (N_6458,N_5269,N_5830);
xnor U6459 (N_6459,N_5387,N_5719);
and U6460 (N_6460,N_5070,N_5289);
and U6461 (N_6461,N_5931,N_5533);
and U6462 (N_6462,N_5010,N_5304);
or U6463 (N_6463,N_5037,N_5745);
or U6464 (N_6464,N_5232,N_5758);
nor U6465 (N_6465,N_5509,N_5820);
or U6466 (N_6466,N_5720,N_5012);
nand U6467 (N_6467,N_5197,N_5560);
nand U6468 (N_6468,N_5347,N_5136);
and U6469 (N_6469,N_5382,N_5523);
and U6470 (N_6470,N_5653,N_5617);
and U6471 (N_6471,N_5547,N_5592);
nor U6472 (N_6472,N_5794,N_5248);
and U6473 (N_6473,N_5815,N_5487);
nand U6474 (N_6474,N_5593,N_5916);
nor U6475 (N_6475,N_5624,N_5499);
nor U6476 (N_6476,N_5472,N_5941);
xor U6477 (N_6477,N_5175,N_5926);
and U6478 (N_6478,N_5287,N_5355);
or U6479 (N_6479,N_5006,N_5908);
and U6480 (N_6480,N_5884,N_5738);
or U6481 (N_6481,N_5630,N_5826);
and U6482 (N_6482,N_5212,N_5101);
or U6483 (N_6483,N_5242,N_5082);
or U6484 (N_6484,N_5551,N_5110);
nand U6485 (N_6485,N_5819,N_5696);
nor U6486 (N_6486,N_5182,N_5920);
xnor U6487 (N_6487,N_5435,N_5960);
nand U6488 (N_6488,N_5335,N_5682);
nor U6489 (N_6489,N_5655,N_5431);
and U6490 (N_6490,N_5892,N_5059);
or U6491 (N_6491,N_5954,N_5567);
nand U6492 (N_6492,N_5167,N_5984);
xnor U6493 (N_6493,N_5784,N_5766);
nand U6494 (N_6494,N_5969,N_5333);
xor U6495 (N_6495,N_5948,N_5502);
and U6496 (N_6496,N_5727,N_5574);
nand U6497 (N_6497,N_5290,N_5583);
and U6498 (N_6498,N_5351,N_5679);
nand U6499 (N_6499,N_5464,N_5362);
nor U6500 (N_6500,N_5490,N_5362);
nand U6501 (N_6501,N_5613,N_5717);
and U6502 (N_6502,N_5728,N_5924);
or U6503 (N_6503,N_5758,N_5455);
or U6504 (N_6504,N_5473,N_5199);
nand U6505 (N_6505,N_5539,N_5849);
or U6506 (N_6506,N_5787,N_5716);
and U6507 (N_6507,N_5527,N_5713);
nand U6508 (N_6508,N_5313,N_5623);
nand U6509 (N_6509,N_5577,N_5495);
and U6510 (N_6510,N_5734,N_5702);
or U6511 (N_6511,N_5364,N_5753);
xnor U6512 (N_6512,N_5731,N_5495);
or U6513 (N_6513,N_5019,N_5160);
or U6514 (N_6514,N_5638,N_5512);
nor U6515 (N_6515,N_5578,N_5553);
xor U6516 (N_6516,N_5704,N_5298);
nand U6517 (N_6517,N_5042,N_5923);
xnor U6518 (N_6518,N_5940,N_5079);
xor U6519 (N_6519,N_5730,N_5364);
nand U6520 (N_6520,N_5228,N_5595);
or U6521 (N_6521,N_5489,N_5354);
and U6522 (N_6522,N_5880,N_5242);
or U6523 (N_6523,N_5689,N_5541);
and U6524 (N_6524,N_5545,N_5883);
and U6525 (N_6525,N_5019,N_5600);
or U6526 (N_6526,N_5134,N_5240);
or U6527 (N_6527,N_5382,N_5305);
nand U6528 (N_6528,N_5591,N_5973);
and U6529 (N_6529,N_5650,N_5655);
and U6530 (N_6530,N_5539,N_5610);
or U6531 (N_6531,N_5168,N_5855);
or U6532 (N_6532,N_5394,N_5343);
nor U6533 (N_6533,N_5865,N_5500);
and U6534 (N_6534,N_5058,N_5931);
and U6535 (N_6535,N_5625,N_5669);
nor U6536 (N_6536,N_5364,N_5980);
xnor U6537 (N_6537,N_5781,N_5579);
xnor U6538 (N_6538,N_5190,N_5947);
nand U6539 (N_6539,N_5956,N_5109);
xnor U6540 (N_6540,N_5048,N_5121);
and U6541 (N_6541,N_5750,N_5491);
xor U6542 (N_6542,N_5567,N_5957);
and U6543 (N_6543,N_5449,N_5743);
nand U6544 (N_6544,N_5185,N_5645);
and U6545 (N_6545,N_5107,N_5422);
or U6546 (N_6546,N_5689,N_5347);
nor U6547 (N_6547,N_5829,N_5512);
nand U6548 (N_6548,N_5457,N_5148);
or U6549 (N_6549,N_5748,N_5571);
or U6550 (N_6550,N_5890,N_5762);
nor U6551 (N_6551,N_5214,N_5621);
or U6552 (N_6552,N_5208,N_5645);
xnor U6553 (N_6553,N_5166,N_5199);
or U6554 (N_6554,N_5266,N_5677);
nand U6555 (N_6555,N_5721,N_5158);
or U6556 (N_6556,N_5859,N_5353);
and U6557 (N_6557,N_5806,N_5171);
nor U6558 (N_6558,N_5003,N_5633);
nor U6559 (N_6559,N_5441,N_5435);
xor U6560 (N_6560,N_5894,N_5131);
and U6561 (N_6561,N_5713,N_5605);
and U6562 (N_6562,N_5246,N_5385);
xor U6563 (N_6563,N_5425,N_5277);
nand U6564 (N_6564,N_5961,N_5772);
xnor U6565 (N_6565,N_5137,N_5457);
nand U6566 (N_6566,N_5003,N_5302);
nor U6567 (N_6567,N_5851,N_5415);
xnor U6568 (N_6568,N_5367,N_5570);
and U6569 (N_6569,N_5275,N_5099);
nor U6570 (N_6570,N_5611,N_5571);
and U6571 (N_6571,N_5087,N_5879);
or U6572 (N_6572,N_5659,N_5874);
nor U6573 (N_6573,N_5812,N_5413);
nand U6574 (N_6574,N_5715,N_5264);
nand U6575 (N_6575,N_5898,N_5145);
xor U6576 (N_6576,N_5392,N_5637);
nand U6577 (N_6577,N_5344,N_5941);
and U6578 (N_6578,N_5190,N_5609);
xnor U6579 (N_6579,N_5158,N_5921);
xnor U6580 (N_6580,N_5120,N_5972);
and U6581 (N_6581,N_5016,N_5047);
and U6582 (N_6582,N_5522,N_5664);
or U6583 (N_6583,N_5322,N_5438);
and U6584 (N_6584,N_5125,N_5600);
xor U6585 (N_6585,N_5246,N_5297);
xnor U6586 (N_6586,N_5414,N_5170);
and U6587 (N_6587,N_5947,N_5729);
nand U6588 (N_6588,N_5410,N_5903);
xor U6589 (N_6589,N_5603,N_5970);
and U6590 (N_6590,N_5539,N_5741);
or U6591 (N_6591,N_5118,N_5507);
nor U6592 (N_6592,N_5820,N_5599);
xnor U6593 (N_6593,N_5789,N_5607);
nand U6594 (N_6594,N_5151,N_5015);
nor U6595 (N_6595,N_5254,N_5375);
nor U6596 (N_6596,N_5105,N_5114);
nand U6597 (N_6597,N_5519,N_5332);
nor U6598 (N_6598,N_5420,N_5558);
nand U6599 (N_6599,N_5178,N_5505);
xnor U6600 (N_6600,N_5289,N_5223);
and U6601 (N_6601,N_5887,N_5391);
or U6602 (N_6602,N_5349,N_5174);
nand U6603 (N_6603,N_5066,N_5608);
nand U6604 (N_6604,N_5924,N_5722);
nand U6605 (N_6605,N_5926,N_5683);
xnor U6606 (N_6606,N_5247,N_5804);
xor U6607 (N_6607,N_5168,N_5064);
nand U6608 (N_6608,N_5059,N_5918);
and U6609 (N_6609,N_5266,N_5091);
or U6610 (N_6610,N_5708,N_5894);
and U6611 (N_6611,N_5681,N_5126);
or U6612 (N_6612,N_5973,N_5890);
nand U6613 (N_6613,N_5604,N_5403);
or U6614 (N_6614,N_5396,N_5193);
nand U6615 (N_6615,N_5003,N_5293);
and U6616 (N_6616,N_5924,N_5742);
nand U6617 (N_6617,N_5775,N_5126);
or U6618 (N_6618,N_5490,N_5667);
nor U6619 (N_6619,N_5471,N_5526);
nor U6620 (N_6620,N_5128,N_5454);
and U6621 (N_6621,N_5970,N_5978);
and U6622 (N_6622,N_5784,N_5255);
nand U6623 (N_6623,N_5843,N_5886);
nand U6624 (N_6624,N_5952,N_5381);
and U6625 (N_6625,N_5797,N_5167);
xor U6626 (N_6626,N_5969,N_5337);
xnor U6627 (N_6627,N_5899,N_5957);
xor U6628 (N_6628,N_5423,N_5559);
and U6629 (N_6629,N_5633,N_5645);
nand U6630 (N_6630,N_5427,N_5861);
nand U6631 (N_6631,N_5918,N_5476);
and U6632 (N_6632,N_5125,N_5417);
and U6633 (N_6633,N_5717,N_5823);
and U6634 (N_6634,N_5392,N_5300);
nand U6635 (N_6635,N_5203,N_5314);
or U6636 (N_6636,N_5827,N_5641);
xor U6637 (N_6637,N_5603,N_5674);
or U6638 (N_6638,N_5421,N_5783);
nand U6639 (N_6639,N_5990,N_5731);
xnor U6640 (N_6640,N_5267,N_5471);
nand U6641 (N_6641,N_5896,N_5314);
nor U6642 (N_6642,N_5228,N_5232);
nor U6643 (N_6643,N_5961,N_5897);
xnor U6644 (N_6644,N_5719,N_5297);
or U6645 (N_6645,N_5856,N_5170);
nor U6646 (N_6646,N_5464,N_5953);
and U6647 (N_6647,N_5639,N_5864);
and U6648 (N_6648,N_5700,N_5766);
and U6649 (N_6649,N_5041,N_5527);
xnor U6650 (N_6650,N_5632,N_5896);
nand U6651 (N_6651,N_5684,N_5653);
nor U6652 (N_6652,N_5705,N_5349);
and U6653 (N_6653,N_5744,N_5375);
xor U6654 (N_6654,N_5255,N_5457);
xor U6655 (N_6655,N_5159,N_5604);
and U6656 (N_6656,N_5648,N_5767);
and U6657 (N_6657,N_5844,N_5967);
nor U6658 (N_6658,N_5435,N_5951);
nand U6659 (N_6659,N_5165,N_5390);
nor U6660 (N_6660,N_5770,N_5156);
nand U6661 (N_6661,N_5185,N_5048);
nor U6662 (N_6662,N_5273,N_5117);
or U6663 (N_6663,N_5028,N_5738);
or U6664 (N_6664,N_5397,N_5859);
nor U6665 (N_6665,N_5950,N_5564);
and U6666 (N_6666,N_5955,N_5154);
nor U6667 (N_6667,N_5025,N_5697);
nand U6668 (N_6668,N_5046,N_5429);
or U6669 (N_6669,N_5196,N_5070);
nand U6670 (N_6670,N_5085,N_5030);
xor U6671 (N_6671,N_5961,N_5679);
xnor U6672 (N_6672,N_5702,N_5233);
xor U6673 (N_6673,N_5080,N_5906);
xor U6674 (N_6674,N_5311,N_5477);
and U6675 (N_6675,N_5743,N_5616);
nand U6676 (N_6676,N_5084,N_5865);
and U6677 (N_6677,N_5347,N_5103);
xor U6678 (N_6678,N_5721,N_5001);
nand U6679 (N_6679,N_5367,N_5023);
nor U6680 (N_6680,N_5339,N_5975);
xor U6681 (N_6681,N_5756,N_5099);
nand U6682 (N_6682,N_5317,N_5917);
xnor U6683 (N_6683,N_5008,N_5620);
or U6684 (N_6684,N_5630,N_5284);
or U6685 (N_6685,N_5389,N_5604);
xnor U6686 (N_6686,N_5331,N_5948);
or U6687 (N_6687,N_5464,N_5891);
and U6688 (N_6688,N_5429,N_5404);
nand U6689 (N_6689,N_5697,N_5786);
nand U6690 (N_6690,N_5092,N_5968);
nand U6691 (N_6691,N_5844,N_5917);
xor U6692 (N_6692,N_5432,N_5634);
xnor U6693 (N_6693,N_5995,N_5190);
and U6694 (N_6694,N_5275,N_5024);
and U6695 (N_6695,N_5961,N_5270);
and U6696 (N_6696,N_5950,N_5937);
nand U6697 (N_6697,N_5538,N_5681);
and U6698 (N_6698,N_5208,N_5067);
xnor U6699 (N_6699,N_5386,N_5286);
and U6700 (N_6700,N_5786,N_5797);
nand U6701 (N_6701,N_5308,N_5804);
nand U6702 (N_6702,N_5706,N_5618);
nand U6703 (N_6703,N_5595,N_5733);
nor U6704 (N_6704,N_5889,N_5851);
nand U6705 (N_6705,N_5681,N_5123);
and U6706 (N_6706,N_5723,N_5516);
xor U6707 (N_6707,N_5708,N_5956);
nand U6708 (N_6708,N_5588,N_5540);
and U6709 (N_6709,N_5847,N_5893);
and U6710 (N_6710,N_5452,N_5068);
nor U6711 (N_6711,N_5781,N_5148);
or U6712 (N_6712,N_5869,N_5911);
and U6713 (N_6713,N_5146,N_5514);
nand U6714 (N_6714,N_5397,N_5061);
and U6715 (N_6715,N_5295,N_5513);
nor U6716 (N_6716,N_5110,N_5332);
nand U6717 (N_6717,N_5175,N_5525);
nor U6718 (N_6718,N_5667,N_5411);
xor U6719 (N_6719,N_5102,N_5328);
nand U6720 (N_6720,N_5046,N_5029);
nand U6721 (N_6721,N_5780,N_5867);
and U6722 (N_6722,N_5457,N_5989);
nand U6723 (N_6723,N_5968,N_5165);
nand U6724 (N_6724,N_5242,N_5501);
or U6725 (N_6725,N_5440,N_5902);
xnor U6726 (N_6726,N_5159,N_5709);
or U6727 (N_6727,N_5164,N_5039);
nor U6728 (N_6728,N_5328,N_5289);
and U6729 (N_6729,N_5632,N_5640);
or U6730 (N_6730,N_5386,N_5774);
or U6731 (N_6731,N_5635,N_5558);
nor U6732 (N_6732,N_5555,N_5560);
or U6733 (N_6733,N_5954,N_5883);
xnor U6734 (N_6734,N_5868,N_5654);
and U6735 (N_6735,N_5234,N_5689);
xor U6736 (N_6736,N_5475,N_5963);
and U6737 (N_6737,N_5545,N_5662);
nor U6738 (N_6738,N_5881,N_5469);
and U6739 (N_6739,N_5711,N_5050);
xnor U6740 (N_6740,N_5432,N_5487);
and U6741 (N_6741,N_5631,N_5751);
and U6742 (N_6742,N_5162,N_5223);
nor U6743 (N_6743,N_5565,N_5718);
xor U6744 (N_6744,N_5929,N_5624);
nor U6745 (N_6745,N_5420,N_5194);
or U6746 (N_6746,N_5099,N_5659);
xnor U6747 (N_6747,N_5868,N_5082);
and U6748 (N_6748,N_5391,N_5362);
nor U6749 (N_6749,N_5259,N_5672);
nor U6750 (N_6750,N_5522,N_5740);
xnor U6751 (N_6751,N_5332,N_5744);
nand U6752 (N_6752,N_5137,N_5081);
and U6753 (N_6753,N_5553,N_5197);
nor U6754 (N_6754,N_5444,N_5975);
nor U6755 (N_6755,N_5948,N_5258);
nor U6756 (N_6756,N_5572,N_5470);
nand U6757 (N_6757,N_5798,N_5039);
and U6758 (N_6758,N_5845,N_5169);
nor U6759 (N_6759,N_5761,N_5141);
or U6760 (N_6760,N_5560,N_5577);
nor U6761 (N_6761,N_5895,N_5950);
nand U6762 (N_6762,N_5465,N_5359);
nor U6763 (N_6763,N_5894,N_5761);
nor U6764 (N_6764,N_5157,N_5239);
and U6765 (N_6765,N_5196,N_5784);
or U6766 (N_6766,N_5560,N_5540);
nand U6767 (N_6767,N_5823,N_5847);
or U6768 (N_6768,N_5478,N_5646);
xor U6769 (N_6769,N_5095,N_5606);
nor U6770 (N_6770,N_5000,N_5348);
or U6771 (N_6771,N_5050,N_5564);
xor U6772 (N_6772,N_5685,N_5961);
nand U6773 (N_6773,N_5035,N_5249);
nor U6774 (N_6774,N_5391,N_5871);
nor U6775 (N_6775,N_5999,N_5584);
nand U6776 (N_6776,N_5688,N_5562);
nor U6777 (N_6777,N_5010,N_5917);
or U6778 (N_6778,N_5366,N_5774);
xor U6779 (N_6779,N_5167,N_5222);
xor U6780 (N_6780,N_5035,N_5504);
xnor U6781 (N_6781,N_5339,N_5475);
or U6782 (N_6782,N_5146,N_5266);
and U6783 (N_6783,N_5964,N_5617);
and U6784 (N_6784,N_5170,N_5283);
nor U6785 (N_6785,N_5528,N_5713);
xnor U6786 (N_6786,N_5253,N_5714);
or U6787 (N_6787,N_5372,N_5345);
and U6788 (N_6788,N_5120,N_5150);
nor U6789 (N_6789,N_5095,N_5537);
or U6790 (N_6790,N_5150,N_5616);
nand U6791 (N_6791,N_5026,N_5348);
and U6792 (N_6792,N_5543,N_5005);
or U6793 (N_6793,N_5269,N_5512);
xor U6794 (N_6794,N_5213,N_5149);
and U6795 (N_6795,N_5544,N_5256);
xnor U6796 (N_6796,N_5092,N_5088);
xnor U6797 (N_6797,N_5343,N_5022);
and U6798 (N_6798,N_5672,N_5588);
nand U6799 (N_6799,N_5360,N_5215);
or U6800 (N_6800,N_5935,N_5835);
or U6801 (N_6801,N_5098,N_5048);
nand U6802 (N_6802,N_5429,N_5494);
and U6803 (N_6803,N_5745,N_5384);
nor U6804 (N_6804,N_5398,N_5637);
nor U6805 (N_6805,N_5662,N_5564);
nand U6806 (N_6806,N_5090,N_5298);
or U6807 (N_6807,N_5851,N_5937);
and U6808 (N_6808,N_5571,N_5551);
or U6809 (N_6809,N_5394,N_5072);
nor U6810 (N_6810,N_5002,N_5733);
and U6811 (N_6811,N_5691,N_5507);
xnor U6812 (N_6812,N_5396,N_5453);
or U6813 (N_6813,N_5636,N_5526);
xor U6814 (N_6814,N_5602,N_5523);
and U6815 (N_6815,N_5389,N_5049);
nor U6816 (N_6816,N_5515,N_5566);
nor U6817 (N_6817,N_5751,N_5581);
nand U6818 (N_6818,N_5703,N_5373);
and U6819 (N_6819,N_5027,N_5600);
xor U6820 (N_6820,N_5698,N_5112);
nor U6821 (N_6821,N_5930,N_5903);
nor U6822 (N_6822,N_5956,N_5032);
or U6823 (N_6823,N_5019,N_5395);
xor U6824 (N_6824,N_5934,N_5035);
xnor U6825 (N_6825,N_5260,N_5044);
nand U6826 (N_6826,N_5658,N_5661);
nor U6827 (N_6827,N_5436,N_5512);
and U6828 (N_6828,N_5801,N_5647);
nand U6829 (N_6829,N_5164,N_5165);
xnor U6830 (N_6830,N_5115,N_5246);
nand U6831 (N_6831,N_5405,N_5649);
nor U6832 (N_6832,N_5516,N_5064);
xnor U6833 (N_6833,N_5093,N_5517);
or U6834 (N_6834,N_5170,N_5348);
xor U6835 (N_6835,N_5653,N_5065);
nand U6836 (N_6836,N_5652,N_5584);
nor U6837 (N_6837,N_5417,N_5664);
xnor U6838 (N_6838,N_5338,N_5249);
or U6839 (N_6839,N_5378,N_5540);
nand U6840 (N_6840,N_5696,N_5465);
xor U6841 (N_6841,N_5635,N_5723);
nor U6842 (N_6842,N_5039,N_5151);
nor U6843 (N_6843,N_5927,N_5118);
xor U6844 (N_6844,N_5916,N_5114);
nand U6845 (N_6845,N_5185,N_5395);
nand U6846 (N_6846,N_5937,N_5521);
and U6847 (N_6847,N_5853,N_5747);
nand U6848 (N_6848,N_5582,N_5500);
nand U6849 (N_6849,N_5798,N_5617);
xor U6850 (N_6850,N_5164,N_5047);
and U6851 (N_6851,N_5792,N_5675);
or U6852 (N_6852,N_5804,N_5362);
xnor U6853 (N_6853,N_5021,N_5295);
or U6854 (N_6854,N_5553,N_5270);
nor U6855 (N_6855,N_5462,N_5114);
nand U6856 (N_6856,N_5246,N_5751);
nand U6857 (N_6857,N_5514,N_5797);
nor U6858 (N_6858,N_5879,N_5974);
nor U6859 (N_6859,N_5664,N_5857);
nand U6860 (N_6860,N_5171,N_5318);
and U6861 (N_6861,N_5160,N_5391);
or U6862 (N_6862,N_5635,N_5161);
or U6863 (N_6863,N_5075,N_5298);
nor U6864 (N_6864,N_5328,N_5907);
nand U6865 (N_6865,N_5473,N_5900);
or U6866 (N_6866,N_5742,N_5331);
and U6867 (N_6867,N_5972,N_5145);
or U6868 (N_6868,N_5736,N_5402);
nor U6869 (N_6869,N_5117,N_5118);
xor U6870 (N_6870,N_5776,N_5643);
xor U6871 (N_6871,N_5884,N_5861);
or U6872 (N_6872,N_5974,N_5517);
and U6873 (N_6873,N_5634,N_5971);
nand U6874 (N_6874,N_5162,N_5917);
nor U6875 (N_6875,N_5738,N_5328);
xor U6876 (N_6876,N_5810,N_5848);
or U6877 (N_6877,N_5592,N_5917);
xnor U6878 (N_6878,N_5287,N_5781);
nand U6879 (N_6879,N_5801,N_5417);
and U6880 (N_6880,N_5112,N_5981);
or U6881 (N_6881,N_5812,N_5271);
nor U6882 (N_6882,N_5494,N_5441);
nand U6883 (N_6883,N_5843,N_5494);
xor U6884 (N_6884,N_5117,N_5532);
nand U6885 (N_6885,N_5298,N_5520);
xor U6886 (N_6886,N_5025,N_5111);
xor U6887 (N_6887,N_5091,N_5276);
nand U6888 (N_6888,N_5231,N_5417);
xor U6889 (N_6889,N_5479,N_5338);
or U6890 (N_6890,N_5994,N_5330);
nor U6891 (N_6891,N_5708,N_5530);
or U6892 (N_6892,N_5791,N_5951);
or U6893 (N_6893,N_5284,N_5865);
nor U6894 (N_6894,N_5684,N_5834);
and U6895 (N_6895,N_5655,N_5640);
and U6896 (N_6896,N_5973,N_5239);
nor U6897 (N_6897,N_5349,N_5578);
or U6898 (N_6898,N_5451,N_5316);
xor U6899 (N_6899,N_5864,N_5997);
nor U6900 (N_6900,N_5043,N_5710);
xnor U6901 (N_6901,N_5966,N_5968);
nand U6902 (N_6902,N_5534,N_5581);
and U6903 (N_6903,N_5505,N_5972);
and U6904 (N_6904,N_5168,N_5837);
nor U6905 (N_6905,N_5362,N_5907);
nand U6906 (N_6906,N_5391,N_5473);
and U6907 (N_6907,N_5363,N_5710);
or U6908 (N_6908,N_5476,N_5877);
or U6909 (N_6909,N_5745,N_5087);
nand U6910 (N_6910,N_5546,N_5993);
and U6911 (N_6911,N_5695,N_5562);
nor U6912 (N_6912,N_5432,N_5183);
nand U6913 (N_6913,N_5864,N_5854);
and U6914 (N_6914,N_5132,N_5118);
xor U6915 (N_6915,N_5062,N_5675);
or U6916 (N_6916,N_5530,N_5816);
nand U6917 (N_6917,N_5573,N_5713);
and U6918 (N_6918,N_5717,N_5877);
or U6919 (N_6919,N_5561,N_5225);
nor U6920 (N_6920,N_5180,N_5162);
or U6921 (N_6921,N_5937,N_5151);
xnor U6922 (N_6922,N_5581,N_5721);
xor U6923 (N_6923,N_5193,N_5483);
nand U6924 (N_6924,N_5463,N_5106);
or U6925 (N_6925,N_5050,N_5567);
nor U6926 (N_6926,N_5323,N_5627);
nor U6927 (N_6927,N_5823,N_5212);
nand U6928 (N_6928,N_5079,N_5809);
nand U6929 (N_6929,N_5466,N_5940);
or U6930 (N_6930,N_5129,N_5689);
or U6931 (N_6931,N_5762,N_5505);
nand U6932 (N_6932,N_5769,N_5775);
xor U6933 (N_6933,N_5943,N_5999);
or U6934 (N_6934,N_5577,N_5971);
xnor U6935 (N_6935,N_5281,N_5920);
and U6936 (N_6936,N_5561,N_5778);
xor U6937 (N_6937,N_5039,N_5693);
nor U6938 (N_6938,N_5123,N_5272);
and U6939 (N_6939,N_5470,N_5404);
and U6940 (N_6940,N_5906,N_5248);
and U6941 (N_6941,N_5655,N_5196);
or U6942 (N_6942,N_5177,N_5964);
xnor U6943 (N_6943,N_5615,N_5589);
and U6944 (N_6944,N_5034,N_5820);
xnor U6945 (N_6945,N_5180,N_5613);
nand U6946 (N_6946,N_5919,N_5867);
nor U6947 (N_6947,N_5643,N_5310);
xnor U6948 (N_6948,N_5810,N_5897);
nor U6949 (N_6949,N_5762,N_5880);
xnor U6950 (N_6950,N_5106,N_5448);
and U6951 (N_6951,N_5199,N_5526);
and U6952 (N_6952,N_5754,N_5914);
xor U6953 (N_6953,N_5511,N_5878);
nor U6954 (N_6954,N_5951,N_5513);
nor U6955 (N_6955,N_5905,N_5274);
and U6956 (N_6956,N_5936,N_5917);
and U6957 (N_6957,N_5812,N_5519);
xor U6958 (N_6958,N_5532,N_5237);
xor U6959 (N_6959,N_5926,N_5229);
and U6960 (N_6960,N_5158,N_5331);
nand U6961 (N_6961,N_5390,N_5440);
nand U6962 (N_6962,N_5330,N_5448);
and U6963 (N_6963,N_5610,N_5781);
nand U6964 (N_6964,N_5615,N_5436);
nor U6965 (N_6965,N_5409,N_5930);
or U6966 (N_6966,N_5937,N_5332);
xnor U6967 (N_6967,N_5333,N_5626);
and U6968 (N_6968,N_5883,N_5132);
nand U6969 (N_6969,N_5344,N_5374);
xor U6970 (N_6970,N_5365,N_5667);
and U6971 (N_6971,N_5524,N_5173);
nand U6972 (N_6972,N_5036,N_5658);
or U6973 (N_6973,N_5535,N_5211);
nand U6974 (N_6974,N_5136,N_5726);
and U6975 (N_6975,N_5935,N_5250);
nand U6976 (N_6976,N_5027,N_5324);
nor U6977 (N_6977,N_5812,N_5815);
nor U6978 (N_6978,N_5685,N_5706);
and U6979 (N_6979,N_5024,N_5096);
nor U6980 (N_6980,N_5778,N_5918);
or U6981 (N_6981,N_5475,N_5274);
or U6982 (N_6982,N_5179,N_5176);
and U6983 (N_6983,N_5890,N_5497);
and U6984 (N_6984,N_5165,N_5125);
nor U6985 (N_6985,N_5908,N_5869);
and U6986 (N_6986,N_5521,N_5728);
nor U6987 (N_6987,N_5885,N_5165);
nor U6988 (N_6988,N_5570,N_5801);
xnor U6989 (N_6989,N_5495,N_5072);
and U6990 (N_6990,N_5574,N_5625);
or U6991 (N_6991,N_5713,N_5254);
and U6992 (N_6992,N_5060,N_5592);
nor U6993 (N_6993,N_5307,N_5900);
and U6994 (N_6994,N_5454,N_5608);
nand U6995 (N_6995,N_5536,N_5921);
and U6996 (N_6996,N_5661,N_5199);
nand U6997 (N_6997,N_5607,N_5060);
nor U6998 (N_6998,N_5564,N_5327);
and U6999 (N_6999,N_5897,N_5947);
xnor U7000 (N_7000,N_6456,N_6748);
nand U7001 (N_7001,N_6611,N_6062);
nor U7002 (N_7002,N_6523,N_6393);
or U7003 (N_7003,N_6047,N_6011);
or U7004 (N_7004,N_6328,N_6213);
nor U7005 (N_7005,N_6740,N_6358);
xor U7006 (N_7006,N_6509,N_6682);
or U7007 (N_7007,N_6940,N_6412);
nand U7008 (N_7008,N_6060,N_6258);
nor U7009 (N_7009,N_6226,N_6561);
or U7010 (N_7010,N_6935,N_6874);
and U7011 (N_7011,N_6096,N_6066);
nor U7012 (N_7012,N_6338,N_6921);
nor U7013 (N_7013,N_6666,N_6477);
and U7014 (N_7014,N_6627,N_6862);
or U7015 (N_7015,N_6608,N_6483);
xor U7016 (N_7016,N_6379,N_6151);
nand U7017 (N_7017,N_6020,N_6661);
xnor U7018 (N_7018,N_6590,N_6339);
or U7019 (N_7019,N_6929,N_6739);
and U7020 (N_7020,N_6735,N_6756);
xnor U7021 (N_7021,N_6606,N_6684);
and U7022 (N_7022,N_6314,N_6922);
nor U7023 (N_7023,N_6734,N_6478);
nand U7024 (N_7024,N_6009,N_6768);
nor U7025 (N_7025,N_6257,N_6090);
nor U7026 (N_7026,N_6521,N_6429);
nand U7027 (N_7027,N_6061,N_6860);
and U7028 (N_7028,N_6941,N_6925);
nor U7029 (N_7029,N_6638,N_6313);
nor U7030 (N_7030,N_6514,N_6037);
or U7031 (N_7031,N_6204,N_6222);
or U7032 (N_7032,N_6091,N_6489);
and U7033 (N_7033,N_6650,N_6100);
and U7034 (N_7034,N_6049,N_6982);
xnor U7035 (N_7035,N_6730,N_6897);
xnor U7036 (N_7036,N_6861,N_6690);
and U7037 (N_7037,N_6882,N_6958);
nand U7038 (N_7038,N_6868,N_6847);
and U7039 (N_7039,N_6769,N_6430);
and U7040 (N_7040,N_6863,N_6946);
xnor U7041 (N_7041,N_6243,N_6828);
or U7042 (N_7042,N_6712,N_6333);
nor U7043 (N_7043,N_6039,N_6557);
and U7044 (N_7044,N_6911,N_6837);
and U7045 (N_7045,N_6706,N_6727);
nand U7046 (N_7046,N_6238,N_6283);
nor U7047 (N_7047,N_6480,N_6779);
or U7048 (N_7048,N_6894,N_6263);
nor U7049 (N_7049,N_6525,N_6449);
nand U7050 (N_7050,N_6033,N_6616);
xnor U7051 (N_7051,N_6629,N_6063);
xnor U7052 (N_7052,N_6494,N_6898);
and U7053 (N_7053,N_6126,N_6369);
or U7054 (N_7054,N_6010,N_6200);
xor U7055 (N_7055,N_6971,N_6174);
nand U7056 (N_7056,N_6366,N_6698);
and U7057 (N_7057,N_6927,N_6839);
nor U7058 (N_7058,N_6107,N_6807);
nor U7059 (N_7059,N_6808,N_6788);
xor U7060 (N_7060,N_6411,N_6830);
xnor U7061 (N_7061,N_6713,N_6256);
xnor U7062 (N_7062,N_6311,N_6332);
and U7063 (N_7063,N_6321,N_6659);
nand U7064 (N_7064,N_6671,N_6424);
nor U7065 (N_7065,N_6645,N_6152);
nand U7066 (N_7066,N_6569,N_6504);
and U7067 (N_7067,N_6915,N_6817);
xor U7068 (N_7068,N_6952,N_6680);
nand U7069 (N_7069,N_6242,N_6092);
nand U7070 (N_7070,N_6545,N_6896);
and U7071 (N_7071,N_6068,N_6065);
xor U7072 (N_7072,N_6472,N_6035);
or U7073 (N_7073,N_6960,N_6133);
nand U7074 (N_7074,N_6121,N_6215);
xnor U7075 (N_7075,N_6932,N_6241);
and U7076 (N_7076,N_6510,N_6754);
and U7077 (N_7077,N_6855,N_6857);
xnor U7078 (N_7078,N_6432,N_6167);
xor U7079 (N_7079,N_6386,N_6655);
nand U7080 (N_7080,N_6284,N_6171);
or U7081 (N_7081,N_6491,N_6440);
and U7082 (N_7082,N_6381,N_6954);
xor U7083 (N_7083,N_6548,N_6324);
or U7084 (N_7084,N_6437,N_6617);
nor U7085 (N_7085,N_6106,N_6064);
nor U7086 (N_7086,N_6715,N_6644);
or U7087 (N_7087,N_6979,N_6452);
nand U7088 (N_7088,N_6672,N_6546);
and U7089 (N_7089,N_6309,N_6775);
and U7090 (N_7090,N_6265,N_6087);
and U7091 (N_7091,N_6205,N_6591);
nand U7092 (N_7092,N_6378,N_6597);
nor U7093 (N_7093,N_6637,N_6741);
or U7094 (N_7094,N_6833,N_6490);
or U7095 (N_7095,N_6155,N_6363);
nand U7096 (N_7096,N_6353,N_6291);
xor U7097 (N_7097,N_6298,N_6574);
nand U7098 (N_7098,N_6325,N_6279);
or U7099 (N_7099,N_6285,N_6781);
xnor U7100 (N_7100,N_6767,N_6850);
and U7101 (N_7101,N_6026,N_6461);
and U7102 (N_7102,N_6813,N_6124);
or U7103 (N_7103,N_6084,N_6519);
nand U7104 (N_7104,N_6917,N_6594);
and U7105 (N_7105,N_6499,N_6919);
or U7106 (N_7106,N_6752,N_6560);
nor U7107 (N_7107,N_6966,N_6446);
xnor U7108 (N_7108,N_6631,N_6914);
nand U7109 (N_7109,N_6145,N_6359);
xor U7110 (N_7110,N_6732,N_6646);
nand U7111 (N_7111,N_6721,N_6602);
and U7112 (N_7112,N_6704,N_6654);
nor U7113 (N_7113,N_6780,N_6007);
nor U7114 (N_7114,N_6433,N_6046);
or U7115 (N_7115,N_6609,N_6178);
nand U7116 (N_7116,N_6231,N_6001);
or U7117 (N_7117,N_6547,N_6635);
or U7118 (N_7118,N_6550,N_6851);
nor U7119 (N_7119,N_6517,N_6259);
or U7120 (N_7120,N_6705,N_6457);
nand U7121 (N_7121,N_6900,N_6697);
or U7122 (N_7122,N_6212,N_6580);
nand U7123 (N_7123,N_6980,N_6108);
nor U7124 (N_7124,N_6392,N_6166);
xor U7125 (N_7125,N_6350,N_6685);
nor U7126 (N_7126,N_6173,N_6190);
and U7127 (N_7127,N_6518,N_6044);
and U7128 (N_7128,N_6239,N_6620);
and U7129 (N_7129,N_6581,N_6370);
or U7130 (N_7130,N_6076,N_6113);
or U7131 (N_7131,N_6636,N_6342);
nor U7132 (N_7132,N_6235,N_6027);
or U7133 (N_7133,N_6567,N_6583);
xor U7134 (N_7134,N_6812,N_6746);
xnor U7135 (N_7135,N_6651,N_6800);
and U7136 (N_7136,N_6251,N_6798);
nor U7137 (N_7137,N_6524,N_6589);
and U7138 (N_7138,N_6928,N_6558);
and U7139 (N_7139,N_6349,N_6199);
nand U7140 (N_7140,N_6520,N_6533);
xnor U7141 (N_7141,N_6649,N_6906);
nand U7142 (N_7142,N_6908,N_6783);
or U7143 (N_7143,N_6832,N_6668);
xor U7144 (N_7144,N_6140,N_6218);
nand U7145 (N_7145,N_6831,N_6623);
nand U7146 (N_7146,N_6972,N_6059);
nand U7147 (N_7147,N_6428,N_6997);
xnor U7148 (N_7148,N_6245,N_6078);
nor U7149 (N_7149,N_6315,N_6431);
nand U7150 (N_7150,N_6612,N_6829);
nor U7151 (N_7151,N_6269,N_6253);
and U7152 (N_7152,N_6120,N_6871);
and U7153 (N_7153,N_6885,N_6738);
xor U7154 (N_7154,N_6728,N_6439);
nor U7155 (N_7155,N_6528,N_6618);
or U7156 (N_7156,N_6080,N_6785);
nand U7157 (N_7157,N_6262,N_6981);
nand U7158 (N_7158,N_6765,N_6395);
nand U7159 (N_7159,N_6968,N_6273);
nand U7160 (N_7160,N_6460,N_6703);
xnor U7161 (N_7161,N_6990,N_6771);
or U7162 (N_7162,N_6067,N_6122);
or U7163 (N_7163,N_6016,N_6289);
xnor U7164 (N_7164,N_6043,N_6916);
nand U7165 (N_7165,N_6965,N_6220);
and U7166 (N_7166,N_6532,N_6913);
nand U7167 (N_7167,N_6694,N_6264);
or U7168 (N_7168,N_6803,N_6744);
nor U7169 (N_7169,N_6209,N_6989);
xor U7170 (N_7170,N_6522,N_6658);
nand U7171 (N_7171,N_6128,N_6942);
and U7172 (N_7172,N_6468,N_6347);
xor U7173 (N_7173,N_6368,N_6938);
nor U7174 (N_7174,N_6419,N_6111);
nor U7175 (N_7175,N_6482,N_6000);
or U7176 (N_7176,N_6867,N_6621);
and U7177 (N_7177,N_6021,N_6400);
nor U7178 (N_7178,N_6642,N_6686);
nor U7179 (N_7179,N_6492,N_6327);
or U7180 (N_7180,N_6986,N_6977);
nor U7181 (N_7181,N_6387,N_6230);
nand U7182 (N_7182,N_6487,N_6710);
nand U7183 (N_7183,N_6041,N_6294);
nand U7184 (N_7184,N_6743,N_6410);
and U7185 (N_7185,N_6474,N_6818);
nand U7186 (N_7186,N_6425,N_6103);
xnor U7187 (N_7187,N_6302,N_6678);
xor U7188 (N_7188,N_6287,N_6409);
and U7189 (N_7189,N_6999,N_6652);
and U7190 (N_7190,N_6605,N_6647);
xor U7191 (N_7191,N_6870,N_6098);
and U7192 (N_7192,N_6054,N_6826);
xnor U7193 (N_7193,N_6513,N_6331);
nor U7194 (N_7194,N_6723,N_6159);
or U7195 (N_7195,N_6607,N_6272);
or U7196 (N_7196,N_6153,N_6516);
nor U7197 (N_7197,N_6290,N_6853);
nand U7198 (N_7198,N_6511,N_6819);
or U7199 (N_7199,N_6232,N_6448);
nor U7200 (N_7200,N_6947,N_6836);
and U7201 (N_7201,N_6416,N_6687);
nor U7202 (N_7202,N_6303,N_6094);
nor U7203 (N_7203,N_6340,N_6210);
xor U7204 (N_7204,N_6714,N_6571);
and U7205 (N_7205,N_6422,N_6604);
xor U7206 (N_7206,N_6471,N_6747);
or U7207 (N_7207,N_6453,N_6426);
or U7208 (N_7208,N_6164,N_6233);
and U7209 (N_7209,N_6790,N_6875);
nand U7210 (N_7210,N_6088,N_6077);
xor U7211 (N_7211,N_6846,N_6268);
nand U7212 (N_7212,N_6130,N_6778);
or U7213 (N_7213,N_6420,N_6329);
xor U7214 (N_7214,N_6013,N_6168);
nor U7215 (N_7215,N_6588,N_6203);
nor U7216 (N_7216,N_6507,N_6444);
and U7217 (N_7217,N_6849,N_6354);
xnor U7218 (N_7218,N_6884,N_6462);
nor U7219 (N_7219,N_6883,N_6967);
and U7220 (N_7220,N_6864,N_6814);
xnor U7221 (N_7221,N_6903,N_6834);
xor U7222 (N_7222,N_6824,N_6282);
nand U7223 (N_7223,N_6249,N_6323);
xnor U7224 (N_7224,N_6475,N_6079);
xnor U7225 (N_7225,N_6751,N_6789);
or U7226 (N_7226,N_6876,N_6689);
xnor U7227 (N_7227,N_6662,N_6719);
and U7228 (N_7228,N_6737,N_6162);
xnor U7229 (N_7229,N_6427,N_6586);
or U7230 (N_7230,N_6148,N_6028);
xnor U7231 (N_7231,N_6726,N_6466);
or U7232 (N_7232,N_6277,N_6699);
or U7233 (N_7233,N_6718,N_6095);
and U7234 (N_7234,N_6415,N_6441);
xor U7235 (N_7235,N_6552,N_6669);
and U7236 (N_7236,N_6074,N_6877);
and U7237 (N_7237,N_6888,N_6809);
xor U7238 (N_7238,N_6539,N_6146);
nand U7239 (N_7239,N_6237,N_6501);
and U7240 (N_7240,N_6530,N_6436);
or U7241 (N_7241,N_6034,N_6592);
nand U7242 (N_7242,N_6464,N_6053);
and U7243 (N_7243,N_6105,N_6673);
and U7244 (N_7244,N_6169,N_6675);
or U7245 (N_7245,N_6144,N_6844);
or U7246 (N_7246,N_6930,N_6840);
nand U7247 (N_7247,N_6086,N_6901);
or U7248 (N_7248,N_6953,N_6984);
or U7249 (N_7249,N_6211,N_6398);
or U7250 (N_7250,N_6700,N_6793);
and U7251 (N_7251,N_6991,N_6810);
nor U7252 (N_7252,N_6307,N_6030);
and U7253 (N_7253,N_6641,N_6936);
nor U7254 (N_7254,N_6599,N_6760);
and U7255 (N_7255,N_6018,N_6795);
xor U7256 (N_7256,N_6656,N_6955);
nand U7257 (N_7257,N_6987,N_6648);
nor U7258 (N_7258,N_6934,N_6485);
nand U7259 (N_7259,N_6562,N_6848);
xor U7260 (N_7260,N_6974,N_6869);
xnor U7261 (N_7261,N_6603,N_6029);
xnor U7262 (N_7262,N_6322,N_6750);
and U7263 (N_7263,N_6051,N_6254);
xor U7264 (N_7264,N_6123,N_6725);
or U7265 (N_7265,N_6383,N_6573);
and U7266 (N_7266,N_6192,N_6318);
and U7267 (N_7267,N_6708,N_6920);
and U7268 (N_7268,N_6390,N_6912);
nor U7269 (N_7269,N_6236,N_6115);
and U7270 (N_7270,N_6676,N_6228);
or U7271 (N_7271,N_6549,N_6188);
and U7272 (N_7272,N_6755,N_6500);
or U7273 (N_7273,N_6216,N_6278);
xnor U7274 (N_7274,N_6119,N_6109);
xnor U7275 (N_7275,N_6172,N_6022);
nor U7276 (N_7276,N_6467,N_6998);
and U7277 (N_7277,N_6380,N_6132);
or U7278 (N_7278,N_6762,N_6255);
and U7279 (N_7279,N_6181,N_6408);
and U7280 (N_7280,N_6615,N_6931);
nand U7281 (N_7281,N_6330,N_6458);
nor U7282 (N_7282,N_6305,N_6266);
nand U7283 (N_7283,N_6702,N_6017);
and U7284 (N_7284,N_6371,N_6841);
nor U7285 (N_7285,N_6292,N_6306);
and U7286 (N_7286,N_6293,N_6729);
nand U7287 (N_7287,N_6250,N_6782);
nand U7288 (N_7288,N_6794,N_6138);
nand U7289 (N_7289,N_6926,N_6886);
nor U7290 (N_7290,N_6820,N_6996);
nand U7291 (N_7291,N_6923,N_6634);
and U7292 (N_7292,N_6014,N_6619);
or U7293 (N_7293,N_6600,N_6568);
xnor U7294 (N_7294,N_6374,N_6455);
xnor U7295 (N_7295,N_6598,N_6512);
and U7296 (N_7296,N_6005,N_6905);
or U7297 (N_7297,N_6413,N_6688);
or U7298 (N_7298,N_6300,N_6023);
and U7299 (N_7299,N_6963,N_6816);
nand U7300 (N_7300,N_6614,N_6731);
nand U7301 (N_7301,N_6799,N_6346);
nand U7302 (N_7302,N_6970,N_6670);
nand U7303 (N_7303,N_6556,N_6206);
nor U7304 (N_7304,N_6842,N_6006);
xnor U7305 (N_7305,N_6918,N_6536);
nand U7306 (N_7306,N_6451,N_6555);
nor U7307 (N_7307,N_6895,N_6459);
and U7308 (N_7308,N_6681,N_6131);
nor U7309 (N_7309,N_6312,N_6160);
and U7310 (N_7310,N_6045,N_6158);
or U7311 (N_7311,N_6101,N_6498);
or U7312 (N_7312,N_6102,N_6057);
nor U7313 (N_7313,N_6667,N_6388);
or U7314 (N_7314,N_6827,N_6949);
nor U7315 (N_7315,N_6048,N_6194);
xor U7316 (N_7316,N_6317,N_6367);
nor U7317 (N_7317,N_6805,N_6075);
and U7318 (N_7318,N_6497,N_6240);
nor U7319 (N_7319,N_6630,N_6773);
xor U7320 (N_7320,N_6529,N_6082);
nor U7321 (N_7321,N_6893,N_6879);
or U7322 (N_7322,N_6985,N_6040);
xor U7323 (N_7323,N_6845,N_6937);
and U7324 (N_7324,N_6657,N_6031);
or U7325 (N_7325,N_6161,N_6450);
nand U7326 (N_7326,N_6653,N_6070);
xor U7327 (N_7327,N_6975,N_6806);
nor U7328 (N_7328,N_6677,N_6632);
or U7329 (N_7329,N_6401,N_6792);
and U7330 (N_7330,N_6357,N_6234);
nor U7331 (N_7331,N_6601,N_6038);
nor U7332 (N_7332,N_6032,N_6149);
or U7333 (N_7333,N_6486,N_6286);
nor U7334 (N_7334,N_6081,N_6186);
and U7335 (N_7335,N_6566,N_6961);
nand U7336 (N_7336,N_6691,N_6180);
or U7337 (N_7337,N_6823,N_6639);
xnor U7338 (N_7338,N_6360,N_6585);
nor U7339 (N_7339,N_6628,N_6973);
xnor U7340 (N_7340,N_6679,N_6247);
nand U7341 (N_7341,N_6304,N_6154);
nor U7342 (N_7342,N_6488,N_6696);
nor U7343 (N_7343,N_6559,N_6904);
nand U7344 (N_7344,N_6469,N_6423);
or U7345 (N_7345,N_6246,N_6711);
and U7346 (N_7346,N_6957,N_6142);
nor U7347 (N_7347,N_6720,N_6320);
or U7348 (N_7348,N_6418,N_6535);
and U7349 (N_7349,N_6177,N_6983);
and U7350 (N_7350,N_6089,N_6008);
and U7351 (N_7351,N_6964,N_6382);
nor U7352 (N_7352,N_6351,N_6992);
or U7353 (N_7353,N_6821,N_6447);
nand U7354 (N_7354,N_6542,N_6165);
or U7355 (N_7355,N_6872,N_6613);
or U7356 (N_7356,N_6856,N_6551);
xor U7357 (N_7357,N_6147,N_6319);
and U7358 (N_7358,N_6036,N_6717);
nand U7359 (N_7359,N_6625,N_6072);
nand U7360 (N_7360,N_6892,N_6626);
or U7361 (N_7361,N_6622,N_6802);
and U7362 (N_7362,N_6344,N_6902);
or U7363 (N_7363,N_6664,N_6110);
nand U7364 (N_7364,N_6179,N_6376);
or U7365 (N_7365,N_6582,N_6252);
nand U7366 (N_7366,N_6384,N_6025);
and U7367 (N_7367,N_6786,N_6660);
and U7368 (N_7368,N_6275,N_6182);
nor U7369 (N_7369,N_6587,N_6407);
or U7370 (N_7370,N_6584,N_6438);
xnor U7371 (N_7371,N_6163,N_6114);
or U7372 (N_7372,N_6099,N_6976);
nand U7373 (N_7373,N_6575,N_6214);
nor U7374 (N_7374,N_6003,N_6310);
xnor U7375 (N_7375,N_6838,N_6024);
or U7376 (N_7376,N_6221,N_6196);
xnor U7377 (N_7377,N_6944,N_6052);
nor U7378 (N_7378,N_6643,N_6707);
nand U7379 (N_7379,N_6337,N_6097);
and U7380 (N_7380,N_6118,N_6508);
and U7381 (N_7381,N_6217,N_6527);
xor U7382 (N_7382,N_6939,N_6742);
nor U7383 (N_7383,N_6207,N_6804);
or U7384 (N_7384,N_6195,N_6276);
and U7385 (N_7385,N_6280,N_6878);
xor U7386 (N_7386,N_6442,N_6825);
nor U7387 (N_7387,N_6633,N_6693);
or U7388 (N_7388,N_6365,N_6175);
nand U7389 (N_7389,N_6399,N_6473);
xor U7390 (N_7390,N_6112,N_6578);
nor U7391 (N_7391,N_6470,N_6336);
nand U7392 (N_7392,N_6722,N_6797);
and U7393 (N_7393,N_6526,N_6537);
and U7394 (N_7394,N_6012,N_6770);
nor U7395 (N_7395,N_6503,N_6610);
and U7396 (N_7396,N_6576,N_6341);
nor U7397 (N_7397,N_6505,N_6881);
xor U7398 (N_7398,N_6889,N_6692);
and U7399 (N_7399,N_6859,N_6201);
nor U7400 (N_7400,N_6766,N_6227);
and U7401 (N_7401,N_6858,N_6579);
nand U7402 (N_7402,N_6377,N_6761);
nand U7403 (N_7403,N_6355,N_6544);
or U7404 (N_7404,N_6184,N_6183);
nand U7405 (N_7405,N_6640,N_6476);
xor U7406 (N_7406,N_6593,N_6297);
or U7407 (N_7407,N_6135,N_6910);
and U7408 (N_7408,N_6811,N_6595);
or U7409 (N_7409,N_6116,N_6443);
and U7410 (N_7410,N_6665,N_6733);
xnor U7411 (N_7411,N_6907,N_6564);
nor U7412 (N_7412,N_6701,N_6695);
nor U7413 (N_7413,N_6758,N_6224);
nand U7414 (N_7414,N_6157,N_6352);
xor U7415 (N_7415,N_6534,N_6141);
or U7416 (N_7416,N_6193,N_6479);
nand U7417 (N_7417,N_6015,N_6801);
xnor U7418 (N_7418,N_6843,N_6299);
or U7419 (N_7419,N_6389,N_6993);
xnor U7420 (N_7420,N_6397,N_6924);
nor U7421 (N_7421,N_6356,N_6865);
and U7422 (N_7422,N_6134,N_6260);
nor U7423 (N_7423,N_6531,N_6073);
or U7424 (N_7424,N_6948,N_6288);
xor U7425 (N_7425,N_6995,N_6434);
nand U7426 (N_7426,N_6002,N_6959);
xor U7427 (N_7427,N_6962,N_6891);
and U7428 (N_7428,N_6301,N_6776);
nor U7429 (N_7429,N_6772,N_6050);
nor U7430 (N_7430,N_6764,N_6267);
and U7431 (N_7431,N_6261,N_6495);
or U7432 (N_7432,N_6663,N_6403);
nand U7433 (N_7433,N_6202,N_6866);
or U7434 (N_7434,N_6815,N_6198);
or U7435 (N_7435,N_6143,N_6085);
or U7436 (N_7436,N_6137,N_6624);
or U7437 (N_7437,N_6326,N_6835);
or U7438 (N_7438,N_6375,N_6136);
and U7439 (N_7439,N_6709,N_6899);
nor U7440 (N_7440,N_6404,N_6270);
or U7441 (N_7441,N_6104,N_6784);
nand U7442 (N_7442,N_6890,N_6056);
and U7443 (N_7443,N_6334,N_6170);
xor U7444 (N_7444,N_6402,N_6873);
xor U7445 (N_7445,N_6553,N_6335);
xnor U7446 (N_7446,N_6308,N_6004);
and U7447 (N_7447,N_6069,N_6796);
or U7448 (N_7448,N_6150,N_6454);
nor U7449 (N_7449,N_6189,N_6345);
and U7450 (N_7450,N_6945,N_6372);
nor U7451 (N_7451,N_6538,N_6348);
nand U7452 (N_7452,N_6093,N_6197);
or U7453 (N_7453,N_6791,N_6125);
nand U7454 (N_7454,N_6343,N_6445);
xor U7455 (N_7455,N_6596,N_6385);
or U7456 (N_7456,N_6570,N_6244);
or U7457 (N_7457,N_6854,N_6055);
or U7458 (N_7458,N_6852,N_6563);
and U7459 (N_7459,N_6435,N_6271);
and U7460 (N_7460,N_6223,N_6745);
nor U7461 (N_7461,N_6724,N_6736);
xor U7462 (N_7462,N_6187,N_6880);
and U7463 (N_7463,N_6019,N_6774);
or U7464 (N_7464,N_6219,N_6281);
nor U7465 (N_7465,N_6208,N_6541);
nor U7466 (N_7466,N_6674,N_6042);
or U7467 (N_7467,N_6496,N_6396);
and U7468 (N_7468,N_6565,N_6943);
and U7469 (N_7469,N_6994,N_6129);
xor U7470 (N_7470,N_6933,N_6951);
nand U7471 (N_7471,N_6361,N_6191);
xor U7472 (N_7472,N_6394,N_6988);
or U7473 (N_7473,N_6083,N_6515);
or U7474 (N_7474,N_6540,N_6417);
nand U7475 (N_7475,N_6777,N_6683);
nor U7476 (N_7476,N_6296,N_6978);
xnor U7477 (N_7477,N_6716,N_6139);
or U7478 (N_7478,N_6543,N_6493);
xnor U7479 (N_7479,N_6909,N_6391);
xor U7480 (N_7480,N_6887,N_6117);
nor U7481 (N_7481,N_6421,N_6414);
nor U7482 (N_7482,N_6406,N_6364);
or U7483 (N_7483,N_6753,N_6127);
and U7484 (N_7484,N_6229,N_6316);
or U7485 (N_7485,N_6554,N_6969);
nor U7486 (N_7486,N_6763,N_6787);
nand U7487 (N_7487,N_6248,N_6484);
and U7488 (N_7488,N_6362,N_6225);
and U7489 (N_7489,N_6506,N_6274);
nor U7490 (N_7490,N_6373,N_6176);
or U7491 (N_7491,N_6749,N_6757);
nand U7492 (N_7492,N_6156,N_6572);
or U7493 (N_7493,N_6405,N_6295);
or U7494 (N_7494,N_6759,N_6463);
nor U7495 (N_7495,N_6481,N_6058);
and U7496 (N_7496,N_6577,N_6822);
xor U7497 (N_7497,N_6185,N_6071);
or U7498 (N_7498,N_6950,N_6465);
nand U7499 (N_7499,N_6502,N_6956);
xor U7500 (N_7500,N_6893,N_6845);
or U7501 (N_7501,N_6469,N_6299);
or U7502 (N_7502,N_6677,N_6121);
or U7503 (N_7503,N_6036,N_6678);
or U7504 (N_7504,N_6376,N_6609);
nor U7505 (N_7505,N_6913,N_6244);
or U7506 (N_7506,N_6060,N_6444);
nor U7507 (N_7507,N_6829,N_6442);
or U7508 (N_7508,N_6679,N_6345);
nor U7509 (N_7509,N_6625,N_6348);
xor U7510 (N_7510,N_6364,N_6266);
or U7511 (N_7511,N_6203,N_6058);
and U7512 (N_7512,N_6676,N_6059);
and U7513 (N_7513,N_6772,N_6630);
nand U7514 (N_7514,N_6610,N_6852);
and U7515 (N_7515,N_6922,N_6363);
and U7516 (N_7516,N_6503,N_6891);
nor U7517 (N_7517,N_6685,N_6773);
or U7518 (N_7518,N_6043,N_6894);
nand U7519 (N_7519,N_6810,N_6805);
xnor U7520 (N_7520,N_6012,N_6208);
and U7521 (N_7521,N_6964,N_6247);
xnor U7522 (N_7522,N_6405,N_6459);
nand U7523 (N_7523,N_6096,N_6609);
and U7524 (N_7524,N_6146,N_6048);
and U7525 (N_7525,N_6126,N_6807);
and U7526 (N_7526,N_6569,N_6988);
nor U7527 (N_7527,N_6387,N_6498);
or U7528 (N_7528,N_6802,N_6405);
nand U7529 (N_7529,N_6463,N_6080);
nor U7530 (N_7530,N_6665,N_6221);
nor U7531 (N_7531,N_6530,N_6174);
or U7532 (N_7532,N_6806,N_6891);
and U7533 (N_7533,N_6629,N_6914);
nor U7534 (N_7534,N_6251,N_6194);
or U7535 (N_7535,N_6239,N_6913);
xnor U7536 (N_7536,N_6325,N_6756);
or U7537 (N_7537,N_6367,N_6113);
xnor U7538 (N_7538,N_6428,N_6535);
nor U7539 (N_7539,N_6495,N_6501);
and U7540 (N_7540,N_6488,N_6453);
nand U7541 (N_7541,N_6726,N_6209);
xor U7542 (N_7542,N_6594,N_6666);
xor U7543 (N_7543,N_6071,N_6018);
nand U7544 (N_7544,N_6679,N_6944);
xor U7545 (N_7545,N_6593,N_6129);
xor U7546 (N_7546,N_6639,N_6326);
nand U7547 (N_7547,N_6656,N_6805);
and U7548 (N_7548,N_6021,N_6994);
and U7549 (N_7549,N_6548,N_6294);
nand U7550 (N_7550,N_6198,N_6995);
and U7551 (N_7551,N_6479,N_6687);
nand U7552 (N_7552,N_6233,N_6047);
and U7553 (N_7553,N_6568,N_6107);
xor U7554 (N_7554,N_6757,N_6694);
and U7555 (N_7555,N_6062,N_6868);
xor U7556 (N_7556,N_6744,N_6908);
xnor U7557 (N_7557,N_6878,N_6938);
nor U7558 (N_7558,N_6690,N_6820);
xor U7559 (N_7559,N_6478,N_6481);
or U7560 (N_7560,N_6084,N_6549);
nor U7561 (N_7561,N_6789,N_6013);
or U7562 (N_7562,N_6895,N_6222);
or U7563 (N_7563,N_6141,N_6776);
xnor U7564 (N_7564,N_6971,N_6669);
and U7565 (N_7565,N_6350,N_6336);
and U7566 (N_7566,N_6184,N_6007);
and U7567 (N_7567,N_6983,N_6141);
nor U7568 (N_7568,N_6707,N_6862);
xor U7569 (N_7569,N_6017,N_6996);
or U7570 (N_7570,N_6895,N_6338);
nor U7571 (N_7571,N_6354,N_6561);
or U7572 (N_7572,N_6735,N_6575);
nor U7573 (N_7573,N_6255,N_6166);
nand U7574 (N_7574,N_6751,N_6132);
or U7575 (N_7575,N_6172,N_6952);
nor U7576 (N_7576,N_6962,N_6154);
nand U7577 (N_7577,N_6875,N_6254);
nand U7578 (N_7578,N_6229,N_6641);
nand U7579 (N_7579,N_6725,N_6111);
nand U7580 (N_7580,N_6722,N_6831);
nor U7581 (N_7581,N_6675,N_6977);
nor U7582 (N_7582,N_6111,N_6288);
nor U7583 (N_7583,N_6037,N_6793);
nand U7584 (N_7584,N_6390,N_6907);
nand U7585 (N_7585,N_6974,N_6445);
xor U7586 (N_7586,N_6572,N_6247);
and U7587 (N_7587,N_6210,N_6167);
nor U7588 (N_7588,N_6368,N_6671);
and U7589 (N_7589,N_6776,N_6092);
or U7590 (N_7590,N_6905,N_6227);
nand U7591 (N_7591,N_6293,N_6801);
and U7592 (N_7592,N_6965,N_6773);
and U7593 (N_7593,N_6674,N_6440);
or U7594 (N_7594,N_6106,N_6357);
or U7595 (N_7595,N_6761,N_6747);
xor U7596 (N_7596,N_6481,N_6377);
nor U7597 (N_7597,N_6044,N_6758);
nand U7598 (N_7598,N_6026,N_6016);
or U7599 (N_7599,N_6961,N_6820);
nand U7600 (N_7600,N_6565,N_6920);
and U7601 (N_7601,N_6606,N_6166);
and U7602 (N_7602,N_6160,N_6694);
xor U7603 (N_7603,N_6136,N_6097);
nor U7604 (N_7604,N_6942,N_6825);
xnor U7605 (N_7605,N_6231,N_6880);
nor U7606 (N_7606,N_6737,N_6774);
xor U7607 (N_7607,N_6722,N_6644);
or U7608 (N_7608,N_6044,N_6276);
nand U7609 (N_7609,N_6754,N_6928);
or U7610 (N_7610,N_6680,N_6564);
nor U7611 (N_7611,N_6183,N_6645);
nand U7612 (N_7612,N_6172,N_6665);
or U7613 (N_7613,N_6553,N_6771);
nand U7614 (N_7614,N_6181,N_6333);
nand U7615 (N_7615,N_6584,N_6295);
and U7616 (N_7616,N_6290,N_6602);
xor U7617 (N_7617,N_6751,N_6463);
and U7618 (N_7618,N_6016,N_6967);
nand U7619 (N_7619,N_6957,N_6525);
or U7620 (N_7620,N_6124,N_6929);
nand U7621 (N_7621,N_6595,N_6610);
nand U7622 (N_7622,N_6080,N_6732);
nand U7623 (N_7623,N_6062,N_6741);
nor U7624 (N_7624,N_6292,N_6594);
and U7625 (N_7625,N_6743,N_6759);
or U7626 (N_7626,N_6562,N_6525);
nand U7627 (N_7627,N_6820,N_6250);
and U7628 (N_7628,N_6628,N_6186);
nor U7629 (N_7629,N_6237,N_6537);
nand U7630 (N_7630,N_6714,N_6381);
and U7631 (N_7631,N_6577,N_6954);
xnor U7632 (N_7632,N_6887,N_6547);
nand U7633 (N_7633,N_6109,N_6531);
xnor U7634 (N_7634,N_6396,N_6940);
xnor U7635 (N_7635,N_6638,N_6620);
and U7636 (N_7636,N_6273,N_6095);
and U7637 (N_7637,N_6755,N_6527);
or U7638 (N_7638,N_6348,N_6035);
and U7639 (N_7639,N_6709,N_6444);
nand U7640 (N_7640,N_6146,N_6376);
or U7641 (N_7641,N_6781,N_6548);
or U7642 (N_7642,N_6688,N_6606);
nor U7643 (N_7643,N_6692,N_6847);
or U7644 (N_7644,N_6059,N_6529);
or U7645 (N_7645,N_6016,N_6730);
or U7646 (N_7646,N_6031,N_6417);
nor U7647 (N_7647,N_6936,N_6239);
nor U7648 (N_7648,N_6999,N_6321);
xor U7649 (N_7649,N_6585,N_6832);
or U7650 (N_7650,N_6920,N_6296);
nor U7651 (N_7651,N_6629,N_6783);
nand U7652 (N_7652,N_6327,N_6064);
or U7653 (N_7653,N_6812,N_6091);
or U7654 (N_7654,N_6107,N_6447);
xnor U7655 (N_7655,N_6368,N_6384);
xor U7656 (N_7656,N_6168,N_6591);
nor U7657 (N_7657,N_6152,N_6144);
and U7658 (N_7658,N_6701,N_6345);
and U7659 (N_7659,N_6232,N_6959);
nor U7660 (N_7660,N_6622,N_6494);
nor U7661 (N_7661,N_6388,N_6100);
and U7662 (N_7662,N_6188,N_6668);
nand U7663 (N_7663,N_6687,N_6533);
nor U7664 (N_7664,N_6341,N_6264);
nor U7665 (N_7665,N_6942,N_6566);
or U7666 (N_7666,N_6466,N_6029);
nand U7667 (N_7667,N_6785,N_6047);
and U7668 (N_7668,N_6266,N_6304);
nand U7669 (N_7669,N_6695,N_6912);
nand U7670 (N_7670,N_6336,N_6274);
nor U7671 (N_7671,N_6045,N_6782);
or U7672 (N_7672,N_6196,N_6335);
and U7673 (N_7673,N_6978,N_6578);
xor U7674 (N_7674,N_6581,N_6433);
nor U7675 (N_7675,N_6917,N_6421);
nor U7676 (N_7676,N_6005,N_6461);
xnor U7677 (N_7677,N_6159,N_6316);
nor U7678 (N_7678,N_6650,N_6192);
xnor U7679 (N_7679,N_6230,N_6331);
and U7680 (N_7680,N_6577,N_6651);
xor U7681 (N_7681,N_6884,N_6057);
and U7682 (N_7682,N_6670,N_6495);
xnor U7683 (N_7683,N_6673,N_6808);
or U7684 (N_7684,N_6617,N_6778);
nor U7685 (N_7685,N_6378,N_6078);
or U7686 (N_7686,N_6256,N_6723);
xnor U7687 (N_7687,N_6779,N_6369);
xnor U7688 (N_7688,N_6190,N_6833);
and U7689 (N_7689,N_6613,N_6121);
xnor U7690 (N_7690,N_6032,N_6204);
or U7691 (N_7691,N_6685,N_6279);
xor U7692 (N_7692,N_6861,N_6520);
xnor U7693 (N_7693,N_6404,N_6327);
nand U7694 (N_7694,N_6116,N_6922);
nand U7695 (N_7695,N_6269,N_6369);
nand U7696 (N_7696,N_6755,N_6237);
nand U7697 (N_7697,N_6671,N_6011);
or U7698 (N_7698,N_6825,N_6072);
nand U7699 (N_7699,N_6288,N_6459);
nand U7700 (N_7700,N_6864,N_6989);
nand U7701 (N_7701,N_6103,N_6447);
and U7702 (N_7702,N_6761,N_6632);
xnor U7703 (N_7703,N_6955,N_6133);
and U7704 (N_7704,N_6543,N_6690);
or U7705 (N_7705,N_6525,N_6396);
or U7706 (N_7706,N_6666,N_6904);
or U7707 (N_7707,N_6978,N_6117);
and U7708 (N_7708,N_6935,N_6882);
xnor U7709 (N_7709,N_6210,N_6956);
xor U7710 (N_7710,N_6429,N_6675);
and U7711 (N_7711,N_6361,N_6193);
xor U7712 (N_7712,N_6560,N_6795);
xor U7713 (N_7713,N_6472,N_6147);
xnor U7714 (N_7714,N_6450,N_6493);
xor U7715 (N_7715,N_6961,N_6169);
and U7716 (N_7716,N_6890,N_6601);
nor U7717 (N_7717,N_6139,N_6013);
or U7718 (N_7718,N_6053,N_6154);
xor U7719 (N_7719,N_6793,N_6806);
xnor U7720 (N_7720,N_6638,N_6425);
nor U7721 (N_7721,N_6238,N_6085);
nand U7722 (N_7722,N_6306,N_6938);
or U7723 (N_7723,N_6138,N_6297);
or U7724 (N_7724,N_6463,N_6847);
nor U7725 (N_7725,N_6455,N_6814);
and U7726 (N_7726,N_6627,N_6850);
xnor U7727 (N_7727,N_6386,N_6363);
and U7728 (N_7728,N_6596,N_6436);
or U7729 (N_7729,N_6319,N_6740);
and U7730 (N_7730,N_6708,N_6578);
nor U7731 (N_7731,N_6392,N_6027);
nor U7732 (N_7732,N_6366,N_6604);
nand U7733 (N_7733,N_6742,N_6057);
xor U7734 (N_7734,N_6792,N_6534);
nand U7735 (N_7735,N_6744,N_6069);
or U7736 (N_7736,N_6623,N_6769);
nor U7737 (N_7737,N_6519,N_6089);
and U7738 (N_7738,N_6314,N_6649);
or U7739 (N_7739,N_6803,N_6704);
nor U7740 (N_7740,N_6671,N_6263);
xnor U7741 (N_7741,N_6324,N_6228);
or U7742 (N_7742,N_6474,N_6643);
and U7743 (N_7743,N_6704,N_6141);
or U7744 (N_7744,N_6958,N_6047);
nand U7745 (N_7745,N_6211,N_6607);
nand U7746 (N_7746,N_6665,N_6901);
nand U7747 (N_7747,N_6931,N_6824);
nand U7748 (N_7748,N_6482,N_6011);
nand U7749 (N_7749,N_6259,N_6709);
or U7750 (N_7750,N_6243,N_6885);
nand U7751 (N_7751,N_6316,N_6742);
nand U7752 (N_7752,N_6864,N_6816);
nand U7753 (N_7753,N_6485,N_6247);
and U7754 (N_7754,N_6341,N_6747);
nand U7755 (N_7755,N_6586,N_6626);
and U7756 (N_7756,N_6414,N_6740);
nor U7757 (N_7757,N_6975,N_6133);
or U7758 (N_7758,N_6399,N_6984);
or U7759 (N_7759,N_6260,N_6157);
and U7760 (N_7760,N_6213,N_6093);
and U7761 (N_7761,N_6974,N_6800);
or U7762 (N_7762,N_6027,N_6006);
and U7763 (N_7763,N_6699,N_6641);
xnor U7764 (N_7764,N_6690,N_6756);
nor U7765 (N_7765,N_6727,N_6526);
or U7766 (N_7766,N_6514,N_6248);
xnor U7767 (N_7767,N_6220,N_6805);
and U7768 (N_7768,N_6691,N_6993);
and U7769 (N_7769,N_6691,N_6802);
and U7770 (N_7770,N_6758,N_6591);
nand U7771 (N_7771,N_6861,N_6283);
xor U7772 (N_7772,N_6720,N_6465);
nand U7773 (N_7773,N_6133,N_6240);
or U7774 (N_7774,N_6613,N_6476);
or U7775 (N_7775,N_6448,N_6493);
xnor U7776 (N_7776,N_6587,N_6322);
nor U7777 (N_7777,N_6799,N_6190);
nor U7778 (N_7778,N_6319,N_6613);
nand U7779 (N_7779,N_6030,N_6809);
nor U7780 (N_7780,N_6893,N_6967);
nand U7781 (N_7781,N_6945,N_6915);
or U7782 (N_7782,N_6143,N_6129);
and U7783 (N_7783,N_6051,N_6009);
and U7784 (N_7784,N_6806,N_6183);
and U7785 (N_7785,N_6798,N_6288);
and U7786 (N_7786,N_6926,N_6024);
nand U7787 (N_7787,N_6781,N_6018);
and U7788 (N_7788,N_6344,N_6917);
nand U7789 (N_7789,N_6007,N_6946);
nand U7790 (N_7790,N_6562,N_6722);
xor U7791 (N_7791,N_6420,N_6840);
xnor U7792 (N_7792,N_6636,N_6816);
or U7793 (N_7793,N_6707,N_6879);
or U7794 (N_7794,N_6994,N_6810);
nor U7795 (N_7795,N_6008,N_6068);
and U7796 (N_7796,N_6928,N_6445);
and U7797 (N_7797,N_6292,N_6467);
xor U7798 (N_7798,N_6545,N_6126);
xor U7799 (N_7799,N_6815,N_6931);
nor U7800 (N_7800,N_6758,N_6493);
or U7801 (N_7801,N_6459,N_6303);
and U7802 (N_7802,N_6940,N_6761);
xor U7803 (N_7803,N_6426,N_6624);
xor U7804 (N_7804,N_6583,N_6540);
and U7805 (N_7805,N_6394,N_6100);
and U7806 (N_7806,N_6875,N_6052);
xnor U7807 (N_7807,N_6771,N_6784);
xor U7808 (N_7808,N_6829,N_6189);
nor U7809 (N_7809,N_6558,N_6468);
and U7810 (N_7810,N_6051,N_6413);
nand U7811 (N_7811,N_6073,N_6167);
and U7812 (N_7812,N_6367,N_6411);
nor U7813 (N_7813,N_6366,N_6800);
or U7814 (N_7814,N_6638,N_6171);
nand U7815 (N_7815,N_6241,N_6603);
nor U7816 (N_7816,N_6020,N_6426);
nand U7817 (N_7817,N_6136,N_6178);
or U7818 (N_7818,N_6929,N_6056);
xnor U7819 (N_7819,N_6855,N_6007);
nor U7820 (N_7820,N_6999,N_6876);
nand U7821 (N_7821,N_6326,N_6319);
nor U7822 (N_7822,N_6983,N_6389);
xor U7823 (N_7823,N_6331,N_6113);
or U7824 (N_7824,N_6876,N_6029);
xnor U7825 (N_7825,N_6751,N_6160);
nor U7826 (N_7826,N_6578,N_6172);
nor U7827 (N_7827,N_6304,N_6143);
xnor U7828 (N_7828,N_6289,N_6640);
xor U7829 (N_7829,N_6097,N_6171);
and U7830 (N_7830,N_6375,N_6095);
or U7831 (N_7831,N_6503,N_6003);
and U7832 (N_7832,N_6352,N_6944);
or U7833 (N_7833,N_6493,N_6407);
nand U7834 (N_7834,N_6658,N_6803);
xnor U7835 (N_7835,N_6193,N_6598);
nor U7836 (N_7836,N_6310,N_6374);
or U7837 (N_7837,N_6939,N_6173);
or U7838 (N_7838,N_6171,N_6841);
nand U7839 (N_7839,N_6641,N_6603);
and U7840 (N_7840,N_6232,N_6257);
xnor U7841 (N_7841,N_6505,N_6801);
and U7842 (N_7842,N_6230,N_6903);
nor U7843 (N_7843,N_6198,N_6051);
nand U7844 (N_7844,N_6222,N_6752);
or U7845 (N_7845,N_6622,N_6935);
xnor U7846 (N_7846,N_6609,N_6592);
nor U7847 (N_7847,N_6196,N_6517);
xnor U7848 (N_7848,N_6895,N_6761);
or U7849 (N_7849,N_6931,N_6466);
and U7850 (N_7850,N_6430,N_6802);
nor U7851 (N_7851,N_6217,N_6518);
nand U7852 (N_7852,N_6812,N_6131);
nand U7853 (N_7853,N_6963,N_6177);
and U7854 (N_7854,N_6922,N_6982);
nor U7855 (N_7855,N_6445,N_6322);
nor U7856 (N_7856,N_6064,N_6768);
xor U7857 (N_7857,N_6413,N_6560);
and U7858 (N_7858,N_6005,N_6682);
and U7859 (N_7859,N_6698,N_6823);
nor U7860 (N_7860,N_6238,N_6355);
xnor U7861 (N_7861,N_6680,N_6446);
nor U7862 (N_7862,N_6914,N_6084);
nor U7863 (N_7863,N_6434,N_6687);
nor U7864 (N_7864,N_6554,N_6392);
and U7865 (N_7865,N_6453,N_6715);
xnor U7866 (N_7866,N_6937,N_6250);
nand U7867 (N_7867,N_6897,N_6272);
and U7868 (N_7868,N_6837,N_6982);
or U7869 (N_7869,N_6841,N_6677);
and U7870 (N_7870,N_6944,N_6613);
or U7871 (N_7871,N_6842,N_6948);
and U7872 (N_7872,N_6511,N_6193);
nand U7873 (N_7873,N_6595,N_6913);
xnor U7874 (N_7874,N_6728,N_6656);
nand U7875 (N_7875,N_6500,N_6935);
or U7876 (N_7876,N_6018,N_6058);
xor U7877 (N_7877,N_6634,N_6554);
or U7878 (N_7878,N_6660,N_6567);
nand U7879 (N_7879,N_6192,N_6904);
or U7880 (N_7880,N_6166,N_6304);
nor U7881 (N_7881,N_6096,N_6475);
nor U7882 (N_7882,N_6037,N_6792);
nand U7883 (N_7883,N_6512,N_6645);
and U7884 (N_7884,N_6677,N_6151);
and U7885 (N_7885,N_6376,N_6356);
nor U7886 (N_7886,N_6630,N_6411);
or U7887 (N_7887,N_6632,N_6407);
or U7888 (N_7888,N_6072,N_6165);
and U7889 (N_7889,N_6478,N_6808);
xor U7890 (N_7890,N_6953,N_6270);
nor U7891 (N_7891,N_6885,N_6170);
and U7892 (N_7892,N_6658,N_6497);
nand U7893 (N_7893,N_6384,N_6081);
nor U7894 (N_7894,N_6945,N_6597);
xnor U7895 (N_7895,N_6962,N_6060);
xor U7896 (N_7896,N_6993,N_6077);
xnor U7897 (N_7897,N_6925,N_6386);
nand U7898 (N_7898,N_6056,N_6314);
xor U7899 (N_7899,N_6828,N_6083);
and U7900 (N_7900,N_6919,N_6806);
or U7901 (N_7901,N_6806,N_6949);
or U7902 (N_7902,N_6291,N_6626);
and U7903 (N_7903,N_6675,N_6763);
nand U7904 (N_7904,N_6184,N_6680);
nand U7905 (N_7905,N_6282,N_6104);
nand U7906 (N_7906,N_6199,N_6789);
nor U7907 (N_7907,N_6033,N_6726);
nor U7908 (N_7908,N_6513,N_6888);
xor U7909 (N_7909,N_6432,N_6040);
nand U7910 (N_7910,N_6727,N_6543);
nor U7911 (N_7911,N_6751,N_6538);
nand U7912 (N_7912,N_6431,N_6738);
or U7913 (N_7913,N_6874,N_6485);
and U7914 (N_7914,N_6380,N_6659);
nand U7915 (N_7915,N_6165,N_6676);
xnor U7916 (N_7916,N_6691,N_6129);
xor U7917 (N_7917,N_6874,N_6755);
or U7918 (N_7918,N_6055,N_6013);
or U7919 (N_7919,N_6109,N_6865);
and U7920 (N_7920,N_6181,N_6394);
and U7921 (N_7921,N_6444,N_6875);
nor U7922 (N_7922,N_6835,N_6539);
nand U7923 (N_7923,N_6935,N_6482);
nor U7924 (N_7924,N_6530,N_6887);
nand U7925 (N_7925,N_6450,N_6550);
nand U7926 (N_7926,N_6310,N_6502);
or U7927 (N_7927,N_6477,N_6577);
nor U7928 (N_7928,N_6566,N_6085);
nand U7929 (N_7929,N_6453,N_6307);
nor U7930 (N_7930,N_6591,N_6183);
and U7931 (N_7931,N_6323,N_6004);
nor U7932 (N_7932,N_6295,N_6213);
nor U7933 (N_7933,N_6748,N_6071);
nor U7934 (N_7934,N_6709,N_6249);
and U7935 (N_7935,N_6932,N_6232);
and U7936 (N_7936,N_6485,N_6725);
xor U7937 (N_7937,N_6718,N_6492);
nor U7938 (N_7938,N_6328,N_6090);
nand U7939 (N_7939,N_6852,N_6668);
and U7940 (N_7940,N_6265,N_6298);
nand U7941 (N_7941,N_6655,N_6612);
nand U7942 (N_7942,N_6786,N_6777);
or U7943 (N_7943,N_6202,N_6723);
nand U7944 (N_7944,N_6419,N_6372);
nor U7945 (N_7945,N_6879,N_6523);
xnor U7946 (N_7946,N_6000,N_6429);
and U7947 (N_7947,N_6117,N_6776);
nor U7948 (N_7948,N_6315,N_6818);
nand U7949 (N_7949,N_6498,N_6241);
nand U7950 (N_7950,N_6971,N_6850);
and U7951 (N_7951,N_6594,N_6511);
nand U7952 (N_7952,N_6701,N_6768);
and U7953 (N_7953,N_6348,N_6487);
nor U7954 (N_7954,N_6427,N_6773);
xnor U7955 (N_7955,N_6630,N_6848);
or U7956 (N_7956,N_6420,N_6457);
and U7957 (N_7957,N_6235,N_6620);
nand U7958 (N_7958,N_6511,N_6814);
xor U7959 (N_7959,N_6558,N_6074);
nor U7960 (N_7960,N_6126,N_6953);
nor U7961 (N_7961,N_6124,N_6851);
or U7962 (N_7962,N_6297,N_6073);
and U7963 (N_7963,N_6302,N_6631);
or U7964 (N_7964,N_6686,N_6809);
and U7965 (N_7965,N_6840,N_6256);
xnor U7966 (N_7966,N_6985,N_6035);
nand U7967 (N_7967,N_6088,N_6113);
or U7968 (N_7968,N_6864,N_6596);
and U7969 (N_7969,N_6044,N_6357);
and U7970 (N_7970,N_6220,N_6137);
and U7971 (N_7971,N_6385,N_6975);
nand U7972 (N_7972,N_6845,N_6336);
nand U7973 (N_7973,N_6333,N_6324);
xor U7974 (N_7974,N_6988,N_6623);
or U7975 (N_7975,N_6709,N_6274);
nor U7976 (N_7976,N_6627,N_6225);
and U7977 (N_7977,N_6763,N_6491);
xor U7978 (N_7978,N_6383,N_6370);
nor U7979 (N_7979,N_6952,N_6106);
and U7980 (N_7980,N_6179,N_6099);
or U7981 (N_7981,N_6154,N_6514);
xor U7982 (N_7982,N_6722,N_6506);
nor U7983 (N_7983,N_6425,N_6215);
or U7984 (N_7984,N_6856,N_6752);
and U7985 (N_7985,N_6782,N_6159);
xor U7986 (N_7986,N_6450,N_6688);
or U7987 (N_7987,N_6087,N_6080);
nor U7988 (N_7988,N_6701,N_6929);
nor U7989 (N_7989,N_6525,N_6193);
or U7990 (N_7990,N_6485,N_6124);
nand U7991 (N_7991,N_6914,N_6123);
and U7992 (N_7992,N_6855,N_6225);
and U7993 (N_7993,N_6800,N_6538);
and U7994 (N_7994,N_6890,N_6370);
nand U7995 (N_7995,N_6987,N_6916);
and U7996 (N_7996,N_6863,N_6342);
or U7997 (N_7997,N_6226,N_6227);
nand U7998 (N_7998,N_6742,N_6605);
nor U7999 (N_7999,N_6250,N_6398);
nand U8000 (N_8000,N_7229,N_7200);
nor U8001 (N_8001,N_7040,N_7533);
nand U8002 (N_8002,N_7561,N_7409);
nor U8003 (N_8003,N_7800,N_7625);
and U8004 (N_8004,N_7001,N_7174);
nor U8005 (N_8005,N_7156,N_7193);
or U8006 (N_8006,N_7120,N_7171);
xor U8007 (N_8007,N_7194,N_7988);
xnor U8008 (N_8008,N_7771,N_7497);
xor U8009 (N_8009,N_7922,N_7687);
nand U8010 (N_8010,N_7935,N_7643);
xnor U8011 (N_8011,N_7803,N_7150);
xor U8012 (N_8012,N_7668,N_7341);
nand U8013 (N_8013,N_7996,N_7874);
and U8014 (N_8014,N_7384,N_7285);
nand U8015 (N_8015,N_7715,N_7936);
nor U8016 (N_8016,N_7818,N_7843);
nand U8017 (N_8017,N_7430,N_7461);
and U8018 (N_8018,N_7439,N_7710);
xnor U8019 (N_8019,N_7196,N_7581);
xor U8020 (N_8020,N_7294,N_7006);
nand U8021 (N_8021,N_7496,N_7751);
nand U8022 (N_8022,N_7722,N_7947);
or U8023 (N_8023,N_7232,N_7280);
and U8024 (N_8024,N_7367,N_7888);
nor U8025 (N_8025,N_7370,N_7420);
and U8026 (N_8026,N_7518,N_7587);
and U8027 (N_8027,N_7291,N_7689);
nor U8028 (N_8028,N_7122,N_7125);
xnor U8029 (N_8029,N_7806,N_7247);
xor U8030 (N_8030,N_7354,N_7113);
or U8031 (N_8031,N_7161,N_7974);
nor U8032 (N_8032,N_7101,N_7071);
xor U8033 (N_8033,N_7024,N_7824);
nor U8034 (N_8034,N_7221,N_7891);
xnor U8035 (N_8035,N_7777,N_7732);
or U8036 (N_8036,N_7433,N_7741);
and U8037 (N_8037,N_7617,N_7240);
xnor U8038 (N_8038,N_7465,N_7223);
xnor U8039 (N_8039,N_7666,N_7269);
and U8040 (N_8040,N_7032,N_7211);
nand U8041 (N_8041,N_7277,N_7117);
and U8042 (N_8042,N_7986,N_7190);
or U8043 (N_8043,N_7956,N_7139);
nor U8044 (N_8044,N_7627,N_7437);
xnor U8045 (N_8045,N_7393,N_7186);
xnor U8046 (N_8046,N_7652,N_7697);
xor U8047 (N_8047,N_7312,N_7353);
nand U8048 (N_8048,N_7245,N_7960);
or U8049 (N_8049,N_7743,N_7281);
nor U8050 (N_8050,N_7736,N_7320);
nand U8051 (N_8051,N_7205,N_7304);
or U8052 (N_8052,N_7417,N_7016);
xnor U8053 (N_8053,N_7178,N_7271);
or U8054 (N_8054,N_7014,N_7940);
and U8055 (N_8055,N_7141,N_7176);
xnor U8056 (N_8056,N_7490,N_7570);
xor U8057 (N_8057,N_7169,N_7943);
or U8058 (N_8058,N_7031,N_7829);
nor U8059 (N_8059,N_7575,N_7415);
xor U8060 (N_8060,N_7334,N_7624);
and U8061 (N_8061,N_7067,N_7614);
xnor U8062 (N_8062,N_7330,N_7840);
nor U8063 (N_8063,N_7758,N_7698);
and U8064 (N_8064,N_7403,N_7089);
nand U8065 (N_8065,N_7337,N_7425);
nand U8066 (N_8066,N_7955,N_7767);
xnor U8067 (N_8067,N_7102,N_7589);
nand U8068 (N_8068,N_7553,N_7939);
or U8069 (N_8069,N_7750,N_7999);
nor U8070 (N_8070,N_7463,N_7686);
and U8071 (N_8071,N_7755,N_7554);
or U8072 (N_8072,N_7607,N_7085);
nand U8073 (N_8073,N_7180,N_7308);
xnor U8074 (N_8074,N_7765,N_7375);
nor U8075 (N_8075,N_7932,N_7363);
nand U8076 (N_8076,N_7987,N_7912);
xor U8077 (N_8077,N_7984,N_7060);
nand U8078 (N_8078,N_7386,N_7339);
nand U8079 (N_8079,N_7526,N_7438);
and U8080 (N_8080,N_7941,N_7458);
and U8081 (N_8081,N_7965,N_7075);
or U8082 (N_8082,N_7459,N_7620);
or U8083 (N_8083,N_7610,N_7557);
nand U8084 (N_8084,N_7709,N_7616);
nor U8085 (N_8085,N_7307,N_7660);
and U8086 (N_8086,N_7931,N_7466);
nor U8087 (N_8087,N_7842,N_7702);
and U8088 (N_8088,N_7725,N_7734);
and U8089 (N_8089,N_7651,N_7305);
or U8090 (N_8090,N_7175,N_7757);
and U8091 (N_8091,N_7055,N_7306);
nor U8092 (N_8092,N_7664,N_7347);
nand U8093 (N_8093,N_7392,N_7880);
xor U8094 (N_8094,N_7914,N_7090);
and U8095 (N_8095,N_7469,N_7527);
nand U8096 (N_8096,N_7213,N_7528);
and U8097 (N_8097,N_7153,N_7388);
or U8098 (N_8098,N_7235,N_7504);
xor U8099 (N_8099,N_7394,N_7064);
and U8100 (N_8100,N_7683,N_7905);
xor U8101 (N_8101,N_7103,N_7236);
xnor U8102 (N_8102,N_7747,N_7712);
and U8103 (N_8103,N_7076,N_7719);
nor U8104 (N_8104,N_7779,N_7704);
nor U8105 (N_8105,N_7980,N_7331);
or U8106 (N_8106,N_7019,N_7047);
nand U8107 (N_8107,N_7756,N_7817);
nand U8108 (N_8108,N_7079,N_7612);
nand U8109 (N_8109,N_7982,N_7883);
and U8110 (N_8110,N_7916,N_7688);
nor U8111 (N_8111,N_7952,N_7789);
or U8112 (N_8112,N_7154,N_7549);
and U8113 (N_8113,N_7477,N_7680);
xnor U8114 (N_8114,N_7866,N_7074);
nand U8115 (N_8115,N_7084,N_7314);
or U8116 (N_8116,N_7547,N_7781);
nor U8117 (N_8117,N_7256,N_7368);
xnor U8118 (N_8118,N_7140,N_7515);
nand U8119 (N_8119,N_7480,N_7954);
xor U8120 (N_8120,N_7691,N_7366);
xor U8121 (N_8121,N_7372,N_7858);
and U8122 (N_8122,N_7721,N_7069);
xnor U8123 (N_8123,N_7682,N_7993);
nand U8124 (N_8124,N_7637,N_7115);
or U8125 (N_8125,N_7656,N_7548);
or U8126 (N_8126,N_7377,N_7413);
or U8127 (N_8127,N_7934,N_7804);
or U8128 (N_8128,N_7718,N_7740);
nand U8129 (N_8129,N_7423,N_7816);
nor U8130 (N_8130,N_7865,N_7565);
and U8131 (N_8131,N_7749,N_7135);
nor U8132 (N_8132,N_7969,N_7784);
or U8133 (N_8133,N_7317,N_7052);
xnor U8134 (N_8134,N_7093,N_7897);
nor U8135 (N_8135,N_7289,N_7631);
nor U8136 (N_8136,N_7975,N_7847);
xor U8137 (N_8137,N_7147,N_7405);
xnor U8138 (N_8138,N_7107,N_7144);
xnor U8139 (N_8139,N_7228,N_7299);
xnor U8140 (N_8140,N_7365,N_7266);
nor U8141 (N_8141,N_7551,N_7673);
nand U8142 (N_8142,N_7907,N_7542);
nor U8143 (N_8143,N_7489,N_7802);
nor U8144 (N_8144,N_7048,N_7857);
and U8145 (N_8145,N_7615,N_7795);
xnor U8146 (N_8146,N_7769,N_7119);
or U8147 (N_8147,N_7894,N_7162);
xor U8148 (N_8148,N_7184,N_7116);
nor U8149 (N_8149,N_7373,N_7644);
and U8150 (N_8150,N_7953,N_7951);
or U8151 (N_8151,N_7825,N_7412);
nor U8152 (N_8152,N_7977,N_7029);
and U8153 (N_8153,N_7177,N_7971);
nand U8154 (N_8154,N_7705,N_7851);
xnor U8155 (N_8155,N_7056,N_7507);
nand U8156 (N_8156,N_7471,N_7219);
or U8157 (N_8157,N_7649,N_7378);
nor U8158 (N_8158,N_7495,N_7853);
and U8159 (N_8159,N_7889,N_7967);
xor U8160 (N_8160,N_7227,N_7435);
nand U8161 (N_8161,N_7634,N_7583);
nand U8162 (N_8162,N_7083,N_7051);
xor U8163 (N_8163,N_7854,N_7142);
and U8164 (N_8164,N_7564,N_7796);
or U8165 (N_8165,N_7904,N_7097);
and U8166 (N_8166,N_7112,N_7622);
or U8167 (N_8167,N_7035,N_7774);
and U8168 (N_8168,N_7920,N_7838);
and U8169 (N_8169,N_7215,N_7185);
xnor U8170 (N_8170,N_7160,N_7836);
or U8171 (N_8171,N_7309,N_7168);
nand U8172 (N_8172,N_7961,N_7399);
nand U8173 (N_8173,N_7500,N_7327);
and U8174 (N_8174,N_7862,N_7559);
nand U8175 (N_8175,N_7319,N_7890);
or U8176 (N_8176,N_7414,N_7994);
nand U8177 (N_8177,N_7131,N_7033);
nand U8178 (N_8178,N_7877,N_7525);
xor U8179 (N_8179,N_7493,N_7761);
or U8180 (N_8180,N_7199,N_7628);
nor U8181 (N_8181,N_7273,N_7510);
and U8182 (N_8182,N_7911,N_7856);
nor U8183 (N_8183,N_7270,N_7716);
or U8184 (N_8184,N_7648,N_7592);
and U8185 (N_8185,N_7577,N_7647);
or U8186 (N_8186,N_7867,N_7241);
xor U8187 (N_8187,N_7663,N_7326);
xnor U8188 (N_8188,N_7580,N_7272);
and U8189 (N_8189,N_7595,N_7487);
or U8190 (N_8190,N_7872,N_7303);
xnor U8191 (N_8191,N_7808,N_7604);
nand U8192 (N_8192,N_7619,N_7517);
or U8193 (N_8193,N_7183,N_7336);
nor U8194 (N_8194,N_7724,N_7224);
nand U8195 (N_8195,N_7809,N_7700);
nor U8196 (N_8196,N_7202,N_7066);
nand U8197 (N_8197,N_7105,N_7950);
xnor U8198 (N_8198,N_7792,N_7424);
xor U8199 (N_8199,N_7195,N_7881);
nor U8200 (N_8200,N_7087,N_7670);
nand U8201 (N_8201,N_7855,N_7030);
and U8202 (N_8202,N_7594,N_7284);
nor U8203 (N_8203,N_7099,N_7310);
and U8204 (N_8204,N_7733,N_7599);
xnor U8205 (N_8205,N_7096,N_7863);
or U8206 (N_8206,N_7930,N_7159);
or U8207 (N_8207,N_7222,N_7778);
and U8208 (N_8208,N_7609,N_7626);
nor U8209 (N_8209,N_7332,N_7204);
xnor U8210 (N_8210,N_7025,N_7927);
or U8211 (N_8211,N_7263,N_7296);
nor U8212 (N_8212,N_7022,N_7027);
nand U8213 (N_8213,N_7203,N_7764);
nor U8214 (N_8214,N_7360,N_7453);
and U8215 (N_8215,N_7072,N_7639);
nor U8216 (N_8216,N_7972,N_7402);
nand U8217 (N_8217,N_7845,N_7913);
or U8218 (N_8218,N_7640,N_7411);
or U8219 (N_8219,N_7748,N_7841);
xnor U8220 (N_8220,N_7288,N_7871);
nand U8221 (N_8221,N_7359,N_7316);
nand U8222 (N_8222,N_7541,N_7369);
nor U8223 (N_8223,N_7449,N_7110);
or U8224 (N_8224,N_7828,N_7835);
nand U8225 (N_8225,N_7552,N_7167);
nand U8226 (N_8226,N_7821,N_7023);
nand U8227 (N_8227,N_7436,N_7418);
or U8228 (N_8228,N_7046,N_7109);
nand U8229 (N_8229,N_7432,N_7638);
nor U8230 (N_8230,N_7082,N_7968);
nand U8231 (N_8231,N_7250,N_7333);
xnor U8232 (N_8232,N_7448,N_7145);
nor U8233 (N_8233,N_7793,N_7545);
xnor U8234 (N_8234,N_7070,N_7293);
nor U8235 (N_8235,N_7282,N_7873);
nor U8236 (N_8236,N_7677,N_7900);
xnor U8237 (N_8237,N_7957,N_7343);
nor U8238 (N_8238,N_7860,N_7283);
and U8239 (N_8239,N_7861,N_7641);
xnor U8240 (N_8240,N_7569,N_7003);
or U8241 (N_8241,N_7529,N_7586);
nand U8242 (N_8242,N_7603,N_7189);
or U8243 (N_8243,N_7279,N_7513);
and U8244 (N_8244,N_7259,N_7717);
xor U8245 (N_8245,N_7864,N_7128);
or U8246 (N_8246,N_7775,N_7606);
nand U8247 (N_8247,N_7410,N_7192);
nand U8248 (N_8248,N_7906,N_7801);
and U8249 (N_8249,N_7532,N_7884);
xor U8250 (N_8250,N_7540,N_7650);
and U8251 (N_8251,N_7268,N_7179);
and U8252 (N_8252,N_7699,N_7512);
xnor U8253 (N_8253,N_7970,N_7483);
or U8254 (N_8254,N_7695,N_7026);
nand U8255 (N_8255,N_7276,N_7735);
or U8256 (N_8256,N_7077,N_7558);
or U8257 (N_8257,N_7440,N_7646);
xor U8258 (N_8258,N_7002,N_7297);
and U8259 (N_8259,N_7218,N_7138);
nor U8260 (N_8260,N_7582,N_7400);
nand U8261 (N_8261,N_7636,N_7539);
xor U8262 (N_8262,N_7530,N_7703);
nor U8263 (N_8263,N_7166,N_7706);
nand U8264 (N_8264,N_7349,N_7254);
and U8265 (N_8265,N_7921,N_7579);
xnor U8266 (N_8266,N_7301,N_7850);
or U8267 (N_8267,N_7267,N_7657);
nor U8268 (N_8268,N_7672,N_7028);
nand U8269 (N_8269,N_7081,N_7992);
nand U8270 (N_8270,N_7859,N_7157);
xnor U8271 (N_8271,N_7476,N_7727);
or U8272 (N_8272,N_7805,N_7694);
nor U8273 (N_8273,N_7944,N_7605);
or U8274 (N_8274,N_7737,N_7182);
nor U8275 (N_8275,N_7121,N_7098);
nor U8276 (N_8276,N_7217,N_7362);
or U8277 (N_8277,N_7519,N_7520);
nand U8278 (N_8278,N_7164,N_7421);
nand U8279 (N_8279,N_7645,N_7908);
nand U8280 (N_8280,N_7300,N_7348);
nor U8281 (N_8281,N_7427,N_7146);
nand U8282 (N_8282,N_7665,N_7264);
xor U8283 (N_8283,N_7964,N_7442);
xnor U8284 (N_8284,N_7601,N_7635);
or U8285 (N_8285,N_7942,N_7242);
nand U8286 (N_8286,N_7878,N_7846);
nand U8287 (N_8287,N_7042,N_7445);
or U8288 (N_8288,N_7172,N_7248);
nor U8289 (N_8289,N_7329,N_7962);
or U8290 (N_8290,N_7018,N_7676);
nor U8291 (N_8291,N_7021,N_7899);
or U8292 (N_8292,N_7562,N_7560);
nand U8293 (N_8293,N_7822,N_7754);
nand U8294 (N_8294,N_7148,N_7536);
or U8295 (N_8295,N_7508,N_7422);
or U8296 (N_8296,N_7322,N_7426);
and U8297 (N_8297,N_7523,N_7443);
nand U8298 (N_8298,N_7623,N_7447);
nor U8299 (N_8299,N_7408,N_7870);
xor U8300 (N_8300,N_7675,N_7742);
xor U8301 (N_8301,N_7265,N_7165);
and U8302 (N_8302,N_7925,N_7342);
xnor U8303 (N_8303,N_7130,N_7133);
nor U8304 (N_8304,N_7197,N_7389);
xor U8305 (N_8305,N_7397,N_7374);
nand U8306 (N_8306,N_7013,N_7578);
xnor U8307 (N_8307,N_7690,N_7929);
nor U8308 (N_8308,N_7902,N_7948);
xor U8309 (N_8309,N_7573,N_7041);
and U8310 (N_8310,N_7711,N_7456);
xnor U8311 (N_8311,N_7849,N_7482);
or U8312 (N_8312,N_7823,N_7618);
xor U8313 (N_8313,N_7550,N_7498);
nand U8314 (N_8314,N_7696,N_7226);
and U8315 (N_8315,N_7132,N_7210);
nor U8316 (N_8316,N_7895,N_7237);
or U8317 (N_8317,N_7134,N_7763);
xor U8318 (N_8318,N_7752,N_7759);
xor U8319 (N_8319,N_7009,N_7387);
nor U8320 (N_8320,N_7600,N_7574);
nor U8321 (N_8321,N_7454,N_7521);
nand U8322 (N_8322,N_7535,N_7662);
xnor U8323 (N_8323,N_7484,N_7830);
or U8324 (N_8324,N_7338,N_7452);
nor U8325 (N_8325,N_7701,N_7509);
or U8326 (N_8326,N_7909,N_7692);
or U8327 (N_8327,N_7446,N_7238);
nand U8328 (N_8328,N_7693,N_7730);
nor U8329 (N_8329,N_7401,N_7669);
or U8330 (N_8330,N_7321,N_7976);
nor U8331 (N_8331,N_7787,N_7658);
nand U8332 (N_8332,N_7278,N_7364);
or U8333 (N_8333,N_7007,N_7045);
xor U8334 (N_8334,N_7744,N_7590);
xor U8335 (N_8335,N_7350,N_7191);
xnor U8336 (N_8336,N_7653,N_7949);
nor U8337 (N_8337,N_7621,N_7839);
and U8338 (N_8338,N_7708,N_7593);
and U8339 (N_8339,N_7261,N_7212);
nor U8340 (N_8340,N_7249,N_7679);
nand U8341 (N_8341,N_7126,N_7479);
and U8342 (N_8342,N_7746,N_7729);
nor U8343 (N_8343,N_7893,N_7505);
or U8344 (N_8344,N_7566,N_7416);
nand U8345 (N_8345,N_7044,N_7813);
or U8346 (N_8346,N_7012,N_7544);
xor U8347 (N_8347,N_7287,N_7555);
xor U8348 (N_8348,N_7492,N_7094);
xnor U8349 (N_8349,N_7837,N_7086);
or U8350 (N_8350,N_7915,N_7831);
nor U8351 (N_8351,N_7151,N_7642);
or U8352 (N_8352,N_7214,N_7501);
xor U8353 (N_8353,N_7567,N_7396);
or U8354 (N_8354,N_7762,N_7819);
or U8355 (N_8355,N_7181,N_7143);
or U8356 (N_8356,N_7659,N_7315);
and U8357 (N_8357,N_7206,N_7596);
and U8358 (N_8358,N_7239,N_7791);
and U8359 (N_8359,N_7344,N_7983);
and U8360 (N_8360,N_7538,N_7661);
and U8361 (N_8361,N_7572,N_7444);
nand U8362 (N_8362,N_7004,N_7464);
or U8363 (N_8363,N_7163,N_7470);
or U8364 (N_8364,N_7457,N_7768);
nor U8365 (N_8365,N_7038,N_7608);
or U8366 (N_8366,N_7058,N_7783);
nand U8367 (N_8367,N_7685,N_7591);
or U8368 (N_8368,N_7371,N_7598);
or U8369 (N_8369,N_7524,N_7770);
and U8370 (N_8370,N_7036,N_7667);
or U8371 (N_8371,N_7460,N_7225);
or U8372 (N_8372,N_7251,N_7923);
and U8373 (N_8373,N_7455,N_7810);
nor U8374 (N_8374,N_7760,N_7882);
nand U8375 (N_8375,N_7158,N_7997);
and U8376 (N_8376,N_7118,N_7833);
nor U8377 (N_8377,N_7137,N_7516);
and U8378 (N_8378,N_7472,N_7629);
nand U8379 (N_8379,N_7313,N_7061);
and U8380 (N_8380,N_7123,N_7379);
xor U8381 (N_8381,N_7991,N_7290);
xor U8382 (N_8382,N_7820,N_7340);
and U8383 (N_8383,N_7188,N_7985);
nand U8384 (N_8384,N_7207,N_7556);
nand U8385 (N_8385,N_7106,N_7785);
nand U8386 (N_8386,N_7848,N_7039);
nor U8387 (N_8387,N_7323,N_7136);
nand U8388 (N_8388,N_7201,N_7978);
and U8389 (N_8389,N_7488,N_7108);
and U8390 (N_8390,N_7358,N_7684);
xnor U8391 (N_8391,N_7346,N_7726);
or U8392 (N_8392,N_7381,N_7275);
nand U8393 (N_8393,N_7246,N_7253);
or U8394 (N_8394,N_7738,N_7357);
nor U8395 (N_8395,N_7678,N_7468);
xnor U8396 (N_8396,N_7361,N_7011);
nand U8397 (N_8397,N_7092,N_7100);
or U8398 (N_8398,N_7017,N_7502);
or U8399 (N_8399,N_7034,N_7352);
or U8400 (N_8400,N_7474,N_7095);
nand U8401 (N_8401,N_7681,N_7208);
or U8402 (N_8402,N_7325,N_7714);
nand U8403 (N_8403,N_7844,N_7990);
and U8404 (N_8404,N_7043,N_7876);
nand U8405 (N_8405,N_7723,N_7473);
or U8406 (N_8406,N_7869,N_7187);
or U8407 (N_8407,N_7963,N_7973);
nand U8408 (N_8408,N_7989,N_7798);
nand U8409 (N_8409,N_7391,N_7998);
xor U8410 (N_8410,N_7630,N_7794);
and U8411 (N_8411,N_7231,N_7938);
nand U8412 (N_8412,N_7576,N_7655);
or U8413 (N_8413,N_7812,N_7753);
xnor U8414 (N_8414,N_7037,N_7707);
nand U8415 (N_8415,N_7903,N_7000);
nor U8416 (N_8416,N_7260,N_7380);
or U8417 (N_8417,N_7395,N_7937);
nand U8418 (N_8418,N_7050,N_7896);
or U8419 (N_8419,N_7979,N_7924);
and U8420 (N_8420,N_7230,N_7129);
nor U8421 (N_8421,N_7886,N_7286);
xnor U8422 (N_8422,N_7946,N_7491);
nor U8423 (N_8423,N_7731,N_7815);
xnor U8424 (N_8424,N_7385,N_7419);
nor U8425 (N_8425,N_7879,N_7534);
nand U8426 (N_8426,N_7173,N_7568);
nor U8427 (N_8427,N_7328,N_7262);
nand U8428 (N_8428,N_7868,N_7068);
xor U8429 (N_8429,N_7811,N_7005);
and U8430 (N_8430,N_7049,N_7780);
and U8431 (N_8431,N_7318,N_7475);
or U8432 (N_8432,N_7486,N_7406);
nor U8433 (N_8433,N_7790,N_7834);
or U8434 (N_8434,N_7407,N_7431);
nor U8435 (N_8435,N_7015,N_7807);
xor U8436 (N_8436,N_7571,N_7020);
and U8437 (N_8437,N_7376,N_7111);
nor U8438 (N_8438,N_7062,N_7739);
or U8439 (N_8439,N_7786,N_7351);
xor U8440 (N_8440,N_7059,N_7917);
xnor U8441 (N_8441,N_7114,N_7345);
and U8442 (N_8442,N_7209,N_7966);
and U8443 (N_8443,N_7543,N_7597);
xnor U8444 (N_8444,N_7632,N_7531);
and U8445 (N_8445,N_7827,N_7633);
nor U8446 (N_8446,N_7233,N_7506);
xnor U8447 (N_8447,N_7485,N_7434);
nand U8448 (N_8448,N_7613,N_7080);
xnor U8449 (N_8449,N_7356,N_7258);
nand U8450 (N_8450,N_7124,N_7451);
nand U8451 (N_8451,N_7584,N_7244);
nand U8452 (N_8452,N_7429,N_7503);
nand U8453 (N_8453,N_7292,N_7243);
or U8454 (N_8454,N_7398,N_7383);
nand U8455 (N_8455,N_7467,N_7390);
nor U8456 (N_8456,N_7745,N_7772);
xnor U8457 (N_8457,N_7234,N_7088);
nand U8458 (N_8458,N_7220,N_7910);
and U8459 (N_8459,N_7252,N_7335);
nand U8460 (N_8460,N_7073,N_7981);
xor U8461 (N_8461,N_7057,N_7008);
nor U8462 (N_8462,N_7852,N_7782);
nand U8463 (N_8463,N_7441,N_7127);
xor U8464 (N_8464,N_7887,N_7149);
xor U8465 (N_8465,N_7311,N_7713);
or U8466 (N_8466,N_7826,N_7918);
nand U8467 (N_8467,N_7933,N_7104);
xnor U8468 (N_8468,N_7674,N_7091);
and U8469 (N_8469,N_7885,N_7324);
or U8470 (N_8470,N_7671,N_7494);
nor U8471 (N_8471,N_7919,N_7537);
xor U8472 (N_8472,N_7295,N_7588);
nand U8473 (N_8473,N_7959,N_7198);
or U8474 (N_8474,N_7355,N_7799);
xnor U8475 (N_8475,N_7462,N_7428);
or U8476 (N_8476,N_7546,N_7928);
xnor U8477 (N_8477,N_7065,N_7892);
or U8478 (N_8478,N_7382,N_7563);
and U8479 (N_8479,N_7602,N_7788);
nor U8480 (N_8480,N_7945,N_7053);
nand U8481 (N_8481,N_7901,N_7898);
or U8482 (N_8482,N_7585,N_7274);
and U8483 (N_8483,N_7995,N_7926);
nor U8484 (N_8484,N_7797,N_7776);
or U8485 (N_8485,N_7010,N_7450);
nor U8486 (N_8486,N_7875,N_7216);
and U8487 (N_8487,N_7958,N_7720);
nor U8488 (N_8488,N_7481,N_7078);
and U8489 (N_8489,N_7054,N_7611);
and U8490 (N_8490,N_7155,N_7255);
nand U8491 (N_8491,N_7832,N_7773);
xor U8492 (N_8492,N_7814,N_7257);
nor U8493 (N_8493,N_7298,N_7152);
and U8494 (N_8494,N_7522,N_7302);
and U8495 (N_8495,N_7499,N_7170);
xor U8496 (N_8496,N_7063,N_7654);
xor U8497 (N_8497,N_7478,N_7514);
and U8498 (N_8498,N_7766,N_7728);
nor U8499 (N_8499,N_7404,N_7511);
and U8500 (N_8500,N_7093,N_7939);
or U8501 (N_8501,N_7513,N_7067);
xor U8502 (N_8502,N_7268,N_7822);
xnor U8503 (N_8503,N_7639,N_7826);
nor U8504 (N_8504,N_7761,N_7883);
xnor U8505 (N_8505,N_7283,N_7317);
or U8506 (N_8506,N_7792,N_7551);
nor U8507 (N_8507,N_7004,N_7344);
nor U8508 (N_8508,N_7453,N_7745);
nand U8509 (N_8509,N_7783,N_7924);
xnor U8510 (N_8510,N_7265,N_7021);
nand U8511 (N_8511,N_7375,N_7102);
and U8512 (N_8512,N_7628,N_7782);
nor U8513 (N_8513,N_7803,N_7736);
xnor U8514 (N_8514,N_7634,N_7467);
nand U8515 (N_8515,N_7973,N_7062);
nand U8516 (N_8516,N_7253,N_7343);
xor U8517 (N_8517,N_7405,N_7869);
and U8518 (N_8518,N_7146,N_7141);
xnor U8519 (N_8519,N_7547,N_7368);
nand U8520 (N_8520,N_7329,N_7577);
and U8521 (N_8521,N_7830,N_7610);
nor U8522 (N_8522,N_7568,N_7014);
nor U8523 (N_8523,N_7250,N_7945);
xor U8524 (N_8524,N_7502,N_7911);
and U8525 (N_8525,N_7745,N_7792);
nor U8526 (N_8526,N_7217,N_7673);
or U8527 (N_8527,N_7660,N_7049);
nor U8528 (N_8528,N_7802,N_7547);
and U8529 (N_8529,N_7202,N_7153);
or U8530 (N_8530,N_7410,N_7838);
xor U8531 (N_8531,N_7996,N_7005);
or U8532 (N_8532,N_7065,N_7914);
xnor U8533 (N_8533,N_7704,N_7262);
and U8534 (N_8534,N_7268,N_7561);
or U8535 (N_8535,N_7793,N_7335);
or U8536 (N_8536,N_7830,N_7957);
nor U8537 (N_8537,N_7958,N_7334);
nor U8538 (N_8538,N_7447,N_7383);
xor U8539 (N_8539,N_7820,N_7495);
xor U8540 (N_8540,N_7352,N_7722);
xnor U8541 (N_8541,N_7190,N_7252);
nand U8542 (N_8542,N_7721,N_7453);
xor U8543 (N_8543,N_7862,N_7802);
or U8544 (N_8544,N_7885,N_7601);
nand U8545 (N_8545,N_7483,N_7113);
nor U8546 (N_8546,N_7624,N_7731);
nand U8547 (N_8547,N_7307,N_7183);
nand U8548 (N_8548,N_7884,N_7746);
xnor U8549 (N_8549,N_7388,N_7303);
and U8550 (N_8550,N_7315,N_7482);
nand U8551 (N_8551,N_7176,N_7273);
xor U8552 (N_8552,N_7696,N_7461);
xnor U8553 (N_8553,N_7337,N_7169);
or U8554 (N_8554,N_7928,N_7573);
nor U8555 (N_8555,N_7760,N_7776);
and U8556 (N_8556,N_7598,N_7475);
xor U8557 (N_8557,N_7540,N_7427);
and U8558 (N_8558,N_7855,N_7058);
xnor U8559 (N_8559,N_7741,N_7091);
and U8560 (N_8560,N_7885,N_7339);
xnor U8561 (N_8561,N_7733,N_7771);
or U8562 (N_8562,N_7561,N_7154);
nand U8563 (N_8563,N_7454,N_7499);
and U8564 (N_8564,N_7928,N_7322);
nor U8565 (N_8565,N_7238,N_7660);
nand U8566 (N_8566,N_7582,N_7343);
xnor U8567 (N_8567,N_7160,N_7116);
and U8568 (N_8568,N_7525,N_7377);
or U8569 (N_8569,N_7034,N_7134);
nand U8570 (N_8570,N_7408,N_7325);
xor U8571 (N_8571,N_7488,N_7490);
or U8572 (N_8572,N_7642,N_7712);
and U8573 (N_8573,N_7159,N_7790);
or U8574 (N_8574,N_7477,N_7361);
or U8575 (N_8575,N_7315,N_7337);
nand U8576 (N_8576,N_7540,N_7169);
or U8577 (N_8577,N_7019,N_7393);
nor U8578 (N_8578,N_7798,N_7513);
and U8579 (N_8579,N_7162,N_7042);
xor U8580 (N_8580,N_7333,N_7779);
or U8581 (N_8581,N_7333,N_7487);
nand U8582 (N_8582,N_7368,N_7097);
or U8583 (N_8583,N_7067,N_7939);
or U8584 (N_8584,N_7078,N_7805);
xor U8585 (N_8585,N_7020,N_7734);
nand U8586 (N_8586,N_7720,N_7920);
xor U8587 (N_8587,N_7979,N_7143);
xnor U8588 (N_8588,N_7145,N_7992);
and U8589 (N_8589,N_7958,N_7307);
or U8590 (N_8590,N_7864,N_7808);
and U8591 (N_8591,N_7736,N_7061);
xnor U8592 (N_8592,N_7632,N_7077);
xor U8593 (N_8593,N_7918,N_7041);
or U8594 (N_8594,N_7390,N_7083);
xor U8595 (N_8595,N_7783,N_7093);
nand U8596 (N_8596,N_7636,N_7820);
nor U8597 (N_8597,N_7019,N_7215);
nor U8598 (N_8598,N_7646,N_7892);
and U8599 (N_8599,N_7518,N_7203);
xor U8600 (N_8600,N_7752,N_7823);
nor U8601 (N_8601,N_7877,N_7558);
xor U8602 (N_8602,N_7336,N_7473);
and U8603 (N_8603,N_7043,N_7372);
xnor U8604 (N_8604,N_7635,N_7093);
and U8605 (N_8605,N_7711,N_7727);
or U8606 (N_8606,N_7710,N_7102);
xor U8607 (N_8607,N_7693,N_7545);
and U8608 (N_8608,N_7003,N_7173);
or U8609 (N_8609,N_7840,N_7952);
nor U8610 (N_8610,N_7163,N_7545);
or U8611 (N_8611,N_7138,N_7176);
xor U8612 (N_8612,N_7690,N_7313);
nand U8613 (N_8613,N_7985,N_7874);
xnor U8614 (N_8614,N_7242,N_7467);
nor U8615 (N_8615,N_7747,N_7791);
nand U8616 (N_8616,N_7470,N_7564);
nor U8617 (N_8617,N_7479,N_7480);
or U8618 (N_8618,N_7711,N_7448);
nor U8619 (N_8619,N_7378,N_7753);
nor U8620 (N_8620,N_7403,N_7405);
xor U8621 (N_8621,N_7514,N_7195);
nor U8622 (N_8622,N_7348,N_7404);
or U8623 (N_8623,N_7834,N_7520);
nor U8624 (N_8624,N_7607,N_7381);
nand U8625 (N_8625,N_7052,N_7768);
nand U8626 (N_8626,N_7103,N_7029);
xnor U8627 (N_8627,N_7668,N_7916);
xnor U8628 (N_8628,N_7588,N_7489);
or U8629 (N_8629,N_7457,N_7124);
nor U8630 (N_8630,N_7257,N_7256);
xnor U8631 (N_8631,N_7910,N_7282);
and U8632 (N_8632,N_7184,N_7134);
nand U8633 (N_8633,N_7071,N_7091);
or U8634 (N_8634,N_7871,N_7013);
nor U8635 (N_8635,N_7711,N_7343);
and U8636 (N_8636,N_7129,N_7626);
and U8637 (N_8637,N_7602,N_7131);
xnor U8638 (N_8638,N_7087,N_7816);
and U8639 (N_8639,N_7858,N_7087);
nand U8640 (N_8640,N_7669,N_7388);
xor U8641 (N_8641,N_7186,N_7586);
and U8642 (N_8642,N_7184,N_7845);
nor U8643 (N_8643,N_7018,N_7182);
xor U8644 (N_8644,N_7719,N_7035);
and U8645 (N_8645,N_7730,N_7532);
xnor U8646 (N_8646,N_7901,N_7766);
and U8647 (N_8647,N_7289,N_7762);
nor U8648 (N_8648,N_7421,N_7602);
and U8649 (N_8649,N_7927,N_7344);
and U8650 (N_8650,N_7060,N_7991);
nand U8651 (N_8651,N_7665,N_7039);
or U8652 (N_8652,N_7274,N_7026);
xor U8653 (N_8653,N_7241,N_7010);
and U8654 (N_8654,N_7886,N_7248);
nand U8655 (N_8655,N_7527,N_7880);
nand U8656 (N_8656,N_7136,N_7460);
and U8657 (N_8657,N_7441,N_7482);
xor U8658 (N_8658,N_7154,N_7436);
nand U8659 (N_8659,N_7875,N_7153);
nand U8660 (N_8660,N_7533,N_7235);
nand U8661 (N_8661,N_7772,N_7378);
and U8662 (N_8662,N_7350,N_7170);
xnor U8663 (N_8663,N_7870,N_7057);
xnor U8664 (N_8664,N_7710,N_7125);
nor U8665 (N_8665,N_7844,N_7065);
or U8666 (N_8666,N_7152,N_7674);
and U8667 (N_8667,N_7160,N_7122);
or U8668 (N_8668,N_7089,N_7895);
and U8669 (N_8669,N_7645,N_7513);
nand U8670 (N_8670,N_7785,N_7597);
nor U8671 (N_8671,N_7331,N_7854);
and U8672 (N_8672,N_7497,N_7331);
or U8673 (N_8673,N_7304,N_7778);
and U8674 (N_8674,N_7386,N_7095);
nand U8675 (N_8675,N_7405,N_7929);
and U8676 (N_8676,N_7143,N_7846);
nor U8677 (N_8677,N_7794,N_7061);
nor U8678 (N_8678,N_7516,N_7165);
and U8679 (N_8679,N_7395,N_7121);
xnor U8680 (N_8680,N_7178,N_7987);
nand U8681 (N_8681,N_7590,N_7799);
nand U8682 (N_8682,N_7955,N_7260);
or U8683 (N_8683,N_7330,N_7379);
and U8684 (N_8684,N_7394,N_7334);
nand U8685 (N_8685,N_7619,N_7387);
nor U8686 (N_8686,N_7715,N_7026);
nor U8687 (N_8687,N_7331,N_7411);
and U8688 (N_8688,N_7455,N_7869);
xor U8689 (N_8689,N_7298,N_7117);
nand U8690 (N_8690,N_7355,N_7917);
xor U8691 (N_8691,N_7533,N_7201);
and U8692 (N_8692,N_7631,N_7849);
xnor U8693 (N_8693,N_7508,N_7074);
nand U8694 (N_8694,N_7893,N_7934);
xnor U8695 (N_8695,N_7821,N_7597);
or U8696 (N_8696,N_7253,N_7221);
xnor U8697 (N_8697,N_7901,N_7803);
xor U8698 (N_8698,N_7249,N_7572);
xnor U8699 (N_8699,N_7062,N_7186);
nor U8700 (N_8700,N_7809,N_7514);
and U8701 (N_8701,N_7313,N_7230);
nor U8702 (N_8702,N_7195,N_7662);
and U8703 (N_8703,N_7600,N_7093);
nand U8704 (N_8704,N_7024,N_7967);
and U8705 (N_8705,N_7020,N_7614);
and U8706 (N_8706,N_7928,N_7673);
xor U8707 (N_8707,N_7057,N_7802);
and U8708 (N_8708,N_7143,N_7478);
nand U8709 (N_8709,N_7574,N_7496);
nand U8710 (N_8710,N_7272,N_7603);
or U8711 (N_8711,N_7867,N_7916);
and U8712 (N_8712,N_7065,N_7234);
nor U8713 (N_8713,N_7967,N_7449);
nor U8714 (N_8714,N_7089,N_7883);
nand U8715 (N_8715,N_7413,N_7786);
nor U8716 (N_8716,N_7116,N_7940);
nor U8717 (N_8717,N_7738,N_7322);
and U8718 (N_8718,N_7962,N_7702);
xor U8719 (N_8719,N_7515,N_7387);
xnor U8720 (N_8720,N_7039,N_7700);
or U8721 (N_8721,N_7811,N_7621);
nor U8722 (N_8722,N_7440,N_7168);
and U8723 (N_8723,N_7806,N_7242);
or U8724 (N_8724,N_7234,N_7846);
and U8725 (N_8725,N_7179,N_7350);
and U8726 (N_8726,N_7298,N_7404);
nand U8727 (N_8727,N_7365,N_7491);
nand U8728 (N_8728,N_7655,N_7701);
or U8729 (N_8729,N_7739,N_7781);
xnor U8730 (N_8730,N_7786,N_7075);
and U8731 (N_8731,N_7491,N_7451);
nand U8732 (N_8732,N_7615,N_7144);
and U8733 (N_8733,N_7460,N_7950);
and U8734 (N_8734,N_7545,N_7478);
or U8735 (N_8735,N_7309,N_7207);
or U8736 (N_8736,N_7632,N_7983);
or U8737 (N_8737,N_7116,N_7958);
or U8738 (N_8738,N_7030,N_7207);
xnor U8739 (N_8739,N_7177,N_7075);
nor U8740 (N_8740,N_7843,N_7907);
or U8741 (N_8741,N_7219,N_7762);
and U8742 (N_8742,N_7414,N_7364);
nor U8743 (N_8743,N_7087,N_7953);
nand U8744 (N_8744,N_7845,N_7987);
xor U8745 (N_8745,N_7045,N_7914);
and U8746 (N_8746,N_7983,N_7386);
nor U8747 (N_8747,N_7717,N_7843);
nor U8748 (N_8748,N_7145,N_7231);
nor U8749 (N_8749,N_7697,N_7298);
nand U8750 (N_8750,N_7419,N_7977);
and U8751 (N_8751,N_7920,N_7310);
and U8752 (N_8752,N_7442,N_7375);
and U8753 (N_8753,N_7302,N_7638);
xor U8754 (N_8754,N_7494,N_7351);
nand U8755 (N_8755,N_7084,N_7270);
nand U8756 (N_8756,N_7980,N_7778);
nor U8757 (N_8757,N_7110,N_7100);
nand U8758 (N_8758,N_7592,N_7899);
or U8759 (N_8759,N_7228,N_7424);
nand U8760 (N_8760,N_7703,N_7188);
and U8761 (N_8761,N_7867,N_7941);
nand U8762 (N_8762,N_7786,N_7249);
nor U8763 (N_8763,N_7668,N_7182);
or U8764 (N_8764,N_7628,N_7617);
xnor U8765 (N_8765,N_7449,N_7045);
and U8766 (N_8766,N_7234,N_7502);
nor U8767 (N_8767,N_7913,N_7552);
or U8768 (N_8768,N_7011,N_7621);
nor U8769 (N_8769,N_7452,N_7548);
or U8770 (N_8770,N_7053,N_7426);
or U8771 (N_8771,N_7948,N_7855);
xnor U8772 (N_8772,N_7745,N_7207);
nand U8773 (N_8773,N_7848,N_7033);
and U8774 (N_8774,N_7360,N_7405);
nor U8775 (N_8775,N_7900,N_7595);
xnor U8776 (N_8776,N_7221,N_7768);
nor U8777 (N_8777,N_7115,N_7571);
and U8778 (N_8778,N_7338,N_7351);
or U8779 (N_8779,N_7520,N_7602);
nor U8780 (N_8780,N_7202,N_7329);
and U8781 (N_8781,N_7190,N_7662);
or U8782 (N_8782,N_7009,N_7403);
xor U8783 (N_8783,N_7908,N_7715);
xor U8784 (N_8784,N_7151,N_7773);
nor U8785 (N_8785,N_7839,N_7959);
nor U8786 (N_8786,N_7799,N_7898);
xor U8787 (N_8787,N_7038,N_7861);
nand U8788 (N_8788,N_7756,N_7642);
nor U8789 (N_8789,N_7380,N_7926);
or U8790 (N_8790,N_7261,N_7133);
nor U8791 (N_8791,N_7287,N_7580);
xor U8792 (N_8792,N_7356,N_7701);
xor U8793 (N_8793,N_7675,N_7044);
xor U8794 (N_8794,N_7585,N_7627);
and U8795 (N_8795,N_7783,N_7031);
nor U8796 (N_8796,N_7564,N_7177);
nand U8797 (N_8797,N_7063,N_7520);
and U8798 (N_8798,N_7145,N_7412);
or U8799 (N_8799,N_7868,N_7158);
and U8800 (N_8800,N_7933,N_7661);
nand U8801 (N_8801,N_7142,N_7088);
nor U8802 (N_8802,N_7441,N_7003);
and U8803 (N_8803,N_7937,N_7229);
nor U8804 (N_8804,N_7987,N_7477);
nand U8805 (N_8805,N_7693,N_7795);
xor U8806 (N_8806,N_7544,N_7469);
nand U8807 (N_8807,N_7837,N_7663);
xnor U8808 (N_8808,N_7567,N_7758);
nor U8809 (N_8809,N_7435,N_7417);
xnor U8810 (N_8810,N_7614,N_7766);
nand U8811 (N_8811,N_7241,N_7176);
xor U8812 (N_8812,N_7560,N_7331);
nor U8813 (N_8813,N_7707,N_7527);
nor U8814 (N_8814,N_7218,N_7410);
xor U8815 (N_8815,N_7908,N_7886);
xnor U8816 (N_8816,N_7436,N_7378);
nand U8817 (N_8817,N_7409,N_7333);
or U8818 (N_8818,N_7776,N_7628);
and U8819 (N_8819,N_7241,N_7348);
and U8820 (N_8820,N_7415,N_7861);
and U8821 (N_8821,N_7010,N_7701);
or U8822 (N_8822,N_7106,N_7922);
or U8823 (N_8823,N_7156,N_7114);
xor U8824 (N_8824,N_7172,N_7760);
or U8825 (N_8825,N_7444,N_7063);
or U8826 (N_8826,N_7731,N_7219);
and U8827 (N_8827,N_7322,N_7156);
and U8828 (N_8828,N_7103,N_7101);
nand U8829 (N_8829,N_7954,N_7304);
and U8830 (N_8830,N_7318,N_7614);
xnor U8831 (N_8831,N_7748,N_7058);
nor U8832 (N_8832,N_7014,N_7081);
xor U8833 (N_8833,N_7744,N_7437);
nand U8834 (N_8834,N_7190,N_7054);
xnor U8835 (N_8835,N_7597,N_7138);
nor U8836 (N_8836,N_7346,N_7702);
nand U8837 (N_8837,N_7032,N_7499);
and U8838 (N_8838,N_7295,N_7052);
nor U8839 (N_8839,N_7183,N_7127);
or U8840 (N_8840,N_7953,N_7868);
nor U8841 (N_8841,N_7712,N_7166);
xor U8842 (N_8842,N_7367,N_7144);
xor U8843 (N_8843,N_7593,N_7766);
nor U8844 (N_8844,N_7664,N_7984);
or U8845 (N_8845,N_7480,N_7708);
or U8846 (N_8846,N_7901,N_7833);
and U8847 (N_8847,N_7035,N_7357);
and U8848 (N_8848,N_7866,N_7314);
or U8849 (N_8849,N_7764,N_7386);
or U8850 (N_8850,N_7675,N_7764);
or U8851 (N_8851,N_7501,N_7820);
or U8852 (N_8852,N_7672,N_7311);
or U8853 (N_8853,N_7911,N_7126);
xor U8854 (N_8854,N_7576,N_7241);
and U8855 (N_8855,N_7489,N_7102);
nand U8856 (N_8856,N_7060,N_7112);
or U8857 (N_8857,N_7897,N_7221);
nand U8858 (N_8858,N_7959,N_7318);
nor U8859 (N_8859,N_7798,N_7951);
nand U8860 (N_8860,N_7438,N_7269);
nand U8861 (N_8861,N_7804,N_7911);
xor U8862 (N_8862,N_7554,N_7675);
nand U8863 (N_8863,N_7079,N_7798);
or U8864 (N_8864,N_7563,N_7431);
or U8865 (N_8865,N_7482,N_7610);
nor U8866 (N_8866,N_7204,N_7036);
xnor U8867 (N_8867,N_7124,N_7860);
nand U8868 (N_8868,N_7211,N_7242);
xor U8869 (N_8869,N_7508,N_7736);
nand U8870 (N_8870,N_7282,N_7837);
nand U8871 (N_8871,N_7532,N_7271);
xnor U8872 (N_8872,N_7016,N_7994);
nand U8873 (N_8873,N_7041,N_7506);
or U8874 (N_8874,N_7984,N_7252);
nor U8875 (N_8875,N_7075,N_7736);
xnor U8876 (N_8876,N_7731,N_7589);
xor U8877 (N_8877,N_7228,N_7020);
and U8878 (N_8878,N_7733,N_7032);
or U8879 (N_8879,N_7757,N_7962);
and U8880 (N_8880,N_7140,N_7601);
or U8881 (N_8881,N_7651,N_7692);
and U8882 (N_8882,N_7323,N_7207);
nor U8883 (N_8883,N_7490,N_7259);
and U8884 (N_8884,N_7759,N_7482);
xnor U8885 (N_8885,N_7844,N_7208);
nor U8886 (N_8886,N_7988,N_7250);
xnor U8887 (N_8887,N_7360,N_7978);
and U8888 (N_8888,N_7548,N_7953);
xnor U8889 (N_8889,N_7964,N_7986);
or U8890 (N_8890,N_7423,N_7669);
nand U8891 (N_8891,N_7646,N_7833);
or U8892 (N_8892,N_7764,N_7960);
xor U8893 (N_8893,N_7758,N_7879);
or U8894 (N_8894,N_7686,N_7471);
or U8895 (N_8895,N_7996,N_7642);
or U8896 (N_8896,N_7736,N_7281);
nor U8897 (N_8897,N_7936,N_7376);
or U8898 (N_8898,N_7611,N_7132);
and U8899 (N_8899,N_7874,N_7106);
nand U8900 (N_8900,N_7260,N_7656);
or U8901 (N_8901,N_7939,N_7625);
or U8902 (N_8902,N_7436,N_7675);
nand U8903 (N_8903,N_7945,N_7101);
xor U8904 (N_8904,N_7963,N_7194);
xnor U8905 (N_8905,N_7008,N_7391);
and U8906 (N_8906,N_7037,N_7837);
nand U8907 (N_8907,N_7597,N_7154);
nand U8908 (N_8908,N_7100,N_7632);
xor U8909 (N_8909,N_7439,N_7267);
nor U8910 (N_8910,N_7526,N_7939);
nor U8911 (N_8911,N_7307,N_7477);
and U8912 (N_8912,N_7256,N_7927);
nor U8913 (N_8913,N_7975,N_7710);
nor U8914 (N_8914,N_7192,N_7913);
nand U8915 (N_8915,N_7291,N_7227);
nor U8916 (N_8916,N_7408,N_7480);
nor U8917 (N_8917,N_7257,N_7940);
and U8918 (N_8918,N_7411,N_7505);
xor U8919 (N_8919,N_7901,N_7878);
xor U8920 (N_8920,N_7663,N_7383);
xnor U8921 (N_8921,N_7213,N_7853);
nor U8922 (N_8922,N_7798,N_7043);
or U8923 (N_8923,N_7955,N_7540);
xnor U8924 (N_8924,N_7893,N_7023);
or U8925 (N_8925,N_7497,N_7749);
xnor U8926 (N_8926,N_7187,N_7858);
xor U8927 (N_8927,N_7183,N_7098);
nand U8928 (N_8928,N_7995,N_7028);
and U8929 (N_8929,N_7422,N_7695);
xor U8930 (N_8930,N_7042,N_7300);
nor U8931 (N_8931,N_7233,N_7165);
and U8932 (N_8932,N_7108,N_7684);
xor U8933 (N_8933,N_7673,N_7961);
or U8934 (N_8934,N_7737,N_7317);
nor U8935 (N_8935,N_7129,N_7539);
xor U8936 (N_8936,N_7472,N_7821);
or U8937 (N_8937,N_7580,N_7947);
nand U8938 (N_8938,N_7782,N_7703);
and U8939 (N_8939,N_7898,N_7262);
xor U8940 (N_8940,N_7107,N_7510);
or U8941 (N_8941,N_7444,N_7332);
nor U8942 (N_8942,N_7419,N_7741);
or U8943 (N_8943,N_7742,N_7150);
nor U8944 (N_8944,N_7842,N_7569);
nor U8945 (N_8945,N_7737,N_7428);
or U8946 (N_8946,N_7573,N_7182);
or U8947 (N_8947,N_7391,N_7185);
xnor U8948 (N_8948,N_7812,N_7609);
and U8949 (N_8949,N_7227,N_7871);
and U8950 (N_8950,N_7280,N_7999);
nand U8951 (N_8951,N_7932,N_7319);
nand U8952 (N_8952,N_7657,N_7363);
nor U8953 (N_8953,N_7328,N_7097);
nand U8954 (N_8954,N_7844,N_7040);
and U8955 (N_8955,N_7944,N_7642);
nor U8956 (N_8956,N_7897,N_7205);
xnor U8957 (N_8957,N_7952,N_7992);
xor U8958 (N_8958,N_7308,N_7420);
xor U8959 (N_8959,N_7174,N_7966);
nand U8960 (N_8960,N_7456,N_7208);
and U8961 (N_8961,N_7940,N_7619);
nand U8962 (N_8962,N_7666,N_7882);
xnor U8963 (N_8963,N_7710,N_7284);
or U8964 (N_8964,N_7850,N_7017);
nor U8965 (N_8965,N_7081,N_7710);
and U8966 (N_8966,N_7570,N_7417);
xor U8967 (N_8967,N_7732,N_7032);
xor U8968 (N_8968,N_7293,N_7163);
or U8969 (N_8969,N_7692,N_7622);
and U8970 (N_8970,N_7800,N_7279);
nor U8971 (N_8971,N_7783,N_7573);
xnor U8972 (N_8972,N_7767,N_7773);
xnor U8973 (N_8973,N_7216,N_7120);
and U8974 (N_8974,N_7165,N_7946);
or U8975 (N_8975,N_7936,N_7758);
nand U8976 (N_8976,N_7980,N_7929);
or U8977 (N_8977,N_7765,N_7579);
and U8978 (N_8978,N_7002,N_7459);
nand U8979 (N_8979,N_7609,N_7195);
and U8980 (N_8980,N_7759,N_7374);
nand U8981 (N_8981,N_7685,N_7818);
or U8982 (N_8982,N_7203,N_7787);
nor U8983 (N_8983,N_7940,N_7520);
or U8984 (N_8984,N_7820,N_7124);
xor U8985 (N_8985,N_7583,N_7523);
nor U8986 (N_8986,N_7811,N_7864);
xnor U8987 (N_8987,N_7473,N_7768);
or U8988 (N_8988,N_7393,N_7447);
or U8989 (N_8989,N_7891,N_7313);
and U8990 (N_8990,N_7464,N_7494);
nand U8991 (N_8991,N_7211,N_7551);
and U8992 (N_8992,N_7271,N_7014);
nand U8993 (N_8993,N_7266,N_7508);
and U8994 (N_8994,N_7382,N_7040);
xor U8995 (N_8995,N_7183,N_7166);
and U8996 (N_8996,N_7189,N_7703);
xor U8997 (N_8997,N_7124,N_7370);
nor U8998 (N_8998,N_7326,N_7419);
nand U8999 (N_8999,N_7039,N_7122);
and U9000 (N_9000,N_8379,N_8014);
and U9001 (N_9001,N_8386,N_8197);
xnor U9002 (N_9002,N_8237,N_8545);
xor U9003 (N_9003,N_8216,N_8271);
nor U9004 (N_9004,N_8221,N_8187);
and U9005 (N_9005,N_8005,N_8891);
and U9006 (N_9006,N_8722,N_8504);
or U9007 (N_9007,N_8611,N_8117);
xor U9008 (N_9008,N_8287,N_8240);
and U9009 (N_9009,N_8487,N_8367);
nand U9010 (N_9010,N_8010,N_8823);
xor U9011 (N_9011,N_8936,N_8046);
xnor U9012 (N_9012,N_8517,N_8736);
xnor U9013 (N_9013,N_8459,N_8508);
and U9014 (N_9014,N_8316,N_8861);
and U9015 (N_9015,N_8866,N_8514);
xor U9016 (N_9016,N_8509,N_8161);
or U9017 (N_9017,N_8338,N_8687);
nand U9018 (N_9018,N_8085,N_8002);
nor U9019 (N_9019,N_8909,N_8147);
and U9020 (N_9020,N_8697,N_8884);
and U9021 (N_9021,N_8908,N_8818);
or U9022 (N_9022,N_8118,N_8346);
nor U9023 (N_9023,N_8901,N_8801);
and U9024 (N_9024,N_8050,N_8232);
xnor U9025 (N_9025,N_8427,N_8448);
nand U9026 (N_9026,N_8036,N_8586);
nand U9027 (N_9027,N_8870,N_8612);
xnor U9028 (N_9028,N_8820,N_8821);
nor U9029 (N_9029,N_8407,N_8279);
xnor U9030 (N_9030,N_8369,N_8879);
nand U9031 (N_9031,N_8443,N_8344);
nand U9032 (N_9032,N_8618,N_8872);
and U9033 (N_9033,N_8852,N_8965);
nand U9034 (N_9034,N_8079,N_8138);
or U9035 (N_9035,N_8315,N_8084);
or U9036 (N_9036,N_8393,N_8871);
or U9037 (N_9037,N_8451,N_8156);
nor U9038 (N_9038,N_8745,N_8293);
or U9039 (N_9039,N_8834,N_8840);
xnor U9040 (N_9040,N_8549,N_8710);
nor U9041 (N_9041,N_8602,N_8247);
or U9042 (N_9042,N_8321,N_8996);
nand U9043 (N_9043,N_8771,N_8806);
xor U9044 (N_9044,N_8000,N_8172);
nor U9045 (N_9045,N_8923,N_8382);
nand U9046 (N_9046,N_8839,N_8640);
and U9047 (N_9047,N_8211,N_8072);
xnor U9048 (N_9048,N_8844,N_8385);
nor U9049 (N_9049,N_8045,N_8998);
and U9050 (N_9050,N_8756,N_8564);
nand U9051 (N_9051,N_8660,N_8658);
or U9052 (N_9052,N_8554,N_8431);
and U9053 (N_9053,N_8828,N_8888);
nor U9054 (N_9054,N_8902,N_8260);
nand U9055 (N_9055,N_8668,N_8097);
xor U9056 (N_9056,N_8935,N_8470);
xor U9057 (N_9057,N_8921,N_8882);
nor U9058 (N_9058,N_8191,N_8966);
nand U9059 (N_9059,N_8850,N_8140);
xnor U9060 (N_9060,N_8467,N_8877);
nand U9061 (N_9061,N_8328,N_8111);
nand U9062 (N_9062,N_8088,N_8686);
and U9063 (N_9063,N_8160,N_8121);
xnor U9064 (N_9064,N_8146,N_8066);
nor U9065 (N_9065,N_8957,N_8536);
nand U9066 (N_9066,N_8592,N_8927);
xor U9067 (N_9067,N_8725,N_8241);
and U9068 (N_9068,N_8265,N_8083);
or U9069 (N_9069,N_8358,N_8974);
nand U9070 (N_9070,N_8842,N_8700);
and U9071 (N_9071,N_8651,N_8123);
or U9072 (N_9072,N_8423,N_8044);
xor U9073 (N_9073,N_8238,N_8661);
xor U9074 (N_9074,N_8062,N_8408);
nor U9075 (N_9075,N_8421,N_8707);
and U9076 (N_9076,N_8254,N_8474);
or U9077 (N_9077,N_8567,N_8009);
and U9078 (N_9078,N_8665,N_8411);
xnor U9079 (N_9079,N_8306,N_8814);
nor U9080 (N_9080,N_8483,N_8028);
xnor U9081 (N_9081,N_8911,N_8772);
xnor U9082 (N_9082,N_8049,N_8548);
xnor U9083 (N_9083,N_8460,N_8994);
and U9084 (N_9084,N_8377,N_8634);
or U9085 (N_9085,N_8750,N_8115);
xnor U9086 (N_9086,N_8414,N_8506);
xor U9087 (N_9087,N_8026,N_8737);
nand U9088 (N_9088,N_8173,N_8288);
xnor U9089 (N_9089,N_8167,N_8067);
and U9090 (N_9090,N_8922,N_8827);
xnor U9091 (N_9091,N_8630,N_8732);
and U9092 (N_9092,N_8071,N_8323);
and U9093 (N_9093,N_8657,N_8712);
and U9094 (N_9094,N_8304,N_8301);
xor U9095 (N_9095,N_8845,N_8929);
nand U9096 (N_9096,N_8094,N_8944);
xor U9097 (N_9097,N_8595,N_8069);
nand U9098 (N_9098,N_8993,N_8533);
nor U9099 (N_9099,N_8142,N_8486);
xor U9100 (N_9100,N_8347,N_8212);
or U9101 (N_9101,N_8859,N_8199);
nand U9102 (N_9102,N_8790,N_8838);
xnor U9103 (N_9103,N_8370,N_8616);
nor U9104 (N_9104,N_8194,N_8125);
and U9105 (N_9105,N_8916,N_8163);
xor U9106 (N_9106,N_8782,N_8724);
or U9107 (N_9107,N_8652,N_8319);
nand U9108 (N_9108,N_8349,N_8610);
nor U9109 (N_9109,N_8468,N_8190);
and U9110 (N_9110,N_8638,N_8366);
nor U9111 (N_9111,N_8777,N_8297);
nor U9112 (N_9112,N_8626,N_8130);
or U9113 (N_9113,N_8149,N_8256);
xor U9114 (N_9114,N_8875,N_8796);
xor U9115 (N_9115,N_8954,N_8720);
and U9116 (N_9116,N_8461,N_8268);
nand U9117 (N_9117,N_8113,N_8792);
and U9118 (N_9118,N_8332,N_8562);
xor U9119 (N_9119,N_8865,N_8357);
nor U9120 (N_9120,N_8734,N_8647);
nor U9121 (N_9121,N_8608,N_8703);
and U9122 (N_9122,N_8495,N_8477);
xnor U9123 (N_9123,N_8698,N_8644);
and U9124 (N_9124,N_8299,N_8598);
nor U9125 (N_9125,N_8885,N_8089);
nand U9126 (N_9126,N_8534,N_8793);
nor U9127 (N_9127,N_8261,N_8699);
nor U9128 (N_9128,N_8714,N_8503);
and U9129 (N_9129,N_8368,N_8206);
nand U9130 (N_9130,N_8995,N_8914);
and U9131 (N_9131,N_8223,N_8109);
xor U9132 (N_9132,N_8807,N_8433);
nor U9133 (N_9133,N_8479,N_8103);
and U9134 (N_9134,N_8339,N_8422);
and U9135 (N_9135,N_8182,N_8532);
nand U9136 (N_9136,N_8258,N_8550);
and U9137 (N_9137,N_8589,N_8677);
xor U9138 (N_9138,N_8526,N_8057);
nand U9139 (N_9139,N_8558,N_8063);
or U9140 (N_9140,N_8091,N_8466);
or U9141 (N_9141,N_8054,N_8680);
xor U9142 (N_9142,N_8544,N_8267);
nor U9143 (N_9143,N_8184,N_8999);
xor U9144 (N_9144,N_8195,N_8437);
xnor U9145 (N_9145,N_8531,N_8711);
nand U9146 (N_9146,N_8308,N_8294);
nand U9147 (N_9147,N_8607,N_8336);
and U9148 (N_9148,N_8624,N_8119);
and U9149 (N_9149,N_8235,N_8799);
and U9150 (N_9150,N_8555,N_8372);
or U9151 (N_9151,N_8900,N_8296);
nand U9152 (N_9152,N_8064,N_8101);
or U9153 (N_9153,N_8579,N_8689);
nand U9154 (N_9154,N_8629,N_8786);
and U9155 (N_9155,N_8869,N_8354);
nor U9156 (N_9156,N_8401,N_8769);
nor U9157 (N_9157,N_8345,N_8748);
nand U9158 (N_9158,N_8484,N_8371);
xor U9159 (N_9159,N_8918,N_8374);
nor U9160 (N_9160,N_8924,N_8501);
nand U9161 (N_9161,N_8632,N_8619);
and U9162 (N_9162,N_8763,N_8383);
nand U9163 (N_9163,N_8179,N_8021);
xnor U9164 (N_9164,N_8874,N_8798);
nand U9165 (N_9165,N_8150,N_8376);
or U9166 (N_9166,N_8243,N_8024);
nand U9167 (N_9167,N_8942,N_8953);
nand U9168 (N_9168,N_8096,N_8389);
nor U9169 (N_9169,N_8655,N_8442);
or U9170 (N_9170,N_8410,N_8982);
or U9171 (N_9171,N_8497,N_8648);
nor U9172 (N_9172,N_8300,N_8810);
nor U9173 (N_9173,N_8073,N_8569);
and U9174 (N_9174,N_8087,N_8694);
nor U9175 (N_9175,N_8858,N_8717);
and U9176 (N_9176,N_8018,N_8582);
or U9177 (N_9177,N_8042,N_8362);
nor U9178 (N_9178,N_8090,N_8963);
and U9179 (N_9179,N_8220,N_8566);
xor U9180 (N_9180,N_8170,N_8473);
and U9181 (N_9181,N_8500,N_8990);
and U9182 (N_9182,N_8100,N_8832);
xnor U9183 (N_9183,N_8975,N_8540);
nor U9184 (N_9184,N_8037,N_8274);
or U9185 (N_9185,N_8812,N_8061);
or U9186 (N_9186,N_8225,N_8269);
xor U9187 (N_9187,N_8127,N_8102);
and U9188 (N_9188,N_8078,N_8785);
and U9189 (N_9189,N_8333,N_8642);
xnor U9190 (N_9190,N_8499,N_8543);
or U9191 (N_9191,N_8637,N_8597);
xor U9192 (N_9192,N_8124,N_8752);
or U9193 (N_9193,N_8754,N_8228);
and U9194 (N_9194,N_8352,N_8721);
nand U9195 (N_9195,N_8104,N_8507);
xnor U9196 (N_9196,N_8378,N_8964);
or U9197 (N_9197,N_8565,N_8709);
nand U9198 (N_9198,N_8848,N_8076);
nand U9199 (N_9199,N_8453,N_8862);
xor U9200 (N_9200,N_8663,N_8255);
or U9201 (N_9201,N_8773,N_8032);
xor U9202 (N_9202,N_8755,N_8588);
xnor U9203 (N_9203,N_8670,N_8390);
and U9204 (N_9204,N_8298,N_8896);
and U9205 (N_9205,N_8281,N_8023);
nand U9206 (N_9206,N_8855,N_8606);
nand U9207 (N_9207,N_8092,N_8641);
or U9208 (N_9208,N_8356,N_8753);
or U9209 (N_9209,N_8106,N_8688);
xor U9210 (N_9210,N_8110,N_8040);
xnor U9211 (N_9211,N_8485,N_8291);
nand U9212 (N_9212,N_8766,N_8518);
or U9213 (N_9213,N_8075,N_8690);
nand U9214 (N_9214,N_8587,N_8892);
nor U9215 (N_9215,N_8757,N_8399);
nor U9216 (N_9216,N_8242,N_8162);
nand U9217 (N_9217,N_8246,N_8133);
xnor U9218 (N_9218,N_8692,N_8528);
or U9219 (N_9219,N_8575,N_8151);
nand U9220 (N_9220,N_8027,N_8977);
nand U9221 (N_9221,N_8988,N_8302);
or U9222 (N_9222,N_8041,N_8968);
nor U9223 (N_9223,N_8047,N_8778);
nand U9224 (N_9224,N_8178,N_8070);
nand U9225 (N_9225,N_8633,N_8449);
nor U9226 (N_9226,N_8765,N_8326);
xor U9227 (N_9227,N_8285,N_8934);
xor U9228 (N_9228,N_8614,N_8020);
and U9229 (N_9229,N_8568,N_8058);
and U9230 (N_9230,N_8920,N_8472);
nor U9231 (N_9231,N_8108,N_8716);
xnor U9232 (N_9232,N_8001,N_8856);
or U9233 (N_9233,N_8404,N_8906);
and U9234 (N_9234,N_8919,N_8599);
nand U9235 (N_9235,N_8955,N_8413);
nand U9236 (N_9236,N_8744,N_8512);
or U9237 (N_9237,N_8959,N_8939);
xnor U9238 (N_9238,N_8552,N_8289);
xor U9239 (N_9239,N_8898,N_8857);
and U9240 (N_9240,N_8337,N_8186);
and U9241 (N_9241,N_8553,N_8463);
and U9242 (N_9242,N_8643,N_8967);
or U9243 (N_9243,N_8135,N_8252);
or U9244 (N_9244,N_8158,N_8120);
xor U9245 (N_9245,N_8131,N_8435);
and U9246 (N_9246,N_8570,N_8415);
nor U9247 (N_9247,N_8649,N_8830);
or U9248 (N_9248,N_8519,N_8405);
or U9249 (N_9249,N_8525,N_8541);
nand U9250 (N_9250,N_8353,N_8873);
or U9251 (N_9251,N_8524,N_8976);
and U9252 (N_9252,N_8019,N_8897);
xnor U9253 (N_9253,N_8718,N_8006);
nand U9254 (N_9254,N_8735,N_8972);
and U9255 (N_9255,N_8334,N_8077);
or U9256 (N_9256,N_8380,N_8189);
and U9257 (N_9257,N_8270,N_8557);
nor U9258 (N_9258,N_8578,N_8985);
and U9259 (N_9259,N_8538,N_8741);
and U9260 (N_9260,N_8895,N_8797);
nand U9261 (N_9261,N_8833,N_8493);
and U9262 (N_9262,N_8715,N_8805);
xor U9263 (N_9263,N_8881,N_8695);
and U9264 (N_9264,N_8946,N_8112);
xor U9265 (N_9265,N_8065,N_8822);
nand U9266 (N_9266,N_8200,N_8155);
and U9267 (N_9267,N_8201,N_8402);
or U9268 (N_9268,N_8476,N_8276);
xor U9269 (N_9269,N_8283,N_8978);
or U9270 (N_9270,N_8529,N_8307);
or U9271 (N_9271,N_8794,N_8945);
xnor U9272 (N_9272,N_8970,N_8465);
xnor U9273 (N_9273,N_8396,N_8751);
and U9274 (N_9274,N_8930,N_8137);
or U9275 (N_9275,N_8726,N_8837);
nand U9276 (N_9276,N_8204,N_8183);
or U9277 (N_9277,N_8636,N_8559);
or U9278 (N_9278,N_8678,N_8312);
nand U9279 (N_9279,N_8282,N_8264);
xor U9280 (N_9280,N_8971,N_8527);
xor U9281 (N_9281,N_8780,N_8253);
or U9282 (N_9282,N_8016,N_8604);
xnor U9283 (N_9283,N_8351,N_8277);
or U9284 (N_9284,N_8248,N_8148);
nor U9285 (N_9285,N_8733,N_8280);
xnor U9286 (N_9286,N_8330,N_8365);
xor U9287 (N_9287,N_8505,N_8876);
nand U9288 (N_9288,N_8788,N_8969);
or U9289 (N_9289,N_8825,N_8444);
and U9290 (N_9290,N_8303,N_8868);
and U9291 (N_9291,N_8341,N_8980);
or U9292 (N_9292,N_8539,N_8853);
nor U9293 (N_9293,N_8284,N_8691);
and U9294 (N_9294,N_8666,N_8207);
nand U9295 (N_9295,N_8886,N_8387);
or U9296 (N_9296,N_8251,N_8795);
nor U9297 (N_9297,N_8650,N_8490);
xor U9298 (N_9298,N_8492,N_8052);
or U9299 (N_9299,N_8925,N_8169);
xor U9300 (N_9300,N_8961,N_8053);
and U9301 (N_9301,N_8730,N_8774);
or U9302 (N_9302,N_8740,N_8391);
nand U9303 (N_9303,N_8452,N_8571);
nand U9304 (N_9304,N_8615,N_8458);
nor U9305 (N_9305,N_8441,N_8464);
nand U9306 (N_9306,N_8854,N_8561);
nor U9307 (N_9307,N_8669,N_8635);
and U9308 (N_9308,N_8841,N_8259);
nor U9309 (N_9309,N_8290,N_8350);
and U9310 (N_9310,N_8904,N_8609);
xor U9311 (N_9311,N_8537,N_8136);
nand U9312 (N_9312,N_8656,N_8502);
xnor U9313 (N_9313,N_8817,N_8813);
and U9314 (N_9314,N_8962,N_8116);
nor U9315 (N_9315,N_8209,N_8584);
xnor U9316 (N_9316,N_8951,N_8318);
and U9317 (N_9317,N_8749,N_8375);
xor U9318 (N_9318,N_8851,N_8932);
and U9319 (N_9319,N_8012,N_8530);
xnor U9320 (N_9320,N_8496,N_8899);
nand U9321 (N_9321,N_8622,N_8613);
nor U9322 (N_9322,N_8779,N_8175);
nor U9323 (N_9323,N_8157,N_8381);
and U9324 (N_9324,N_8804,N_8960);
nand U9325 (N_9325,N_8174,N_8627);
nand U9326 (N_9326,N_8679,N_8154);
or U9327 (N_9327,N_8489,N_8491);
xnor U9328 (N_9328,N_8245,N_8593);
nor U9329 (N_9329,N_8917,N_8789);
nor U9330 (N_9330,N_8436,N_8943);
and U9331 (N_9331,N_8198,N_8938);
nor U9332 (N_9332,N_8266,N_8580);
nand U9333 (N_9333,N_8542,N_8572);
nor U9334 (N_9334,N_8286,N_8702);
nand U9335 (N_9335,N_8098,N_8229);
or U9336 (N_9336,N_8165,N_8438);
xnor U9337 (N_9337,N_8193,N_8787);
and U9338 (N_9338,N_8342,N_8941);
nor U9339 (N_9339,N_8646,N_8218);
nand U9340 (N_9340,N_8456,N_8093);
xor U9341 (N_9341,N_8309,N_8800);
nand U9342 (N_9342,N_8992,N_8956);
nor U9343 (N_9343,N_8192,N_8516);
nand U9344 (N_9344,N_8590,N_8122);
or U9345 (N_9345,N_8494,N_8671);
nor U9346 (N_9346,N_8556,N_8469);
and U9347 (N_9347,N_8912,N_8250);
or U9348 (N_9348,N_8141,N_8498);
nand U9349 (N_9349,N_8324,N_8355);
nand U9350 (N_9350,N_8719,N_8171);
xor U9351 (N_9351,N_8205,N_8145);
xor U9352 (N_9352,N_8620,N_8728);
and U9353 (N_9353,N_8819,N_8105);
nand U9354 (N_9354,N_8989,N_8653);
nand U9355 (N_9355,N_8803,N_8392);
nand U9356 (N_9356,N_8674,N_8729);
or U9357 (N_9357,N_8776,N_8585);
xor U9358 (N_9358,N_8217,N_8887);
xor U9359 (N_9359,N_8706,N_8114);
nand U9360 (N_9360,N_8080,N_8029);
nand U9361 (N_9361,N_8907,N_8563);
nor U9362 (N_9362,N_8747,N_8030);
xor U9363 (N_9363,N_8581,N_8462);
nand U9364 (N_9364,N_8673,N_8340);
or U9365 (N_9365,N_8577,N_8034);
nand U9366 (N_9366,N_8188,N_8095);
nor U9367 (N_9367,N_8180,N_8676);
or U9368 (N_9368,N_8181,N_8654);
and U9369 (N_9369,N_8824,N_8406);
xnor U9370 (N_9370,N_8547,N_8952);
nand U9371 (N_9371,N_8625,N_8987);
or U9372 (N_9372,N_8867,N_8126);
and U9373 (N_9373,N_8997,N_8783);
nor U9374 (N_9374,N_8546,N_8395);
nand U9375 (N_9375,N_8428,N_8055);
nand U9376 (N_9376,N_8836,N_8236);
or U9377 (N_9377,N_8081,N_8981);
nor U9378 (N_9378,N_8059,N_8915);
and U9379 (N_9379,N_8535,N_8768);
nor U9380 (N_9380,N_8033,N_8511);
nor U9381 (N_9381,N_8523,N_8683);
and U9382 (N_9382,N_8322,N_8398);
nor U9383 (N_9383,N_8905,N_8457);
nor U9384 (N_9384,N_8048,N_8928);
nand U9385 (N_9385,N_8416,N_8166);
nor U9386 (N_9386,N_8685,N_8475);
nand U9387 (N_9387,N_8086,N_8940);
nor U9388 (N_9388,N_8903,N_8835);
xor U9389 (N_9389,N_8424,N_8883);
nor U9390 (N_9390,N_8429,N_8600);
nor U9391 (N_9391,N_8947,N_8292);
nand U9392 (N_9392,N_8662,N_8177);
nor U9393 (N_9393,N_8278,N_8164);
nor U9394 (N_9394,N_8446,N_8979);
or U9395 (N_9395,N_8134,N_8313);
xnor U9396 (N_9396,N_8623,N_8521);
and U9397 (N_9397,N_8224,N_8215);
xnor U9398 (N_9398,N_8601,N_8471);
and U9399 (N_9399,N_8015,N_8481);
or U9400 (N_9400,N_8325,N_8482);
or U9401 (N_9401,N_8878,N_8843);
and U9402 (N_9402,N_8373,N_8143);
and U9403 (N_9403,N_8628,N_8360);
nor U9404 (N_9404,N_8826,N_8013);
nand U9405 (N_9405,N_8176,N_8025);
or U9406 (N_9406,N_8684,N_8210);
or U9407 (N_9407,N_8152,N_8573);
xnor U9408 (N_9408,N_8203,N_8758);
or U9409 (N_9409,N_8426,N_8639);
nor U9410 (N_9410,N_8257,N_8388);
or U9411 (N_9411,N_8208,N_8051);
and U9412 (N_9412,N_8560,N_8331);
nand U9413 (N_9413,N_8450,N_8731);
or U9414 (N_9414,N_8983,N_8617);
or U9415 (N_9415,N_8860,N_8007);
xor U9416 (N_9416,N_8764,N_8348);
nor U9417 (N_9417,N_8738,N_8011);
or U9418 (N_9418,N_8272,N_8327);
nand U9419 (N_9419,N_8226,N_8403);
or U9420 (N_9420,N_8359,N_8039);
or U9421 (N_9421,N_8984,N_8335);
or U9422 (N_9422,N_8038,N_8035);
and U9423 (N_9423,N_8659,N_8767);
nor U9424 (N_9424,N_8551,N_8222);
or U9425 (N_9425,N_8890,N_8031);
xor U9426 (N_9426,N_8770,N_8933);
nand U9427 (N_9427,N_8185,N_8488);
nand U9428 (N_9428,N_8664,N_8394);
nand U9429 (N_9429,N_8675,N_8829);
nand U9430 (N_9430,N_8846,N_8060);
nand U9431 (N_9431,N_8227,N_8230);
nand U9432 (N_9432,N_8742,N_8434);
nand U9433 (N_9433,N_8412,N_8384);
nor U9434 (N_9434,N_8986,N_8594);
xor U9435 (N_9435,N_8202,N_8681);
nand U9436 (N_9436,N_8311,N_8950);
or U9437 (N_9437,N_8008,N_8831);
and U9438 (N_9438,N_8305,N_8849);
or U9439 (N_9439,N_8239,N_8591);
nor U9440 (N_9440,N_8004,N_8522);
nor U9441 (N_9441,N_8701,N_8132);
or U9442 (N_9442,N_8913,N_8515);
and U9443 (N_9443,N_8759,N_8275);
nor U9444 (N_9444,N_8363,N_8418);
and U9445 (N_9445,N_8310,N_8958);
or U9446 (N_9446,N_8672,N_8262);
and U9447 (N_9447,N_8364,N_8603);
or U9448 (N_9448,N_8168,N_8708);
and U9449 (N_9449,N_8705,N_8219);
or U9450 (N_9450,N_8863,N_8704);
and U9451 (N_9451,N_8513,N_8809);
xnor U9452 (N_9452,N_8739,N_8847);
and U9453 (N_9453,N_8894,N_8864);
xnor U9454 (N_9454,N_8454,N_8781);
nor U9455 (N_9455,N_8937,N_8419);
nand U9456 (N_9456,N_8727,N_8397);
xnor U9457 (N_9457,N_8273,N_8439);
nor U9458 (N_9458,N_8107,N_8693);
and U9459 (N_9459,N_8743,N_8455);
or U9460 (N_9460,N_8263,N_8017);
nor U9461 (N_9461,N_8417,N_8784);
nor U9462 (N_9462,N_8880,N_8214);
nand U9463 (N_9463,N_8926,N_8760);
xnor U9464 (N_9464,N_8713,N_8576);
nand U9465 (N_9465,N_8320,N_8295);
or U9466 (N_9466,N_8948,N_8425);
and U9467 (N_9467,N_8068,N_8022);
xnor U9468 (N_9468,N_8510,N_8682);
xnor U9469 (N_9469,N_8645,N_8478);
or U9470 (N_9470,N_8056,N_8583);
and U9471 (N_9471,N_8082,N_8233);
nor U9472 (N_9472,N_8409,N_8128);
and U9473 (N_9473,N_8213,N_8889);
or U9474 (N_9474,N_8480,N_8667);
and U9475 (N_9475,N_8621,N_8445);
and U9476 (N_9476,N_8249,N_8343);
nor U9477 (N_9477,N_8520,N_8762);
xnor U9478 (N_9478,N_8816,N_8099);
xnor U9479 (N_9479,N_8432,N_8074);
nand U9480 (N_9480,N_8775,N_8802);
or U9481 (N_9481,N_8949,N_8159);
nand U9482 (N_9482,N_8420,N_8574);
and U9483 (N_9483,N_8723,N_8815);
xnor U9484 (N_9484,N_8440,N_8791);
nand U9485 (N_9485,N_8893,N_8761);
or U9486 (N_9486,N_8746,N_8361);
nor U9487 (N_9487,N_8153,N_8043);
xor U9488 (N_9488,N_8605,N_8973);
xnor U9489 (N_9489,N_8430,N_8631);
and U9490 (N_9490,N_8139,N_8129);
nor U9491 (N_9491,N_8931,N_8696);
xnor U9492 (N_9492,N_8244,N_8003);
nand U9493 (N_9493,N_8596,N_8910);
xor U9494 (N_9494,N_8314,N_8811);
and U9495 (N_9495,N_8196,N_8231);
and U9496 (N_9496,N_8329,N_8808);
nor U9497 (N_9497,N_8234,N_8447);
xnor U9498 (N_9498,N_8991,N_8400);
nor U9499 (N_9499,N_8317,N_8144);
and U9500 (N_9500,N_8620,N_8429);
xnor U9501 (N_9501,N_8069,N_8488);
nor U9502 (N_9502,N_8716,N_8803);
and U9503 (N_9503,N_8921,N_8108);
nor U9504 (N_9504,N_8662,N_8911);
nor U9505 (N_9505,N_8990,N_8639);
or U9506 (N_9506,N_8449,N_8555);
and U9507 (N_9507,N_8853,N_8785);
or U9508 (N_9508,N_8837,N_8783);
nor U9509 (N_9509,N_8581,N_8143);
nor U9510 (N_9510,N_8534,N_8207);
nand U9511 (N_9511,N_8608,N_8054);
nand U9512 (N_9512,N_8544,N_8505);
nor U9513 (N_9513,N_8183,N_8490);
xnor U9514 (N_9514,N_8195,N_8545);
or U9515 (N_9515,N_8291,N_8337);
and U9516 (N_9516,N_8350,N_8448);
xor U9517 (N_9517,N_8205,N_8448);
xnor U9518 (N_9518,N_8368,N_8568);
or U9519 (N_9519,N_8521,N_8395);
xnor U9520 (N_9520,N_8743,N_8876);
nor U9521 (N_9521,N_8880,N_8280);
nor U9522 (N_9522,N_8103,N_8765);
nand U9523 (N_9523,N_8213,N_8443);
or U9524 (N_9524,N_8962,N_8967);
nand U9525 (N_9525,N_8714,N_8319);
xor U9526 (N_9526,N_8164,N_8957);
xnor U9527 (N_9527,N_8155,N_8859);
nor U9528 (N_9528,N_8942,N_8170);
or U9529 (N_9529,N_8956,N_8888);
or U9530 (N_9530,N_8028,N_8231);
and U9531 (N_9531,N_8207,N_8118);
and U9532 (N_9532,N_8943,N_8772);
and U9533 (N_9533,N_8579,N_8856);
nor U9534 (N_9534,N_8544,N_8521);
nor U9535 (N_9535,N_8172,N_8406);
or U9536 (N_9536,N_8467,N_8315);
and U9537 (N_9537,N_8233,N_8543);
and U9538 (N_9538,N_8029,N_8892);
nor U9539 (N_9539,N_8410,N_8175);
or U9540 (N_9540,N_8392,N_8550);
nor U9541 (N_9541,N_8745,N_8913);
nand U9542 (N_9542,N_8282,N_8223);
nor U9543 (N_9543,N_8429,N_8319);
xnor U9544 (N_9544,N_8172,N_8931);
xnor U9545 (N_9545,N_8709,N_8113);
and U9546 (N_9546,N_8854,N_8626);
or U9547 (N_9547,N_8118,N_8396);
nor U9548 (N_9548,N_8396,N_8594);
xor U9549 (N_9549,N_8722,N_8436);
and U9550 (N_9550,N_8681,N_8300);
xnor U9551 (N_9551,N_8707,N_8158);
xor U9552 (N_9552,N_8503,N_8832);
xor U9553 (N_9553,N_8234,N_8618);
xor U9554 (N_9554,N_8155,N_8781);
xor U9555 (N_9555,N_8688,N_8063);
xor U9556 (N_9556,N_8603,N_8784);
xor U9557 (N_9557,N_8089,N_8724);
nor U9558 (N_9558,N_8219,N_8335);
nor U9559 (N_9559,N_8456,N_8323);
and U9560 (N_9560,N_8048,N_8321);
or U9561 (N_9561,N_8529,N_8524);
nor U9562 (N_9562,N_8160,N_8997);
nor U9563 (N_9563,N_8555,N_8473);
and U9564 (N_9564,N_8067,N_8420);
xor U9565 (N_9565,N_8148,N_8197);
nand U9566 (N_9566,N_8201,N_8414);
nor U9567 (N_9567,N_8925,N_8992);
or U9568 (N_9568,N_8692,N_8150);
nand U9569 (N_9569,N_8895,N_8270);
xnor U9570 (N_9570,N_8610,N_8611);
xnor U9571 (N_9571,N_8077,N_8965);
xnor U9572 (N_9572,N_8208,N_8506);
nor U9573 (N_9573,N_8068,N_8295);
nor U9574 (N_9574,N_8545,N_8636);
or U9575 (N_9575,N_8070,N_8816);
or U9576 (N_9576,N_8229,N_8790);
nand U9577 (N_9577,N_8868,N_8256);
and U9578 (N_9578,N_8794,N_8801);
and U9579 (N_9579,N_8825,N_8837);
nor U9580 (N_9580,N_8537,N_8853);
nor U9581 (N_9581,N_8593,N_8486);
xor U9582 (N_9582,N_8689,N_8543);
and U9583 (N_9583,N_8749,N_8160);
xor U9584 (N_9584,N_8418,N_8413);
nor U9585 (N_9585,N_8979,N_8248);
nor U9586 (N_9586,N_8095,N_8839);
xnor U9587 (N_9587,N_8003,N_8112);
or U9588 (N_9588,N_8283,N_8417);
and U9589 (N_9589,N_8926,N_8405);
nor U9590 (N_9590,N_8015,N_8078);
xor U9591 (N_9591,N_8090,N_8068);
or U9592 (N_9592,N_8915,N_8701);
nor U9593 (N_9593,N_8154,N_8093);
and U9594 (N_9594,N_8913,N_8829);
and U9595 (N_9595,N_8267,N_8583);
nand U9596 (N_9596,N_8524,N_8071);
nor U9597 (N_9597,N_8546,N_8756);
xnor U9598 (N_9598,N_8785,N_8101);
nand U9599 (N_9599,N_8091,N_8355);
and U9600 (N_9600,N_8957,N_8626);
and U9601 (N_9601,N_8951,N_8265);
nor U9602 (N_9602,N_8702,N_8694);
nor U9603 (N_9603,N_8135,N_8333);
nand U9604 (N_9604,N_8110,N_8177);
xor U9605 (N_9605,N_8604,N_8993);
or U9606 (N_9606,N_8575,N_8694);
xnor U9607 (N_9607,N_8035,N_8327);
xnor U9608 (N_9608,N_8160,N_8807);
nand U9609 (N_9609,N_8530,N_8853);
nor U9610 (N_9610,N_8781,N_8375);
nor U9611 (N_9611,N_8605,N_8958);
or U9612 (N_9612,N_8461,N_8822);
or U9613 (N_9613,N_8519,N_8332);
xor U9614 (N_9614,N_8301,N_8139);
xnor U9615 (N_9615,N_8085,N_8283);
nand U9616 (N_9616,N_8661,N_8138);
and U9617 (N_9617,N_8106,N_8342);
and U9618 (N_9618,N_8241,N_8193);
xor U9619 (N_9619,N_8257,N_8714);
xnor U9620 (N_9620,N_8099,N_8511);
and U9621 (N_9621,N_8134,N_8123);
or U9622 (N_9622,N_8902,N_8966);
xor U9623 (N_9623,N_8525,N_8538);
xor U9624 (N_9624,N_8511,N_8483);
nand U9625 (N_9625,N_8245,N_8767);
xnor U9626 (N_9626,N_8742,N_8707);
nor U9627 (N_9627,N_8181,N_8500);
xnor U9628 (N_9628,N_8819,N_8340);
nand U9629 (N_9629,N_8523,N_8960);
nand U9630 (N_9630,N_8355,N_8667);
or U9631 (N_9631,N_8198,N_8116);
and U9632 (N_9632,N_8340,N_8142);
xnor U9633 (N_9633,N_8538,N_8226);
nand U9634 (N_9634,N_8852,N_8655);
nor U9635 (N_9635,N_8874,N_8980);
or U9636 (N_9636,N_8488,N_8471);
and U9637 (N_9637,N_8170,N_8872);
xor U9638 (N_9638,N_8977,N_8724);
xor U9639 (N_9639,N_8727,N_8851);
nor U9640 (N_9640,N_8266,N_8632);
or U9641 (N_9641,N_8159,N_8699);
xnor U9642 (N_9642,N_8201,N_8910);
xor U9643 (N_9643,N_8848,N_8251);
or U9644 (N_9644,N_8320,N_8757);
or U9645 (N_9645,N_8735,N_8498);
nor U9646 (N_9646,N_8111,N_8428);
xnor U9647 (N_9647,N_8267,N_8517);
or U9648 (N_9648,N_8632,N_8259);
xor U9649 (N_9649,N_8598,N_8256);
xnor U9650 (N_9650,N_8843,N_8578);
nor U9651 (N_9651,N_8910,N_8366);
and U9652 (N_9652,N_8513,N_8432);
nor U9653 (N_9653,N_8631,N_8763);
and U9654 (N_9654,N_8452,N_8002);
nand U9655 (N_9655,N_8407,N_8287);
or U9656 (N_9656,N_8384,N_8420);
nor U9657 (N_9657,N_8742,N_8523);
nor U9658 (N_9658,N_8588,N_8560);
nand U9659 (N_9659,N_8820,N_8226);
nand U9660 (N_9660,N_8331,N_8376);
and U9661 (N_9661,N_8423,N_8109);
nand U9662 (N_9662,N_8125,N_8882);
nand U9663 (N_9663,N_8288,N_8993);
and U9664 (N_9664,N_8343,N_8502);
or U9665 (N_9665,N_8391,N_8989);
nor U9666 (N_9666,N_8958,N_8850);
and U9667 (N_9667,N_8311,N_8166);
nor U9668 (N_9668,N_8748,N_8264);
xor U9669 (N_9669,N_8572,N_8863);
nor U9670 (N_9670,N_8292,N_8204);
or U9671 (N_9671,N_8210,N_8317);
xor U9672 (N_9672,N_8320,N_8624);
or U9673 (N_9673,N_8095,N_8402);
or U9674 (N_9674,N_8322,N_8482);
or U9675 (N_9675,N_8739,N_8852);
or U9676 (N_9676,N_8826,N_8715);
xor U9677 (N_9677,N_8882,N_8709);
and U9678 (N_9678,N_8079,N_8052);
xnor U9679 (N_9679,N_8696,N_8629);
xor U9680 (N_9680,N_8540,N_8747);
xnor U9681 (N_9681,N_8872,N_8783);
and U9682 (N_9682,N_8344,N_8039);
or U9683 (N_9683,N_8273,N_8097);
xor U9684 (N_9684,N_8780,N_8863);
or U9685 (N_9685,N_8848,N_8017);
nor U9686 (N_9686,N_8460,N_8303);
xor U9687 (N_9687,N_8169,N_8536);
and U9688 (N_9688,N_8118,N_8883);
xnor U9689 (N_9689,N_8780,N_8911);
or U9690 (N_9690,N_8208,N_8264);
xnor U9691 (N_9691,N_8953,N_8556);
xor U9692 (N_9692,N_8913,N_8932);
and U9693 (N_9693,N_8272,N_8586);
xor U9694 (N_9694,N_8443,N_8661);
nor U9695 (N_9695,N_8644,N_8926);
or U9696 (N_9696,N_8565,N_8303);
nand U9697 (N_9697,N_8609,N_8887);
and U9698 (N_9698,N_8628,N_8604);
xnor U9699 (N_9699,N_8569,N_8444);
or U9700 (N_9700,N_8685,N_8775);
nor U9701 (N_9701,N_8942,N_8098);
or U9702 (N_9702,N_8821,N_8222);
nor U9703 (N_9703,N_8962,N_8707);
or U9704 (N_9704,N_8638,N_8555);
nor U9705 (N_9705,N_8861,N_8699);
or U9706 (N_9706,N_8612,N_8209);
xor U9707 (N_9707,N_8292,N_8162);
and U9708 (N_9708,N_8052,N_8851);
and U9709 (N_9709,N_8423,N_8027);
nor U9710 (N_9710,N_8540,N_8551);
nor U9711 (N_9711,N_8388,N_8484);
nand U9712 (N_9712,N_8194,N_8401);
xnor U9713 (N_9713,N_8232,N_8193);
or U9714 (N_9714,N_8838,N_8119);
or U9715 (N_9715,N_8763,N_8302);
nor U9716 (N_9716,N_8273,N_8148);
nand U9717 (N_9717,N_8405,N_8623);
nor U9718 (N_9718,N_8518,N_8432);
nor U9719 (N_9719,N_8215,N_8229);
nor U9720 (N_9720,N_8779,N_8517);
nand U9721 (N_9721,N_8540,N_8157);
nand U9722 (N_9722,N_8369,N_8717);
xor U9723 (N_9723,N_8863,N_8399);
or U9724 (N_9724,N_8458,N_8830);
xnor U9725 (N_9725,N_8781,N_8505);
nor U9726 (N_9726,N_8744,N_8308);
nor U9727 (N_9727,N_8265,N_8899);
or U9728 (N_9728,N_8935,N_8237);
nor U9729 (N_9729,N_8456,N_8277);
nand U9730 (N_9730,N_8971,N_8738);
or U9731 (N_9731,N_8147,N_8863);
nand U9732 (N_9732,N_8503,N_8034);
or U9733 (N_9733,N_8155,N_8502);
or U9734 (N_9734,N_8823,N_8826);
nand U9735 (N_9735,N_8972,N_8673);
and U9736 (N_9736,N_8299,N_8932);
nor U9737 (N_9737,N_8054,N_8921);
or U9738 (N_9738,N_8771,N_8323);
xor U9739 (N_9739,N_8077,N_8865);
xor U9740 (N_9740,N_8474,N_8539);
or U9741 (N_9741,N_8758,N_8732);
and U9742 (N_9742,N_8605,N_8212);
and U9743 (N_9743,N_8213,N_8278);
or U9744 (N_9744,N_8856,N_8026);
xor U9745 (N_9745,N_8965,N_8015);
xor U9746 (N_9746,N_8229,N_8721);
or U9747 (N_9747,N_8472,N_8891);
nand U9748 (N_9748,N_8584,N_8743);
nand U9749 (N_9749,N_8816,N_8194);
nor U9750 (N_9750,N_8137,N_8197);
nor U9751 (N_9751,N_8427,N_8690);
xnor U9752 (N_9752,N_8493,N_8363);
nor U9753 (N_9753,N_8561,N_8006);
nand U9754 (N_9754,N_8571,N_8472);
nand U9755 (N_9755,N_8740,N_8767);
nand U9756 (N_9756,N_8816,N_8962);
xor U9757 (N_9757,N_8627,N_8124);
and U9758 (N_9758,N_8098,N_8676);
nor U9759 (N_9759,N_8594,N_8250);
xnor U9760 (N_9760,N_8249,N_8410);
nand U9761 (N_9761,N_8144,N_8517);
nand U9762 (N_9762,N_8789,N_8334);
nand U9763 (N_9763,N_8934,N_8532);
xnor U9764 (N_9764,N_8525,N_8615);
xor U9765 (N_9765,N_8044,N_8648);
and U9766 (N_9766,N_8383,N_8397);
nor U9767 (N_9767,N_8818,N_8097);
nor U9768 (N_9768,N_8056,N_8376);
nand U9769 (N_9769,N_8804,N_8241);
nor U9770 (N_9770,N_8933,N_8717);
or U9771 (N_9771,N_8853,N_8771);
and U9772 (N_9772,N_8110,N_8291);
xor U9773 (N_9773,N_8729,N_8326);
nand U9774 (N_9774,N_8864,N_8565);
xor U9775 (N_9775,N_8414,N_8268);
and U9776 (N_9776,N_8513,N_8360);
xor U9777 (N_9777,N_8250,N_8941);
xor U9778 (N_9778,N_8206,N_8347);
or U9779 (N_9779,N_8188,N_8144);
or U9780 (N_9780,N_8240,N_8965);
xor U9781 (N_9781,N_8409,N_8088);
and U9782 (N_9782,N_8828,N_8679);
xnor U9783 (N_9783,N_8874,N_8853);
or U9784 (N_9784,N_8563,N_8117);
nor U9785 (N_9785,N_8923,N_8289);
and U9786 (N_9786,N_8405,N_8768);
nor U9787 (N_9787,N_8530,N_8457);
nand U9788 (N_9788,N_8812,N_8430);
and U9789 (N_9789,N_8736,N_8440);
nand U9790 (N_9790,N_8496,N_8343);
and U9791 (N_9791,N_8959,N_8111);
nor U9792 (N_9792,N_8471,N_8503);
xor U9793 (N_9793,N_8677,N_8808);
or U9794 (N_9794,N_8548,N_8990);
xnor U9795 (N_9795,N_8567,N_8990);
and U9796 (N_9796,N_8244,N_8739);
nor U9797 (N_9797,N_8442,N_8827);
and U9798 (N_9798,N_8821,N_8520);
nor U9799 (N_9799,N_8436,N_8274);
xor U9800 (N_9800,N_8699,N_8125);
nor U9801 (N_9801,N_8390,N_8411);
or U9802 (N_9802,N_8586,N_8616);
and U9803 (N_9803,N_8847,N_8355);
and U9804 (N_9804,N_8849,N_8275);
xor U9805 (N_9805,N_8531,N_8548);
nand U9806 (N_9806,N_8553,N_8001);
xor U9807 (N_9807,N_8544,N_8475);
nor U9808 (N_9808,N_8267,N_8229);
or U9809 (N_9809,N_8365,N_8316);
nand U9810 (N_9810,N_8818,N_8003);
nor U9811 (N_9811,N_8606,N_8345);
or U9812 (N_9812,N_8543,N_8521);
nand U9813 (N_9813,N_8077,N_8407);
nor U9814 (N_9814,N_8745,N_8804);
and U9815 (N_9815,N_8500,N_8530);
xor U9816 (N_9816,N_8330,N_8012);
nor U9817 (N_9817,N_8895,N_8824);
or U9818 (N_9818,N_8674,N_8776);
xor U9819 (N_9819,N_8973,N_8961);
xnor U9820 (N_9820,N_8630,N_8762);
nand U9821 (N_9821,N_8345,N_8389);
nor U9822 (N_9822,N_8955,N_8219);
or U9823 (N_9823,N_8319,N_8332);
xor U9824 (N_9824,N_8621,N_8737);
or U9825 (N_9825,N_8848,N_8084);
and U9826 (N_9826,N_8714,N_8769);
nand U9827 (N_9827,N_8577,N_8552);
or U9828 (N_9828,N_8337,N_8239);
and U9829 (N_9829,N_8477,N_8611);
or U9830 (N_9830,N_8424,N_8081);
or U9831 (N_9831,N_8434,N_8250);
or U9832 (N_9832,N_8272,N_8243);
or U9833 (N_9833,N_8038,N_8994);
xnor U9834 (N_9834,N_8956,N_8679);
and U9835 (N_9835,N_8562,N_8681);
xnor U9836 (N_9836,N_8626,N_8922);
nor U9837 (N_9837,N_8086,N_8911);
and U9838 (N_9838,N_8075,N_8795);
and U9839 (N_9839,N_8285,N_8676);
or U9840 (N_9840,N_8577,N_8602);
or U9841 (N_9841,N_8514,N_8760);
and U9842 (N_9842,N_8590,N_8803);
xnor U9843 (N_9843,N_8230,N_8337);
xor U9844 (N_9844,N_8529,N_8362);
nor U9845 (N_9845,N_8019,N_8275);
nor U9846 (N_9846,N_8572,N_8650);
nor U9847 (N_9847,N_8172,N_8886);
xnor U9848 (N_9848,N_8855,N_8721);
and U9849 (N_9849,N_8332,N_8003);
nand U9850 (N_9850,N_8970,N_8836);
or U9851 (N_9851,N_8323,N_8766);
or U9852 (N_9852,N_8180,N_8782);
or U9853 (N_9853,N_8620,N_8628);
nor U9854 (N_9854,N_8823,N_8003);
and U9855 (N_9855,N_8822,N_8577);
xnor U9856 (N_9856,N_8346,N_8921);
nor U9857 (N_9857,N_8805,N_8993);
xor U9858 (N_9858,N_8331,N_8519);
nand U9859 (N_9859,N_8066,N_8681);
nor U9860 (N_9860,N_8377,N_8542);
nor U9861 (N_9861,N_8660,N_8402);
and U9862 (N_9862,N_8454,N_8678);
and U9863 (N_9863,N_8323,N_8194);
xnor U9864 (N_9864,N_8929,N_8410);
or U9865 (N_9865,N_8167,N_8780);
or U9866 (N_9866,N_8707,N_8399);
and U9867 (N_9867,N_8472,N_8290);
nand U9868 (N_9868,N_8817,N_8404);
nand U9869 (N_9869,N_8663,N_8661);
xor U9870 (N_9870,N_8637,N_8548);
nor U9871 (N_9871,N_8639,N_8276);
or U9872 (N_9872,N_8716,N_8356);
xnor U9873 (N_9873,N_8318,N_8641);
nand U9874 (N_9874,N_8755,N_8150);
nand U9875 (N_9875,N_8605,N_8755);
nand U9876 (N_9876,N_8006,N_8984);
xnor U9877 (N_9877,N_8785,N_8800);
nand U9878 (N_9878,N_8328,N_8643);
nand U9879 (N_9879,N_8815,N_8735);
xor U9880 (N_9880,N_8483,N_8512);
or U9881 (N_9881,N_8244,N_8885);
and U9882 (N_9882,N_8622,N_8456);
nor U9883 (N_9883,N_8586,N_8910);
or U9884 (N_9884,N_8630,N_8208);
or U9885 (N_9885,N_8172,N_8254);
and U9886 (N_9886,N_8146,N_8398);
nor U9887 (N_9887,N_8164,N_8868);
nand U9888 (N_9888,N_8956,N_8624);
nand U9889 (N_9889,N_8525,N_8146);
and U9890 (N_9890,N_8932,N_8248);
xnor U9891 (N_9891,N_8867,N_8292);
or U9892 (N_9892,N_8644,N_8075);
nand U9893 (N_9893,N_8540,N_8097);
or U9894 (N_9894,N_8584,N_8961);
or U9895 (N_9895,N_8956,N_8874);
nor U9896 (N_9896,N_8246,N_8587);
xnor U9897 (N_9897,N_8404,N_8637);
nor U9898 (N_9898,N_8978,N_8834);
and U9899 (N_9899,N_8642,N_8787);
and U9900 (N_9900,N_8216,N_8596);
nor U9901 (N_9901,N_8894,N_8911);
nand U9902 (N_9902,N_8107,N_8773);
or U9903 (N_9903,N_8206,N_8063);
xnor U9904 (N_9904,N_8905,N_8910);
nor U9905 (N_9905,N_8439,N_8777);
nand U9906 (N_9906,N_8044,N_8884);
nor U9907 (N_9907,N_8054,N_8417);
nand U9908 (N_9908,N_8040,N_8176);
and U9909 (N_9909,N_8458,N_8834);
xnor U9910 (N_9910,N_8284,N_8485);
nor U9911 (N_9911,N_8288,N_8279);
xor U9912 (N_9912,N_8230,N_8447);
nand U9913 (N_9913,N_8134,N_8936);
and U9914 (N_9914,N_8828,N_8822);
xnor U9915 (N_9915,N_8088,N_8547);
xor U9916 (N_9916,N_8902,N_8338);
or U9917 (N_9917,N_8094,N_8387);
nand U9918 (N_9918,N_8043,N_8045);
nand U9919 (N_9919,N_8304,N_8302);
nor U9920 (N_9920,N_8855,N_8799);
and U9921 (N_9921,N_8814,N_8101);
nor U9922 (N_9922,N_8793,N_8075);
nand U9923 (N_9923,N_8183,N_8215);
nand U9924 (N_9924,N_8460,N_8515);
nand U9925 (N_9925,N_8028,N_8085);
or U9926 (N_9926,N_8452,N_8614);
xor U9927 (N_9927,N_8819,N_8740);
or U9928 (N_9928,N_8641,N_8662);
xnor U9929 (N_9929,N_8842,N_8441);
nor U9930 (N_9930,N_8172,N_8724);
nand U9931 (N_9931,N_8999,N_8209);
or U9932 (N_9932,N_8512,N_8634);
xor U9933 (N_9933,N_8302,N_8215);
or U9934 (N_9934,N_8282,N_8556);
nor U9935 (N_9935,N_8374,N_8792);
or U9936 (N_9936,N_8859,N_8328);
nand U9937 (N_9937,N_8045,N_8265);
nor U9938 (N_9938,N_8266,N_8802);
and U9939 (N_9939,N_8130,N_8734);
or U9940 (N_9940,N_8542,N_8395);
or U9941 (N_9941,N_8682,N_8616);
nor U9942 (N_9942,N_8390,N_8140);
or U9943 (N_9943,N_8976,N_8720);
or U9944 (N_9944,N_8439,N_8859);
xor U9945 (N_9945,N_8800,N_8043);
or U9946 (N_9946,N_8370,N_8691);
and U9947 (N_9947,N_8951,N_8670);
xor U9948 (N_9948,N_8100,N_8252);
xnor U9949 (N_9949,N_8869,N_8987);
nand U9950 (N_9950,N_8554,N_8571);
xnor U9951 (N_9951,N_8915,N_8375);
and U9952 (N_9952,N_8401,N_8245);
nand U9953 (N_9953,N_8682,N_8707);
nand U9954 (N_9954,N_8277,N_8066);
nand U9955 (N_9955,N_8336,N_8398);
nor U9956 (N_9956,N_8367,N_8648);
or U9957 (N_9957,N_8371,N_8830);
nand U9958 (N_9958,N_8302,N_8407);
nor U9959 (N_9959,N_8959,N_8299);
nand U9960 (N_9960,N_8304,N_8020);
and U9961 (N_9961,N_8652,N_8153);
or U9962 (N_9962,N_8838,N_8002);
xor U9963 (N_9963,N_8823,N_8845);
and U9964 (N_9964,N_8728,N_8749);
nand U9965 (N_9965,N_8989,N_8445);
nor U9966 (N_9966,N_8671,N_8448);
and U9967 (N_9967,N_8290,N_8323);
and U9968 (N_9968,N_8976,N_8612);
and U9969 (N_9969,N_8329,N_8807);
nand U9970 (N_9970,N_8689,N_8490);
xnor U9971 (N_9971,N_8765,N_8873);
and U9972 (N_9972,N_8063,N_8062);
xor U9973 (N_9973,N_8485,N_8558);
or U9974 (N_9974,N_8517,N_8696);
nor U9975 (N_9975,N_8056,N_8668);
nand U9976 (N_9976,N_8703,N_8439);
nand U9977 (N_9977,N_8027,N_8805);
or U9978 (N_9978,N_8408,N_8635);
nand U9979 (N_9979,N_8749,N_8640);
or U9980 (N_9980,N_8240,N_8422);
nor U9981 (N_9981,N_8923,N_8907);
nand U9982 (N_9982,N_8788,N_8448);
and U9983 (N_9983,N_8685,N_8695);
or U9984 (N_9984,N_8746,N_8438);
xnor U9985 (N_9985,N_8090,N_8275);
and U9986 (N_9986,N_8057,N_8254);
or U9987 (N_9987,N_8194,N_8730);
xnor U9988 (N_9988,N_8818,N_8175);
nand U9989 (N_9989,N_8685,N_8894);
nor U9990 (N_9990,N_8529,N_8406);
or U9991 (N_9991,N_8101,N_8374);
or U9992 (N_9992,N_8298,N_8963);
or U9993 (N_9993,N_8860,N_8295);
or U9994 (N_9994,N_8032,N_8858);
nor U9995 (N_9995,N_8843,N_8541);
or U9996 (N_9996,N_8767,N_8372);
xor U9997 (N_9997,N_8439,N_8279);
nor U9998 (N_9998,N_8742,N_8509);
xor U9999 (N_9999,N_8454,N_8787);
nand UO_0 (O_0,N_9671,N_9602);
and UO_1 (O_1,N_9272,N_9415);
or UO_2 (O_2,N_9144,N_9243);
or UO_3 (O_3,N_9895,N_9716);
and UO_4 (O_4,N_9531,N_9119);
and UO_5 (O_5,N_9141,N_9528);
nand UO_6 (O_6,N_9041,N_9870);
or UO_7 (O_7,N_9394,N_9814);
or UO_8 (O_8,N_9817,N_9952);
nand UO_9 (O_9,N_9588,N_9223);
nand UO_10 (O_10,N_9884,N_9309);
nand UO_11 (O_11,N_9927,N_9562);
and UO_12 (O_12,N_9084,N_9063);
and UO_13 (O_13,N_9167,N_9400);
nand UO_14 (O_14,N_9023,N_9827);
or UO_15 (O_15,N_9964,N_9821);
nand UO_16 (O_16,N_9247,N_9692);
and UO_17 (O_17,N_9168,N_9442);
xnor UO_18 (O_18,N_9347,N_9199);
and UO_19 (O_19,N_9398,N_9926);
and UO_20 (O_20,N_9031,N_9914);
nand UO_21 (O_21,N_9738,N_9457);
and UO_22 (O_22,N_9380,N_9685);
nand UO_23 (O_23,N_9291,N_9941);
nor UO_24 (O_24,N_9687,N_9592);
xor UO_25 (O_25,N_9440,N_9581);
nor UO_26 (O_26,N_9973,N_9064);
or UO_27 (O_27,N_9226,N_9274);
nor UO_28 (O_28,N_9128,N_9633);
or UO_29 (O_29,N_9570,N_9049);
nor UO_30 (O_30,N_9536,N_9495);
nor UO_31 (O_31,N_9136,N_9338);
nor UO_32 (O_32,N_9950,N_9391);
and UO_33 (O_33,N_9478,N_9789);
nand UO_34 (O_34,N_9346,N_9868);
and UO_35 (O_35,N_9138,N_9542);
and UO_36 (O_36,N_9148,N_9636);
and UO_37 (O_37,N_9578,N_9635);
nand UO_38 (O_38,N_9087,N_9651);
or UO_39 (O_39,N_9967,N_9285);
or UO_40 (O_40,N_9159,N_9170);
xor UO_41 (O_41,N_9307,N_9587);
nand UO_42 (O_42,N_9426,N_9677);
or UO_43 (O_43,N_9175,N_9683);
xnor UO_44 (O_44,N_9509,N_9147);
nor UO_45 (O_45,N_9874,N_9378);
xnor UO_46 (O_46,N_9767,N_9854);
and UO_47 (O_47,N_9310,N_9918);
nor UO_48 (O_48,N_9251,N_9920);
xnor UO_49 (O_49,N_9813,N_9277);
or UO_50 (O_50,N_9344,N_9999);
and UO_51 (O_51,N_9704,N_9404);
or UO_52 (O_52,N_9376,N_9011);
xnor UO_53 (O_53,N_9909,N_9235);
or UO_54 (O_54,N_9244,N_9334);
or UO_55 (O_55,N_9688,N_9682);
and UO_56 (O_56,N_9286,N_9406);
and UO_57 (O_57,N_9858,N_9872);
nand UO_58 (O_58,N_9497,N_9327);
nand UO_59 (O_59,N_9493,N_9900);
nor UO_60 (O_60,N_9254,N_9490);
nand UO_61 (O_61,N_9844,N_9585);
or UO_62 (O_62,N_9358,N_9712);
and UO_63 (O_63,N_9473,N_9553);
nor UO_64 (O_64,N_9545,N_9289);
or UO_65 (O_65,N_9997,N_9150);
nor UO_66 (O_66,N_9943,N_9444);
xor UO_67 (O_67,N_9968,N_9607);
nor UO_68 (O_68,N_9778,N_9705);
nand UO_69 (O_69,N_9043,N_9919);
or UO_70 (O_70,N_9666,N_9451);
or UO_71 (O_71,N_9122,N_9510);
xnor UO_72 (O_72,N_9019,N_9463);
or UO_73 (O_73,N_9220,N_9686);
or UO_74 (O_74,N_9186,N_9988);
nand UO_75 (O_75,N_9187,N_9593);
nand UO_76 (O_76,N_9349,N_9328);
or UO_77 (O_77,N_9676,N_9776);
nand UO_78 (O_78,N_9402,N_9539);
and UO_79 (O_79,N_9202,N_9977);
nand UO_80 (O_80,N_9308,N_9629);
or UO_81 (O_81,N_9046,N_9631);
nor UO_82 (O_82,N_9236,N_9832);
nor UO_83 (O_83,N_9230,N_9184);
nor UO_84 (O_84,N_9355,N_9998);
or UO_85 (O_85,N_9760,N_9969);
xor UO_86 (O_86,N_9921,N_9595);
xnor UO_87 (O_87,N_9154,N_9924);
nor UO_88 (O_88,N_9555,N_9322);
xnor UO_89 (O_89,N_9375,N_9461);
nor UO_90 (O_90,N_9743,N_9548);
and UO_91 (O_91,N_9320,N_9978);
or UO_92 (O_92,N_9204,N_9248);
nand UO_93 (O_93,N_9030,N_9020);
and UO_94 (O_94,N_9362,N_9381);
nand UO_95 (O_95,N_9646,N_9925);
nor UO_96 (O_96,N_9241,N_9456);
nand UO_97 (O_97,N_9042,N_9881);
nor UO_98 (O_98,N_9282,N_9123);
or UO_99 (O_99,N_9034,N_9260);
and UO_100 (O_100,N_9650,N_9661);
and UO_101 (O_101,N_9865,N_9133);
nor UO_102 (O_102,N_9949,N_9418);
nor UO_103 (O_103,N_9145,N_9219);
nor UO_104 (O_104,N_9169,N_9519);
nor UO_105 (O_105,N_9829,N_9281);
xor UO_106 (O_106,N_9546,N_9574);
or UO_107 (O_107,N_9229,N_9601);
nand UO_108 (O_108,N_9113,N_9847);
nand UO_109 (O_109,N_9499,N_9526);
or UO_110 (O_110,N_9200,N_9234);
nor UO_111 (O_111,N_9431,N_9037);
or UO_112 (O_112,N_9935,N_9240);
nand UO_113 (O_113,N_9742,N_9162);
nor UO_114 (O_114,N_9665,N_9916);
nor UO_115 (O_115,N_9675,N_9565);
nor UO_116 (O_116,N_9799,N_9547);
nand UO_117 (O_117,N_9283,N_9433);
xor UO_118 (O_118,N_9749,N_9024);
or UO_119 (O_119,N_9855,N_9589);
xor UO_120 (O_120,N_9785,N_9937);
nand UO_121 (O_121,N_9560,N_9667);
nor UO_122 (O_122,N_9314,N_9656);
xnor UO_123 (O_123,N_9231,N_9901);
xor UO_124 (O_124,N_9954,N_9970);
nor UO_125 (O_125,N_9753,N_9852);
and UO_126 (O_126,N_9411,N_9794);
nand UO_127 (O_127,N_9225,N_9896);
nand UO_128 (O_128,N_9691,N_9641);
nand UO_129 (O_129,N_9085,N_9820);
or UO_130 (O_130,N_9538,N_9904);
or UO_131 (O_131,N_9905,N_9730);
xor UO_132 (O_132,N_9191,N_9965);
and UO_133 (O_133,N_9628,N_9211);
nand UO_134 (O_134,N_9318,N_9718);
or UO_135 (O_135,N_9193,N_9010);
nor UO_136 (O_136,N_9093,N_9487);
nand UO_137 (O_137,N_9535,N_9080);
nand UO_138 (O_138,N_9563,N_9157);
or UO_139 (O_139,N_9216,N_9597);
nand UO_140 (O_140,N_9819,N_9525);
and UO_141 (O_141,N_9354,N_9891);
nand UO_142 (O_142,N_9069,N_9898);
xor UO_143 (O_143,N_9364,N_9611);
nand UO_144 (O_144,N_9953,N_9757);
and UO_145 (O_145,N_9811,N_9383);
nor UO_146 (O_146,N_9714,N_9130);
xor UO_147 (O_147,N_9771,N_9003);
nand UO_148 (O_148,N_9680,N_9025);
and UO_149 (O_149,N_9933,N_9207);
and UO_150 (O_150,N_9072,N_9805);
nand UO_151 (O_151,N_9479,N_9609);
nand UO_152 (O_152,N_9335,N_9996);
nand UO_153 (O_153,N_9894,N_9419);
nor UO_154 (O_154,N_9496,N_9494);
or UO_155 (O_155,N_9971,N_9002);
or UO_156 (O_156,N_9125,N_9224);
nand UO_157 (O_157,N_9985,N_9527);
or UO_158 (O_158,N_9534,N_9054);
nand UO_159 (O_159,N_9252,N_9784);
nand UO_160 (O_160,N_9139,N_9561);
nor UO_161 (O_161,N_9625,N_9302);
xor UO_162 (O_162,N_9627,N_9506);
and UO_163 (O_163,N_9336,N_9114);
or UO_164 (O_164,N_9903,N_9246);
and UO_165 (O_165,N_9082,N_9387);
nand UO_166 (O_166,N_9780,N_9893);
and UO_167 (O_167,N_9339,N_9039);
or UO_168 (O_168,N_9174,N_9569);
and UO_169 (O_169,N_9779,N_9867);
or UO_170 (O_170,N_9746,N_9837);
and UO_171 (O_171,N_9810,N_9151);
xor UO_172 (O_172,N_9099,N_9710);
nand UO_173 (O_173,N_9348,N_9057);
and UO_174 (O_174,N_9679,N_9214);
nor UO_175 (O_175,N_9115,N_9700);
nand UO_176 (O_176,N_9443,N_9511);
nand UO_177 (O_177,N_9363,N_9135);
nand UO_178 (O_178,N_9986,N_9566);
nand UO_179 (O_179,N_9763,N_9630);
xor UO_180 (O_180,N_9075,N_9834);
and UO_181 (O_181,N_9153,N_9212);
nor UO_182 (O_182,N_9374,N_9594);
or UO_183 (O_183,N_9180,N_9963);
and UO_184 (O_184,N_9556,N_9198);
nand UO_185 (O_185,N_9098,N_9612);
nand UO_186 (O_186,N_9040,N_9100);
xor UO_187 (O_187,N_9915,N_9222);
nor UO_188 (O_188,N_9856,N_9001);
xnor UO_189 (O_189,N_9412,N_9196);
and UO_190 (O_190,N_9709,N_9257);
nor UO_191 (O_191,N_9055,N_9341);
nand UO_192 (O_192,N_9360,N_9873);
and UO_193 (O_193,N_9853,N_9544);
xor UO_194 (O_194,N_9637,N_9849);
nand UO_195 (O_195,N_9579,N_9410);
or UO_196 (O_196,N_9770,N_9864);
or UO_197 (O_197,N_9836,N_9568);
or UO_198 (O_198,N_9504,N_9689);
or UO_199 (O_199,N_9584,N_9599);
xnor UO_200 (O_200,N_9861,N_9713);
and UO_201 (O_201,N_9888,N_9270);
nand UO_202 (O_202,N_9724,N_9524);
xnor UO_203 (O_203,N_9660,N_9397);
and UO_204 (O_204,N_9467,N_9598);
xor UO_205 (O_205,N_9365,N_9802);
and UO_206 (O_206,N_9294,N_9902);
or UO_207 (O_207,N_9695,N_9179);
or UO_208 (O_208,N_9824,N_9181);
or UO_209 (O_209,N_9908,N_9500);
nand UO_210 (O_210,N_9727,N_9720);
nor UO_211 (O_211,N_9726,N_9583);
and UO_212 (O_212,N_9751,N_9481);
xor UO_213 (O_213,N_9729,N_9137);
and UO_214 (O_214,N_9006,N_9731);
nand UO_215 (O_215,N_9027,N_9863);
or UO_216 (O_216,N_9803,N_9543);
nand UO_217 (O_217,N_9475,N_9317);
nor UO_218 (O_218,N_9879,N_9129);
xnor UO_219 (O_219,N_9319,N_9477);
nor UO_220 (O_220,N_9089,N_9045);
or UO_221 (O_221,N_9796,N_9717);
or UO_222 (O_222,N_9668,N_9203);
or UO_223 (O_223,N_9871,N_9155);
and UO_224 (O_224,N_9752,N_9541);
xor UO_225 (O_225,N_9897,N_9409);
xnor UO_226 (O_226,N_9848,N_9697);
and UO_227 (O_227,N_9103,N_9576);
and UO_228 (O_228,N_9250,N_9368);
and UO_229 (O_229,N_9945,N_9210);
and UO_230 (O_230,N_9065,N_9851);
xor UO_231 (O_231,N_9036,N_9177);
or UO_232 (O_232,N_9498,N_9617);
nand UO_233 (O_233,N_9206,N_9425);
or UO_234 (O_234,N_9333,N_9590);
nand UO_235 (O_235,N_9761,N_9176);
xnor UO_236 (O_236,N_9640,N_9357);
nand UO_237 (O_237,N_9452,N_9422);
xor UO_238 (O_238,N_9552,N_9102);
nand UO_239 (O_239,N_9423,N_9468);
or UO_240 (O_240,N_9816,N_9373);
or UO_241 (O_241,N_9066,N_9058);
or UO_242 (O_242,N_9392,N_9060);
xnor UO_243 (O_243,N_9809,N_9619);
nor UO_244 (O_244,N_9306,N_9804);
nand UO_245 (O_245,N_9690,N_9134);
or UO_246 (O_246,N_9118,N_9981);
xor UO_247 (O_247,N_9068,N_9446);
or UO_248 (O_248,N_9350,N_9684);
and UO_249 (O_249,N_9655,N_9911);
and UO_250 (O_250,N_9735,N_9429);
nor UO_251 (O_251,N_9140,N_9416);
xnor UO_252 (O_252,N_9649,N_9812);
and UO_253 (O_253,N_9994,N_9258);
nor UO_254 (O_254,N_9958,N_9448);
xor UO_255 (O_255,N_9715,N_9875);
nand UO_256 (O_256,N_9377,N_9790);
nand UO_257 (O_257,N_9737,N_9614);
nor UO_258 (O_258,N_9866,N_9604);
or UO_259 (O_259,N_9267,N_9886);
and UO_260 (O_260,N_9626,N_9501);
xnor UO_261 (O_261,N_9882,N_9505);
nand UO_262 (O_262,N_9488,N_9559);
nor UO_263 (O_263,N_9741,N_9944);
xor UO_264 (O_264,N_9182,N_9765);
nor UO_265 (O_265,N_9116,N_9736);
xor UO_266 (O_266,N_9917,N_9417);
xnor UO_267 (O_267,N_9472,N_9342);
xor UO_268 (O_268,N_9421,N_9728);
or UO_269 (O_269,N_9664,N_9722);
and UO_270 (O_270,N_9303,N_9474);
nand UO_271 (O_271,N_9750,N_9414);
or UO_272 (O_272,N_9259,N_9793);
or UO_273 (O_273,N_9470,N_9669);
and UO_274 (O_274,N_9255,N_9610);
nor UO_275 (O_275,N_9095,N_9907);
nor UO_276 (O_276,N_9194,N_9486);
nand UO_277 (O_277,N_9842,N_9242);
xnor UO_278 (O_278,N_9432,N_9185);
nor UO_279 (O_279,N_9201,N_9015);
or UO_280 (O_280,N_9466,N_9449);
xor UO_281 (O_281,N_9465,N_9663);
and UO_282 (O_282,N_9645,N_9554);
xor UO_283 (O_283,N_9990,N_9239);
xor UO_284 (O_284,N_9022,N_9183);
xor UO_285 (O_285,N_9939,N_9846);
or UO_286 (O_286,N_9883,N_9476);
nor UO_287 (O_287,N_9922,N_9507);
xor UO_288 (O_288,N_9517,N_9453);
or UO_289 (O_289,N_9192,N_9615);
xor UO_290 (O_290,N_9980,N_9104);
xnor UO_291 (O_291,N_9221,N_9390);
nor UO_292 (O_292,N_9766,N_9838);
nor UO_293 (O_293,N_9026,N_9081);
nand UO_294 (O_294,N_9420,N_9021);
nand UO_295 (O_295,N_9616,N_9938);
xnor UO_296 (O_296,N_9483,N_9056);
or UO_297 (O_297,N_9271,N_9067);
and UO_298 (O_298,N_9826,N_9957);
or UO_299 (O_299,N_9698,N_9263);
or UO_300 (O_300,N_9862,N_9092);
xor UO_301 (O_301,N_9156,N_9121);
nor UO_302 (O_302,N_9946,N_9047);
nand UO_303 (O_303,N_9877,N_9295);
or UO_304 (O_304,N_9781,N_9108);
or UO_305 (O_305,N_9618,N_9127);
and UO_306 (O_306,N_9083,N_9132);
nand UO_307 (O_307,N_9723,N_9029);
or UO_308 (O_308,N_9438,N_9332);
nand UO_309 (O_309,N_9936,N_9343);
nor UO_310 (O_310,N_9979,N_9190);
nand UO_311 (O_311,N_9351,N_9312);
nor UO_312 (O_312,N_9460,N_9052);
nand UO_313 (O_313,N_9575,N_9105);
and UO_314 (O_314,N_9995,N_9454);
xor UO_315 (O_315,N_9783,N_9632);
xor UO_316 (O_316,N_9831,N_9050);
and UO_317 (O_317,N_9644,N_9384);
and UO_318 (O_318,N_9993,N_9401);
or UO_319 (O_319,N_9480,N_9004);
nor UO_320 (O_320,N_9513,N_9197);
nor UO_321 (O_321,N_9120,N_9984);
xnor UO_322 (O_322,N_9428,N_9253);
and UO_323 (O_323,N_9131,N_9016);
or UO_324 (O_324,N_9489,N_9928);
nor UO_325 (O_325,N_9828,N_9966);
nor UO_326 (O_326,N_9395,N_9035);
xor UO_327 (O_327,N_9323,N_9773);
xnor UO_328 (O_328,N_9218,N_9393);
xnor UO_329 (O_329,N_9279,N_9117);
or UO_330 (O_330,N_9931,N_9366);
nor UO_331 (O_331,N_9078,N_9951);
or UO_332 (O_332,N_9972,N_9857);
and UO_333 (O_333,N_9424,N_9955);
nand UO_334 (O_334,N_9975,N_9352);
and UO_335 (O_335,N_9007,N_9711);
nand UO_336 (O_336,N_9839,N_9642);
nor UO_337 (O_337,N_9795,N_9379);
nand UO_338 (O_338,N_9324,N_9573);
or UO_339 (O_339,N_9305,N_9013);
nand UO_340 (O_340,N_9292,N_9297);
nor UO_341 (O_341,N_9106,N_9876);
xor UO_342 (O_342,N_9076,N_9755);
and UO_343 (O_343,N_9090,N_9734);
nand UO_344 (O_344,N_9189,N_9808);
and UO_345 (O_345,N_9540,N_9699);
nor UO_346 (O_346,N_9208,N_9906);
and UO_347 (O_347,N_9899,N_9516);
or UO_348 (O_348,N_9772,N_9840);
xor UO_349 (O_349,N_9005,N_9503);
xnor UO_350 (O_350,N_9437,N_9992);
and UO_351 (O_351,N_9396,N_9747);
nor UO_352 (O_352,N_9732,N_9329);
nor UO_353 (O_353,N_9471,N_9659);
or UO_354 (O_354,N_9149,N_9678);
nand UO_355 (O_355,N_9800,N_9096);
xnor UO_356 (O_356,N_9791,N_9797);
or UO_357 (O_357,N_9051,N_9608);
xor UO_358 (O_358,N_9386,N_9708);
or UO_359 (O_359,N_9833,N_9215);
or UO_360 (O_360,N_9529,N_9721);
nor UO_361 (O_361,N_9643,N_9245);
xor UO_362 (O_362,N_9662,N_9681);
or UO_363 (O_363,N_9316,N_9389);
and UO_364 (O_364,N_9786,N_9033);
nor UO_365 (O_365,N_9124,N_9754);
nor UO_366 (O_366,N_9464,N_9408);
nor UO_367 (O_367,N_9088,N_9603);
or UO_368 (O_368,N_9775,N_9976);
nor UO_369 (O_369,N_9172,N_9549);
and UO_370 (O_370,N_9508,N_9077);
or UO_371 (O_371,N_9275,N_9340);
nand UO_372 (O_372,N_9702,N_9450);
and UO_373 (O_373,N_9537,N_9654);
nand UO_374 (O_374,N_9053,N_9158);
xor UO_375 (O_375,N_9522,N_9337);
or UO_376 (O_376,N_9606,N_9445);
nand UO_377 (O_377,N_9094,N_9325);
nand UO_378 (O_378,N_9195,N_9237);
xnor UO_379 (O_379,N_9515,N_9798);
or UO_380 (O_380,N_9719,N_9097);
and UO_381 (O_381,N_9012,N_9359);
nand UO_382 (O_382,N_9205,N_9758);
xor UO_383 (O_383,N_9913,N_9371);
and UO_384 (O_384,N_9407,N_9841);
xnor UO_385 (O_385,N_9382,N_9605);
or UO_386 (O_386,N_9345,N_9107);
and UO_387 (O_387,N_9441,N_9948);
xor UO_388 (O_388,N_9620,N_9652);
nand UO_389 (O_389,N_9768,N_9582);
nor UO_390 (O_390,N_9962,N_9326);
or UO_391 (O_391,N_9032,N_9694);
nor UO_392 (O_392,N_9188,N_9178);
or UO_393 (O_393,N_9956,N_9238);
or UO_394 (O_394,N_9523,N_9311);
nand UO_395 (O_395,N_9028,N_9693);
xnor UO_396 (O_396,N_9764,N_9923);
xor UO_397 (O_397,N_9672,N_9586);
and UO_398 (O_398,N_9430,N_9835);
and UO_399 (O_399,N_9017,N_9367);
or UO_400 (O_400,N_9290,N_9745);
nand UO_401 (O_401,N_9878,N_9934);
nand UO_402 (O_402,N_9280,N_9447);
and UO_403 (O_403,N_9073,N_9171);
nand UO_404 (O_404,N_9707,N_9091);
nor UO_405 (O_405,N_9596,N_9142);
or UO_406 (O_406,N_9788,N_9213);
xnor UO_407 (O_407,N_9166,N_9653);
xnor UO_408 (O_408,N_9300,N_9845);
xor UO_409 (O_409,N_9982,N_9930);
or UO_410 (O_410,N_9143,N_9111);
or UO_411 (O_411,N_9462,N_9613);
nand UO_412 (O_412,N_9885,N_9502);
or UO_413 (O_413,N_9759,N_9571);
nor UO_414 (O_414,N_9388,N_9491);
nor UO_415 (O_415,N_9657,N_9321);
and UO_416 (O_416,N_9278,N_9774);
xor UO_417 (O_417,N_9580,N_9815);
nor UO_418 (O_418,N_9869,N_9146);
xnor UO_419 (O_419,N_9126,N_9860);
and UO_420 (O_420,N_9304,N_9009);
or UO_421 (O_421,N_9109,N_9014);
nand UO_422 (O_422,N_9634,N_9287);
or UO_423 (O_423,N_9674,N_9288);
or UO_424 (O_424,N_9520,N_9947);
nor UO_425 (O_425,N_9806,N_9859);
and UO_426 (O_426,N_9370,N_9173);
nor UO_427 (O_427,N_9638,N_9960);
or UO_428 (O_428,N_9777,N_9353);
nand UO_429 (O_429,N_9455,N_9807);
xnor UO_430 (O_430,N_9706,N_9313);
nand UO_431 (O_431,N_9284,N_9163);
or UO_432 (O_432,N_9086,N_9880);
nand UO_433 (O_433,N_9696,N_9910);
or UO_434 (O_434,N_9492,N_9762);
nand UO_435 (O_435,N_9264,N_9434);
nor UO_436 (O_436,N_9110,N_9298);
or UO_437 (O_437,N_9929,N_9639);
nand UO_438 (O_438,N_9273,N_9801);
and UO_439 (O_439,N_9739,N_9818);
nand UO_440 (O_440,N_9331,N_9112);
or UO_441 (O_441,N_9427,N_9725);
nand UO_442 (O_442,N_9413,N_9769);
or UO_443 (O_443,N_9070,N_9621);
xnor UO_444 (O_444,N_9482,N_9059);
nor UO_445 (O_445,N_9228,N_9782);
and UO_446 (O_446,N_9161,N_9061);
nand UO_447 (O_447,N_9701,N_9458);
xnor UO_448 (O_448,N_9044,N_9843);
xor UO_449 (O_449,N_9436,N_9227);
and UO_450 (O_450,N_9940,N_9887);
nand UO_451 (O_451,N_9330,N_9521);
or UO_452 (O_452,N_9624,N_9484);
nand UO_453 (O_453,N_9648,N_9296);
or UO_454 (O_454,N_9459,N_9792);
and UO_455 (O_455,N_9101,N_9038);
nand UO_456 (O_456,N_9822,N_9748);
and UO_457 (O_457,N_9823,N_9372);
nor UO_458 (O_458,N_9164,N_9160);
or UO_459 (O_459,N_9018,N_9600);
nand UO_460 (O_460,N_9293,N_9233);
or UO_461 (O_461,N_9567,N_9399);
nand UO_462 (O_462,N_9892,N_9825);
xor UO_463 (O_463,N_9830,N_9262);
xor UO_464 (O_464,N_9991,N_9673);
xor UO_465 (O_465,N_9550,N_9266);
xor UO_466 (O_466,N_9744,N_9989);
xor UO_467 (O_467,N_9959,N_9572);
nand UO_468 (O_468,N_9369,N_9932);
and UO_469 (O_469,N_9961,N_9008);
xnor UO_470 (O_470,N_9385,N_9558);
and UO_471 (O_471,N_9532,N_9756);
and UO_472 (O_472,N_9512,N_9623);
and UO_473 (O_473,N_9974,N_9533);
xnor UO_474 (O_474,N_9850,N_9889);
or UO_475 (O_475,N_9485,N_9530);
xnor UO_476 (O_476,N_9276,N_9079);
xnor UO_477 (O_477,N_9439,N_9256);
nand UO_478 (O_478,N_9265,N_9658);
xor UO_479 (O_479,N_9405,N_9000);
xor UO_480 (O_480,N_9518,N_9622);
xnor UO_481 (O_481,N_9435,N_9890);
nand UO_482 (O_482,N_9469,N_9048);
nand UO_483 (O_483,N_9165,N_9209);
and UO_484 (O_484,N_9577,N_9062);
nand UO_485 (O_485,N_9912,N_9403);
or UO_486 (O_486,N_9315,N_9361);
or UO_487 (O_487,N_9356,N_9299);
xor UO_488 (O_488,N_9301,N_9564);
and UO_489 (O_489,N_9268,N_9557);
or UO_490 (O_490,N_9942,N_9787);
and UO_491 (O_491,N_9670,N_9152);
nor UO_492 (O_492,N_9733,N_9249);
nor UO_493 (O_493,N_9647,N_9217);
nor UO_494 (O_494,N_9987,N_9740);
nor UO_495 (O_495,N_9269,N_9591);
nor UO_496 (O_496,N_9983,N_9514);
nor UO_497 (O_497,N_9703,N_9261);
or UO_498 (O_498,N_9074,N_9071);
and UO_499 (O_499,N_9551,N_9232);
nor UO_500 (O_500,N_9025,N_9435);
xnor UO_501 (O_501,N_9057,N_9826);
or UO_502 (O_502,N_9143,N_9478);
or UO_503 (O_503,N_9874,N_9107);
nand UO_504 (O_504,N_9462,N_9285);
and UO_505 (O_505,N_9669,N_9868);
or UO_506 (O_506,N_9064,N_9756);
xnor UO_507 (O_507,N_9989,N_9943);
and UO_508 (O_508,N_9757,N_9072);
xnor UO_509 (O_509,N_9944,N_9615);
xnor UO_510 (O_510,N_9051,N_9537);
xor UO_511 (O_511,N_9049,N_9566);
xor UO_512 (O_512,N_9111,N_9783);
nor UO_513 (O_513,N_9191,N_9019);
xor UO_514 (O_514,N_9635,N_9355);
and UO_515 (O_515,N_9994,N_9927);
nand UO_516 (O_516,N_9573,N_9370);
xnor UO_517 (O_517,N_9377,N_9572);
and UO_518 (O_518,N_9430,N_9770);
xnor UO_519 (O_519,N_9709,N_9154);
nor UO_520 (O_520,N_9651,N_9603);
xor UO_521 (O_521,N_9491,N_9608);
nor UO_522 (O_522,N_9865,N_9205);
nor UO_523 (O_523,N_9493,N_9039);
xor UO_524 (O_524,N_9049,N_9158);
xnor UO_525 (O_525,N_9479,N_9407);
nand UO_526 (O_526,N_9092,N_9909);
xor UO_527 (O_527,N_9549,N_9658);
nand UO_528 (O_528,N_9238,N_9174);
xor UO_529 (O_529,N_9836,N_9292);
nor UO_530 (O_530,N_9657,N_9207);
xor UO_531 (O_531,N_9457,N_9723);
nor UO_532 (O_532,N_9790,N_9903);
nor UO_533 (O_533,N_9949,N_9313);
nand UO_534 (O_534,N_9554,N_9872);
xnor UO_535 (O_535,N_9918,N_9408);
or UO_536 (O_536,N_9475,N_9959);
or UO_537 (O_537,N_9037,N_9724);
nand UO_538 (O_538,N_9169,N_9758);
and UO_539 (O_539,N_9192,N_9349);
and UO_540 (O_540,N_9038,N_9263);
nand UO_541 (O_541,N_9311,N_9353);
nand UO_542 (O_542,N_9324,N_9256);
and UO_543 (O_543,N_9359,N_9639);
and UO_544 (O_544,N_9374,N_9405);
or UO_545 (O_545,N_9714,N_9848);
nor UO_546 (O_546,N_9656,N_9153);
or UO_547 (O_547,N_9154,N_9963);
nor UO_548 (O_548,N_9515,N_9227);
and UO_549 (O_549,N_9247,N_9213);
nor UO_550 (O_550,N_9994,N_9975);
or UO_551 (O_551,N_9398,N_9567);
nand UO_552 (O_552,N_9681,N_9521);
xnor UO_553 (O_553,N_9009,N_9398);
xor UO_554 (O_554,N_9407,N_9513);
nand UO_555 (O_555,N_9180,N_9841);
nor UO_556 (O_556,N_9454,N_9268);
nor UO_557 (O_557,N_9757,N_9566);
nor UO_558 (O_558,N_9401,N_9794);
and UO_559 (O_559,N_9553,N_9917);
and UO_560 (O_560,N_9712,N_9822);
xor UO_561 (O_561,N_9621,N_9883);
or UO_562 (O_562,N_9658,N_9885);
xor UO_563 (O_563,N_9810,N_9800);
nand UO_564 (O_564,N_9687,N_9398);
or UO_565 (O_565,N_9836,N_9657);
or UO_566 (O_566,N_9957,N_9806);
or UO_567 (O_567,N_9077,N_9175);
nand UO_568 (O_568,N_9290,N_9278);
or UO_569 (O_569,N_9083,N_9733);
nor UO_570 (O_570,N_9146,N_9052);
nor UO_571 (O_571,N_9818,N_9381);
nand UO_572 (O_572,N_9718,N_9030);
nor UO_573 (O_573,N_9700,N_9087);
or UO_574 (O_574,N_9210,N_9655);
and UO_575 (O_575,N_9190,N_9464);
nand UO_576 (O_576,N_9725,N_9115);
and UO_577 (O_577,N_9626,N_9929);
nor UO_578 (O_578,N_9772,N_9640);
nand UO_579 (O_579,N_9489,N_9875);
nor UO_580 (O_580,N_9733,N_9595);
nor UO_581 (O_581,N_9512,N_9862);
or UO_582 (O_582,N_9001,N_9339);
or UO_583 (O_583,N_9113,N_9891);
xnor UO_584 (O_584,N_9391,N_9184);
nand UO_585 (O_585,N_9843,N_9674);
or UO_586 (O_586,N_9739,N_9058);
and UO_587 (O_587,N_9316,N_9831);
and UO_588 (O_588,N_9052,N_9377);
nor UO_589 (O_589,N_9668,N_9917);
xnor UO_590 (O_590,N_9510,N_9893);
and UO_591 (O_591,N_9463,N_9200);
nor UO_592 (O_592,N_9549,N_9312);
and UO_593 (O_593,N_9737,N_9032);
nand UO_594 (O_594,N_9738,N_9485);
and UO_595 (O_595,N_9554,N_9707);
xor UO_596 (O_596,N_9748,N_9187);
nor UO_597 (O_597,N_9241,N_9969);
nor UO_598 (O_598,N_9197,N_9799);
xor UO_599 (O_599,N_9141,N_9640);
xnor UO_600 (O_600,N_9999,N_9220);
nand UO_601 (O_601,N_9355,N_9066);
nand UO_602 (O_602,N_9419,N_9389);
xnor UO_603 (O_603,N_9367,N_9268);
nand UO_604 (O_604,N_9225,N_9649);
or UO_605 (O_605,N_9219,N_9856);
nand UO_606 (O_606,N_9137,N_9895);
nor UO_607 (O_607,N_9487,N_9625);
or UO_608 (O_608,N_9013,N_9256);
nand UO_609 (O_609,N_9008,N_9950);
nor UO_610 (O_610,N_9506,N_9326);
nand UO_611 (O_611,N_9423,N_9070);
xor UO_612 (O_612,N_9027,N_9590);
nand UO_613 (O_613,N_9438,N_9156);
xor UO_614 (O_614,N_9360,N_9818);
xor UO_615 (O_615,N_9322,N_9049);
nand UO_616 (O_616,N_9255,N_9308);
nand UO_617 (O_617,N_9600,N_9418);
nor UO_618 (O_618,N_9641,N_9237);
nor UO_619 (O_619,N_9848,N_9358);
nand UO_620 (O_620,N_9940,N_9793);
nand UO_621 (O_621,N_9808,N_9456);
and UO_622 (O_622,N_9753,N_9361);
and UO_623 (O_623,N_9022,N_9790);
and UO_624 (O_624,N_9695,N_9841);
nand UO_625 (O_625,N_9607,N_9760);
nand UO_626 (O_626,N_9583,N_9047);
or UO_627 (O_627,N_9259,N_9968);
or UO_628 (O_628,N_9009,N_9242);
and UO_629 (O_629,N_9616,N_9039);
and UO_630 (O_630,N_9540,N_9281);
xnor UO_631 (O_631,N_9115,N_9429);
or UO_632 (O_632,N_9828,N_9154);
nor UO_633 (O_633,N_9168,N_9543);
or UO_634 (O_634,N_9760,N_9965);
xor UO_635 (O_635,N_9964,N_9086);
nor UO_636 (O_636,N_9634,N_9024);
nor UO_637 (O_637,N_9549,N_9061);
xnor UO_638 (O_638,N_9105,N_9607);
and UO_639 (O_639,N_9592,N_9737);
or UO_640 (O_640,N_9866,N_9326);
xor UO_641 (O_641,N_9668,N_9026);
or UO_642 (O_642,N_9140,N_9810);
or UO_643 (O_643,N_9176,N_9738);
or UO_644 (O_644,N_9555,N_9991);
xnor UO_645 (O_645,N_9141,N_9597);
or UO_646 (O_646,N_9506,N_9125);
nand UO_647 (O_647,N_9664,N_9549);
nor UO_648 (O_648,N_9978,N_9003);
xnor UO_649 (O_649,N_9179,N_9998);
nor UO_650 (O_650,N_9104,N_9893);
and UO_651 (O_651,N_9581,N_9386);
or UO_652 (O_652,N_9023,N_9338);
or UO_653 (O_653,N_9066,N_9785);
or UO_654 (O_654,N_9848,N_9520);
or UO_655 (O_655,N_9879,N_9313);
or UO_656 (O_656,N_9676,N_9665);
xnor UO_657 (O_657,N_9910,N_9721);
xor UO_658 (O_658,N_9914,N_9849);
xor UO_659 (O_659,N_9868,N_9055);
and UO_660 (O_660,N_9401,N_9636);
and UO_661 (O_661,N_9526,N_9318);
nand UO_662 (O_662,N_9163,N_9950);
nand UO_663 (O_663,N_9671,N_9273);
nor UO_664 (O_664,N_9734,N_9315);
or UO_665 (O_665,N_9151,N_9318);
xor UO_666 (O_666,N_9848,N_9855);
nand UO_667 (O_667,N_9964,N_9874);
or UO_668 (O_668,N_9547,N_9488);
nor UO_669 (O_669,N_9954,N_9526);
and UO_670 (O_670,N_9397,N_9137);
nor UO_671 (O_671,N_9885,N_9856);
or UO_672 (O_672,N_9958,N_9639);
and UO_673 (O_673,N_9629,N_9619);
nor UO_674 (O_674,N_9074,N_9918);
nor UO_675 (O_675,N_9060,N_9004);
nand UO_676 (O_676,N_9166,N_9847);
nand UO_677 (O_677,N_9384,N_9169);
nand UO_678 (O_678,N_9299,N_9148);
xnor UO_679 (O_679,N_9651,N_9974);
or UO_680 (O_680,N_9585,N_9517);
or UO_681 (O_681,N_9694,N_9468);
nor UO_682 (O_682,N_9120,N_9297);
nor UO_683 (O_683,N_9734,N_9718);
or UO_684 (O_684,N_9064,N_9819);
nor UO_685 (O_685,N_9520,N_9648);
and UO_686 (O_686,N_9542,N_9076);
nor UO_687 (O_687,N_9395,N_9495);
xor UO_688 (O_688,N_9229,N_9789);
nand UO_689 (O_689,N_9501,N_9700);
or UO_690 (O_690,N_9122,N_9457);
nor UO_691 (O_691,N_9194,N_9507);
or UO_692 (O_692,N_9810,N_9294);
nand UO_693 (O_693,N_9955,N_9877);
or UO_694 (O_694,N_9888,N_9922);
and UO_695 (O_695,N_9123,N_9860);
or UO_696 (O_696,N_9591,N_9333);
or UO_697 (O_697,N_9328,N_9653);
nand UO_698 (O_698,N_9534,N_9375);
or UO_699 (O_699,N_9275,N_9667);
nand UO_700 (O_700,N_9408,N_9878);
nor UO_701 (O_701,N_9781,N_9237);
nand UO_702 (O_702,N_9177,N_9303);
nor UO_703 (O_703,N_9861,N_9386);
nand UO_704 (O_704,N_9756,N_9856);
nor UO_705 (O_705,N_9507,N_9422);
nand UO_706 (O_706,N_9106,N_9648);
or UO_707 (O_707,N_9603,N_9849);
nor UO_708 (O_708,N_9565,N_9186);
nor UO_709 (O_709,N_9784,N_9489);
nor UO_710 (O_710,N_9663,N_9761);
and UO_711 (O_711,N_9259,N_9476);
or UO_712 (O_712,N_9837,N_9433);
or UO_713 (O_713,N_9278,N_9306);
and UO_714 (O_714,N_9820,N_9679);
xnor UO_715 (O_715,N_9644,N_9413);
or UO_716 (O_716,N_9023,N_9556);
nand UO_717 (O_717,N_9794,N_9063);
xnor UO_718 (O_718,N_9847,N_9954);
nand UO_719 (O_719,N_9077,N_9577);
xnor UO_720 (O_720,N_9548,N_9155);
or UO_721 (O_721,N_9078,N_9929);
nor UO_722 (O_722,N_9180,N_9552);
and UO_723 (O_723,N_9443,N_9227);
xnor UO_724 (O_724,N_9714,N_9340);
or UO_725 (O_725,N_9273,N_9234);
nor UO_726 (O_726,N_9223,N_9543);
or UO_727 (O_727,N_9399,N_9504);
xnor UO_728 (O_728,N_9656,N_9908);
nand UO_729 (O_729,N_9978,N_9218);
nor UO_730 (O_730,N_9886,N_9412);
or UO_731 (O_731,N_9189,N_9702);
xnor UO_732 (O_732,N_9616,N_9802);
nor UO_733 (O_733,N_9495,N_9203);
and UO_734 (O_734,N_9205,N_9791);
and UO_735 (O_735,N_9881,N_9754);
and UO_736 (O_736,N_9458,N_9371);
nand UO_737 (O_737,N_9749,N_9211);
nor UO_738 (O_738,N_9723,N_9028);
or UO_739 (O_739,N_9552,N_9982);
and UO_740 (O_740,N_9222,N_9560);
or UO_741 (O_741,N_9555,N_9318);
and UO_742 (O_742,N_9674,N_9722);
and UO_743 (O_743,N_9485,N_9512);
or UO_744 (O_744,N_9084,N_9952);
or UO_745 (O_745,N_9567,N_9823);
xor UO_746 (O_746,N_9587,N_9014);
nor UO_747 (O_747,N_9108,N_9956);
or UO_748 (O_748,N_9212,N_9032);
nor UO_749 (O_749,N_9630,N_9170);
xor UO_750 (O_750,N_9924,N_9961);
and UO_751 (O_751,N_9542,N_9994);
or UO_752 (O_752,N_9190,N_9347);
nor UO_753 (O_753,N_9413,N_9605);
nor UO_754 (O_754,N_9254,N_9759);
xnor UO_755 (O_755,N_9925,N_9444);
nand UO_756 (O_756,N_9243,N_9276);
and UO_757 (O_757,N_9335,N_9298);
and UO_758 (O_758,N_9033,N_9417);
nand UO_759 (O_759,N_9821,N_9956);
xor UO_760 (O_760,N_9327,N_9351);
and UO_761 (O_761,N_9949,N_9877);
or UO_762 (O_762,N_9535,N_9149);
nand UO_763 (O_763,N_9394,N_9014);
nand UO_764 (O_764,N_9316,N_9242);
or UO_765 (O_765,N_9622,N_9564);
nor UO_766 (O_766,N_9679,N_9551);
nor UO_767 (O_767,N_9624,N_9518);
nand UO_768 (O_768,N_9143,N_9435);
nand UO_769 (O_769,N_9396,N_9124);
xnor UO_770 (O_770,N_9186,N_9378);
nor UO_771 (O_771,N_9236,N_9048);
or UO_772 (O_772,N_9216,N_9810);
and UO_773 (O_773,N_9411,N_9134);
xor UO_774 (O_774,N_9251,N_9760);
or UO_775 (O_775,N_9422,N_9894);
and UO_776 (O_776,N_9339,N_9765);
or UO_777 (O_777,N_9594,N_9274);
nor UO_778 (O_778,N_9603,N_9497);
and UO_779 (O_779,N_9580,N_9578);
nand UO_780 (O_780,N_9526,N_9919);
nor UO_781 (O_781,N_9461,N_9011);
and UO_782 (O_782,N_9856,N_9775);
nor UO_783 (O_783,N_9822,N_9910);
nor UO_784 (O_784,N_9705,N_9977);
nor UO_785 (O_785,N_9412,N_9948);
nor UO_786 (O_786,N_9377,N_9205);
nand UO_787 (O_787,N_9848,N_9837);
nor UO_788 (O_788,N_9973,N_9405);
nand UO_789 (O_789,N_9896,N_9411);
or UO_790 (O_790,N_9596,N_9634);
or UO_791 (O_791,N_9992,N_9091);
nor UO_792 (O_792,N_9085,N_9339);
nor UO_793 (O_793,N_9806,N_9043);
nor UO_794 (O_794,N_9875,N_9618);
and UO_795 (O_795,N_9344,N_9349);
nor UO_796 (O_796,N_9870,N_9181);
xnor UO_797 (O_797,N_9208,N_9458);
nand UO_798 (O_798,N_9160,N_9678);
nand UO_799 (O_799,N_9685,N_9556);
and UO_800 (O_800,N_9170,N_9995);
nor UO_801 (O_801,N_9611,N_9535);
nor UO_802 (O_802,N_9873,N_9971);
nor UO_803 (O_803,N_9766,N_9933);
nor UO_804 (O_804,N_9400,N_9611);
and UO_805 (O_805,N_9216,N_9545);
and UO_806 (O_806,N_9757,N_9767);
nor UO_807 (O_807,N_9985,N_9194);
and UO_808 (O_808,N_9535,N_9956);
and UO_809 (O_809,N_9844,N_9058);
nand UO_810 (O_810,N_9119,N_9677);
and UO_811 (O_811,N_9232,N_9955);
nand UO_812 (O_812,N_9643,N_9192);
xor UO_813 (O_813,N_9097,N_9805);
nand UO_814 (O_814,N_9532,N_9533);
or UO_815 (O_815,N_9573,N_9623);
nor UO_816 (O_816,N_9474,N_9716);
or UO_817 (O_817,N_9684,N_9682);
nor UO_818 (O_818,N_9904,N_9309);
nor UO_819 (O_819,N_9916,N_9378);
nand UO_820 (O_820,N_9411,N_9639);
xor UO_821 (O_821,N_9652,N_9344);
nand UO_822 (O_822,N_9908,N_9974);
xor UO_823 (O_823,N_9543,N_9070);
nand UO_824 (O_824,N_9304,N_9189);
xor UO_825 (O_825,N_9593,N_9074);
nor UO_826 (O_826,N_9303,N_9904);
nand UO_827 (O_827,N_9515,N_9029);
and UO_828 (O_828,N_9691,N_9567);
nor UO_829 (O_829,N_9554,N_9184);
xor UO_830 (O_830,N_9844,N_9613);
nand UO_831 (O_831,N_9668,N_9357);
nand UO_832 (O_832,N_9109,N_9913);
nor UO_833 (O_833,N_9054,N_9145);
nor UO_834 (O_834,N_9432,N_9007);
nor UO_835 (O_835,N_9659,N_9356);
nor UO_836 (O_836,N_9954,N_9360);
and UO_837 (O_837,N_9971,N_9275);
or UO_838 (O_838,N_9776,N_9043);
nor UO_839 (O_839,N_9014,N_9875);
nor UO_840 (O_840,N_9222,N_9260);
xor UO_841 (O_841,N_9607,N_9835);
nand UO_842 (O_842,N_9458,N_9856);
nand UO_843 (O_843,N_9675,N_9648);
nor UO_844 (O_844,N_9613,N_9700);
or UO_845 (O_845,N_9090,N_9695);
and UO_846 (O_846,N_9171,N_9749);
nor UO_847 (O_847,N_9492,N_9494);
nand UO_848 (O_848,N_9874,N_9495);
or UO_849 (O_849,N_9515,N_9278);
or UO_850 (O_850,N_9397,N_9554);
nand UO_851 (O_851,N_9406,N_9175);
nor UO_852 (O_852,N_9572,N_9631);
nand UO_853 (O_853,N_9118,N_9754);
or UO_854 (O_854,N_9446,N_9940);
and UO_855 (O_855,N_9772,N_9698);
nand UO_856 (O_856,N_9287,N_9631);
nand UO_857 (O_857,N_9272,N_9243);
nand UO_858 (O_858,N_9997,N_9828);
nand UO_859 (O_859,N_9473,N_9795);
or UO_860 (O_860,N_9986,N_9878);
nor UO_861 (O_861,N_9970,N_9187);
or UO_862 (O_862,N_9867,N_9143);
nor UO_863 (O_863,N_9238,N_9938);
nor UO_864 (O_864,N_9154,N_9350);
nor UO_865 (O_865,N_9786,N_9366);
xnor UO_866 (O_866,N_9556,N_9961);
xnor UO_867 (O_867,N_9508,N_9018);
nor UO_868 (O_868,N_9297,N_9643);
nor UO_869 (O_869,N_9331,N_9214);
nor UO_870 (O_870,N_9942,N_9355);
xor UO_871 (O_871,N_9798,N_9503);
nand UO_872 (O_872,N_9248,N_9279);
xor UO_873 (O_873,N_9349,N_9179);
xnor UO_874 (O_874,N_9014,N_9538);
and UO_875 (O_875,N_9289,N_9772);
and UO_876 (O_876,N_9004,N_9141);
nand UO_877 (O_877,N_9849,N_9832);
nor UO_878 (O_878,N_9773,N_9873);
or UO_879 (O_879,N_9832,N_9926);
and UO_880 (O_880,N_9886,N_9827);
and UO_881 (O_881,N_9530,N_9310);
nand UO_882 (O_882,N_9654,N_9028);
nand UO_883 (O_883,N_9042,N_9197);
nor UO_884 (O_884,N_9613,N_9198);
xnor UO_885 (O_885,N_9290,N_9907);
xnor UO_886 (O_886,N_9507,N_9505);
and UO_887 (O_887,N_9518,N_9672);
xor UO_888 (O_888,N_9680,N_9625);
or UO_889 (O_889,N_9529,N_9664);
nand UO_890 (O_890,N_9103,N_9752);
xor UO_891 (O_891,N_9860,N_9561);
xnor UO_892 (O_892,N_9212,N_9196);
and UO_893 (O_893,N_9571,N_9667);
nor UO_894 (O_894,N_9186,N_9455);
and UO_895 (O_895,N_9709,N_9406);
or UO_896 (O_896,N_9269,N_9368);
and UO_897 (O_897,N_9937,N_9587);
or UO_898 (O_898,N_9288,N_9824);
nor UO_899 (O_899,N_9025,N_9695);
and UO_900 (O_900,N_9221,N_9462);
nor UO_901 (O_901,N_9730,N_9789);
and UO_902 (O_902,N_9542,N_9636);
and UO_903 (O_903,N_9985,N_9091);
or UO_904 (O_904,N_9723,N_9138);
and UO_905 (O_905,N_9786,N_9852);
or UO_906 (O_906,N_9109,N_9127);
nand UO_907 (O_907,N_9214,N_9091);
nor UO_908 (O_908,N_9662,N_9620);
nand UO_909 (O_909,N_9120,N_9784);
xnor UO_910 (O_910,N_9000,N_9517);
nor UO_911 (O_911,N_9898,N_9974);
and UO_912 (O_912,N_9767,N_9770);
or UO_913 (O_913,N_9900,N_9301);
and UO_914 (O_914,N_9708,N_9158);
xnor UO_915 (O_915,N_9760,N_9401);
nand UO_916 (O_916,N_9794,N_9832);
or UO_917 (O_917,N_9497,N_9904);
nor UO_918 (O_918,N_9542,N_9823);
and UO_919 (O_919,N_9354,N_9262);
xor UO_920 (O_920,N_9647,N_9410);
xnor UO_921 (O_921,N_9285,N_9686);
xor UO_922 (O_922,N_9863,N_9417);
xnor UO_923 (O_923,N_9437,N_9330);
xor UO_924 (O_924,N_9055,N_9298);
nor UO_925 (O_925,N_9938,N_9428);
xor UO_926 (O_926,N_9811,N_9232);
nor UO_927 (O_927,N_9995,N_9196);
nor UO_928 (O_928,N_9961,N_9329);
or UO_929 (O_929,N_9563,N_9932);
or UO_930 (O_930,N_9748,N_9475);
or UO_931 (O_931,N_9830,N_9826);
nand UO_932 (O_932,N_9605,N_9652);
or UO_933 (O_933,N_9192,N_9411);
and UO_934 (O_934,N_9535,N_9230);
and UO_935 (O_935,N_9012,N_9226);
nor UO_936 (O_936,N_9626,N_9619);
nor UO_937 (O_937,N_9784,N_9088);
nand UO_938 (O_938,N_9718,N_9540);
and UO_939 (O_939,N_9080,N_9262);
nor UO_940 (O_940,N_9997,N_9677);
nor UO_941 (O_941,N_9024,N_9037);
xnor UO_942 (O_942,N_9253,N_9631);
xor UO_943 (O_943,N_9720,N_9632);
nand UO_944 (O_944,N_9078,N_9956);
and UO_945 (O_945,N_9217,N_9188);
or UO_946 (O_946,N_9031,N_9521);
xnor UO_947 (O_947,N_9089,N_9792);
and UO_948 (O_948,N_9168,N_9568);
nor UO_949 (O_949,N_9991,N_9307);
nor UO_950 (O_950,N_9941,N_9200);
nand UO_951 (O_951,N_9240,N_9126);
nor UO_952 (O_952,N_9821,N_9333);
xor UO_953 (O_953,N_9017,N_9256);
and UO_954 (O_954,N_9717,N_9105);
nor UO_955 (O_955,N_9585,N_9094);
or UO_956 (O_956,N_9191,N_9883);
or UO_957 (O_957,N_9826,N_9041);
and UO_958 (O_958,N_9602,N_9067);
nand UO_959 (O_959,N_9796,N_9504);
xnor UO_960 (O_960,N_9553,N_9734);
xor UO_961 (O_961,N_9881,N_9065);
and UO_962 (O_962,N_9230,N_9799);
xor UO_963 (O_963,N_9028,N_9228);
nor UO_964 (O_964,N_9983,N_9356);
nand UO_965 (O_965,N_9926,N_9351);
xnor UO_966 (O_966,N_9473,N_9446);
nand UO_967 (O_967,N_9365,N_9113);
or UO_968 (O_968,N_9997,N_9774);
and UO_969 (O_969,N_9277,N_9645);
nor UO_970 (O_970,N_9717,N_9373);
or UO_971 (O_971,N_9349,N_9949);
and UO_972 (O_972,N_9679,N_9381);
and UO_973 (O_973,N_9535,N_9919);
or UO_974 (O_974,N_9102,N_9193);
xnor UO_975 (O_975,N_9340,N_9578);
xor UO_976 (O_976,N_9567,N_9568);
or UO_977 (O_977,N_9318,N_9344);
and UO_978 (O_978,N_9952,N_9531);
and UO_979 (O_979,N_9262,N_9113);
nand UO_980 (O_980,N_9151,N_9918);
nand UO_981 (O_981,N_9321,N_9464);
or UO_982 (O_982,N_9621,N_9010);
and UO_983 (O_983,N_9379,N_9327);
and UO_984 (O_984,N_9199,N_9310);
nand UO_985 (O_985,N_9355,N_9650);
xnor UO_986 (O_986,N_9393,N_9162);
or UO_987 (O_987,N_9826,N_9465);
xnor UO_988 (O_988,N_9062,N_9972);
nand UO_989 (O_989,N_9981,N_9892);
and UO_990 (O_990,N_9910,N_9392);
or UO_991 (O_991,N_9822,N_9171);
or UO_992 (O_992,N_9657,N_9720);
and UO_993 (O_993,N_9308,N_9696);
nor UO_994 (O_994,N_9058,N_9329);
nor UO_995 (O_995,N_9579,N_9414);
nor UO_996 (O_996,N_9695,N_9219);
nor UO_997 (O_997,N_9983,N_9986);
xor UO_998 (O_998,N_9544,N_9005);
or UO_999 (O_999,N_9879,N_9210);
xnor UO_1000 (O_1000,N_9148,N_9904);
and UO_1001 (O_1001,N_9034,N_9532);
xnor UO_1002 (O_1002,N_9509,N_9054);
or UO_1003 (O_1003,N_9545,N_9824);
or UO_1004 (O_1004,N_9475,N_9589);
nand UO_1005 (O_1005,N_9540,N_9935);
and UO_1006 (O_1006,N_9820,N_9273);
or UO_1007 (O_1007,N_9141,N_9551);
nand UO_1008 (O_1008,N_9075,N_9270);
nand UO_1009 (O_1009,N_9489,N_9845);
nand UO_1010 (O_1010,N_9600,N_9614);
or UO_1011 (O_1011,N_9570,N_9999);
or UO_1012 (O_1012,N_9409,N_9427);
nor UO_1013 (O_1013,N_9621,N_9932);
or UO_1014 (O_1014,N_9338,N_9815);
xor UO_1015 (O_1015,N_9514,N_9441);
nand UO_1016 (O_1016,N_9639,N_9887);
and UO_1017 (O_1017,N_9100,N_9470);
or UO_1018 (O_1018,N_9040,N_9235);
and UO_1019 (O_1019,N_9620,N_9012);
and UO_1020 (O_1020,N_9415,N_9509);
xnor UO_1021 (O_1021,N_9531,N_9782);
nand UO_1022 (O_1022,N_9842,N_9313);
xnor UO_1023 (O_1023,N_9091,N_9478);
xnor UO_1024 (O_1024,N_9792,N_9130);
nand UO_1025 (O_1025,N_9895,N_9764);
or UO_1026 (O_1026,N_9303,N_9240);
or UO_1027 (O_1027,N_9507,N_9787);
and UO_1028 (O_1028,N_9787,N_9946);
and UO_1029 (O_1029,N_9575,N_9768);
xnor UO_1030 (O_1030,N_9185,N_9594);
nor UO_1031 (O_1031,N_9527,N_9871);
nor UO_1032 (O_1032,N_9196,N_9088);
xnor UO_1033 (O_1033,N_9067,N_9166);
xnor UO_1034 (O_1034,N_9950,N_9647);
xnor UO_1035 (O_1035,N_9923,N_9672);
nor UO_1036 (O_1036,N_9861,N_9818);
nor UO_1037 (O_1037,N_9329,N_9124);
xor UO_1038 (O_1038,N_9237,N_9741);
or UO_1039 (O_1039,N_9987,N_9517);
xnor UO_1040 (O_1040,N_9690,N_9093);
xor UO_1041 (O_1041,N_9132,N_9215);
or UO_1042 (O_1042,N_9934,N_9862);
nor UO_1043 (O_1043,N_9151,N_9529);
or UO_1044 (O_1044,N_9791,N_9248);
xnor UO_1045 (O_1045,N_9857,N_9258);
and UO_1046 (O_1046,N_9437,N_9723);
nor UO_1047 (O_1047,N_9425,N_9034);
and UO_1048 (O_1048,N_9786,N_9905);
and UO_1049 (O_1049,N_9710,N_9251);
xor UO_1050 (O_1050,N_9814,N_9970);
nor UO_1051 (O_1051,N_9392,N_9111);
or UO_1052 (O_1052,N_9354,N_9467);
xnor UO_1053 (O_1053,N_9090,N_9304);
and UO_1054 (O_1054,N_9774,N_9735);
and UO_1055 (O_1055,N_9656,N_9145);
and UO_1056 (O_1056,N_9945,N_9306);
xnor UO_1057 (O_1057,N_9756,N_9515);
or UO_1058 (O_1058,N_9301,N_9440);
nor UO_1059 (O_1059,N_9528,N_9145);
nor UO_1060 (O_1060,N_9951,N_9492);
xor UO_1061 (O_1061,N_9970,N_9357);
nand UO_1062 (O_1062,N_9302,N_9085);
xor UO_1063 (O_1063,N_9844,N_9598);
xor UO_1064 (O_1064,N_9645,N_9123);
nand UO_1065 (O_1065,N_9013,N_9779);
nand UO_1066 (O_1066,N_9920,N_9254);
or UO_1067 (O_1067,N_9306,N_9617);
and UO_1068 (O_1068,N_9949,N_9906);
xor UO_1069 (O_1069,N_9498,N_9330);
nand UO_1070 (O_1070,N_9649,N_9114);
xnor UO_1071 (O_1071,N_9207,N_9663);
nand UO_1072 (O_1072,N_9317,N_9014);
or UO_1073 (O_1073,N_9431,N_9508);
xor UO_1074 (O_1074,N_9412,N_9272);
and UO_1075 (O_1075,N_9394,N_9090);
nand UO_1076 (O_1076,N_9303,N_9010);
nand UO_1077 (O_1077,N_9621,N_9321);
and UO_1078 (O_1078,N_9201,N_9159);
nand UO_1079 (O_1079,N_9826,N_9636);
nor UO_1080 (O_1080,N_9621,N_9476);
nand UO_1081 (O_1081,N_9993,N_9842);
or UO_1082 (O_1082,N_9812,N_9582);
nor UO_1083 (O_1083,N_9902,N_9871);
and UO_1084 (O_1084,N_9190,N_9918);
and UO_1085 (O_1085,N_9795,N_9429);
or UO_1086 (O_1086,N_9705,N_9308);
or UO_1087 (O_1087,N_9685,N_9533);
nor UO_1088 (O_1088,N_9600,N_9489);
xnor UO_1089 (O_1089,N_9500,N_9255);
xnor UO_1090 (O_1090,N_9437,N_9385);
xor UO_1091 (O_1091,N_9949,N_9419);
nand UO_1092 (O_1092,N_9456,N_9964);
nand UO_1093 (O_1093,N_9112,N_9999);
xnor UO_1094 (O_1094,N_9405,N_9830);
and UO_1095 (O_1095,N_9801,N_9145);
nor UO_1096 (O_1096,N_9237,N_9100);
xnor UO_1097 (O_1097,N_9616,N_9055);
or UO_1098 (O_1098,N_9608,N_9028);
xnor UO_1099 (O_1099,N_9872,N_9617);
xor UO_1100 (O_1100,N_9238,N_9416);
nor UO_1101 (O_1101,N_9310,N_9848);
or UO_1102 (O_1102,N_9076,N_9281);
nand UO_1103 (O_1103,N_9428,N_9209);
nand UO_1104 (O_1104,N_9219,N_9084);
nand UO_1105 (O_1105,N_9276,N_9719);
xor UO_1106 (O_1106,N_9626,N_9711);
nor UO_1107 (O_1107,N_9219,N_9131);
nor UO_1108 (O_1108,N_9892,N_9070);
and UO_1109 (O_1109,N_9635,N_9190);
and UO_1110 (O_1110,N_9819,N_9429);
nor UO_1111 (O_1111,N_9967,N_9503);
or UO_1112 (O_1112,N_9953,N_9433);
nand UO_1113 (O_1113,N_9983,N_9446);
nand UO_1114 (O_1114,N_9314,N_9105);
and UO_1115 (O_1115,N_9765,N_9178);
nor UO_1116 (O_1116,N_9134,N_9427);
nand UO_1117 (O_1117,N_9695,N_9658);
nand UO_1118 (O_1118,N_9592,N_9061);
and UO_1119 (O_1119,N_9098,N_9794);
nand UO_1120 (O_1120,N_9203,N_9518);
nand UO_1121 (O_1121,N_9739,N_9717);
and UO_1122 (O_1122,N_9899,N_9218);
or UO_1123 (O_1123,N_9289,N_9476);
nor UO_1124 (O_1124,N_9435,N_9402);
or UO_1125 (O_1125,N_9368,N_9644);
nor UO_1126 (O_1126,N_9311,N_9154);
nand UO_1127 (O_1127,N_9605,N_9240);
nand UO_1128 (O_1128,N_9768,N_9626);
nor UO_1129 (O_1129,N_9825,N_9633);
and UO_1130 (O_1130,N_9962,N_9989);
xnor UO_1131 (O_1131,N_9696,N_9154);
xor UO_1132 (O_1132,N_9027,N_9749);
nand UO_1133 (O_1133,N_9799,N_9981);
nand UO_1134 (O_1134,N_9891,N_9448);
and UO_1135 (O_1135,N_9244,N_9322);
and UO_1136 (O_1136,N_9510,N_9392);
nand UO_1137 (O_1137,N_9988,N_9823);
and UO_1138 (O_1138,N_9048,N_9731);
or UO_1139 (O_1139,N_9894,N_9348);
nand UO_1140 (O_1140,N_9293,N_9848);
nand UO_1141 (O_1141,N_9790,N_9708);
nand UO_1142 (O_1142,N_9073,N_9619);
nor UO_1143 (O_1143,N_9932,N_9101);
xor UO_1144 (O_1144,N_9095,N_9563);
nand UO_1145 (O_1145,N_9891,N_9651);
nand UO_1146 (O_1146,N_9359,N_9625);
nor UO_1147 (O_1147,N_9160,N_9272);
nor UO_1148 (O_1148,N_9739,N_9068);
or UO_1149 (O_1149,N_9996,N_9916);
or UO_1150 (O_1150,N_9184,N_9658);
nand UO_1151 (O_1151,N_9703,N_9295);
and UO_1152 (O_1152,N_9386,N_9317);
or UO_1153 (O_1153,N_9006,N_9548);
nor UO_1154 (O_1154,N_9283,N_9660);
nand UO_1155 (O_1155,N_9454,N_9397);
and UO_1156 (O_1156,N_9978,N_9001);
nor UO_1157 (O_1157,N_9678,N_9357);
or UO_1158 (O_1158,N_9086,N_9697);
nor UO_1159 (O_1159,N_9886,N_9816);
or UO_1160 (O_1160,N_9521,N_9489);
xor UO_1161 (O_1161,N_9884,N_9742);
and UO_1162 (O_1162,N_9665,N_9580);
xnor UO_1163 (O_1163,N_9896,N_9327);
and UO_1164 (O_1164,N_9595,N_9455);
nor UO_1165 (O_1165,N_9538,N_9858);
and UO_1166 (O_1166,N_9001,N_9784);
xor UO_1167 (O_1167,N_9599,N_9783);
nor UO_1168 (O_1168,N_9462,N_9174);
nor UO_1169 (O_1169,N_9251,N_9009);
or UO_1170 (O_1170,N_9317,N_9185);
nand UO_1171 (O_1171,N_9737,N_9940);
and UO_1172 (O_1172,N_9526,N_9466);
nor UO_1173 (O_1173,N_9690,N_9508);
or UO_1174 (O_1174,N_9998,N_9475);
xor UO_1175 (O_1175,N_9209,N_9382);
nor UO_1176 (O_1176,N_9655,N_9620);
nand UO_1177 (O_1177,N_9238,N_9253);
or UO_1178 (O_1178,N_9935,N_9100);
nor UO_1179 (O_1179,N_9162,N_9888);
nand UO_1180 (O_1180,N_9848,N_9594);
and UO_1181 (O_1181,N_9196,N_9220);
and UO_1182 (O_1182,N_9131,N_9187);
and UO_1183 (O_1183,N_9498,N_9466);
and UO_1184 (O_1184,N_9551,N_9955);
nand UO_1185 (O_1185,N_9488,N_9602);
and UO_1186 (O_1186,N_9203,N_9022);
nand UO_1187 (O_1187,N_9569,N_9338);
and UO_1188 (O_1188,N_9147,N_9384);
nand UO_1189 (O_1189,N_9550,N_9771);
nor UO_1190 (O_1190,N_9107,N_9307);
xnor UO_1191 (O_1191,N_9435,N_9430);
xor UO_1192 (O_1192,N_9837,N_9656);
or UO_1193 (O_1193,N_9500,N_9769);
xnor UO_1194 (O_1194,N_9337,N_9019);
xor UO_1195 (O_1195,N_9988,N_9531);
and UO_1196 (O_1196,N_9014,N_9087);
or UO_1197 (O_1197,N_9851,N_9405);
xor UO_1198 (O_1198,N_9337,N_9569);
xnor UO_1199 (O_1199,N_9305,N_9012);
xor UO_1200 (O_1200,N_9730,N_9438);
nor UO_1201 (O_1201,N_9786,N_9216);
xor UO_1202 (O_1202,N_9763,N_9235);
nor UO_1203 (O_1203,N_9763,N_9467);
and UO_1204 (O_1204,N_9820,N_9062);
nor UO_1205 (O_1205,N_9810,N_9715);
xor UO_1206 (O_1206,N_9087,N_9358);
or UO_1207 (O_1207,N_9798,N_9862);
nand UO_1208 (O_1208,N_9383,N_9360);
and UO_1209 (O_1209,N_9482,N_9931);
xnor UO_1210 (O_1210,N_9825,N_9309);
nand UO_1211 (O_1211,N_9860,N_9480);
xor UO_1212 (O_1212,N_9301,N_9261);
or UO_1213 (O_1213,N_9434,N_9143);
or UO_1214 (O_1214,N_9210,N_9706);
or UO_1215 (O_1215,N_9329,N_9470);
or UO_1216 (O_1216,N_9529,N_9392);
xor UO_1217 (O_1217,N_9934,N_9422);
xnor UO_1218 (O_1218,N_9301,N_9342);
nor UO_1219 (O_1219,N_9585,N_9516);
nor UO_1220 (O_1220,N_9322,N_9423);
nor UO_1221 (O_1221,N_9265,N_9724);
xnor UO_1222 (O_1222,N_9988,N_9885);
xnor UO_1223 (O_1223,N_9202,N_9610);
or UO_1224 (O_1224,N_9377,N_9799);
nor UO_1225 (O_1225,N_9566,N_9283);
xor UO_1226 (O_1226,N_9134,N_9150);
and UO_1227 (O_1227,N_9297,N_9531);
nand UO_1228 (O_1228,N_9875,N_9903);
xor UO_1229 (O_1229,N_9041,N_9021);
and UO_1230 (O_1230,N_9060,N_9271);
and UO_1231 (O_1231,N_9586,N_9482);
or UO_1232 (O_1232,N_9176,N_9475);
nand UO_1233 (O_1233,N_9876,N_9989);
and UO_1234 (O_1234,N_9865,N_9206);
nand UO_1235 (O_1235,N_9168,N_9051);
xnor UO_1236 (O_1236,N_9854,N_9998);
nand UO_1237 (O_1237,N_9860,N_9979);
or UO_1238 (O_1238,N_9763,N_9054);
nand UO_1239 (O_1239,N_9992,N_9732);
nand UO_1240 (O_1240,N_9396,N_9763);
and UO_1241 (O_1241,N_9611,N_9815);
nor UO_1242 (O_1242,N_9732,N_9659);
nand UO_1243 (O_1243,N_9055,N_9292);
and UO_1244 (O_1244,N_9250,N_9810);
nand UO_1245 (O_1245,N_9831,N_9882);
or UO_1246 (O_1246,N_9097,N_9308);
or UO_1247 (O_1247,N_9167,N_9882);
or UO_1248 (O_1248,N_9570,N_9006);
nor UO_1249 (O_1249,N_9454,N_9507);
or UO_1250 (O_1250,N_9331,N_9134);
nor UO_1251 (O_1251,N_9955,N_9921);
nor UO_1252 (O_1252,N_9409,N_9431);
nand UO_1253 (O_1253,N_9826,N_9067);
nor UO_1254 (O_1254,N_9445,N_9485);
and UO_1255 (O_1255,N_9029,N_9164);
or UO_1256 (O_1256,N_9020,N_9779);
or UO_1257 (O_1257,N_9586,N_9848);
nand UO_1258 (O_1258,N_9133,N_9766);
or UO_1259 (O_1259,N_9621,N_9798);
nor UO_1260 (O_1260,N_9729,N_9611);
or UO_1261 (O_1261,N_9149,N_9695);
nand UO_1262 (O_1262,N_9759,N_9987);
xnor UO_1263 (O_1263,N_9477,N_9867);
nor UO_1264 (O_1264,N_9020,N_9081);
or UO_1265 (O_1265,N_9993,N_9835);
and UO_1266 (O_1266,N_9925,N_9019);
xnor UO_1267 (O_1267,N_9639,N_9098);
nand UO_1268 (O_1268,N_9747,N_9155);
nor UO_1269 (O_1269,N_9508,N_9888);
xor UO_1270 (O_1270,N_9915,N_9209);
or UO_1271 (O_1271,N_9913,N_9303);
xnor UO_1272 (O_1272,N_9466,N_9512);
nor UO_1273 (O_1273,N_9480,N_9372);
and UO_1274 (O_1274,N_9300,N_9449);
and UO_1275 (O_1275,N_9555,N_9711);
or UO_1276 (O_1276,N_9296,N_9874);
nand UO_1277 (O_1277,N_9854,N_9473);
nor UO_1278 (O_1278,N_9952,N_9563);
xnor UO_1279 (O_1279,N_9374,N_9172);
nor UO_1280 (O_1280,N_9018,N_9696);
and UO_1281 (O_1281,N_9058,N_9516);
nor UO_1282 (O_1282,N_9126,N_9665);
or UO_1283 (O_1283,N_9559,N_9560);
xor UO_1284 (O_1284,N_9113,N_9886);
or UO_1285 (O_1285,N_9117,N_9194);
and UO_1286 (O_1286,N_9557,N_9512);
or UO_1287 (O_1287,N_9160,N_9826);
and UO_1288 (O_1288,N_9752,N_9304);
or UO_1289 (O_1289,N_9046,N_9578);
and UO_1290 (O_1290,N_9208,N_9773);
or UO_1291 (O_1291,N_9128,N_9325);
nor UO_1292 (O_1292,N_9901,N_9728);
or UO_1293 (O_1293,N_9517,N_9310);
nor UO_1294 (O_1294,N_9289,N_9170);
or UO_1295 (O_1295,N_9626,N_9832);
nand UO_1296 (O_1296,N_9543,N_9139);
or UO_1297 (O_1297,N_9428,N_9028);
and UO_1298 (O_1298,N_9185,N_9899);
nand UO_1299 (O_1299,N_9254,N_9202);
xnor UO_1300 (O_1300,N_9965,N_9447);
or UO_1301 (O_1301,N_9228,N_9541);
or UO_1302 (O_1302,N_9469,N_9560);
or UO_1303 (O_1303,N_9357,N_9301);
nor UO_1304 (O_1304,N_9199,N_9241);
and UO_1305 (O_1305,N_9398,N_9738);
or UO_1306 (O_1306,N_9811,N_9270);
and UO_1307 (O_1307,N_9461,N_9589);
nand UO_1308 (O_1308,N_9730,N_9292);
or UO_1309 (O_1309,N_9579,N_9537);
nor UO_1310 (O_1310,N_9487,N_9194);
nor UO_1311 (O_1311,N_9831,N_9287);
and UO_1312 (O_1312,N_9456,N_9699);
and UO_1313 (O_1313,N_9669,N_9231);
nand UO_1314 (O_1314,N_9965,N_9594);
nor UO_1315 (O_1315,N_9276,N_9522);
and UO_1316 (O_1316,N_9258,N_9930);
xnor UO_1317 (O_1317,N_9303,N_9282);
nand UO_1318 (O_1318,N_9494,N_9245);
xor UO_1319 (O_1319,N_9054,N_9613);
nand UO_1320 (O_1320,N_9436,N_9877);
nand UO_1321 (O_1321,N_9911,N_9684);
nand UO_1322 (O_1322,N_9077,N_9224);
or UO_1323 (O_1323,N_9661,N_9929);
nor UO_1324 (O_1324,N_9883,N_9032);
and UO_1325 (O_1325,N_9549,N_9973);
nand UO_1326 (O_1326,N_9935,N_9481);
xor UO_1327 (O_1327,N_9132,N_9799);
nand UO_1328 (O_1328,N_9522,N_9896);
xor UO_1329 (O_1329,N_9082,N_9089);
nor UO_1330 (O_1330,N_9738,N_9594);
or UO_1331 (O_1331,N_9167,N_9492);
nor UO_1332 (O_1332,N_9322,N_9941);
and UO_1333 (O_1333,N_9080,N_9176);
or UO_1334 (O_1334,N_9172,N_9291);
or UO_1335 (O_1335,N_9608,N_9006);
and UO_1336 (O_1336,N_9390,N_9972);
nor UO_1337 (O_1337,N_9956,N_9199);
xor UO_1338 (O_1338,N_9870,N_9784);
nand UO_1339 (O_1339,N_9291,N_9351);
nor UO_1340 (O_1340,N_9510,N_9927);
xnor UO_1341 (O_1341,N_9045,N_9508);
or UO_1342 (O_1342,N_9750,N_9181);
nor UO_1343 (O_1343,N_9087,N_9093);
nand UO_1344 (O_1344,N_9396,N_9974);
or UO_1345 (O_1345,N_9929,N_9926);
xnor UO_1346 (O_1346,N_9701,N_9688);
xnor UO_1347 (O_1347,N_9080,N_9168);
and UO_1348 (O_1348,N_9663,N_9229);
xnor UO_1349 (O_1349,N_9519,N_9089);
and UO_1350 (O_1350,N_9943,N_9386);
xor UO_1351 (O_1351,N_9087,N_9577);
xor UO_1352 (O_1352,N_9658,N_9024);
xor UO_1353 (O_1353,N_9180,N_9044);
nor UO_1354 (O_1354,N_9852,N_9937);
or UO_1355 (O_1355,N_9073,N_9807);
and UO_1356 (O_1356,N_9181,N_9032);
nand UO_1357 (O_1357,N_9979,N_9117);
nand UO_1358 (O_1358,N_9329,N_9936);
nand UO_1359 (O_1359,N_9016,N_9602);
nor UO_1360 (O_1360,N_9608,N_9327);
nand UO_1361 (O_1361,N_9546,N_9014);
or UO_1362 (O_1362,N_9805,N_9908);
and UO_1363 (O_1363,N_9118,N_9878);
nand UO_1364 (O_1364,N_9011,N_9746);
nor UO_1365 (O_1365,N_9218,N_9030);
and UO_1366 (O_1366,N_9761,N_9821);
nand UO_1367 (O_1367,N_9356,N_9844);
or UO_1368 (O_1368,N_9657,N_9746);
or UO_1369 (O_1369,N_9843,N_9224);
nand UO_1370 (O_1370,N_9999,N_9840);
nand UO_1371 (O_1371,N_9829,N_9595);
nand UO_1372 (O_1372,N_9267,N_9855);
nand UO_1373 (O_1373,N_9149,N_9362);
and UO_1374 (O_1374,N_9491,N_9835);
or UO_1375 (O_1375,N_9654,N_9073);
nor UO_1376 (O_1376,N_9962,N_9149);
nor UO_1377 (O_1377,N_9066,N_9239);
xnor UO_1378 (O_1378,N_9614,N_9147);
and UO_1379 (O_1379,N_9808,N_9310);
nand UO_1380 (O_1380,N_9579,N_9924);
nand UO_1381 (O_1381,N_9581,N_9229);
xnor UO_1382 (O_1382,N_9065,N_9629);
xnor UO_1383 (O_1383,N_9250,N_9680);
or UO_1384 (O_1384,N_9631,N_9284);
xnor UO_1385 (O_1385,N_9660,N_9172);
nand UO_1386 (O_1386,N_9030,N_9026);
and UO_1387 (O_1387,N_9829,N_9869);
or UO_1388 (O_1388,N_9730,N_9454);
nand UO_1389 (O_1389,N_9968,N_9927);
or UO_1390 (O_1390,N_9023,N_9706);
nand UO_1391 (O_1391,N_9791,N_9523);
nor UO_1392 (O_1392,N_9821,N_9363);
xnor UO_1393 (O_1393,N_9519,N_9650);
or UO_1394 (O_1394,N_9400,N_9446);
nand UO_1395 (O_1395,N_9688,N_9355);
xnor UO_1396 (O_1396,N_9630,N_9136);
and UO_1397 (O_1397,N_9835,N_9014);
and UO_1398 (O_1398,N_9511,N_9418);
nand UO_1399 (O_1399,N_9659,N_9199);
and UO_1400 (O_1400,N_9522,N_9679);
nand UO_1401 (O_1401,N_9970,N_9007);
nand UO_1402 (O_1402,N_9561,N_9207);
nor UO_1403 (O_1403,N_9568,N_9623);
xnor UO_1404 (O_1404,N_9900,N_9982);
nand UO_1405 (O_1405,N_9005,N_9330);
nor UO_1406 (O_1406,N_9081,N_9591);
and UO_1407 (O_1407,N_9023,N_9492);
nand UO_1408 (O_1408,N_9856,N_9473);
and UO_1409 (O_1409,N_9359,N_9745);
nor UO_1410 (O_1410,N_9203,N_9990);
xor UO_1411 (O_1411,N_9835,N_9742);
nand UO_1412 (O_1412,N_9880,N_9363);
nor UO_1413 (O_1413,N_9732,N_9552);
and UO_1414 (O_1414,N_9161,N_9784);
nand UO_1415 (O_1415,N_9724,N_9761);
nor UO_1416 (O_1416,N_9654,N_9093);
xnor UO_1417 (O_1417,N_9360,N_9553);
nor UO_1418 (O_1418,N_9727,N_9567);
xor UO_1419 (O_1419,N_9573,N_9271);
nand UO_1420 (O_1420,N_9354,N_9025);
and UO_1421 (O_1421,N_9751,N_9562);
and UO_1422 (O_1422,N_9054,N_9689);
or UO_1423 (O_1423,N_9847,N_9741);
or UO_1424 (O_1424,N_9254,N_9382);
or UO_1425 (O_1425,N_9448,N_9476);
or UO_1426 (O_1426,N_9712,N_9995);
and UO_1427 (O_1427,N_9857,N_9105);
and UO_1428 (O_1428,N_9007,N_9987);
and UO_1429 (O_1429,N_9840,N_9042);
nand UO_1430 (O_1430,N_9205,N_9628);
and UO_1431 (O_1431,N_9784,N_9416);
or UO_1432 (O_1432,N_9939,N_9078);
nand UO_1433 (O_1433,N_9589,N_9245);
nand UO_1434 (O_1434,N_9571,N_9222);
nor UO_1435 (O_1435,N_9317,N_9300);
or UO_1436 (O_1436,N_9769,N_9745);
and UO_1437 (O_1437,N_9077,N_9017);
and UO_1438 (O_1438,N_9799,N_9680);
nand UO_1439 (O_1439,N_9087,N_9486);
or UO_1440 (O_1440,N_9415,N_9819);
or UO_1441 (O_1441,N_9986,N_9392);
or UO_1442 (O_1442,N_9390,N_9962);
or UO_1443 (O_1443,N_9109,N_9277);
xor UO_1444 (O_1444,N_9382,N_9173);
xor UO_1445 (O_1445,N_9774,N_9939);
nor UO_1446 (O_1446,N_9632,N_9446);
or UO_1447 (O_1447,N_9551,N_9198);
nor UO_1448 (O_1448,N_9357,N_9889);
nor UO_1449 (O_1449,N_9278,N_9452);
and UO_1450 (O_1450,N_9918,N_9451);
xnor UO_1451 (O_1451,N_9891,N_9461);
nand UO_1452 (O_1452,N_9109,N_9293);
nor UO_1453 (O_1453,N_9313,N_9179);
and UO_1454 (O_1454,N_9328,N_9187);
nor UO_1455 (O_1455,N_9485,N_9544);
nor UO_1456 (O_1456,N_9068,N_9537);
xnor UO_1457 (O_1457,N_9770,N_9887);
and UO_1458 (O_1458,N_9189,N_9822);
nand UO_1459 (O_1459,N_9093,N_9238);
nor UO_1460 (O_1460,N_9292,N_9198);
xor UO_1461 (O_1461,N_9483,N_9223);
and UO_1462 (O_1462,N_9827,N_9883);
xnor UO_1463 (O_1463,N_9893,N_9964);
nand UO_1464 (O_1464,N_9391,N_9050);
xor UO_1465 (O_1465,N_9374,N_9480);
xor UO_1466 (O_1466,N_9182,N_9174);
nor UO_1467 (O_1467,N_9801,N_9762);
nand UO_1468 (O_1468,N_9172,N_9672);
xnor UO_1469 (O_1469,N_9133,N_9471);
nand UO_1470 (O_1470,N_9068,N_9604);
xor UO_1471 (O_1471,N_9420,N_9387);
xor UO_1472 (O_1472,N_9644,N_9503);
xnor UO_1473 (O_1473,N_9244,N_9608);
or UO_1474 (O_1474,N_9068,N_9120);
nor UO_1475 (O_1475,N_9392,N_9066);
or UO_1476 (O_1476,N_9049,N_9900);
nor UO_1477 (O_1477,N_9033,N_9629);
nand UO_1478 (O_1478,N_9266,N_9804);
nand UO_1479 (O_1479,N_9465,N_9796);
xor UO_1480 (O_1480,N_9698,N_9832);
xor UO_1481 (O_1481,N_9556,N_9206);
or UO_1482 (O_1482,N_9715,N_9046);
xor UO_1483 (O_1483,N_9479,N_9440);
xnor UO_1484 (O_1484,N_9224,N_9645);
nor UO_1485 (O_1485,N_9566,N_9168);
nand UO_1486 (O_1486,N_9715,N_9956);
or UO_1487 (O_1487,N_9017,N_9313);
xor UO_1488 (O_1488,N_9208,N_9427);
or UO_1489 (O_1489,N_9236,N_9079);
nand UO_1490 (O_1490,N_9780,N_9959);
and UO_1491 (O_1491,N_9787,N_9872);
or UO_1492 (O_1492,N_9956,N_9948);
and UO_1493 (O_1493,N_9871,N_9458);
xor UO_1494 (O_1494,N_9391,N_9473);
nand UO_1495 (O_1495,N_9140,N_9248);
nor UO_1496 (O_1496,N_9540,N_9041);
nor UO_1497 (O_1497,N_9805,N_9207);
nor UO_1498 (O_1498,N_9081,N_9407);
nor UO_1499 (O_1499,N_9855,N_9299);
endmodule