module basic_2000_20000_2500_4_levels_1xor_2(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999;
or U0 (N_0,In_150,In_378);
and U1 (N_1,In_1462,In_1495);
nor U2 (N_2,In_1506,In_546);
nor U3 (N_3,In_1617,In_909);
nand U4 (N_4,In_1902,In_46);
nand U5 (N_5,In_1421,In_1610);
or U6 (N_6,In_826,In_122);
or U7 (N_7,In_369,In_1535);
xor U8 (N_8,In_932,In_544);
or U9 (N_9,In_960,In_217);
nand U10 (N_10,In_259,In_836);
nor U11 (N_11,In_1956,In_1991);
and U12 (N_12,In_1411,In_1728);
nand U13 (N_13,In_509,In_1623);
nor U14 (N_14,In_1512,In_1584);
and U15 (N_15,In_72,In_481);
and U16 (N_16,In_1268,In_1895);
nor U17 (N_17,In_375,In_1081);
nor U18 (N_18,In_1191,In_1447);
and U19 (N_19,In_1550,In_356);
or U20 (N_20,In_336,In_283);
and U21 (N_21,In_109,In_1739);
nand U22 (N_22,In_348,In_799);
or U23 (N_23,In_1139,In_1492);
nand U24 (N_24,In_947,In_1886);
nand U25 (N_25,In_434,In_1430);
or U26 (N_26,In_950,In_271);
nand U27 (N_27,In_151,In_1939);
and U28 (N_28,In_115,In_535);
and U29 (N_29,In_1523,In_408);
or U30 (N_30,In_769,In_1515);
or U31 (N_31,In_738,In_765);
and U32 (N_32,In_508,In_442);
or U33 (N_33,In_1772,In_1799);
or U34 (N_34,In_1432,In_1793);
and U35 (N_35,In_315,In_444);
nand U36 (N_36,In_937,In_1358);
nand U37 (N_37,In_76,In_349);
or U38 (N_38,In_1625,In_170);
or U39 (N_39,In_1582,In_1273);
nor U40 (N_40,In_1213,In_1392);
and U41 (N_41,In_1335,In_404);
nand U42 (N_42,In_1169,In_751);
and U43 (N_43,In_865,In_8);
and U44 (N_44,In_298,In_541);
and U45 (N_45,In_1572,In_207);
and U46 (N_46,In_1732,In_1463);
or U47 (N_47,In_629,In_1877);
and U48 (N_48,In_1456,In_618);
and U49 (N_49,In_1442,In_301);
nor U50 (N_50,In_563,In_938);
nor U51 (N_51,In_665,In_1056);
xor U52 (N_52,In_126,In_44);
and U53 (N_53,In_286,In_80);
nor U54 (N_54,In_174,In_986);
and U55 (N_55,In_1669,In_1344);
nand U56 (N_56,In_427,In_319);
nor U57 (N_57,In_391,In_1935);
nand U58 (N_58,In_1321,In_658);
nor U59 (N_59,In_995,In_1600);
nor U60 (N_60,In_1223,In_48);
or U61 (N_61,In_1088,In_1755);
nor U62 (N_62,In_467,In_575);
or U63 (N_63,In_1901,In_307);
and U64 (N_64,In_29,In_1745);
nor U65 (N_65,In_1657,In_700);
nand U66 (N_66,In_915,In_609);
nand U67 (N_67,In_979,In_141);
and U68 (N_68,In_1632,In_308);
nor U69 (N_69,In_204,In_1685);
or U70 (N_70,In_884,In_1178);
nand U71 (N_71,In_1468,In_441);
nor U72 (N_72,In_1194,In_1561);
or U73 (N_73,In_334,In_1687);
or U74 (N_74,In_1014,In_709);
or U75 (N_75,In_859,In_1326);
nand U76 (N_76,In_635,In_985);
and U77 (N_77,In_1378,In_1848);
or U78 (N_78,In_1148,In_1385);
nor U79 (N_79,In_1648,In_214);
or U80 (N_80,In_1470,In_129);
nand U81 (N_81,In_1706,In_764);
nor U82 (N_82,In_1634,In_523);
and U83 (N_83,In_341,In_233);
or U84 (N_84,In_1283,In_579);
nand U85 (N_85,In_279,In_412);
or U86 (N_86,In_1481,In_23);
or U87 (N_87,In_1845,In_1419);
nand U88 (N_88,In_1309,In_149);
nor U89 (N_89,In_147,In_1949);
nor U90 (N_90,In_838,In_978);
and U91 (N_91,In_388,In_191);
and U92 (N_92,In_847,In_89);
nor U93 (N_93,In_1409,In_90);
or U94 (N_94,In_976,In_1460);
or U95 (N_95,In_866,In_1620);
nand U96 (N_96,In_1133,In_990);
or U97 (N_97,In_1597,In_379);
nand U98 (N_98,In_921,In_1237);
nor U99 (N_99,In_768,In_241);
or U100 (N_100,In_262,In_250);
or U101 (N_101,In_697,In_1444);
and U102 (N_102,In_1143,In_1259);
nor U103 (N_103,In_657,In_1461);
or U104 (N_104,In_1814,In_186);
or U105 (N_105,In_1067,In_649);
nand U106 (N_106,In_57,In_456);
or U107 (N_107,In_1812,In_132);
nand U108 (N_108,In_144,In_1227);
nor U109 (N_109,In_1406,In_519);
nor U110 (N_110,In_1941,In_719);
nor U111 (N_111,In_1693,In_1068);
nor U112 (N_112,In_1182,In_1719);
and U113 (N_113,In_1538,In_928);
nor U114 (N_114,In_748,In_722);
or U115 (N_115,In_1602,In_430);
and U116 (N_116,In_874,In_585);
nand U117 (N_117,In_1472,In_1490);
nor U118 (N_118,In_1501,In_892);
or U119 (N_119,In_531,In_1542);
nor U120 (N_120,In_1342,In_1959);
nand U121 (N_121,In_1498,In_184);
and U122 (N_122,In_1312,In_1170);
or U123 (N_123,In_1705,In_1933);
nor U124 (N_124,In_1675,In_1818);
or U125 (N_125,In_428,In_426);
or U126 (N_126,In_1063,In_86);
nand U127 (N_127,In_1496,In_1080);
nor U128 (N_128,In_196,In_824);
nor U129 (N_129,In_257,In_1744);
or U130 (N_130,In_295,In_1436);
and U131 (N_131,In_490,In_347);
and U132 (N_132,In_782,In_1164);
or U133 (N_133,In_888,In_1806);
and U134 (N_134,In_1244,In_1373);
nor U135 (N_135,In_302,In_1938);
nand U136 (N_136,In_91,In_1709);
nor U137 (N_137,In_1364,In_202);
and U138 (N_138,In_1219,In_708);
nor U139 (N_139,In_1296,In_294);
and U140 (N_140,In_1779,In_1811);
or U141 (N_141,In_561,In_371);
nor U142 (N_142,In_226,In_1547);
and U143 (N_143,In_623,In_676);
and U144 (N_144,In_63,In_724);
nor U145 (N_145,In_612,In_1489);
nand U146 (N_146,In_203,In_1165);
nor U147 (N_147,In_613,In_1817);
and U148 (N_148,In_1784,In_1688);
or U149 (N_149,In_1246,In_1270);
and U150 (N_150,In_1382,In_580);
and U151 (N_151,In_1247,In_1915);
nand U152 (N_152,In_515,In_367);
and U153 (N_153,In_1149,In_447);
and U154 (N_154,In_582,In_199);
nand U155 (N_155,In_377,In_694);
nand U156 (N_156,In_479,In_660);
and U157 (N_157,In_1345,In_1913);
nand U158 (N_158,In_567,In_1986);
or U159 (N_159,In_886,In_1328);
and U160 (N_160,In_1885,In_1236);
and U161 (N_161,In_125,In_1960);
nand U162 (N_162,In_1307,In_1361);
nor U163 (N_163,In_1887,In_1850);
and U164 (N_164,In_641,In_1950);
or U165 (N_165,In_1565,In_789);
nand U166 (N_166,In_60,In_58);
nand U167 (N_167,In_1588,In_930);
nor U168 (N_168,In_1137,In_1519);
nor U169 (N_169,In_926,In_633);
nand U170 (N_170,In_754,In_1104);
and U171 (N_171,In_1131,In_1847);
or U172 (N_172,In_1184,In_1423);
and U173 (N_173,In_1961,In_972);
or U174 (N_174,In_1062,In_1893);
nor U175 (N_175,In_1931,In_79);
nand U176 (N_176,In_807,In_1537);
nor U177 (N_177,In_1993,In_472);
or U178 (N_178,In_1973,In_1029);
or U179 (N_179,In_445,In_981);
nor U180 (N_180,In_1408,In_1243);
nand U181 (N_181,In_1039,In_105);
nand U182 (N_182,In_1381,In_464);
nor U183 (N_183,In_1253,In_1510);
nor U184 (N_184,In_520,In_1690);
and U185 (N_185,In_1614,In_646);
nor U186 (N_186,In_1872,In_363);
or U187 (N_187,In_1770,In_1022);
nor U188 (N_188,In_1658,In_999);
nand U189 (N_189,In_954,In_1952);
and U190 (N_190,In_1252,In_331);
and U191 (N_191,In_462,In_620);
nand U192 (N_192,In_992,In_1372);
nand U193 (N_193,In_1028,In_1504);
nand U194 (N_194,In_1094,In_143);
or U195 (N_195,In_1676,In_1593);
nor U196 (N_196,In_1999,In_1867);
or U197 (N_197,In_316,In_848);
or U198 (N_198,In_664,In_589);
nand U199 (N_199,In_452,In_154);
nand U200 (N_200,In_1718,In_94);
nor U201 (N_201,In_1396,In_550);
or U202 (N_202,In_800,In_415);
and U203 (N_203,In_291,In_1363);
or U204 (N_204,In_1909,In_417);
nand U205 (N_205,In_374,In_153);
or U206 (N_206,In_1533,In_1248);
nand U207 (N_207,In_1526,In_77);
nor U208 (N_208,In_1633,In_1558);
nor U209 (N_209,In_1813,In_525);
and U210 (N_210,In_1391,In_1486);
nor U211 (N_211,In_698,In_624);
nor U212 (N_212,In_1666,In_970);
nor U213 (N_213,In_35,In_1107);
or U214 (N_214,In_1226,In_306);
nor U215 (N_215,In_766,In_1305);
nor U216 (N_216,In_268,In_1857);
and U217 (N_217,In_574,In_1790);
or U218 (N_218,In_1616,In_84);
nand U219 (N_219,In_1796,In_171);
nand U220 (N_220,In_484,In_1458);
nor U221 (N_221,In_514,In_1323);
or U222 (N_222,In_50,In_1077);
nor U223 (N_223,In_1032,In_1948);
or U224 (N_224,In_1794,In_1389);
nor U225 (N_225,In_872,In_1776);
and U226 (N_226,In_1860,In_1311);
nor U227 (N_227,In_453,In_1769);
or U228 (N_228,In_736,In_1734);
nor U229 (N_229,In_1866,In_267);
or U230 (N_230,In_1507,In_1890);
and U231 (N_231,In_1701,In_335);
nand U232 (N_232,In_617,In_263);
and U233 (N_233,In_1166,In_409);
nor U234 (N_234,In_1645,In_9);
and U235 (N_235,In_743,In_54);
or U236 (N_236,In_1635,In_1762);
nand U237 (N_237,In_1609,In_1820);
nor U238 (N_238,In_364,In_1724);
nor U239 (N_239,In_1232,In_1439);
and U240 (N_240,In_1211,In_1575);
nor U241 (N_241,In_1332,In_390);
nand U242 (N_242,In_1092,In_1167);
nor U243 (N_243,In_64,In_1228);
nand U244 (N_244,In_465,In_43);
nor U245 (N_245,In_123,In_964);
nor U246 (N_246,In_1318,In_1262);
nor U247 (N_247,In_1066,In_1831);
or U248 (N_248,In_1070,In_1892);
nand U249 (N_249,In_1919,In_616);
or U250 (N_250,In_784,In_366);
nand U251 (N_251,In_25,In_440);
nor U252 (N_252,In_56,In_1752);
and U253 (N_253,In_1402,In_1074);
or U254 (N_254,In_274,In_1388);
xor U255 (N_255,In_1543,In_41);
and U256 (N_256,In_1753,In_399);
nand U257 (N_257,In_931,In_1578);
and U258 (N_258,In_463,In_1454);
and U259 (N_259,In_177,In_678);
and U260 (N_260,In_429,In_1007);
nor U261 (N_261,In_1929,In_1521);
nor U262 (N_262,In_1301,In_1132);
nor U263 (N_263,In_540,In_1789);
nand U264 (N_264,In_1216,In_1638);
nand U265 (N_265,In_1006,In_548);
or U266 (N_266,In_1837,In_1716);
or U267 (N_267,In_1240,In_1466);
or U268 (N_268,In_673,In_672);
nand U269 (N_269,In_292,In_1004);
and U270 (N_270,In_1873,In_881);
and U271 (N_271,In_1256,In_1299);
nand U272 (N_272,In_1862,In_967);
nor U273 (N_273,In_1766,In_137);
nand U274 (N_274,In_1955,In_730);
and U275 (N_275,In_1390,In_275);
or U276 (N_276,In_398,In_1918);
nor U277 (N_277,In_750,In_1355);
or U278 (N_278,In_1261,In_1671);
nand U279 (N_279,In_342,In_804);
and U280 (N_280,In_242,In_1703);
nor U281 (N_281,In_1138,In_1413);
nand U282 (N_282,In_49,In_1613);
or U283 (N_283,In_725,In_278);
nand U284 (N_284,In_901,In_338);
nor U285 (N_285,In_209,In_1978);
or U286 (N_286,In_1567,In_1069);
or U287 (N_287,In_1589,In_1276);
and U288 (N_288,In_7,In_433);
nor U289 (N_289,In_785,In_818);
nand U290 (N_290,In_449,In_584);
nor U291 (N_291,In_1591,In_1469);
and U292 (N_292,In_1383,In_707);
xnor U293 (N_293,In_1655,In_1522);
nand U294 (N_294,In_1225,In_1025);
or U295 (N_295,In_1883,In_1241);
nor U296 (N_296,In_1829,In_1109);
or U297 (N_297,In_1083,In_436);
nand U298 (N_298,In_756,In_194);
nand U299 (N_299,In_1622,In_438);
nor U300 (N_300,In_1827,In_419);
nand U301 (N_301,In_510,In_1921);
or U302 (N_302,In_236,In_912);
nand U303 (N_303,In_1084,In_1947);
and U304 (N_304,In_368,In_1038);
nor U305 (N_305,In_1042,In_1962);
or U306 (N_306,In_1023,In_1146);
nand U307 (N_307,In_1816,In_1096);
nor U308 (N_308,In_1097,In_1422);
or U309 (N_309,In_640,In_47);
nand U310 (N_310,In_88,In_831);
or U311 (N_311,In_1995,In_66);
and U312 (N_312,In_834,In_1863);
and U313 (N_313,In_588,In_1777);
or U314 (N_314,In_647,In_537);
nor U315 (N_315,In_1128,In_1833);
nor U316 (N_316,In_713,In_324);
and U317 (N_317,In_1677,In_1568);
and U318 (N_318,In_993,In_396);
nand U319 (N_319,In_1606,In_99);
nor U320 (N_320,In_1375,In_536);
and U321 (N_321,In_835,In_98);
nand U322 (N_322,In_1729,In_1387);
and U323 (N_323,In_1541,In_936);
nand U324 (N_324,In_1682,In_1087);
and U325 (N_325,In_1041,In_997);
nand U326 (N_326,In_1912,In_968);
nand U327 (N_327,In_205,In_503);
nor U328 (N_328,In_1304,In_1015);
nand U329 (N_329,In_1369,In_1162);
xor U330 (N_330,In_1297,In_1204);
nor U331 (N_331,In_1187,In_944);
nand U332 (N_332,In_630,In_95);
or U333 (N_333,In_586,In_593);
or U334 (N_334,In_1819,In_432);
or U335 (N_335,In_220,In_1545);
and U336 (N_336,In_1186,In_254);
or U337 (N_337,In_1446,In_116);
nor U338 (N_338,In_1577,In_849);
and U339 (N_339,In_1516,In_1269);
nor U340 (N_340,In_1053,In_735);
and U341 (N_341,In_1574,In_1539);
or U342 (N_342,In_989,In_919);
and U343 (N_343,In_437,In_712);
nor U344 (N_344,In_505,In_1267);
or U345 (N_345,In_1631,In_684);
nand U346 (N_346,In_1731,In_1856);
nand U347 (N_347,In_1198,In_1058);
nor U348 (N_348,In_1122,In_382);
or U349 (N_349,In_829,In_1977);
nand U350 (N_350,In_656,In_330);
or U351 (N_351,In_857,In_114);
or U352 (N_352,In_1713,In_1778);
nand U353 (N_353,In_1880,In_140);
and U354 (N_354,In_1764,In_1985);
and U355 (N_355,In_1156,In_603);
or U356 (N_356,In_1964,In_104);
and U357 (N_357,In_1019,In_309);
nand U358 (N_358,In_975,In_1659);
nand U359 (N_359,In_100,In_1548);
and U360 (N_360,In_1319,In_1502);
and U361 (N_361,In_1113,In_329);
nor U362 (N_362,In_558,In_1882);
nor U363 (N_363,In_1479,In_1888);
nand U364 (N_364,In_1289,In_1599);
nor U365 (N_365,In_1802,In_1485);
and U366 (N_366,In_1168,In_887);
or U367 (N_367,In_1736,In_496);
or U368 (N_368,In_853,In_1836);
and U369 (N_369,In_67,In_569);
nand U370 (N_370,In_475,In_1528);
or U371 (N_371,In_1377,In_1281);
xnor U372 (N_372,In_512,In_1740);
nand U373 (N_373,In_247,In_1043);
and U374 (N_374,In_552,In_457);
nor U375 (N_375,In_1288,In_661);
nand U376 (N_376,In_825,In_353);
nor U377 (N_377,In_811,In_1425);
or U378 (N_378,In_255,In_922);
nand U379 (N_379,In_1927,In_819);
or U380 (N_380,In_1086,In_1242);
nand U381 (N_381,In_855,In_1989);
nand U382 (N_382,In_1354,In_1551);
or U383 (N_383,In_42,In_957);
or U384 (N_384,In_1210,In_1202);
nand U385 (N_385,In_1220,In_1171);
or U386 (N_386,In_1988,In_918);
nand U387 (N_387,In_1556,In_328);
nor U388 (N_388,In_17,In_28);
nor U389 (N_389,In_790,In_393);
or U390 (N_390,In_636,In_1636);
and U391 (N_391,In_1293,In_160);
nor U392 (N_392,In_211,In_1735);
or U393 (N_393,In_1870,In_333);
nand U394 (N_394,In_1160,In_699);
or U395 (N_395,In_1742,In_394);
nor U396 (N_396,In_461,In_856);
and U397 (N_397,In_1386,In_326);
nor U398 (N_398,In_833,In_1130);
nor U399 (N_399,In_682,In_591);
or U400 (N_400,In_411,In_1982);
or U401 (N_401,In_424,In_459);
and U402 (N_402,In_622,In_714);
nor U403 (N_403,In_680,In_343);
or U404 (N_404,In_1590,In_1426);
nand U405 (N_405,In_945,In_534);
and U406 (N_406,In_860,In_1157);
nor U407 (N_407,In_1608,In_704);
and U408 (N_408,In_1177,In_1928);
or U409 (N_409,In_573,In_1452);
nor U410 (N_410,In_1975,In_282);
or U411 (N_411,In_1457,In_499);
nor U412 (N_412,In_1530,In_1708);
and U413 (N_413,In_1493,In_1260);
nor U414 (N_414,In_1410,In_837);
nand U415 (N_415,In_594,In_1050);
and U416 (N_416,In_923,In_1864);
and U417 (N_417,In_1559,In_621);
nor U418 (N_418,In_953,In_1840);
or U419 (N_419,In_1250,In_733);
or U420 (N_420,In_71,In_1680);
nor U421 (N_421,In_16,In_101);
and U422 (N_422,In_1844,In_677);
and U423 (N_423,In_1189,In_1005);
nand U424 (N_424,In_361,In_1771);
or U425 (N_425,In_683,In_1180);
nand U426 (N_426,In_1757,In_788);
or U427 (N_427,In_1224,In_1427);
or U428 (N_428,In_1945,In_120);
nor U429 (N_429,In_281,In_21);
nor U430 (N_430,In_1418,In_1879);
nand U431 (N_431,In_1103,In_1925);
and U432 (N_432,In_767,In_898);
or U433 (N_433,In_1615,In_20);
nor U434 (N_434,In_1774,In_1111);
and U435 (N_435,In_1641,In_169);
nor U436 (N_436,In_1271,In_270);
nor U437 (N_437,In_688,In_1197);
nand U438 (N_438,In_476,In_1370);
and U439 (N_439,In_1183,In_1518);
or U440 (N_440,In_600,In_1403);
nor U441 (N_441,In_1839,In_200);
nor U442 (N_442,In_422,In_1531);
nor U443 (N_443,In_572,In_373);
nor U444 (N_444,In_1483,In_1804);
and U445 (N_445,In_372,In_1822);
or U446 (N_446,In_1116,In_245);
or U447 (N_447,In_181,In_131);
nor U448 (N_448,In_69,In_178);
or U449 (N_449,In_1497,In_414);
nor U450 (N_450,In_1765,In_235);
nand U451 (N_451,In_1044,In_528);
or U452 (N_452,In_491,In_486);
nand U453 (N_453,In_397,In_1749);
and U454 (N_454,In_108,In_1937);
nand U455 (N_455,In_296,In_867);
nor U456 (N_456,In_6,In_1333);
or U457 (N_457,In_244,In_781);
nor U458 (N_458,In_1562,In_1917);
nand U459 (N_459,In_24,In_431);
and U460 (N_460,In_1192,In_1153);
or U461 (N_461,In_631,In_345);
and U462 (N_462,In_466,In_1683);
nand U463 (N_463,In_1594,In_304);
or U464 (N_464,In_1871,In_1637);
nand U465 (N_465,In_1453,In_210);
xnor U466 (N_466,In_213,In_1027);
and U467 (N_467,In_741,In_1320);
and U468 (N_468,In_74,In_581);
and U469 (N_469,In_1722,In_933);
and U470 (N_470,In_159,In_1121);
and U471 (N_471,In_272,In_606);
and U472 (N_472,In_1287,In_206);
nor U473 (N_473,In_300,In_1815);
nor U474 (N_474,In_13,In_805);
nor U475 (N_475,In_1958,In_1595);
nor U476 (N_476,In_317,In_1112);
nand U477 (N_477,In_70,In_798);
and U478 (N_478,In_899,In_1400);
and U479 (N_479,In_451,In_493);
or U480 (N_480,In_142,In_500);
or U481 (N_481,In_1583,In_1906);
nand U482 (N_482,In_365,In_942);
nand U483 (N_483,In_1546,In_906);
and U484 (N_484,In_82,In_470);
nand U485 (N_485,In_1117,In_998);
and U486 (N_486,In_823,In_1026);
nor U487 (N_487,In_1957,In_4);
and U488 (N_488,In_1329,In_1334);
or U489 (N_489,In_1003,In_547);
or U490 (N_490,In_1415,In_1254);
or U491 (N_491,In_1348,In_792);
nor U492 (N_492,In_1758,In_1011);
and U493 (N_493,In_1279,In_22);
or U494 (N_494,In_1911,In_1351);
and U495 (N_495,In_1689,In_951);
nand U496 (N_496,In_744,In_655);
and U497 (N_497,In_717,In_1336);
nand U498 (N_498,In_182,In_1517);
or U499 (N_499,In_1030,In_775);
nand U500 (N_500,In_243,In_1141);
nand U501 (N_501,In_1163,In_1394);
or U502 (N_502,In_1048,In_237);
nand U503 (N_503,In_1549,In_305);
nand U504 (N_504,In_198,In_354);
nand U505 (N_505,In_776,In_1896);
xor U506 (N_506,In_321,In_794);
nor U507 (N_507,In_956,In_1313);
and U508 (N_508,In_1711,In_1298);
nor U509 (N_509,In_1748,In_1580);
nor U510 (N_510,In_1897,In_1098);
and U511 (N_511,In_1073,In_1316);
and U512 (N_512,In_1598,In_763);
nor U513 (N_513,In_340,In_62);
or U514 (N_514,In_851,In_614);
nand U515 (N_515,In_1476,In_996);
nand U516 (N_516,In_1859,In_966);
or U517 (N_517,In_1434,In_844);
nor U518 (N_518,In_723,In_359);
and U519 (N_519,In_1868,In_891);
nand U520 (N_520,In_504,In_346);
nand U521 (N_521,In_1759,In_1398);
or U522 (N_522,In_113,In_1437);
and U523 (N_523,In_1308,In_1205);
nand U524 (N_524,In_1324,In_1071);
or U525 (N_525,In_1079,In_727);
nand U526 (N_526,In_124,In_135);
and U527 (N_527,In_809,In_1773);
or U528 (N_528,In_796,In_1662);
or U529 (N_529,In_1105,In_566);
and U530 (N_530,In_1478,In_1215);
and U531 (N_531,In_1020,In_941);
nand U532 (N_532,In_1035,In_1554);
nor U533 (N_533,In_994,In_925);
nor U534 (N_534,In_1294,In_869);
or U535 (N_535,In_1951,In_770);
nor U536 (N_536,In_188,In_1723);
nand U537 (N_537,In_1717,In_1756);
and U538 (N_538,In_51,In_895);
or U539 (N_539,In_1557,In_908);
nor U540 (N_540,In_92,In_420);
and U541 (N_541,In_1953,In_940);
xnor U542 (N_542,In_659,In_55);
and U543 (N_543,In_403,In_1810);
or U544 (N_544,In_1401,In_93);
and U545 (N_545,In_916,In_690);
or U546 (N_546,In_786,In_197);
and U547 (N_547,In_0,In_1399);
and U548 (N_548,In_1229,In_1331);
nand U549 (N_549,In_1946,In_667);
and U550 (N_550,In_252,In_1278);
nor U551 (N_551,In_1,In_290);
nand U552 (N_552,In_497,In_1359);
nand U553 (N_553,In_1586,In_386);
or U554 (N_554,In_1272,In_842);
or U555 (N_555,In_1181,In_128);
nor U556 (N_556,In_1926,In_1852);
nand U557 (N_557,In_1788,In_224);
and U558 (N_558,In_1916,In_896);
and U559 (N_559,In_1750,In_1983);
or U560 (N_560,In_774,In_1529);
and U561 (N_561,In_1987,In_795);
nor U562 (N_562,In_1291,In_545);
nand U563 (N_563,In_1894,In_1563);
or U564 (N_564,In_1057,In_653);
and U565 (N_565,In_965,In_38);
and U566 (N_566,In_1093,In_33);
nor U567 (N_567,In_1930,In_679);
or U568 (N_568,In_734,In_1553);
and U569 (N_569,In_982,In_1341);
nand U570 (N_570,In_1125,In_75);
nor U571 (N_571,In_1440,In_1037);
or U572 (N_572,In_392,In_332);
nor U573 (N_573,In_991,In_1825);
or U574 (N_574,In_527,In_1905);
xnor U575 (N_575,In_1830,In_1159);
and U576 (N_576,In_533,In_894);
and U577 (N_577,In_1222,In_1646);
nor U578 (N_578,In_1823,In_1161);
or U579 (N_579,In_877,In_1998);
or U580 (N_580,In_1325,In_1801);
nor U581 (N_581,In_557,In_549);
nand U582 (N_582,In_350,In_195);
and U583 (N_583,In_180,In_1208);
and U584 (N_584,In_1448,In_755);
and U585 (N_585,In_914,In_266);
nor U586 (N_586,In_362,In_376);
or U587 (N_587,In_726,In_1809);
or U588 (N_588,In_1621,In_1257);
nand U589 (N_589,In_863,In_1420);
and U590 (N_590,In_828,In_1624);
and U591 (N_591,In_1738,In_793);
nor U592 (N_592,In_1746,In_360);
nand U593 (N_593,In_753,In_78);
and U594 (N_594,In_639,In_858);
nor U595 (N_595,In_1349,In_1834);
and U596 (N_596,In_1842,In_1644);
nand U597 (N_597,In_1564,In_1994);
nor U598 (N_598,In_761,In_903);
and U599 (N_599,In_228,In_1480);
and U600 (N_600,In_448,In_249);
nand U601 (N_601,In_791,In_1775);
nor U602 (N_602,In_1040,In_779);
and U603 (N_603,In_783,In_477);
nand U604 (N_604,In_1878,In_1710);
or U605 (N_605,In_1969,In_662);
nor U606 (N_606,In_406,In_185);
or U607 (N_607,In_1433,In_1861);
nand U608 (N_608,In_880,In_1142);
and U609 (N_609,In_615,In_1154);
and U610 (N_610,In_605,In_1200);
and U611 (N_611,In_1932,In_1049);
nor U612 (N_612,In_1763,In_175);
xor U613 (N_613,In_821,In_402);
nor U614 (N_614,In_568,In_889);
nand U615 (N_615,In_1119,In_1797);
nand U616 (N_616,In_216,In_839);
nor U617 (N_617,In_1924,In_166);
or U618 (N_618,In_383,In_1158);
and U619 (N_619,In_1838,In_1395);
and U620 (N_620,In_560,In_1136);
nand U621 (N_621,In_701,In_161);
or U622 (N_622,In_551,In_1347);
or U623 (N_623,In_1376,In_961);
and U624 (N_624,In_421,In_111);
or U625 (N_625,In_506,In_1630);
nand U626 (N_626,In_102,In_1571);
or U627 (N_627,In_1235,In_758);
nor U628 (N_628,In_1920,In_1832);
nand U629 (N_629,In_1715,In_480);
nand U630 (N_630,In_1108,In_1465);
nand U631 (N_631,In_642,In_1371);
nor U632 (N_632,In_974,In_1397);
nand U633 (N_633,In_1781,In_320);
and U634 (N_634,In_787,In_529);
or U635 (N_635,In_269,In_1876);
nand U636 (N_636,In_273,In_1099);
or U637 (N_637,In_1033,In_1127);
nand U638 (N_638,In_873,In_1356);
nand U639 (N_639,In_742,In_797);
or U640 (N_640,In_310,In_1218);
nand U641 (N_641,In_777,In_1743);
or U642 (N_642,In_760,In_820);
nand U643 (N_643,In_778,In_1449);
and U644 (N_644,In_543,In_927);
and U645 (N_645,In_870,In_37);
or U646 (N_646,In_423,In_1000);
and U647 (N_647,In_1340,In_1670);
nand U648 (N_648,In_223,In_458);
and U649 (N_649,In_1209,In_893);
or U650 (N_650,In_1101,In_910);
and U651 (N_651,In_729,In_1665);
or U652 (N_652,In_1274,In_577);
and U653 (N_653,In_643,In_1536);
nor U654 (N_654,In_1686,In_1700);
nor U655 (N_655,In_619,In_602);
nand U656 (N_656,In_854,In_1314);
nand U657 (N_657,In_815,In_1914);
nand U658 (N_658,In_1315,In_323);
or U659 (N_659,In_1607,In_232);
or U660 (N_660,In_1255,In_1265);
or U661 (N_661,In_1234,In_11);
and U662 (N_662,In_1730,In_318);
nand U663 (N_663,In_176,In_1714);
or U664 (N_664,In_1429,In_39);
and U665 (N_665,In_780,In_1016);
nor U666 (N_666,In_474,In_948);
xor U667 (N_667,In_261,In_671);
and U668 (N_668,In_1508,In_1482);
nor U669 (N_669,In_148,In_644);
or U670 (N_670,In_634,In_1725);
nand U671 (N_671,In_68,In_507);
nand U672 (N_672,In_1805,In_1110);
or U673 (N_673,In_1212,In_952);
or U674 (N_674,In_483,In_229);
and U675 (N_675,In_1140,In_1795);
nand U676 (N_676,In_813,In_587);
or U677 (N_677,In_136,In_1514);
and U678 (N_678,In_739,In_139);
and U679 (N_679,In_1702,In_1884);
and U680 (N_680,In_1627,In_806);
or U681 (N_681,In_1691,In_1875);
nor U682 (N_682,In_1980,In_1652);
nand U683 (N_683,In_1560,In_1707);
or U684 (N_684,In_1199,In_1065);
or U685 (N_685,In_583,In_1695);
or U686 (N_686,In_1855,In_977);
nand U687 (N_687,In_1152,In_3);
or U688 (N_688,In_439,In_721);
nand U689 (N_689,In_822,In_817);
and U690 (N_690,In_521,In_1459);
nor U691 (N_691,In_30,In_668);
nand U692 (N_692,In_920,In_1090);
nor U693 (N_693,In_1339,In_215);
and U694 (N_694,In_460,In_885);
or U695 (N_695,In_1761,In_234);
nand U696 (N_696,In_1954,In_1503);
xnor U697 (N_697,In_542,In_757);
and U698 (N_698,In_1656,In_576);
nor U699 (N_699,In_1100,In_1123);
or U700 (N_700,In_1172,In_1963);
nor U701 (N_701,In_312,In_189);
or U702 (N_702,In_337,In_118);
nor U703 (N_703,In_1366,In_648);
or U704 (N_704,In_110,In_1660);
nor U705 (N_705,In_222,In_1942);
and U706 (N_706,In_715,In_929);
or U707 (N_707,In_187,In_1474);
or U708 (N_708,In_1532,In_1970);
and U709 (N_709,In_1384,In_212);
nor U710 (N_710,In_645,In_158);
nand U711 (N_711,In_1185,In_1380);
or U712 (N_712,In_288,In_969);
nor U713 (N_713,In_1405,In_1534);
nor U714 (N_714,In_1800,In_845);
or U715 (N_715,In_1367,In_1106);
nand U716 (N_716,In_578,In_1407);
nand U717 (N_717,In_1190,In_897);
xor U718 (N_718,In_801,In_955);
nor U719 (N_719,In_1826,In_935);
or U720 (N_720,In_36,In_1233);
nor U721 (N_721,In_1338,In_485);
or U722 (N_722,In_27,In_384);
or U723 (N_723,In_1672,In_351);
and U724 (N_724,In_1494,In_674);
nand U725 (N_725,In_1145,In_1673);
nand U726 (N_726,In_248,In_1484);
nand U727 (N_727,In_604,In_339);
and U728 (N_728,In_1013,In_1017);
nand U729 (N_729,In_1908,In_172);
and U730 (N_730,In_85,In_1174);
and U731 (N_731,In_702,In_454);
or U732 (N_732,In_883,In_1821);
nor U733 (N_733,In_596,In_1697);
and U734 (N_734,In_1118,In_538);
and U735 (N_735,In_1653,In_357);
nand U736 (N_736,In_1450,In_10);
xor U737 (N_737,In_260,In_1966);
and U738 (N_738,In_225,In_165);
and U739 (N_739,In_1135,In_1511);
and U740 (N_740,In_52,In_284);
xnor U741 (N_741,In_1726,In_32);
nor U742 (N_742,In_138,In_1196);
and U743 (N_743,In_1552,In_156);
or U744 (N_744,In_687,In_1054);
nor U745 (N_745,In_626,In_946);
and U746 (N_746,In_1667,In_1431);
or U747 (N_747,In_1741,In_1712);
or U748 (N_748,In_1747,In_258);
nand U749 (N_749,In_443,In_251);
and U750 (N_750,In_902,In_238);
and U751 (N_751,In_1684,In_1214);
nor U752 (N_752,In_1643,In_1604);
nor U753 (N_753,In_890,In_1513);
and U754 (N_754,In_344,In_1475);
or U755 (N_755,In_1891,In_692);
nand U756 (N_756,In_227,In_1285);
nor U757 (N_757,In_1720,In_1155);
and U758 (N_758,In_1188,In_112);
or U759 (N_759,In_413,In_1642);
and U760 (N_760,In_1803,In_1031);
or U761 (N_761,In_168,In_1612);
nand U762 (N_762,In_410,In_1981);
nand U763 (N_763,In_1592,In_1596);
and U764 (N_764,In_1661,In_559);
and U765 (N_765,In_1322,In_1302);
and U766 (N_766,In_1195,In_1992);
nor U767 (N_767,In_864,In_1611);
and U768 (N_768,In_1417,In_650);
or U769 (N_769,In_1075,In_1102);
nor U770 (N_770,In_19,In_498);
nor U771 (N_771,In_1733,In_939);
nor U772 (N_772,In_1144,In_1780);
or U773 (N_773,In_163,In_1692);
nand U774 (N_774,In_314,In_1649);
and U775 (N_775,In_1441,In_1854);
nor U776 (N_776,In_313,In_1835);
nor U777 (N_777,In_598,In_1990);
nor U778 (N_778,In_1907,In_1576);
nand U779 (N_779,In_1783,In_595);
nand U780 (N_780,In_868,In_1768);
and U781 (N_781,In_638,In_913);
nor U782 (N_782,In_73,In_285);
or U783 (N_783,In_571,In_40);
or U784 (N_784,In_1491,In_522);
nand U785 (N_785,In_435,In_904);
nor U786 (N_786,In_827,In_1176);
or U787 (N_787,In_87,In_1619);
or U788 (N_788,In_1527,In_487);
and U789 (N_789,In_1264,In_1605);
or U790 (N_790,In_1059,In_1786);
nand U791 (N_791,In_1488,In_83);
nor U792 (N_792,In_1899,In_1051);
nand U793 (N_793,In_1072,In_219);
nand U794 (N_794,In_762,In_1060);
or U795 (N_795,In_1651,In_1721);
nor U796 (N_796,In_1904,In_164);
and U797 (N_797,In_814,In_1674);
and U798 (N_798,In_1085,In_1303);
or U799 (N_799,In_155,In_405);
or U800 (N_800,In_14,In_601);
and U801 (N_801,In_737,In_231);
nor U802 (N_802,In_322,In_1275);
nand U803 (N_803,In_425,In_1008);
nand U804 (N_804,In_1694,In_26);
nor U805 (N_805,In_119,In_1965);
or U806 (N_806,In_1414,In_1664);
nand U807 (N_807,In_1996,In_370);
nand U808 (N_808,In_1628,In_663);
and U809 (N_809,In_759,In_917);
xor U810 (N_810,In_488,In_1754);
nand U811 (N_811,In_446,In_812);
nand U812 (N_812,In_752,In_1327);
nand U813 (N_813,In_1362,In_121);
or U814 (N_814,In_179,In_716);
nand U815 (N_815,In_5,In_1471);
and U816 (N_816,In_494,In_695);
and U817 (N_817,In_1064,In_731);
nand U818 (N_818,In_1151,In_299);
and U819 (N_819,In_1647,In_15);
xnor U820 (N_820,In_1934,In_1681);
and U821 (N_821,In_53,In_1509);
nor U822 (N_822,In_1095,In_1438);
xnor U823 (N_823,In_81,In_934);
and U824 (N_824,In_1076,In_12);
or U825 (N_825,In_924,In_167);
nor U826 (N_826,In_1179,In_962);
and U827 (N_827,In_1520,In_1357);
and U828 (N_828,In_949,In_1024);
nand U829 (N_829,In_1782,In_1350);
nor U830 (N_830,In_218,In_772);
and U831 (N_831,In_1922,In_876);
and U832 (N_832,In_455,In_1865);
and U833 (N_833,In_256,In_311);
or U834 (N_834,In_61,In_416);
or U835 (N_835,In_117,In_1435);
and U836 (N_836,In_852,In_840);
or U837 (N_837,In_1266,In_592);
nor U838 (N_838,In_1629,In_246);
nor U839 (N_839,In_162,In_516);
nor U840 (N_840,In_554,In_1290);
nor U841 (N_841,In_478,In_1858);
nand U842 (N_842,In_1126,In_675);
and U843 (N_843,In_832,In_1078);
and U844 (N_844,In_1581,In_878);
nand U845 (N_845,In_1846,In_1284);
and U846 (N_846,In_1849,In_230);
and U847 (N_847,In_152,In_1668);
nor U848 (N_848,In_1585,In_276);
nor U849 (N_849,In_1147,In_693);
nor U850 (N_850,In_1045,In_720);
nand U851 (N_851,In_740,In_1540);
or U852 (N_852,In_705,In_495);
and U853 (N_853,In_1696,In_599);
nand U854 (N_854,In_1115,In_303);
or U855 (N_855,In_771,In_611);
or U856 (N_856,In_1346,In_1258);
or U857 (N_857,In_524,In_1851);
and U858 (N_858,In_1968,In_562);
or U859 (N_859,In_1052,In_1343);
nor U860 (N_860,In_1091,In_1286);
nand U861 (N_861,In_173,In_1238);
and U862 (N_862,In_1451,In_1245);
nand U863 (N_863,In_1698,In_489);
or U864 (N_864,In_34,In_1500);
nor U865 (N_865,In_1374,In_1455);
nor U866 (N_866,In_239,In_1910);
and U867 (N_867,In_65,In_130);
nand U868 (N_868,In_1277,In_830);
nor U869 (N_869,In_387,In_1787);
nand U870 (N_870,In_1404,In_808);
nor U871 (N_871,In_1047,In_1843);
and U872 (N_872,In_651,In_1082);
or U873 (N_873,In_1828,In_632);
or U874 (N_874,In_983,In_1573);
and U875 (N_875,In_681,In_565);
and U876 (N_876,In_608,In_473);
or U877 (N_877,In_1330,In_570);
and U878 (N_878,In_1001,In_146);
or U879 (N_879,In_418,In_728);
nor U880 (N_880,In_1566,In_352);
and U881 (N_881,In_1249,In_747);
nor U882 (N_882,In_482,In_407);
nand U883 (N_883,In_670,In_190);
nor U884 (N_884,In_590,In_846);
and U885 (N_885,In_518,In_1663);
nor U886 (N_886,In_861,In_1569);
nor U887 (N_887,In_133,In_1881);
or U888 (N_888,In_1936,In_530);
nand U889 (N_889,In_1036,In_1808);
nand U890 (N_890,In_1114,In_1231);
and U891 (N_891,In_1785,In_564);
and U892 (N_892,In_2,In_1292);
and U893 (N_893,In_297,In_277);
nand U894 (N_894,In_843,In_201);
and U895 (N_895,In_1737,In_1654);
nand U896 (N_896,In_502,In_841);
and U897 (N_897,In_1678,In_959);
nand U898 (N_898,In_1601,In_289);
and U899 (N_899,In_654,In_1979);
and U900 (N_900,In_327,In_1306);
or U901 (N_901,In_532,In_287);
and U902 (N_902,In_627,In_597);
or U903 (N_903,In_1173,In_1874);
and U904 (N_904,In_746,In_958);
and U905 (N_905,In_1587,In_732);
or U906 (N_906,In_1055,In_526);
or U907 (N_907,In_1544,In_1889);
or U908 (N_908,In_1428,In_963);
nand U909 (N_909,In_803,In_1807);
and U910 (N_910,In_1555,In_1251);
nor U911 (N_911,In_264,In_1704);
nor U912 (N_912,In_183,In_1009);
nand U913 (N_913,In_1193,In_1944);
and U914 (N_914,In_652,In_607);
or U915 (N_915,In_1976,In_905);
and U916 (N_916,In_971,In_1310);
and U917 (N_917,In_208,In_325);
or U918 (N_918,In_1984,In_1603);
or U919 (N_919,In_1570,In_1824);
nor U920 (N_920,In_469,In_1012);
nor U921 (N_921,In_1639,In_1134);
or U922 (N_922,In_1792,In_395);
nor U923 (N_923,In_637,In_293);
nand U924 (N_924,In_380,In_1445);
and U925 (N_925,In_1120,In_810);
nand U926 (N_926,In_103,In_1353);
nand U927 (N_927,In_1201,In_802);
or U928 (N_928,In_221,In_1221);
nand U929 (N_929,In_1368,In_871);
or U930 (N_930,In_1002,In_240);
nand U931 (N_931,In_265,In_1900);
and U932 (N_932,In_1903,In_107);
and U933 (N_933,In_1524,In_468);
and U934 (N_934,In_1967,In_145);
nand U935 (N_935,In_1798,In_943);
nand U936 (N_936,In_696,In_1473);
nand U937 (N_937,In_1295,In_666);
nor U938 (N_938,In_689,In_45);
nand U939 (N_939,In_1943,In_1443);
nand U940 (N_940,In_1393,In_1505);
nor U941 (N_941,In_710,In_1853);
and U942 (N_942,In_1010,In_1207);
nand U943 (N_943,In_628,In_192);
nand U944 (N_944,In_1869,In_1477);
nand U945 (N_945,In_157,In_385);
or U946 (N_946,In_1974,In_879);
and U947 (N_947,In_1416,In_355);
nand U948 (N_948,In_1129,In_1280);
or U949 (N_949,In_1791,In_127);
nor U950 (N_950,In_511,In_749);
or U951 (N_951,In_1217,In_1499);
nand U952 (N_952,In_280,In_1337);
nand U953 (N_953,In_1972,In_513);
nand U954 (N_954,In_97,In_850);
nand U955 (N_955,In_389,In_1923);
nand U956 (N_956,In_1898,In_882);
nand U957 (N_957,In_1767,In_553);
and U958 (N_958,In_517,In_1203);
nand U959 (N_959,In_1940,In_1727);
nor U960 (N_960,In_1379,In_106);
and U961 (N_961,In_1841,In_1525);
xor U962 (N_962,In_686,In_1230);
or U963 (N_963,In_1300,In_1626);
and U964 (N_964,In_900,In_501);
xnor U965 (N_965,In_1061,In_1971);
and U966 (N_966,In_1760,In_691);
and U967 (N_967,In_1263,In_816);
nand U968 (N_968,In_450,In_555);
nand U969 (N_969,In_492,In_1650);
nor U970 (N_970,In_610,In_1579);
nor U971 (N_971,In_625,In_984);
and U972 (N_972,In_1282,In_669);
nand U973 (N_973,In_1175,In_875);
nand U974 (N_974,In_1412,In_31);
nand U975 (N_975,In_1997,In_1640);
or U976 (N_976,In_1360,In_862);
nor U977 (N_977,In_18,In_703);
or U978 (N_978,In_1679,In_1317);
nor U979 (N_979,In_1046,In_1487);
and U980 (N_980,In_706,In_973);
nor U981 (N_981,In_556,In_1618);
nand U982 (N_982,In_907,In_980);
and U983 (N_983,In_911,In_745);
nand U984 (N_984,In_1751,In_1239);
and U985 (N_985,In_1021,In_988);
and U986 (N_986,In_1089,In_1699);
and U987 (N_987,In_381,In_193);
and U988 (N_988,In_1150,In_1206);
or U989 (N_989,In_987,In_1034);
or U990 (N_990,In_1365,In_1352);
nor U991 (N_991,In_685,In_539);
nand U992 (N_992,In_773,In_718);
nor U993 (N_993,In_400,In_253);
and U994 (N_994,In_1018,In_1124);
or U995 (N_995,In_1464,In_711);
and U996 (N_996,In_59,In_401);
and U997 (N_997,In_1424,In_471);
or U998 (N_998,In_134,In_1467);
nor U999 (N_999,In_96,In_358);
nand U1000 (N_1000,In_362,In_1545);
or U1001 (N_1001,In_1599,In_611);
nand U1002 (N_1002,In_1376,In_29);
or U1003 (N_1003,In_1259,In_871);
and U1004 (N_1004,In_73,In_584);
or U1005 (N_1005,In_977,In_1392);
xor U1006 (N_1006,In_417,In_364);
nor U1007 (N_1007,In_491,In_1375);
xor U1008 (N_1008,In_73,In_395);
nor U1009 (N_1009,In_611,In_1277);
and U1010 (N_1010,In_1233,In_1846);
nand U1011 (N_1011,In_1400,In_287);
nand U1012 (N_1012,In_1339,In_553);
and U1013 (N_1013,In_806,In_215);
or U1014 (N_1014,In_23,In_1316);
or U1015 (N_1015,In_1113,In_585);
and U1016 (N_1016,In_813,In_455);
nand U1017 (N_1017,In_1841,In_1252);
xor U1018 (N_1018,In_1942,In_795);
or U1019 (N_1019,In_1908,In_1279);
nand U1020 (N_1020,In_1550,In_704);
nor U1021 (N_1021,In_64,In_721);
nor U1022 (N_1022,In_1317,In_1884);
nand U1023 (N_1023,In_918,In_1126);
and U1024 (N_1024,In_1858,In_893);
nor U1025 (N_1025,In_198,In_983);
or U1026 (N_1026,In_886,In_1801);
or U1027 (N_1027,In_1527,In_1137);
and U1028 (N_1028,In_626,In_1383);
and U1029 (N_1029,In_1619,In_43);
or U1030 (N_1030,In_942,In_919);
nor U1031 (N_1031,In_1093,In_998);
or U1032 (N_1032,In_64,In_1649);
nor U1033 (N_1033,In_816,In_1072);
nand U1034 (N_1034,In_295,In_1632);
and U1035 (N_1035,In_278,In_695);
or U1036 (N_1036,In_1068,In_1498);
and U1037 (N_1037,In_677,In_255);
and U1038 (N_1038,In_97,In_986);
nand U1039 (N_1039,In_601,In_146);
or U1040 (N_1040,In_1469,In_1096);
and U1041 (N_1041,In_1484,In_1866);
or U1042 (N_1042,In_1751,In_416);
or U1043 (N_1043,In_1548,In_507);
nor U1044 (N_1044,In_1917,In_172);
nor U1045 (N_1045,In_1352,In_1155);
nand U1046 (N_1046,In_383,In_920);
nand U1047 (N_1047,In_1554,In_643);
nand U1048 (N_1048,In_1798,In_1770);
nand U1049 (N_1049,In_189,In_1116);
nor U1050 (N_1050,In_1725,In_90);
and U1051 (N_1051,In_1926,In_138);
nor U1052 (N_1052,In_475,In_45);
nand U1053 (N_1053,In_425,In_23);
nand U1054 (N_1054,In_286,In_1583);
and U1055 (N_1055,In_675,In_455);
and U1056 (N_1056,In_225,In_650);
nor U1057 (N_1057,In_737,In_460);
or U1058 (N_1058,In_478,In_1760);
and U1059 (N_1059,In_539,In_1509);
and U1060 (N_1060,In_1438,In_1602);
or U1061 (N_1061,In_405,In_1900);
and U1062 (N_1062,In_1017,In_1729);
and U1063 (N_1063,In_1476,In_1262);
or U1064 (N_1064,In_669,In_1301);
nand U1065 (N_1065,In_1836,In_286);
nand U1066 (N_1066,In_1638,In_911);
xor U1067 (N_1067,In_656,In_471);
and U1068 (N_1068,In_385,In_130);
nor U1069 (N_1069,In_544,In_1074);
nand U1070 (N_1070,In_564,In_778);
nor U1071 (N_1071,In_562,In_381);
nand U1072 (N_1072,In_349,In_71);
and U1073 (N_1073,In_1607,In_70);
or U1074 (N_1074,In_794,In_987);
and U1075 (N_1075,In_95,In_576);
nand U1076 (N_1076,In_974,In_18);
and U1077 (N_1077,In_1563,In_776);
or U1078 (N_1078,In_1342,In_1860);
and U1079 (N_1079,In_1947,In_896);
nor U1080 (N_1080,In_1305,In_868);
nor U1081 (N_1081,In_1680,In_624);
and U1082 (N_1082,In_939,In_1076);
and U1083 (N_1083,In_467,In_867);
or U1084 (N_1084,In_931,In_912);
and U1085 (N_1085,In_28,In_1452);
or U1086 (N_1086,In_51,In_1811);
nand U1087 (N_1087,In_1415,In_801);
nand U1088 (N_1088,In_265,In_1311);
nand U1089 (N_1089,In_1568,In_220);
nor U1090 (N_1090,In_1507,In_1661);
or U1091 (N_1091,In_974,In_1091);
nor U1092 (N_1092,In_312,In_1065);
or U1093 (N_1093,In_792,In_1938);
nand U1094 (N_1094,In_207,In_448);
or U1095 (N_1095,In_1650,In_1199);
nand U1096 (N_1096,In_568,In_1468);
and U1097 (N_1097,In_992,In_1659);
nor U1098 (N_1098,In_840,In_935);
nand U1099 (N_1099,In_551,In_361);
or U1100 (N_1100,In_1667,In_1597);
nor U1101 (N_1101,In_1635,In_748);
and U1102 (N_1102,In_1893,In_338);
nand U1103 (N_1103,In_502,In_1143);
and U1104 (N_1104,In_1961,In_65);
nor U1105 (N_1105,In_1475,In_912);
or U1106 (N_1106,In_1198,In_358);
or U1107 (N_1107,In_684,In_1339);
or U1108 (N_1108,In_1622,In_1294);
nand U1109 (N_1109,In_20,In_189);
and U1110 (N_1110,In_103,In_975);
nand U1111 (N_1111,In_1367,In_995);
xnor U1112 (N_1112,In_1438,In_1160);
and U1113 (N_1113,In_938,In_41);
or U1114 (N_1114,In_1971,In_1034);
nand U1115 (N_1115,In_351,In_676);
nor U1116 (N_1116,In_1167,In_1779);
and U1117 (N_1117,In_1630,In_408);
and U1118 (N_1118,In_1868,In_1205);
nand U1119 (N_1119,In_1559,In_1691);
nand U1120 (N_1120,In_1681,In_1242);
and U1121 (N_1121,In_373,In_1570);
nor U1122 (N_1122,In_1849,In_1282);
nand U1123 (N_1123,In_1814,In_1576);
nor U1124 (N_1124,In_431,In_1284);
nor U1125 (N_1125,In_1610,In_1293);
nor U1126 (N_1126,In_1724,In_96);
and U1127 (N_1127,In_1566,In_297);
nor U1128 (N_1128,In_1403,In_1255);
or U1129 (N_1129,In_1749,In_1704);
and U1130 (N_1130,In_1959,In_1773);
nor U1131 (N_1131,In_767,In_17);
nor U1132 (N_1132,In_585,In_1893);
nand U1133 (N_1133,In_1953,In_391);
nand U1134 (N_1134,In_1134,In_590);
and U1135 (N_1135,In_1765,In_699);
and U1136 (N_1136,In_1532,In_915);
or U1137 (N_1137,In_1873,In_264);
and U1138 (N_1138,In_804,In_1662);
and U1139 (N_1139,In_729,In_819);
nor U1140 (N_1140,In_84,In_635);
or U1141 (N_1141,In_135,In_533);
nor U1142 (N_1142,In_1230,In_577);
and U1143 (N_1143,In_35,In_1571);
or U1144 (N_1144,In_58,In_667);
or U1145 (N_1145,In_1391,In_1840);
nor U1146 (N_1146,In_640,In_100);
nand U1147 (N_1147,In_683,In_92);
or U1148 (N_1148,In_1700,In_1820);
nand U1149 (N_1149,In_1404,In_1142);
nand U1150 (N_1150,In_1559,In_830);
or U1151 (N_1151,In_1202,In_148);
or U1152 (N_1152,In_165,In_1639);
and U1153 (N_1153,In_1347,In_1119);
nand U1154 (N_1154,In_1921,In_1344);
and U1155 (N_1155,In_354,In_933);
and U1156 (N_1156,In_1095,In_199);
or U1157 (N_1157,In_1047,In_1428);
nor U1158 (N_1158,In_730,In_1555);
nand U1159 (N_1159,In_186,In_768);
nand U1160 (N_1160,In_758,In_248);
or U1161 (N_1161,In_1608,In_15);
nor U1162 (N_1162,In_1171,In_1149);
nor U1163 (N_1163,In_1293,In_567);
nor U1164 (N_1164,In_1436,In_1997);
nor U1165 (N_1165,In_288,In_396);
or U1166 (N_1166,In_357,In_1592);
nand U1167 (N_1167,In_1472,In_583);
and U1168 (N_1168,In_637,In_236);
and U1169 (N_1169,In_421,In_1413);
nor U1170 (N_1170,In_780,In_853);
or U1171 (N_1171,In_1712,In_1346);
or U1172 (N_1172,In_747,In_1587);
nand U1173 (N_1173,In_942,In_441);
nor U1174 (N_1174,In_1395,In_1869);
and U1175 (N_1175,In_1899,In_426);
nor U1176 (N_1176,In_1506,In_229);
nor U1177 (N_1177,In_967,In_853);
nand U1178 (N_1178,In_1869,In_575);
or U1179 (N_1179,In_1387,In_497);
and U1180 (N_1180,In_1059,In_688);
nor U1181 (N_1181,In_1791,In_294);
nand U1182 (N_1182,In_1820,In_1002);
or U1183 (N_1183,In_1993,In_1531);
or U1184 (N_1184,In_818,In_316);
nand U1185 (N_1185,In_1487,In_638);
or U1186 (N_1186,In_1267,In_653);
or U1187 (N_1187,In_1561,In_705);
or U1188 (N_1188,In_1193,In_1329);
nand U1189 (N_1189,In_559,In_677);
nand U1190 (N_1190,In_1823,In_953);
nor U1191 (N_1191,In_1574,In_551);
nor U1192 (N_1192,In_1472,In_1320);
nand U1193 (N_1193,In_122,In_1128);
and U1194 (N_1194,In_1824,In_745);
nor U1195 (N_1195,In_1992,In_36);
and U1196 (N_1196,In_1805,In_1324);
or U1197 (N_1197,In_768,In_999);
and U1198 (N_1198,In_1584,In_397);
and U1199 (N_1199,In_1901,In_1330);
nor U1200 (N_1200,In_1167,In_1313);
or U1201 (N_1201,In_683,In_603);
nor U1202 (N_1202,In_1070,In_1201);
and U1203 (N_1203,In_1278,In_552);
or U1204 (N_1204,In_194,In_1842);
nor U1205 (N_1205,In_1328,In_1414);
nor U1206 (N_1206,In_1326,In_1580);
or U1207 (N_1207,In_1244,In_824);
nand U1208 (N_1208,In_1499,In_1365);
nand U1209 (N_1209,In_1404,In_233);
nand U1210 (N_1210,In_1255,In_940);
nor U1211 (N_1211,In_376,In_1208);
or U1212 (N_1212,In_374,In_1511);
nor U1213 (N_1213,In_1853,In_346);
and U1214 (N_1214,In_697,In_1489);
nand U1215 (N_1215,In_1570,In_239);
nand U1216 (N_1216,In_23,In_979);
or U1217 (N_1217,In_1434,In_590);
xnor U1218 (N_1218,In_487,In_1324);
nand U1219 (N_1219,In_134,In_151);
nand U1220 (N_1220,In_716,In_688);
nand U1221 (N_1221,In_1760,In_835);
nor U1222 (N_1222,In_69,In_512);
and U1223 (N_1223,In_1416,In_1456);
nor U1224 (N_1224,In_375,In_1404);
or U1225 (N_1225,In_472,In_1001);
or U1226 (N_1226,In_784,In_438);
nand U1227 (N_1227,In_1057,In_1049);
and U1228 (N_1228,In_1686,In_1521);
and U1229 (N_1229,In_275,In_738);
nor U1230 (N_1230,In_70,In_1173);
nand U1231 (N_1231,In_1991,In_970);
or U1232 (N_1232,In_411,In_381);
and U1233 (N_1233,In_1356,In_591);
nor U1234 (N_1234,In_1751,In_1195);
nor U1235 (N_1235,In_812,In_1178);
nand U1236 (N_1236,In_928,In_392);
or U1237 (N_1237,In_1786,In_1842);
nand U1238 (N_1238,In_805,In_1816);
nand U1239 (N_1239,In_1073,In_1537);
xor U1240 (N_1240,In_501,In_1152);
or U1241 (N_1241,In_1675,In_403);
nand U1242 (N_1242,In_1349,In_384);
nor U1243 (N_1243,In_601,In_1986);
nor U1244 (N_1244,In_768,In_1830);
or U1245 (N_1245,In_6,In_547);
nor U1246 (N_1246,In_1283,In_1079);
nand U1247 (N_1247,In_800,In_121);
nand U1248 (N_1248,In_791,In_392);
and U1249 (N_1249,In_192,In_1825);
or U1250 (N_1250,In_130,In_1381);
or U1251 (N_1251,In_834,In_477);
nand U1252 (N_1252,In_1834,In_672);
or U1253 (N_1253,In_475,In_1846);
and U1254 (N_1254,In_17,In_232);
or U1255 (N_1255,In_1548,In_1296);
and U1256 (N_1256,In_461,In_390);
nor U1257 (N_1257,In_71,In_1898);
nor U1258 (N_1258,In_1907,In_1705);
and U1259 (N_1259,In_1375,In_236);
and U1260 (N_1260,In_607,In_123);
or U1261 (N_1261,In_1192,In_1676);
nand U1262 (N_1262,In_435,In_202);
nand U1263 (N_1263,In_1292,In_472);
and U1264 (N_1264,In_1632,In_139);
or U1265 (N_1265,In_40,In_15);
and U1266 (N_1266,In_1617,In_558);
or U1267 (N_1267,In_457,In_1844);
nand U1268 (N_1268,In_1965,In_588);
or U1269 (N_1269,In_1005,In_1597);
nand U1270 (N_1270,In_1695,In_300);
or U1271 (N_1271,In_767,In_1167);
or U1272 (N_1272,In_546,In_505);
nor U1273 (N_1273,In_299,In_1521);
nand U1274 (N_1274,In_1523,In_1505);
or U1275 (N_1275,In_206,In_1295);
and U1276 (N_1276,In_255,In_718);
and U1277 (N_1277,In_1312,In_920);
and U1278 (N_1278,In_1713,In_1647);
nand U1279 (N_1279,In_1741,In_454);
nand U1280 (N_1280,In_1424,In_428);
nand U1281 (N_1281,In_1507,In_1725);
or U1282 (N_1282,In_847,In_1315);
or U1283 (N_1283,In_1853,In_58);
xor U1284 (N_1284,In_1457,In_409);
or U1285 (N_1285,In_168,In_1602);
nor U1286 (N_1286,In_221,In_571);
nand U1287 (N_1287,In_1993,In_947);
and U1288 (N_1288,In_268,In_1160);
or U1289 (N_1289,In_515,In_1580);
nand U1290 (N_1290,In_1197,In_975);
or U1291 (N_1291,In_44,In_138);
and U1292 (N_1292,In_1481,In_1330);
or U1293 (N_1293,In_1825,In_186);
and U1294 (N_1294,In_1560,In_387);
nor U1295 (N_1295,In_1931,In_12);
and U1296 (N_1296,In_1524,In_1999);
nand U1297 (N_1297,In_1532,In_482);
and U1298 (N_1298,In_1270,In_1151);
nand U1299 (N_1299,In_1564,In_1396);
or U1300 (N_1300,In_199,In_756);
or U1301 (N_1301,In_1125,In_1399);
or U1302 (N_1302,In_1049,In_191);
and U1303 (N_1303,In_421,In_697);
or U1304 (N_1304,In_1108,In_19);
nor U1305 (N_1305,In_1583,In_794);
and U1306 (N_1306,In_1155,In_846);
or U1307 (N_1307,In_1478,In_295);
and U1308 (N_1308,In_1627,In_1648);
and U1309 (N_1309,In_51,In_474);
or U1310 (N_1310,In_1312,In_129);
xnor U1311 (N_1311,In_1264,In_894);
nand U1312 (N_1312,In_1104,In_589);
or U1313 (N_1313,In_33,In_1072);
nand U1314 (N_1314,In_548,In_1993);
nor U1315 (N_1315,In_1911,In_904);
and U1316 (N_1316,In_1,In_324);
and U1317 (N_1317,In_1527,In_1971);
or U1318 (N_1318,In_1907,In_369);
and U1319 (N_1319,In_341,In_1278);
or U1320 (N_1320,In_1063,In_331);
nand U1321 (N_1321,In_1520,In_1997);
nand U1322 (N_1322,In_628,In_1253);
or U1323 (N_1323,In_197,In_1635);
nor U1324 (N_1324,In_1624,In_1805);
nor U1325 (N_1325,In_1337,In_423);
nand U1326 (N_1326,In_1074,In_1305);
nor U1327 (N_1327,In_29,In_827);
nor U1328 (N_1328,In_1935,In_1477);
or U1329 (N_1329,In_703,In_1304);
or U1330 (N_1330,In_1054,In_1899);
or U1331 (N_1331,In_576,In_1895);
nor U1332 (N_1332,In_1401,In_112);
or U1333 (N_1333,In_1489,In_241);
or U1334 (N_1334,In_1928,In_717);
nor U1335 (N_1335,In_219,In_434);
nand U1336 (N_1336,In_239,In_1937);
nor U1337 (N_1337,In_1481,In_1724);
nand U1338 (N_1338,In_797,In_478);
nand U1339 (N_1339,In_1686,In_1656);
nand U1340 (N_1340,In_1528,In_1084);
nor U1341 (N_1341,In_1319,In_872);
nor U1342 (N_1342,In_1531,In_961);
and U1343 (N_1343,In_890,In_1214);
xor U1344 (N_1344,In_1495,In_1350);
nand U1345 (N_1345,In_913,In_140);
or U1346 (N_1346,In_1521,In_1348);
and U1347 (N_1347,In_652,In_398);
nand U1348 (N_1348,In_899,In_1605);
or U1349 (N_1349,In_1592,In_1659);
or U1350 (N_1350,In_95,In_433);
and U1351 (N_1351,In_434,In_761);
or U1352 (N_1352,In_1093,In_14);
or U1353 (N_1353,In_1601,In_163);
or U1354 (N_1354,In_1415,In_143);
and U1355 (N_1355,In_1134,In_1002);
nor U1356 (N_1356,In_751,In_624);
nand U1357 (N_1357,In_1678,In_961);
or U1358 (N_1358,In_650,In_378);
or U1359 (N_1359,In_1811,In_1483);
and U1360 (N_1360,In_1768,In_856);
nand U1361 (N_1361,In_1363,In_355);
and U1362 (N_1362,In_1787,In_101);
nor U1363 (N_1363,In_17,In_1921);
nor U1364 (N_1364,In_1815,In_1531);
nand U1365 (N_1365,In_984,In_1248);
or U1366 (N_1366,In_555,In_960);
nand U1367 (N_1367,In_374,In_1773);
nand U1368 (N_1368,In_213,In_1096);
or U1369 (N_1369,In_549,In_1203);
nor U1370 (N_1370,In_1504,In_955);
nand U1371 (N_1371,In_1096,In_1812);
nor U1372 (N_1372,In_80,In_1852);
or U1373 (N_1373,In_214,In_491);
and U1374 (N_1374,In_1318,In_1970);
and U1375 (N_1375,In_1745,In_1999);
and U1376 (N_1376,In_621,In_516);
and U1377 (N_1377,In_1839,In_966);
or U1378 (N_1378,In_1060,In_440);
nand U1379 (N_1379,In_1431,In_368);
nand U1380 (N_1380,In_290,In_421);
or U1381 (N_1381,In_415,In_1650);
nand U1382 (N_1382,In_1570,In_1395);
or U1383 (N_1383,In_1005,In_249);
nor U1384 (N_1384,In_1826,In_693);
and U1385 (N_1385,In_1437,In_800);
or U1386 (N_1386,In_1231,In_1788);
nor U1387 (N_1387,In_1312,In_703);
or U1388 (N_1388,In_522,In_1397);
nand U1389 (N_1389,In_1481,In_583);
and U1390 (N_1390,In_246,In_1152);
nand U1391 (N_1391,In_1963,In_752);
and U1392 (N_1392,In_821,In_908);
or U1393 (N_1393,In_1799,In_962);
or U1394 (N_1394,In_989,In_1509);
or U1395 (N_1395,In_1006,In_297);
nor U1396 (N_1396,In_57,In_1883);
xnor U1397 (N_1397,In_229,In_1009);
nand U1398 (N_1398,In_142,In_436);
or U1399 (N_1399,In_570,In_1583);
or U1400 (N_1400,In_488,In_1259);
nor U1401 (N_1401,In_767,In_1573);
nor U1402 (N_1402,In_1113,In_1335);
nor U1403 (N_1403,In_1808,In_1674);
nand U1404 (N_1404,In_123,In_1196);
nand U1405 (N_1405,In_982,In_875);
nor U1406 (N_1406,In_60,In_884);
nor U1407 (N_1407,In_1755,In_1644);
and U1408 (N_1408,In_476,In_407);
nand U1409 (N_1409,In_1593,In_457);
nor U1410 (N_1410,In_111,In_1328);
nor U1411 (N_1411,In_1818,In_988);
and U1412 (N_1412,In_849,In_1028);
or U1413 (N_1413,In_133,In_457);
nand U1414 (N_1414,In_1522,In_478);
nor U1415 (N_1415,In_705,In_944);
nand U1416 (N_1416,In_41,In_1547);
or U1417 (N_1417,In_14,In_548);
nor U1418 (N_1418,In_82,In_533);
and U1419 (N_1419,In_312,In_1486);
nor U1420 (N_1420,In_1683,In_714);
nand U1421 (N_1421,In_1236,In_768);
and U1422 (N_1422,In_1296,In_1614);
and U1423 (N_1423,In_8,In_484);
nand U1424 (N_1424,In_1273,In_144);
nor U1425 (N_1425,In_395,In_1600);
and U1426 (N_1426,In_430,In_1003);
and U1427 (N_1427,In_1264,In_1760);
nand U1428 (N_1428,In_883,In_1537);
nor U1429 (N_1429,In_1638,In_436);
or U1430 (N_1430,In_867,In_1336);
or U1431 (N_1431,In_580,In_319);
and U1432 (N_1432,In_1250,In_1529);
and U1433 (N_1433,In_1593,In_1997);
or U1434 (N_1434,In_109,In_305);
and U1435 (N_1435,In_1611,In_81);
nor U1436 (N_1436,In_55,In_213);
and U1437 (N_1437,In_1033,In_1195);
and U1438 (N_1438,In_1384,In_1792);
and U1439 (N_1439,In_48,In_701);
nand U1440 (N_1440,In_1358,In_1333);
nand U1441 (N_1441,In_1475,In_925);
or U1442 (N_1442,In_306,In_1034);
or U1443 (N_1443,In_9,In_622);
nand U1444 (N_1444,In_297,In_1400);
nand U1445 (N_1445,In_284,In_354);
nand U1446 (N_1446,In_1272,In_487);
nand U1447 (N_1447,In_994,In_1508);
nand U1448 (N_1448,In_1945,In_952);
or U1449 (N_1449,In_1904,In_1867);
nand U1450 (N_1450,In_1894,In_488);
and U1451 (N_1451,In_735,In_1114);
and U1452 (N_1452,In_155,In_1726);
and U1453 (N_1453,In_635,In_1442);
or U1454 (N_1454,In_672,In_1300);
nor U1455 (N_1455,In_249,In_654);
nor U1456 (N_1456,In_659,In_936);
nand U1457 (N_1457,In_633,In_445);
and U1458 (N_1458,In_1576,In_1746);
or U1459 (N_1459,In_1764,In_360);
nand U1460 (N_1460,In_809,In_754);
nor U1461 (N_1461,In_1342,In_616);
and U1462 (N_1462,In_1450,In_1182);
and U1463 (N_1463,In_1101,In_640);
nand U1464 (N_1464,In_694,In_454);
nand U1465 (N_1465,In_1552,In_45);
nor U1466 (N_1466,In_695,In_361);
nand U1467 (N_1467,In_1558,In_1534);
nand U1468 (N_1468,In_983,In_451);
or U1469 (N_1469,In_1848,In_938);
nor U1470 (N_1470,In_1103,In_1858);
nand U1471 (N_1471,In_1412,In_1743);
nand U1472 (N_1472,In_950,In_1180);
and U1473 (N_1473,In_1560,In_1767);
or U1474 (N_1474,In_1949,In_71);
nor U1475 (N_1475,In_1889,In_702);
or U1476 (N_1476,In_274,In_1061);
nor U1477 (N_1477,In_677,In_1946);
or U1478 (N_1478,In_807,In_1228);
and U1479 (N_1479,In_1770,In_1882);
nand U1480 (N_1480,In_1050,In_1206);
and U1481 (N_1481,In_435,In_1618);
nor U1482 (N_1482,In_344,In_453);
and U1483 (N_1483,In_1748,In_1317);
nor U1484 (N_1484,In_1912,In_1562);
and U1485 (N_1485,In_1777,In_695);
and U1486 (N_1486,In_1382,In_958);
or U1487 (N_1487,In_1544,In_1448);
nand U1488 (N_1488,In_262,In_1348);
nand U1489 (N_1489,In_1383,In_391);
nand U1490 (N_1490,In_606,In_842);
or U1491 (N_1491,In_7,In_40);
or U1492 (N_1492,In_504,In_1756);
nand U1493 (N_1493,In_1905,In_1949);
nand U1494 (N_1494,In_343,In_1235);
and U1495 (N_1495,In_51,In_1016);
and U1496 (N_1496,In_346,In_563);
nand U1497 (N_1497,In_1362,In_1093);
and U1498 (N_1498,In_1482,In_1702);
nor U1499 (N_1499,In_909,In_1156);
or U1500 (N_1500,In_840,In_429);
nor U1501 (N_1501,In_946,In_1199);
or U1502 (N_1502,In_665,In_1561);
nand U1503 (N_1503,In_80,In_473);
nor U1504 (N_1504,In_1201,In_1864);
and U1505 (N_1505,In_728,In_1267);
and U1506 (N_1506,In_471,In_722);
nor U1507 (N_1507,In_1379,In_715);
or U1508 (N_1508,In_814,In_61);
and U1509 (N_1509,In_1333,In_284);
and U1510 (N_1510,In_1513,In_679);
or U1511 (N_1511,In_1515,In_1876);
nand U1512 (N_1512,In_1073,In_556);
and U1513 (N_1513,In_949,In_1089);
nor U1514 (N_1514,In_1726,In_921);
nand U1515 (N_1515,In_1589,In_1432);
or U1516 (N_1516,In_396,In_860);
nor U1517 (N_1517,In_399,In_532);
and U1518 (N_1518,In_761,In_665);
nand U1519 (N_1519,In_1274,In_1793);
or U1520 (N_1520,In_1197,In_1991);
nand U1521 (N_1521,In_78,In_1160);
nor U1522 (N_1522,In_246,In_350);
nor U1523 (N_1523,In_1246,In_1675);
nor U1524 (N_1524,In_728,In_1195);
nand U1525 (N_1525,In_1019,In_382);
and U1526 (N_1526,In_229,In_748);
and U1527 (N_1527,In_764,In_484);
and U1528 (N_1528,In_904,In_1719);
nor U1529 (N_1529,In_1484,In_1970);
or U1530 (N_1530,In_1968,In_1939);
nand U1531 (N_1531,In_1508,In_961);
and U1532 (N_1532,In_771,In_1704);
and U1533 (N_1533,In_255,In_1591);
nor U1534 (N_1534,In_799,In_409);
nor U1535 (N_1535,In_545,In_753);
nor U1536 (N_1536,In_547,In_492);
nand U1537 (N_1537,In_1377,In_1357);
nand U1538 (N_1538,In_1338,In_1905);
or U1539 (N_1539,In_511,In_1098);
nand U1540 (N_1540,In_689,In_1984);
nand U1541 (N_1541,In_1917,In_135);
nand U1542 (N_1542,In_216,In_573);
or U1543 (N_1543,In_358,In_887);
or U1544 (N_1544,In_743,In_1672);
nand U1545 (N_1545,In_1227,In_1162);
nand U1546 (N_1546,In_1734,In_1839);
nor U1547 (N_1547,In_1763,In_1703);
or U1548 (N_1548,In_342,In_354);
or U1549 (N_1549,In_899,In_1140);
nand U1550 (N_1550,In_1953,In_1744);
or U1551 (N_1551,In_1047,In_538);
and U1552 (N_1552,In_1965,In_587);
and U1553 (N_1553,In_252,In_671);
and U1554 (N_1554,In_1037,In_1424);
nor U1555 (N_1555,In_526,In_809);
or U1556 (N_1556,In_1741,In_759);
nor U1557 (N_1557,In_432,In_554);
nand U1558 (N_1558,In_892,In_1814);
xor U1559 (N_1559,In_528,In_653);
nand U1560 (N_1560,In_1975,In_342);
or U1561 (N_1561,In_403,In_145);
and U1562 (N_1562,In_1168,In_574);
nand U1563 (N_1563,In_587,In_1549);
or U1564 (N_1564,In_862,In_1423);
or U1565 (N_1565,In_1509,In_1236);
and U1566 (N_1566,In_1863,In_1413);
nor U1567 (N_1567,In_822,In_324);
nor U1568 (N_1568,In_511,In_773);
nor U1569 (N_1569,In_426,In_61);
nor U1570 (N_1570,In_1903,In_1337);
nor U1571 (N_1571,In_1553,In_881);
nor U1572 (N_1572,In_1470,In_51);
nand U1573 (N_1573,In_1219,In_775);
or U1574 (N_1574,In_30,In_251);
or U1575 (N_1575,In_1079,In_1420);
nor U1576 (N_1576,In_453,In_138);
nand U1577 (N_1577,In_1563,In_974);
and U1578 (N_1578,In_1814,In_272);
and U1579 (N_1579,In_1728,In_257);
and U1580 (N_1580,In_1921,In_1524);
and U1581 (N_1581,In_1282,In_704);
nand U1582 (N_1582,In_351,In_1092);
and U1583 (N_1583,In_342,In_1225);
xnor U1584 (N_1584,In_1259,In_1185);
and U1585 (N_1585,In_13,In_622);
or U1586 (N_1586,In_302,In_102);
or U1587 (N_1587,In_598,In_955);
or U1588 (N_1588,In_1691,In_695);
and U1589 (N_1589,In_658,In_1891);
and U1590 (N_1590,In_73,In_1441);
nand U1591 (N_1591,In_1389,In_1201);
nor U1592 (N_1592,In_568,In_1078);
or U1593 (N_1593,In_1503,In_682);
xnor U1594 (N_1594,In_362,In_959);
and U1595 (N_1595,In_544,In_938);
or U1596 (N_1596,In_1184,In_1088);
nor U1597 (N_1597,In_32,In_119);
and U1598 (N_1598,In_240,In_20);
nor U1599 (N_1599,In_385,In_482);
or U1600 (N_1600,In_946,In_175);
nor U1601 (N_1601,In_758,In_2);
and U1602 (N_1602,In_865,In_1105);
nor U1603 (N_1603,In_500,In_1203);
nor U1604 (N_1604,In_158,In_633);
nor U1605 (N_1605,In_1586,In_582);
or U1606 (N_1606,In_1170,In_1514);
and U1607 (N_1607,In_1683,In_135);
and U1608 (N_1608,In_398,In_1731);
or U1609 (N_1609,In_1635,In_94);
and U1610 (N_1610,In_594,In_30);
or U1611 (N_1611,In_1150,In_1686);
nor U1612 (N_1612,In_804,In_1363);
nand U1613 (N_1613,In_931,In_1977);
nor U1614 (N_1614,In_1177,In_513);
or U1615 (N_1615,In_836,In_1682);
nor U1616 (N_1616,In_1368,In_1494);
nand U1617 (N_1617,In_1809,In_343);
xnor U1618 (N_1618,In_160,In_320);
or U1619 (N_1619,In_979,In_923);
nand U1620 (N_1620,In_1031,In_1761);
nand U1621 (N_1621,In_1158,In_193);
nor U1622 (N_1622,In_1526,In_254);
or U1623 (N_1623,In_797,In_1230);
or U1624 (N_1624,In_700,In_1447);
nand U1625 (N_1625,In_1229,In_54);
nand U1626 (N_1626,In_733,In_426);
or U1627 (N_1627,In_1494,In_517);
or U1628 (N_1628,In_1691,In_1317);
or U1629 (N_1629,In_1056,In_753);
nor U1630 (N_1630,In_156,In_702);
or U1631 (N_1631,In_513,In_1644);
or U1632 (N_1632,In_1959,In_1288);
or U1633 (N_1633,In_962,In_1585);
or U1634 (N_1634,In_1522,In_591);
nand U1635 (N_1635,In_1560,In_98);
nand U1636 (N_1636,In_1475,In_1811);
nand U1637 (N_1637,In_468,In_1935);
nor U1638 (N_1638,In_884,In_1439);
nor U1639 (N_1639,In_825,In_815);
and U1640 (N_1640,In_636,In_587);
or U1641 (N_1641,In_1088,In_1952);
nand U1642 (N_1642,In_1049,In_585);
nor U1643 (N_1643,In_860,In_328);
nand U1644 (N_1644,In_1020,In_1448);
and U1645 (N_1645,In_1127,In_1643);
nand U1646 (N_1646,In_447,In_837);
or U1647 (N_1647,In_1728,In_769);
or U1648 (N_1648,In_942,In_439);
nand U1649 (N_1649,In_130,In_207);
or U1650 (N_1650,In_553,In_725);
or U1651 (N_1651,In_956,In_986);
nor U1652 (N_1652,In_945,In_104);
nand U1653 (N_1653,In_111,In_1565);
nor U1654 (N_1654,In_1799,In_339);
nor U1655 (N_1655,In_1605,In_1952);
and U1656 (N_1656,In_859,In_889);
and U1657 (N_1657,In_1967,In_471);
and U1658 (N_1658,In_644,In_1389);
nand U1659 (N_1659,In_1962,In_1995);
nand U1660 (N_1660,In_1875,In_1684);
nor U1661 (N_1661,In_180,In_53);
nor U1662 (N_1662,In_335,In_756);
nor U1663 (N_1663,In_847,In_1877);
and U1664 (N_1664,In_1644,In_1009);
and U1665 (N_1665,In_1103,In_1501);
nand U1666 (N_1666,In_1396,In_1493);
nand U1667 (N_1667,In_1957,In_1852);
or U1668 (N_1668,In_798,In_1204);
and U1669 (N_1669,In_1006,In_562);
nor U1670 (N_1670,In_279,In_1805);
nand U1671 (N_1671,In_242,In_182);
or U1672 (N_1672,In_1331,In_306);
or U1673 (N_1673,In_742,In_1775);
nand U1674 (N_1674,In_933,In_1762);
or U1675 (N_1675,In_1568,In_1974);
or U1676 (N_1676,In_111,In_1911);
and U1677 (N_1677,In_485,In_625);
nor U1678 (N_1678,In_913,In_1027);
nor U1679 (N_1679,In_1991,In_1941);
nor U1680 (N_1680,In_1889,In_584);
and U1681 (N_1681,In_1045,In_1922);
nand U1682 (N_1682,In_446,In_1271);
nor U1683 (N_1683,In_131,In_297);
nor U1684 (N_1684,In_1304,In_121);
nand U1685 (N_1685,In_379,In_851);
nand U1686 (N_1686,In_983,In_1382);
nand U1687 (N_1687,In_889,In_1279);
or U1688 (N_1688,In_162,In_649);
and U1689 (N_1689,In_718,In_115);
and U1690 (N_1690,In_346,In_633);
and U1691 (N_1691,In_620,In_1496);
or U1692 (N_1692,In_1949,In_677);
and U1693 (N_1693,In_986,In_589);
and U1694 (N_1694,In_1736,In_289);
or U1695 (N_1695,In_1961,In_1330);
nand U1696 (N_1696,In_199,In_871);
nand U1697 (N_1697,In_327,In_1599);
nor U1698 (N_1698,In_1275,In_426);
nand U1699 (N_1699,In_1080,In_1829);
xnor U1700 (N_1700,In_1337,In_699);
or U1701 (N_1701,In_1313,In_1110);
nor U1702 (N_1702,In_175,In_725);
nor U1703 (N_1703,In_1957,In_90);
nor U1704 (N_1704,In_1367,In_1180);
or U1705 (N_1705,In_1047,In_356);
nand U1706 (N_1706,In_1204,In_1312);
or U1707 (N_1707,In_1654,In_1000);
or U1708 (N_1708,In_1169,In_1315);
and U1709 (N_1709,In_1495,In_558);
and U1710 (N_1710,In_180,In_997);
nand U1711 (N_1711,In_108,In_878);
and U1712 (N_1712,In_1477,In_1124);
and U1713 (N_1713,In_166,In_1779);
nor U1714 (N_1714,In_1032,In_92);
nor U1715 (N_1715,In_1420,In_1556);
nor U1716 (N_1716,In_201,In_1297);
and U1717 (N_1717,In_1712,In_865);
and U1718 (N_1718,In_1490,In_1660);
and U1719 (N_1719,In_1253,In_1833);
nand U1720 (N_1720,In_1845,In_1218);
or U1721 (N_1721,In_1341,In_354);
nor U1722 (N_1722,In_399,In_1077);
or U1723 (N_1723,In_173,In_535);
nor U1724 (N_1724,In_1840,In_1606);
nand U1725 (N_1725,In_523,In_961);
and U1726 (N_1726,In_1901,In_1850);
and U1727 (N_1727,In_771,In_1134);
or U1728 (N_1728,In_1020,In_528);
nand U1729 (N_1729,In_134,In_807);
or U1730 (N_1730,In_958,In_376);
nand U1731 (N_1731,In_1843,In_1969);
or U1732 (N_1732,In_91,In_642);
or U1733 (N_1733,In_361,In_256);
nor U1734 (N_1734,In_560,In_411);
or U1735 (N_1735,In_321,In_478);
or U1736 (N_1736,In_191,In_1880);
or U1737 (N_1737,In_1596,In_738);
nand U1738 (N_1738,In_880,In_1119);
nor U1739 (N_1739,In_322,In_886);
or U1740 (N_1740,In_1249,In_1444);
and U1741 (N_1741,In_1666,In_1084);
or U1742 (N_1742,In_224,In_918);
and U1743 (N_1743,In_810,In_306);
nor U1744 (N_1744,In_697,In_1154);
and U1745 (N_1745,In_604,In_230);
nand U1746 (N_1746,In_430,In_667);
nor U1747 (N_1747,In_1265,In_1781);
nand U1748 (N_1748,In_1290,In_1101);
nor U1749 (N_1749,In_525,In_387);
nor U1750 (N_1750,In_1002,In_1041);
nor U1751 (N_1751,In_712,In_360);
nand U1752 (N_1752,In_141,In_1823);
nand U1753 (N_1753,In_477,In_992);
nand U1754 (N_1754,In_722,In_1627);
nand U1755 (N_1755,In_1359,In_1157);
nor U1756 (N_1756,In_1989,In_839);
nand U1757 (N_1757,In_688,In_878);
or U1758 (N_1758,In_1017,In_142);
nor U1759 (N_1759,In_309,In_254);
and U1760 (N_1760,In_1351,In_262);
and U1761 (N_1761,In_926,In_1367);
and U1762 (N_1762,In_1242,In_722);
nor U1763 (N_1763,In_1597,In_76);
and U1764 (N_1764,In_466,In_1816);
nand U1765 (N_1765,In_1487,In_1581);
or U1766 (N_1766,In_1413,In_1012);
or U1767 (N_1767,In_1861,In_946);
nand U1768 (N_1768,In_1350,In_976);
and U1769 (N_1769,In_26,In_758);
or U1770 (N_1770,In_470,In_1669);
nand U1771 (N_1771,In_1095,In_1679);
or U1772 (N_1772,In_293,In_599);
or U1773 (N_1773,In_795,In_1869);
or U1774 (N_1774,In_782,In_1523);
and U1775 (N_1775,In_1508,In_786);
nor U1776 (N_1776,In_307,In_441);
or U1777 (N_1777,In_1885,In_1692);
or U1778 (N_1778,In_875,In_321);
or U1779 (N_1779,In_1804,In_676);
or U1780 (N_1780,In_485,In_667);
or U1781 (N_1781,In_945,In_1743);
nor U1782 (N_1782,In_1695,In_1555);
nand U1783 (N_1783,In_330,In_581);
xnor U1784 (N_1784,In_421,In_1401);
nor U1785 (N_1785,In_1023,In_806);
and U1786 (N_1786,In_545,In_1426);
and U1787 (N_1787,In_1195,In_1416);
nor U1788 (N_1788,In_1940,In_1045);
and U1789 (N_1789,In_469,In_1919);
xnor U1790 (N_1790,In_1592,In_1452);
xor U1791 (N_1791,In_789,In_1428);
nor U1792 (N_1792,In_944,In_1586);
nand U1793 (N_1793,In_291,In_1078);
or U1794 (N_1794,In_1663,In_643);
or U1795 (N_1795,In_1370,In_1301);
and U1796 (N_1796,In_1301,In_1079);
nand U1797 (N_1797,In_506,In_839);
nand U1798 (N_1798,In_617,In_1307);
nor U1799 (N_1799,In_642,In_760);
or U1800 (N_1800,In_520,In_807);
and U1801 (N_1801,In_1666,In_537);
nor U1802 (N_1802,In_1842,In_1143);
nor U1803 (N_1803,In_678,In_919);
nor U1804 (N_1804,In_1916,In_1535);
and U1805 (N_1805,In_868,In_467);
nand U1806 (N_1806,In_1903,In_1116);
and U1807 (N_1807,In_436,In_1979);
or U1808 (N_1808,In_1502,In_1859);
nor U1809 (N_1809,In_814,In_1536);
or U1810 (N_1810,In_801,In_128);
and U1811 (N_1811,In_1928,In_826);
or U1812 (N_1812,In_1288,In_1077);
nand U1813 (N_1813,In_1130,In_508);
nand U1814 (N_1814,In_912,In_34);
nor U1815 (N_1815,In_711,In_440);
nand U1816 (N_1816,In_481,In_607);
nand U1817 (N_1817,In_1903,In_376);
and U1818 (N_1818,In_1603,In_1738);
and U1819 (N_1819,In_210,In_1114);
nor U1820 (N_1820,In_550,In_259);
nand U1821 (N_1821,In_1408,In_1557);
or U1822 (N_1822,In_750,In_1582);
nor U1823 (N_1823,In_961,In_1435);
xnor U1824 (N_1824,In_337,In_223);
nand U1825 (N_1825,In_72,In_1019);
or U1826 (N_1826,In_597,In_1360);
nor U1827 (N_1827,In_1946,In_352);
and U1828 (N_1828,In_1235,In_901);
and U1829 (N_1829,In_501,In_712);
nand U1830 (N_1830,In_732,In_736);
and U1831 (N_1831,In_1595,In_309);
nor U1832 (N_1832,In_814,In_1350);
nor U1833 (N_1833,In_911,In_1493);
nand U1834 (N_1834,In_881,In_1596);
and U1835 (N_1835,In_3,In_585);
nor U1836 (N_1836,In_643,In_1061);
nor U1837 (N_1837,In_453,In_1747);
nand U1838 (N_1838,In_1935,In_1432);
or U1839 (N_1839,In_1789,In_324);
or U1840 (N_1840,In_1656,In_1440);
or U1841 (N_1841,In_261,In_1631);
nor U1842 (N_1842,In_1019,In_952);
or U1843 (N_1843,In_1390,In_368);
nor U1844 (N_1844,In_1262,In_335);
and U1845 (N_1845,In_1498,In_1332);
or U1846 (N_1846,In_1155,In_1051);
nand U1847 (N_1847,In_63,In_36);
nand U1848 (N_1848,In_508,In_613);
and U1849 (N_1849,In_1737,In_4);
nor U1850 (N_1850,In_1190,In_504);
and U1851 (N_1851,In_684,In_187);
and U1852 (N_1852,In_1817,In_852);
and U1853 (N_1853,In_1528,In_309);
and U1854 (N_1854,In_1409,In_1401);
or U1855 (N_1855,In_6,In_770);
nand U1856 (N_1856,In_1214,In_1313);
nor U1857 (N_1857,In_1949,In_1933);
or U1858 (N_1858,In_1216,In_1312);
nor U1859 (N_1859,In_575,In_1161);
nor U1860 (N_1860,In_1774,In_1929);
nor U1861 (N_1861,In_1693,In_1356);
or U1862 (N_1862,In_610,In_823);
and U1863 (N_1863,In_1593,In_1025);
nand U1864 (N_1864,In_1193,In_1651);
nor U1865 (N_1865,In_345,In_991);
nor U1866 (N_1866,In_1143,In_519);
and U1867 (N_1867,In_1416,In_571);
nor U1868 (N_1868,In_284,In_1777);
or U1869 (N_1869,In_614,In_654);
and U1870 (N_1870,In_1135,In_1016);
nand U1871 (N_1871,In_683,In_149);
or U1872 (N_1872,In_277,In_1928);
nand U1873 (N_1873,In_1015,In_210);
nor U1874 (N_1874,In_592,In_301);
or U1875 (N_1875,In_1508,In_1783);
and U1876 (N_1876,In_150,In_1461);
nor U1877 (N_1877,In_1810,In_1862);
nand U1878 (N_1878,In_793,In_1859);
or U1879 (N_1879,In_65,In_454);
nand U1880 (N_1880,In_1052,In_558);
nor U1881 (N_1881,In_1104,In_1260);
nor U1882 (N_1882,In_1497,In_1035);
and U1883 (N_1883,In_839,In_1568);
nand U1884 (N_1884,In_1008,In_823);
nor U1885 (N_1885,In_894,In_860);
nand U1886 (N_1886,In_1234,In_1033);
or U1887 (N_1887,In_1516,In_512);
or U1888 (N_1888,In_156,In_6);
or U1889 (N_1889,In_182,In_851);
nand U1890 (N_1890,In_951,In_843);
or U1891 (N_1891,In_311,In_1855);
or U1892 (N_1892,In_1706,In_1076);
nand U1893 (N_1893,In_775,In_501);
nor U1894 (N_1894,In_487,In_687);
nor U1895 (N_1895,In_1319,In_453);
nor U1896 (N_1896,In_1087,In_1209);
and U1897 (N_1897,In_696,In_400);
nand U1898 (N_1898,In_1139,In_1694);
and U1899 (N_1899,In_973,In_1482);
nor U1900 (N_1900,In_117,In_1004);
or U1901 (N_1901,In_1928,In_1190);
or U1902 (N_1902,In_806,In_1832);
nor U1903 (N_1903,In_754,In_6);
or U1904 (N_1904,In_282,In_1234);
nor U1905 (N_1905,In_1518,In_389);
nor U1906 (N_1906,In_1249,In_802);
and U1907 (N_1907,In_1973,In_412);
or U1908 (N_1908,In_349,In_1022);
nand U1909 (N_1909,In_269,In_251);
or U1910 (N_1910,In_927,In_364);
nand U1911 (N_1911,In_1988,In_1318);
and U1912 (N_1912,In_1910,In_415);
and U1913 (N_1913,In_1887,In_677);
and U1914 (N_1914,In_135,In_259);
or U1915 (N_1915,In_685,In_941);
nor U1916 (N_1916,In_1430,In_1573);
nand U1917 (N_1917,In_1004,In_801);
and U1918 (N_1918,In_1599,In_1457);
nand U1919 (N_1919,In_77,In_1576);
nand U1920 (N_1920,In_1134,In_981);
and U1921 (N_1921,In_202,In_1097);
nor U1922 (N_1922,In_259,In_240);
nand U1923 (N_1923,In_1872,In_1161);
nor U1924 (N_1924,In_539,In_632);
nor U1925 (N_1925,In_1902,In_1539);
or U1926 (N_1926,In_969,In_948);
xor U1927 (N_1927,In_1168,In_1623);
and U1928 (N_1928,In_1447,In_1379);
and U1929 (N_1929,In_421,In_1381);
nor U1930 (N_1930,In_1141,In_98);
nor U1931 (N_1931,In_1333,In_1318);
nor U1932 (N_1932,In_1676,In_1315);
or U1933 (N_1933,In_888,In_1459);
nand U1934 (N_1934,In_882,In_827);
nor U1935 (N_1935,In_227,In_69);
nand U1936 (N_1936,In_389,In_7);
nand U1937 (N_1937,In_585,In_808);
nand U1938 (N_1938,In_446,In_1890);
xor U1939 (N_1939,In_619,In_1463);
nand U1940 (N_1940,In_240,In_664);
nor U1941 (N_1941,In_1864,In_513);
nor U1942 (N_1942,In_1244,In_450);
nand U1943 (N_1943,In_635,In_1086);
nor U1944 (N_1944,In_1677,In_879);
nand U1945 (N_1945,In_1592,In_1645);
nand U1946 (N_1946,In_1665,In_406);
nand U1947 (N_1947,In_1841,In_1990);
nand U1948 (N_1948,In_1388,In_1326);
nand U1949 (N_1949,In_1495,In_807);
and U1950 (N_1950,In_380,In_1349);
nor U1951 (N_1951,In_1297,In_359);
nand U1952 (N_1952,In_1448,In_40);
and U1953 (N_1953,In_92,In_692);
or U1954 (N_1954,In_1093,In_697);
and U1955 (N_1955,In_399,In_66);
or U1956 (N_1956,In_1216,In_1357);
and U1957 (N_1957,In_19,In_763);
nor U1958 (N_1958,In_426,In_632);
and U1959 (N_1959,In_401,In_284);
nand U1960 (N_1960,In_1934,In_1259);
and U1961 (N_1961,In_1484,In_1483);
or U1962 (N_1962,In_1447,In_1591);
or U1963 (N_1963,In_1622,In_527);
and U1964 (N_1964,In_1288,In_173);
or U1965 (N_1965,In_1227,In_258);
nor U1966 (N_1966,In_1197,In_1615);
and U1967 (N_1967,In_1317,In_1053);
and U1968 (N_1968,In_621,In_1272);
or U1969 (N_1969,In_264,In_1280);
and U1970 (N_1970,In_1144,In_878);
and U1971 (N_1971,In_1662,In_1926);
or U1972 (N_1972,In_165,In_1558);
nand U1973 (N_1973,In_120,In_764);
nor U1974 (N_1974,In_1144,In_1237);
and U1975 (N_1975,In_873,In_1022);
nor U1976 (N_1976,In_1349,In_1133);
nand U1977 (N_1977,In_1592,In_1523);
and U1978 (N_1978,In_1270,In_522);
and U1979 (N_1979,In_315,In_823);
nor U1980 (N_1980,In_1721,In_858);
or U1981 (N_1981,In_861,In_7);
or U1982 (N_1982,In_418,In_1159);
and U1983 (N_1983,In_790,In_1527);
and U1984 (N_1984,In_1934,In_40);
nand U1985 (N_1985,In_1484,In_1014);
and U1986 (N_1986,In_1961,In_1870);
nor U1987 (N_1987,In_257,In_1307);
nor U1988 (N_1988,In_1642,In_1758);
and U1989 (N_1989,In_388,In_1550);
xor U1990 (N_1990,In_907,In_344);
nor U1991 (N_1991,In_1013,In_1269);
nand U1992 (N_1992,In_965,In_1682);
or U1993 (N_1993,In_1706,In_1046);
nand U1994 (N_1994,In_1884,In_882);
nand U1995 (N_1995,In_1052,In_1694);
nor U1996 (N_1996,In_1829,In_984);
nand U1997 (N_1997,In_272,In_1128);
nor U1998 (N_1998,In_48,In_1939);
or U1999 (N_1999,In_1647,In_1316);
or U2000 (N_2000,In_141,In_1738);
and U2001 (N_2001,In_789,In_809);
nand U2002 (N_2002,In_1221,In_758);
or U2003 (N_2003,In_786,In_1427);
and U2004 (N_2004,In_846,In_1672);
and U2005 (N_2005,In_1663,In_819);
nand U2006 (N_2006,In_1939,In_1121);
nand U2007 (N_2007,In_402,In_383);
and U2008 (N_2008,In_1344,In_1145);
nor U2009 (N_2009,In_1620,In_695);
nand U2010 (N_2010,In_1367,In_347);
nand U2011 (N_2011,In_511,In_421);
nor U2012 (N_2012,In_895,In_896);
and U2013 (N_2013,In_1697,In_1631);
and U2014 (N_2014,In_491,In_1874);
and U2015 (N_2015,In_1236,In_830);
nor U2016 (N_2016,In_564,In_230);
nor U2017 (N_2017,In_824,In_493);
and U2018 (N_2018,In_609,In_1998);
nand U2019 (N_2019,In_745,In_765);
and U2020 (N_2020,In_1425,In_848);
or U2021 (N_2021,In_304,In_1327);
and U2022 (N_2022,In_737,In_1955);
or U2023 (N_2023,In_1467,In_246);
and U2024 (N_2024,In_735,In_625);
or U2025 (N_2025,In_408,In_640);
nand U2026 (N_2026,In_1994,In_337);
nand U2027 (N_2027,In_923,In_739);
and U2028 (N_2028,In_1008,In_38);
nor U2029 (N_2029,In_1603,In_701);
or U2030 (N_2030,In_1285,In_512);
and U2031 (N_2031,In_1874,In_1267);
nand U2032 (N_2032,In_529,In_1870);
or U2033 (N_2033,In_1714,In_1349);
or U2034 (N_2034,In_1623,In_951);
nand U2035 (N_2035,In_1007,In_1190);
or U2036 (N_2036,In_888,In_1632);
nor U2037 (N_2037,In_698,In_1554);
nand U2038 (N_2038,In_916,In_845);
and U2039 (N_2039,In_1615,In_646);
or U2040 (N_2040,In_156,In_658);
and U2041 (N_2041,In_1576,In_1430);
or U2042 (N_2042,In_275,In_195);
and U2043 (N_2043,In_202,In_62);
and U2044 (N_2044,In_136,In_1593);
or U2045 (N_2045,In_287,In_858);
nor U2046 (N_2046,In_1497,In_1742);
or U2047 (N_2047,In_108,In_1362);
and U2048 (N_2048,In_477,In_1830);
or U2049 (N_2049,In_613,In_1651);
nor U2050 (N_2050,In_856,In_960);
and U2051 (N_2051,In_971,In_1757);
nand U2052 (N_2052,In_1145,In_759);
nand U2053 (N_2053,In_1338,In_1162);
nor U2054 (N_2054,In_148,In_1567);
and U2055 (N_2055,In_1963,In_424);
nor U2056 (N_2056,In_1095,In_1349);
and U2057 (N_2057,In_706,In_1412);
or U2058 (N_2058,In_442,In_200);
nand U2059 (N_2059,In_1234,In_796);
nor U2060 (N_2060,In_1476,In_1666);
nand U2061 (N_2061,In_522,In_1765);
or U2062 (N_2062,In_1535,In_1850);
and U2063 (N_2063,In_44,In_831);
nand U2064 (N_2064,In_279,In_1098);
and U2065 (N_2065,In_1492,In_1948);
or U2066 (N_2066,In_1918,In_47);
nand U2067 (N_2067,In_405,In_1955);
nand U2068 (N_2068,In_1320,In_1270);
or U2069 (N_2069,In_1038,In_1226);
and U2070 (N_2070,In_68,In_1306);
or U2071 (N_2071,In_1890,In_304);
nand U2072 (N_2072,In_894,In_1203);
and U2073 (N_2073,In_1766,In_1412);
and U2074 (N_2074,In_131,In_394);
nor U2075 (N_2075,In_2,In_796);
nand U2076 (N_2076,In_1142,In_1991);
or U2077 (N_2077,In_827,In_1203);
and U2078 (N_2078,In_1280,In_1344);
and U2079 (N_2079,In_1815,In_1544);
or U2080 (N_2080,In_1373,In_1848);
or U2081 (N_2081,In_1113,In_665);
nand U2082 (N_2082,In_1495,In_673);
and U2083 (N_2083,In_1904,In_1595);
or U2084 (N_2084,In_1273,In_1002);
nor U2085 (N_2085,In_1751,In_138);
nor U2086 (N_2086,In_1638,In_479);
nand U2087 (N_2087,In_1287,In_1927);
nand U2088 (N_2088,In_285,In_1706);
xnor U2089 (N_2089,In_1310,In_1048);
nand U2090 (N_2090,In_418,In_1485);
or U2091 (N_2091,In_565,In_421);
nor U2092 (N_2092,In_1589,In_508);
and U2093 (N_2093,In_1066,In_1581);
and U2094 (N_2094,In_10,In_1798);
xor U2095 (N_2095,In_528,In_773);
nor U2096 (N_2096,In_706,In_726);
nor U2097 (N_2097,In_1076,In_1140);
nand U2098 (N_2098,In_1123,In_518);
and U2099 (N_2099,In_1712,In_695);
or U2100 (N_2100,In_1857,In_1867);
and U2101 (N_2101,In_1436,In_1783);
and U2102 (N_2102,In_842,In_1415);
nand U2103 (N_2103,In_98,In_1194);
nand U2104 (N_2104,In_713,In_346);
or U2105 (N_2105,In_1517,In_1919);
and U2106 (N_2106,In_354,In_1433);
nand U2107 (N_2107,In_991,In_1167);
xor U2108 (N_2108,In_1557,In_1204);
nand U2109 (N_2109,In_1774,In_1832);
nand U2110 (N_2110,In_624,In_850);
nor U2111 (N_2111,In_1786,In_1165);
or U2112 (N_2112,In_590,In_1017);
nor U2113 (N_2113,In_323,In_18);
and U2114 (N_2114,In_1958,In_1475);
nand U2115 (N_2115,In_790,In_506);
and U2116 (N_2116,In_545,In_566);
and U2117 (N_2117,In_315,In_653);
and U2118 (N_2118,In_1167,In_1949);
and U2119 (N_2119,In_1685,In_1232);
and U2120 (N_2120,In_245,In_232);
or U2121 (N_2121,In_1647,In_1655);
or U2122 (N_2122,In_43,In_738);
nor U2123 (N_2123,In_959,In_1162);
nor U2124 (N_2124,In_1945,In_714);
or U2125 (N_2125,In_80,In_1667);
or U2126 (N_2126,In_1480,In_1688);
nand U2127 (N_2127,In_947,In_152);
nor U2128 (N_2128,In_28,In_1450);
nand U2129 (N_2129,In_966,In_967);
and U2130 (N_2130,In_1193,In_124);
nand U2131 (N_2131,In_1856,In_1928);
and U2132 (N_2132,In_1484,In_1139);
nor U2133 (N_2133,In_216,In_873);
or U2134 (N_2134,In_982,In_1003);
nor U2135 (N_2135,In_1520,In_1726);
and U2136 (N_2136,In_1064,In_293);
and U2137 (N_2137,In_1219,In_1021);
and U2138 (N_2138,In_1379,In_264);
nor U2139 (N_2139,In_498,In_215);
nor U2140 (N_2140,In_594,In_1744);
nor U2141 (N_2141,In_941,In_495);
nand U2142 (N_2142,In_94,In_1885);
nand U2143 (N_2143,In_180,In_1285);
and U2144 (N_2144,In_1715,In_1827);
and U2145 (N_2145,In_762,In_1139);
nor U2146 (N_2146,In_558,In_1070);
and U2147 (N_2147,In_605,In_1613);
nand U2148 (N_2148,In_1042,In_388);
nor U2149 (N_2149,In_1019,In_644);
and U2150 (N_2150,In_797,In_414);
nor U2151 (N_2151,In_109,In_960);
nand U2152 (N_2152,In_362,In_413);
nor U2153 (N_2153,In_196,In_1963);
nand U2154 (N_2154,In_1788,In_895);
nor U2155 (N_2155,In_722,In_1784);
xor U2156 (N_2156,In_526,In_1624);
or U2157 (N_2157,In_1551,In_71);
and U2158 (N_2158,In_1003,In_853);
nor U2159 (N_2159,In_643,In_961);
nand U2160 (N_2160,In_102,In_1852);
nand U2161 (N_2161,In_1425,In_1597);
nor U2162 (N_2162,In_1503,In_954);
and U2163 (N_2163,In_910,In_1401);
and U2164 (N_2164,In_731,In_252);
and U2165 (N_2165,In_188,In_560);
or U2166 (N_2166,In_1366,In_832);
nand U2167 (N_2167,In_1558,In_1783);
or U2168 (N_2168,In_1856,In_1723);
and U2169 (N_2169,In_1120,In_559);
nand U2170 (N_2170,In_935,In_1939);
nor U2171 (N_2171,In_1896,In_102);
xnor U2172 (N_2172,In_1719,In_1538);
nor U2173 (N_2173,In_419,In_1638);
nor U2174 (N_2174,In_1690,In_245);
nor U2175 (N_2175,In_1314,In_395);
or U2176 (N_2176,In_726,In_126);
nand U2177 (N_2177,In_700,In_1594);
nand U2178 (N_2178,In_290,In_786);
or U2179 (N_2179,In_124,In_1898);
or U2180 (N_2180,In_370,In_135);
or U2181 (N_2181,In_966,In_1816);
nand U2182 (N_2182,In_1726,In_703);
or U2183 (N_2183,In_1351,In_1024);
and U2184 (N_2184,In_877,In_1744);
and U2185 (N_2185,In_1328,In_1771);
nand U2186 (N_2186,In_420,In_1653);
and U2187 (N_2187,In_1189,In_460);
or U2188 (N_2188,In_663,In_1243);
or U2189 (N_2189,In_1813,In_938);
nor U2190 (N_2190,In_873,In_487);
nand U2191 (N_2191,In_302,In_1544);
nor U2192 (N_2192,In_1876,In_1392);
nor U2193 (N_2193,In_235,In_209);
or U2194 (N_2194,In_978,In_790);
nor U2195 (N_2195,In_771,In_280);
nand U2196 (N_2196,In_258,In_1236);
nand U2197 (N_2197,In_66,In_878);
nand U2198 (N_2198,In_568,In_1597);
and U2199 (N_2199,In_1980,In_1496);
and U2200 (N_2200,In_1200,In_214);
or U2201 (N_2201,In_1410,In_824);
or U2202 (N_2202,In_1968,In_575);
nor U2203 (N_2203,In_1400,In_1563);
and U2204 (N_2204,In_1043,In_1241);
or U2205 (N_2205,In_43,In_1355);
nor U2206 (N_2206,In_373,In_912);
or U2207 (N_2207,In_1562,In_1775);
nor U2208 (N_2208,In_148,In_1260);
nand U2209 (N_2209,In_1035,In_1091);
or U2210 (N_2210,In_1683,In_487);
nand U2211 (N_2211,In_1381,In_1543);
and U2212 (N_2212,In_786,In_1177);
and U2213 (N_2213,In_1969,In_175);
nor U2214 (N_2214,In_369,In_401);
and U2215 (N_2215,In_292,In_1630);
nor U2216 (N_2216,In_1192,In_1948);
nand U2217 (N_2217,In_1366,In_814);
or U2218 (N_2218,In_1112,In_1603);
or U2219 (N_2219,In_40,In_896);
or U2220 (N_2220,In_496,In_1158);
or U2221 (N_2221,In_775,In_1171);
and U2222 (N_2222,In_134,In_680);
nor U2223 (N_2223,In_321,In_1440);
nor U2224 (N_2224,In_869,In_161);
nor U2225 (N_2225,In_1974,In_1689);
and U2226 (N_2226,In_1604,In_210);
nor U2227 (N_2227,In_1276,In_1972);
and U2228 (N_2228,In_553,In_483);
nand U2229 (N_2229,In_350,In_670);
nand U2230 (N_2230,In_1070,In_1925);
nand U2231 (N_2231,In_1039,In_710);
nor U2232 (N_2232,In_1776,In_927);
nor U2233 (N_2233,In_1276,In_1139);
nand U2234 (N_2234,In_261,In_1441);
nor U2235 (N_2235,In_929,In_1976);
nand U2236 (N_2236,In_1805,In_216);
or U2237 (N_2237,In_143,In_1755);
nor U2238 (N_2238,In_1342,In_648);
and U2239 (N_2239,In_1153,In_174);
nor U2240 (N_2240,In_827,In_1961);
nor U2241 (N_2241,In_810,In_1636);
or U2242 (N_2242,In_1517,In_865);
or U2243 (N_2243,In_1629,In_1592);
nor U2244 (N_2244,In_546,In_1811);
nor U2245 (N_2245,In_1381,In_1304);
or U2246 (N_2246,In_60,In_1482);
or U2247 (N_2247,In_1797,In_1066);
and U2248 (N_2248,In_1550,In_0);
nand U2249 (N_2249,In_1442,In_1507);
or U2250 (N_2250,In_1168,In_1166);
or U2251 (N_2251,In_929,In_1966);
nor U2252 (N_2252,In_411,In_1265);
nand U2253 (N_2253,In_1698,In_1312);
and U2254 (N_2254,In_1566,In_936);
nand U2255 (N_2255,In_357,In_538);
nor U2256 (N_2256,In_728,In_1791);
and U2257 (N_2257,In_1780,In_1554);
or U2258 (N_2258,In_1081,In_271);
or U2259 (N_2259,In_302,In_1593);
or U2260 (N_2260,In_339,In_1556);
and U2261 (N_2261,In_1433,In_457);
and U2262 (N_2262,In_1341,In_1826);
or U2263 (N_2263,In_1492,In_1450);
or U2264 (N_2264,In_1346,In_880);
or U2265 (N_2265,In_113,In_1449);
and U2266 (N_2266,In_87,In_994);
and U2267 (N_2267,In_533,In_432);
nor U2268 (N_2268,In_1190,In_651);
and U2269 (N_2269,In_1874,In_1575);
nor U2270 (N_2270,In_415,In_1536);
and U2271 (N_2271,In_1812,In_154);
nand U2272 (N_2272,In_1521,In_144);
and U2273 (N_2273,In_368,In_1801);
and U2274 (N_2274,In_1805,In_28);
nand U2275 (N_2275,In_806,In_1586);
and U2276 (N_2276,In_202,In_198);
nor U2277 (N_2277,In_1643,In_1828);
nand U2278 (N_2278,In_1315,In_1955);
or U2279 (N_2279,In_348,In_179);
and U2280 (N_2280,In_1381,In_1669);
and U2281 (N_2281,In_796,In_1110);
and U2282 (N_2282,In_531,In_804);
or U2283 (N_2283,In_1555,In_1608);
xor U2284 (N_2284,In_905,In_566);
nor U2285 (N_2285,In_360,In_1938);
and U2286 (N_2286,In_1769,In_370);
nor U2287 (N_2287,In_363,In_263);
and U2288 (N_2288,In_1918,In_581);
nand U2289 (N_2289,In_331,In_1461);
or U2290 (N_2290,In_1863,In_1359);
and U2291 (N_2291,In_799,In_65);
or U2292 (N_2292,In_992,In_1067);
nor U2293 (N_2293,In_730,In_1840);
nand U2294 (N_2294,In_464,In_324);
xnor U2295 (N_2295,In_1115,In_1349);
nand U2296 (N_2296,In_9,In_1845);
nand U2297 (N_2297,In_1395,In_725);
and U2298 (N_2298,In_1914,In_392);
and U2299 (N_2299,In_322,In_514);
or U2300 (N_2300,In_862,In_1527);
nor U2301 (N_2301,In_1282,In_1719);
or U2302 (N_2302,In_1646,In_1029);
nand U2303 (N_2303,In_444,In_203);
nand U2304 (N_2304,In_562,In_1064);
nand U2305 (N_2305,In_1059,In_1459);
nor U2306 (N_2306,In_1345,In_101);
or U2307 (N_2307,In_1342,In_132);
nor U2308 (N_2308,In_1614,In_1131);
nand U2309 (N_2309,In_1559,In_925);
nor U2310 (N_2310,In_1920,In_20);
nor U2311 (N_2311,In_1817,In_313);
and U2312 (N_2312,In_1959,In_1650);
and U2313 (N_2313,In_1495,In_1772);
nand U2314 (N_2314,In_1038,In_203);
nand U2315 (N_2315,In_436,In_891);
nand U2316 (N_2316,In_223,In_440);
nand U2317 (N_2317,In_1376,In_1411);
nand U2318 (N_2318,In_707,In_1108);
xor U2319 (N_2319,In_460,In_1699);
and U2320 (N_2320,In_920,In_1493);
nor U2321 (N_2321,In_494,In_923);
and U2322 (N_2322,In_1788,In_1371);
nor U2323 (N_2323,In_1528,In_813);
or U2324 (N_2324,In_1119,In_1156);
nor U2325 (N_2325,In_1422,In_1461);
or U2326 (N_2326,In_904,In_251);
nor U2327 (N_2327,In_1006,In_503);
nand U2328 (N_2328,In_166,In_102);
and U2329 (N_2329,In_1943,In_661);
or U2330 (N_2330,In_731,In_1177);
nor U2331 (N_2331,In_901,In_1158);
or U2332 (N_2332,In_16,In_216);
nor U2333 (N_2333,In_1275,In_24);
and U2334 (N_2334,In_583,In_11);
nand U2335 (N_2335,In_678,In_299);
nand U2336 (N_2336,In_1960,In_761);
nand U2337 (N_2337,In_301,In_1846);
nor U2338 (N_2338,In_1214,In_1831);
nor U2339 (N_2339,In_1609,In_1999);
nand U2340 (N_2340,In_1519,In_742);
and U2341 (N_2341,In_503,In_459);
nand U2342 (N_2342,In_1180,In_1255);
or U2343 (N_2343,In_1173,In_362);
nand U2344 (N_2344,In_774,In_1154);
nand U2345 (N_2345,In_133,In_1703);
or U2346 (N_2346,In_1090,In_134);
or U2347 (N_2347,In_548,In_1651);
nor U2348 (N_2348,In_394,In_196);
and U2349 (N_2349,In_1914,In_757);
or U2350 (N_2350,In_537,In_1843);
or U2351 (N_2351,In_318,In_1992);
or U2352 (N_2352,In_206,In_307);
nand U2353 (N_2353,In_1870,In_93);
nor U2354 (N_2354,In_1334,In_603);
and U2355 (N_2355,In_1828,In_85);
nor U2356 (N_2356,In_1096,In_1602);
and U2357 (N_2357,In_736,In_179);
nand U2358 (N_2358,In_663,In_1357);
or U2359 (N_2359,In_1284,In_1787);
nand U2360 (N_2360,In_593,In_1129);
and U2361 (N_2361,In_711,In_398);
and U2362 (N_2362,In_1640,In_1131);
or U2363 (N_2363,In_1747,In_985);
and U2364 (N_2364,In_1976,In_105);
nand U2365 (N_2365,In_1840,In_460);
nor U2366 (N_2366,In_538,In_1834);
nand U2367 (N_2367,In_368,In_584);
nand U2368 (N_2368,In_73,In_1947);
and U2369 (N_2369,In_1110,In_338);
or U2370 (N_2370,In_1647,In_643);
and U2371 (N_2371,In_1392,In_98);
nor U2372 (N_2372,In_43,In_1474);
or U2373 (N_2373,In_1310,In_1507);
nor U2374 (N_2374,In_934,In_327);
and U2375 (N_2375,In_212,In_761);
or U2376 (N_2376,In_273,In_1258);
nand U2377 (N_2377,In_141,In_1890);
nor U2378 (N_2378,In_1851,In_917);
nand U2379 (N_2379,In_252,In_166);
or U2380 (N_2380,In_1914,In_1100);
nor U2381 (N_2381,In_1794,In_686);
or U2382 (N_2382,In_180,In_1953);
or U2383 (N_2383,In_1973,In_1890);
nor U2384 (N_2384,In_1543,In_400);
or U2385 (N_2385,In_368,In_663);
or U2386 (N_2386,In_856,In_1054);
or U2387 (N_2387,In_1930,In_735);
nor U2388 (N_2388,In_1230,In_1159);
nor U2389 (N_2389,In_1725,In_1316);
and U2390 (N_2390,In_977,In_1096);
or U2391 (N_2391,In_321,In_479);
and U2392 (N_2392,In_1687,In_562);
nand U2393 (N_2393,In_1447,In_886);
and U2394 (N_2394,In_1872,In_335);
or U2395 (N_2395,In_768,In_49);
nor U2396 (N_2396,In_635,In_102);
and U2397 (N_2397,In_831,In_972);
nor U2398 (N_2398,In_1501,In_1079);
or U2399 (N_2399,In_751,In_437);
and U2400 (N_2400,In_1633,In_548);
and U2401 (N_2401,In_284,In_1954);
nand U2402 (N_2402,In_1789,In_151);
nor U2403 (N_2403,In_34,In_930);
or U2404 (N_2404,In_455,In_1557);
nand U2405 (N_2405,In_694,In_1838);
nand U2406 (N_2406,In_1839,In_1585);
nand U2407 (N_2407,In_90,In_1765);
nand U2408 (N_2408,In_1198,In_1837);
nand U2409 (N_2409,In_377,In_566);
nand U2410 (N_2410,In_1734,In_574);
nand U2411 (N_2411,In_1540,In_1118);
and U2412 (N_2412,In_1435,In_1958);
nand U2413 (N_2413,In_1692,In_840);
nor U2414 (N_2414,In_295,In_1525);
nand U2415 (N_2415,In_193,In_330);
nor U2416 (N_2416,In_951,In_1728);
or U2417 (N_2417,In_240,In_475);
and U2418 (N_2418,In_73,In_1335);
nand U2419 (N_2419,In_1111,In_1863);
nor U2420 (N_2420,In_218,In_955);
and U2421 (N_2421,In_1797,In_1479);
nor U2422 (N_2422,In_1164,In_1918);
nor U2423 (N_2423,In_1325,In_943);
nor U2424 (N_2424,In_957,In_742);
or U2425 (N_2425,In_1319,In_891);
and U2426 (N_2426,In_1260,In_1712);
or U2427 (N_2427,In_559,In_737);
nor U2428 (N_2428,In_10,In_1050);
or U2429 (N_2429,In_1608,In_619);
or U2430 (N_2430,In_1521,In_1299);
and U2431 (N_2431,In_728,In_568);
or U2432 (N_2432,In_1478,In_1225);
nor U2433 (N_2433,In_929,In_1201);
or U2434 (N_2434,In_1935,In_1335);
and U2435 (N_2435,In_851,In_822);
or U2436 (N_2436,In_705,In_277);
nor U2437 (N_2437,In_902,In_1442);
or U2438 (N_2438,In_172,In_632);
nand U2439 (N_2439,In_1070,In_1185);
nor U2440 (N_2440,In_868,In_927);
nor U2441 (N_2441,In_1256,In_1972);
and U2442 (N_2442,In_1009,In_1591);
xnor U2443 (N_2443,In_1118,In_3);
nor U2444 (N_2444,In_1999,In_1476);
or U2445 (N_2445,In_1155,In_751);
or U2446 (N_2446,In_1333,In_1566);
and U2447 (N_2447,In_256,In_1247);
and U2448 (N_2448,In_1399,In_775);
nand U2449 (N_2449,In_1871,In_1150);
and U2450 (N_2450,In_2,In_1359);
nand U2451 (N_2451,In_592,In_1526);
or U2452 (N_2452,In_1505,In_1686);
or U2453 (N_2453,In_1174,In_1008);
and U2454 (N_2454,In_394,In_949);
or U2455 (N_2455,In_1099,In_1438);
nand U2456 (N_2456,In_1611,In_441);
and U2457 (N_2457,In_992,In_355);
or U2458 (N_2458,In_1488,In_738);
nand U2459 (N_2459,In_1299,In_679);
nand U2460 (N_2460,In_1284,In_1600);
nand U2461 (N_2461,In_823,In_1926);
nor U2462 (N_2462,In_564,In_360);
and U2463 (N_2463,In_806,In_45);
and U2464 (N_2464,In_1464,In_230);
or U2465 (N_2465,In_717,In_1561);
and U2466 (N_2466,In_42,In_1073);
nand U2467 (N_2467,In_1628,In_961);
nand U2468 (N_2468,In_891,In_979);
and U2469 (N_2469,In_819,In_1733);
or U2470 (N_2470,In_527,In_1692);
and U2471 (N_2471,In_1372,In_1597);
nor U2472 (N_2472,In_1849,In_1403);
nor U2473 (N_2473,In_1932,In_826);
or U2474 (N_2474,In_1854,In_1114);
nand U2475 (N_2475,In_13,In_904);
and U2476 (N_2476,In_1196,In_112);
nand U2477 (N_2477,In_1909,In_292);
or U2478 (N_2478,In_103,In_581);
nor U2479 (N_2479,In_1274,In_303);
nand U2480 (N_2480,In_1388,In_970);
and U2481 (N_2481,In_203,In_1067);
nor U2482 (N_2482,In_1796,In_773);
and U2483 (N_2483,In_379,In_1295);
and U2484 (N_2484,In_697,In_1677);
nor U2485 (N_2485,In_415,In_496);
or U2486 (N_2486,In_1265,In_758);
or U2487 (N_2487,In_1283,In_1148);
and U2488 (N_2488,In_1995,In_1606);
nand U2489 (N_2489,In_236,In_1939);
and U2490 (N_2490,In_537,In_1793);
or U2491 (N_2491,In_202,In_525);
and U2492 (N_2492,In_1901,In_50);
and U2493 (N_2493,In_1987,In_549);
nand U2494 (N_2494,In_579,In_1883);
nor U2495 (N_2495,In_208,In_1687);
and U2496 (N_2496,In_111,In_1713);
nor U2497 (N_2497,In_1245,In_1846);
nand U2498 (N_2498,In_380,In_1609);
or U2499 (N_2499,In_1146,In_702);
or U2500 (N_2500,In_309,In_974);
nand U2501 (N_2501,In_1133,In_545);
nor U2502 (N_2502,In_1442,In_1896);
and U2503 (N_2503,In_1687,In_119);
or U2504 (N_2504,In_1742,In_755);
xnor U2505 (N_2505,In_1529,In_780);
and U2506 (N_2506,In_1696,In_226);
nand U2507 (N_2507,In_1457,In_140);
or U2508 (N_2508,In_1253,In_181);
nand U2509 (N_2509,In_1460,In_190);
and U2510 (N_2510,In_1956,In_785);
or U2511 (N_2511,In_551,In_1697);
and U2512 (N_2512,In_1389,In_971);
or U2513 (N_2513,In_762,In_1051);
or U2514 (N_2514,In_764,In_68);
and U2515 (N_2515,In_555,In_1818);
and U2516 (N_2516,In_353,In_1346);
nor U2517 (N_2517,In_630,In_1082);
nor U2518 (N_2518,In_1283,In_375);
nor U2519 (N_2519,In_1051,In_1426);
or U2520 (N_2520,In_811,In_273);
nand U2521 (N_2521,In_1289,In_369);
or U2522 (N_2522,In_1385,In_630);
nor U2523 (N_2523,In_401,In_1366);
or U2524 (N_2524,In_1477,In_102);
and U2525 (N_2525,In_474,In_325);
nor U2526 (N_2526,In_38,In_1530);
and U2527 (N_2527,In_1951,In_1489);
and U2528 (N_2528,In_458,In_8);
and U2529 (N_2529,In_1336,In_1741);
or U2530 (N_2530,In_763,In_1759);
or U2531 (N_2531,In_1838,In_126);
nand U2532 (N_2532,In_1194,In_179);
nand U2533 (N_2533,In_732,In_1409);
and U2534 (N_2534,In_670,In_789);
nand U2535 (N_2535,In_1586,In_846);
and U2536 (N_2536,In_1440,In_342);
or U2537 (N_2537,In_1994,In_1171);
or U2538 (N_2538,In_155,In_578);
or U2539 (N_2539,In_129,In_815);
nand U2540 (N_2540,In_649,In_929);
or U2541 (N_2541,In_1341,In_1307);
or U2542 (N_2542,In_292,In_1412);
nor U2543 (N_2543,In_1465,In_633);
nand U2544 (N_2544,In_639,In_1620);
nand U2545 (N_2545,In_1600,In_184);
and U2546 (N_2546,In_1966,In_891);
or U2547 (N_2547,In_133,In_958);
and U2548 (N_2548,In_185,In_1163);
nor U2549 (N_2549,In_64,In_1634);
and U2550 (N_2550,In_521,In_1087);
nand U2551 (N_2551,In_75,In_534);
or U2552 (N_2552,In_1186,In_1162);
nand U2553 (N_2553,In_1702,In_1791);
nand U2554 (N_2554,In_803,In_1052);
nand U2555 (N_2555,In_1451,In_1114);
or U2556 (N_2556,In_1301,In_776);
and U2557 (N_2557,In_1647,In_143);
nor U2558 (N_2558,In_224,In_505);
nand U2559 (N_2559,In_739,In_1341);
and U2560 (N_2560,In_1677,In_1292);
nand U2561 (N_2561,In_703,In_548);
nand U2562 (N_2562,In_443,In_573);
and U2563 (N_2563,In_32,In_1421);
xnor U2564 (N_2564,In_1213,In_727);
nor U2565 (N_2565,In_1206,In_1119);
or U2566 (N_2566,In_1350,In_1773);
or U2567 (N_2567,In_1343,In_1728);
and U2568 (N_2568,In_158,In_576);
nand U2569 (N_2569,In_1495,In_736);
nor U2570 (N_2570,In_760,In_883);
or U2571 (N_2571,In_232,In_552);
or U2572 (N_2572,In_308,In_1080);
xor U2573 (N_2573,In_716,In_91);
nand U2574 (N_2574,In_1593,In_1137);
and U2575 (N_2575,In_1294,In_1585);
or U2576 (N_2576,In_744,In_1734);
or U2577 (N_2577,In_1250,In_1219);
or U2578 (N_2578,In_1569,In_12);
nor U2579 (N_2579,In_894,In_839);
nand U2580 (N_2580,In_158,In_1473);
nand U2581 (N_2581,In_313,In_1688);
and U2582 (N_2582,In_1350,In_1186);
nand U2583 (N_2583,In_376,In_601);
and U2584 (N_2584,In_91,In_1488);
nand U2585 (N_2585,In_1453,In_655);
nand U2586 (N_2586,In_1701,In_190);
and U2587 (N_2587,In_1622,In_59);
nand U2588 (N_2588,In_916,In_1020);
or U2589 (N_2589,In_1085,In_600);
nand U2590 (N_2590,In_275,In_353);
nor U2591 (N_2591,In_574,In_835);
or U2592 (N_2592,In_1528,In_496);
and U2593 (N_2593,In_450,In_536);
nor U2594 (N_2594,In_423,In_1405);
and U2595 (N_2595,In_203,In_1977);
xor U2596 (N_2596,In_1278,In_1550);
or U2597 (N_2597,In_1156,In_885);
nand U2598 (N_2598,In_1542,In_1765);
and U2599 (N_2599,In_1531,In_451);
and U2600 (N_2600,In_1515,In_1007);
nor U2601 (N_2601,In_103,In_81);
and U2602 (N_2602,In_1824,In_1032);
and U2603 (N_2603,In_1822,In_31);
or U2604 (N_2604,In_593,In_18);
or U2605 (N_2605,In_1886,In_1033);
and U2606 (N_2606,In_678,In_740);
and U2607 (N_2607,In_1943,In_1022);
or U2608 (N_2608,In_667,In_1134);
and U2609 (N_2609,In_1779,In_1000);
and U2610 (N_2610,In_1597,In_1684);
and U2611 (N_2611,In_1146,In_1989);
and U2612 (N_2612,In_547,In_1125);
and U2613 (N_2613,In_409,In_1332);
nand U2614 (N_2614,In_1776,In_1495);
or U2615 (N_2615,In_261,In_1219);
nor U2616 (N_2616,In_1637,In_714);
nor U2617 (N_2617,In_702,In_887);
nand U2618 (N_2618,In_1765,In_515);
nand U2619 (N_2619,In_178,In_1930);
and U2620 (N_2620,In_1259,In_1301);
or U2621 (N_2621,In_1578,In_888);
and U2622 (N_2622,In_629,In_1810);
nor U2623 (N_2623,In_1763,In_679);
nor U2624 (N_2624,In_1700,In_221);
and U2625 (N_2625,In_584,In_404);
nand U2626 (N_2626,In_69,In_934);
nand U2627 (N_2627,In_797,In_914);
or U2628 (N_2628,In_979,In_1587);
nor U2629 (N_2629,In_1532,In_1423);
nand U2630 (N_2630,In_435,In_733);
and U2631 (N_2631,In_1274,In_773);
and U2632 (N_2632,In_207,In_1235);
and U2633 (N_2633,In_678,In_1029);
and U2634 (N_2634,In_625,In_1951);
and U2635 (N_2635,In_448,In_1027);
or U2636 (N_2636,In_1861,In_1121);
nor U2637 (N_2637,In_941,In_1030);
nand U2638 (N_2638,In_733,In_1838);
nand U2639 (N_2639,In_387,In_1555);
nand U2640 (N_2640,In_1840,In_301);
or U2641 (N_2641,In_1833,In_1883);
or U2642 (N_2642,In_1448,In_1786);
or U2643 (N_2643,In_1892,In_1716);
nor U2644 (N_2644,In_1959,In_926);
and U2645 (N_2645,In_1025,In_1020);
nand U2646 (N_2646,In_1536,In_1197);
nand U2647 (N_2647,In_957,In_744);
and U2648 (N_2648,In_1470,In_1233);
nor U2649 (N_2649,In_1119,In_1896);
or U2650 (N_2650,In_1120,In_907);
nand U2651 (N_2651,In_112,In_107);
nand U2652 (N_2652,In_1045,In_435);
or U2653 (N_2653,In_1662,In_1710);
nand U2654 (N_2654,In_1710,In_1177);
nor U2655 (N_2655,In_1633,In_1652);
nor U2656 (N_2656,In_1111,In_697);
nand U2657 (N_2657,In_1759,In_844);
nand U2658 (N_2658,In_1381,In_1720);
or U2659 (N_2659,In_502,In_998);
and U2660 (N_2660,In_1408,In_1580);
or U2661 (N_2661,In_1054,In_1981);
and U2662 (N_2662,In_1514,In_963);
and U2663 (N_2663,In_1401,In_1204);
or U2664 (N_2664,In_260,In_1800);
nand U2665 (N_2665,In_1160,In_1161);
nand U2666 (N_2666,In_857,In_1503);
or U2667 (N_2667,In_257,In_398);
nand U2668 (N_2668,In_1202,In_383);
nand U2669 (N_2669,In_104,In_1894);
and U2670 (N_2670,In_1275,In_423);
or U2671 (N_2671,In_908,In_451);
nor U2672 (N_2672,In_872,In_1405);
and U2673 (N_2673,In_1219,In_828);
nor U2674 (N_2674,In_959,In_518);
or U2675 (N_2675,In_1984,In_59);
or U2676 (N_2676,In_756,In_213);
or U2677 (N_2677,In_328,In_973);
and U2678 (N_2678,In_659,In_1539);
nor U2679 (N_2679,In_1084,In_34);
and U2680 (N_2680,In_1569,In_1300);
and U2681 (N_2681,In_1198,In_1923);
nor U2682 (N_2682,In_1596,In_918);
nor U2683 (N_2683,In_1876,In_1592);
nor U2684 (N_2684,In_1885,In_1727);
or U2685 (N_2685,In_195,In_1859);
nor U2686 (N_2686,In_1795,In_1981);
and U2687 (N_2687,In_705,In_831);
or U2688 (N_2688,In_343,In_1823);
nand U2689 (N_2689,In_672,In_744);
nor U2690 (N_2690,In_30,In_260);
nor U2691 (N_2691,In_994,In_1451);
nand U2692 (N_2692,In_469,In_1740);
nand U2693 (N_2693,In_40,In_1368);
or U2694 (N_2694,In_1165,In_1554);
nand U2695 (N_2695,In_382,In_1725);
nor U2696 (N_2696,In_102,In_402);
or U2697 (N_2697,In_678,In_439);
and U2698 (N_2698,In_1344,In_1715);
nand U2699 (N_2699,In_286,In_1197);
nor U2700 (N_2700,In_1572,In_1522);
nor U2701 (N_2701,In_1995,In_1089);
or U2702 (N_2702,In_1831,In_1925);
nand U2703 (N_2703,In_1720,In_514);
nor U2704 (N_2704,In_1397,In_420);
or U2705 (N_2705,In_1414,In_174);
and U2706 (N_2706,In_1009,In_365);
and U2707 (N_2707,In_887,In_1816);
or U2708 (N_2708,In_888,In_1467);
and U2709 (N_2709,In_889,In_621);
and U2710 (N_2710,In_1768,In_1075);
and U2711 (N_2711,In_488,In_552);
and U2712 (N_2712,In_385,In_1826);
nand U2713 (N_2713,In_1980,In_839);
or U2714 (N_2714,In_1612,In_1962);
xnor U2715 (N_2715,In_323,In_414);
nand U2716 (N_2716,In_199,In_1337);
and U2717 (N_2717,In_1700,In_1987);
or U2718 (N_2718,In_753,In_505);
and U2719 (N_2719,In_257,In_1358);
and U2720 (N_2720,In_829,In_1009);
and U2721 (N_2721,In_1341,In_535);
nand U2722 (N_2722,In_35,In_115);
nand U2723 (N_2723,In_244,In_41);
or U2724 (N_2724,In_956,In_1746);
nor U2725 (N_2725,In_1438,In_644);
nor U2726 (N_2726,In_560,In_1654);
nand U2727 (N_2727,In_637,In_554);
nor U2728 (N_2728,In_226,In_21);
nand U2729 (N_2729,In_931,In_1553);
nand U2730 (N_2730,In_1528,In_1906);
and U2731 (N_2731,In_1701,In_894);
or U2732 (N_2732,In_1103,In_1269);
or U2733 (N_2733,In_939,In_1306);
nor U2734 (N_2734,In_648,In_1760);
nand U2735 (N_2735,In_1401,In_146);
nor U2736 (N_2736,In_1785,In_177);
and U2737 (N_2737,In_192,In_1861);
and U2738 (N_2738,In_27,In_1111);
nor U2739 (N_2739,In_498,In_613);
or U2740 (N_2740,In_1253,In_77);
and U2741 (N_2741,In_1636,In_1265);
or U2742 (N_2742,In_521,In_1954);
nand U2743 (N_2743,In_1466,In_1404);
nand U2744 (N_2744,In_1950,In_276);
or U2745 (N_2745,In_1586,In_1047);
nor U2746 (N_2746,In_1980,In_1725);
and U2747 (N_2747,In_360,In_1769);
nor U2748 (N_2748,In_4,In_1437);
nor U2749 (N_2749,In_1344,In_823);
or U2750 (N_2750,In_1177,In_1294);
and U2751 (N_2751,In_1518,In_889);
nand U2752 (N_2752,In_192,In_1297);
or U2753 (N_2753,In_1729,In_1985);
or U2754 (N_2754,In_343,In_1933);
nand U2755 (N_2755,In_770,In_166);
or U2756 (N_2756,In_1677,In_762);
and U2757 (N_2757,In_242,In_733);
nand U2758 (N_2758,In_83,In_1802);
nor U2759 (N_2759,In_881,In_108);
nor U2760 (N_2760,In_993,In_207);
or U2761 (N_2761,In_243,In_1162);
or U2762 (N_2762,In_925,In_297);
nor U2763 (N_2763,In_1671,In_1053);
and U2764 (N_2764,In_1120,In_1643);
nor U2765 (N_2765,In_116,In_323);
nand U2766 (N_2766,In_877,In_837);
nand U2767 (N_2767,In_650,In_43);
and U2768 (N_2768,In_1374,In_750);
or U2769 (N_2769,In_1191,In_298);
and U2770 (N_2770,In_1633,In_1092);
nor U2771 (N_2771,In_1884,In_1860);
nor U2772 (N_2772,In_1980,In_1441);
nor U2773 (N_2773,In_1742,In_1208);
nor U2774 (N_2774,In_42,In_510);
nor U2775 (N_2775,In_402,In_1588);
and U2776 (N_2776,In_869,In_1457);
nor U2777 (N_2777,In_984,In_917);
nand U2778 (N_2778,In_870,In_1289);
nand U2779 (N_2779,In_826,In_71);
nand U2780 (N_2780,In_754,In_1444);
and U2781 (N_2781,In_1783,In_1403);
nor U2782 (N_2782,In_1412,In_406);
nand U2783 (N_2783,In_1651,In_1006);
nand U2784 (N_2784,In_625,In_600);
or U2785 (N_2785,In_1857,In_1628);
or U2786 (N_2786,In_1301,In_174);
nor U2787 (N_2787,In_751,In_1129);
and U2788 (N_2788,In_1670,In_345);
nand U2789 (N_2789,In_1794,In_1480);
or U2790 (N_2790,In_471,In_104);
or U2791 (N_2791,In_942,In_477);
or U2792 (N_2792,In_557,In_1880);
nor U2793 (N_2793,In_1574,In_68);
nor U2794 (N_2794,In_161,In_1898);
or U2795 (N_2795,In_464,In_1008);
and U2796 (N_2796,In_1566,In_1904);
and U2797 (N_2797,In_1781,In_1322);
nor U2798 (N_2798,In_703,In_1649);
nor U2799 (N_2799,In_1362,In_1001);
or U2800 (N_2800,In_615,In_1750);
nand U2801 (N_2801,In_1325,In_1070);
and U2802 (N_2802,In_270,In_1772);
nand U2803 (N_2803,In_1658,In_81);
nor U2804 (N_2804,In_1272,In_672);
and U2805 (N_2805,In_1081,In_1327);
nor U2806 (N_2806,In_1066,In_982);
and U2807 (N_2807,In_429,In_1511);
or U2808 (N_2808,In_829,In_36);
nor U2809 (N_2809,In_899,In_1507);
nand U2810 (N_2810,In_1083,In_845);
nor U2811 (N_2811,In_275,In_270);
nand U2812 (N_2812,In_296,In_1676);
nand U2813 (N_2813,In_1319,In_534);
and U2814 (N_2814,In_306,In_1156);
and U2815 (N_2815,In_96,In_1496);
and U2816 (N_2816,In_606,In_1200);
nand U2817 (N_2817,In_1659,In_1597);
nor U2818 (N_2818,In_110,In_396);
nor U2819 (N_2819,In_1279,In_548);
and U2820 (N_2820,In_1151,In_1122);
or U2821 (N_2821,In_1772,In_449);
nand U2822 (N_2822,In_1505,In_1725);
nand U2823 (N_2823,In_273,In_484);
or U2824 (N_2824,In_1042,In_1619);
or U2825 (N_2825,In_113,In_1946);
or U2826 (N_2826,In_238,In_1269);
or U2827 (N_2827,In_1253,In_533);
and U2828 (N_2828,In_1632,In_618);
nor U2829 (N_2829,In_1355,In_1420);
nand U2830 (N_2830,In_1842,In_1361);
nand U2831 (N_2831,In_787,In_1118);
or U2832 (N_2832,In_278,In_824);
nand U2833 (N_2833,In_1327,In_503);
or U2834 (N_2834,In_1622,In_288);
and U2835 (N_2835,In_1133,In_25);
nand U2836 (N_2836,In_201,In_1861);
and U2837 (N_2837,In_1979,In_80);
and U2838 (N_2838,In_340,In_1100);
and U2839 (N_2839,In_775,In_1984);
or U2840 (N_2840,In_911,In_547);
and U2841 (N_2841,In_380,In_249);
and U2842 (N_2842,In_1945,In_819);
nand U2843 (N_2843,In_52,In_43);
and U2844 (N_2844,In_1073,In_1884);
and U2845 (N_2845,In_1506,In_109);
and U2846 (N_2846,In_1341,In_22);
nand U2847 (N_2847,In_876,In_737);
and U2848 (N_2848,In_1423,In_1982);
nor U2849 (N_2849,In_828,In_194);
nand U2850 (N_2850,In_248,In_1108);
nor U2851 (N_2851,In_1137,In_1020);
nand U2852 (N_2852,In_1402,In_1084);
nor U2853 (N_2853,In_1493,In_1945);
and U2854 (N_2854,In_1135,In_1055);
nand U2855 (N_2855,In_460,In_1245);
and U2856 (N_2856,In_758,In_237);
nand U2857 (N_2857,In_1951,In_1151);
or U2858 (N_2858,In_100,In_626);
nand U2859 (N_2859,In_1638,In_1925);
or U2860 (N_2860,In_873,In_553);
nand U2861 (N_2861,In_1008,In_106);
nand U2862 (N_2862,In_871,In_307);
or U2863 (N_2863,In_1904,In_1520);
and U2864 (N_2864,In_1715,In_408);
or U2865 (N_2865,In_1626,In_1679);
nor U2866 (N_2866,In_1369,In_1650);
nor U2867 (N_2867,In_805,In_1466);
or U2868 (N_2868,In_238,In_1204);
and U2869 (N_2869,In_539,In_1349);
nor U2870 (N_2870,In_389,In_1655);
nand U2871 (N_2871,In_1155,In_330);
and U2872 (N_2872,In_582,In_97);
nor U2873 (N_2873,In_102,In_1210);
and U2874 (N_2874,In_407,In_1901);
or U2875 (N_2875,In_1473,In_1721);
nor U2876 (N_2876,In_1221,In_163);
and U2877 (N_2877,In_1885,In_1779);
and U2878 (N_2878,In_1202,In_894);
nand U2879 (N_2879,In_1720,In_25);
and U2880 (N_2880,In_721,In_7);
xor U2881 (N_2881,In_131,In_970);
nand U2882 (N_2882,In_1598,In_1349);
or U2883 (N_2883,In_1775,In_1931);
nand U2884 (N_2884,In_120,In_1465);
or U2885 (N_2885,In_318,In_1156);
nor U2886 (N_2886,In_543,In_861);
or U2887 (N_2887,In_1264,In_569);
and U2888 (N_2888,In_1484,In_263);
or U2889 (N_2889,In_164,In_80);
nor U2890 (N_2890,In_1348,In_285);
nand U2891 (N_2891,In_1099,In_12);
and U2892 (N_2892,In_1331,In_690);
or U2893 (N_2893,In_584,In_364);
nand U2894 (N_2894,In_455,In_1812);
nand U2895 (N_2895,In_1675,In_1231);
nand U2896 (N_2896,In_851,In_1568);
nand U2897 (N_2897,In_114,In_535);
nand U2898 (N_2898,In_1289,In_2);
and U2899 (N_2899,In_782,In_1040);
nor U2900 (N_2900,In_1908,In_1594);
and U2901 (N_2901,In_1132,In_1932);
and U2902 (N_2902,In_1654,In_192);
nand U2903 (N_2903,In_1375,In_428);
nand U2904 (N_2904,In_1500,In_878);
or U2905 (N_2905,In_1406,In_1490);
nor U2906 (N_2906,In_1912,In_229);
nand U2907 (N_2907,In_301,In_1128);
or U2908 (N_2908,In_1858,In_273);
nand U2909 (N_2909,In_602,In_1322);
or U2910 (N_2910,In_1537,In_358);
or U2911 (N_2911,In_287,In_1270);
nor U2912 (N_2912,In_906,In_1124);
nor U2913 (N_2913,In_982,In_1189);
nand U2914 (N_2914,In_1764,In_1577);
nor U2915 (N_2915,In_988,In_865);
and U2916 (N_2916,In_1044,In_967);
and U2917 (N_2917,In_635,In_1420);
nor U2918 (N_2918,In_1601,In_1974);
or U2919 (N_2919,In_1377,In_1368);
nand U2920 (N_2920,In_1142,In_1765);
nand U2921 (N_2921,In_1358,In_1103);
nand U2922 (N_2922,In_588,In_817);
and U2923 (N_2923,In_1854,In_777);
xor U2924 (N_2924,In_1369,In_1415);
nor U2925 (N_2925,In_14,In_1467);
or U2926 (N_2926,In_1024,In_1858);
nand U2927 (N_2927,In_268,In_1596);
nor U2928 (N_2928,In_1211,In_885);
or U2929 (N_2929,In_1764,In_699);
or U2930 (N_2930,In_1636,In_1593);
nand U2931 (N_2931,In_1716,In_1922);
and U2932 (N_2932,In_442,In_995);
nor U2933 (N_2933,In_690,In_906);
nand U2934 (N_2934,In_1008,In_315);
nor U2935 (N_2935,In_824,In_1587);
or U2936 (N_2936,In_326,In_1425);
and U2937 (N_2937,In_137,In_50);
and U2938 (N_2938,In_1064,In_1901);
nor U2939 (N_2939,In_1786,In_1320);
or U2940 (N_2940,In_26,In_1346);
nor U2941 (N_2941,In_1648,In_1045);
nor U2942 (N_2942,In_988,In_1353);
nand U2943 (N_2943,In_1218,In_300);
nor U2944 (N_2944,In_1280,In_633);
or U2945 (N_2945,In_477,In_1441);
or U2946 (N_2946,In_1098,In_856);
nor U2947 (N_2947,In_703,In_1529);
and U2948 (N_2948,In_303,In_647);
and U2949 (N_2949,In_1974,In_295);
nor U2950 (N_2950,In_1462,In_1354);
and U2951 (N_2951,In_1690,In_1813);
xnor U2952 (N_2952,In_1269,In_1914);
nor U2953 (N_2953,In_255,In_1631);
nand U2954 (N_2954,In_1370,In_186);
and U2955 (N_2955,In_1362,In_1327);
and U2956 (N_2956,In_1923,In_371);
nand U2957 (N_2957,In_15,In_405);
nand U2958 (N_2958,In_70,In_1890);
or U2959 (N_2959,In_1977,In_1286);
nand U2960 (N_2960,In_401,In_756);
or U2961 (N_2961,In_1429,In_1528);
or U2962 (N_2962,In_312,In_1329);
nand U2963 (N_2963,In_1418,In_1025);
nor U2964 (N_2964,In_725,In_464);
nor U2965 (N_2965,In_1269,In_303);
nor U2966 (N_2966,In_1455,In_564);
and U2967 (N_2967,In_891,In_170);
or U2968 (N_2968,In_997,In_1475);
nor U2969 (N_2969,In_1511,In_125);
and U2970 (N_2970,In_656,In_1572);
nand U2971 (N_2971,In_1988,In_604);
or U2972 (N_2972,In_1409,In_1402);
or U2973 (N_2973,In_1335,In_652);
or U2974 (N_2974,In_108,In_1248);
nand U2975 (N_2975,In_1641,In_889);
or U2976 (N_2976,In_816,In_892);
nand U2977 (N_2977,In_1242,In_45);
nand U2978 (N_2978,In_585,In_1734);
nand U2979 (N_2979,In_1405,In_461);
or U2980 (N_2980,In_242,In_1264);
nand U2981 (N_2981,In_962,In_503);
or U2982 (N_2982,In_1971,In_207);
or U2983 (N_2983,In_1468,In_1246);
and U2984 (N_2984,In_242,In_662);
nor U2985 (N_2985,In_367,In_1636);
nor U2986 (N_2986,In_1650,In_814);
or U2987 (N_2987,In_1928,In_452);
nand U2988 (N_2988,In_652,In_73);
nor U2989 (N_2989,In_1961,In_606);
nand U2990 (N_2990,In_1942,In_1678);
nor U2991 (N_2991,In_1741,In_1014);
or U2992 (N_2992,In_1522,In_1840);
nand U2993 (N_2993,In_1119,In_339);
nand U2994 (N_2994,In_1846,In_812);
nand U2995 (N_2995,In_1977,In_1766);
and U2996 (N_2996,In_486,In_1227);
or U2997 (N_2997,In_246,In_1790);
nor U2998 (N_2998,In_1382,In_499);
and U2999 (N_2999,In_444,In_1601);
nand U3000 (N_3000,In_1653,In_295);
nand U3001 (N_3001,In_634,In_449);
or U3002 (N_3002,In_508,In_1819);
and U3003 (N_3003,In_701,In_1322);
and U3004 (N_3004,In_332,In_532);
and U3005 (N_3005,In_1743,In_871);
nor U3006 (N_3006,In_59,In_42);
nand U3007 (N_3007,In_157,In_357);
and U3008 (N_3008,In_979,In_67);
nand U3009 (N_3009,In_56,In_1525);
nor U3010 (N_3010,In_1963,In_599);
nand U3011 (N_3011,In_468,In_5);
nand U3012 (N_3012,In_1757,In_1234);
nand U3013 (N_3013,In_1881,In_26);
nor U3014 (N_3014,In_1927,In_339);
or U3015 (N_3015,In_1321,In_120);
and U3016 (N_3016,In_232,In_415);
or U3017 (N_3017,In_1025,In_1124);
nor U3018 (N_3018,In_901,In_1095);
or U3019 (N_3019,In_628,In_1773);
nor U3020 (N_3020,In_1051,In_515);
or U3021 (N_3021,In_723,In_330);
or U3022 (N_3022,In_560,In_1416);
nor U3023 (N_3023,In_1293,In_369);
nor U3024 (N_3024,In_425,In_143);
nor U3025 (N_3025,In_1562,In_65);
or U3026 (N_3026,In_385,In_1397);
nand U3027 (N_3027,In_943,In_1468);
nor U3028 (N_3028,In_947,In_524);
nand U3029 (N_3029,In_940,In_1148);
nand U3030 (N_3030,In_1505,In_1377);
or U3031 (N_3031,In_1782,In_194);
nand U3032 (N_3032,In_582,In_1774);
or U3033 (N_3033,In_217,In_1806);
and U3034 (N_3034,In_1214,In_257);
and U3035 (N_3035,In_469,In_1698);
nand U3036 (N_3036,In_29,In_545);
nor U3037 (N_3037,In_342,In_1384);
nor U3038 (N_3038,In_1119,In_773);
nor U3039 (N_3039,In_1751,In_1593);
nor U3040 (N_3040,In_1764,In_1002);
xnor U3041 (N_3041,In_1429,In_1562);
and U3042 (N_3042,In_1623,In_1231);
and U3043 (N_3043,In_221,In_775);
and U3044 (N_3044,In_1276,In_250);
nor U3045 (N_3045,In_1458,In_1925);
and U3046 (N_3046,In_210,In_698);
nand U3047 (N_3047,In_634,In_270);
and U3048 (N_3048,In_1726,In_1076);
and U3049 (N_3049,In_535,In_258);
nor U3050 (N_3050,In_1727,In_603);
and U3051 (N_3051,In_114,In_1709);
xnor U3052 (N_3052,In_884,In_1045);
nand U3053 (N_3053,In_659,In_1393);
or U3054 (N_3054,In_1875,In_170);
nand U3055 (N_3055,In_1387,In_1483);
nand U3056 (N_3056,In_523,In_1787);
nor U3057 (N_3057,In_1816,In_901);
or U3058 (N_3058,In_1624,In_1552);
nor U3059 (N_3059,In_255,In_52);
and U3060 (N_3060,In_475,In_1084);
and U3061 (N_3061,In_1013,In_1962);
and U3062 (N_3062,In_716,In_108);
and U3063 (N_3063,In_1437,In_1224);
and U3064 (N_3064,In_1834,In_351);
and U3065 (N_3065,In_1344,In_1805);
and U3066 (N_3066,In_66,In_711);
and U3067 (N_3067,In_635,In_871);
or U3068 (N_3068,In_1570,In_1940);
nand U3069 (N_3069,In_941,In_1420);
nand U3070 (N_3070,In_799,In_516);
nand U3071 (N_3071,In_1155,In_339);
nor U3072 (N_3072,In_1534,In_1207);
nand U3073 (N_3073,In_1663,In_1055);
nand U3074 (N_3074,In_1362,In_831);
and U3075 (N_3075,In_1273,In_1893);
or U3076 (N_3076,In_1064,In_616);
and U3077 (N_3077,In_1149,In_1474);
nor U3078 (N_3078,In_1632,In_53);
and U3079 (N_3079,In_1693,In_580);
and U3080 (N_3080,In_1754,In_496);
nand U3081 (N_3081,In_1112,In_1951);
and U3082 (N_3082,In_880,In_1024);
nor U3083 (N_3083,In_1964,In_1399);
and U3084 (N_3084,In_1879,In_1449);
or U3085 (N_3085,In_935,In_175);
nor U3086 (N_3086,In_494,In_1217);
nor U3087 (N_3087,In_1497,In_1462);
nor U3088 (N_3088,In_1555,In_348);
nor U3089 (N_3089,In_1114,In_1494);
or U3090 (N_3090,In_1633,In_1218);
nand U3091 (N_3091,In_1157,In_1363);
nand U3092 (N_3092,In_1877,In_1043);
and U3093 (N_3093,In_258,In_1507);
nor U3094 (N_3094,In_369,In_1513);
nand U3095 (N_3095,In_1778,In_1941);
nor U3096 (N_3096,In_1376,In_815);
or U3097 (N_3097,In_395,In_654);
nand U3098 (N_3098,In_2,In_1431);
or U3099 (N_3099,In_1304,In_274);
nand U3100 (N_3100,In_1295,In_1799);
and U3101 (N_3101,In_1432,In_1762);
nor U3102 (N_3102,In_1933,In_1554);
nand U3103 (N_3103,In_1492,In_532);
and U3104 (N_3104,In_153,In_1602);
nand U3105 (N_3105,In_1803,In_844);
nor U3106 (N_3106,In_1326,In_131);
or U3107 (N_3107,In_1525,In_1731);
nor U3108 (N_3108,In_1351,In_958);
nor U3109 (N_3109,In_1161,In_4);
nor U3110 (N_3110,In_1223,In_1194);
and U3111 (N_3111,In_1370,In_1293);
or U3112 (N_3112,In_1819,In_50);
nand U3113 (N_3113,In_1579,In_1680);
nor U3114 (N_3114,In_208,In_1096);
nor U3115 (N_3115,In_1375,In_1453);
nand U3116 (N_3116,In_239,In_1713);
nor U3117 (N_3117,In_1735,In_1447);
nand U3118 (N_3118,In_1620,In_824);
nand U3119 (N_3119,In_581,In_92);
and U3120 (N_3120,In_71,In_572);
nor U3121 (N_3121,In_440,In_408);
nand U3122 (N_3122,In_866,In_193);
and U3123 (N_3123,In_978,In_1273);
nand U3124 (N_3124,In_713,In_1997);
nor U3125 (N_3125,In_855,In_1526);
nor U3126 (N_3126,In_411,In_716);
or U3127 (N_3127,In_1834,In_909);
or U3128 (N_3128,In_1128,In_482);
and U3129 (N_3129,In_524,In_1668);
nor U3130 (N_3130,In_1013,In_1449);
nand U3131 (N_3131,In_1521,In_1850);
and U3132 (N_3132,In_1044,In_827);
and U3133 (N_3133,In_1922,In_1513);
nor U3134 (N_3134,In_1933,In_1342);
and U3135 (N_3135,In_1523,In_900);
and U3136 (N_3136,In_1824,In_316);
and U3137 (N_3137,In_68,In_669);
or U3138 (N_3138,In_941,In_575);
nand U3139 (N_3139,In_1231,In_1956);
and U3140 (N_3140,In_527,In_1274);
nand U3141 (N_3141,In_829,In_1544);
or U3142 (N_3142,In_788,In_309);
and U3143 (N_3143,In_1763,In_1060);
or U3144 (N_3144,In_674,In_296);
or U3145 (N_3145,In_1705,In_26);
nand U3146 (N_3146,In_638,In_1157);
nand U3147 (N_3147,In_48,In_755);
and U3148 (N_3148,In_223,In_1899);
or U3149 (N_3149,In_1158,In_1465);
nand U3150 (N_3150,In_461,In_1639);
or U3151 (N_3151,In_715,In_1926);
xor U3152 (N_3152,In_224,In_643);
nor U3153 (N_3153,In_877,In_1350);
or U3154 (N_3154,In_727,In_1074);
nand U3155 (N_3155,In_1234,In_1687);
nand U3156 (N_3156,In_672,In_963);
nor U3157 (N_3157,In_921,In_1130);
and U3158 (N_3158,In_741,In_239);
or U3159 (N_3159,In_128,In_447);
nand U3160 (N_3160,In_1042,In_1183);
or U3161 (N_3161,In_1729,In_411);
or U3162 (N_3162,In_1560,In_741);
or U3163 (N_3163,In_1023,In_93);
nand U3164 (N_3164,In_1402,In_404);
or U3165 (N_3165,In_1977,In_463);
and U3166 (N_3166,In_1143,In_1754);
or U3167 (N_3167,In_1960,In_1242);
nor U3168 (N_3168,In_1782,In_460);
nand U3169 (N_3169,In_1428,In_869);
nor U3170 (N_3170,In_1523,In_1478);
nor U3171 (N_3171,In_114,In_1740);
nor U3172 (N_3172,In_1300,In_916);
and U3173 (N_3173,In_1982,In_681);
nor U3174 (N_3174,In_1964,In_410);
or U3175 (N_3175,In_1616,In_1760);
nand U3176 (N_3176,In_1150,In_754);
and U3177 (N_3177,In_1709,In_344);
or U3178 (N_3178,In_512,In_1673);
and U3179 (N_3179,In_1973,In_278);
and U3180 (N_3180,In_302,In_216);
nor U3181 (N_3181,In_1175,In_1055);
and U3182 (N_3182,In_536,In_610);
or U3183 (N_3183,In_806,In_1086);
nand U3184 (N_3184,In_1577,In_1256);
nand U3185 (N_3185,In_750,In_1122);
and U3186 (N_3186,In_1637,In_541);
or U3187 (N_3187,In_1442,In_1213);
and U3188 (N_3188,In_1690,In_1027);
nor U3189 (N_3189,In_409,In_1183);
and U3190 (N_3190,In_1098,In_1476);
or U3191 (N_3191,In_242,In_368);
nand U3192 (N_3192,In_1905,In_783);
or U3193 (N_3193,In_491,In_678);
or U3194 (N_3194,In_25,In_191);
and U3195 (N_3195,In_269,In_262);
and U3196 (N_3196,In_898,In_1645);
xor U3197 (N_3197,In_1454,In_1508);
or U3198 (N_3198,In_73,In_1360);
and U3199 (N_3199,In_1236,In_1189);
and U3200 (N_3200,In_1784,In_955);
and U3201 (N_3201,In_508,In_588);
and U3202 (N_3202,In_701,In_621);
or U3203 (N_3203,In_644,In_1365);
nor U3204 (N_3204,In_1419,In_1136);
nor U3205 (N_3205,In_283,In_1489);
and U3206 (N_3206,In_1050,In_1862);
nor U3207 (N_3207,In_1365,In_614);
nor U3208 (N_3208,In_99,In_1931);
nand U3209 (N_3209,In_701,In_1388);
or U3210 (N_3210,In_1078,In_1558);
nand U3211 (N_3211,In_1750,In_1957);
nand U3212 (N_3212,In_1532,In_1685);
or U3213 (N_3213,In_1959,In_284);
or U3214 (N_3214,In_538,In_1248);
nor U3215 (N_3215,In_1536,In_1861);
or U3216 (N_3216,In_956,In_63);
and U3217 (N_3217,In_1805,In_906);
nor U3218 (N_3218,In_356,In_1094);
nor U3219 (N_3219,In_377,In_785);
or U3220 (N_3220,In_1005,In_175);
nor U3221 (N_3221,In_215,In_193);
nor U3222 (N_3222,In_576,In_1057);
and U3223 (N_3223,In_119,In_823);
or U3224 (N_3224,In_547,In_446);
and U3225 (N_3225,In_1667,In_1368);
nand U3226 (N_3226,In_1962,In_241);
and U3227 (N_3227,In_814,In_710);
nand U3228 (N_3228,In_1635,In_707);
and U3229 (N_3229,In_1166,In_1474);
or U3230 (N_3230,In_919,In_1786);
nand U3231 (N_3231,In_1134,In_1075);
and U3232 (N_3232,In_163,In_567);
and U3233 (N_3233,In_829,In_527);
and U3234 (N_3234,In_958,In_1443);
nand U3235 (N_3235,In_515,In_1801);
and U3236 (N_3236,In_209,In_1833);
nor U3237 (N_3237,In_1315,In_1931);
nor U3238 (N_3238,In_96,In_1650);
or U3239 (N_3239,In_354,In_748);
or U3240 (N_3240,In_340,In_1792);
nor U3241 (N_3241,In_851,In_1456);
nand U3242 (N_3242,In_1765,In_1);
and U3243 (N_3243,In_1852,In_1115);
and U3244 (N_3244,In_1435,In_48);
nand U3245 (N_3245,In_963,In_569);
nor U3246 (N_3246,In_79,In_1825);
or U3247 (N_3247,In_1291,In_1774);
nand U3248 (N_3248,In_34,In_85);
and U3249 (N_3249,In_208,In_1779);
or U3250 (N_3250,In_1247,In_156);
and U3251 (N_3251,In_1331,In_917);
nand U3252 (N_3252,In_1364,In_262);
and U3253 (N_3253,In_1965,In_1573);
or U3254 (N_3254,In_1302,In_882);
and U3255 (N_3255,In_758,In_1307);
nand U3256 (N_3256,In_750,In_1380);
or U3257 (N_3257,In_479,In_1640);
and U3258 (N_3258,In_667,In_788);
or U3259 (N_3259,In_1462,In_943);
or U3260 (N_3260,In_927,In_872);
or U3261 (N_3261,In_731,In_307);
nand U3262 (N_3262,In_1567,In_1590);
or U3263 (N_3263,In_1272,In_748);
nand U3264 (N_3264,In_705,In_1067);
nand U3265 (N_3265,In_1824,In_170);
and U3266 (N_3266,In_820,In_1627);
nor U3267 (N_3267,In_203,In_364);
nor U3268 (N_3268,In_1250,In_1893);
and U3269 (N_3269,In_1553,In_579);
and U3270 (N_3270,In_449,In_290);
and U3271 (N_3271,In_1983,In_1277);
nand U3272 (N_3272,In_1738,In_96);
or U3273 (N_3273,In_1332,In_1345);
xor U3274 (N_3274,In_54,In_1482);
nor U3275 (N_3275,In_1675,In_633);
or U3276 (N_3276,In_398,In_242);
and U3277 (N_3277,In_1719,In_1631);
and U3278 (N_3278,In_1429,In_1686);
nor U3279 (N_3279,In_211,In_585);
nor U3280 (N_3280,In_1915,In_1710);
nor U3281 (N_3281,In_1399,In_29);
and U3282 (N_3282,In_1555,In_1328);
nand U3283 (N_3283,In_790,In_894);
or U3284 (N_3284,In_1791,In_530);
nor U3285 (N_3285,In_535,In_362);
nor U3286 (N_3286,In_1536,In_832);
or U3287 (N_3287,In_208,In_607);
nor U3288 (N_3288,In_1636,In_245);
nand U3289 (N_3289,In_1268,In_1136);
nand U3290 (N_3290,In_1658,In_854);
or U3291 (N_3291,In_1422,In_92);
nor U3292 (N_3292,In_94,In_677);
xnor U3293 (N_3293,In_1873,In_1041);
and U3294 (N_3294,In_262,In_1779);
nand U3295 (N_3295,In_1369,In_1489);
and U3296 (N_3296,In_1708,In_597);
or U3297 (N_3297,In_1075,In_1702);
xor U3298 (N_3298,In_499,In_1991);
nand U3299 (N_3299,In_229,In_80);
or U3300 (N_3300,In_990,In_987);
nand U3301 (N_3301,In_1879,In_1792);
and U3302 (N_3302,In_1543,In_866);
or U3303 (N_3303,In_1147,In_421);
or U3304 (N_3304,In_12,In_1310);
or U3305 (N_3305,In_532,In_1246);
or U3306 (N_3306,In_623,In_1734);
or U3307 (N_3307,In_855,In_183);
and U3308 (N_3308,In_1323,In_1051);
or U3309 (N_3309,In_66,In_1260);
nand U3310 (N_3310,In_1918,In_702);
and U3311 (N_3311,In_1703,In_153);
nor U3312 (N_3312,In_744,In_1512);
and U3313 (N_3313,In_1585,In_425);
or U3314 (N_3314,In_307,In_424);
nand U3315 (N_3315,In_1945,In_626);
and U3316 (N_3316,In_1703,In_484);
nand U3317 (N_3317,In_1617,In_670);
or U3318 (N_3318,In_1001,In_340);
or U3319 (N_3319,In_1270,In_13);
or U3320 (N_3320,In_1741,In_678);
nand U3321 (N_3321,In_1266,In_120);
and U3322 (N_3322,In_1877,In_1576);
nor U3323 (N_3323,In_948,In_572);
or U3324 (N_3324,In_926,In_499);
nand U3325 (N_3325,In_1001,In_120);
or U3326 (N_3326,In_336,In_955);
nand U3327 (N_3327,In_34,In_1313);
and U3328 (N_3328,In_1682,In_1661);
nand U3329 (N_3329,In_1692,In_1679);
nand U3330 (N_3330,In_1260,In_1894);
nand U3331 (N_3331,In_192,In_650);
nand U3332 (N_3332,In_1858,In_958);
or U3333 (N_3333,In_1616,In_1453);
nand U3334 (N_3334,In_1553,In_1540);
nand U3335 (N_3335,In_1780,In_427);
or U3336 (N_3336,In_1522,In_1499);
and U3337 (N_3337,In_1354,In_1615);
or U3338 (N_3338,In_241,In_905);
nor U3339 (N_3339,In_944,In_1923);
or U3340 (N_3340,In_262,In_1366);
nand U3341 (N_3341,In_1525,In_854);
nand U3342 (N_3342,In_273,In_1500);
nor U3343 (N_3343,In_371,In_1903);
nand U3344 (N_3344,In_957,In_671);
nand U3345 (N_3345,In_143,In_1375);
and U3346 (N_3346,In_606,In_114);
or U3347 (N_3347,In_100,In_1271);
and U3348 (N_3348,In_1078,In_514);
or U3349 (N_3349,In_471,In_1200);
or U3350 (N_3350,In_1091,In_234);
or U3351 (N_3351,In_503,In_883);
nor U3352 (N_3352,In_300,In_1322);
and U3353 (N_3353,In_1616,In_325);
nand U3354 (N_3354,In_1113,In_1124);
nand U3355 (N_3355,In_582,In_1016);
or U3356 (N_3356,In_1029,In_949);
nand U3357 (N_3357,In_212,In_1893);
nor U3358 (N_3358,In_500,In_932);
nor U3359 (N_3359,In_1897,In_1082);
nand U3360 (N_3360,In_293,In_1989);
or U3361 (N_3361,In_139,In_935);
nand U3362 (N_3362,In_617,In_485);
nor U3363 (N_3363,In_87,In_1931);
nor U3364 (N_3364,In_948,In_19);
or U3365 (N_3365,In_1001,In_266);
and U3366 (N_3366,In_1245,In_282);
or U3367 (N_3367,In_1928,In_1032);
or U3368 (N_3368,In_991,In_152);
or U3369 (N_3369,In_1644,In_1610);
or U3370 (N_3370,In_1637,In_173);
nor U3371 (N_3371,In_1307,In_178);
and U3372 (N_3372,In_275,In_845);
nand U3373 (N_3373,In_683,In_1373);
and U3374 (N_3374,In_173,In_569);
nand U3375 (N_3375,In_1964,In_1540);
or U3376 (N_3376,In_1849,In_758);
nand U3377 (N_3377,In_675,In_1622);
and U3378 (N_3378,In_186,In_1201);
nand U3379 (N_3379,In_70,In_1515);
nor U3380 (N_3380,In_1517,In_1213);
and U3381 (N_3381,In_797,In_1914);
nand U3382 (N_3382,In_1881,In_1749);
nor U3383 (N_3383,In_573,In_728);
nor U3384 (N_3384,In_857,In_77);
nand U3385 (N_3385,In_145,In_958);
or U3386 (N_3386,In_1219,In_706);
nor U3387 (N_3387,In_388,In_330);
nor U3388 (N_3388,In_851,In_1227);
or U3389 (N_3389,In_1989,In_47);
or U3390 (N_3390,In_828,In_134);
xnor U3391 (N_3391,In_1796,In_1963);
or U3392 (N_3392,In_276,In_1963);
nor U3393 (N_3393,In_298,In_1106);
nor U3394 (N_3394,In_574,In_1454);
or U3395 (N_3395,In_1265,In_1916);
nor U3396 (N_3396,In_432,In_358);
nor U3397 (N_3397,In_221,In_933);
and U3398 (N_3398,In_661,In_704);
nand U3399 (N_3399,In_1211,In_319);
nand U3400 (N_3400,In_1490,In_1387);
nor U3401 (N_3401,In_65,In_1515);
or U3402 (N_3402,In_101,In_632);
nand U3403 (N_3403,In_1301,In_1615);
nor U3404 (N_3404,In_689,In_974);
and U3405 (N_3405,In_1965,In_1639);
nor U3406 (N_3406,In_364,In_40);
and U3407 (N_3407,In_569,In_1145);
nand U3408 (N_3408,In_919,In_535);
or U3409 (N_3409,In_88,In_1030);
or U3410 (N_3410,In_209,In_511);
nand U3411 (N_3411,In_1056,In_1680);
or U3412 (N_3412,In_1886,In_836);
nor U3413 (N_3413,In_941,In_1994);
nand U3414 (N_3414,In_355,In_1098);
or U3415 (N_3415,In_301,In_995);
nand U3416 (N_3416,In_1535,In_297);
and U3417 (N_3417,In_888,In_1541);
nand U3418 (N_3418,In_382,In_431);
nand U3419 (N_3419,In_1113,In_1941);
or U3420 (N_3420,In_212,In_1389);
nand U3421 (N_3421,In_442,In_654);
and U3422 (N_3422,In_1537,In_262);
and U3423 (N_3423,In_910,In_369);
and U3424 (N_3424,In_312,In_779);
or U3425 (N_3425,In_1016,In_962);
nand U3426 (N_3426,In_1273,In_971);
nand U3427 (N_3427,In_1101,In_1986);
and U3428 (N_3428,In_1488,In_225);
nor U3429 (N_3429,In_992,In_534);
or U3430 (N_3430,In_1450,In_810);
or U3431 (N_3431,In_1467,In_1200);
nand U3432 (N_3432,In_1802,In_1573);
nand U3433 (N_3433,In_1296,In_709);
nor U3434 (N_3434,In_387,In_25);
nor U3435 (N_3435,In_219,In_639);
nand U3436 (N_3436,In_1578,In_1759);
nor U3437 (N_3437,In_481,In_500);
nor U3438 (N_3438,In_1049,In_700);
or U3439 (N_3439,In_912,In_493);
and U3440 (N_3440,In_1851,In_1234);
nand U3441 (N_3441,In_89,In_671);
nand U3442 (N_3442,In_266,In_1440);
nand U3443 (N_3443,In_1338,In_1331);
or U3444 (N_3444,In_894,In_1686);
nand U3445 (N_3445,In_972,In_634);
nor U3446 (N_3446,In_768,In_646);
nor U3447 (N_3447,In_1951,In_847);
nor U3448 (N_3448,In_1533,In_1156);
nor U3449 (N_3449,In_1802,In_78);
nand U3450 (N_3450,In_610,In_1678);
and U3451 (N_3451,In_1651,In_933);
nand U3452 (N_3452,In_1197,In_1051);
nor U3453 (N_3453,In_276,In_1631);
nor U3454 (N_3454,In_901,In_715);
or U3455 (N_3455,In_1,In_330);
nor U3456 (N_3456,In_1957,In_1324);
nand U3457 (N_3457,In_675,In_1118);
and U3458 (N_3458,In_818,In_60);
nand U3459 (N_3459,In_1907,In_64);
nand U3460 (N_3460,In_1775,In_739);
and U3461 (N_3461,In_749,In_1730);
and U3462 (N_3462,In_1835,In_516);
and U3463 (N_3463,In_1722,In_1546);
nor U3464 (N_3464,In_1995,In_1771);
nor U3465 (N_3465,In_42,In_786);
nand U3466 (N_3466,In_1695,In_326);
or U3467 (N_3467,In_19,In_1283);
or U3468 (N_3468,In_1939,In_878);
nor U3469 (N_3469,In_1394,In_1331);
nand U3470 (N_3470,In_569,In_1909);
and U3471 (N_3471,In_208,In_389);
or U3472 (N_3472,In_988,In_107);
and U3473 (N_3473,In_469,In_462);
or U3474 (N_3474,In_1356,In_1244);
nor U3475 (N_3475,In_984,In_380);
nor U3476 (N_3476,In_198,In_769);
or U3477 (N_3477,In_875,In_973);
nand U3478 (N_3478,In_70,In_150);
xor U3479 (N_3479,In_1124,In_696);
and U3480 (N_3480,In_1027,In_1181);
nor U3481 (N_3481,In_1035,In_1210);
nor U3482 (N_3482,In_1992,In_921);
or U3483 (N_3483,In_1019,In_1639);
nor U3484 (N_3484,In_1413,In_1165);
nor U3485 (N_3485,In_1618,In_304);
nor U3486 (N_3486,In_1892,In_1622);
nor U3487 (N_3487,In_985,In_485);
and U3488 (N_3488,In_1479,In_1298);
nor U3489 (N_3489,In_115,In_1802);
nor U3490 (N_3490,In_783,In_410);
nor U3491 (N_3491,In_1390,In_1693);
and U3492 (N_3492,In_1105,In_1899);
and U3493 (N_3493,In_1785,In_974);
nor U3494 (N_3494,In_1357,In_812);
nand U3495 (N_3495,In_495,In_1794);
nand U3496 (N_3496,In_1541,In_1056);
or U3497 (N_3497,In_1319,In_1828);
nor U3498 (N_3498,In_503,In_694);
and U3499 (N_3499,In_286,In_254);
nand U3500 (N_3500,In_1985,In_1859);
nor U3501 (N_3501,In_972,In_1933);
nand U3502 (N_3502,In_496,In_1971);
nand U3503 (N_3503,In_1837,In_1127);
nand U3504 (N_3504,In_1766,In_1145);
nand U3505 (N_3505,In_969,In_944);
or U3506 (N_3506,In_1467,In_897);
and U3507 (N_3507,In_1722,In_139);
nor U3508 (N_3508,In_48,In_11);
nor U3509 (N_3509,In_1975,In_193);
and U3510 (N_3510,In_1937,In_1978);
xnor U3511 (N_3511,In_1636,In_1296);
nor U3512 (N_3512,In_1767,In_1568);
nor U3513 (N_3513,In_1177,In_1365);
nand U3514 (N_3514,In_1943,In_1825);
or U3515 (N_3515,In_2,In_1833);
and U3516 (N_3516,In_1657,In_880);
or U3517 (N_3517,In_1668,In_317);
and U3518 (N_3518,In_1556,In_1966);
and U3519 (N_3519,In_878,In_1231);
nand U3520 (N_3520,In_1963,In_602);
nand U3521 (N_3521,In_612,In_60);
nand U3522 (N_3522,In_1337,In_813);
xor U3523 (N_3523,In_841,In_1842);
nor U3524 (N_3524,In_1221,In_1267);
or U3525 (N_3525,In_1202,In_1676);
or U3526 (N_3526,In_108,In_1868);
nor U3527 (N_3527,In_1959,In_333);
or U3528 (N_3528,In_595,In_391);
or U3529 (N_3529,In_323,In_112);
or U3530 (N_3530,In_878,In_1724);
nor U3531 (N_3531,In_1300,In_109);
nand U3532 (N_3532,In_1911,In_869);
nor U3533 (N_3533,In_1718,In_628);
nand U3534 (N_3534,In_490,In_1512);
nand U3535 (N_3535,In_1404,In_1726);
nand U3536 (N_3536,In_910,In_1286);
and U3537 (N_3537,In_1749,In_1413);
or U3538 (N_3538,In_852,In_1301);
or U3539 (N_3539,In_1246,In_1488);
and U3540 (N_3540,In_1474,In_1535);
and U3541 (N_3541,In_1572,In_440);
nand U3542 (N_3542,In_575,In_1866);
nand U3543 (N_3543,In_1904,In_34);
or U3544 (N_3544,In_883,In_538);
or U3545 (N_3545,In_643,In_786);
and U3546 (N_3546,In_180,In_250);
nor U3547 (N_3547,In_160,In_1705);
and U3548 (N_3548,In_510,In_10);
nor U3549 (N_3549,In_48,In_627);
and U3550 (N_3550,In_1237,In_67);
nor U3551 (N_3551,In_1089,In_615);
nor U3552 (N_3552,In_1552,In_877);
nor U3553 (N_3553,In_1662,In_204);
and U3554 (N_3554,In_1766,In_730);
nand U3555 (N_3555,In_1058,In_216);
nor U3556 (N_3556,In_1164,In_1375);
nor U3557 (N_3557,In_1224,In_142);
nor U3558 (N_3558,In_728,In_1737);
or U3559 (N_3559,In_1494,In_1586);
nor U3560 (N_3560,In_79,In_806);
xor U3561 (N_3561,In_1796,In_240);
or U3562 (N_3562,In_871,In_666);
or U3563 (N_3563,In_1954,In_212);
nand U3564 (N_3564,In_885,In_345);
or U3565 (N_3565,In_1514,In_1231);
nand U3566 (N_3566,In_1093,In_1836);
or U3567 (N_3567,In_527,In_1379);
or U3568 (N_3568,In_704,In_1131);
and U3569 (N_3569,In_1632,In_16);
and U3570 (N_3570,In_1107,In_127);
and U3571 (N_3571,In_1976,In_1623);
and U3572 (N_3572,In_382,In_468);
nor U3573 (N_3573,In_352,In_491);
xnor U3574 (N_3574,In_1477,In_313);
and U3575 (N_3575,In_1719,In_364);
xnor U3576 (N_3576,In_260,In_1814);
and U3577 (N_3577,In_1964,In_627);
nor U3578 (N_3578,In_1134,In_1656);
xor U3579 (N_3579,In_1499,In_225);
and U3580 (N_3580,In_1501,In_841);
nor U3581 (N_3581,In_1157,In_1758);
nor U3582 (N_3582,In_1703,In_1504);
and U3583 (N_3583,In_1301,In_1998);
nand U3584 (N_3584,In_528,In_365);
and U3585 (N_3585,In_389,In_854);
or U3586 (N_3586,In_541,In_454);
or U3587 (N_3587,In_1410,In_405);
and U3588 (N_3588,In_1237,In_181);
nor U3589 (N_3589,In_678,In_979);
or U3590 (N_3590,In_1153,In_844);
nand U3591 (N_3591,In_1993,In_225);
nor U3592 (N_3592,In_77,In_1045);
nand U3593 (N_3593,In_914,In_767);
nand U3594 (N_3594,In_1989,In_1299);
and U3595 (N_3595,In_378,In_1666);
nor U3596 (N_3596,In_159,In_1113);
nand U3597 (N_3597,In_919,In_957);
or U3598 (N_3598,In_1225,In_1834);
or U3599 (N_3599,In_722,In_1062);
nor U3600 (N_3600,In_1659,In_1745);
and U3601 (N_3601,In_470,In_947);
or U3602 (N_3602,In_784,In_424);
nor U3603 (N_3603,In_1769,In_1736);
nand U3604 (N_3604,In_1766,In_136);
or U3605 (N_3605,In_1842,In_1654);
or U3606 (N_3606,In_1318,In_1562);
nor U3607 (N_3607,In_1843,In_458);
or U3608 (N_3608,In_1290,In_455);
nand U3609 (N_3609,In_1228,In_1527);
or U3610 (N_3610,In_356,In_1741);
nor U3611 (N_3611,In_1658,In_707);
and U3612 (N_3612,In_1679,In_754);
nand U3613 (N_3613,In_1715,In_223);
and U3614 (N_3614,In_1096,In_848);
nand U3615 (N_3615,In_1624,In_1279);
and U3616 (N_3616,In_425,In_176);
nor U3617 (N_3617,In_630,In_1179);
nor U3618 (N_3618,In_1821,In_1848);
or U3619 (N_3619,In_1866,In_491);
nor U3620 (N_3620,In_243,In_54);
nand U3621 (N_3621,In_838,In_895);
or U3622 (N_3622,In_917,In_724);
nor U3623 (N_3623,In_1277,In_1076);
or U3624 (N_3624,In_1329,In_1242);
nand U3625 (N_3625,In_1879,In_938);
and U3626 (N_3626,In_1748,In_1381);
nand U3627 (N_3627,In_1885,In_1577);
and U3628 (N_3628,In_1650,In_1928);
xnor U3629 (N_3629,In_576,In_1169);
or U3630 (N_3630,In_1332,In_1223);
nor U3631 (N_3631,In_215,In_187);
nor U3632 (N_3632,In_91,In_626);
nor U3633 (N_3633,In_1225,In_1601);
nor U3634 (N_3634,In_1655,In_1963);
or U3635 (N_3635,In_401,In_341);
nand U3636 (N_3636,In_1613,In_507);
nor U3637 (N_3637,In_1259,In_415);
nor U3638 (N_3638,In_546,In_1479);
and U3639 (N_3639,In_1302,In_191);
nor U3640 (N_3640,In_646,In_1377);
nand U3641 (N_3641,In_126,In_1494);
nand U3642 (N_3642,In_145,In_767);
or U3643 (N_3643,In_574,In_973);
nand U3644 (N_3644,In_960,In_1873);
nor U3645 (N_3645,In_1913,In_1240);
and U3646 (N_3646,In_1352,In_1906);
or U3647 (N_3647,In_1583,In_1879);
nor U3648 (N_3648,In_1472,In_1168);
nand U3649 (N_3649,In_645,In_1241);
nand U3650 (N_3650,In_678,In_25);
and U3651 (N_3651,In_1573,In_1314);
nor U3652 (N_3652,In_772,In_376);
nor U3653 (N_3653,In_1008,In_875);
nor U3654 (N_3654,In_1981,In_982);
nor U3655 (N_3655,In_313,In_1841);
or U3656 (N_3656,In_1504,In_1737);
nand U3657 (N_3657,In_1880,In_670);
and U3658 (N_3658,In_607,In_628);
nor U3659 (N_3659,In_189,In_1651);
nand U3660 (N_3660,In_1275,In_549);
and U3661 (N_3661,In_1993,In_312);
and U3662 (N_3662,In_1525,In_1088);
nor U3663 (N_3663,In_1691,In_1750);
and U3664 (N_3664,In_1401,In_463);
nand U3665 (N_3665,In_1793,In_355);
and U3666 (N_3666,In_1753,In_831);
or U3667 (N_3667,In_1781,In_713);
nand U3668 (N_3668,In_722,In_1963);
nor U3669 (N_3669,In_972,In_1729);
nand U3670 (N_3670,In_543,In_1792);
and U3671 (N_3671,In_225,In_322);
nand U3672 (N_3672,In_764,In_689);
nor U3673 (N_3673,In_725,In_1262);
nand U3674 (N_3674,In_1417,In_443);
nor U3675 (N_3675,In_1650,In_974);
or U3676 (N_3676,In_1558,In_387);
or U3677 (N_3677,In_1546,In_180);
or U3678 (N_3678,In_1053,In_1939);
nand U3679 (N_3679,In_1160,In_1649);
nor U3680 (N_3680,In_683,In_278);
or U3681 (N_3681,In_304,In_1486);
and U3682 (N_3682,In_1522,In_737);
nor U3683 (N_3683,In_1830,In_522);
nor U3684 (N_3684,In_163,In_1278);
nand U3685 (N_3685,In_694,In_484);
or U3686 (N_3686,In_561,In_1929);
or U3687 (N_3687,In_1282,In_1227);
or U3688 (N_3688,In_95,In_86);
nand U3689 (N_3689,In_1131,In_1021);
or U3690 (N_3690,In_26,In_225);
nand U3691 (N_3691,In_1178,In_233);
and U3692 (N_3692,In_1586,In_128);
nand U3693 (N_3693,In_1992,In_505);
nor U3694 (N_3694,In_1909,In_1138);
nor U3695 (N_3695,In_1115,In_78);
nor U3696 (N_3696,In_1707,In_1672);
nand U3697 (N_3697,In_1143,In_86);
and U3698 (N_3698,In_89,In_1185);
nor U3699 (N_3699,In_1759,In_369);
nor U3700 (N_3700,In_579,In_991);
nand U3701 (N_3701,In_760,In_1913);
nor U3702 (N_3702,In_1137,In_1079);
and U3703 (N_3703,In_1597,In_12);
nor U3704 (N_3704,In_1270,In_350);
nor U3705 (N_3705,In_211,In_1023);
nor U3706 (N_3706,In_1764,In_534);
nand U3707 (N_3707,In_1546,In_1693);
nor U3708 (N_3708,In_914,In_882);
and U3709 (N_3709,In_1534,In_17);
or U3710 (N_3710,In_869,In_252);
nor U3711 (N_3711,In_1703,In_1893);
and U3712 (N_3712,In_351,In_880);
nand U3713 (N_3713,In_652,In_1084);
or U3714 (N_3714,In_1937,In_1336);
nand U3715 (N_3715,In_898,In_1007);
and U3716 (N_3716,In_1719,In_1870);
nand U3717 (N_3717,In_960,In_1762);
nand U3718 (N_3718,In_1100,In_156);
nand U3719 (N_3719,In_1232,In_998);
and U3720 (N_3720,In_344,In_359);
or U3721 (N_3721,In_358,In_33);
nand U3722 (N_3722,In_721,In_1176);
nand U3723 (N_3723,In_1948,In_285);
nand U3724 (N_3724,In_907,In_316);
nor U3725 (N_3725,In_1049,In_936);
nor U3726 (N_3726,In_743,In_508);
or U3727 (N_3727,In_180,In_404);
or U3728 (N_3728,In_26,In_527);
and U3729 (N_3729,In_412,In_313);
nor U3730 (N_3730,In_1442,In_874);
and U3731 (N_3731,In_1922,In_310);
or U3732 (N_3732,In_1699,In_880);
or U3733 (N_3733,In_295,In_72);
and U3734 (N_3734,In_1194,In_1447);
or U3735 (N_3735,In_471,In_602);
nor U3736 (N_3736,In_239,In_1557);
and U3737 (N_3737,In_1030,In_1914);
or U3738 (N_3738,In_930,In_742);
xnor U3739 (N_3739,In_769,In_1267);
or U3740 (N_3740,In_1672,In_571);
nor U3741 (N_3741,In_853,In_985);
nand U3742 (N_3742,In_1822,In_1069);
nor U3743 (N_3743,In_1658,In_1485);
nand U3744 (N_3744,In_346,In_660);
nand U3745 (N_3745,In_1481,In_1474);
and U3746 (N_3746,In_1235,In_473);
or U3747 (N_3747,In_1382,In_182);
xnor U3748 (N_3748,In_933,In_1765);
and U3749 (N_3749,In_1705,In_959);
or U3750 (N_3750,In_1972,In_1289);
nand U3751 (N_3751,In_1772,In_1486);
nand U3752 (N_3752,In_72,In_757);
or U3753 (N_3753,In_1731,In_969);
nand U3754 (N_3754,In_1124,In_1457);
or U3755 (N_3755,In_1285,In_132);
nor U3756 (N_3756,In_1589,In_479);
and U3757 (N_3757,In_986,In_913);
nor U3758 (N_3758,In_1586,In_1548);
nand U3759 (N_3759,In_696,In_1092);
nand U3760 (N_3760,In_1807,In_1482);
nand U3761 (N_3761,In_1824,In_1379);
and U3762 (N_3762,In_1566,In_1970);
or U3763 (N_3763,In_154,In_1976);
nor U3764 (N_3764,In_1900,In_885);
and U3765 (N_3765,In_558,In_1473);
or U3766 (N_3766,In_1970,In_820);
nor U3767 (N_3767,In_1197,In_1640);
and U3768 (N_3768,In_25,In_1633);
nor U3769 (N_3769,In_380,In_577);
and U3770 (N_3770,In_1546,In_1345);
or U3771 (N_3771,In_858,In_221);
nor U3772 (N_3772,In_622,In_1620);
and U3773 (N_3773,In_813,In_279);
or U3774 (N_3774,In_652,In_983);
and U3775 (N_3775,In_1056,In_1681);
nand U3776 (N_3776,In_1832,In_1040);
and U3777 (N_3777,In_715,In_961);
and U3778 (N_3778,In_420,In_425);
or U3779 (N_3779,In_111,In_1333);
nor U3780 (N_3780,In_494,In_311);
and U3781 (N_3781,In_64,In_743);
and U3782 (N_3782,In_144,In_1720);
or U3783 (N_3783,In_598,In_813);
and U3784 (N_3784,In_476,In_1052);
nand U3785 (N_3785,In_1010,In_1434);
and U3786 (N_3786,In_894,In_896);
or U3787 (N_3787,In_9,In_69);
nor U3788 (N_3788,In_1216,In_985);
nand U3789 (N_3789,In_1814,In_1980);
nor U3790 (N_3790,In_1156,In_1993);
or U3791 (N_3791,In_598,In_1012);
nand U3792 (N_3792,In_223,In_1543);
nor U3793 (N_3793,In_1708,In_1059);
xnor U3794 (N_3794,In_742,In_311);
or U3795 (N_3795,In_278,In_480);
and U3796 (N_3796,In_93,In_972);
nor U3797 (N_3797,In_114,In_1511);
or U3798 (N_3798,In_854,In_1227);
and U3799 (N_3799,In_644,In_393);
nor U3800 (N_3800,In_1882,In_779);
nand U3801 (N_3801,In_641,In_1247);
or U3802 (N_3802,In_1061,In_697);
nor U3803 (N_3803,In_1428,In_223);
nand U3804 (N_3804,In_1992,In_1424);
nand U3805 (N_3805,In_859,In_1038);
nor U3806 (N_3806,In_741,In_377);
nor U3807 (N_3807,In_965,In_114);
nor U3808 (N_3808,In_1977,In_1094);
and U3809 (N_3809,In_1598,In_169);
nor U3810 (N_3810,In_954,In_518);
and U3811 (N_3811,In_419,In_300);
or U3812 (N_3812,In_844,In_1056);
nand U3813 (N_3813,In_859,In_14);
nor U3814 (N_3814,In_102,In_415);
nand U3815 (N_3815,In_50,In_1287);
nand U3816 (N_3816,In_1451,In_321);
nand U3817 (N_3817,In_244,In_427);
nor U3818 (N_3818,In_1994,In_1749);
nor U3819 (N_3819,In_1469,In_1219);
nor U3820 (N_3820,In_1279,In_1840);
nand U3821 (N_3821,In_1456,In_498);
or U3822 (N_3822,In_1289,In_1729);
nor U3823 (N_3823,In_185,In_903);
and U3824 (N_3824,In_570,In_1579);
or U3825 (N_3825,In_1979,In_88);
and U3826 (N_3826,In_1147,In_1389);
nor U3827 (N_3827,In_340,In_1464);
nand U3828 (N_3828,In_1679,In_729);
nand U3829 (N_3829,In_1155,In_1924);
and U3830 (N_3830,In_47,In_603);
and U3831 (N_3831,In_1580,In_1075);
and U3832 (N_3832,In_1787,In_278);
or U3833 (N_3833,In_1516,In_291);
nand U3834 (N_3834,In_980,In_1237);
nor U3835 (N_3835,In_478,In_192);
nor U3836 (N_3836,In_270,In_1894);
nand U3837 (N_3837,In_469,In_1137);
or U3838 (N_3838,In_1695,In_543);
nor U3839 (N_3839,In_877,In_1968);
nor U3840 (N_3840,In_236,In_651);
nor U3841 (N_3841,In_1312,In_475);
nor U3842 (N_3842,In_1442,In_1769);
or U3843 (N_3843,In_163,In_364);
and U3844 (N_3844,In_630,In_1076);
nor U3845 (N_3845,In_1551,In_885);
and U3846 (N_3846,In_613,In_668);
nand U3847 (N_3847,In_1625,In_442);
or U3848 (N_3848,In_1533,In_197);
nand U3849 (N_3849,In_854,In_1471);
nand U3850 (N_3850,In_784,In_951);
nor U3851 (N_3851,In_1685,In_912);
nor U3852 (N_3852,In_852,In_620);
and U3853 (N_3853,In_1929,In_304);
nand U3854 (N_3854,In_309,In_242);
nand U3855 (N_3855,In_1373,In_1092);
and U3856 (N_3856,In_283,In_1817);
nand U3857 (N_3857,In_1468,In_95);
and U3858 (N_3858,In_629,In_193);
or U3859 (N_3859,In_1105,In_1527);
nor U3860 (N_3860,In_1397,In_1874);
nor U3861 (N_3861,In_981,In_1303);
nor U3862 (N_3862,In_641,In_1736);
nand U3863 (N_3863,In_1451,In_1175);
and U3864 (N_3864,In_925,In_1596);
or U3865 (N_3865,In_448,In_1535);
nor U3866 (N_3866,In_229,In_1977);
nor U3867 (N_3867,In_731,In_250);
and U3868 (N_3868,In_294,In_1508);
or U3869 (N_3869,In_542,In_883);
or U3870 (N_3870,In_19,In_846);
and U3871 (N_3871,In_1571,In_398);
or U3872 (N_3872,In_1009,In_558);
nand U3873 (N_3873,In_309,In_1439);
xnor U3874 (N_3874,In_376,In_1674);
nand U3875 (N_3875,In_86,In_1963);
nand U3876 (N_3876,In_1492,In_961);
nand U3877 (N_3877,In_730,In_837);
nor U3878 (N_3878,In_1523,In_662);
nand U3879 (N_3879,In_806,In_670);
nand U3880 (N_3880,In_641,In_1747);
and U3881 (N_3881,In_1487,In_1520);
xor U3882 (N_3882,In_1843,In_488);
xnor U3883 (N_3883,In_481,In_1110);
nand U3884 (N_3884,In_532,In_1432);
or U3885 (N_3885,In_1881,In_1535);
or U3886 (N_3886,In_1770,In_2);
nor U3887 (N_3887,In_136,In_1327);
or U3888 (N_3888,In_208,In_1028);
and U3889 (N_3889,In_819,In_1457);
and U3890 (N_3890,In_335,In_903);
nor U3891 (N_3891,In_890,In_1177);
or U3892 (N_3892,In_255,In_1843);
nand U3893 (N_3893,In_1562,In_261);
nand U3894 (N_3894,In_1815,In_1361);
nand U3895 (N_3895,In_568,In_777);
nor U3896 (N_3896,In_816,In_1970);
and U3897 (N_3897,In_351,In_636);
and U3898 (N_3898,In_1879,In_83);
nor U3899 (N_3899,In_1174,In_1689);
or U3900 (N_3900,In_1652,In_350);
nand U3901 (N_3901,In_711,In_1471);
or U3902 (N_3902,In_1000,In_932);
or U3903 (N_3903,In_1265,In_1164);
or U3904 (N_3904,In_987,In_1893);
and U3905 (N_3905,In_891,In_994);
or U3906 (N_3906,In_1899,In_689);
and U3907 (N_3907,In_1949,In_1486);
or U3908 (N_3908,In_1467,In_1324);
or U3909 (N_3909,In_182,In_546);
and U3910 (N_3910,In_1084,In_541);
xnor U3911 (N_3911,In_8,In_138);
and U3912 (N_3912,In_959,In_1250);
nand U3913 (N_3913,In_1553,In_1284);
nor U3914 (N_3914,In_741,In_645);
or U3915 (N_3915,In_890,In_356);
and U3916 (N_3916,In_260,In_471);
nand U3917 (N_3917,In_222,In_462);
and U3918 (N_3918,In_1545,In_333);
nor U3919 (N_3919,In_788,In_359);
nand U3920 (N_3920,In_429,In_1870);
and U3921 (N_3921,In_330,In_508);
or U3922 (N_3922,In_1861,In_1706);
nand U3923 (N_3923,In_1781,In_538);
xnor U3924 (N_3924,In_1647,In_1430);
and U3925 (N_3925,In_1526,In_1822);
nor U3926 (N_3926,In_458,In_405);
nor U3927 (N_3927,In_1551,In_497);
nand U3928 (N_3928,In_723,In_452);
or U3929 (N_3929,In_164,In_743);
or U3930 (N_3930,In_1887,In_873);
nand U3931 (N_3931,In_571,In_519);
nand U3932 (N_3932,In_573,In_42);
or U3933 (N_3933,In_1656,In_741);
nand U3934 (N_3934,In_980,In_1981);
nor U3935 (N_3935,In_681,In_261);
nor U3936 (N_3936,In_1747,In_148);
and U3937 (N_3937,In_1974,In_1208);
nor U3938 (N_3938,In_542,In_707);
nand U3939 (N_3939,In_185,In_1476);
or U3940 (N_3940,In_1785,In_100);
or U3941 (N_3941,In_1187,In_885);
or U3942 (N_3942,In_1905,In_1507);
or U3943 (N_3943,In_258,In_1148);
or U3944 (N_3944,In_1367,In_1072);
and U3945 (N_3945,In_1131,In_1392);
or U3946 (N_3946,In_1066,In_1064);
nor U3947 (N_3947,In_246,In_612);
and U3948 (N_3948,In_955,In_144);
or U3949 (N_3949,In_352,In_381);
or U3950 (N_3950,In_1309,In_435);
and U3951 (N_3951,In_1678,In_242);
nand U3952 (N_3952,In_1885,In_1624);
nor U3953 (N_3953,In_812,In_1664);
nor U3954 (N_3954,In_140,In_269);
nor U3955 (N_3955,In_243,In_1709);
and U3956 (N_3956,In_1143,In_228);
or U3957 (N_3957,In_1733,In_236);
nand U3958 (N_3958,In_837,In_1740);
and U3959 (N_3959,In_1929,In_1246);
nor U3960 (N_3960,In_1542,In_503);
nor U3961 (N_3961,In_224,In_1531);
or U3962 (N_3962,In_1332,In_1690);
nor U3963 (N_3963,In_1802,In_761);
nor U3964 (N_3964,In_962,In_1321);
and U3965 (N_3965,In_817,In_409);
or U3966 (N_3966,In_1613,In_1334);
and U3967 (N_3967,In_187,In_845);
nand U3968 (N_3968,In_1590,In_33);
and U3969 (N_3969,In_1713,In_912);
or U3970 (N_3970,In_1425,In_586);
nand U3971 (N_3971,In_943,In_1659);
nand U3972 (N_3972,In_1655,In_742);
and U3973 (N_3973,In_1620,In_1400);
or U3974 (N_3974,In_1629,In_1340);
nand U3975 (N_3975,In_1826,In_844);
or U3976 (N_3976,In_1759,In_830);
and U3977 (N_3977,In_484,In_1839);
and U3978 (N_3978,In_449,In_13);
or U3979 (N_3979,In_1243,In_1321);
nor U3980 (N_3980,In_327,In_1664);
and U3981 (N_3981,In_1089,In_1220);
nand U3982 (N_3982,In_555,In_602);
nand U3983 (N_3983,In_1756,In_325);
nor U3984 (N_3984,In_1793,In_998);
or U3985 (N_3985,In_1727,In_701);
nor U3986 (N_3986,In_410,In_349);
or U3987 (N_3987,In_1799,In_1947);
nand U3988 (N_3988,In_204,In_1384);
nand U3989 (N_3989,In_1073,In_801);
nor U3990 (N_3990,In_1238,In_652);
nand U3991 (N_3991,In_782,In_761);
and U3992 (N_3992,In_1767,In_910);
and U3993 (N_3993,In_268,In_1519);
nand U3994 (N_3994,In_10,In_899);
and U3995 (N_3995,In_216,In_1238);
and U3996 (N_3996,In_865,In_1893);
and U3997 (N_3997,In_1355,In_1805);
or U3998 (N_3998,In_807,In_1712);
or U3999 (N_3999,In_1438,In_1852);
and U4000 (N_4000,In_117,In_830);
or U4001 (N_4001,In_225,In_790);
and U4002 (N_4002,In_1332,In_71);
or U4003 (N_4003,In_1317,In_348);
or U4004 (N_4004,In_1131,In_930);
and U4005 (N_4005,In_691,In_1046);
or U4006 (N_4006,In_904,In_1832);
and U4007 (N_4007,In_311,In_553);
or U4008 (N_4008,In_1249,In_1419);
nand U4009 (N_4009,In_594,In_1805);
xor U4010 (N_4010,In_1051,In_569);
or U4011 (N_4011,In_1055,In_329);
and U4012 (N_4012,In_1851,In_1196);
and U4013 (N_4013,In_1820,In_1591);
nand U4014 (N_4014,In_1520,In_1284);
nand U4015 (N_4015,In_713,In_1824);
nor U4016 (N_4016,In_1297,In_856);
nor U4017 (N_4017,In_1291,In_676);
nand U4018 (N_4018,In_1675,In_691);
and U4019 (N_4019,In_115,In_820);
and U4020 (N_4020,In_1017,In_100);
nand U4021 (N_4021,In_832,In_1176);
nand U4022 (N_4022,In_1837,In_1290);
nand U4023 (N_4023,In_781,In_439);
nor U4024 (N_4024,In_222,In_1374);
xor U4025 (N_4025,In_1426,In_802);
or U4026 (N_4026,In_275,In_306);
nor U4027 (N_4027,In_1205,In_1263);
nand U4028 (N_4028,In_1477,In_1852);
nor U4029 (N_4029,In_1493,In_1698);
or U4030 (N_4030,In_997,In_1400);
or U4031 (N_4031,In_776,In_946);
or U4032 (N_4032,In_53,In_1636);
and U4033 (N_4033,In_1584,In_1449);
and U4034 (N_4034,In_660,In_368);
and U4035 (N_4035,In_591,In_1929);
nand U4036 (N_4036,In_1351,In_1609);
or U4037 (N_4037,In_1132,In_756);
and U4038 (N_4038,In_1709,In_1637);
or U4039 (N_4039,In_1089,In_158);
or U4040 (N_4040,In_91,In_616);
and U4041 (N_4041,In_796,In_629);
nand U4042 (N_4042,In_311,In_412);
and U4043 (N_4043,In_480,In_192);
and U4044 (N_4044,In_144,In_1943);
and U4045 (N_4045,In_1811,In_1138);
or U4046 (N_4046,In_138,In_1523);
and U4047 (N_4047,In_404,In_864);
nor U4048 (N_4048,In_266,In_832);
nand U4049 (N_4049,In_385,In_1509);
nor U4050 (N_4050,In_240,In_1559);
and U4051 (N_4051,In_1107,In_1553);
and U4052 (N_4052,In_1453,In_965);
nand U4053 (N_4053,In_380,In_454);
nand U4054 (N_4054,In_181,In_748);
nand U4055 (N_4055,In_66,In_1542);
nor U4056 (N_4056,In_1202,In_1178);
or U4057 (N_4057,In_1605,In_1277);
and U4058 (N_4058,In_104,In_1458);
nand U4059 (N_4059,In_973,In_1509);
or U4060 (N_4060,In_918,In_1351);
nand U4061 (N_4061,In_547,In_1663);
nand U4062 (N_4062,In_1405,In_24);
xor U4063 (N_4063,In_59,In_962);
nor U4064 (N_4064,In_986,In_935);
nand U4065 (N_4065,In_78,In_874);
or U4066 (N_4066,In_1085,In_342);
nor U4067 (N_4067,In_170,In_476);
nand U4068 (N_4068,In_396,In_971);
nor U4069 (N_4069,In_1371,In_658);
and U4070 (N_4070,In_1279,In_100);
and U4071 (N_4071,In_1687,In_1602);
and U4072 (N_4072,In_1189,In_286);
nor U4073 (N_4073,In_682,In_1088);
nor U4074 (N_4074,In_1599,In_1842);
nor U4075 (N_4075,In_243,In_291);
nor U4076 (N_4076,In_1610,In_229);
or U4077 (N_4077,In_596,In_1998);
nor U4078 (N_4078,In_1857,In_246);
and U4079 (N_4079,In_87,In_1093);
nand U4080 (N_4080,In_1859,In_1843);
nor U4081 (N_4081,In_411,In_1962);
nand U4082 (N_4082,In_468,In_337);
nor U4083 (N_4083,In_86,In_1878);
and U4084 (N_4084,In_314,In_108);
and U4085 (N_4085,In_1029,In_1837);
or U4086 (N_4086,In_134,In_1604);
nor U4087 (N_4087,In_1641,In_431);
nor U4088 (N_4088,In_819,In_1397);
and U4089 (N_4089,In_181,In_805);
or U4090 (N_4090,In_189,In_836);
nand U4091 (N_4091,In_535,In_228);
or U4092 (N_4092,In_512,In_459);
or U4093 (N_4093,In_1951,In_1326);
or U4094 (N_4094,In_1906,In_1824);
and U4095 (N_4095,In_1892,In_862);
nor U4096 (N_4096,In_1133,In_1423);
and U4097 (N_4097,In_1445,In_1720);
or U4098 (N_4098,In_1316,In_1748);
nand U4099 (N_4099,In_860,In_1948);
and U4100 (N_4100,In_1743,In_437);
nor U4101 (N_4101,In_1976,In_1196);
and U4102 (N_4102,In_723,In_167);
or U4103 (N_4103,In_954,In_1095);
or U4104 (N_4104,In_411,In_500);
nor U4105 (N_4105,In_1281,In_129);
nor U4106 (N_4106,In_1582,In_1734);
and U4107 (N_4107,In_1220,In_90);
and U4108 (N_4108,In_1564,In_1372);
nor U4109 (N_4109,In_930,In_1264);
or U4110 (N_4110,In_904,In_1649);
or U4111 (N_4111,In_420,In_965);
nor U4112 (N_4112,In_1804,In_1447);
xnor U4113 (N_4113,In_25,In_1103);
and U4114 (N_4114,In_1441,In_175);
nand U4115 (N_4115,In_1507,In_1706);
or U4116 (N_4116,In_1550,In_1274);
nor U4117 (N_4117,In_287,In_259);
nor U4118 (N_4118,In_1546,In_415);
and U4119 (N_4119,In_1174,In_532);
nand U4120 (N_4120,In_1134,In_845);
or U4121 (N_4121,In_283,In_348);
and U4122 (N_4122,In_632,In_1415);
or U4123 (N_4123,In_279,In_1154);
nor U4124 (N_4124,In_1166,In_1992);
and U4125 (N_4125,In_1069,In_396);
nand U4126 (N_4126,In_1612,In_104);
nand U4127 (N_4127,In_670,In_895);
nand U4128 (N_4128,In_1581,In_912);
nor U4129 (N_4129,In_547,In_1636);
nor U4130 (N_4130,In_433,In_90);
or U4131 (N_4131,In_1980,In_1617);
nand U4132 (N_4132,In_744,In_1594);
nor U4133 (N_4133,In_1822,In_526);
or U4134 (N_4134,In_127,In_591);
or U4135 (N_4135,In_1680,In_1960);
or U4136 (N_4136,In_1579,In_1456);
and U4137 (N_4137,In_640,In_516);
and U4138 (N_4138,In_216,In_1443);
nor U4139 (N_4139,In_1577,In_809);
and U4140 (N_4140,In_1380,In_937);
nand U4141 (N_4141,In_974,In_1462);
nand U4142 (N_4142,In_1770,In_188);
or U4143 (N_4143,In_533,In_969);
or U4144 (N_4144,In_889,In_61);
xnor U4145 (N_4145,In_345,In_214);
and U4146 (N_4146,In_1685,In_1551);
or U4147 (N_4147,In_138,In_211);
xor U4148 (N_4148,In_440,In_1415);
or U4149 (N_4149,In_138,In_10);
and U4150 (N_4150,In_1650,In_35);
or U4151 (N_4151,In_1733,In_570);
xor U4152 (N_4152,In_902,In_611);
or U4153 (N_4153,In_1931,In_139);
and U4154 (N_4154,In_1209,In_1845);
or U4155 (N_4155,In_1604,In_812);
nand U4156 (N_4156,In_639,In_954);
or U4157 (N_4157,In_759,In_1155);
and U4158 (N_4158,In_1179,In_1928);
and U4159 (N_4159,In_1710,In_1872);
and U4160 (N_4160,In_1187,In_829);
and U4161 (N_4161,In_711,In_1720);
or U4162 (N_4162,In_1591,In_380);
nand U4163 (N_4163,In_1530,In_241);
nand U4164 (N_4164,In_994,In_1393);
nand U4165 (N_4165,In_331,In_1280);
nand U4166 (N_4166,In_1873,In_1162);
nand U4167 (N_4167,In_198,In_997);
nand U4168 (N_4168,In_1608,In_871);
or U4169 (N_4169,In_1444,In_535);
nand U4170 (N_4170,In_558,In_1465);
or U4171 (N_4171,In_1427,In_1008);
nand U4172 (N_4172,In_1086,In_1029);
and U4173 (N_4173,In_1146,In_1877);
and U4174 (N_4174,In_597,In_814);
nand U4175 (N_4175,In_1711,In_504);
or U4176 (N_4176,In_1856,In_121);
nor U4177 (N_4177,In_210,In_816);
nand U4178 (N_4178,In_992,In_1440);
nor U4179 (N_4179,In_680,In_253);
nand U4180 (N_4180,In_1350,In_1408);
nand U4181 (N_4181,In_1265,In_938);
and U4182 (N_4182,In_1728,In_181);
nor U4183 (N_4183,In_877,In_1796);
or U4184 (N_4184,In_338,In_319);
and U4185 (N_4185,In_716,In_1026);
and U4186 (N_4186,In_354,In_833);
nor U4187 (N_4187,In_1689,In_1028);
and U4188 (N_4188,In_346,In_927);
and U4189 (N_4189,In_447,In_1980);
nor U4190 (N_4190,In_1806,In_1959);
nand U4191 (N_4191,In_1981,In_1212);
and U4192 (N_4192,In_110,In_456);
and U4193 (N_4193,In_1143,In_1765);
nor U4194 (N_4194,In_856,In_1399);
and U4195 (N_4195,In_553,In_1765);
nand U4196 (N_4196,In_1772,In_558);
nand U4197 (N_4197,In_40,In_1233);
nor U4198 (N_4198,In_1335,In_71);
nand U4199 (N_4199,In_153,In_751);
nor U4200 (N_4200,In_179,In_605);
nor U4201 (N_4201,In_1436,In_376);
or U4202 (N_4202,In_1435,In_1543);
or U4203 (N_4203,In_252,In_1043);
and U4204 (N_4204,In_344,In_1987);
and U4205 (N_4205,In_1617,In_589);
nor U4206 (N_4206,In_736,In_1271);
or U4207 (N_4207,In_55,In_1456);
nor U4208 (N_4208,In_758,In_1702);
nor U4209 (N_4209,In_1559,In_46);
and U4210 (N_4210,In_834,In_720);
nor U4211 (N_4211,In_1095,In_179);
and U4212 (N_4212,In_89,In_1929);
nor U4213 (N_4213,In_165,In_388);
nor U4214 (N_4214,In_1493,In_1275);
nand U4215 (N_4215,In_1741,In_166);
or U4216 (N_4216,In_962,In_1677);
nand U4217 (N_4217,In_1834,In_1108);
and U4218 (N_4218,In_1147,In_799);
nand U4219 (N_4219,In_398,In_0);
nand U4220 (N_4220,In_1618,In_833);
nand U4221 (N_4221,In_859,In_613);
or U4222 (N_4222,In_72,In_1168);
and U4223 (N_4223,In_513,In_1149);
nor U4224 (N_4224,In_1782,In_1443);
nand U4225 (N_4225,In_1810,In_648);
nand U4226 (N_4226,In_1413,In_426);
or U4227 (N_4227,In_584,In_758);
and U4228 (N_4228,In_1871,In_130);
xnor U4229 (N_4229,In_258,In_1505);
or U4230 (N_4230,In_1689,In_510);
or U4231 (N_4231,In_956,In_1837);
or U4232 (N_4232,In_1480,In_1226);
nand U4233 (N_4233,In_1939,In_453);
and U4234 (N_4234,In_88,In_1497);
nand U4235 (N_4235,In_1948,In_338);
and U4236 (N_4236,In_1554,In_1490);
or U4237 (N_4237,In_822,In_190);
nor U4238 (N_4238,In_1282,In_227);
nand U4239 (N_4239,In_1251,In_1322);
and U4240 (N_4240,In_1833,In_1550);
and U4241 (N_4241,In_1126,In_312);
nor U4242 (N_4242,In_35,In_684);
nand U4243 (N_4243,In_1150,In_1066);
nor U4244 (N_4244,In_1466,In_466);
nor U4245 (N_4245,In_898,In_1202);
nor U4246 (N_4246,In_150,In_182);
xnor U4247 (N_4247,In_966,In_220);
or U4248 (N_4248,In_127,In_38);
nand U4249 (N_4249,In_1364,In_1494);
nor U4250 (N_4250,In_166,In_599);
nor U4251 (N_4251,In_404,In_542);
nor U4252 (N_4252,In_264,In_1087);
or U4253 (N_4253,In_1239,In_35);
nor U4254 (N_4254,In_1533,In_1630);
and U4255 (N_4255,In_795,In_617);
or U4256 (N_4256,In_1535,In_1057);
or U4257 (N_4257,In_1111,In_654);
or U4258 (N_4258,In_896,In_719);
or U4259 (N_4259,In_1451,In_1552);
nor U4260 (N_4260,In_870,In_1728);
and U4261 (N_4261,In_1644,In_643);
nor U4262 (N_4262,In_1288,In_102);
and U4263 (N_4263,In_1718,In_149);
nor U4264 (N_4264,In_933,In_829);
or U4265 (N_4265,In_202,In_199);
and U4266 (N_4266,In_1425,In_1992);
or U4267 (N_4267,In_1053,In_1331);
nand U4268 (N_4268,In_1782,In_1504);
and U4269 (N_4269,In_1968,In_1989);
nand U4270 (N_4270,In_203,In_1677);
or U4271 (N_4271,In_347,In_892);
nor U4272 (N_4272,In_1638,In_617);
and U4273 (N_4273,In_566,In_1097);
nor U4274 (N_4274,In_961,In_709);
xnor U4275 (N_4275,In_1407,In_1969);
nor U4276 (N_4276,In_1065,In_1528);
or U4277 (N_4277,In_1343,In_1936);
or U4278 (N_4278,In_1800,In_1606);
nor U4279 (N_4279,In_455,In_467);
nand U4280 (N_4280,In_642,In_672);
or U4281 (N_4281,In_1660,In_1624);
or U4282 (N_4282,In_1799,In_578);
or U4283 (N_4283,In_91,In_1255);
and U4284 (N_4284,In_1242,In_1299);
or U4285 (N_4285,In_356,In_1351);
and U4286 (N_4286,In_1159,In_460);
or U4287 (N_4287,In_1774,In_776);
nor U4288 (N_4288,In_85,In_1975);
nor U4289 (N_4289,In_1784,In_1675);
nand U4290 (N_4290,In_1273,In_1611);
or U4291 (N_4291,In_485,In_383);
and U4292 (N_4292,In_948,In_1813);
nand U4293 (N_4293,In_183,In_1073);
nand U4294 (N_4294,In_698,In_1115);
and U4295 (N_4295,In_894,In_755);
or U4296 (N_4296,In_397,In_711);
nand U4297 (N_4297,In_42,In_166);
and U4298 (N_4298,In_90,In_170);
nor U4299 (N_4299,In_635,In_1777);
nand U4300 (N_4300,In_869,In_476);
xnor U4301 (N_4301,In_532,In_1476);
nand U4302 (N_4302,In_576,In_980);
or U4303 (N_4303,In_1868,In_1854);
nand U4304 (N_4304,In_782,In_1461);
and U4305 (N_4305,In_920,In_1819);
or U4306 (N_4306,In_889,In_1401);
and U4307 (N_4307,In_565,In_1192);
or U4308 (N_4308,In_297,In_599);
nand U4309 (N_4309,In_1146,In_829);
xor U4310 (N_4310,In_1072,In_1745);
nand U4311 (N_4311,In_1347,In_160);
nor U4312 (N_4312,In_636,In_1817);
and U4313 (N_4313,In_1711,In_501);
nand U4314 (N_4314,In_386,In_310);
or U4315 (N_4315,In_1564,In_1981);
nor U4316 (N_4316,In_428,In_964);
and U4317 (N_4317,In_271,In_104);
and U4318 (N_4318,In_1996,In_1591);
and U4319 (N_4319,In_113,In_418);
nor U4320 (N_4320,In_1180,In_618);
or U4321 (N_4321,In_1908,In_1451);
nor U4322 (N_4322,In_171,In_1242);
nand U4323 (N_4323,In_113,In_1535);
nor U4324 (N_4324,In_1132,In_1473);
nand U4325 (N_4325,In_1957,In_418);
and U4326 (N_4326,In_283,In_1526);
and U4327 (N_4327,In_1259,In_38);
or U4328 (N_4328,In_684,In_1852);
and U4329 (N_4329,In_605,In_1828);
nor U4330 (N_4330,In_1701,In_1318);
nor U4331 (N_4331,In_926,In_658);
nand U4332 (N_4332,In_507,In_1392);
and U4333 (N_4333,In_1208,In_1661);
nand U4334 (N_4334,In_862,In_856);
nand U4335 (N_4335,In_434,In_1289);
nor U4336 (N_4336,In_244,In_1203);
or U4337 (N_4337,In_665,In_420);
nor U4338 (N_4338,In_1590,In_1708);
nand U4339 (N_4339,In_1757,In_1458);
nor U4340 (N_4340,In_1367,In_1004);
nand U4341 (N_4341,In_816,In_937);
nand U4342 (N_4342,In_503,In_1855);
nor U4343 (N_4343,In_206,In_128);
or U4344 (N_4344,In_985,In_1753);
nor U4345 (N_4345,In_193,In_1151);
or U4346 (N_4346,In_287,In_979);
and U4347 (N_4347,In_1380,In_455);
nor U4348 (N_4348,In_1954,In_589);
or U4349 (N_4349,In_1330,In_1421);
xor U4350 (N_4350,In_1696,In_1811);
or U4351 (N_4351,In_325,In_1339);
or U4352 (N_4352,In_1897,In_1157);
or U4353 (N_4353,In_157,In_1834);
and U4354 (N_4354,In_1566,In_407);
nand U4355 (N_4355,In_1853,In_985);
and U4356 (N_4356,In_300,In_41);
or U4357 (N_4357,In_899,In_285);
and U4358 (N_4358,In_945,In_996);
and U4359 (N_4359,In_678,In_618);
nor U4360 (N_4360,In_1437,In_1409);
nor U4361 (N_4361,In_1699,In_1164);
nor U4362 (N_4362,In_1097,In_303);
xnor U4363 (N_4363,In_926,In_367);
xnor U4364 (N_4364,In_290,In_1928);
or U4365 (N_4365,In_162,In_1032);
nor U4366 (N_4366,In_937,In_1003);
and U4367 (N_4367,In_1718,In_562);
and U4368 (N_4368,In_691,In_606);
and U4369 (N_4369,In_1964,In_644);
and U4370 (N_4370,In_807,In_233);
nand U4371 (N_4371,In_898,In_347);
or U4372 (N_4372,In_863,In_711);
nand U4373 (N_4373,In_594,In_1107);
or U4374 (N_4374,In_418,In_789);
nor U4375 (N_4375,In_1452,In_634);
nor U4376 (N_4376,In_1174,In_187);
and U4377 (N_4377,In_1368,In_502);
or U4378 (N_4378,In_1578,In_364);
nand U4379 (N_4379,In_1856,In_1494);
nor U4380 (N_4380,In_1381,In_203);
or U4381 (N_4381,In_1434,In_1206);
and U4382 (N_4382,In_1554,In_896);
or U4383 (N_4383,In_1360,In_1809);
nor U4384 (N_4384,In_557,In_1361);
nand U4385 (N_4385,In_1569,In_1211);
and U4386 (N_4386,In_1338,In_1395);
nor U4387 (N_4387,In_207,In_464);
nor U4388 (N_4388,In_6,In_661);
nand U4389 (N_4389,In_1311,In_1752);
and U4390 (N_4390,In_46,In_689);
nor U4391 (N_4391,In_821,In_1525);
or U4392 (N_4392,In_1272,In_1558);
nand U4393 (N_4393,In_1902,In_139);
nor U4394 (N_4394,In_1564,In_1311);
nand U4395 (N_4395,In_1134,In_1678);
nor U4396 (N_4396,In_199,In_1983);
and U4397 (N_4397,In_198,In_381);
nor U4398 (N_4398,In_619,In_1484);
nand U4399 (N_4399,In_454,In_1312);
or U4400 (N_4400,In_1170,In_994);
nor U4401 (N_4401,In_517,In_659);
nor U4402 (N_4402,In_375,In_865);
or U4403 (N_4403,In_515,In_869);
nand U4404 (N_4404,In_1772,In_1489);
nor U4405 (N_4405,In_1580,In_1343);
or U4406 (N_4406,In_1752,In_143);
nor U4407 (N_4407,In_1815,In_212);
nand U4408 (N_4408,In_1542,In_99);
or U4409 (N_4409,In_119,In_1552);
nor U4410 (N_4410,In_752,In_1488);
nand U4411 (N_4411,In_1303,In_402);
and U4412 (N_4412,In_921,In_412);
and U4413 (N_4413,In_182,In_1089);
nor U4414 (N_4414,In_1294,In_246);
and U4415 (N_4415,In_61,In_1982);
nor U4416 (N_4416,In_682,In_1517);
and U4417 (N_4417,In_1521,In_1124);
and U4418 (N_4418,In_1358,In_1901);
nand U4419 (N_4419,In_179,In_1983);
nor U4420 (N_4420,In_1093,In_1705);
nand U4421 (N_4421,In_1708,In_1110);
nor U4422 (N_4422,In_532,In_1647);
nand U4423 (N_4423,In_107,In_425);
or U4424 (N_4424,In_1505,In_1824);
or U4425 (N_4425,In_1721,In_1580);
and U4426 (N_4426,In_180,In_203);
nand U4427 (N_4427,In_733,In_822);
or U4428 (N_4428,In_61,In_513);
nor U4429 (N_4429,In_1184,In_169);
nor U4430 (N_4430,In_344,In_234);
or U4431 (N_4431,In_882,In_897);
nor U4432 (N_4432,In_1275,In_706);
and U4433 (N_4433,In_1117,In_441);
or U4434 (N_4434,In_1437,In_5);
and U4435 (N_4435,In_512,In_438);
nand U4436 (N_4436,In_1839,In_1040);
or U4437 (N_4437,In_1774,In_1893);
and U4438 (N_4438,In_696,In_1293);
and U4439 (N_4439,In_1141,In_1023);
and U4440 (N_4440,In_38,In_1715);
nor U4441 (N_4441,In_272,In_1427);
or U4442 (N_4442,In_733,In_1789);
nor U4443 (N_4443,In_1703,In_1165);
nand U4444 (N_4444,In_586,In_94);
nand U4445 (N_4445,In_1027,In_1750);
and U4446 (N_4446,In_400,In_841);
nand U4447 (N_4447,In_611,In_696);
xor U4448 (N_4448,In_409,In_243);
and U4449 (N_4449,In_253,In_18);
nor U4450 (N_4450,In_1332,In_295);
and U4451 (N_4451,In_685,In_1461);
nand U4452 (N_4452,In_649,In_1778);
or U4453 (N_4453,In_1230,In_573);
and U4454 (N_4454,In_1164,In_1065);
nand U4455 (N_4455,In_1251,In_94);
or U4456 (N_4456,In_1711,In_1345);
and U4457 (N_4457,In_466,In_1179);
nor U4458 (N_4458,In_1610,In_498);
nand U4459 (N_4459,In_1745,In_567);
or U4460 (N_4460,In_446,In_965);
nand U4461 (N_4461,In_285,In_898);
nand U4462 (N_4462,In_151,In_918);
nand U4463 (N_4463,In_214,In_1576);
or U4464 (N_4464,In_1415,In_1393);
nor U4465 (N_4465,In_1349,In_1256);
nor U4466 (N_4466,In_1292,In_1547);
nand U4467 (N_4467,In_973,In_1034);
and U4468 (N_4468,In_150,In_1440);
nor U4469 (N_4469,In_1610,In_315);
nor U4470 (N_4470,In_1142,In_669);
xnor U4471 (N_4471,In_1651,In_1862);
and U4472 (N_4472,In_28,In_245);
or U4473 (N_4473,In_1518,In_1730);
nand U4474 (N_4474,In_382,In_1750);
nand U4475 (N_4475,In_888,In_1999);
nand U4476 (N_4476,In_1081,In_1328);
or U4477 (N_4477,In_453,In_811);
nor U4478 (N_4478,In_80,In_1283);
nand U4479 (N_4479,In_653,In_1538);
nand U4480 (N_4480,In_1718,In_1630);
nor U4481 (N_4481,In_1538,In_1);
and U4482 (N_4482,In_1925,In_1077);
nor U4483 (N_4483,In_608,In_90);
or U4484 (N_4484,In_942,In_107);
nor U4485 (N_4485,In_781,In_1533);
nand U4486 (N_4486,In_365,In_1941);
nor U4487 (N_4487,In_1988,In_1773);
nand U4488 (N_4488,In_601,In_1018);
or U4489 (N_4489,In_1113,In_834);
nand U4490 (N_4490,In_800,In_1898);
nand U4491 (N_4491,In_191,In_382);
nor U4492 (N_4492,In_1044,In_184);
nand U4493 (N_4493,In_1318,In_529);
or U4494 (N_4494,In_1869,In_153);
and U4495 (N_4495,In_601,In_1684);
and U4496 (N_4496,In_213,In_1239);
and U4497 (N_4497,In_1773,In_31);
and U4498 (N_4498,In_1254,In_357);
nor U4499 (N_4499,In_1494,In_448);
and U4500 (N_4500,In_1243,In_1983);
xor U4501 (N_4501,In_840,In_212);
and U4502 (N_4502,In_586,In_907);
or U4503 (N_4503,In_1737,In_617);
or U4504 (N_4504,In_764,In_389);
nand U4505 (N_4505,In_133,In_948);
and U4506 (N_4506,In_420,In_718);
or U4507 (N_4507,In_417,In_471);
nor U4508 (N_4508,In_357,In_657);
nand U4509 (N_4509,In_1115,In_1235);
and U4510 (N_4510,In_1509,In_1877);
nand U4511 (N_4511,In_1264,In_1676);
and U4512 (N_4512,In_1031,In_1782);
or U4513 (N_4513,In_316,In_939);
nor U4514 (N_4514,In_1920,In_1855);
and U4515 (N_4515,In_1176,In_416);
and U4516 (N_4516,In_1262,In_1257);
nor U4517 (N_4517,In_1237,In_214);
nand U4518 (N_4518,In_1774,In_19);
nor U4519 (N_4519,In_289,In_1321);
and U4520 (N_4520,In_1115,In_1939);
nor U4521 (N_4521,In_1180,In_452);
nand U4522 (N_4522,In_1583,In_833);
nor U4523 (N_4523,In_100,In_257);
and U4524 (N_4524,In_1484,In_1924);
nand U4525 (N_4525,In_839,In_1755);
or U4526 (N_4526,In_1050,In_1072);
and U4527 (N_4527,In_600,In_437);
or U4528 (N_4528,In_2,In_1190);
nand U4529 (N_4529,In_681,In_1770);
or U4530 (N_4530,In_1117,In_81);
nor U4531 (N_4531,In_1454,In_37);
nand U4532 (N_4532,In_997,In_176);
nand U4533 (N_4533,In_762,In_127);
or U4534 (N_4534,In_247,In_846);
and U4535 (N_4535,In_1040,In_761);
and U4536 (N_4536,In_1808,In_873);
and U4537 (N_4537,In_1437,In_1679);
or U4538 (N_4538,In_861,In_1379);
and U4539 (N_4539,In_1330,In_1030);
nand U4540 (N_4540,In_669,In_613);
nor U4541 (N_4541,In_1019,In_1297);
nand U4542 (N_4542,In_1780,In_1009);
nor U4543 (N_4543,In_55,In_46);
nor U4544 (N_4544,In_1383,In_621);
nand U4545 (N_4545,In_1831,In_1761);
nand U4546 (N_4546,In_1625,In_1105);
nand U4547 (N_4547,In_1670,In_504);
and U4548 (N_4548,In_1469,In_939);
or U4549 (N_4549,In_1867,In_592);
nor U4550 (N_4550,In_1330,In_1692);
nor U4551 (N_4551,In_390,In_1649);
nor U4552 (N_4552,In_1578,In_1654);
or U4553 (N_4553,In_847,In_886);
nor U4554 (N_4554,In_1194,In_838);
nor U4555 (N_4555,In_1025,In_1705);
nor U4556 (N_4556,In_1487,In_1890);
nor U4557 (N_4557,In_189,In_1732);
nand U4558 (N_4558,In_854,In_1004);
and U4559 (N_4559,In_1679,In_630);
nand U4560 (N_4560,In_1701,In_928);
nor U4561 (N_4561,In_1789,In_1481);
or U4562 (N_4562,In_695,In_368);
nor U4563 (N_4563,In_1671,In_997);
and U4564 (N_4564,In_1525,In_156);
nor U4565 (N_4565,In_268,In_882);
and U4566 (N_4566,In_1500,In_1236);
nand U4567 (N_4567,In_457,In_829);
nor U4568 (N_4568,In_1906,In_614);
and U4569 (N_4569,In_690,In_592);
and U4570 (N_4570,In_1399,In_784);
nor U4571 (N_4571,In_1965,In_536);
or U4572 (N_4572,In_1392,In_1998);
or U4573 (N_4573,In_233,In_1840);
or U4574 (N_4574,In_599,In_1254);
and U4575 (N_4575,In_334,In_165);
and U4576 (N_4576,In_1491,In_1726);
and U4577 (N_4577,In_239,In_1487);
and U4578 (N_4578,In_1637,In_413);
or U4579 (N_4579,In_663,In_771);
and U4580 (N_4580,In_287,In_511);
nor U4581 (N_4581,In_1617,In_1581);
or U4582 (N_4582,In_1718,In_1365);
nand U4583 (N_4583,In_221,In_1016);
and U4584 (N_4584,In_263,In_1795);
and U4585 (N_4585,In_1295,In_1931);
or U4586 (N_4586,In_1330,In_1424);
or U4587 (N_4587,In_1761,In_604);
or U4588 (N_4588,In_1675,In_613);
xor U4589 (N_4589,In_1824,In_115);
nor U4590 (N_4590,In_625,In_1066);
or U4591 (N_4591,In_1747,In_869);
or U4592 (N_4592,In_995,In_462);
nand U4593 (N_4593,In_1317,In_692);
or U4594 (N_4594,In_898,In_1691);
or U4595 (N_4595,In_1254,In_1722);
and U4596 (N_4596,In_587,In_425);
and U4597 (N_4597,In_38,In_1137);
nand U4598 (N_4598,In_32,In_363);
or U4599 (N_4599,In_143,In_163);
nand U4600 (N_4600,In_706,In_37);
and U4601 (N_4601,In_681,In_310);
nand U4602 (N_4602,In_374,In_247);
or U4603 (N_4603,In_58,In_701);
nor U4604 (N_4604,In_1113,In_1220);
nor U4605 (N_4605,In_794,In_348);
nand U4606 (N_4606,In_1308,In_1356);
or U4607 (N_4607,In_1948,In_1495);
or U4608 (N_4608,In_827,In_182);
nor U4609 (N_4609,In_1077,In_828);
nor U4610 (N_4610,In_1647,In_713);
or U4611 (N_4611,In_1322,In_1673);
nand U4612 (N_4612,In_651,In_1932);
nand U4613 (N_4613,In_710,In_327);
nor U4614 (N_4614,In_1071,In_1925);
and U4615 (N_4615,In_1795,In_789);
or U4616 (N_4616,In_62,In_1805);
or U4617 (N_4617,In_1532,In_586);
nand U4618 (N_4618,In_1542,In_955);
nor U4619 (N_4619,In_1023,In_1197);
nor U4620 (N_4620,In_423,In_1468);
nor U4621 (N_4621,In_1239,In_1047);
nand U4622 (N_4622,In_756,In_604);
or U4623 (N_4623,In_1370,In_181);
nor U4624 (N_4624,In_204,In_1324);
or U4625 (N_4625,In_56,In_1344);
and U4626 (N_4626,In_171,In_1482);
nor U4627 (N_4627,In_460,In_776);
and U4628 (N_4628,In_1709,In_237);
nand U4629 (N_4629,In_380,In_1573);
nand U4630 (N_4630,In_806,In_1994);
or U4631 (N_4631,In_1968,In_1980);
or U4632 (N_4632,In_1852,In_1258);
and U4633 (N_4633,In_1977,In_1113);
nor U4634 (N_4634,In_1357,In_1274);
nand U4635 (N_4635,In_488,In_1707);
nand U4636 (N_4636,In_1240,In_23);
or U4637 (N_4637,In_1210,In_1312);
nand U4638 (N_4638,In_1499,In_1201);
or U4639 (N_4639,In_1851,In_22);
or U4640 (N_4640,In_602,In_283);
nand U4641 (N_4641,In_1150,In_768);
nand U4642 (N_4642,In_1717,In_1834);
and U4643 (N_4643,In_507,In_1006);
or U4644 (N_4644,In_1146,In_1818);
nor U4645 (N_4645,In_411,In_926);
nand U4646 (N_4646,In_363,In_1034);
or U4647 (N_4647,In_978,In_592);
nor U4648 (N_4648,In_1807,In_941);
nand U4649 (N_4649,In_1365,In_847);
nand U4650 (N_4650,In_486,In_62);
or U4651 (N_4651,In_258,In_815);
nor U4652 (N_4652,In_624,In_1643);
nor U4653 (N_4653,In_591,In_1336);
or U4654 (N_4654,In_1313,In_54);
nand U4655 (N_4655,In_1829,In_221);
or U4656 (N_4656,In_652,In_472);
or U4657 (N_4657,In_1312,In_513);
nand U4658 (N_4658,In_1050,In_148);
nand U4659 (N_4659,In_1500,In_1833);
or U4660 (N_4660,In_382,In_373);
and U4661 (N_4661,In_820,In_1719);
nand U4662 (N_4662,In_1796,In_1640);
and U4663 (N_4663,In_1036,In_1438);
and U4664 (N_4664,In_105,In_859);
or U4665 (N_4665,In_1090,In_824);
and U4666 (N_4666,In_314,In_141);
nor U4667 (N_4667,In_909,In_844);
or U4668 (N_4668,In_928,In_1356);
nor U4669 (N_4669,In_80,In_669);
nand U4670 (N_4670,In_1697,In_1943);
or U4671 (N_4671,In_67,In_1124);
or U4672 (N_4672,In_429,In_243);
or U4673 (N_4673,In_1265,In_1444);
nand U4674 (N_4674,In_1365,In_1899);
xor U4675 (N_4675,In_1310,In_1822);
nand U4676 (N_4676,In_1231,In_142);
nand U4677 (N_4677,In_925,In_759);
or U4678 (N_4678,In_541,In_1818);
and U4679 (N_4679,In_1170,In_1969);
or U4680 (N_4680,In_393,In_289);
and U4681 (N_4681,In_333,In_71);
nor U4682 (N_4682,In_74,In_370);
and U4683 (N_4683,In_1931,In_1617);
and U4684 (N_4684,In_1926,In_1478);
and U4685 (N_4685,In_758,In_1337);
or U4686 (N_4686,In_1914,In_611);
and U4687 (N_4687,In_1909,In_517);
nand U4688 (N_4688,In_742,In_339);
or U4689 (N_4689,In_1336,In_74);
nor U4690 (N_4690,In_1590,In_305);
xnor U4691 (N_4691,In_523,In_964);
nor U4692 (N_4692,In_1468,In_1823);
nand U4693 (N_4693,In_1705,In_976);
and U4694 (N_4694,In_1007,In_1260);
nor U4695 (N_4695,In_343,In_51);
or U4696 (N_4696,In_610,In_273);
nor U4697 (N_4697,In_1850,In_193);
nand U4698 (N_4698,In_55,In_540);
and U4699 (N_4699,In_695,In_326);
nand U4700 (N_4700,In_76,In_1591);
nor U4701 (N_4701,In_1409,In_410);
nor U4702 (N_4702,In_671,In_315);
nor U4703 (N_4703,In_1325,In_1454);
nand U4704 (N_4704,In_1892,In_1337);
nor U4705 (N_4705,In_1234,In_1388);
and U4706 (N_4706,In_950,In_914);
and U4707 (N_4707,In_1947,In_1194);
nand U4708 (N_4708,In_696,In_139);
and U4709 (N_4709,In_671,In_1715);
or U4710 (N_4710,In_1018,In_316);
and U4711 (N_4711,In_1227,In_172);
nor U4712 (N_4712,In_807,In_1866);
or U4713 (N_4713,In_938,In_596);
nand U4714 (N_4714,In_1434,In_31);
nor U4715 (N_4715,In_1287,In_1840);
nand U4716 (N_4716,In_764,In_155);
nor U4717 (N_4717,In_796,In_1210);
nor U4718 (N_4718,In_287,In_1529);
and U4719 (N_4719,In_621,In_1249);
nor U4720 (N_4720,In_181,In_1717);
or U4721 (N_4721,In_398,In_1151);
nand U4722 (N_4722,In_212,In_429);
nand U4723 (N_4723,In_1352,In_1952);
and U4724 (N_4724,In_697,In_326);
or U4725 (N_4725,In_365,In_780);
and U4726 (N_4726,In_1717,In_1917);
and U4727 (N_4727,In_1796,In_400);
and U4728 (N_4728,In_951,In_1753);
nand U4729 (N_4729,In_994,In_1893);
or U4730 (N_4730,In_1489,In_1418);
nand U4731 (N_4731,In_1689,In_360);
nand U4732 (N_4732,In_1572,In_1236);
nand U4733 (N_4733,In_1040,In_328);
or U4734 (N_4734,In_998,In_1323);
nand U4735 (N_4735,In_1566,In_1687);
or U4736 (N_4736,In_219,In_1795);
nand U4737 (N_4737,In_1272,In_1115);
nor U4738 (N_4738,In_1777,In_367);
or U4739 (N_4739,In_623,In_659);
or U4740 (N_4740,In_435,In_843);
and U4741 (N_4741,In_1919,In_1678);
nor U4742 (N_4742,In_1687,In_1843);
nand U4743 (N_4743,In_286,In_1188);
or U4744 (N_4744,In_13,In_112);
nor U4745 (N_4745,In_636,In_1261);
xor U4746 (N_4746,In_571,In_1709);
nand U4747 (N_4747,In_120,In_243);
nor U4748 (N_4748,In_1437,In_1045);
nor U4749 (N_4749,In_1303,In_1794);
and U4750 (N_4750,In_539,In_333);
nor U4751 (N_4751,In_821,In_897);
nor U4752 (N_4752,In_846,In_305);
nand U4753 (N_4753,In_1665,In_343);
nor U4754 (N_4754,In_1409,In_770);
and U4755 (N_4755,In_1649,In_789);
nand U4756 (N_4756,In_519,In_154);
nand U4757 (N_4757,In_1644,In_162);
or U4758 (N_4758,In_1503,In_1748);
nor U4759 (N_4759,In_1191,In_469);
and U4760 (N_4760,In_1343,In_349);
or U4761 (N_4761,In_133,In_1115);
and U4762 (N_4762,In_790,In_332);
nor U4763 (N_4763,In_384,In_1001);
or U4764 (N_4764,In_797,In_1604);
or U4765 (N_4765,In_746,In_202);
nor U4766 (N_4766,In_1051,In_1163);
and U4767 (N_4767,In_1706,In_275);
nand U4768 (N_4768,In_343,In_1710);
nor U4769 (N_4769,In_1925,In_1543);
nand U4770 (N_4770,In_29,In_1281);
nand U4771 (N_4771,In_1459,In_1441);
nand U4772 (N_4772,In_824,In_1039);
and U4773 (N_4773,In_1295,In_482);
nor U4774 (N_4774,In_1877,In_943);
nand U4775 (N_4775,In_1186,In_766);
nand U4776 (N_4776,In_988,In_1133);
and U4777 (N_4777,In_1799,In_705);
nand U4778 (N_4778,In_996,In_874);
nand U4779 (N_4779,In_151,In_1679);
and U4780 (N_4780,In_592,In_1695);
and U4781 (N_4781,In_1198,In_1210);
or U4782 (N_4782,In_1055,In_1575);
nor U4783 (N_4783,In_1619,In_154);
or U4784 (N_4784,In_1488,In_1992);
nor U4785 (N_4785,In_486,In_180);
nand U4786 (N_4786,In_1949,In_944);
nand U4787 (N_4787,In_808,In_1888);
nor U4788 (N_4788,In_647,In_627);
nand U4789 (N_4789,In_332,In_1914);
nor U4790 (N_4790,In_1440,In_845);
and U4791 (N_4791,In_778,In_910);
or U4792 (N_4792,In_1294,In_1743);
xor U4793 (N_4793,In_524,In_1788);
and U4794 (N_4794,In_1918,In_1331);
nand U4795 (N_4795,In_132,In_295);
nand U4796 (N_4796,In_1372,In_900);
or U4797 (N_4797,In_537,In_1997);
or U4798 (N_4798,In_123,In_971);
or U4799 (N_4799,In_830,In_927);
nand U4800 (N_4800,In_489,In_1772);
nor U4801 (N_4801,In_178,In_1450);
nand U4802 (N_4802,In_582,In_1682);
and U4803 (N_4803,In_944,In_1398);
or U4804 (N_4804,In_1961,In_306);
or U4805 (N_4805,In_1377,In_76);
nor U4806 (N_4806,In_1853,In_943);
and U4807 (N_4807,In_1121,In_1813);
or U4808 (N_4808,In_614,In_1392);
nor U4809 (N_4809,In_866,In_1699);
nand U4810 (N_4810,In_434,In_1792);
or U4811 (N_4811,In_1081,In_1586);
nor U4812 (N_4812,In_548,In_1748);
nor U4813 (N_4813,In_274,In_1541);
nor U4814 (N_4814,In_572,In_209);
and U4815 (N_4815,In_640,In_1538);
or U4816 (N_4816,In_1516,In_1520);
and U4817 (N_4817,In_349,In_1908);
nor U4818 (N_4818,In_1435,In_1948);
or U4819 (N_4819,In_574,In_1266);
or U4820 (N_4820,In_693,In_907);
nand U4821 (N_4821,In_441,In_948);
and U4822 (N_4822,In_199,In_1385);
and U4823 (N_4823,In_542,In_1815);
or U4824 (N_4824,In_579,In_1182);
nor U4825 (N_4825,In_1583,In_1939);
or U4826 (N_4826,In_1831,In_1416);
nand U4827 (N_4827,In_599,In_926);
nand U4828 (N_4828,In_367,In_1663);
nor U4829 (N_4829,In_728,In_1332);
nor U4830 (N_4830,In_1860,In_1561);
or U4831 (N_4831,In_1614,In_1386);
xnor U4832 (N_4832,In_1920,In_1418);
nand U4833 (N_4833,In_1644,In_1385);
or U4834 (N_4834,In_799,In_684);
xnor U4835 (N_4835,In_873,In_744);
nand U4836 (N_4836,In_1070,In_11);
and U4837 (N_4837,In_797,In_640);
and U4838 (N_4838,In_507,In_801);
nor U4839 (N_4839,In_995,In_1120);
or U4840 (N_4840,In_875,In_192);
xnor U4841 (N_4841,In_355,In_850);
nor U4842 (N_4842,In_1914,In_905);
and U4843 (N_4843,In_81,In_1184);
and U4844 (N_4844,In_74,In_1114);
or U4845 (N_4845,In_1107,In_72);
and U4846 (N_4846,In_1780,In_1104);
or U4847 (N_4847,In_1524,In_166);
nand U4848 (N_4848,In_1510,In_123);
or U4849 (N_4849,In_1228,In_190);
nand U4850 (N_4850,In_1811,In_1893);
or U4851 (N_4851,In_934,In_746);
or U4852 (N_4852,In_1639,In_721);
and U4853 (N_4853,In_1971,In_844);
nor U4854 (N_4854,In_1643,In_381);
nor U4855 (N_4855,In_274,In_847);
and U4856 (N_4856,In_402,In_1129);
nand U4857 (N_4857,In_1665,In_1731);
or U4858 (N_4858,In_872,In_1652);
nor U4859 (N_4859,In_215,In_1418);
or U4860 (N_4860,In_1664,In_1372);
nand U4861 (N_4861,In_1993,In_1983);
or U4862 (N_4862,In_1082,In_1603);
xnor U4863 (N_4863,In_122,In_999);
nor U4864 (N_4864,In_416,In_634);
and U4865 (N_4865,In_87,In_964);
nor U4866 (N_4866,In_1054,In_127);
nand U4867 (N_4867,In_1318,In_991);
nor U4868 (N_4868,In_1430,In_1605);
or U4869 (N_4869,In_1394,In_1073);
nand U4870 (N_4870,In_1541,In_416);
or U4871 (N_4871,In_323,In_1321);
or U4872 (N_4872,In_1873,In_433);
nor U4873 (N_4873,In_1060,In_1191);
nor U4874 (N_4874,In_657,In_722);
nand U4875 (N_4875,In_854,In_74);
and U4876 (N_4876,In_1303,In_44);
nand U4877 (N_4877,In_1924,In_1792);
nand U4878 (N_4878,In_1570,In_1510);
nand U4879 (N_4879,In_635,In_1065);
or U4880 (N_4880,In_1161,In_653);
nor U4881 (N_4881,In_993,In_470);
nor U4882 (N_4882,In_403,In_693);
and U4883 (N_4883,In_1701,In_411);
nor U4884 (N_4884,In_971,In_611);
nand U4885 (N_4885,In_655,In_1373);
nand U4886 (N_4886,In_734,In_1767);
or U4887 (N_4887,In_1106,In_302);
or U4888 (N_4888,In_1582,In_273);
and U4889 (N_4889,In_972,In_1146);
xnor U4890 (N_4890,In_1257,In_99);
nor U4891 (N_4891,In_1750,In_817);
and U4892 (N_4892,In_974,In_483);
nor U4893 (N_4893,In_226,In_69);
and U4894 (N_4894,In_1138,In_97);
nand U4895 (N_4895,In_805,In_1804);
nor U4896 (N_4896,In_702,In_1320);
nor U4897 (N_4897,In_1229,In_1953);
and U4898 (N_4898,In_181,In_639);
and U4899 (N_4899,In_122,In_175);
and U4900 (N_4900,In_724,In_1639);
and U4901 (N_4901,In_1666,In_1183);
or U4902 (N_4902,In_500,In_1802);
nand U4903 (N_4903,In_867,In_264);
nor U4904 (N_4904,In_336,In_1127);
nor U4905 (N_4905,In_423,In_1739);
and U4906 (N_4906,In_1160,In_305);
and U4907 (N_4907,In_15,In_818);
nand U4908 (N_4908,In_456,In_760);
or U4909 (N_4909,In_368,In_350);
xnor U4910 (N_4910,In_73,In_44);
or U4911 (N_4911,In_735,In_1585);
and U4912 (N_4912,In_1729,In_397);
or U4913 (N_4913,In_1267,In_1689);
nor U4914 (N_4914,In_434,In_1856);
or U4915 (N_4915,In_1704,In_1778);
nor U4916 (N_4916,In_1112,In_268);
nor U4917 (N_4917,In_955,In_1470);
and U4918 (N_4918,In_1592,In_508);
nor U4919 (N_4919,In_313,In_809);
and U4920 (N_4920,In_1068,In_424);
nand U4921 (N_4921,In_1013,In_1080);
and U4922 (N_4922,In_1184,In_645);
nor U4923 (N_4923,In_1723,In_1951);
or U4924 (N_4924,In_171,In_1081);
nand U4925 (N_4925,In_344,In_485);
nor U4926 (N_4926,In_1915,In_747);
or U4927 (N_4927,In_1919,In_954);
or U4928 (N_4928,In_1429,In_0);
and U4929 (N_4929,In_1877,In_549);
and U4930 (N_4930,In_1211,In_1103);
and U4931 (N_4931,In_396,In_1853);
nor U4932 (N_4932,In_1630,In_1784);
and U4933 (N_4933,In_397,In_36);
or U4934 (N_4934,In_340,In_1164);
or U4935 (N_4935,In_228,In_1027);
and U4936 (N_4936,In_8,In_1055);
nand U4937 (N_4937,In_1831,In_889);
or U4938 (N_4938,In_1149,In_880);
or U4939 (N_4939,In_1312,In_263);
nor U4940 (N_4940,In_809,In_1079);
nor U4941 (N_4941,In_1948,In_1505);
or U4942 (N_4942,In_676,In_386);
and U4943 (N_4943,In_974,In_880);
nand U4944 (N_4944,In_548,In_1070);
or U4945 (N_4945,In_900,In_183);
nor U4946 (N_4946,In_1534,In_1171);
or U4947 (N_4947,In_1042,In_39);
nand U4948 (N_4948,In_718,In_1666);
nor U4949 (N_4949,In_439,In_1567);
nor U4950 (N_4950,In_1528,In_488);
or U4951 (N_4951,In_595,In_1171);
and U4952 (N_4952,In_175,In_954);
or U4953 (N_4953,In_1349,In_1678);
nand U4954 (N_4954,In_46,In_1402);
nand U4955 (N_4955,In_1556,In_1042);
nor U4956 (N_4956,In_1343,In_1786);
nor U4957 (N_4957,In_1887,In_1044);
nor U4958 (N_4958,In_876,In_1249);
or U4959 (N_4959,In_167,In_896);
and U4960 (N_4960,In_1016,In_910);
nand U4961 (N_4961,In_445,In_1968);
nand U4962 (N_4962,In_1220,In_1262);
nor U4963 (N_4963,In_1029,In_298);
xor U4964 (N_4964,In_1681,In_1000);
nand U4965 (N_4965,In_646,In_21);
nand U4966 (N_4966,In_1262,In_963);
or U4967 (N_4967,In_604,In_913);
and U4968 (N_4968,In_1217,In_1086);
and U4969 (N_4969,In_880,In_1319);
or U4970 (N_4970,In_1483,In_1202);
nand U4971 (N_4971,In_627,In_1041);
nor U4972 (N_4972,In_1942,In_1999);
nand U4973 (N_4973,In_575,In_231);
xnor U4974 (N_4974,In_1783,In_71);
nor U4975 (N_4975,In_72,In_686);
nor U4976 (N_4976,In_957,In_492);
nor U4977 (N_4977,In_404,In_1837);
nand U4978 (N_4978,In_1270,In_1768);
or U4979 (N_4979,In_1428,In_1771);
or U4980 (N_4980,In_974,In_1359);
or U4981 (N_4981,In_314,In_1414);
nand U4982 (N_4982,In_1102,In_1498);
nand U4983 (N_4983,In_730,In_635);
and U4984 (N_4984,In_437,In_127);
nor U4985 (N_4985,In_1832,In_653);
nand U4986 (N_4986,In_674,In_192);
nor U4987 (N_4987,In_1299,In_305);
or U4988 (N_4988,In_1719,In_1855);
and U4989 (N_4989,In_179,In_1600);
and U4990 (N_4990,In_1374,In_1902);
nand U4991 (N_4991,In_1195,In_761);
nand U4992 (N_4992,In_1011,In_2);
nand U4993 (N_4993,In_971,In_1866);
or U4994 (N_4994,In_1706,In_115);
nand U4995 (N_4995,In_638,In_1029);
and U4996 (N_4996,In_1965,In_1525);
or U4997 (N_4997,In_1652,In_1052);
or U4998 (N_4998,In_1011,In_1662);
nor U4999 (N_4999,In_529,In_1054);
nand U5000 (N_5000,N_41,N_708);
nor U5001 (N_5001,N_4500,N_2287);
and U5002 (N_5002,N_1147,N_3308);
and U5003 (N_5003,N_2925,N_4310);
or U5004 (N_5004,N_4198,N_3728);
or U5005 (N_5005,N_4559,N_1953);
or U5006 (N_5006,N_418,N_2856);
nand U5007 (N_5007,N_2327,N_2362);
nor U5008 (N_5008,N_399,N_4738);
nand U5009 (N_5009,N_3012,N_468);
or U5010 (N_5010,N_900,N_4524);
or U5011 (N_5011,N_74,N_1739);
nor U5012 (N_5012,N_1322,N_1639);
nand U5013 (N_5013,N_40,N_2740);
nand U5014 (N_5014,N_4272,N_3478);
and U5015 (N_5015,N_3972,N_4718);
nor U5016 (N_5016,N_3790,N_3178);
or U5017 (N_5017,N_4337,N_2315);
or U5018 (N_5018,N_727,N_58);
nand U5019 (N_5019,N_454,N_1348);
nor U5020 (N_5020,N_4857,N_389);
nor U5021 (N_5021,N_4065,N_3207);
or U5022 (N_5022,N_1551,N_1959);
nor U5023 (N_5023,N_4583,N_4465);
or U5024 (N_5024,N_3668,N_17);
and U5025 (N_5025,N_2797,N_2804);
or U5026 (N_5026,N_2401,N_4746);
and U5027 (N_5027,N_3936,N_4810);
and U5028 (N_5028,N_3442,N_209);
nand U5029 (N_5029,N_4792,N_3887);
nor U5030 (N_5030,N_4029,N_2744);
nand U5031 (N_5031,N_2483,N_2523);
nor U5032 (N_5032,N_3835,N_1766);
nand U5033 (N_5033,N_2558,N_4459);
and U5034 (N_5034,N_4182,N_1400);
nor U5035 (N_5035,N_4507,N_2695);
nand U5036 (N_5036,N_375,N_382);
and U5037 (N_5037,N_1564,N_1656);
nor U5038 (N_5038,N_1346,N_4160);
nand U5039 (N_5039,N_3256,N_3624);
nand U5040 (N_5040,N_4973,N_2490);
and U5041 (N_5041,N_110,N_612);
or U5042 (N_5042,N_506,N_398);
nand U5043 (N_5043,N_3919,N_4052);
and U5044 (N_5044,N_2493,N_4613);
or U5045 (N_5045,N_3409,N_2444);
nor U5046 (N_5046,N_1485,N_4118);
and U5047 (N_5047,N_1506,N_324);
and U5048 (N_5048,N_2267,N_4388);
nand U5049 (N_5049,N_4868,N_2606);
or U5050 (N_5050,N_1242,N_2528);
and U5051 (N_5051,N_899,N_2424);
or U5052 (N_5052,N_2369,N_2177);
or U5053 (N_5053,N_2752,N_1516);
or U5054 (N_5054,N_4938,N_1978);
nand U5055 (N_5055,N_96,N_1100);
or U5056 (N_5056,N_66,N_2978);
or U5057 (N_5057,N_689,N_3038);
or U5058 (N_5058,N_503,N_4887);
nand U5059 (N_5059,N_3385,N_1889);
or U5060 (N_5060,N_3903,N_2847);
or U5061 (N_5061,N_812,N_2060);
nand U5062 (N_5062,N_1136,N_3413);
nand U5063 (N_5063,N_917,N_3736);
and U5064 (N_5064,N_4414,N_488);
nor U5065 (N_5065,N_1626,N_122);
nand U5066 (N_5066,N_576,N_1713);
and U5067 (N_5067,N_2828,N_1880);
and U5068 (N_5068,N_825,N_3960);
and U5069 (N_5069,N_4540,N_4333);
or U5070 (N_5070,N_3269,N_587);
and U5071 (N_5071,N_68,N_3040);
and U5072 (N_5072,N_1772,N_477);
nand U5073 (N_5073,N_3306,N_244);
nor U5074 (N_5074,N_3904,N_4428);
nor U5075 (N_5075,N_712,N_307);
or U5076 (N_5076,N_1567,N_2090);
nand U5077 (N_5077,N_410,N_4783);
xor U5078 (N_5078,N_1177,N_2512);
or U5079 (N_5079,N_891,N_139);
or U5080 (N_5080,N_2015,N_3803);
nor U5081 (N_5081,N_4297,N_4257);
and U5082 (N_5082,N_730,N_3459);
nor U5083 (N_5083,N_2831,N_1861);
or U5084 (N_5084,N_2049,N_889);
nand U5085 (N_5085,N_3174,N_502);
nand U5086 (N_5086,N_3161,N_43);
nand U5087 (N_5087,N_1935,N_4377);
and U5088 (N_5088,N_1795,N_4822);
or U5089 (N_5089,N_4349,N_2076);
or U5090 (N_5090,N_3741,N_1926);
nor U5091 (N_5091,N_1972,N_2452);
or U5092 (N_5092,N_2781,N_759);
nand U5093 (N_5093,N_1513,N_2890);
nor U5094 (N_5094,N_572,N_844);
or U5095 (N_5095,N_4749,N_4617);
and U5096 (N_5096,N_1051,N_950);
or U5097 (N_5097,N_4867,N_4237);
nor U5098 (N_5098,N_3110,N_2999);
nand U5099 (N_5099,N_3824,N_4138);
and U5100 (N_5100,N_4744,N_1759);
and U5101 (N_5101,N_733,N_141);
nor U5102 (N_5102,N_811,N_2190);
or U5103 (N_5103,N_1503,N_3751);
and U5104 (N_5104,N_3495,N_4979);
xor U5105 (N_5105,N_2281,N_2866);
nand U5106 (N_5106,N_3299,N_1356);
nand U5107 (N_5107,N_872,N_3830);
nand U5108 (N_5108,N_2078,N_813);
nor U5109 (N_5109,N_4233,N_2586);
nand U5110 (N_5110,N_2485,N_510);
and U5111 (N_5111,N_2081,N_3928);
and U5112 (N_5112,N_4195,N_1657);
nand U5113 (N_5113,N_540,N_764);
nand U5114 (N_5114,N_3358,N_1716);
nand U5115 (N_5115,N_4519,N_2111);
nor U5116 (N_5116,N_4274,N_1520);
nand U5117 (N_5117,N_4823,N_1291);
or U5118 (N_5118,N_3967,N_4485);
or U5119 (N_5119,N_3193,N_4186);
nand U5120 (N_5120,N_4036,N_3220);
and U5121 (N_5121,N_2768,N_884);
nor U5122 (N_5122,N_284,N_1612);
or U5123 (N_5123,N_2141,N_1080);
or U5124 (N_5124,N_4134,N_1295);
and U5125 (N_5125,N_3167,N_4099);
nand U5126 (N_5126,N_3428,N_990);
nor U5127 (N_5127,N_2554,N_2378);
or U5128 (N_5128,N_4703,N_3056);
and U5129 (N_5129,N_1003,N_586);
and U5130 (N_5130,N_2535,N_634);
nor U5131 (N_5131,N_1034,N_3147);
nor U5132 (N_5132,N_600,N_4173);
or U5133 (N_5133,N_1509,N_3411);
or U5134 (N_5134,N_4796,N_456);
nor U5135 (N_5135,N_2165,N_1575);
and U5136 (N_5136,N_4102,N_1380);
nand U5137 (N_5137,N_2318,N_1462);
nand U5138 (N_5138,N_2114,N_36);
nor U5139 (N_5139,N_3732,N_2214);
nor U5140 (N_5140,N_2537,N_4053);
nor U5141 (N_5141,N_3241,N_3456);
nand U5142 (N_5142,N_1860,N_2839);
and U5143 (N_5143,N_4714,N_2851);
nor U5144 (N_5144,N_408,N_1001);
nor U5145 (N_5145,N_1667,N_3700);
nand U5146 (N_5146,N_3592,N_2749);
nand U5147 (N_5147,N_2548,N_2718);
nand U5148 (N_5148,N_896,N_4832);
nor U5149 (N_5149,N_3807,N_4410);
or U5150 (N_5150,N_1311,N_4244);
nand U5151 (N_5151,N_479,N_1105);
nand U5152 (N_5152,N_3452,N_2331);
and U5153 (N_5153,N_2805,N_534);
nor U5154 (N_5154,N_533,N_1222);
and U5155 (N_5155,N_2745,N_2320);
and U5156 (N_5156,N_3627,N_2884);
or U5157 (N_5157,N_3543,N_2024);
or U5158 (N_5158,N_2158,N_121);
and U5159 (N_5159,N_939,N_839);
or U5160 (N_5160,N_2034,N_3432);
and U5161 (N_5161,N_3712,N_1542);
or U5162 (N_5162,N_3158,N_3378);
nor U5163 (N_5163,N_2373,N_4022);
nand U5164 (N_5164,N_341,N_1533);
or U5165 (N_5165,N_3572,N_1473);
or U5166 (N_5166,N_3343,N_4179);
nor U5167 (N_5167,N_4123,N_1908);
nor U5168 (N_5168,N_3076,N_1998);
nor U5169 (N_5169,N_2511,N_329);
nand U5170 (N_5170,N_3801,N_752);
nand U5171 (N_5171,N_4656,N_911);
or U5172 (N_5172,N_1009,N_1176);
and U5173 (N_5173,N_1951,N_2432);
or U5174 (N_5174,N_1298,N_2868);
nand U5175 (N_5175,N_3598,N_471);
and U5176 (N_5176,N_535,N_613);
nand U5177 (N_5177,N_627,N_34);
nor U5178 (N_5178,N_304,N_4340);
nand U5179 (N_5179,N_625,N_3516);
nor U5180 (N_5180,N_3840,N_1099);
nor U5181 (N_5181,N_1022,N_4861);
nor U5182 (N_5182,N_3705,N_2118);
or U5183 (N_5183,N_2365,N_1749);
and U5184 (N_5184,N_4983,N_1263);
nor U5185 (N_5185,N_430,N_2233);
and U5186 (N_5186,N_2889,N_4026);
and U5187 (N_5187,N_832,N_4343);
and U5188 (N_5188,N_660,N_4227);
nor U5189 (N_5189,N_1026,N_303);
and U5190 (N_5190,N_3953,N_4907);
and U5191 (N_5191,N_4927,N_4460);
nand U5192 (N_5192,N_3512,N_2599);
nand U5193 (N_5193,N_4416,N_2017);
or U5194 (N_5194,N_2492,N_3978);
nand U5195 (N_5195,N_2617,N_1011);
or U5196 (N_5196,N_3657,N_1056);
nor U5197 (N_5197,N_2882,N_317);
nor U5198 (N_5198,N_3695,N_3421);
or U5199 (N_5199,N_1521,N_4178);
nand U5200 (N_5200,N_1044,N_1832);
nor U5201 (N_5201,N_3743,N_4588);
nand U5202 (N_5202,N_3944,N_365);
and U5203 (N_5203,N_658,N_4710);
nand U5204 (N_5204,N_871,N_2035);
or U5205 (N_5205,N_3414,N_2992);
or U5206 (N_5206,N_357,N_2756);
or U5207 (N_5207,N_1031,N_1901);
nor U5208 (N_5208,N_3877,N_1801);
and U5209 (N_5209,N_4968,N_3001);
and U5210 (N_5210,N_2443,N_895);
nor U5211 (N_5211,N_3286,N_1725);
or U5212 (N_5212,N_1124,N_1215);
nand U5213 (N_5213,N_4042,N_2008);
and U5214 (N_5214,N_2569,N_3727);
and U5215 (N_5215,N_4715,N_1275);
nor U5216 (N_5216,N_1864,N_519);
nor U5217 (N_5217,N_1399,N_1198);
nor U5218 (N_5218,N_1108,N_3433);
and U5219 (N_5219,N_1386,N_33);
nor U5220 (N_5220,N_308,N_4466);
and U5221 (N_5221,N_3121,N_1777);
and U5222 (N_5222,N_1754,N_2716);
or U5223 (N_5223,N_145,N_2089);
nand U5224 (N_5224,N_3391,N_646);
nand U5225 (N_5225,N_1878,N_1942);
and U5226 (N_5226,N_1152,N_2830);
nor U5227 (N_5227,N_72,N_3331);
nor U5228 (N_5228,N_4276,N_3329);
and U5229 (N_5229,N_1774,N_1184);
or U5230 (N_5230,N_3262,N_269);
or U5231 (N_5231,N_2607,N_311);
nand U5232 (N_5232,N_492,N_4578);
or U5233 (N_5233,N_1599,N_669);
nor U5234 (N_5234,N_3218,N_4152);
or U5235 (N_5235,N_4669,N_3441);
and U5236 (N_5236,N_273,N_3896);
or U5237 (N_5237,N_2396,N_2213);
nand U5238 (N_5238,N_4113,N_1094);
nor U5239 (N_5239,N_3263,N_1363);
or U5240 (N_5240,N_2074,N_1057);
or U5241 (N_5241,N_4797,N_4862);
nor U5242 (N_5242,N_2042,N_2522);
or U5243 (N_5243,N_2789,N_2926);
and U5244 (N_5244,N_4158,N_670);
nor U5245 (N_5245,N_1893,N_491);
nand U5246 (N_5246,N_4811,N_4933);
and U5247 (N_5247,N_2225,N_496);
nor U5248 (N_5248,N_306,N_4441);
nand U5249 (N_5249,N_3231,N_1272);
or U5250 (N_5250,N_2229,N_4708);
nor U5251 (N_5251,N_87,N_3011);
nand U5252 (N_5252,N_3104,N_4433);
nor U5253 (N_5253,N_803,N_4269);
nor U5254 (N_5254,N_1494,N_3485);
nand U5255 (N_5255,N_743,N_2767);
nand U5256 (N_5256,N_1091,N_4896);
and U5257 (N_5257,N_4334,N_3984);
or U5258 (N_5258,N_3142,N_2426);
and U5259 (N_5259,N_2096,N_4328);
nor U5260 (N_5260,N_2525,N_3622);
nor U5261 (N_5261,N_421,N_469);
nand U5262 (N_5262,N_1426,N_4000);
nand U5263 (N_5263,N_4883,N_4982);
and U5264 (N_5264,N_937,N_1857);
nor U5265 (N_5265,N_2397,N_3791);
nand U5266 (N_5266,N_3025,N_1151);
nand U5267 (N_5267,N_964,N_3515);
and U5268 (N_5268,N_2316,N_725);
or U5269 (N_5269,N_1512,N_155);
nor U5270 (N_5270,N_3044,N_3628);
or U5271 (N_5271,N_4697,N_2025);
nand U5272 (N_5272,N_980,N_3188);
or U5273 (N_5273,N_1197,N_4590);
or U5274 (N_5274,N_299,N_4087);
and U5275 (N_5275,N_509,N_2390);
nand U5276 (N_5276,N_4643,N_1069);
nor U5277 (N_5277,N_4322,N_2314);
or U5278 (N_5278,N_256,N_4112);
nor U5279 (N_5279,N_3612,N_3711);
nor U5280 (N_5280,N_583,N_787);
nor U5281 (N_5281,N_4769,N_4060);
nand U5282 (N_5282,N_628,N_2033);
nor U5283 (N_5283,N_2794,N_4183);
or U5284 (N_5284,N_3879,N_4326);
nor U5285 (N_5285,N_2590,N_2960);
nand U5286 (N_5286,N_4737,N_2787);
or U5287 (N_5287,N_279,N_4775);
nor U5288 (N_5288,N_2971,N_1032);
and U5289 (N_5289,N_4603,N_2986);
nand U5290 (N_5290,N_3394,N_2904);
nor U5291 (N_5291,N_2997,N_3046);
or U5292 (N_5292,N_2109,N_4365);
nand U5293 (N_5293,N_4128,N_629);
or U5294 (N_5294,N_4437,N_3006);
nand U5295 (N_5295,N_1737,N_1427);
nor U5296 (N_5296,N_4920,N_2625);
nand U5297 (N_5297,N_4033,N_2638);
or U5298 (N_5298,N_53,N_3560);
nor U5299 (N_5299,N_3393,N_741);
nor U5300 (N_5300,N_425,N_3533);
or U5301 (N_5301,N_2338,N_3914);
and U5302 (N_5302,N_3386,N_1540);
nor U5303 (N_5303,N_3435,N_1876);
or U5304 (N_5304,N_3664,N_223);
nor U5305 (N_5305,N_4536,N_1392);
nand U5306 (N_5306,N_3647,N_1405);
nor U5307 (N_5307,N_4230,N_478);
nor U5308 (N_5308,N_3809,N_3603);
nor U5309 (N_5309,N_2572,N_1681);
and U5310 (N_5310,N_3125,N_4374);
nand U5311 (N_5311,N_3725,N_1345);
and U5312 (N_5312,N_626,N_4597);
or U5313 (N_5313,N_1852,N_2179);
nand U5314 (N_5314,N_930,N_236);
nor U5315 (N_5315,N_4552,N_580);
or U5316 (N_5316,N_618,N_1634);
nor U5317 (N_5317,N_3945,N_3510);
and U5318 (N_5318,N_277,N_361);
nand U5319 (N_5319,N_1622,N_4948);
and U5320 (N_5320,N_3010,N_3768);
nor U5321 (N_5321,N_4172,N_1382);
nand U5322 (N_5322,N_4440,N_3307);
and U5323 (N_5323,N_1178,N_1803);
or U5324 (N_5324,N_3030,N_4355);
nor U5325 (N_5325,N_2352,N_2888);
and U5326 (N_5326,N_489,N_4457);
and U5327 (N_5327,N_2878,N_4580);
and U5328 (N_5328,N_1007,N_2463);
nand U5329 (N_5329,N_1378,N_562);
nand U5330 (N_5330,N_2310,N_3986);
nor U5331 (N_5331,N_3527,N_4111);
and U5332 (N_5332,N_4692,N_4455);
nor U5333 (N_5333,N_3183,N_107);
or U5334 (N_5334,N_4731,N_4288);
or U5335 (N_5335,N_568,N_2486);
and U5336 (N_5336,N_2726,N_1219);
nor U5337 (N_5337,N_2880,N_1074);
or U5338 (N_5338,N_4924,N_3399);
nor U5339 (N_5339,N_176,N_1922);
and U5340 (N_5340,N_3078,N_245);
and U5341 (N_5341,N_2095,N_2683);
nor U5342 (N_5342,N_2429,N_4311);
or U5343 (N_5343,N_1186,N_3004);
and U5344 (N_5344,N_3426,N_2050);
nand U5345 (N_5345,N_2143,N_2786);
or U5346 (N_5346,N_3818,N_154);
nor U5347 (N_5347,N_3999,N_2791);
or U5348 (N_5348,N_958,N_2083);
nor U5349 (N_5349,N_1967,N_4481);
nand U5350 (N_5350,N_386,N_3787);
and U5351 (N_5351,N_2404,N_4280);
nand U5352 (N_5352,N_3720,N_1562);
nor U5353 (N_5353,N_965,N_131);
nand U5354 (N_5354,N_1471,N_757);
and U5355 (N_5355,N_2510,N_855);
and U5356 (N_5356,N_4035,N_546);
or U5357 (N_5357,N_4001,N_359);
nor U5358 (N_5358,N_2296,N_728);
or U5359 (N_5359,N_1897,N_3245);
or U5360 (N_5360,N_1297,N_3446);
and U5361 (N_5361,N_3529,N_3095);
and U5362 (N_5362,N_1835,N_3785);
or U5363 (N_5363,N_1673,N_4772);
nor U5364 (N_5364,N_758,N_152);
nor U5365 (N_5365,N_4962,N_1456);
nor U5366 (N_5366,N_2005,N_1588);
and U5367 (N_5367,N_619,N_1005);
and U5368 (N_5368,N_1847,N_1255);
nand U5369 (N_5369,N_4729,N_3205);
or U5370 (N_5370,N_3,N_4259);
nor U5371 (N_5371,N_4814,N_4495);
or U5372 (N_5372,N_2923,N_3609);
or U5373 (N_5373,N_3092,N_207);
xor U5374 (N_5374,N_1885,N_2843);
nand U5375 (N_5375,N_4425,N_4287);
nor U5376 (N_5376,N_4961,N_4030);
nor U5377 (N_5377,N_2000,N_1243);
or U5378 (N_5378,N_104,N_156);
nor U5379 (N_5379,N_1154,N_2755);
nand U5380 (N_5380,N_1790,N_2680);
nor U5381 (N_5381,N_2441,N_696);
nand U5382 (N_5382,N_621,N_3355);
nand U5383 (N_5383,N_853,N_1609);
and U5384 (N_5384,N_9,N_2280);
and U5385 (N_5385,N_523,N_4126);
nand U5386 (N_5386,N_1067,N_1507);
nand U5387 (N_5387,N_4479,N_4594);
nand U5388 (N_5388,N_734,N_4252);
nand U5389 (N_5389,N_4864,N_1684);
or U5390 (N_5390,N_545,N_1413);
and U5391 (N_5391,N_3596,N_2700);
and U5392 (N_5392,N_4127,N_2153);
nand U5393 (N_5393,N_1979,N_2527);
nor U5394 (N_5394,N_3623,N_158);
or U5395 (N_5395,N_1496,N_2023);
nor U5396 (N_5396,N_2466,N_3767);
nand U5397 (N_5397,N_4409,N_3739);
and U5398 (N_5398,N_1407,N_1251);
and U5399 (N_5399,N_3156,N_3671);
or U5400 (N_5400,N_2711,N_3150);
or U5401 (N_5401,N_1931,N_3918);
nand U5402 (N_5402,N_2907,N_1203);
nor U5403 (N_5403,N_2857,N_3293);
and U5404 (N_5404,N_1472,N_674);
nand U5405 (N_5405,N_2,N_2655);
nand U5406 (N_5406,N_1334,N_3539);
nand U5407 (N_5407,N_3105,N_2210);
nor U5408 (N_5408,N_4503,N_4599);
nand U5409 (N_5409,N_4665,N_4967);
nand U5410 (N_5410,N_883,N_3228);
or U5411 (N_5411,N_3261,N_3356);
nand U5412 (N_5412,N_2286,N_1464);
nor U5413 (N_5413,N_2136,N_3017);
nor U5414 (N_5414,N_4605,N_4068);
nor U5415 (N_5415,N_3766,N_2021);
and U5416 (N_5416,N_4490,N_1581);
nor U5417 (N_5417,N_406,N_711);
and U5418 (N_5418,N_1064,N_906);
or U5419 (N_5419,N_925,N_3362);
or U5420 (N_5420,N_2909,N_162);
nor U5421 (N_5421,N_3534,N_4284);
nor U5422 (N_5422,N_3828,N_3200);
or U5423 (N_5423,N_2826,N_3584);
and U5424 (N_5424,N_3496,N_4830);
or U5425 (N_5425,N_1220,N_1404);
nand U5426 (N_5426,N_1989,N_2657);
nor U5427 (N_5427,N_1875,N_642);
and U5428 (N_5428,N_902,N_1349);
and U5429 (N_5429,N_391,N_1693);
and U5430 (N_5430,N_2254,N_1361);
nand U5431 (N_5431,N_4002,N_3058);
and U5432 (N_5432,N_4494,N_3112);
nand U5433 (N_5433,N_4105,N_1580);
nor U5434 (N_5434,N_1528,N_4820);
or U5435 (N_5435,N_544,N_2272);
and U5436 (N_5436,N_3649,N_3471);
and U5437 (N_5437,N_684,N_1752);
xor U5438 (N_5438,N_1325,N_1577);
and U5439 (N_5439,N_2253,N_3157);
nor U5440 (N_5440,N_1422,N_638);
nand U5441 (N_5441,N_1711,N_2499);
nand U5442 (N_5442,N_3748,N_2829);
or U5443 (N_5443,N_1375,N_3244);
nand U5444 (N_5444,N_4641,N_3694);
nand U5445 (N_5445,N_3651,N_2354);
or U5446 (N_5446,N_3875,N_440);
and U5447 (N_5447,N_1585,N_3611);
or U5448 (N_5448,N_1663,N_3804);
or U5449 (N_5449,N_3648,N_1715);
nor U5450 (N_5450,N_4696,N_2104);
and U5451 (N_5451,N_1319,N_4194);
and U5452 (N_5452,N_2113,N_1850);
nand U5453 (N_5453,N_718,N_717);
nor U5454 (N_5454,N_1985,N_3955);
or U5455 (N_5455,N_2688,N_179);
or U5456 (N_5456,N_2167,N_2603);
nor U5457 (N_5457,N_849,N_3374);
nand U5458 (N_5458,N_1025,N_1213);
nor U5459 (N_5459,N_511,N_4319);
nor U5460 (N_5460,N_4579,N_1424);
or U5461 (N_5461,N_3087,N_4037);
nor U5462 (N_5462,N_1808,N_2447);
nor U5463 (N_5463,N_3264,N_3202);
nand U5464 (N_5464,N_451,N_1731);
nand U5465 (N_5465,N_1140,N_4724);
and U5466 (N_5466,N_4682,N_3505);
nor U5467 (N_5467,N_1065,N_3680);
and U5468 (N_5468,N_1260,N_144);
or U5469 (N_5469,N_782,N_637);
and U5470 (N_5470,N_4200,N_4591);
nor U5471 (N_5471,N_1717,N_4686);
nor U5472 (N_5472,N_4639,N_1317);
and U5473 (N_5473,N_3844,N_2555);
and U5474 (N_5474,N_4743,N_3724);
nor U5475 (N_5475,N_3698,N_735);
nor U5476 (N_5476,N_2181,N_4196);
and U5477 (N_5477,N_1401,N_904);
or U5478 (N_5478,N_2988,N_881);
nor U5479 (N_5479,N_4004,N_4740);
and U5480 (N_5480,N_22,N_1651);
nand U5481 (N_5481,N_944,N_2051);
nand U5482 (N_5482,N_2328,N_1055);
and U5483 (N_5483,N_850,N_3016);
nor U5484 (N_5484,N_2387,N_840);
nor U5485 (N_5485,N_2955,N_1434);
and U5486 (N_5486,N_2516,N_27);
nor U5487 (N_5487,N_1654,N_103);
or U5488 (N_5488,N_4824,N_4906);
nor U5489 (N_5489,N_3942,N_1710);
and U5490 (N_5490,N_1463,N_3295);
and U5491 (N_5491,N_1780,N_3235);
and U5492 (N_5492,N_532,N_933);
and U5493 (N_5493,N_683,N_2707);
and U5494 (N_5494,N_4338,N_1264);
nor U5495 (N_5495,N_4051,N_2952);
nor U5496 (N_5496,N_1038,N_3891);
or U5497 (N_5497,N_2693,N_3898);
nor U5498 (N_5498,N_4403,N_1840);
and U5499 (N_5499,N_3062,N_3722);
nand U5500 (N_5500,N_520,N_3277);
nand U5501 (N_5501,N_1445,N_1906);
and U5502 (N_5502,N_404,N_3225);
nand U5503 (N_5503,N_443,N_2344);
nand U5504 (N_5504,N_4438,N_4190);
nor U5505 (N_5505,N_995,N_2340);
or U5506 (N_5506,N_4504,N_3699);
and U5507 (N_5507,N_4185,N_731);
nor U5508 (N_5508,N_1262,N_4260);
and U5509 (N_5509,N_2380,N_2129);
or U5510 (N_5510,N_4401,N_4191);
nand U5511 (N_5511,N_1570,N_4532);
or U5512 (N_5512,N_2840,N_2985);
nand U5513 (N_5513,N_3445,N_3650);
and U5514 (N_5514,N_1975,N_615);
and U5515 (N_5515,N_4064,N_3814);
or U5516 (N_5516,N_1493,N_2285);
nand U5517 (N_5517,N_4828,N_4056);
nand U5518 (N_5518,N_3947,N_4290);
nand U5519 (N_5519,N_75,N_348);
nor U5520 (N_5520,N_1465,N_4895);
and U5521 (N_5521,N_639,N_3783);
nor U5522 (N_5522,N_4601,N_4626);
and U5523 (N_5523,N_4329,N_2053);
and U5524 (N_5524,N_192,N_4380);
or U5525 (N_5525,N_2014,N_1157);
nand U5526 (N_5526,N_3614,N_700);
nor U5527 (N_5527,N_2779,N_589);
nand U5528 (N_5528,N_161,N_321);
nor U5529 (N_5529,N_3806,N_3401);
and U5530 (N_5530,N_1054,N_4932);
or U5531 (N_5531,N_4705,N_3943);
and U5532 (N_5532,N_1226,N_92);
nor U5533 (N_5533,N_1239,N_4413);
nor U5534 (N_5534,N_1126,N_1824);
and U5535 (N_5535,N_2295,N_3486);
nand U5536 (N_5536,N_1863,N_1561);
and U5537 (N_5537,N_821,N_4347);
nand U5538 (N_5538,N_1645,N_1867);
nand U5539 (N_5539,N_3162,N_3372);
or U5540 (N_5540,N_4071,N_885);
or U5541 (N_5541,N_1237,N_3477);
and U5542 (N_5542,N_219,N_2611);
and U5543 (N_5543,N_555,N_4395);
nand U5544 (N_5544,N_4751,N_1160);
or U5545 (N_5545,N_822,N_333);
or U5546 (N_5546,N_4249,N_3153);
or U5547 (N_5547,N_1111,N_1411);
xor U5548 (N_5548,N_2891,N_914);
nor U5549 (N_5549,N_1796,N_1578);
nand U5550 (N_5550,N_3765,N_824);
nor U5551 (N_5551,N_4050,N_1266);
nand U5552 (N_5552,N_3557,N_2827);
nand U5553 (N_5553,N_2775,N_4034);
nand U5554 (N_5554,N_3171,N_2972);
and U5555 (N_5555,N_1598,N_4197);
and U5556 (N_5556,N_2319,N_1703);
nand U5557 (N_5557,N_1983,N_4393);
nor U5558 (N_5558,N_2940,N_4398);
nor U5559 (N_5559,N_3885,N_2530);
nor U5560 (N_5560,N_2433,N_3581);
nand U5561 (N_5561,N_4847,N_3865);
and U5562 (N_5562,N_4396,N_3652);
and U5563 (N_5563,N_1461,N_1193);
nand U5564 (N_5564,N_1474,N_3206);
nand U5565 (N_5565,N_3132,N_2676);
nand U5566 (N_5566,N_2596,N_666);
and U5567 (N_5567,N_290,N_3473);
nor U5568 (N_5568,N_4406,N_1128);
and U5569 (N_5569,N_3689,N_1398);
nand U5570 (N_5570,N_2788,N_754);
or U5571 (N_5571,N_2848,N_435);
nor U5572 (N_5572,N_841,N_4376);
or U5573 (N_5573,N_2746,N_1419);
and U5574 (N_5574,N_3310,N_4587);
xnor U5575 (N_5575,N_1560,N_2292);
or U5576 (N_5576,N_170,N_1958);
nand U5577 (N_5577,N_1344,N_420);
or U5578 (N_5578,N_1918,N_1601);
nor U5579 (N_5579,N_1604,N_2157);
or U5580 (N_5580,N_1650,N_2066);
or U5581 (N_5581,N_2576,N_897);
or U5582 (N_5582,N_2626,N_4510);
nor U5583 (N_5583,N_63,N_1522);
nand U5584 (N_5584,N_2532,N_1130);
or U5585 (N_5585,N_3798,N_2560);
nor U5586 (N_5586,N_424,N_4638);
or U5587 (N_5587,N_1279,N_163);
and U5588 (N_5588,N_2124,N_83);
nand U5589 (N_5589,N_2047,N_704);
nand U5590 (N_5590,N_4012,N_3168);
nor U5591 (N_5591,N_2038,N_1881);
nor U5592 (N_5592,N_4140,N_1534);
nand U5593 (N_5593,N_4728,N_2774);
nor U5594 (N_5594,N_2705,N_4032);
nor U5595 (N_5595,N_1793,N_4308);
nor U5596 (N_5596,N_3996,N_1523);
or U5597 (N_5597,N_785,N_4095);
and U5598 (N_5598,N_1469,N_2079);
nor U5599 (N_5599,N_798,N_246);
and U5600 (N_5600,N_4684,N_1050);
and U5601 (N_5601,N_3966,N_780);
and U5602 (N_5602,N_1823,N_73);
nand U5603 (N_5603,N_3068,N_3196);
or U5604 (N_5604,N_1467,N_2413);
and U5605 (N_5605,N_3370,N_2162);
or U5606 (N_5606,N_2133,N_4901);
nor U5607 (N_5607,N_4859,N_3998);
nor U5608 (N_5608,N_127,N_3666);
or U5609 (N_5609,N_1195,N_1515);
nand U5610 (N_5610,N_1934,N_1433);
or U5611 (N_5611,N_3014,N_4537);
or U5612 (N_5612,N_3463,N_542);
nor U5613 (N_5613,N_1783,N_1018);
or U5614 (N_5614,N_3642,N_1726);
xor U5615 (N_5615,N_1149,N_3388);
or U5616 (N_5616,N_11,N_2168);
or U5617 (N_5617,N_2730,N_4752);
nand U5618 (N_5618,N_2313,N_4411);
nor U5619 (N_5619,N_2967,N_1743);
and U5620 (N_5620,N_3332,N_184);
nor U5621 (N_5621,N_2761,N_4716);
or U5622 (N_5622,N_3855,N_2620);
and U5623 (N_5623,N_302,N_1535);
nor U5624 (N_5624,N_1153,N_2563);
nor U5625 (N_5625,N_3619,N_3550);
or U5626 (N_5626,N_793,N_2149);
or U5627 (N_5627,N_3279,N_3907);
or U5628 (N_5628,N_1182,N_3103);
or U5629 (N_5629,N_1117,N_1301);
and U5630 (N_5630,N_4006,N_19);
nand U5631 (N_5631,N_1955,N_1756);
nor U5632 (N_5632,N_255,N_1909);
and U5633 (N_5633,N_4644,N_2724);
nand U5634 (N_5634,N_1084,N_3757);
nor U5635 (N_5635,N_3802,N_250);
nor U5636 (N_5636,N_2612,N_123);
nand U5637 (N_5637,N_167,N_2252);
or U5638 (N_5638,N_1919,N_659);
nand U5639 (N_5639,N_2834,N_3416);
or U5640 (N_5640,N_1049,N_870);
nand U5641 (N_5641,N_55,N_1145);
and U5642 (N_5642,N_536,N_6);
nand U5643 (N_5643,N_3015,N_1910);
nor U5644 (N_5644,N_4452,N_2844);
nand U5645 (N_5645,N_4909,N_3831);
nor U5646 (N_5646,N_912,N_4549);
or U5647 (N_5647,N_2577,N_2166);
nand U5648 (N_5648,N_295,N_1676);
and U5649 (N_5649,N_330,N_1035);
nor U5650 (N_5650,N_4464,N_4637);
nor U5651 (N_5651,N_1458,N_4782);
xor U5652 (N_5652,N_2115,N_1937);
nor U5653 (N_5653,N_2211,N_4013);
nand U5654 (N_5654,N_3583,N_4668);
nor U5655 (N_5655,N_327,N_4487);
or U5656 (N_5656,N_113,N_4592);
nand U5657 (N_5657,N_3561,N_3975);
and U5658 (N_5658,N_537,N_2913);
and U5659 (N_5659,N_2640,N_4606);
nand U5660 (N_5660,N_2743,N_3980);
nor U5661 (N_5661,N_2559,N_4218);
nand U5662 (N_5662,N_2148,N_3954);
nor U5663 (N_5663,N_2932,N_3469);
and U5664 (N_5664,N_1372,N_1646);
nand U5665 (N_5665,N_1475,N_276);
nand U5666 (N_5666,N_1093,N_1092);
or U5667 (N_5667,N_486,N_4755);
nor U5668 (N_5668,N_466,N_4489);
nor U5669 (N_5669,N_1158,N_476);
nand U5670 (N_5670,N_3730,N_3069);
nand U5671 (N_5671,N_1293,N_4672);
nor U5672 (N_5672,N_4561,N_1928);
or U5673 (N_5673,N_4954,N_3997);
nor U5674 (N_5674,N_1261,N_753);
or U5675 (N_5675,N_132,N_2241);
or U5676 (N_5676,N_4720,N_2505);
and U5677 (N_5677,N_2150,N_242);
or U5678 (N_5678,N_676,N_3133);
and U5679 (N_5679,N_2842,N_4664);
and U5680 (N_5680,N_3608,N_1688);
and U5681 (N_5681,N_3424,N_1815);
nor U5682 (N_5682,N_3740,N_3771);
or U5683 (N_5683,N_166,N_3227);
and U5684 (N_5684,N_3983,N_1884);
nor U5685 (N_5685,N_2508,N_4066);
nand U5686 (N_5686,N_4091,N_3759);
nand U5687 (N_5687,N_1053,N_1905);
or U5688 (N_5688,N_1685,N_3457);
nor U5689 (N_5689,N_1956,N_550);
or U5690 (N_5690,N_4941,N_1402);
or U5691 (N_5691,N_3061,N_913);
or U5692 (N_5692,N_2542,N_4408);
nand U5693 (N_5693,N_2531,N_4085);
or U5694 (N_5694,N_4739,N_4477);
nand U5695 (N_5695,N_3742,N_1697);
nor U5696 (N_5696,N_3169,N_1043);
or U5697 (N_5697,N_3109,N_4880);
nor U5698 (N_5698,N_147,N_2474);
nor U5699 (N_5699,N_4912,N_102);
nand U5700 (N_5700,N_3620,N_3154);
and U5701 (N_5701,N_4330,N_4846);
nand U5702 (N_5702,N_852,N_4345);
nor U5703 (N_5703,N_4516,N_1029);
nand U5704 (N_5704,N_1555,N_2442);
nand U5705 (N_5705,N_1008,N_4840);
nor U5706 (N_5706,N_3250,N_2482);
nand U5707 (N_5707,N_2742,N_2533);
and U5708 (N_5708,N_1315,N_4934);
or U5709 (N_5709,N_903,N_847);
nand U5710 (N_5710,N_3952,N_1666);
nor U5711 (N_5711,N_4488,N_3049);
or U5712 (N_5712,N_3950,N_1171);
or U5713 (N_5713,N_1761,N_1077);
or U5714 (N_5714,N_1818,N_1);
or U5715 (N_5715,N_2758,N_2628);
nor U5716 (N_5716,N_4097,N_2864);
and U5717 (N_5717,N_3847,N_4542);
nor U5718 (N_5718,N_3637,N_4086);
nand U5719 (N_5719,N_1963,N_3899);
or U5720 (N_5720,N_282,N_4131);
nor U5721 (N_5721,N_251,N_809);
or U5722 (N_5722,N_164,N_483);
and U5723 (N_5723,N_2350,N_4204);
and U5724 (N_5724,N_3528,N_472);
and U5725 (N_5725,N_1596,N_1527);
and U5726 (N_5726,N_3462,N_1874);
nand U5727 (N_5727,N_3282,N_2125);
nand U5728 (N_5728,N_1957,N_1118);
or U5729 (N_5729,N_2507,N_3003);
or U5730 (N_5730,N_2304,N_3418);
and U5731 (N_5731,N_4972,N_663);
or U5732 (N_5732,N_2037,N_1862);
or U5733 (N_5733,N_4640,N_1207);
nor U5734 (N_5734,N_1791,N_1786);
and U5735 (N_5735,N_3799,N_4693);
nor U5736 (N_5736,N_407,N_602);
nand U5737 (N_5737,N_2391,N_2498);
nor U5738 (N_5738,N_4707,N_3843);
or U5739 (N_5739,N_3568,N_3686);
or U5740 (N_5740,N_2183,N_3634);
or U5741 (N_5741,N_2246,N_4381);
nor U5742 (N_5742,N_1584,N_1627);
nand U5743 (N_5743,N_4798,N_4077);
nor U5744 (N_5744,N_3034,N_1016);
nor U5745 (N_5745,N_3811,N_1628);
and U5746 (N_5746,N_2916,N_1886);
nor U5747 (N_5747,N_1059,N_4897);
and U5748 (N_5748,N_2421,N_1618);
and U5749 (N_5749,N_1339,N_241);
nand U5750 (N_5750,N_1409,N_3000);
and U5751 (N_5751,N_2894,N_4611);
nand U5752 (N_5752,N_898,N_3272);
or U5753 (N_5753,N_2710,N_4916);
and U5754 (N_5754,N_3813,N_2132);
nand U5755 (N_5755,N_2887,N_3352);
nand U5756 (N_5756,N_2469,N_1668);
or U5757 (N_5757,N_2480,N_1211);
and U5758 (N_5758,N_2959,N_1377);
and U5759 (N_5759,N_2093,N_2029);
or U5760 (N_5760,N_3908,N_1294);
nand U5761 (N_5761,N_233,N_1190);
nor U5762 (N_5762,N_3860,N_2147);
nand U5763 (N_5763,N_1450,N_1449);
and U5764 (N_5764,N_1966,N_2239);
nor U5765 (N_5765,N_2193,N_959);
or U5766 (N_5766,N_2386,N_986);
and U5767 (N_5767,N_4292,N_1682);
nor U5768 (N_5768,N_1359,N_1416);
and U5769 (N_5769,N_4754,N_200);
nor U5770 (N_5770,N_1131,N_3963);
nor U5771 (N_5771,N_2722,N_3921);
nand U5772 (N_5772,N_240,N_2598);
nor U5773 (N_5773,N_1484,N_1167);
and U5774 (N_5774,N_3536,N_4307);
and U5775 (N_5775,N_3229,N_108);
nand U5776 (N_5776,N_1383,N_4557);
or U5777 (N_5777,N_4243,N_3455);
or U5778 (N_5778,N_2906,N_1748);
or U5779 (N_5779,N_3252,N_4882);
or U5780 (N_5780,N_1040,N_3714);
nor U5781 (N_5781,N_3364,N_1787);
nand U5782 (N_5782,N_1917,N_4825);
nor U5783 (N_5783,N_171,N_186);
nor U5784 (N_5784,N_3599,N_1308);
and U5785 (N_5785,N_291,N_4991);
nor U5786 (N_5786,N_3335,N_1997);
and U5787 (N_5787,N_4221,N_205);
and U5788 (N_5788,N_2341,N_1892);
nand U5789 (N_5789,N_3351,N_742);
nand U5790 (N_5790,N_2568,N_4563);
and U5791 (N_5791,N_1642,N_2455);
or U5792 (N_5792,N_4826,N_678);
or U5793 (N_5793,N_3091,N_584);
or U5794 (N_5794,N_4216,N_2099);
nand U5795 (N_5795,N_3769,N_632);
nand U5796 (N_5796,N_2958,N_4848);
or U5797 (N_5797,N_1730,N_921);
nand U5798 (N_5798,N_2041,N_2833);
nor U5799 (N_5799,N_1246,N_3190);
nand U5800 (N_5800,N_288,N_4585);
nand U5801 (N_5801,N_2968,N_3621);
nand U5802 (N_5802,N_376,N_835);
nor U5803 (N_5803,N_3434,N_3797);
or U5804 (N_5804,N_971,N_3367);
or U5805 (N_5805,N_1999,N_4980);
and U5806 (N_5806,N_4429,N_559);
nand U5807 (N_5807,N_862,N_436);
nand U5808 (N_5808,N_1877,N_1629);
nand U5809 (N_5809,N_1127,N_340);
nor U5810 (N_5810,N_1851,N_4156);
nand U5811 (N_5811,N_1891,N_3981);
and U5812 (N_5812,N_3866,N_4110);
or U5813 (N_5813,N_3600,N_2813);
or U5814 (N_5814,N_378,N_4046);
and U5815 (N_5815,N_3906,N_4316);
nand U5816 (N_5816,N_4683,N_3638);
nand U5817 (N_5817,N_1898,N_1511);
nor U5818 (N_5818,N_2564,N_1593);
and U5819 (N_5819,N_4366,N_3558);
nand U5820 (N_5820,N_558,N_2347);
nand U5821 (N_5821,N_3738,N_1252);
nand U5822 (N_5822,N_4475,N_4662);
or U5823 (N_5823,N_254,N_1318);
nand U5824 (N_5824,N_4472,N_2030);
or U5825 (N_5825,N_918,N_1350);
xnor U5826 (N_5826,N_3460,N_474);
and U5827 (N_5827,N_2363,N_3029);
nand U5828 (N_5828,N_2116,N_4384);
nand U5829 (N_5829,N_3663,N_2189);
nand U5830 (N_5830,N_1284,N_2440);
or U5831 (N_5831,N_3958,N_4908);
and U5832 (N_5832,N_3005,N_823);
nand U5833 (N_5833,N_3048,N_716);
and U5834 (N_5834,N_447,N_505);
or U5835 (N_5835,N_2656,N_814);
or U5836 (N_5836,N_763,N_2431);
or U5837 (N_5837,N_1299,N_3412);
or U5838 (N_5838,N_2458,N_116);
nand U5839 (N_5839,N_3971,N_3526);
nor U5840 (N_5840,N_2896,N_1700);
nand U5841 (N_5841,N_3131,N_2825);
or U5842 (N_5842,N_2026,N_2580);
nor U5843 (N_5843,N_4154,N_1075);
or U5844 (N_5844,N_4513,N_2760);
nand U5845 (N_5845,N_4247,N_3692);
and U5846 (N_5846,N_679,N_3451);
and U5847 (N_5847,N_1855,N_2202);
and U5848 (N_5848,N_362,N_522);
nand U5849 (N_5849,N_322,N_292);
or U5850 (N_5850,N_1229,N_1313);
or U5851 (N_5851,N_79,N_1543);
nand U5852 (N_5852,N_3415,N_2659);
nor U5853 (N_5853,N_60,N_37);
and U5854 (N_5854,N_4645,N_1352);
and U5855 (N_5855,N_3672,N_4193);
and U5856 (N_5856,N_126,N_2870);
nand U5857 (N_5857,N_3823,N_2260);
and U5858 (N_5858,N_4850,N_2098);
and U5859 (N_5859,N_65,N_614);
or U5860 (N_5860,N_383,N_2273);
nor U5861 (N_5861,N_4142,N_854);
nor U5862 (N_5862,N_216,N_880);
or U5863 (N_5863,N_3602,N_3579);
nor U5864 (N_5864,N_794,N_206);
nor U5865 (N_5865,N_3554,N_1286);
nand U5866 (N_5866,N_2302,N_2645);
nand U5867 (N_5867,N_1765,N_4514);
or U5868 (N_5868,N_723,N_417);
nor U5869 (N_5869,N_3319,N_2725);
nor U5870 (N_5870,N_1204,N_645);
nor U5871 (N_5871,N_1788,N_3886);
nor U5872 (N_5872,N_4813,N_3931);
nor U5873 (N_5873,N_458,N_4295);
and U5874 (N_5874,N_3487,N_4177);
and U5875 (N_5875,N_1015,N_461);
and U5876 (N_5876,N_3882,N_3039);
nand U5877 (N_5877,N_2991,N_3318);
and U5878 (N_5878,N_1396,N_1856);
nand U5879 (N_5879,N_2072,N_3857);
or U5880 (N_5880,N_4081,N_4531);
and U5881 (N_5881,N_877,N_1276);
and U5882 (N_5882,N_42,N_1457);
nand U5883 (N_5883,N_3357,N_4533);
or U5884 (N_5884,N_4750,N_2366);
and U5885 (N_5885,N_4873,N_4630);
nor U5886 (N_5886,N_1695,N_3859);
nor U5887 (N_5887,N_3881,N_4449);
nor U5888 (N_5888,N_4283,N_953);
nand U5889 (N_5889,N_218,N_1524);
xnor U5890 (N_5890,N_3564,N_2618);
and U5891 (N_5891,N_3576,N_2266);
nand U5892 (N_5892,N_274,N_2112);
nand U5893 (N_5893,N_4443,N_1326);
nand U5894 (N_5894,N_3280,N_1394);
or U5895 (N_5895,N_1495,N_3114);
nor U5896 (N_5896,N_1828,N_2690);
and U5897 (N_5897,N_2339,N_2420);
nor U5898 (N_5898,N_148,N_3084);
or U5899 (N_5899,N_2159,N_4761);
nor U5900 (N_5900,N_761,N_4327);
and U5901 (N_5901,N_4610,N_681);
or U5902 (N_5902,N_2106,N_698);
nand U5903 (N_5903,N_3640,N_817);
nor U5904 (N_5904,N_4212,N_3080);
or U5905 (N_5905,N_2931,N_374);
nand U5906 (N_5906,N_915,N_2820);
or U5907 (N_5907,N_1658,N_1968);
and U5908 (N_5908,N_1712,N_1929);
nor U5909 (N_5909,N_2639,N_1973);
nand U5910 (N_5910,N_1592,N_2644);
and U5911 (N_5911,N_1722,N_4405);
nor U5912 (N_5912,N_776,N_2223);
and U5913 (N_5913,N_4827,N_1683);
or U5914 (N_5914,N_2717,N_1309);
nand U5915 (N_5915,N_608,N_1231);
nand U5916 (N_5916,N_2616,N_1845);
nor U5917 (N_5917,N_4698,N_3719);
or U5918 (N_5918,N_4987,N_160);
or U5919 (N_5919,N_1270,N_2462);
and U5920 (N_5920,N_4009,N_1547);
nor U5921 (N_5921,N_2583,N_1376);
nor U5922 (N_5922,N_2080,N_4721);
nor U5923 (N_5923,N_2536,N_4058);
nand U5924 (N_5924,N_2332,N_4049);
or U5925 (N_5925,N_195,N_1655);
xor U5926 (N_5926,N_2630,N_606);
or U5927 (N_5927,N_4809,N_2964);
and U5928 (N_5928,N_4299,N_3760);
nand U5929 (N_5929,N_1133,N_2356);
nand U5930 (N_5930,N_3549,N_2235);
nand U5931 (N_5931,N_1804,N_4174);
nor U5932 (N_5932,N_2070,N_1915);
or U5933 (N_5933,N_4926,N_3927);
nor U5934 (N_5934,N_2497,N_4952);
nor U5935 (N_5935,N_1776,N_3965);
or U5936 (N_5936,N_3488,N_992);
or U5937 (N_5937,N_4663,N_3697);
and U5938 (N_5938,N_4346,N_919);
nor U5939 (N_5939,N_1163,N_591);
and U5940 (N_5940,N_1621,N_2308);
and U5941 (N_5941,N_4144,N_3098);
nor U5942 (N_5942,N_1106,N_2471);
and U5943 (N_5943,N_4492,N_3509);
or U5944 (N_5944,N_2773,N_4985);
and U5945 (N_5945,N_604,N_2914);
nand U5946 (N_5946,N_999,N_4239);
nand U5947 (N_5947,N_3165,N_2105);
nor U5948 (N_5948,N_2370,N_3126);
nor U5949 (N_5949,N_2258,N_3234);
or U5950 (N_5950,N_2624,N_3135);
and U5951 (N_5951,N_4890,N_3934);
and U5952 (N_5952,N_2990,N_622);
and U5953 (N_5953,N_1174,N_4902);
nor U5954 (N_5954,N_4956,N_1122);
and U5955 (N_5955,N_3693,N_1071);
nor U5956 (N_5956,N_3969,N_1414);
or U5957 (N_5957,N_4819,N_2137);
and U5958 (N_5958,N_1762,N_35);
or U5959 (N_5959,N_412,N_3873);
or U5960 (N_5960,N_3880,N_4390);
nor U5961 (N_5961,N_573,N_744);
and U5962 (N_5962,N_3490,N_1179);
or U5963 (N_5963,N_3336,N_3492);
or U5964 (N_5964,N_3186,N_3829);
nand U5965 (N_5965,N_3681,N_4757);
and U5966 (N_5966,N_2892,N_4378);
xor U5967 (N_5967,N_4018,N_3779);
and U5968 (N_5968,N_2086,N_189);
or U5969 (N_5969,N_3938,N_4869);
nand U5970 (N_5970,N_2238,N_2262);
nor U5971 (N_5971,N_2407,N_2418);
and U5972 (N_5972,N_2100,N_3586);
or U5973 (N_5973,N_51,N_1283);
nor U5974 (N_5974,N_4192,N_1141);
nand U5975 (N_5975,N_1391,N_1771);
and U5976 (N_5976,N_1321,N_1519);
or U5977 (N_5977,N_908,N_993);
nand U5978 (N_5978,N_4432,N_1623);
nor U5979 (N_5979,N_3763,N_395);
or U5980 (N_5980,N_1557,N_3531);
nand U5981 (N_5981,N_657,N_4028);
nor U5982 (N_5982,N_2936,N_3658);
nor U5983 (N_5983,N_449,N_543);
nor U5984 (N_5984,N_2648,N_1342);
nor U5985 (N_5985,N_969,N_1811);
or U5986 (N_5986,N_4208,N_1573);
or U5987 (N_5987,N_3497,N_415);
or U5988 (N_5988,N_2835,N_649);
or U5989 (N_5989,N_3350,N_2770);
nand U5990 (N_5990,N_1421,N_3530);
nor U5991 (N_5991,N_2585,N_4270);
nor U5992 (N_5992,N_426,N_4804);
or U5993 (N_5993,N_1843,N_2058);
nor U5994 (N_5994,N_3140,N_1872);
nor U5995 (N_5995,N_4486,N_3708);
and U5996 (N_5996,N_1490,N_2650);
or U5997 (N_5997,N_4007,N_2068);
nand U5998 (N_5998,N_4622,N_338);
and U5999 (N_5999,N_2741,N_1225);
nand U6000 (N_6000,N_4124,N_2994);
or U6001 (N_6001,N_4666,N_351);
nor U6002 (N_6002,N_4165,N_3524);
nor U6003 (N_6003,N_1982,N_3715);
or U6004 (N_6004,N_3594,N_3354);
and U6005 (N_6005,N_4805,N_2769);
nand U6006 (N_6006,N_4960,N_4296);
nor U6007 (N_6007,N_3690,N_119);
nor U6008 (N_6008,N_2244,N_778);
or U6009 (N_6009,N_4706,N_4278);
and U6010 (N_6010,N_3239,N_4789);
or U6011 (N_6011,N_4690,N_319);
xnor U6012 (N_6012,N_653,N_4581);
nor U6013 (N_6013,N_513,N_2282);
nand U6014 (N_6014,N_1571,N_2123);
and U6015 (N_6015,N_4677,N_1660);
nand U6016 (N_6016,N_2675,N_2795);
nor U6017 (N_6017,N_2855,N_2216);
or U6018 (N_6018,N_2589,N_3064);
nand U6019 (N_6019,N_2393,N_1630);
or U6020 (N_6020,N_1837,N_4354);
and U6021 (N_6021,N_3778,N_4083);
and U6022 (N_6022,N_3826,N_4246);
nand U6023 (N_6023,N_4114,N_243);
and U6024 (N_6024,N_457,N_4511);
nor U6025 (N_6025,N_4763,N_3498);
nand U6026 (N_6026,N_4469,N_4852);
nor U6027 (N_6027,N_2846,N_1340);
nor U6028 (N_6028,N_1789,N_4369);
and U6029 (N_6029,N_1155,N_3344);
nor U6030 (N_6030,N_932,N_188);
or U6031 (N_6031,N_4631,N_4236);
and U6032 (N_6032,N_2002,N_1329);
nor U6033 (N_6033,N_1572,N_3298);
nand U6034 (N_6034,N_3575,N_2473);
nand U6035 (N_6035,N_3317,N_1489);
and U6036 (N_6036,N_962,N_484);
or U6037 (N_6037,N_1941,N_4115);
nor U6038 (N_6038,N_633,N_3935);
nand U6039 (N_6039,N_128,N_3501);
or U6040 (N_6040,N_2361,N_1347);
nand U6041 (N_6041,N_498,N_2721);
or U6042 (N_6042,N_1289,N_3618);
or U6043 (N_6043,N_1699,N_3894);
nor U6044 (N_6044,N_3376,N_2454);
or U6045 (N_6045,N_4726,N_1900);
or U6046 (N_6046,N_3591,N_4448);
and U6047 (N_6047,N_4412,N_4776);
and U6048 (N_6048,N_4795,N_563);
nor U6049 (N_6049,N_2557,N_4874);
nand U6050 (N_6050,N_3291,N_4523);
nand U6051 (N_6051,N_4893,N_829);
and U6052 (N_6052,N_2288,N_970);
or U6053 (N_6053,N_1510,N_869);
or U6054 (N_6054,N_2706,N_807);
nand U6055 (N_6055,N_2709,N_3377);
or U6056 (N_6056,N_1649,N_442);
nor U6057 (N_6057,N_3585,N_2392);
and U6058 (N_6058,N_507,N_3436);
nor U6059 (N_6059,N_271,N_3099);
or U6060 (N_6060,N_3134,N_2311);
nor U6061 (N_6061,N_4431,N_4397);
or U6062 (N_6062,N_4430,N_777);
nor U6063 (N_6063,N_3781,N_3041);
or U6064 (N_6064,N_3300,N_3817);
and U6065 (N_6065,N_1257,N_4831);
nand U6066 (N_6066,N_3493,N_3822);
or U6067 (N_6067,N_4482,N_4509);
or U6068 (N_6068,N_819,N_2643);
or U6069 (N_6069,N_3517,N_4747);
nand U6070 (N_6070,N_2969,N_2372);
and U6071 (N_6071,N_4202,N_2547);
nand U6072 (N_6072,N_786,N_2364);
nand U6073 (N_6073,N_1273,N_4992);
nor U6074 (N_6074,N_1019,N_3258);
and U6075 (N_6075,N_799,N_3195);
or U6076 (N_6076,N_3065,N_2698);
nor U6077 (N_6077,N_4568,N_2275);
nand U6078 (N_6078,N_3271,N_2763);
nor U6079 (N_6079,N_3653,N_3247);
and U6080 (N_6080,N_44,N_2912);
or U6081 (N_6081,N_4844,N_1088);
nand U6082 (N_6082,N_623,N_3949);
nor U6083 (N_6083,N_699,N_373);
nand U6084 (N_6084,N_4894,N_7);
nor U6085 (N_6085,N_259,N_1720);
and U6086 (N_6086,N_3974,N_1508);
nor U6087 (N_6087,N_2966,N_4341);
nand U6088 (N_6088,N_4787,N_1191);
nand U6089 (N_6089,N_1045,N_111);
or U6090 (N_6090,N_3461,N_4418);
and U6091 (N_6091,N_1635,N_2224);
nor U6092 (N_6092,N_748,N_2427);
and U6093 (N_6093,N_4422,N_2578);
and U6094 (N_6094,N_2600,N_3273);
xor U6095 (N_6095,N_1098,N_1608);
or U6096 (N_6096,N_4989,N_4543);
nand U6097 (N_6097,N_2472,N_3117);
or U6098 (N_6098,N_428,N_4104);
and U6099 (N_6099,N_1687,N_4702);
or U6100 (N_6100,N_4995,N_1768);
nand U6101 (N_6101,N_2065,N_1202);
or U6102 (N_6102,N_876,N_2139);
nor U6103 (N_6103,N_4615,N_2324);
and U6104 (N_6104,N_682,N_779);
xor U6105 (N_6105,N_3100,N_1991);
and U6106 (N_6106,N_1081,N_4554);
or U6107 (N_6107,N_961,N_4586);
nand U6108 (N_6108,N_309,N_570);
or U6109 (N_6109,N_4661,N_1671);
or U6110 (N_6110,N_32,N_3662);
nand U6111 (N_6111,N_524,N_1104);
or U6112 (N_6112,N_783,N_3869);
nor U6113 (N_6113,N_3129,N_5);
nor U6114 (N_6114,N_4569,N_1691);
nand U6115 (N_6115,N_3535,N_526);
nor U6116 (N_6116,N_2778,N_749);
or U6117 (N_6117,N_2409,N_3381);
and U6118 (N_6118,N_3155,N_90);
and U6119 (N_6119,N_769,N_1498);
and U6120 (N_6120,N_4442,N_2334);
and U6121 (N_6121,N_2681,N_1894);
nor U6122 (N_6122,N_1740,N_1139);
and U6123 (N_6123,N_1258,N_239);
and U6124 (N_6124,N_1491,N_3074);
and U6125 (N_6125,N_4262,N_4062);
or U6126 (N_6126,N_816,N_1904);
or U6127 (N_6127,N_3122,N_2869);
and U6128 (N_6128,N_2799,N_2946);
or U6129 (N_6129,N_2939,N_2475);
or U6130 (N_6130,N_3888,N_4370);
and U6131 (N_6131,N_1809,N_2712);
nor U6132 (N_6132,N_1123,N_377);
and U6133 (N_6133,N_190,N_225);
and U6134 (N_6134,N_1954,N_1451);
nand U6135 (N_6135,N_729,N_705);
nand U6136 (N_6136,N_101,N_3567);
and U6137 (N_6137,N_2494,N_3825);
and U6138 (N_6138,N_4958,N_924);
nand U6139 (N_6139,N_1698,N_4090);
nor U6140 (N_6140,N_4905,N_1614);
nand U6141 (N_6141,N_4476,N_2231);
or U6142 (N_6142,N_2915,N_2694);
or U6143 (N_6143,N_384,N_1734);
nor U6144 (N_6144,N_3764,N_985);
nor U6145 (N_6145,N_4267,N_2691);
and U6146 (N_6146,N_3547,N_2071);
nor U6147 (N_6147,N_4371,N_124);
nor U6148 (N_6148,N_1278,N_3120);
and U6149 (N_6149,N_1162,N_4801);
and U6150 (N_6150,N_931,N_1086);
or U6151 (N_6151,N_3805,N_1310);
and U6152 (N_6152,N_4674,N_1014);
or U6153 (N_6153,N_2668,N_2581);
nor U6154 (N_6154,N_3223,N_4800);
or U6155 (N_6155,N_4915,N_3136);
nand U6156 (N_6156,N_354,N_575);
and U6157 (N_6157,N_1943,N_4551);
and U6158 (N_6158,N_4463,N_1374);
nand U6159 (N_6159,N_427,N_150);
and U6160 (N_6160,N_2938,N_1438);
and U6161 (N_6161,N_1582,N_1589);
nor U6162 (N_6162,N_2832,N_4541);
nor U6163 (N_6163,N_1694,N_1675);
or U6164 (N_6164,N_4119,N_2219);
or U6165 (N_6165,N_528,N_2860);
or U6166 (N_6166,N_4923,N_198);
or U6167 (N_6167,N_401,N_2259);
and U6168 (N_6168,N_3733,N_2028);
nand U6169 (N_6169,N_3808,N_140);
nor U6170 (N_6170,N_257,N_4965);
nor U6171 (N_6171,N_1206,N_318);
and U6172 (N_6172,N_1914,N_2317);
nor U6173 (N_6173,N_3948,N_4990);
nor U6174 (N_6174,N_2336,N_392);
or U6175 (N_6175,N_2594,N_651);
or U6176 (N_6176,N_2200,N_1782);
nor U6177 (N_6177,N_2552,N_1550);
nand U6178 (N_6178,N_2173,N_52);
or U6179 (N_6179,N_3870,N_3410);
and U6180 (N_6180,N_2283,N_2622);
nor U6181 (N_6181,N_2297,N_3260);
or U6182 (N_6182,N_1879,N_804);
nand U6183 (N_6183,N_118,N_1102);
and U6184 (N_6184,N_4748,N_1802);
or U6185 (N_6185,N_4450,N_3774);
and U6186 (N_6186,N_2128,N_4163);
or U6187 (N_6187,N_701,N_3511);
nor U6188 (N_6188,N_2858,N_4019);
and U6189 (N_6189,N_2853,N_1505);
nand U6190 (N_6190,N_2984,N_388);
and U6191 (N_6191,N_1338,N_2367);
or U6192 (N_6192,N_4709,N_1821);
nor U6193 (N_6193,N_3542,N_266);
or U6194 (N_6194,N_3696,N_773);
nor U6195 (N_6195,N_3701,N_968);
or U6196 (N_6196,N_2646,N_2151);
and U6197 (N_6197,N_3276,N_3872);
nor U6198 (N_6198,N_3683,N_4271);
nand U6199 (N_6199,N_1970,N_4222);
or U6200 (N_6200,N_4802,N_1750);
nand U6201 (N_6201,N_864,N_347);
nor U6202 (N_6202,N_3716,N_4527);
and U6203 (N_6203,N_2764,N_54);
or U6204 (N_6204,N_4454,N_1442);
nor U6205 (N_6205,N_4079,N_185);
and U6206 (N_6206,N_45,N_1412);
nor U6207 (N_6207,N_2130,N_737);
nand U6208 (N_6208,N_394,N_3379);
nor U6209 (N_6209,N_4774,N_2948);
and U6210 (N_6210,N_4957,N_1357);
or U6211 (N_6211,N_556,N_1706);
or U6212 (N_6212,N_1046,N_4646);
and U6213 (N_6213,N_4913,N_316);
or U6214 (N_6214,N_4220,N_4620);
and U6215 (N_6215,N_2545,N_2020);
nor U6216 (N_6216,N_4671,N_3819);
and U6217 (N_6217,N_393,N_3674);
or U6218 (N_6218,N_3447,N_4072);
nand U6219 (N_6219,N_3198,N_983);
and U6220 (N_6220,N_2045,N_21);
nor U6221 (N_6221,N_3281,N_846);
or U6222 (N_6222,N_3837,N_1744);
and U6223 (N_6223,N_387,N_1428);
or U6224 (N_6224,N_703,N_3387);
nand U6225 (N_6225,N_1549,N_781);
and U6226 (N_6226,N_2785,N_1678);
and U6227 (N_6227,N_2230,N_2011);
nand U6228 (N_6228,N_3789,N_1068);
nor U6229 (N_6229,N_3951,N_4263);
and U6230 (N_6230,N_1962,N_713);
nor U6231 (N_6231,N_413,N_1070);
and U6232 (N_6232,N_770,N_423);
nand U6233 (N_6233,N_1633,N_2570);
nor U6234 (N_6234,N_494,N_4067);
nor U6235 (N_6235,N_1826,N_2551);
and U6236 (N_6236,N_3884,N_1271);
nand U6237 (N_6237,N_3970,N_650);
and U6238 (N_6238,N_265,N_4678);
nand U6239 (N_6239,N_202,N_3660);
or U6240 (N_6240,N_1142,N_2204);
nor U6241 (N_6241,N_3776,N_4016);
and U6242 (N_6242,N_2439,N_2765);
or U6243 (N_6243,N_4911,N_2279);
nor U6244 (N_6244,N_3745,N_2422);
nor U6245 (N_6245,N_893,N_2465);
or U6246 (N_6246,N_1063,N_2642);
nor U6247 (N_6247,N_213,N_4473);
or U6248 (N_6248,N_788,N_300);
and U6249 (N_6249,N_4529,N_1974);
and U6250 (N_6250,N_569,N_861);
or U6251 (N_6251,N_2541,N_882);
nor U6252 (N_6252,N_1388,N_4922);
nand U6253 (N_6253,N_4470,N_448);
nor U6254 (N_6254,N_475,N_1488);
nor U6255 (N_6255,N_1188,N_1288);
nor U6256 (N_6256,N_1597,N_3661);
or U6257 (N_6257,N_1912,N_2198);
or U6258 (N_6258,N_2562,N_4944);
and U6259 (N_6259,N_2063,N_750);
or U6260 (N_6260,N_966,N_88);
nand U6261 (N_6261,N_1702,N_790);
or U6262 (N_6262,N_994,N_2883);
or U6263 (N_6263,N_3398,N_183);
or U6264 (N_6264,N_736,N_4003);
nor U6265 (N_6265,N_874,N_3792);
nor U6266 (N_6266,N_2539,N_3072);
nor U6267 (N_6267,N_4888,N_3390);
or U6268 (N_6268,N_527,N_1830);
nand U6269 (N_6269,N_129,N_1960);
nand U6270 (N_6270,N_796,N_3278);
or U6271 (N_6271,N_1735,N_3941);
nand U6272 (N_6272,N_1420,N_2965);
nor U6273 (N_6273,N_1090,N_2172);
nand U6274 (N_6274,N_2739,N_1545);
and U6275 (N_6275,N_2662,N_1138);
nand U6276 (N_6276,N_2477,N_2092);
and U6277 (N_6277,N_1233,N_372);
nor U6278 (N_6278,N_4577,N_2107);
nand U6279 (N_6279,N_677,N_739);
nand U6280 (N_6280,N_3812,N_2504);
or U6281 (N_6281,N_3184,N_4946);
nand U6282 (N_6282,N_4878,N_2905);
and U6283 (N_6283,N_4017,N_310);
and U6284 (N_6284,N_485,N_1337);
nand U6285 (N_6285,N_3553,N_1052);
nor U6286 (N_6286,N_4602,N_910);
nand U6287 (N_6287,N_3912,N_1353);
nand U6288 (N_6288,N_2631,N_3177);
nor U6289 (N_6289,N_3968,N_12);
nand U6290 (N_6290,N_516,N_3962);
and U6291 (N_6291,N_1644,N_1965);
or U6292 (N_6292,N_1033,N_339);
and U6293 (N_6293,N_4139,N_1314);
nand U6294 (N_6294,N_4143,N_2423);
nand U6295 (N_6295,N_2801,N_2343);
and U6296 (N_6296,N_3541,N_594);
and U6297 (N_6297,N_4770,N_539);
nor U6298 (N_6298,N_3375,N_106);
nor U6299 (N_6299,N_1478,N_3075);
or U6300 (N_6300,N_2412,N_4420);
nand U6301 (N_6301,N_396,N_4556);
and U6302 (N_6302,N_1320,N_298);
nand U6303 (N_6303,N_3213,N_1665);
nor U6304 (N_6304,N_4550,N_3197);
nor U6305 (N_6305,N_4986,N_3302);
nor U6306 (N_6306,N_529,N_93);
or U6307 (N_6307,N_2814,N_747);
and U6308 (N_6308,N_2750,N_845);
or U6309 (N_6309,N_3365,N_3371);
or U6310 (N_6310,N_2629,N_2453);
nor U6311 (N_6311,N_2389,N_4546);
and U6312 (N_6312,N_2004,N_2385);
and U6313 (N_6313,N_551,N_4435);
nand U6314 (N_6314,N_3900,N_1579);
nor U6315 (N_6315,N_4141,N_4351);
nand U6316 (N_6316,N_1101,N_4794);
and U6317 (N_6317,N_4596,N_579);
nor U6318 (N_6318,N_480,N_344);
nor U6319 (N_6319,N_2144,N_643);
nand U6320 (N_6320,N_571,N_3992);
and U6321 (N_6321,N_4628,N_2097);
nor U6322 (N_6322,N_2627,N_1328);
and U6323 (N_6323,N_2771,N_2345);
nor U6324 (N_6324,N_4609,N_989);
nand U6325 (N_6325,N_574,N_1085);
nor U6326 (N_6326,N_332,N_2291);
nor U6327 (N_6327,N_4447,N_3506);
nor U6328 (N_6328,N_4891,N_1165);
nor U6329 (N_6329,N_709,N_4242);
nor U6330 (N_6330,N_3625,N_4779);
or U6331 (N_6331,N_1216,N_1076);
nor U6332 (N_6332,N_181,N_4534);
and U6333 (N_6333,N_1986,N_4005);
nor U6334 (N_6334,N_3669,N_2961);
nor U6335 (N_6335,N_2067,N_3328);
nand U6336 (N_6336,N_1662,N_3977);
nand U6337 (N_6337,N_2256,N_2817);
or U6338 (N_6338,N_4942,N_4031);
nor U6339 (N_6339,N_2660,N_2687);
and U6340 (N_6340,N_3523,N_1810);
and U6341 (N_6341,N_4424,N_2674);
and U6342 (N_6342,N_857,N_977);
and U6343 (N_6343,N_3182,N_2191);
or U6344 (N_6344,N_687,N_4279);
or U6345 (N_6345,N_3656,N_314);
or U6346 (N_6346,N_3108,N_1590);
nand U6347 (N_6347,N_2619,N_3189);
or U6348 (N_6348,N_887,N_508);
or U6349 (N_6349,N_2636,N_3522);
nor U6350 (N_6350,N_2337,N_2873);
or U6351 (N_6351,N_3704,N_3124);
or U6352 (N_6352,N_936,N_1816);
or U6353 (N_6353,N_2975,N_1536);
and U6354 (N_6354,N_3097,N_2255);
or U6355 (N_6355,N_596,N_3373);
nand U6356 (N_6356,N_1846,N_467);
nor U6357 (N_6357,N_1479,N_1223);
or U6358 (N_6358,N_3755,N_3794);
and U6359 (N_6359,N_2064,N_973);
and U6360 (N_6360,N_1300,N_3472);
nor U6361 (N_6361,N_774,N_4654);
and U6362 (N_6362,N_3314,N_1241);
nor U6363 (N_6363,N_4866,N_293);
nor U6364 (N_6364,N_2610,N_3571);
nor U6365 (N_6365,N_4229,N_2806);
nand U6366 (N_6366,N_3500,N_1736);
and U6367 (N_6367,N_4277,N_3976);
nor U6368 (N_6368,N_1946,N_2759);
and U6369 (N_6369,N_2732,N_4535);
and U6370 (N_6370,N_2479,N_4318);
and U6371 (N_6371,N_3607,N_2333);
nand U6372 (N_6372,N_3721,N_1403);
nor U6373 (N_6373,N_16,N_3616);
nor U6374 (N_6374,N_1969,N_1994);
and U6375 (N_6375,N_2175,N_504);
and U6376 (N_6376,N_2006,N_1849);
nor U6377 (N_6377,N_2747,N_3226);
and U6378 (N_6378,N_335,N_3569);
and U6379 (N_6379,N_143,N_1992);
or U6380 (N_6380,N_3238,N_2298);
and U6381 (N_6381,N_3111,N_2448);
or U6382 (N_6382,N_605,N_3224);
or U6383 (N_6383,N_3933,N_1613);
nor U6384 (N_6384,N_3540,N_3876);
nor U6385 (N_6385,N_2951,N_2001);
or U6386 (N_6386,N_2182,N_3659);
or U6387 (N_6387,N_2425,N_1964);
nand U6388 (N_6388,N_1733,N_197);
nor U6389 (N_6389,N_3266,N_975);
nor U6390 (N_6390,N_722,N_1603);
or U6391 (N_6391,N_270,N_2859);
nor U6392 (N_6392,N_3160,N_210);
nand U6393 (N_6393,N_1679,N_3449);
or U6394 (N_6394,N_3901,N_675);
and U6395 (N_6395,N_2405,N_4758);
or U6396 (N_6396,N_4421,N_4955);
nand U6397 (N_6397,N_1006,N_3444);
or U6398 (N_6398,N_4659,N_2403);
or U6399 (N_6399,N_655,N_2658);
nand U6400 (N_6400,N_221,N_4930);
or U6401 (N_6401,N_2515,N_1143);
nand U6402 (N_6402,N_2022,N_833);
and U6403 (N_6403,N_4231,N_1607);
nor U6404 (N_6404,N_1173,N_2274);
and U6405 (N_6405,N_1865,N_3717);
or U6406 (N_6406,N_4305,N_3222);
or U6407 (N_6407,N_2476,N_2032);
or U6408 (N_6408,N_4904,N_1938);
or U6409 (N_6409,N_2754,N_2221);
nand U6410 (N_6410,N_2176,N_1468);
nand U6411 (N_6411,N_2415,N_2036);
nand U6412 (N_6412,N_142,N_3145);
or U6413 (N_6413,N_2342,N_828);
and U6414 (N_6414,N_1010,N_4011);
and U6415 (N_6415,N_115,N_3315);
and U6416 (N_6416,N_2977,N_630);
nor U6417 (N_6417,N_287,N_979);
or U6418 (N_6418,N_2496,N_2595);
nand U6419 (N_6419,N_802,N_3297);
and U6420 (N_6420,N_3673,N_419);
nand U6421 (N_6421,N_1274,N_3185);
or U6422 (N_6422,N_1980,N_1831);
and U6423 (N_6423,N_1741,N_4576);
or U6424 (N_6424,N_3342,N_3383);
nand U6425 (N_6425,N_3458,N_2731);
nand U6426 (N_6426,N_3465,N_4352);
nor U6427 (N_6427,N_3861,N_4181);
nand U6428 (N_6428,N_3752,N_2417);
nand U6429 (N_6429,N_3589,N_4109);
or U6430 (N_6430,N_837,N_182);
xnor U6431 (N_6431,N_2543,N_4984);
nor U6432 (N_6432,N_4695,N_4162);
nand U6433 (N_6433,N_3159,N_2845);
nor U6434 (N_6434,N_4993,N_2934);
nor U6435 (N_6435,N_1647,N_2040);
or U6436 (N_6436,N_3334,N_2850);
or U6437 (N_6437,N_4812,N_2861);
nand U6438 (N_6438,N_4073,N_1838);
nand U6439 (N_6439,N_3402,N_3641);
nor U6440 (N_6440,N_4314,N_117);
nor U6441 (N_6441,N_3116,N_4701);
or U6442 (N_6442,N_1976,N_1355);
nor U6443 (N_6443,N_3045,N_549);
nand U6444 (N_6444,N_3191,N_1146);
or U6445 (N_6445,N_818,N_4170);
or U6446 (N_6446,N_3026,N_2696);
nand U6447 (N_6447,N_4089,N_1827);
or U6448 (N_6448,N_720,N_2654);
nor U6449 (N_6449,N_336,N_1384);
and U6450 (N_6450,N_4474,N_2360);
nand U6451 (N_6451,N_2301,N_1869);
or U6452 (N_6452,N_3233,N_1169);
or U6453 (N_6453,N_1452,N_3909);
and U6454 (N_6454,N_77,N_3149);
or U6455 (N_6455,N_350,N_4248);
nor U6456 (N_6456,N_1115,N_4621);
nand U6457 (N_6457,N_4876,N_2218);
and U6458 (N_6458,N_972,N_3874);
nor U6459 (N_6459,N_1439,N_4298);
or U6460 (N_6460,N_1020,N_4321);
nand U6461 (N_6461,N_3643,N_610);
nor U6462 (N_6462,N_4723,N_1659);
nor U6463 (N_6463,N_3556,N_4241);
or U6464 (N_6464,N_151,N_1727);
or U6465 (N_6465,N_867,N_3210);
and U6466 (N_6466,N_2085,N_2459);
nand U6467 (N_6467,N_3204,N_2488);
or U6468 (N_6468,N_4076,N_2534);
nand U6469 (N_6469,N_2901,N_2277);
nor U6470 (N_6470,N_3758,N_3353);
nor U6471 (N_6471,N_191,N_2154);
nor U6472 (N_6472,N_2184,N_2783);
nor U6473 (N_6473,N_4108,N_1708);
and U6474 (N_6474,N_3236,N_2164);
or U6475 (N_6475,N_1296,N_3023);
nand U6476 (N_6476,N_756,N_3548);
nor U6477 (N_6477,N_3427,N_3304);
nand U6478 (N_6478,N_928,N_952);
nand U6479 (N_6479,N_1066,N_4502);
or U6480 (N_6480,N_3082,N_3035);
and U6481 (N_6481,N_3146,N_3667);
or U6482 (N_6482,N_3389,N_2236);
nand U6483 (N_6483,N_3864,N_1887);
nor U6484 (N_6484,N_4255,N_3685);
or U6485 (N_6485,N_3054,N_4520);
and U6486 (N_6486,N_3249,N_4629);
and U6487 (N_6487,N_1574,N_4171);
nand U6488 (N_6488,N_1012,N_3408);
and U6489 (N_6489,N_4939,N_3684);
and U6490 (N_6490,N_3780,N_173);
nand U6491 (N_6491,N_3066,N_2145);
nand U6492 (N_6492,N_4803,N_1692);
nor U6493 (N_6493,N_3532,N_3311);
or U6494 (N_6494,N_1690,N_1902);
or U6495 (N_6495,N_4070,N_2419);
nand U6496 (N_6496,N_3359,N_4836);
and U6497 (N_6497,N_1677,N_1541);
and U6498 (N_6498,N_848,N_4063);
and U6499 (N_6499,N_1430,N_4025);
or U6500 (N_6500,N_662,N_2461);
nand U6501 (N_6501,N_815,N_1728);
and U6502 (N_6502,N_3361,N_2007);
and U6503 (N_6503,N_4132,N_1250);
and U6504 (N_6504,N_3027,N_1212);
nand U6505 (N_6505,N_3582,N_4505);
and U6506 (N_6506,N_4027,N_827);
xnor U6507 (N_6507,N_4816,N_1554);
or U6508 (N_6508,N_249,N_2501);
xnor U6509 (N_6509,N_2205,N_3994);
nand U6510 (N_6510,N_3729,N_3610);
and U6511 (N_6511,N_3989,N_1358);
and U6512 (N_6512,N_4694,N_949);
nand U6513 (N_6513,N_4275,N_459);
nor U6514 (N_6514,N_4254,N_4164);
and U6515 (N_6515,N_403,N_3820);
nor U6516 (N_6516,N_2312,N_3821);
or U6517 (N_6517,N_1569,N_438);
nand U6518 (N_6518,N_381,N_1460);
nor U6519 (N_6519,N_3323,N_1395);
nor U6520 (N_6520,N_1137,N_4203);
or U6521 (N_6521,N_3143,N_988);
or U6522 (N_6522,N_1408,N_2903);
nor U6523 (N_6523,N_2220,N_3216);
nand U6524 (N_6524,N_4146,N_3330);
nand U6525 (N_6525,N_2661,N_4103);
or U6526 (N_6526,N_873,N_3088);
nor U6527 (N_6527,N_4689,N_2209);
nand U6528 (N_6528,N_566,N_2719);
nor U6529 (N_6529,N_1030,N_1888);
or U6530 (N_6530,N_4571,N_2284);
or U6531 (N_6531,N_1335,N_3605);
nor U6532 (N_6532,N_1004,N_3194);
and U6533 (N_6533,N_409,N_4760);
nor U6534 (N_6534,N_1247,N_441);
xnor U6535 (N_6535,N_481,N_4574);
nor U6536 (N_6536,N_640,N_3420);
nand U6537 (N_6537,N_740,N_4959);
and U6538 (N_6538,N_560,N_1078);
or U6539 (N_6539,N_2062,N_2529);
or U6540 (N_6540,N_3713,N_907);
and U6541 (N_6541,N_211,N_1853);
nand U6542 (N_6542,N_3032,N_109);
and U6543 (N_6543,N_3588,N_4539);
and U6544 (N_6544,N_3544,N_1209);
and U6545 (N_6545,N_624,N_38);
nor U6546 (N_6546,N_4963,N_4206);
and U6547 (N_6547,N_4919,N_922);
and U6548 (N_6548,N_2348,N_1150);
nor U6549 (N_6549,N_4780,N_3453);
nor U6550 (N_6550,N_1587,N_4642);
xnor U6551 (N_6551,N_3057,N_1595);
or U6552 (N_6552,N_1285,N_2467);
and U6553 (N_6553,N_2679,N_4382);
or U6554 (N_6554,N_2013,N_4771);
or U6555 (N_6555,N_3305,N_3313);
or U6556 (N_6556,N_2550,N_3284);
nor U6557 (N_6557,N_1187,N_1373);
or U6558 (N_6558,N_1230,N_3795);
or U6559 (N_6559,N_2865,N_3670);
and U6560 (N_6560,N_595,N_4223);
and U6561 (N_6561,N_1709,N_3406);
nor U6562 (N_6562,N_1689,N_3924);
nor U6563 (N_6563,N_165,N_926);
nand U6564 (N_6564,N_4344,N_3217);
and U6565 (N_6565,N_564,N_4713);
or U6566 (N_6566,N_2088,N_3288);
or U6567 (N_6567,N_4936,N_3275);
nand U6568 (N_6568,N_2265,N_1028);
and U6569 (N_6569,N_4966,N_385);
and U6570 (N_6570,N_4155,N_1704);
nor U6571 (N_6571,N_4525,N_1981);
and U6572 (N_6572,N_2796,N_3333);
or U6573 (N_6573,N_57,N_3022);
nand U6574 (N_6574,N_680,N_1836);
or U6575 (N_6575,N_31,N_3123);
xnor U6576 (N_6576,N_2772,N_3285);
nand U6577 (N_6577,N_2970,N_2556);
and U6578 (N_6578,N_434,N_39);
nand U6579 (N_6579,N_4225,N_4815);
nor U6580 (N_6580,N_1447,N_2227);
or U6581 (N_6581,N_14,N_2263);
nor U6582 (N_6582,N_1061,N_4400);
and U6583 (N_6583,N_1911,N_3617);
and U6584 (N_6584,N_1619,N_4735);
or U6585 (N_6585,N_4655,N_2379);
or U6586 (N_6586,N_4817,N_4324);
nand U6587 (N_6587,N_230,N_2927);
and U6588 (N_6588,N_3081,N_1624);
nand U6589 (N_6589,N_2226,N_4008);
nor U6590 (N_6590,N_2388,N_2751);
nand U6591 (N_6591,N_4699,N_2723);
nor U6592 (N_6592,N_3636,N_4148);
or U6593 (N_6593,N_2837,N_2981);
or U6594 (N_6594,N_1371,N_47);
or U6595 (N_6595,N_2101,N_2016);
nand U6596 (N_6596,N_1087,N_3946);
or U6597 (N_6597,N_4575,N_792);
nor U6598 (N_6598,N_358,N_2487);
and U6599 (N_6599,N_1625,N_4332);
or U6600 (N_6600,N_414,N_4419);
and U6601 (N_6601,N_4315,N_1936);
and U6602 (N_6602,N_452,N_1114);
nand U6603 (N_6603,N_984,N_960);
nand U6604 (N_6604,N_4407,N_3400);
or U6605 (N_6605,N_4166,N_732);
and U6606 (N_6606,N_2538,N_4302);
or U6607 (N_6607,N_4362,N_2091);
or U6608 (N_6608,N_1600,N_4618);
nor U6609 (N_6609,N_3138,N_4176);
nor U6610 (N_6610,N_4061,N_4940);
or U6611 (N_6611,N_3369,N_901);
nand U6612 (N_6612,N_3851,N_1324);
nor U6613 (N_6613,N_1470,N_4205);
nor U6614 (N_6614,N_4736,N_2194);
or U6615 (N_6615,N_2812,N_590);
and U6616 (N_6616,N_3270,N_2995);
nor U6617 (N_6617,N_1185,N_97);
and U6618 (N_6618,N_3324,N_1306);
and U6619 (N_6619,N_3537,N_1436);
nand U6620 (N_6620,N_4793,N_345);
nor U6621 (N_6621,N_547,N_1805);
nor U6622 (N_6622,N_1245,N_1638);
nand U6623 (N_6623,N_512,N_1021);
and U6624 (N_6624,N_224,N_1799);
nor U6625 (N_6625,N_4506,N_3985);
and U6626 (N_6626,N_941,N_3267);
nor U6627 (N_6627,N_616,N_4313);
and U6628 (N_6628,N_1594,N_3009);
or U6629 (N_6629,N_2943,N_2588);
and U6630 (N_6630,N_3940,N_3930);
nor U6631 (N_6631,N_1996,N_940);
and U6632 (N_6632,N_1027,N_3961);
or U6633 (N_6633,N_4635,N_2766);
and U6634 (N_6634,N_2673,N_4943);
nand U6635 (N_6635,N_3604,N_29);
nand U6636 (N_6636,N_3838,N_2408);
or U6637 (N_6637,N_656,N_2521);
and U6638 (N_6638,N_134,N_947);
or U6639 (N_6639,N_2519,N_1290);
and U6640 (N_6640,N_3929,N_2871);
or U6641 (N_6641,N_1721,N_2435);
nor U6642 (N_6642,N_3152,N_2171);
nor U6643 (N_6643,N_3979,N_4945);
and U6644 (N_6644,N_1062,N_3788);
nor U6645 (N_6645,N_3679,N_585);
or U6646 (N_6646,N_1192,N_4226);
or U6647 (N_6647,N_4881,N_4);
or U6648 (N_6648,N_2489,N_379);
or U6649 (N_6649,N_2094,N_2456);
nor U6650 (N_6650,N_751,N_2974);
and U6651 (N_6651,N_4730,N_2816);
or U6652 (N_6652,N_4808,N_3793);
or U6653 (N_6653,N_578,N_3467);
nand U6654 (N_6654,N_4521,N_3565);
and U6655 (N_6655,N_2305,N_3052);
nand U6656 (N_6656,N_1871,N_4317);
or U6657 (N_6657,N_120,N_2852);
nor U6658 (N_6658,N_81,N_4851);
nand U6659 (N_6659,N_397,N_3474);
nor U6660 (N_6660,N_4970,N_4619);
or U6661 (N_6661,N_1714,N_3268);
or U6662 (N_6662,N_4679,N_4975);
nor U6663 (N_6663,N_2651,N_3211);
nand U6664 (N_6664,N_1859,N_370);
nand U6665 (N_6665,N_1454,N_1913);
or U6666 (N_6666,N_3028,N_4566);
or U6667 (N_6667,N_1039,N_1477);
or U6668 (N_6668,N_1047,N_1343);
and U6669 (N_6669,N_3514,N_2838);
nor U6670 (N_6670,N_2178,N_3956);
or U6671 (N_6671,N_3848,N_1369);
or U6672 (N_6672,N_2197,N_3782);
nand U6673 (N_6673,N_1425,N_1602);
or U6674 (N_6674,N_772,N_4928);
or U6675 (N_6675,N_1670,N_2039);
nor U6676 (N_6676,N_217,N_1779);
and U6677 (N_6677,N_4232,N_3858);
nor U6678 (N_6678,N_3737,N_1538);
and U6679 (N_6679,N_2637,N_1079);
and U6680 (N_6680,N_446,N_3470);
and U6681 (N_6681,N_4117,N_3021);
or U6682 (N_6682,N_599,N_360);
nor U6683 (N_6683,N_4918,N_3703);
and U6684 (N_6684,N_2502,N_3993);
or U6685 (N_6685,N_4600,N_1729);
nor U6686 (N_6686,N_227,N_482);
nand U6687 (N_6687,N_1525,N_3396);
nand U6688 (N_6688,N_4353,N_1987);
and U6689 (N_6689,N_4884,N_672);
nand U6690 (N_6690,N_2671,N_1531);
or U6691 (N_6691,N_315,N_3916);
nor U6692 (N_6692,N_1180,N_3181);
nor U6693 (N_6693,N_2949,N_3917);
or U6694 (N_6694,N_2862,N_4261);
or U6695 (N_6695,N_3630,N_2122);
and U6696 (N_6696,N_538,N_3499);
or U6697 (N_6697,N_3852,N_2579);
nor U6698 (N_6698,N_1302,N_775);
nor U6699 (N_6699,N_2881,N_2406);
nor U6700 (N_6700,N_3910,N_4595);
or U6701 (N_6701,N_252,N_4807);
and U6702 (N_6702,N_2757,N_3180);
or U6703 (N_6703,N_4675,N_2809);
nor U6704 (N_6704,N_4325,N_2950);
or U6705 (N_6705,N_4201,N_3071);
nand U6706 (N_6706,N_2929,N_4994);
and U6707 (N_6707,N_268,N_1236);
or U6708 (N_6708,N_253,N_3746);
or U6709 (N_6709,N_3836,N_1119);
and U6710 (N_6710,N_3494,N_875);
nor U6711 (N_6711,N_834,N_13);
and U6712 (N_6712,N_4363,N_3849);
or U6713 (N_6713,N_2506,N_2685);
nor U6714 (N_6714,N_4094,N_3644);
nand U6715 (N_6715,N_1423,N_2956);
nor U6716 (N_6716,N_153,N_4917);
nor U6717 (N_6717,N_3107,N_548);
nand U6718 (N_6718,N_2800,N_935);
or U6719 (N_6719,N_4350,N_3187);
nand U6720 (N_6720,N_2872,N_1784);
and U6721 (N_6721,N_4116,N_3731);
xnor U6722 (N_6722,N_2513,N_4491);
nand U6723 (N_6723,N_4385,N_4839);
and U6724 (N_6724,N_4791,N_4712);
and U6725 (N_6725,N_493,N_1196);
and U6726 (N_6726,N_4870,N_4462);
or U6727 (N_6727,N_4790,N_2937);
and U6728 (N_6728,N_2782,N_2917);
nand U6729 (N_6729,N_1920,N_3166);
nand U6730 (N_6730,N_2325,N_1218);
or U6731 (N_6731,N_4210,N_2349);
or U6732 (N_6732,N_364,N_4838);
nand U6733 (N_6733,N_3545,N_1903);
or U6734 (N_6734,N_3655,N_2902);
nor U6735 (N_6735,N_1553,N_105);
nand U6736 (N_6736,N_2436,N_3403);
nor U6737 (N_6737,N_328,N_593);
or U6738 (N_6738,N_1839,N_2161);
or U6739 (N_6739,N_2735,N_4627);
and U6740 (N_6740,N_99,N_263);
nor U6741 (N_6741,N_4767,N_1444);
or U6742 (N_6742,N_4069,N_3775);
and U6743 (N_6743,N_214,N_8);
nor U6744 (N_6744,N_1546,N_1632);
nor U6745 (N_6745,N_3615,N_405);
or U6746 (N_6746,N_1287,N_4285);
xor U6747 (N_6747,N_3772,N_2138);
nor U6748 (N_6748,N_1183,N_2808);
nand U6749 (N_6749,N_3292,N_2689);
or U6750 (N_6750,N_525,N_1539);
or U6751 (N_6751,N_2199,N_2573);
nor U6752 (N_6752,N_1254,N_3337);
and U6753 (N_6753,N_2728,N_1364);
nand U6754 (N_6754,N_851,N_4951);
or U6755 (N_6755,N_2669,N_4461);
nand U6756 (N_6756,N_4187,N_3212);
and U6757 (N_6757,N_2670,N_1036);
and U6758 (N_6758,N_4335,N_1591);
or U6759 (N_6759,N_2140,N_4357);
or U6760 (N_6760,N_3067,N_2699);
or U6761 (N_6761,N_664,N_3856);
and U6762 (N_6762,N_61,N_3289);
or U6763 (N_6763,N_609,N_138);
and U6764 (N_6764,N_2792,N_2701);
nand U6765 (N_6765,N_84,N_1548);
and U6766 (N_6766,N_1483,N_2738);
nor U6767 (N_6767,N_2793,N_2666);
and U6768 (N_6768,N_836,N_4373);
and U6769 (N_6769,N_2278,N_4323);
nand U6770 (N_6770,N_4293,N_927);
or U6771 (N_6771,N_1995,N_4670);
nand U6772 (N_6772,N_431,N_208);
and U6773 (N_6773,N_2575,N_654);
or U6774 (N_6774,N_349,N_3507);
and U6775 (N_6775,N_2885,N_3053);
nor U6776 (N_6776,N_3020,N_4727);
or U6777 (N_6777,N_4265,N_3504);
or U6778 (N_6778,N_3597,N_702);
nor U6779 (N_6779,N_3201,N_285);
or U6780 (N_6780,N_174,N_789);
or U6781 (N_6781,N_289,N_2935);
nand U6782 (N_6782,N_1487,N_2918);
and U6783 (N_6783,N_3079,N_3042);
nand U6784 (N_6784,N_2715,N_724);
nand U6785 (N_6785,N_1002,N_3777);
nor U6786 (N_6786,N_4258,N_2632);
nor U6787 (N_6787,N_1921,N_237);
and U6788 (N_6788,N_1265,N_187);
and U6789 (N_6789,N_172,N_3255);
and U6790 (N_6790,N_3479,N_2156);
or U6791 (N_6791,N_1486,N_4773);
nor U6792 (N_6792,N_331,N_1990);
nor U6793 (N_6793,N_4530,N_2924);
and U6794 (N_6794,N_1764,N_3450);
nand U6795 (N_6795,N_3106,N_2163);
or U6796 (N_6796,N_3850,N_1116);
nand U6797 (N_6797,N_3570,N_3563);
nor U6798 (N_6798,N_3546,N_3762);
nand U6799 (N_6799,N_82,N_1806);
nor U6800 (N_6800,N_1529,N_4047);
nor U6801 (N_6801,N_4125,N_1648);
and U6802 (N_6802,N_3484,N_4997);
nand U6803 (N_6803,N_1586,N_4681);
or U6804 (N_6804,N_951,N_2609);
or U6805 (N_6805,N_954,N_1882);
nor U6806 (N_6806,N_3815,N_4608);
or U6807 (N_6807,N_2520,N_3294);
and U6808 (N_6808,N_3481,N_4593);
nor U6809 (N_6809,N_3172,N_1636);
and U6810 (N_6810,N_929,N_746);
nor U6811 (N_6811,N_2919,N_3939);
nand U6812 (N_6812,N_199,N_688);
nand U6813 (N_6813,N_1144,N_4931);
nor U6814 (N_6814,N_1429,N_4136);
nand U6815 (N_6815,N_4331,N_1365);
nand U6816 (N_6816,N_157,N_1605);
xnor U6817 (N_6817,N_4885,N_2242);
or U6818 (N_6818,N_1950,N_1518);
or U6819 (N_6819,N_2228,N_2566);
and U6820 (N_6820,N_1362,N_3839);
nand U6821 (N_6821,N_2734,N_641);
nor U6822 (N_6822,N_1410,N_4921);
and U6823 (N_6823,N_2933,N_4835);
nor U6824 (N_6824,N_2544,N_4122);
nor U6825 (N_6825,N_4766,N_4508);
nor U6826 (N_6826,N_3059,N_2044);
and U6827 (N_6827,N_842,N_905);
or U6828 (N_6828,N_4167,N_3151);
nor U6829 (N_6829,N_1825,N_1501);
nor U6830 (N_6830,N_429,N_1746);
nand U6831 (N_6831,N_2188,N_4175);
nor U6832 (N_6832,N_453,N_4786);
nor U6833 (N_6833,N_2930,N_685);
or U6834 (N_6834,N_2908,N_1753);
or U6835 (N_6835,N_1249,N_212);
and U6836 (N_6836,N_2692,N_2375);
or U6837 (N_6837,N_286,N_3639);
nor U6838 (N_6838,N_4303,N_98);
nand U6839 (N_6839,N_4680,N_3093);
or U6840 (N_6840,N_2597,N_2187);
nand U6841 (N_6841,N_2414,N_557);
nor U6842 (N_6842,N_4865,N_1988);
nor U6843 (N_6843,N_4045,N_1234);
nand U6844 (N_6844,N_2430,N_1459);
nor U6845 (N_6845,N_3707,N_1259);
or U6846 (N_6846,N_2108,N_1201);
nor U6847 (N_6847,N_1829,N_2306);
nor U6848 (N_6848,N_2567,N_2445);
and U6849 (N_6849,N_2438,N_4209);
nand U6850 (N_6850,N_4892,N_963);
or U6851 (N_6851,N_1332,N_2135);
or U6852 (N_6852,N_2614,N_4632);
and U6853 (N_6853,N_3863,N_2398);
and U6854 (N_6854,N_4224,N_4829);
and U6855 (N_6855,N_2877,N_4458);
or U6856 (N_6856,N_565,N_2672);
nand U6857 (N_6857,N_920,N_3257);
or U6858 (N_6858,N_4725,N_863);
or U6859 (N_6859,N_220,N_3890);
and U6860 (N_6860,N_2437,N_582);
nor U6861 (N_6861,N_3735,N_2980);
nor U6862 (N_6862,N_1432,N_2941);
and U6863 (N_6863,N_3063,N_2170);
and U6864 (N_6864,N_4974,N_3382);
or U6865 (N_6865,N_368,N_2075);
nand U6866 (N_6866,N_4356,N_3422);
nand U6867 (N_6867,N_3423,N_4021);
nor U6868 (N_6868,N_2875,N_1794);
nand U6869 (N_6869,N_2518,N_3796);
and U6870 (N_6870,N_1500,N_4149);
nor U6871 (N_6871,N_2056,N_4517);
nor U6872 (N_6872,N_3380,N_1227);
and U6873 (N_6873,N_2591,N_2329);
xnor U6874 (N_6874,N_4497,N_4217);
and U6875 (N_6875,N_2897,N_997);
and U6876 (N_6876,N_2703,N_4010);
or U6877 (N_6877,N_4444,N_4704);
nor U6878 (N_6878,N_4286,N_2358);
nor U6879 (N_6879,N_10,N_4673);
nor U6880 (N_6880,N_369,N_2102);
or U6881 (N_6881,N_1817,N_4268);
and U6882 (N_6882,N_4039,N_3846);
or U6883 (N_6883,N_2601,N_4251);
nor U6884 (N_6884,N_946,N_2818);
or U6885 (N_6885,N_1331,N_3466);
nor U6886 (N_6886,N_1559,N_3148);
and U6887 (N_6887,N_3339,N_991);
or U6888 (N_6888,N_4300,N_3677);
nor U6889 (N_6889,N_3274,N_46);
or U6890 (N_6890,N_3346,N_3520);
or U6891 (N_6891,N_3601,N_4080);
or U6892 (N_6892,N_967,N_3341);
and U6893 (N_6893,N_552,N_1701);
or U6894 (N_6894,N_2886,N_1732);
nand U6895 (N_6895,N_694,N_690);
nor U6896 (N_6896,N_3878,N_2879);
and U6897 (N_6897,N_1281,N_3905);
or U6898 (N_6898,N_272,N_974);
or U6899 (N_6899,N_3926,N_2867);
nand U6900 (N_6900,N_2077,N_1755);
or U6901 (N_6901,N_4059,N_607);
or U6902 (N_6902,N_4925,N_4624);
and U6903 (N_6903,N_297,N_1674);
or U6904 (N_6904,N_231,N_2874);
nor U6905 (N_6905,N_1232,N_4391);
nand U6906 (N_6906,N_353,N_1417);
or U6907 (N_6907,N_4312,N_3552);
nor U6908 (N_6908,N_1907,N_4471);
xnor U6909 (N_6909,N_3709,N_581);
and U6910 (N_6910,N_4020,N_3024);
nand U6911 (N_6911,N_3368,N_470);
nand U6912 (N_6912,N_4493,N_3083);
nand U6913 (N_6913,N_4837,N_2400);
or U6914 (N_6914,N_2055,N_706);
nor U6915 (N_6915,N_1333,N_4375);
nand U6916 (N_6916,N_4445,N_878);
and U6917 (N_6917,N_4304,N_4806);
and U6918 (N_6918,N_4238,N_1616);
nor U6919 (N_6919,N_2987,N_1952);
nor U6920 (N_6920,N_2714,N_3987);
nand U6921 (N_6921,N_3710,N_2571);
and U6922 (N_6922,N_4120,N_2802);
and U6923 (N_6923,N_644,N_1159);
nor U6924 (N_6924,N_4903,N_1530);
and U6925 (N_6925,N_1437,N_3340);
nand U6926 (N_6926,N_3101,N_3141);
and U6927 (N_6927,N_3973,N_4649);
or U6928 (N_6928,N_4753,N_3932);
or U6929 (N_6929,N_4456,N_215);
and U6930 (N_6930,N_3209,N_2634);
and U6931 (N_6931,N_4676,N_3246);
nand U6932 (N_6932,N_1440,N_1208);
nor U6933 (N_6933,N_4914,N_691);
nor U6934 (N_6934,N_28,N_4858);
and U6935 (N_6935,N_416,N_0);
or U6936 (N_6936,N_1770,N_2384);
nor U6937 (N_6937,N_3301,N_1366);
and U6938 (N_6938,N_1883,N_3580);
nand U6939 (N_6939,N_3892,N_3395);
and U6940 (N_6940,N_4367,N_4788);
or U6941 (N_6941,N_1330,N_3253);
and U6942 (N_6942,N_4732,N_4768);
or U6943 (N_6943,N_762,N_1686);
nor U6944 (N_6944,N_2565,N_3749);
nor U6945 (N_6945,N_3327,N_3008);
and U6946 (N_6946,N_2665,N_3192);
or U6947 (N_6947,N_697,N_196);
nor U6948 (N_6948,N_260,N_1172);
nand U6949 (N_6949,N_3559,N_261);
nand U6950 (N_6950,N_886,N_366);
xnor U6951 (N_6951,N_2633,N_2237);
or U6952 (N_6952,N_4092,N_1923);
or U6953 (N_6953,N_4762,N_2411);
nor U6954 (N_6954,N_1083,N_85);
xnor U6955 (N_6955,N_3895,N_4392);
or U6956 (N_6956,N_3902,N_2973);
nor U6957 (N_6957,N_2470,N_3754);
nand U6958 (N_6958,N_4211,N_2134);
nor U6959 (N_6959,N_4057,N_3468);
or U6960 (N_6960,N_3259,N_3338);
nor U6961 (N_6961,N_4582,N_1705);
and U6962 (N_6962,N_114,N_1041);
or U6963 (N_6963,N_859,N_501);
or U6964 (N_6964,N_3051,N_4700);
nand U6965 (N_6965,N_3404,N_2500);
or U6966 (N_6966,N_1042,N_945);
and U6967 (N_6967,N_4074,N_2381);
or U6968 (N_6968,N_3085,N_2374);
and U6969 (N_6969,N_2394,N_4879);
or U6970 (N_6970,N_4687,N_1441);
and U6971 (N_6971,N_4953,N_352);
nand U6972 (N_6972,N_3214,N_4833);
nand U6973 (N_6973,N_2807,N_4652);
and U6974 (N_6974,N_20,N_4853);
nor U6975 (N_6975,N_4402,N_1164);
nand U6976 (N_6976,N_1129,N_1481);
nand U6977 (N_6977,N_1448,N_2824);
nor U6978 (N_6978,N_2810,N_2359);
and U6979 (N_6979,N_1431,N_3595);
and U6980 (N_6980,N_1175,N_4616);
nand U6981 (N_6981,N_808,N_3893);
nand U6982 (N_6982,N_601,N_1615);
nor U6983 (N_6983,N_916,N_4399);
nand U6984 (N_6984,N_1556,N_3675);
nand U6985 (N_6985,N_3345,N_2957);
or U6986 (N_6986,N_490,N_3179);
nand U6987 (N_6987,N_2117,N_4981);
or U6988 (N_6988,N_4364,N_4572);
nand U6989 (N_6989,N_647,N_2822);
and U6990 (N_6990,N_4871,N_4950);
and U6991 (N_6991,N_4784,N_465);
or U6992 (N_6992,N_3170,N_3678);
nor U6993 (N_6993,N_1718,N_4650);
nand U6994 (N_6994,N_4733,N_1082);
xor U6995 (N_6995,N_1253,N_30);
nor U6996 (N_6996,N_4910,N_715);
and U6997 (N_6997,N_2481,N_1499);
xnor U6998 (N_6998,N_3482,N_3770);
nand U6999 (N_6999,N_3833,N_4107);
nand U7000 (N_7000,N_2357,N_2131);
nor U7001 (N_7001,N_4048,N_2009);
nand U7002 (N_7002,N_1653,N_1446);
nor U7003 (N_7003,N_497,N_1336);
nor U7004 (N_7004,N_3094,N_1813);
nand U7005 (N_7005,N_450,N_4040);
or U7006 (N_7006,N_860,N_4159);
nor U7007 (N_7007,N_2582,N_2942);
nor U7008 (N_7008,N_3606,N_222);
nand U7009 (N_7009,N_2841,N_2911);
nor U7010 (N_7010,N_892,N_76);
nor U7011 (N_7011,N_1719,N_2059);
or U7012 (N_7012,N_1819,N_422);
nand U7013 (N_7013,N_3920,N_1504);
nand U7014 (N_7014,N_3508,N_2018);
nand U7015 (N_7015,N_3440,N_838);
nor U7016 (N_7016,N_3518,N_3360);
or U7017 (N_7017,N_4570,N_2146);
and U7018 (N_7018,N_204,N_177);
nor U7019 (N_7019,N_1696,N_175);
nor U7020 (N_7020,N_2944,N_3827);
and U7021 (N_7021,N_3203,N_4612);
nand U7022 (N_7022,N_2416,N_3991);
and U7023 (N_7023,N_455,N_3480);
and U7024 (N_7024,N_247,N_4207);
or U7025 (N_7025,N_4555,N_4404);
xor U7026 (N_7026,N_326,N_3867);
nand U7027 (N_7027,N_894,N_2663);
and U7028 (N_7028,N_4856,N_3889);
nor U7029 (N_7029,N_3018,N_238);
nor U7030 (N_7030,N_228,N_2377);
nand U7031 (N_7031,N_1763,N_1397);
and U7032 (N_7032,N_2998,N_2222);
or U7033 (N_7033,N_2110,N_2261);
nor U7034 (N_7034,N_4234,N_1387);
and U7035 (N_7035,N_3265,N_2729);
nand U7036 (N_7036,N_2003,N_4137);
xor U7037 (N_7037,N_15,N_1060);
nor U7038 (N_7038,N_2160,N_4964);
nand U7039 (N_7039,N_4093,N_4372);
nor U7040 (N_7040,N_2276,N_652);
nor U7041 (N_7041,N_3525,N_1933);
or U7042 (N_7042,N_3439,N_3747);
and U7043 (N_7043,N_80,N_283);
nor U7044 (N_7044,N_3800,N_4055);
or U7045 (N_7045,N_4169,N_4741);
and U7046 (N_7046,N_146,N_2269);
or U7047 (N_7047,N_2899,N_2450);
nor U7048 (N_7048,N_831,N_178);
or U7049 (N_7049,N_665,N_1393);
and U7050 (N_7050,N_4625,N_4387);
nor U7051 (N_7051,N_2921,N_4044);
or U7052 (N_7052,N_2584,N_1110);
or U7053 (N_7053,N_710,N_4415);
nor U7054 (N_7054,N_948,N_1125);
nor U7055 (N_7055,N_69,N_2720);
nor U7056 (N_7056,N_2247,N_3562);
nor U7057 (N_7057,N_3691,N_1807);
or U7058 (N_7058,N_2621,N_346);
and U7059 (N_7059,N_411,N_4685);
nor U7060 (N_7060,N_70,N_3102);
or U7061 (N_7061,N_1848,N_1256);
nand U7062 (N_7062,N_1895,N_856);
nor U7063 (N_7063,N_2155,N_3593);
nand U7064 (N_7064,N_3036,N_2268);
nor U7065 (N_7065,N_1072,N_3988);
nor U7066 (N_7066,N_1048,N_4359);
and U7067 (N_7067,N_2979,N_2054);
nand U7068 (N_7068,N_797,N_1228);
nand U7069 (N_7069,N_2652,N_3502);
nor U7070 (N_7070,N_1517,N_4834);
nand U7071 (N_7071,N_760,N_620);
or U7072 (N_7072,N_4014,N_2468);
nand U7073 (N_7073,N_553,N_4228);
or U7074 (N_7074,N_3430,N_4785);
or U7075 (N_7075,N_1406,N_4717);
and U7076 (N_7076,N_3283,N_4899);
xor U7077 (N_7077,N_3163,N_2048);
and U7078 (N_7078,N_826,N_2484);
and U7079 (N_7079,N_439,N_3911);
and U7080 (N_7080,N_3476,N_3626);
and U7081 (N_7081,N_879,N_2376);
and U7082 (N_7082,N_1199,N_2410);
or U7083 (N_7083,N_4188,N_943);
or U7084 (N_7084,N_4291,N_1724);
nand U7085 (N_7085,N_1769,N_1868);
and U7086 (N_7086,N_229,N_4054);
and U7087 (N_7087,N_2201,N_1747);
and U7088 (N_7088,N_1354,N_371);
nand U7089 (N_7089,N_2250,N_4294);
or U7090 (N_7090,N_1664,N_4937);
or U7091 (N_7091,N_2196,N_1323);
and U7092 (N_7092,N_1415,N_301);
or U7093 (N_7093,N_554,N_2289);
nor U7094 (N_7094,N_2922,N_2251);
and U7095 (N_7095,N_1000,N_4711);
nand U7096 (N_7096,N_363,N_50);
or U7097 (N_7097,N_791,N_4383);
nor U7098 (N_7098,N_2514,N_180);
or U7099 (N_7099,N_2082,N_1097);
nor U7100 (N_7100,N_3073,N_1312);
nand U7101 (N_7101,N_2509,N_294);
nand U7102 (N_7102,N_4799,N_1930);
nor U7103 (N_7103,N_2245,N_3348);
nor U7104 (N_7104,N_1944,N_495);
nor U7105 (N_7105,N_3871,N_4849);
nand U7106 (N_7106,N_2823,N_3013);
nand U7107 (N_7107,N_4339,N_3845);
and U7108 (N_7108,N_25,N_858);
nor U7109 (N_7109,N_3629,N_4078);
or U7110 (N_7110,N_367,N_1822);
and U7111 (N_7111,N_2895,N_4544);
nor U7112 (N_7112,N_2351,N_4301);
and U7113 (N_7113,N_1583,N_437);
nor U7114 (N_7114,N_3937,N_4379);
nand U7115 (N_7115,N_1107,N_487);
or U7116 (N_7116,N_325,N_334);
nor U7117 (N_7117,N_2330,N_3089);
or U7118 (N_7118,N_1833,N_1751);
and U7119 (N_7119,N_4129,N_135);
and U7120 (N_7120,N_1316,N_3555);
or U7121 (N_7121,N_686,N_4900);
nand U7122 (N_7122,N_3090,N_3290);
nand U7123 (N_7123,N_3417,N_707);
and U7124 (N_7124,N_1949,N_3173);
and U7125 (N_7125,N_2664,N_617);
nor U7126 (N_7126,N_3425,N_1924);
and U7127 (N_7127,N_2103,N_4872);
or U7128 (N_7128,N_1916,N_1109);
xnor U7129 (N_7129,N_3688,N_4253);
nand U7130 (N_7130,N_262,N_2517);
nand U7131 (N_7131,N_2126,N_1205);
or U7132 (N_7132,N_4564,N_767);
or U7133 (N_7133,N_942,N_3832);
nand U7134 (N_7134,N_2120,N_2945);
or U7135 (N_7135,N_2174,N_1792);
nor U7136 (N_7136,N_3287,N_3419);
nor U7137 (N_7137,N_2309,N_3519);
nand U7138 (N_7138,N_1971,N_1238);
nor U7139 (N_7139,N_1367,N_668);
nor U7140 (N_7140,N_4573,N_3055);
nor U7141 (N_7141,N_567,N_1189);
nor U7142 (N_7142,N_62,N_4082);
or U7143 (N_7143,N_4969,N_3665);
xnor U7144 (N_7144,N_4147,N_1194);
or U7145 (N_7145,N_4978,N_1778);
or U7146 (N_7146,N_3366,N_3841);
nor U7147 (N_7147,N_1775,N_3007);
or U7148 (N_7148,N_2713,N_281);
and U7149 (N_7149,N_4633,N_3443);
or U7150 (N_7150,N_2983,N_4219);
nor U7151 (N_7151,N_56,N_3296);
or U7152 (N_7152,N_3454,N_1389);
or U7153 (N_7153,N_3922,N_4998);
or U7154 (N_7154,N_2524,N_1652);
nand U7155 (N_7155,N_4976,N_1565);
nor U7156 (N_7156,N_978,N_3031);
or U7157 (N_7157,N_2215,N_768);
or U7158 (N_7158,N_1492,N_938);
nand U7159 (N_7159,N_4898,N_3392);
or U7160 (N_7160,N_2303,N_3990);
nand U7161 (N_7161,N_4478,N_3219);
nand U7162 (N_7162,N_4098,N_2954);
nand U7163 (N_7163,N_4636,N_169);
and U7164 (N_7164,N_4282,N_59);
and U7165 (N_7165,N_3503,N_1643);
and U7166 (N_7166,N_1641,N_4821);
or U7167 (N_7167,N_4434,N_4498);
nand U7168 (N_7168,N_1945,N_518);
or U7169 (N_7169,N_4394,N_26);
and U7170 (N_7170,N_1089,N_432);
or U7171 (N_7171,N_159,N_3483);
nor U7172 (N_7172,N_4436,N_3437);
or U7173 (N_7173,N_631,N_648);
or U7174 (N_7174,N_112,N_4841);
and U7175 (N_7175,N_2127,N_1221);
and U7176 (N_7176,N_1723,N_4106);
nor U7177 (N_7177,N_1476,N_1842);
nand U7178 (N_7178,N_2593,N_981);
and U7179 (N_7179,N_1798,N_4161);
and U7180 (N_7180,N_4189,N_2993);
and U7181 (N_7181,N_94,N_2010);
nand U7182 (N_7182,N_2326,N_1482);
nor U7183 (N_7183,N_3215,N_843);
nand U7184 (N_7184,N_3753,N_2248);
and U7185 (N_7185,N_755,N_3577);
or U7186 (N_7186,N_3309,N_1277);
and U7187 (N_7187,N_1385,N_1303);
nor U7188 (N_7188,N_3130,N_3913);
or U7189 (N_7189,N_1617,N_2371);
or U7190 (N_7190,N_1497,N_4553);
or U7191 (N_7191,N_2574,N_4320);
nand U7192 (N_7192,N_765,N_2217);
nand U7193 (N_7193,N_4256,N_3070);
nand U7194 (N_7194,N_3676,N_3431);
and U7195 (N_7195,N_4389,N_168);
nor U7196 (N_7196,N_390,N_4977);
nand U7197 (N_7197,N_4657,N_1267);
or U7198 (N_7198,N_1210,N_1947);
nor U7199 (N_7199,N_1890,N_3645);
nand U7200 (N_7200,N_3349,N_1282);
or U7201 (N_7201,N_4863,N_3551);
or U7202 (N_7202,N_3448,N_100);
and U7203 (N_7203,N_957,N_3429);
nor U7204 (N_7204,N_4855,N_531);
nand U7205 (N_7205,N_2819,N_1435);
nor U7206 (N_7206,N_4281,N_2206);
nand U7207 (N_7207,N_1620,N_4499);
and U7208 (N_7208,N_4215,N_2451);
nand U7209 (N_7209,N_320,N_3086);
nand U7210 (N_7210,N_890,N_3816);
nor U7211 (N_7211,N_1304,N_2270);
or U7212 (N_7212,N_3316,N_2863);
nor U7213 (N_7213,N_2057,N_2383);
and U7214 (N_7214,N_4240,N_3631);
nor U7215 (N_7215,N_1680,N_2186);
and U7216 (N_7216,N_4348,N_1844);
or U7217 (N_7217,N_4719,N_2928);
nand U7218 (N_7218,N_3633,N_258);
nor U7219 (N_7219,N_4515,N_888);
or U7220 (N_7220,N_1870,N_4818);
or U7221 (N_7221,N_996,N_305);
and U7222 (N_7222,N_2635,N_2294);
or U7223 (N_7223,N_2777,N_1268);
nor U7224 (N_7224,N_1341,N_4935);
or U7225 (N_7225,N_3230,N_2736);
and U7226 (N_7226,N_2353,N_3176);
or U7227 (N_7227,N_463,N_635);
nand U7228 (N_7228,N_2457,N_1132);
and U7229 (N_7229,N_4145,N_517);
nand U7230 (N_7230,N_4483,N_2180);
nor U7231 (N_7231,N_4842,N_2682);
nor U7232 (N_7232,N_3574,N_1611);
nand U7233 (N_7233,N_2271,N_2495);
or U7234 (N_7234,N_4658,N_3959);
nor U7235 (N_7235,N_49,N_2012);
and U7236 (N_7236,N_4446,N_4745);
nand U7237 (N_7237,N_342,N_695);
or U7238 (N_7238,N_3915,N_2684);
or U7239 (N_7239,N_275,N_3240);
and U7240 (N_7240,N_2989,N_2073);
nand U7241 (N_7241,N_865,N_1181);
and U7242 (N_7242,N_1351,N_4133);
and U7243 (N_7243,N_4417,N_2667);
nand U7244 (N_7244,N_3325,N_3208);
nand U7245 (N_7245,N_2784,N_3862);
or U7246 (N_7246,N_721,N_2299);
nand U7247 (N_7247,N_3322,N_2195);
nor U7248 (N_7248,N_4971,N_464);
or U7249 (N_7249,N_4875,N_2623);
and U7250 (N_7250,N_3756,N_462);
and U7251 (N_7251,N_1240,N_4096);
and U7252 (N_7252,N_2647,N_4691);
or U7253 (N_7253,N_323,N_2920);
xnor U7254 (N_7254,N_3464,N_3723);
or U7255 (N_7255,N_2382,N_2322);
nand U7256 (N_7256,N_1368,N_3326);
nand U7257 (N_7257,N_1017,N_1896);
or U7258 (N_7258,N_3243,N_4889);
nor U7259 (N_7259,N_2293,N_78);
nor U7260 (N_7260,N_2169,N_2748);
nand U7261 (N_7261,N_203,N_806);
and U7262 (N_7262,N_2300,N_137);
nand U7263 (N_7263,N_402,N_2264);
nand U7264 (N_7264,N_1820,N_2119);
nand U7265 (N_7265,N_1023,N_4886);
nand U7266 (N_7266,N_133,N_2996);
and U7267 (N_7267,N_2733,N_3868);
or U7268 (N_7268,N_2790,N_2395);
nand U7269 (N_7269,N_1514,N_4360);
nor U7270 (N_7270,N_1814,N_3995);
nor U7271 (N_7271,N_4496,N_1418);
and U7272 (N_7272,N_4547,N_4589);
or U7273 (N_7273,N_2649,N_4199);
nor U7274 (N_7274,N_4756,N_1610);
and U7275 (N_7275,N_2290,N_3734);
nor U7276 (N_7276,N_4180,N_1096);
nand U7277 (N_7277,N_976,N_956);
nor U7278 (N_7278,N_1558,N_3923);
nor U7279 (N_7279,N_3232,N_1977);
and U7280 (N_7280,N_3475,N_1773);
nor U7281 (N_7281,N_2753,N_810);
nand U7282 (N_7282,N_2031,N_24);
nand U7283 (N_7283,N_598,N_1757);
nor U7284 (N_7284,N_4101,N_4467);
and U7285 (N_7285,N_4245,N_313);
and U7286 (N_7286,N_4742,N_91);
and U7287 (N_7287,N_343,N_2240);
nor U7288 (N_7288,N_3144,N_2613);
or U7289 (N_7289,N_1037,N_248);
and U7290 (N_7290,N_4567,N_71);
nor U7291 (N_7291,N_3397,N_3784);
and U7292 (N_7292,N_4023,N_2815);
nor U7293 (N_7293,N_561,N_1073);
or U7294 (N_7294,N_4439,N_4947);
nor U7295 (N_7295,N_193,N_1280);
and U7296 (N_7296,N_4623,N_611);
and U7297 (N_7297,N_4468,N_2449);
nand U7298 (N_7298,N_1927,N_866);
nand U7299 (N_7299,N_3347,N_226);
nor U7300 (N_7300,N_3242,N_1939);
and U7301 (N_7301,N_2402,N_2203);
nand U7302 (N_7302,N_3115,N_2355);
or U7303 (N_7303,N_2849,N_3513);
nand U7304 (N_7304,N_4250,N_1381);
xor U7305 (N_7305,N_4667,N_3050);
and U7306 (N_7306,N_4184,N_1637);
and U7307 (N_7307,N_2428,N_521);
and U7308 (N_7308,N_3407,N_1925);
and U7309 (N_7309,N_1168,N_541);
xnor U7310 (N_7310,N_400,N_2608);
and U7311 (N_7311,N_1932,N_2561);
nand U7312 (N_7312,N_86,N_3750);
or U7313 (N_7313,N_1166,N_194);
and U7314 (N_7314,N_4845,N_2207);
nor U7315 (N_7315,N_3566,N_1640);
nor U7316 (N_7316,N_1112,N_1834);
and U7317 (N_7317,N_955,N_1544);
or U7318 (N_7318,N_2019,N_4213);
nor U7319 (N_7319,N_2321,N_4151);
nor U7320 (N_7320,N_784,N_337);
and U7321 (N_7321,N_909,N_23);
and U7322 (N_7322,N_2549,N_3363);
nand U7323 (N_7323,N_2587,N_3384);
and U7324 (N_7324,N_445,N_2185);
or U7325 (N_7325,N_592,N_4854);
or U7326 (N_7326,N_3897,N_2762);
or U7327 (N_7327,N_603,N_4560);
nand U7328 (N_7328,N_4075,N_2697);
and U7329 (N_7329,N_1758,N_4289);
or U7330 (N_7330,N_3128,N_4157);
and U7331 (N_7331,N_4342,N_4512);
nor U7332 (N_7332,N_4451,N_2910);
or U7333 (N_7333,N_515,N_201);
nand U7334 (N_7334,N_1453,N_4153);
or U7335 (N_7335,N_2368,N_4528);
or U7336 (N_7336,N_64,N_2653);
and U7337 (N_7337,N_1502,N_1120);
nand U7338 (N_7338,N_1899,N_4361);
and U7339 (N_7339,N_130,N_4386);
nor U7340 (N_7340,N_636,N_4584);
nor U7341 (N_7341,N_3118,N_444);
and U7342 (N_7342,N_4368,N_2704);
nand U7343 (N_7343,N_1103,N_1537);
and U7344 (N_7344,N_4988,N_4648);
or U7345 (N_7345,N_2346,N_667);
and U7346 (N_7346,N_2052,N_3964);
or U7347 (N_7347,N_3175,N_1993);
nor U7348 (N_7348,N_4765,N_3060);
nand U7349 (N_7349,N_235,N_4306);
nor U7350 (N_7350,N_923,N_1785);
and U7351 (N_7351,N_4084,N_2947);
or U7352 (N_7352,N_4604,N_1121);
nor U7353 (N_7353,N_1200,N_2460);
nand U7354 (N_7354,N_4778,N_1058);
or U7355 (N_7355,N_1984,N_3854);
and U7356 (N_7356,N_3654,N_3883);
or U7357 (N_7357,N_2737,N_1024);
nor U7358 (N_7358,N_1866,N_2434);
and U7359 (N_7359,N_499,N_4653);
nor U7360 (N_7360,N_280,N_3957);
or U7361 (N_7361,N_3489,N_530);
or U7362 (N_7362,N_4423,N_4426);
nor U7363 (N_7363,N_3635,N_4121);
nand U7364 (N_7364,N_4538,N_693);
or U7365 (N_7365,N_2836,N_4764);
nor U7366 (N_7366,N_3682,N_4038);
nand U7367 (N_7367,N_2027,N_4024);
xnor U7368 (N_7368,N_1661,N_4877);
and U7369 (N_7369,N_577,N_1669);
nor U7370 (N_7370,N_3726,N_4427);
and U7371 (N_7371,N_726,N_356);
and U7372 (N_7372,N_4949,N_1742);
nand U7373 (N_7373,N_2043,N_2780);
nand U7374 (N_7374,N_433,N_2503);
nor U7375 (N_7375,N_2592,N_3047);
and U7376 (N_7376,N_1797,N_136);
and U7377 (N_7377,N_2702,N_738);
or U7378 (N_7378,N_3320,N_1224);
or U7379 (N_7379,N_1244,N_232);
nand U7380 (N_7380,N_1948,N_2727);
nor U7381 (N_7381,N_2900,N_2087);
and U7382 (N_7382,N_4522,N_1013);
and U7383 (N_7383,N_4545,N_1235);
nand U7384 (N_7384,N_805,N_671);
nor U7385 (N_7385,N_1443,N_2446);
and U7386 (N_7386,N_2982,N_149);
and U7387 (N_7387,N_2803,N_3687);
nand U7388 (N_7388,N_514,N_4929);
or U7389 (N_7389,N_3521,N_1217);
nand U7390 (N_7390,N_1873,N_1841);
and U7391 (N_7391,N_801,N_95);
nand U7392 (N_7392,N_1156,N_1305);
nand U7393 (N_7393,N_820,N_3303);
nor U7394 (N_7394,N_3438,N_4088);
and U7395 (N_7395,N_3405,N_4518);
and U7396 (N_7396,N_3578,N_4688);
nand U7397 (N_7397,N_4651,N_2686);
nand U7398 (N_7398,N_473,N_2084);
nand U7399 (N_7399,N_2399,N_2192);
and U7400 (N_7400,N_1858,N_267);
or U7401 (N_7401,N_1161,N_1379);
nor U7402 (N_7402,N_1781,N_2821);
and U7403 (N_7403,N_1526,N_278);
and U7404 (N_7404,N_1466,N_3033);
and U7405 (N_7405,N_4273,N_3251);
and U7406 (N_7406,N_868,N_795);
or U7407 (N_7407,N_2257,N_4135);
nand U7408 (N_7408,N_673,N_2121);
or U7409 (N_7409,N_4777,N_3096);
or U7410 (N_7410,N_2677,N_1566);
nor U7411 (N_7411,N_1170,N_2152);
and U7412 (N_7412,N_1480,N_4480);
nor U7413 (N_7413,N_771,N_1552);
nand U7414 (N_7414,N_2478,N_18);
nand U7415 (N_7415,N_3164,N_1135);
and U7416 (N_7416,N_2323,N_3842);
or U7417 (N_7417,N_2708,N_3538);
and U7418 (N_7418,N_1568,N_3248);
or U7419 (N_7419,N_1738,N_2232);
nand U7420 (N_7420,N_89,N_3786);
nand U7421 (N_7421,N_2540,N_1269);
or U7422 (N_7422,N_3002,N_745);
nand U7423 (N_7423,N_3491,N_3632);
nand U7424 (N_7424,N_3077,N_588);
and U7425 (N_7425,N_4562,N_2798);
nor U7426 (N_7426,N_2898,N_3019);
and U7427 (N_7427,N_460,N_3613);
nor U7428 (N_7428,N_2212,N_987);
nor U7429 (N_7429,N_4634,N_4843);
nand U7430 (N_7430,N_661,N_2876);
nor U7431 (N_7431,N_597,N_48);
or U7432 (N_7432,N_3119,N_4781);
and U7433 (N_7433,N_4722,N_2963);
nand U7434 (N_7434,N_4565,N_2307);
nor U7435 (N_7435,N_2962,N_1095);
nand U7436 (N_7436,N_2602,N_4015);
and U7437 (N_7437,N_4358,N_1214);
or U7438 (N_7438,N_830,N_2234);
nor U7439 (N_7439,N_2142,N_1248);
and U7440 (N_7440,N_1854,N_1390);
or U7441 (N_7441,N_3702,N_1134);
nand U7442 (N_7442,N_2243,N_4607);
nor U7443 (N_7443,N_998,N_982);
nor U7444 (N_7444,N_4614,N_3810);
nand U7445 (N_7445,N_4996,N_312);
or U7446 (N_7446,N_3773,N_692);
or U7447 (N_7447,N_3834,N_3925);
and U7448 (N_7448,N_1148,N_1631);
nand U7449 (N_7449,N_264,N_766);
nor U7450 (N_7450,N_4526,N_2546);
and U7451 (N_7451,N_3139,N_4558);
nand U7452 (N_7452,N_4100,N_1812);
or U7453 (N_7453,N_2491,N_4734);
nand U7454 (N_7454,N_3321,N_1767);
or U7455 (N_7455,N_4501,N_1307);
nand U7456 (N_7456,N_4309,N_4150);
or U7457 (N_7457,N_2335,N_2605);
and U7458 (N_7458,N_2854,N_1940);
nor U7459 (N_7459,N_1360,N_3590);
and U7460 (N_7460,N_1672,N_2976);
or U7461 (N_7461,N_3587,N_3573);
or U7462 (N_7462,N_2776,N_3254);
nor U7463 (N_7463,N_355,N_719);
and U7464 (N_7464,N_2069,N_3237);
nor U7465 (N_7465,N_2553,N_1455);
nand U7466 (N_7466,N_1113,N_4041);
nor U7467 (N_7467,N_4336,N_4168);
or U7468 (N_7468,N_4860,N_2046);
nor U7469 (N_7469,N_3199,N_4214);
and U7470 (N_7470,N_4043,N_4647);
and U7471 (N_7471,N_714,N_1532);
or U7472 (N_7472,N_125,N_4264);
xnor U7473 (N_7473,N_1760,N_2061);
nand U7474 (N_7474,N_4759,N_380);
and U7475 (N_7475,N_2526,N_2678);
nand U7476 (N_7476,N_4235,N_4548);
nand U7477 (N_7477,N_1327,N_4660);
nor U7478 (N_7478,N_2893,N_500);
and U7479 (N_7479,N_2604,N_1606);
and U7480 (N_7480,N_1370,N_2208);
nor U7481 (N_7481,N_1292,N_3646);
and U7482 (N_7482,N_1745,N_3853);
and U7483 (N_7483,N_800,N_3982);
and U7484 (N_7484,N_3221,N_3137);
nand U7485 (N_7485,N_2464,N_1576);
nor U7486 (N_7486,N_4484,N_1707);
and U7487 (N_7487,N_3127,N_3043);
nor U7488 (N_7488,N_3037,N_296);
nor U7489 (N_7489,N_2811,N_3312);
and U7490 (N_7490,N_4130,N_67);
and U7491 (N_7491,N_3761,N_4453);
or U7492 (N_7492,N_4598,N_2249);
and U7493 (N_7493,N_3113,N_3744);
or U7494 (N_7494,N_934,N_3706);
xor U7495 (N_7495,N_2615,N_4266);
or U7496 (N_7496,N_1961,N_2953);
nand U7497 (N_7497,N_3718,N_1800);
or U7498 (N_7498,N_1563,N_2641);
and U7499 (N_7499,N_234,N_4999);
xnor U7500 (N_7500,N_3338,N_2382);
nand U7501 (N_7501,N_3992,N_2706);
or U7502 (N_7502,N_314,N_2756);
nor U7503 (N_7503,N_3550,N_3975);
or U7504 (N_7504,N_3477,N_1702);
or U7505 (N_7505,N_3562,N_249);
nor U7506 (N_7506,N_3098,N_2193);
or U7507 (N_7507,N_3373,N_4990);
nor U7508 (N_7508,N_620,N_3267);
nand U7509 (N_7509,N_1947,N_2894);
or U7510 (N_7510,N_3684,N_3110);
nor U7511 (N_7511,N_3317,N_4549);
xnor U7512 (N_7512,N_3536,N_1391);
or U7513 (N_7513,N_590,N_556);
or U7514 (N_7514,N_3945,N_3706);
nor U7515 (N_7515,N_4192,N_1970);
and U7516 (N_7516,N_3857,N_3194);
and U7517 (N_7517,N_2285,N_4640);
and U7518 (N_7518,N_3138,N_769);
nor U7519 (N_7519,N_2579,N_4957);
nor U7520 (N_7520,N_3605,N_3741);
nand U7521 (N_7521,N_3069,N_2107);
nand U7522 (N_7522,N_4625,N_4324);
nor U7523 (N_7523,N_460,N_1024);
or U7524 (N_7524,N_1600,N_3943);
nor U7525 (N_7525,N_4951,N_3381);
nand U7526 (N_7526,N_24,N_4714);
or U7527 (N_7527,N_22,N_2902);
and U7528 (N_7528,N_209,N_3935);
and U7529 (N_7529,N_485,N_777);
or U7530 (N_7530,N_1494,N_850);
or U7531 (N_7531,N_274,N_213);
nor U7532 (N_7532,N_1850,N_607);
and U7533 (N_7533,N_2224,N_3725);
nand U7534 (N_7534,N_4775,N_2395);
or U7535 (N_7535,N_3338,N_850);
or U7536 (N_7536,N_4664,N_1637);
nor U7537 (N_7537,N_368,N_4762);
nand U7538 (N_7538,N_1426,N_1984);
and U7539 (N_7539,N_1399,N_1950);
or U7540 (N_7540,N_4846,N_4758);
and U7541 (N_7541,N_3544,N_2194);
and U7542 (N_7542,N_4212,N_838);
or U7543 (N_7543,N_2206,N_861);
or U7544 (N_7544,N_3115,N_3615);
nor U7545 (N_7545,N_3830,N_4235);
and U7546 (N_7546,N_2010,N_4945);
nand U7547 (N_7547,N_564,N_3919);
or U7548 (N_7548,N_4699,N_3394);
or U7549 (N_7549,N_1174,N_1634);
nor U7550 (N_7550,N_3994,N_3348);
or U7551 (N_7551,N_3639,N_242);
or U7552 (N_7552,N_2394,N_3943);
and U7553 (N_7553,N_2488,N_1731);
nor U7554 (N_7554,N_2141,N_4267);
nor U7555 (N_7555,N_4923,N_2326);
nor U7556 (N_7556,N_456,N_3522);
nand U7557 (N_7557,N_4155,N_4720);
and U7558 (N_7558,N_351,N_1541);
nand U7559 (N_7559,N_4786,N_2859);
or U7560 (N_7560,N_2385,N_778);
and U7561 (N_7561,N_1262,N_4077);
nand U7562 (N_7562,N_1470,N_3478);
nor U7563 (N_7563,N_4532,N_3631);
and U7564 (N_7564,N_3266,N_779);
nand U7565 (N_7565,N_2551,N_369);
xor U7566 (N_7566,N_1014,N_3114);
nand U7567 (N_7567,N_2198,N_3874);
nand U7568 (N_7568,N_4655,N_1388);
xnor U7569 (N_7569,N_1079,N_4220);
nand U7570 (N_7570,N_3803,N_1544);
nand U7571 (N_7571,N_1294,N_769);
or U7572 (N_7572,N_873,N_567);
and U7573 (N_7573,N_834,N_2810);
nor U7574 (N_7574,N_2461,N_4032);
and U7575 (N_7575,N_4720,N_3219);
nor U7576 (N_7576,N_3170,N_3771);
nor U7577 (N_7577,N_4671,N_2248);
nor U7578 (N_7578,N_1644,N_4083);
and U7579 (N_7579,N_917,N_1374);
nand U7580 (N_7580,N_4121,N_3688);
and U7581 (N_7581,N_3610,N_3222);
nor U7582 (N_7582,N_3517,N_1806);
or U7583 (N_7583,N_3458,N_3641);
nand U7584 (N_7584,N_1912,N_4374);
and U7585 (N_7585,N_1111,N_2896);
or U7586 (N_7586,N_220,N_2166);
and U7587 (N_7587,N_3169,N_1742);
or U7588 (N_7588,N_2272,N_462);
nand U7589 (N_7589,N_3757,N_4765);
nand U7590 (N_7590,N_3420,N_208);
nor U7591 (N_7591,N_3157,N_3183);
and U7592 (N_7592,N_1695,N_3318);
nor U7593 (N_7593,N_3347,N_1846);
and U7594 (N_7594,N_2099,N_4662);
nor U7595 (N_7595,N_1897,N_434);
and U7596 (N_7596,N_2158,N_1983);
nand U7597 (N_7597,N_1698,N_628);
nand U7598 (N_7598,N_4533,N_1796);
or U7599 (N_7599,N_1710,N_1866);
and U7600 (N_7600,N_3031,N_4782);
nor U7601 (N_7601,N_1478,N_377);
nor U7602 (N_7602,N_440,N_796);
or U7603 (N_7603,N_4343,N_486);
nor U7604 (N_7604,N_2765,N_26);
or U7605 (N_7605,N_949,N_2734);
or U7606 (N_7606,N_2852,N_1998);
nand U7607 (N_7607,N_285,N_4218);
nand U7608 (N_7608,N_2942,N_893);
and U7609 (N_7609,N_4233,N_1571);
nor U7610 (N_7610,N_4703,N_963);
and U7611 (N_7611,N_2886,N_495);
nor U7612 (N_7612,N_2210,N_1420);
and U7613 (N_7613,N_4820,N_3947);
nand U7614 (N_7614,N_4243,N_1066);
or U7615 (N_7615,N_1505,N_1478);
or U7616 (N_7616,N_209,N_926);
and U7617 (N_7617,N_2755,N_841);
or U7618 (N_7618,N_2036,N_1477);
nand U7619 (N_7619,N_1690,N_4898);
nor U7620 (N_7620,N_3745,N_4802);
nor U7621 (N_7621,N_3099,N_3459);
nand U7622 (N_7622,N_385,N_4057);
nor U7623 (N_7623,N_4700,N_2084);
or U7624 (N_7624,N_3978,N_68);
or U7625 (N_7625,N_2967,N_4257);
nor U7626 (N_7626,N_2711,N_1598);
nand U7627 (N_7627,N_2737,N_3052);
and U7628 (N_7628,N_3989,N_3532);
and U7629 (N_7629,N_711,N_2992);
nand U7630 (N_7630,N_3842,N_4176);
nand U7631 (N_7631,N_1907,N_4942);
or U7632 (N_7632,N_2199,N_4210);
or U7633 (N_7633,N_3384,N_3517);
or U7634 (N_7634,N_2480,N_67);
nor U7635 (N_7635,N_4483,N_1264);
nand U7636 (N_7636,N_1878,N_586);
nand U7637 (N_7637,N_2992,N_1036);
nor U7638 (N_7638,N_3773,N_1325);
nand U7639 (N_7639,N_3718,N_4987);
and U7640 (N_7640,N_4813,N_1401);
or U7641 (N_7641,N_2258,N_3942);
or U7642 (N_7642,N_3824,N_1767);
or U7643 (N_7643,N_3746,N_3790);
nand U7644 (N_7644,N_3519,N_4511);
and U7645 (N_7645,N_1570,N_1351);
nand U7646 (N_7646,N_1121,N_1069);
or U7647 (N_7647,N_1357,N_2235);
nor U7648 (N_7648,N_3699,N_3516);
or U7649 (N_7649,N_4219,N_891);
and U7650 (N_7650,N_264,N_1305);
and U7651 (N_7651,N_2181,N_337);
and U7652 (N_7652,N_3218,N_319);
or U7653 (N_7653,N_3986,N_2123);
nor U7654 (N_7654,N_361,N_864);
nand U7655 (N_7655,N_3927,N_3980);
nand U7656 (N_7656,N_3550,N_4684);
or U7657 (N_7657,N_4081,N_1843);
and U7658 (N_7658,N_1992,N_2991);
nand U7659 (N_7659,N_3741,N_902);
nor U7660 (N_7660,N_4730,N_555);
or U7661 (N_7661,N_2477,N_4362);
xor U7662 (N_7662,N_3532,N_3087);
nand U7663 (N_7663,N_1396,N_780);
or U7664 (N_7664,N_4957,N_3302);
nor U7665 (N_7665,N_1434,N_2053);
nand U7666 (N_7666,N_489,N_2177);
or U7667 (N_7667,N_4059,N_2495);
nand U7668 (N_7668,N_2479,N_4788);
or U7669 (N_7669,N_3568,N_4092);
xnor U7670 (N_7670,N_917,N_1792);
nor U7671 (N_7671,N_3873,N_594);
nor U7672 (N_7672,N_4458,N_3668);
or U7673 (N_7673,N_152,N_4826);
or U7674 (N_7674,N_3636,N_488);
and U7675 (N_7675,N_1610,N_2957);
nand U7676 (N_7676,N_3475,N_3439);
nand U7677 (N_7677,N_3136,N_1747);
xnor U7678 (N_7678,N_2432,N_546);
nand U7679 (N_7679,N_3651,N_4723);
or U7680 (N_7680,N_3061,N_2405);
nor U7681 (N_7681,N_4007,N_3824);
and U7682 (N_7682,N_3512,N_1920);
and U7683 (N_7683,N_3758,N_3311);
and U7684 (N_7684,N_1078,N_792);
and U7685 (N_7685,N_2999,N_574);
or U7686 (N_7686,N_1288,N_3653);
or U7687 (N_7687,N_939,N_540);
and U7688 (N_7688,N_3817,N_3791);
or U7689 (N_7689,N_336,N_4920);
or U7690 (N_7690,N_2171,N_2067);
nor U7691 (N_7691,N_2721,N_1251);
or U7692 (N_7692,N_4323,N_2037);
or U7693 (N_7693,N_1459,N_2605);
and U7694 (N_7694,N_795,N_3421);
nor U7695 (N_7695,N_4662,N_3221);
nand U7696 (N_7696,N_1613,N_2112);
and U7697 (N_7697,N_767,N_3700);
or U7698 (N_7698,N_1525,N_1886);
nor U7699 (N_7699,N_3067,N_424);
and U7700 (N_7700,N_1824,N_4707);
xnor U7701 (N_7701,N_3121,N_4688);
and U7702 (N_7702,N_885,N_3865);
nor U7703 (N_7703,N_2112,N_2457);
and U7704 (N_7704,N_1318,N_4340);
or U7705 (N_7705,N_4117,N_2448);
and U7706 (N_7706,N_4125,N_4547);
and U7707 (N_7707,N_2831,N_955);
nand U7708 (N_7708,N_479,N_4904);
and U7709 (N_7709,N_4339,N_1103);
nand U7710 (N_7710,N_1232,N_4419);
and U7711 (N_7711,N_1400,N_3181);
nor U7712 (N_7712,N_1875,N_2502);
and U7713 (N_7713,N_3737,N_926);
or U7714 (N_7714,N_1547,N_3208);
nand U7715 (N_7715,N_4450,N_4207);
nand U7716 (N_7716,N_2865,N_50);
nand U7717 (N_7717,N_2849,N_1917);
or U7718 (N_7718,N_849,N_1144);
nor U7719 (N_7719,N_1753,N_3765);
nor U7720 (N_7720,N_1884,N_4301);
and U7721 (N_7721,N_1155,N_72);
nand U7722 (N_7722,N_3946,N_3382);
or U7723 (N_7723,N_854,N_1671);
or U7724 (N_7724,N_177,N_276);
or U7725 (N_7725,N_2026,N_1307);
nand U7726 (N_7726,N_3901,N_2017);
or U7727 (N_7727,N_4612,N_2405);
nand U7728 (N_7728,N_4817,N_4865);
nand U7729 (N_7729,N_1730,N_1677);
or U7730 (N_7730,N_4623,N_4094);
nand U7731 (N_7731,N_4857,N_1572);
xor U7732 (N_7732,N_1236,N_310);
nor U7733 (N_7733,N_3158,N_4143);
or U7734 (N_7734,N_3543,N_1584);
or U7735 (N_7735,N_3321,N_3638);
nand U7736 (N_7736,N_2604,N_256);
nand U7737 (N_7737,N_4044,N_2700);
and U7738 (N_7738,N_1532,N_2421);
and U7739 (N_7739,N_614,N_3882);
nor U7740 (N_7740,N_3535,N_4946);
and U7741 (N_7741,N_3554,N_2966);
nor U7742 (N_7742,N_4360,N_2825);
nand U7743 (N_7743,N_3630,N_990);
or U7744 (N_7744,N_3483,N_1397);
xor U7745 (N_7745,N_4896,N_1641);
nor U7746 (N_7746,N_2744,N_2518);
or U7747 (N_7747,N_1693,N_3763);
and U7748 (N_7748,N_1404,N_1234);
nand U7749 (N_7749,N_3089,N_2818);
nor U7750 (N_7750,N_4460,N_3425);
or U7751 (N_7751,N_442,N_2912);
nor U7752 (N_7752,N_1665,N_1737);
or U7753 (N_7753,N_3105,N_2748);
nor U7754 (N_7754,N_4862,N_3866);
nand U7755 (N_7755,N_591,N_3223);
nor U7756 (N_7756,N_871,N_1231);
nand U7757 (N_7757,N_3808,N_3134);
nand U7758 (N_7758,N_950,N_3362);
nand U7759 (N_7759,N_4795,N_3967);
or U7760 (N_7760,N_383,N_2342);
and U7761 (N_7761,N_1259,N_3400);
or U7762 (N_7762,N_1078,N_1460);
or U7763 (N_7763,N_2467,N_1789);
or U7764 (N_7764,N_3422,N_1753);
nand U7765 (N_7765,N_1565,N_1762);
and U7766 (N_7766,N_4385,N_1438);
nand U7767 (N_7767,N_302,N_2973);
nand U7768 (N_7768,N_2608,N_1910);
nand U7769 (N_7769,N_3474,N_3089);
nor U7770 (N_7770,N_4341,N_3962);
or U7771 (N_7771,N_216,N_19);
nand U7772 (N_7772,N_4535,N_81);
or U7773 (N_7773,N_3625,N_1218);
or U7774 (N_7774,N_1024,N_2528);
nand U7775 (N_7775,N_462,N_98);
and U7776 (N_7776,N_4456,N_3839);
and U7777 (N_7777,N_3476,N_1848);
or U7778 (N_7778,N_4461,N_3873);
or U7779 (N_7779,N_3199,N_3600);
nor U7780 (N_7780,N_336,N_3325);
or U7781 (N_7781,N_4292,N_1776);
and U7782 (N_7782,N_54,N_4900);
nor U7783 (N_7783,N_2174,N_2886);
nor U7784 (N_7784,N_2984,N_2119);
nor U7785 (N_7785,N_3918,N_3471);
nor U7786 (N_7786,N_1768,N_1007);
nor U7787 (N_7787,N_4358,N_3016);
nor U7788 (N_7788,N_2075,N_1016);
nor U7789 (N_7789,N_2312,N_4685);
and U7790 (N_7790,N_3085,N_2642);
or U7791 (N_7791,N_3759,N_2267);
or U7792 (N_7792,N_3053,N_3690);
nand U7793 (N_7793,N_589,N_3058);
or U7794 (N_7794,N_2726,N_1538);
and U7795 (N_7795,N_3129,N_4041);
nor U7796 (N_7796,N_2811,N_2590);
or U7797 (N_7797,N_4959,N_3278);
nor U7798 (N_7798,N_2516,N_3847);
and U7799 (N_7799,N_2501,N_2735);
nor U7800 (N_7800,N_163,N_3644);
nor U7801 (N_7801,N_1444,N_4700);
nor U7802 (N_7802,N_3630,N_3044);
nand U7803 (N_7803,N_1878,N_716);
and U7804 (N_7804,N_4034,N_4412);
nor U7805 (N_7805,N_1740,N_2970);
and U7806 (N_7806,N_773,N_2800);
and U7807 (N_7807,N_3550,N_286);
or U7808 (N_7808,N_1348,N_1746);
or U7809 (N_7809,N_868,N_3014);
nand U7810 (N_7810,N_3441,N_4386);
and U7811 (N_7811,N_2011,N_1200);
or U7812 (N_7812,N_2382,N_510);
nand U7813 (N_7813,N_3433,N_2142);
and U7814 (N_7814,N_477,N_1614);
or U7815 (N_7815,N_2231,N_3171);
and U7816 (N_7816,N_565,N_3139);
and U7817 (N_7817,N_3059,N_4837);
xor U7818 (N_7818,N_726,N_4226);
nand U7819 (N_7819,N_2766,N_3928);
and U7820 (N_7820,N_4405,N_3494);
nand U7821 (N_7821,N_335,N_4388);
or U7822 (N_7822,N_3,N_1973);
nor U7823 (N_7823,N_2493,N_348);
or U7824 (N_7824,N_4273,N_3121);
or U7825 (N_7825,N_2136,N_4361);
nand U7826 (N_7826,N_4292,N_3606);
nor U7827 (N_7827,N_1621,N_1523);
or U7828 (N_7828,N_387,N_1119);
nor U7829 (N_7829,N_613,N_3119);
and U7830 (N_7830,N_619,N_4773);
nand U7831 (N_7831,N_3660,N_1157);
or U7832 (N_7832,N_3793,N_2829);
and U7833 (N_7833,N_658,N_144);
nand U7834 (N_7834,N_3087,N_1499);
or U7835 (N_7835,N_3668,N_230);
nor U7836 (N_7836,N_1831,N_4720);
or U7837 (N_7837,N_1614,N_2795);
nor U7838 (N_7838,N_779,N_1083);
nand U7839 (N_7839,N_1891,N_2632);
nand U7840 (N_7840,N_1679,N_2502);
and U7841 (N_7841,N_3585,N_3300);
nand U7842 (N_7842,N_538,N_2396);
and U7843 (N_7843,N_3944,N_1105);
nor U7844 (N_7844,N_3712,N_4892);
nand U7845 (N_7845,N_3007,N_879);
nand U7846 (N_7846,N_2928,N_2177);
nand U7847 (N_7847,N_3461,N_4823);
nor U7848 (N_7848,N_3991,N_1694);
and U7849 (N_7849,N_1672,N_3599);
or U7850 (N_7850,N_2894,N_1294);
or U7851 (N_7851,N_1594,N_345);
nand U7852 (N_7852,N_3519,N_520);
nand U7853 (N_7853,N_4236,N_1794);
xnor U7854 (N_7854,N_1773,N_3518);
nand U7855 (N_7855,N_2186,N_3079);
or U7856 (N_7856,N_776,N_4781);
nand U7857 (N_7857,N_799,N_1948);
xnor U7858 (N_7858,N_124,N_2966);
nor U7859 (N_7859,N_1709,N_2588);
or U7860 (N_7860,N_4094,N_2162);
nor U7861 (N_7861,N_3466,N_1687);
and U7862 (N_7862,N_2961,N_1872);
or U7863 (N_7863,N_3115,N_4017);
nand U7864 (N_7864,N_3409,N_1150);
and U7865 (N_7865,N_1836,N_1893);
or U7866 (N_7866,N_78,N_2558);
nor U7867 (N_7867,N_1824,N_2607);
nor U7868 (N_7868,N_3107,N_1497);
and U7869 (N_7869,N_822,N_3459);
nand U7870 (N_7870,N_2398,N_3009);
or U7871 (N_7871,N_2679,N_4329);
nor U7872 (N_7872,N_103,N_3075);
nor U7873 (N_7873,N_3640,N_2176);
and U7874 (N_7874,N_3030,N_1266);
nand U7875 (N_7875,N_3051,N_1722);
and U7876 (N_7876,N_2835,N_3625);
and U7877 (N_7877,N_700,N_3010);
and U7878 (N_7878,N_90,N_626);
and U7879 (N_7879,N_878,N_2277);
nor U7880 (N_7880,N_397,N_3748);
or U7881 (N_7881,N_1129,N_2570);
and U7882 (N_7882,N_2930,N_4325);
nand U7883 (N_7883,N_3257,N_2273);
or U7884 (N_7884,N_1822,N_591);
nand U7885 (N_7885,N_3122,N_2550);
or U7886 (N_7886,N_3881,N_3221);
nor U7887 (N_7887,N_3860,N_2966);
and U7888 (N_7888,N_3370,N_3686);
nand U7889 (N_7889,N_4661,N_3203);
and U7890 (N_7890,N_3416,N_3534);
and U7891 (N_7891,N_3645,N_2068);
nand U7892 (N_7892,N_2278,N_4227);
and U7893 (N_7893,N_1920,N_568);
or U7894 (N_7894,N_831,N_3777);
or U7895 (N_7895,N_3906,N_4491);
nor U7896 (N_7896,N_3997,N_4302);
or U7897 (N_7897,N_774,N_2168);
nand U7898 (N_7898,N_2939,N_2684);
or U7899 (N_7899,N_1337,N_2644);
and U7900 (N_7900,N_419,N_2272);
nand U7901 (N_7901,N_3230,N_2362);
nand U7902 (N_7902,N_4253,N_872);
nor U7903 (N_7903,N_2896,N_3162);
or U7904 (N_7904,N_1056,N_4859);
nand U7905 (N_7905,N_2119,N_3965);
nor U7906 (N_7906,N_3877,N_3237);
or U7907 (N_7907,N_4509,N_307);
nor U7908 (N_7908,N_845,N_3081);
nand U7909 (N_7909,N_398,N_4816);
nor U7910 (N_7910,N_4225,N_4931);
and U7911 (N_7911,N_412,N_2733);
nor U7912 (N_7912,N_519,N_1944);
nor U7913 (N_7913,N_3389,N_4662);
nand U7914 (N_7914,N_4260,N_1018);
and U7915 (N_7915,N_1137,N_4278);
nand U7916 (N_7916,N_229,N_2546);
and U7917 (N_7917,N_2534,N_2479);
nor U7918 (N_7918,N_2652,N_3169);
and U7919 (N_7919,N_4756,N_2984);
nand U7920 (N_7920,N_3450,N_1776);
nor U7921 (N_7921,N_1952,N_2644);
and U7922 (N_7922,N_1320,N_2888);
nor U7923 (N_7923,N_4540,N_2367);
or U7924 (N_7924,N_1630,N_4648);
nor U7925 (N_7925,N_2460,N_3857);
or U7926 (N_7926,N_3354,N_1553);
nor U7927 (N_7927,N_763,N_2581);
nor U7928 (N_7928,N_3415,N_375);
or U7929 (N_7929,N_2285,N_1245);
nor U7930 (N_7930,N_558,N_2036);
or U7931 (N_7931,N_786,N_617);
nor U7932 (N_7932,N_4572,N_2818);
or U7933 (N_7933,N_3149,N_1315);
nor U7934 (N_7934,N_704,N_2117);
nand U7935 (N_7935,N_3817,N_2711);
nand U7936 (N_7936,N_2702,N_732);
nand U7937 (N_7937,N_2560,N_4128);
nor U7938 (N_7938,N_879,N_1974);
or U7939 (N_7939,N_2896,N_3588);
or U7940 (N_7940,N_1673,N_1555);
nor U7941 (N_7941,N_1511,N_1802);
nor U7942 (N_7942,N_3242,N_430);
or U7943 (N_7943,N_1844,N_1068);
or U7944 (N_7944,N_2536,N_2942);
nand U7945 (N_7945,N_4445,N_2285);
and U7946 (N_7946,N_230,N_1716);
nand U7947 (N_7947,N_1582,N_3323);
or U7948 (N_7948,N_1264,N_981);
nor U7949 (N_7949,N_1582,N_190);
nor U7950 (N_7950,N_1679,N_4531);
nor U7951 (N_7951,N_1960,N_3195);
xnor U7952 (N_7952,N_262,N_585);
nand U7953 (N_7953,N_1035,N_4753);
nor U7954 (N_7954,N_4400,N_4539);
and U7955 (N_7955,N_829,N_4633);
nor U7956 (N_7956,N_3630,N_1810);
nand U7957 (N_7957,N_3995,N_1713);
and U7958 (N_7958,N_259,N_2637);
nor U7959 (N_7959,N_4827,N_832);
and U7960 (N_7960,N_2662,N_3796);
nor U7961 (N_7961,N_3843,N_4333);
or U7962 (N_7962,N_2311,N_4771);
and U7963 (N_7963,N_1920,N_2335);
nor U7964 (N_7964,N_3346,N_1250);
and U7965 (N_7965,N_843,N_4186);
nor U7966 (N_7966,N_3215,N_3072);
nand U7967 (N_7967,N_4259,N_4220);
and U7968 (N_7968,N_2115,N_2176);
nor U7969 (N_7969,N_3227,N_3090);
and U7970 (N_7970,N_1586,N_3742);
nand U7971 (N_7971,N_413,N_3164);
nand U7972 (N_7972,N_2387,N_4198);
nor U7973 (N_7973,N_4487,N_421);
nor U7974 (N_7974,N_3254,N_2100);
and U7975 (N_7975,N_2470,N_3843);
or U7976 (N_7976,N_1737,N_2280);
nor U7977 (N_7977,N_3089,N_1235);
and U7978 (N_7978,N_4162,N_4793);
nor U7979 (N_7979,N_2635,N_3599);
or U7980 (N_7980,N_4274,N_2182);
or U7981 (N_7981,N_120,N_276);
or U7982 (N_7982,N_2653,N_1583);
or U7983 (N_7983,N_804,N_2112);
and U7984 (N_7984,N_1779,N_4431);
and U7985 (N_7985,N_3973,N_3308);
nor U7986 (N_7986,N_2135,N_3258);
nor U7987 (N_7987,N_4569,N_2997);
nor U7988 (N_7988,N_4606,N_95);
nor U7989 (N_7989,N_4734,N_3747);
and U7990 (N_7990,N_4333,N_1544);
or U7991 (N_7991,N_4554,N_3747);
and U7992 (N_7992,N_2494,N_1826);
or U7993 (N_7993,N_4810,N_1523);
nand U7994 (N_7994,N_2699,N_4262);
or U7995 (N_7995,N_261,N_4698);
and U7996 (N_7996,N_4890,N_1423);
nor U7997 (N_7997,N_4497,N_170);
or U7998 (N_7998,N_3137,N_1453);
nand U7999 (N_7999,N_4484,N_2044);
and U8000 (N_8000,N_1193,N_4332);
and U8001 (N_8001,N_1718,N_271);
nand U8002 (N_8002,N_1657,N_2288);
and U8003 (N_8003,N_809,N_4905);
nor U8004 (N_8004,N_2607,N_455);
nand U8005 (N_8005,N_639,N_2476);
and U8006 (N_8006,N_116,N_4008);
nor U8007 (N_8007,N_1383,N_4663);
and U8008 (N_8008,N_2781,N_1084);
and U8009 (N_8009,N_2246,N_1647);
and U8010 (N_8010,N_4382,N_277);
nand U8011 (N_8011,N_2262,N_3966);
nor U8012 (N_8012,N_1359,N_336);
nor U8013 (N_8013,N_3581,N_4357);
and U8014 (N_8014,N_2090,N_4363);
nand U8015 (N_8015,N_2519,N_2417);
nor U8016 (N_8016,N_4270,N_1087);
and U8017 (N_8017,N_2201,N_3968);
and U8018 (N_8018,N_135,N_995);
nand U8019 (N_8019,N_2271,N_4436);
nand U8020 (N_8020,N_4719,N_890);
nor U8021 (N_8021,N_1584,N_2062);
or U8022 (N_8022,N_2345,N_4509);
nand U8023 (N_8023,N_2123,N_161);
nand U8024 (N_8024,N_2250,N_3278);
and U8025 (N_8025,N_3266,N_1329);
and U8026 (N_8026,N_2549,N_2274);
nand U8027 (N_8027,N_4294,N_3502);
or U8028 (N_8028,N_357,N_2794);
nand U8029 (N_8029,N_3424,N_3925);
nand U8030 (N_8030,N_4132,N_371);
nand U8031 (N_8031,N_4800,N_4121);
nand U8032 (N_8032,N_3703,N_3726);
nor U8033 (N_8033,N_412,N_863);
or U8034 (N_8034,N_1409,N_3262);
nand U8035 (N_8035,N_4271,N_3470);
and U8036 (N_8036,N_2138,N_4922);
or U8037 (N_8037,N_3302,N_1418);
or U8038 (N_8038,N_2601,N_660);
and U8039 (N_8039,N_2088,N_1647);
nand U8040 (N_8040,N_1860,N_3977);
nor U8041 (N_8041,N_42,N_2523);
and U8042 (N_8042,N_1622,N_2555);
nand U8043 (N_8043,N_4743,N_4629);
or U8044 (N_8044,N_3013,N_3796);
nor U8045 (N_8045,N_2908,N_1660);
nor U8046 (N_8046,N_749,N_114);
and U8047 (N_8047,N_2038,N_589);
nand U8048 (N_8048,N_2110,N_4203);
nor U8049 (N_8049,N_887,N_3077);
nor U8050 (N_8050,N_987,N_1647);
nor U8051 (N_8051,N_4771,N_509);
and U8052 (N_8052,N_2881,N_2110);
or U8053 (N_8053,N_2240,N_809);
or U8054 (N_8054,N_1640,N_2632);
or U8055 (N_8055,N_3226,N_3665);
and U8056 (N_8056,N_917,N_4204);
or U8057 (N_8057,N_4348,N_4613);
nor U8058 (N_8058,N_1522,N_9);
nand U8059 (N_8059,N_418,N_537);
and U8060 (N_8060,N_3521,N_3509);
nand U8061 (N_8061,N_680,N_349);
nand U8062 (N_8062,N_3679,N_4938);
or U8063 (N_8063,N_3733,N_3853);
or U8064 (N_8064,N_1809,N_3425);
and U8065 (N_8065,N_3086,N_3424);
nand U8066 (N_8066,N_836,N_3774);
and U8067 (N_8067,N_994,N_3671);
nand U8068 (N_8068,N_1750,N_4412);
and U8069 (N_8069,N_668,N_56);
or U8070 (N_8070,N_4217,N_4226);
or U8071 (N_8071,N_3091,N_419);
or U8072 (N_8072,N_483,N_4012);
nand U8073 (N_8073,N_4364,N_3467);
or U8074 (N_8074,N_2185,N_653);
or U8075 (N_8075,N_3626,N_297);
nor U8076 (N_8076,N_1174,N_445);
and U8077 (N_8077,N_1675,N_4602);
nand U8078 (N_8078,N_1595,N_214);
nor U8079 (N_8079,N_3946,N_3133);
nand U8080 (N_8080,N_4989,N_4873);
or U8081 (N_8081,N_2578,N_2022);
nand U8082 (N_8082,N_1751,N_2240);
nor U8083 (N_8083,N_4071,N_1728);
or U8084 (N_8084,N_2729,N_2394);
xor U8085 (N_8085,N_4256,N_2311);
nand U8086 (N_8086,N_3409,N_2918);
nand U8087 (N_8087,N_3537,N_1088);
nand U8088 (N_8088,N_1197,N_2920);
or U8089 (N_8089,N_1119,N_4226);
nor U8090 (N_8090,N_4967,N_634);
and U8091 (N_8091,N_3600,N_3);
and U8092 (N_8092,N_2505,N_2150);
and U8093 (N_8093,N_1418,N_1823);
nor U8094 (N_8094,N_1492,N_3418);
and U8095 (N_8095,N_2781,N_680);
or U8096 (N_8096,N_2121,N_4057);
nand U8097 (N_8097,N_4190,N_741);
xor U8098 (N_8098,N_3708,N_4207);
nand U8099 (N_8099,N_1787,N_758);
or U8100 (N_8100,N_3181,N_1145);
or U8101 (N_8101,N_3825,N_1195);
nand U8102 (N_8102,N_3675,N_2815);
or U8103 (N_8103,N_984,N_4775);
or U8104 (N_8104,N_2520,N_1895);
and U8105 (N_8105,N_3728,N_3117);
nand U8106 (N_8106,N_4305,N_3489);
and U8107 (N_8107,N_3782,N_3329);
nor U8108 (N_8108,N_2962,N_1894);
and U8109 (N_8109,N_3666,N_4038);
or U8110 (N_8110,N_3615,N_1648);
nand U8111 (N_8111,N_970,N_1723);
nor U8112 (N_8112,N_1621,N_2810);
nand U8113 (N_8113,N_2664,N_1494);
nor U8114 (N_8114,N_2547,N_1764);
or U8115 (N_8115,N_2985,N_1018);
or U8116 (N_8116,N_3703,N_929);
and U8117 (N_8117,N_2325,N_3888);
nor U8118 (N_8118,N_2798,N_1148);
nand U8119 (N_8119,N_1492,N_3374);
or U8120 (N_8120,N_4535,N_1147);
and U8121 (N_8121,N_2514,N_3360);
and U8122 (N_8122,N_4844,N_891);
or U8123 (N_8123,N_1222,N_1146);
and U8124 (N_8124,N_3218,N_2918);
or U8125 (N_8125,N_2373,N_3398);
nand U8126 (N_8126,N_4501,N_4697);
or U8127 (N_8127,N_544,N_2397);
and U8128 (N_8128,N_2934,N_4880);
and U8129 (N_8129,N_263,N_1606);
nand U8130 (N_8130,N_4209,N_805);
or U8131 (N_8131,N_2718,N_4527);
or U8132 (N_8132,N_2236,N_3659);
nor U8133 (N_8133,N_1480,N_3438);
and U8134 (N_8134,N_3963,N_33);
and U8135 (N_8135,N_2157,N_3368);
and U8136 (N_8136,N_332,N_4730);
nand U8137 (N_8137,N_4522,N_4312);
and U8138 (N_8138,N_954,N_3560);
or U8139 (N_8139,N_1773,N_2586);
nor U8140 (N_8140,N_3747,N_4313);
xor U8141 (N_8141,N_7,N_1871);
nand U8142 (N_8142,N_1158,N_3905);
or U8143 (N_8143,N_4709,N_4351);
nand U8144 (N_8144,N_151,N_3466);
and U8145 (N_8145,N_3787,N_2352);
or U8146 (N_8146,N_3120,N_4405);
and U8147 (N_8147,N_3656,N_3538);
and U8148 (N_8148,N_3743,N_361);
or U8149 (N_8149,N_1907,N_898);
nor U8150 (N_8150,N_524,N_2271);
nand U8151 (N_8151,N_4568,N_961);
and U8152 (N_8152,N_2703,N_1668);
and U8153 (N_8153,N_1665,N_3683);
nand U8154 (N_8154,N_3333,N_3002);
or U8155 (N_8155,N_2609,N_3317);
nand U8156 (N_8156,N_3998,N_3277);
and U8157 (N_8157,N_3424,N_1981);
and U8158 (N_8158,N_3809,N_2907);
and U8159 (N_8159,N_3279,N_4171);
nor U8160 (N_8160,N_2114,N_4996);
nor U8161 (N_8161,N_4501,N_2221);
and U8162 (N_8162,N_3236,N_1687);
or U8163 (N_8163,N_3642,N_4908);
or U8164 (N_8164,N_4064,N_3705);
or U8165 (N_8165,N_3833,N_1432);
or U8166 (N_8166,N_3361,N_2731);
nor U8167 (N_8167,N_4502,N_625);
nand U8168 (N_8168,N_2548,N_4534);
or U8169 (N_8169,N_1874,N_4237);
nand U8170 (N_8170,N_3157,N_3796);
nor U8171 (N_8171,N_747,N_1454);
nand U8172 (N_8172,N_2909,N_2274);
and U8173 (N_8173,N_448,N_1514);
nand U8174 (N_8174,N_2347,N_3328);
nor U8175 (N_8175,N_1600,N_900);
or U8176 (N_8176,N_722,N_835);
nand U8177 (N_8177,N_3736,N_293);
nor U8178 (N_8178,N_1177,N_4381);
nor U8179 (N_8179,N_1931,N_3181);
nand U8180 (N_8180,N_1651,N_4973);
and U8181 (N_8181,N_4772,N_2354);
and U8182 (N_8182,N_2670,N_1908);
nor U8183 (N_8183,N_584,N_4423);
and U8184 (N_8184,N_2945,N_4552);
or U8185 (N_8185,N_299,N_3596);
xnor U8186 (N_8186,N_4700,N_1966);
or U8187 (N_8187,N_3305,N_3187);
xnor U8188 (N_8188,N_1844,N_3313);
nand U8189 (N_8189,N_1512,N_2191);
or U8190 (N_8190,N_2118,N_3473);
nand U8191 (N_8191,N_4773,N_887);
or U8192 (N_8192,N_3665,N_824);
nor U8193 (N_8193,N_4836,N_1897);
or U8194 (N_8194,N_716,N_4498);
nor U8195 (N_8195,N_778,N_2301);
nand U8196 (N_8196,N_166,N_3807);
or U8197 (N_8197,N_1548,N_4296);
or U8198 (N_8198,N_4159,N_327);
and U8199 (N_8199,N_2412,N_1408);
and U8200 (N_8200,N_2388,N_4298);
nand U8201 (N_8201,N_1287,N_3111);
nand U8202 (N_8202,N_380,N_4981);
and U8203 (N_8203,N_4402,N_3534);
and U8204 (N_8204,N_238,N_4802);
or U8205 (N_8205,N_536,N_1814);
nand U8206 (N_8206,N_1549,N_3839);
xor U8207 (N_8207,N_1568,N_3197);
and U8208 (N_8208,N_4106,N_2241);
nor U8209 (N_8209,N_117,N_464);
or U8210 (N_8210,N_2673,N_905);
xor U8211 (N_8211,N_4617,N_1830);
and U8212 (N_8212,N_4288,N_2663);
nor U8213 (N_8213,N_4152,N_2029);
and U8214 (N_8214,N_2961,N_3665);
nor U8215 (N_8215,N_3466,N_272);
nor U8216 (N_8216,N_942,N_4694);
and U8217 (N_8217,N_2622,N_4620);
nor U8218 (N_8218,N_3336,N_3752);
or U8219 (N_8219,N_2918,N_628);
nand U8220 (N_8220,N_689,N_1294);
nand U8221 (N_8221,N_4811,N_3755);
xor U8222 (N_8222,N_1329,N_928);
nor U8223 (N_8223,N_2853,N_3976);
and U8224 (N_8224,N_1027,N_540);
xnor U8225 (N_8225,N_1556,N_1922);
or U8226 (N_8226,N_912,N_3669);
or U8227 (N_8227,N_1879,N_379);
and U8228 (N_8228,N_4931,N_2384);
and U8229 (N_8229,N_2378,N_3011);
and U8230 (N_8230,N_4863,N_3627);
nor U8231 (N_8231,N_745,N_1253);
and U8232 (N_8232,N_4397,N_3034);
nor U8233 (N_8233,N_2215,N_4138);
nor U8234 (N_8234,N_989,N_2480);
nor U8235 (N_8235,N_913,N_1251);
nor U8236 (N_8236,N_1075,N_1327);
and U8237 (N_8237,N_3342,N_1711);
and U8238 (N_8238,N_2510,N_2372);
nor U8239 (N_8239,N_4566,N_3579);
and U8240 (N_8240,N_936,N_3270);
nand U8241 (N_8241,N_4121,N_3167);
or U8242 (N_8242,N_4158,N_4673);
nor U8243 (N_8243,N_1360,N_1116);
and U8244 (N_8244,N_685,N_2527);
nand U8245 (N_8245,N_4378,N_434);
nand U8246 (N_8246,N_1484,N_266);
nand U8247 (N_8247,N_3092,N_1123);
nor U8248 (N_8248,N_2428,N_4378);
or U8249 (N_8249,N_2241,N_3645);
nor U8250 (N_8250,N_664,N_2088);
nor U8251 (N_8251,N_1343,N_4755);
nand U8252 (N_8252,N_2893,N_201);
or U8253 (N_8253,N_376,N_3574);
or U8254 (N_8254,N_3176,N_2351);
and U8255 (N_8255,N_3502,N_2147);
nor U8256 (N_8256,N_3890,N_4032);
and U8257 (N_8257,N_2734,N_4274);
nand U8258 (N_8258,N_4578,N_1827);
nand U8259 (N_8259,N_4661,N_4373);
nand U8260 (N_8260,N_1491,N_3269);
nor U8261 (N_8261,N_3325,N_608);
and U8262 (N_8262,N_174,N_38);
nand U8263 (N_8263,N_863,N_207);
or U8264 (N_8264,N_2371,N_2342);
and U8265 (N_8265,N_235,N_1532);
xor U8266 (N_8266,N_3238,N_2269);
nor U8267 (N_8267,N_1005,N_4922);
and U8268 (N_8268,N_4458,N_2194);
nor U8269 (N_8269,N_3147,N_1023);
and U8270 (N_8270,N_4319,N_707);
or U8271 (N_8271,N_1931,N_2482);
and U8272 (N_8272,N_1303,N_4412);
and U8273 (N_8273,N_3921,N_4803);
nand U8274 (N_8274,N_225,N_3765);
nand U8275 (N_8275,N_3464,N_3174);
or U8276 (N_8276,N_3686,N_2368);
and U8277 (N_8277,N_113,N_3387);
or U8278 (N_8278,N_211,N_2234);
nand U8279 (N_8279,N_774,N_3626);
or U8280 (N_8280,N_109,N_367);
nand U8281 (N_8281,N_1675,N_4469);
and U8282 (N_8282,N_2242,N_4519);
and U8283 (N_8283,N_3786,N_3709);
and U8284 (N_8284,N_4624,N_1347);
nor U8285 (N_8285,N_3075,N_4451);
or U8286 (N_8286,N_4247,N_1764);
nor U8287 (N_8287,N_893,N_2760);
and U8288 (N_8288,N_2590,N_4841);
nand U8289 (N_8289,N_3529,N_3522);
or U8290 (N_8290,N_3830,N_1564);
and U8291 (N_8291,N_2372,N_760);
nor U8292 (N_8292,N_3228,N_2174);
or U8293 (N_8293,N_3430,N_2140);
or U8294 (N_8294,N_2453,N_4548);
nand U8295 (N_8295,N_5,N_4199);
or U8296 (N_8296,N_2937,N_3540);
nand U8297 (N_8297,N_4918,N_47);
nand U8298 (N_8298,N_1514,N_524);
nor U8299 (N_8299,N_1858,N_4789);
or U8300 (N_8300,N_2632,N_3330);
or U8301 (N_8301,N_4458,N_2052);
nand U8302 (N_8302,N_2386,N_3011);
and U8303 (N_8303,N_4647,N_4728);
nand U8304 (N_8304,N_3497,N_3296);
nand U8305 (N_8305,N_4017,N_4161);
or U8306 (N_8306,N_2312,N_1497);
nand U8307 (N_8307,N_748,N_772);
or U8308 (N_8308,N_4612,N_1651);
or U8309 (N_8309,N_678,N_3410);
or U8310 (N_8310,N_3732,N_2470);
nand U8311 (N_8311,N_4864,N_219);
nor U8312 (N_8312,N_2829,N_2051);
or U8313 (N_8313,N_3545,N_2591);
or U8314 (N_8314,N_2810,N_4338);
and U8315 (N_8315,N_2274,N_3243);
and U8316 (N_8316,N_4466,N_4846);
and U8317 (N_8317,N_1745,N_2045);
nor U8318 (N_8318,N_2238,N_376);
or U8319 (N_8319,N_248,N_4586);
nand U8320 (N_8320,N_3741,N_989);
or U8321 (N_8321,N_508,N_3839);
or U8322 (N_8322,N_910,N_3123);
or U8323 (N_8323,N_333,N_942);
or U8324 (N_8324,N_420,N_3254);
or U8325 (N_8325,N_590,N_1439);
or U8326 (N_8326,N_349,N_3422);
nand U8327 (N_8327,N_803,N_457);
nand U8328 (N_8328,N_3777,N_890);
nand U8329 (N_8329,N_2009,N_1446);
nor U8330 (N_8330,N_2131,N_1118);
nand U8331 (N_8331,N_1680,N_3653);
or U8332 (N_8332,N_2253,N_2852);
and U8333 (N_8333,N_4697,N_653);
nand U8334 (N_8334,N_1037,N_3019);
or U8335 (N_8335,N_2028,N_2206);
nand U8336 (N_8336,N_3892,N_2175);
and U8337 (N_8337,N_3602,N_4176);
or U8338 (N_8338,N_311,N_151);
and U8339 (N_8339,N_1691,N_4665);
or U8340 (N_8340,N_816,N_1389);
or U8341 (N_8341,N_1742,N_4471);
and U8342 (N_8342,N_575,N_1730);
nand U8343 (N_8343,N_4640,N_30);
nor U8344 (N_8344,N_145,N_4649);
and U8345 (N_8345,N_1034,N_2827);
and U8346 (N_8346,N_2759,N_2429);
nand U8347 (N_8347,N_539,N_2042);
nor U8348 (N_8348,N_3249,N_379);
and U8349 (N_8349,N_293,N_3036);
nand U8350 (N_8350,N_3850,N_4683);
and U8351 (N_8351,N_4239,N_4985);
nand U8352 (N_8352,N_312,N_1022);
nor U8353 (N_8353,N_590,N_3355);
nand U8354 (N_8354,N_2252,N_1533);
nor U8355 (N_8355,N_4521,N_1506);
and U8356 (N_8356,N_1644,N_1473);
nand U8357 (N_8357,N_4058,N_1470);
nand U8358 (N_8358,N_3598,N_4132);
nor U8359 (N_8359,N_1906,N_4519);
or U8360 (N_8360,N_2805,N_92);
and U8361 (N_8361,N_1170,N_530);
or U8362 (N_8362,N_3698,N_255);
nor U8363 (N_8363,N_543,N_2368);
nand U8364 (N_8364,N_2610,N_2850);
nor U8365 (N_8365,N_4399,N_739);
and U8366 (N_8366,N_4483,N_305);
or U8367 (N_8367,N_698,N_242);
or U8368 (N_8368,N_838,N_4026);
nand U8369 (N_8369,N_1866,N_2650);
and U8370 (N_8370,N_937,N_3078);
and U8371 (N_8371,N_3440,N_2387);
or U8372 (N_8372,N_38,N_848);
and U8373 (N_8373,N_617,N_3453);
nand U8374 (N_8374,N_2572,N_54);
nand U8375 (N_8375,N_3713,N_1649);
or U8376 (N_8376,N_3762,N_3019);
nand U8377 (N_8377,N_896,N_1834);
or U8378 (N_8378,N_4262,N_2349);
and U8379 (N_8379,N_586,N_2991);
or U8380 (N_8380,N_967,N_464);
and U8381 (N_8381,N_1928,N_2750);
or U8382 (N_8382,N_458,N_3691);
nor U8383 (N_8383,N_199,N_4803);
nand U8384 (N_8384,N_2814,N_3402);
nor U8385 (N_8385,N_1999,N_924);
nand U8386 (N_8386,N_4762,N_1830);
or U8387 (N_8387,N_4114,N_2709);
and U8388 (N_8388,N_3603,N_4473);
nand U8389 (N_8389,N_4345,N_3882);
or U8390 (N_8390,N_1779,N_1868);
nor U8391 (N_8391,N_4145,N_1569);
and U8392 (N_8392,N_4577,N_1284);
or U8393 (N_8393,N_4299,N_2470);
and U8394 (N_8394,N_334,N_3608);
and U8395 (N_8395,N_2468,N_128);
and U8396 (N_8396,N_2742,N_3989);
and U8397 (N_8397,N_3759,N_2588);
nor U8398 (N_8398,N_4682,N_2700);
and U8399 (N_8399,N_3726,N_692);
and U8400 (N_8400,N_2972,N_3373);
nor U8401 (N_8401,N_957,N_1080);
nor U8402 (N_8402,N_4966,N_3654);
and U8403 (N_8403,N_639,N_1716);
or U8404 (N_8404,N_1943,N_1985);
or U8405 (N_8405,N_3268,N_4886);
and U8406 (N_8406,N_1586,N_917);
nand U8407 (N_8407,N_4469,N_4996);
or U8408 (N_8408,N_1207,N_4092);
nor U8409 (N_8409,N_2808,N_3042);
nor U8410 (N_8410,N_4436,N_679);
nor U8411 (N_8411,N_3586,N_1389);
nor U8412 (N_8412,N_4822,N_2206);
and U8413 (N_8413,N_2753,N_1349);
or U8414 (N_8414,N_4499,N_1375);
nand U8415 (N_8415,N_3241,N_3326);
nand U8416 (N_8416,N_3964,N_57);
or U8417 (N_8417,N_2055,N_2754);
nand U8418 (N_8418,N_3417,N_2667);
and U8419 (N_8419,N_660,N_4178);
or U8420 (N_8420,N_1273,N_588);
and U8421 (N_8421,N_2817,N_732);
nor U8422 (N_8422,N_4857,N_2918);
nand U8423 (N_8423,N_260,N_779);
and U8424 (N_8424,N_3857,N_465);
nor U8425 (N_8425,N_4352,N_2626);
nand U8426 (N_8426,N_3549,N_4097);
nand U8427 (N_8427,N_1738,N_3063);
and U8428 (N_8428,N_1810,N_2844);
and U8429 (N_8429,N_4600,N_4541);
nor U8430 (N_8430,N_79,N_3015);
nor U8431 (N_8431,N_1701,N_1488);
nor U8432 (N_8432,N_4101,N_4775);
or U8433 (N_8433,N_3296,N_3985);
nand U8434 (N_8434,N_1247,N_2644);
nand U8435 (N_8435,N_3146,N_133);
nand U8436 (N_8436,N_3013,N_3670);
and U8437 (N_8437,N_2699,N_4748);
nand U8438 (N_8438,N_412,N_3350);
and U8439 (N_8439,N_2587,N_1702);
nor U8440 (N_8440,N_1807,N_131);
nor U8441 (N_8441,N_1064,N_2287);
or U8442 (N_8442,N_79,N_2320);
nand U8443 (N_8443,N_2283,N_319);
or U8444 (N_8444,N_2874,N_1033);
and U8445 (N_8445,N_4809,N_3536);
nand U8446 (N_8446,N_1988,N_1854);
and U8447 (N_8447,N_738,N_4661);
or U8448 (N_8448,N_3177,N_1220);
nand U8449 (N_8449,N_610,N_4498);
nand U8450 (N_8450,N_2415,N_1139);
nand U8451 (N_8451,N_3541,N_3060);
or U8452 (N_8452,N_3798,N_3702);
nor U8453 (N_8453,N_3925,N_373);
nand U8454 (N_8454,N_757,N_1672);
and U8455 (N_8455,N_3177,N_529);
or U8456 (N_8456,N_1952,N_4199);
and U8457 (N_8457,N_695,N_3049);
and U8458 (N_8458,N_1219,N_2295);
nor U8459 (N_8459,N_2619,N_3431);
or U8460 (N_8460,N_2311,N_3309);
and U8461 (N_8461,N_4753,N_4486);
nor U8462 (N_8462,N_4570,N_3838);
nand U8463 (N_8463,N_1729,N_893);
or U8464 (N_8464,N_2479,N_1002);
or U8465 (N_8465,N_4593,N_4878);
and U8466 (N_8466,N_1238,N_1707);
xor U8467 (N_8467,N_1872,N_2142);
nand U8468 (N_8468,N_172,N_1399);
nor U8469 (N_8469,N_1569,N_3667);
nand U8470 (N_8470,N_4997,N_2352);
nand U8471 (N_8471,N_3169,N_4351);
or U8472 (N_8472,N_3438,N_3683);
or U8473 (N_8473,N_4236,N_124);
nor U8474 (N_8474,N_404,N_4517);
xnor U8475 (N_8475,N_3799,N_137);
or U8476 (N_8476,N_2278,N_2188);
or U8477 (N_8477,N_3204,N_4368);
xor U8478 (N_8478,N_2521,N_4118);
nand U8479 (N_8479,N_2084,N_3147);
nand U8480 (N_8480,N_79,N_2553);
or U8481 (N_8481,N_190,N_2492);
and U8482 (N_8482,N_1999,N_4304);
nand U8483 (N_8483,N_1951,N_4710);
and U8484 (N_8484,N_2446,N_2042);
or U8485 (N_8485,N_3028,N_3917);
nand U8486 (N_8486,N_185,N_542);
nor U8487 (N_8487,N_3059,N_787);
nor U8488 (N_8488,N_4017,N_1818);
or U8489 (N_8489,N_1753,N_3606);
nand U8490 (N_8490,N_594,N_3304);
and U8491 (N_8491,N_358,N_420);
and U8492 (N_8492,N_1410,N_1447);
and U8493 (N_8493,N_4882,N_3400);
and U8494 (N_8494,N_4759,N_3869);
nand U8495 (N_8495,N_1005,N_1625);
nand U8496 (N_8496,N_2461,N_1632);
nor U8497 (N_8497,N_3363,N_2470);
and U8498 (N_8498,N_4858,N_4392);
nor U8499 (N_8499,N_2103,N_4549);
and U8500 (N_8500,N_3594,N_3223);
nand U8501 (N_8501,N_1719,N_2269);
and U8502 (N_8502,N_4736,N_2961);
nand U8503 (N_8503,N_3272,N_438);
nand U8504 (N_8504,N_2973,N_4569);
nor U8505 (N_8505,N_4212,N_3186);
nor U8506 (N_8506,N_3072,N_1898);
nand U8507 (N_8507,N_3019,N_139);
nand U8508 (N_8508,N_3437,N_2006);
nand U8509 (N_8509,N_3735,N_2784);
nand U8510 (N_8510,N_3733,N_3384);
or U8511 (N_8511,N_3085,N_4631);
nand U8512 (N_8512,N_294,N_1097);
and U8513 (N_8513,N_3225,N_3744);
nor U8514 (N_8514,N_3539,N_2769);
and U8515 (N_8515,N_3574,N_1600);
nor U8516 (N_8516,N_2048,N_2516);
or U8517 (N_8517,N_787,N_4879);
nand U8518 (N_8518,N_4206,N_3790);
and U8519 (N_8519,N_2991,N_505);
or U8520 (N_8520,N_4265,N_409);
or U8521 (N_8521,N_1058,N_1666);
nor U8522 (N_8522,N_1834,N_3014);
or U8523 (N_8523,N_2153,N_748);
nor U8524 (N_8524,N_3349,N_517);
nor U8525 (N_8525,N_2253,N_1154);
or U8526 (N_8526,N_4015,N_1032);
and U8527 (N_8527,N_3404,N_4822);
and U8528 (N_8528,N_3487,N_1004);
and U8529 (N_8529,N_1408,N_4403);
or U8530 (N_8530,N_4227,N_1035);
or U8531 (N_8531,N_2339,N_668);
nand U8532 (N_8532,N_3349,N_2912);
or U8533 (N_8533,N_330,N_173);
nor U8534 (N_8534,N_4627,N_4252);
nand U8535 (N_8535,N_2045,N_4368);
nor U8536 (N_8536,N_672,N_2770);
nor U8537 (N_8537,N_4100,N_196);
nor U8538 (N_8538,N_922,N_3141);
nor U8539 (N_8539,N_4240,N_1265);
and U8540 (N_8540,N_4069,N_4816);
nor U8541 (N_8541,N_679,N_1108);
or U8542 (N_8542,N_567,N_3617);
or U8543 (N_8543,N_704,N_3048);
or U8544 (N_8544,N_1544,N_4180);
or U8545 (N_8545,N_1752,N_3013);
nor U8546 (N_8546,N_3099,N_829);
nand U8547 (N_8547,N_1936,N_2945);
or U8548 (N_8548,N_2347,N_2216);
and U8549 (N_8549,N_316,N_2928);
nor U8550 (N_8550,N_2308,N_4068);
nand U8551 (N_8551,N_3332,N_2104);
or U8552 (N_8552,N_3938,N_3841);
or U8553 (N_8553,N_1787,N_3108);
nand U8554 (N_8554,N_236,N_2054);
or U8555 (N_8555,N_3328,N_2641);
or U8556 (N_8556,N_1901,N_4120);
or U8557 (N_8557,N_608,N_4749);
or U8558 (N_8558,N_1146,N_2097);
or U8559 (N_8559,N_764,N_438);
nor U8560 (N_8560,N_4170,N_4951);
or U8561 (N_8561,N_1818,N_2187);
xor U8562 (N_8562,N_2548,N_3507);
nor U8563 (N_8563,N_1418,N_14);
nand U8564 (N_8564,N_2170,N_3563);
and U8565 (N_8565,N_2817,N_1997);
nand U8566 (N_8566,N_4626,N_3451);
nor U8567 (N_8567,N_948,N_4955);
and U8568 (N_8568,N_2171,N_2086);
or U8569 (N_8569,N_2756,N_4402);
nor U8570 (N_8570,N_1451,N_1907);
or U8571 (N_8571,N_4309,N_96);
nand U8572 (N_8572,N_4838,N_2775);
and U8573 (N_8573,N_3644,N_4721);
nor U8574 (N_8574,N_2767,N_3197);
or U8575 (N_8575,N_939,N_942);
and U8576 (N_8576,N_4011,N_4880);
nand U8577 (N_8577,N_384,N_1940);
nand U8578 (N_8578,N_3138,N_4562);
or U8579 (N_8579,N_524,N_101);
nor U8580 (N_8580,N_4295,N_3422);
or U8581 (N_8581,N_3580,N_565);
nor U8582 (N_8582,N_436,N_2864);
nor U8583 (N_8583,N_3097,N_4819);
nand U8584 (N_8584,N_3138,N_1720);
or U8585 (N_8585,N_2847,N_20);
and U8586 (N_8586,N_4943,N_4891);
and U8587 (N_8587,N_351,N_1762);
nor U8588 (N_8588,N_3068,N_2585);
nand U8589 (N_8589,N_3131,N_117);
and U8590 (N_8590,N_294,N_2906);
and U8591 (N_8591,N_376,N_1928);
nand U8592 (N_8592,N_138,N_55);
nand U8593 (N_8593,N_2528,N_3723);
or U8594 (N_8594,N_2648,N_3858);
nor U8595 (N_8595,N_3561,N_2442);
and U8596 (N_8596,N_21,N_4811);
or U8597 (N_8597,N_3078,N_886);
nor U8598 (N_8598,N_1895,N_4033);
nand U8599 (N_8599,N_1614,N_146);
or U8600 (N_8600,N_2566,N_2372);
and U8601 (N_8601,N_4578,N_1603);
and U8602 (N_8602,N_1372,N_2133);
and U8603 (N_8603,N_1643,N_1324);
nand U8604 (N_8604,N_166,N_2942);
or U8605 (N_8605,N_91,N_3535);
nand U8606 (N_8606,N_438,N_3887);
nor U8607 (N_8607,N_3853,N_770);
and U8608 (N_8608,N_3513,N_4426);
nor U8609 (N_8609,N_103,N_3047);
nand U8610 (N_8610,N_4667,N_323);
nor U8611 (N_8611,N_3704,N_4582);
nor U8612 (N_8612,N_446,N_4751);
nor U8613 (N_8613,N_583,N_4835);
nor U8614 (N_8614,N_602,N_4555);
or U8615 (N_8615,N_4079,N_1888);
nor U8616 (N_8616,N_421,N_2049);
nor U8617 (N_8617,N_1515,N_4891);
or U8618 (N_8618,N_1125,N_156);
nor U8619 (N_8619,N_2418,N_4188);
or U8620 (N_8620,N_2400,N_2865);
nand U8621 (N_8621,N_1141,N_1185);
nand U8622 (N_8622,N_2334,N_1543);
nor U8623 (N_8623,N_1507,N_2201);
nor U8624 (N_8624,N_168,N_3569);
and U8625 (N_8625,N_3232,N_4378);
nand U8626 (N_8626,N_3620,N_1372);
nand U8627 (N_8627,N_2587,N_4896);
or U8628 (N_8628,N_1609,N_1132);
and U8629 (N_8629,N_689,N_449);
and U8630 (N_8630,N_1632,N_2950);
nand U8631 (N_8631,N_2686,N_3618);
nand U8632 (N_8632,N_3327,N_3321);
xnor U8633 (N_8633,N_1583,N_3107);
nand U8634 (N_8634,N_4576,N_3405);
and U8635 (N_8635,N_3946,N_3810);
xor U8636 (N_8636,N_2904,N_2442);
or U8637 (N_8637,N_34,N_2297);
nand U8638 (N_8638,N_4552,N_3385);
or U8639 (N_8639,N_3804,N_3925);
or U8640 (N_8640,N_2280,N_4355);
or U8641 (N_8641,N_2602,N_1982);
or U8642 (N_8642,N_1478,N_2529);
nand U8643 (N_8643,N_1820,N_575);
nor U8644 (N_8644,N_3470,N_4895);
or U8645 (N_8645,N_628,N_2795);
or U8646 (N_8646,N_2313,N_4079);
nor U8647 (N_8647,N_2070,N_4221);
nand U8648 (N_8648,N_1630,N_4612);
nand U8649 (N_8649,N_3310,N_236);
nor U8650 (N_8650,N_76,N_1765);
nand U8651 (N_8651,N_1752,N_2206);
or U8652 (N_8652,N_43,N_1381);
nand U8653 (N_8653,N_4401,N_2049);
nand U8654 (N_8654,N_3827,N_3177);
and U8655 (N_8655,N_1501,N_4253);
nand U8656 (N_8656,N_4990,N_3565);
nor U8657 (N_8657,N_1721,N_233);
nor U8658 (N_8658,N_2051,N_1340);
and U8659 (N_8659,N_2063,N_420);
nor U8660 (N_8660,N_2575,N_2612);
nor U8661 (N_8661,N_4190,N_4202);
nand U8662 (N_8662,N_2117,N_3790);
nor U8663 (N_8663,N_345,N_3479);
nand U8664 (N_8664,N_2385,N_2200);
or U8665 (N_8665,N_2788,N_2272);
or U8666 (N_8666,N_2221,N_3809);
nand U8667 (N_8667,N_1106,N_445);
and U8668 (N_8668,N_490,N_1634);
nor U8669 (N_8669,N_3520,N_1172);
or U8670 (N_8670,N_2838,N_3845);
and U8671 (N_8671,N_4530,N_167);
and U8672 (N_8672,N_3783,N_1246);
nand U8673 (N_8673,N_4251,N_293);
nand U8674 (N_8674,N_2439,N_1695);
nor U8675 (N_8675,N_1785,N_1739);
nand U8676 (N_8676,N_288,N_4330);
and U8677 (N_8677,N_2836,N_3776);
and U8678 (N_8678,N_3413,N_2095);
or U8679 (N_8679,N_2157,N_2006);
or U8680 (N_8680,N_892,N_2747);
nor U8681 (N_8681,N_2580,N_4911);
nand U8682 (N_8682,N_1325,N_3347);
nor U8683 (N_8683,N_3623,N_2745);
or U8684 (N_8684,N_3655,N_89);
nor U8685 (N_8685,N_1467,N_1555);
and U8686 (N_8686,N_379,N_4730);
nor U8687 (N_8687,N_2061,N_2308);
or U8688 (N_8688,N_1933,N_1875);
and U8689 (N_8689,N_2138,N_3146);
nand U8690 (N_8690,N_1941,N_585);
and U8691 (N_8691,N_21,N_206);
and U8692 (N_8692,N_3652,N_530);
or U8693 (N_8693,N_3269,N_370);
and U8694 (N_8694,N_217,N_4718);
or U8695 (N_8695,N_4258,N_525);
nand U8696 (N_8696,N_4873,N_2657);
or U8697 (N_8697,N_1935,N_541);
nor U8698 (N_8698,N_3245,N_4555);
nor U8699 (N_8699,N_3814,N_2951);
and U8700 (N_8700,N_530,N_370);
nor U8701 (N_8701,N_2408,N_1238);
nor U8702 (N_8702,N_4732,N_4996);
or U8703 (N_8703,N_1456,N_3691);
nor U8704 (N_8704,N_2819,N_2935);
or U8705 (N_8705,N_1463,N_2683);
and U8706 (N_8706,N_1749,N_4352);
and U8707 (N_8707,N_346,N_2708);
nand U8708 (N_8708,N_1109,N_722);
and U8709 (N_8709,N_2573,N_3455);
nor U8710 (N_8710,N_869,N_4925);
or U8711 (N_8711,N_507,N_3891);
and U8712 (N_8712,N_4771,N_4554);
or U8713 (N_8713,N_2045,N_3306);
nand U8714 (N_8714,N_3453,N_2055);
nor U8715 (N_8715,N_707,N_3912);
and U8716 (N_8716,N_941,N_1782);
or U8717 (N_8717,N_2751,N_1722);
nor U8718 (N_8718,N_4395,N_2581);
or U8719 (N_8719,N_3336,N_3378);
or U8720 (N_8720,N_362,N_3961);
nand U8721 (N_8721,N_2330,N_4656);
and U8722 (N_8722,N_4041,N_361);
or U8723 (N_8723,N_4142,N_4181);
or U8724 (N_8724,N_2848,N_2882);
nor U8725 (N_8725,N_1603,N_3484);
nand U8726 (N_8726,N_3557,N_2073);
or U8727 (N_8727,N_714,N_1173);
nor U8728 (N_8728,N_37,N_3684);
and U8729 (N_8729,N_1164,N_202);
and U8730 (N_8730,N_3013,N_2655);
nand U8731 (N_8731,N_2623,N_4647);
and U8732 (N_8732,N_3371,N_758);
nor U8733 (N_8733,N_2158,N_873);
nor U8734 (N_8734,N_4118,N_2756);
nor U8735 (N_8735,N_1582,N_158);
nor U8736 (N_8736,N_4344,N_4521);
nor U8737 (N_8737,N_2701,N_4680);
and U8738 (N_8738,N_2419,N_34);
and U8739 (N_8739,N_3459,N_1700);
or U8740 (N_8740,N_4979,N_590);
nor U8741 (N_8741,N_2670,N_1636);
or U8742 (N_8742,N_3295,N_144);
and U8743 (N_8743,N_4950,N_483);
and U8744 (N_8744,N_2404,N_3835);
nor U8745 (N_8745,N_2909,N_928);
nand U8746 (N_8746,N_3709,N_3000);
and U8747 (N_8747,N_2620,N_3620);
or U8748 (N_8748,N_3896,N_4459);
or U8749 (N_8749,N_3535,N_2030);
or U8750 (N_8750,N_4434,N_4967);
nor U8751 (N_8751,N_511,N_4657);
nor U8752 (N_8752,N_4099,N_4386);
or U8753 (N_8753,N_2395,N_1850);
and U8754 (N_8754,N_3299,N_4329);
nand U8755 (N_8755,N_4051,N_1951);
nor U8756 (N_8756,N_2862,N_1550);
nand U8757 (N_8757,N_4789,N_2867);
or U8758 (N_8758,N_3861,N_1998);
or U8759 (N_8759,N_3365,N_2341);
nor U8760 (N_8760,N_4129,N_998);
or U8761 (N_8761,N_4235,N_2232);
nor U8762 (N_8762,N_3432,N_841);
nand U8763 (N_8763,N_4313,N_4010);
and U8764 (N_8764,N_2571,N_1545);
and U8765 (N_8765,N_2938,N_2596);
nand U8766 (N_8766,N_4696,N_4605);
or U8767 (N_8767,N_45,N_2575);
or U8768 (N_8768,N_714,N_4919);
and U8769 (N_8769,N_3359,N_3161);
and U8770 (N_8770,N_2276,N_4421);
and U8771 (N_8771,N_2267,N_2835);
nor U8772 (N_8772,N_3847,N_4834);
or U8773 (N_8773,N_4891,N_3325);
and U8774 (N_8774,N_3042,N_3026);
or U8775 (N_8775,N_4966,N_4608);
or U8776 (N_8776,N_2467,N_1026);
or U8777 (N_8777,N_2366,N_4923);
or U8778 (N_8778,N_2718,N_4386);
and U8779 (N_8779,N_2038,N_3185);
and U8780 (N_8780,N_2416,N_910);
and U8781 (N_8781,N_3566,N_2402);
or U8782 (N_8782,N_4664,N_1923);
nor U8783 (N_8783,N_434,N_839);
or U8784 (N_8784,N_341,N_406);
nand U8785 (N_8785,N_3230,N_3875);
nand U8786 (N_8786,N_4165,N_3256);
nand U8787 (N_8787,N_815,N_580);
and U8788 (N_8788,N_491,N_3787);
nand U8789 (N_8789,N_1533,N_2075);
nand U8790 (N_8790,N_1668,N_670);
and U8791 (N_8791,N_644,N_2304);
nand U8792 (N_8792,N_2374,N_3327);
and U8793 (N_8793,N_3607,N_462);
nand U8794 (N_8794,N_848,N_1395);
or U8795 (N_8795,N_2165,N_3670);
and U8796 (N_8796,N_3112,N_3214);
nor U8797 (N_8797,N_311,N_2340);
nor U8798 (N_8798,N_2574,N_2456);
and U8799 (N_8799,N_637,N_3569);
nor U8800 (N_8800,N_1259,N_4211);
nor U8801 (N_8801,N_2277,N_3792);
and U8802 (N_8802,N_4437,N_295);
nand U8803 (N_8803,N_1689,N_194);
nand U8804 (N_8804,N_4815,N_3256);
and U8805 (N_8805,N_2578,N_2967);
or U8806 (N_8806,N_4905,N_4880);
and U8807 (N_8807,N_2488,N_871);
or U8808 (N_8808,N_2708,N_1917);
and U8809 (N_8809,N_821,N_1059);
nand U8810 (N_8810,N_3582,N_253);
and U8811 (N_8811,N_3926,N_3606);
nand U8812 (N_8812,N_3724,N_4960);
nor U8813 (N_8813,N_330,N_3892);
nand U8814 (N_8814,N_2638,N_1579);
nand U8815 (N_8815,N_500,N_2022);
or U8816 (N_8816,N_1730,N_907);
and U8817 (N_8817,N_3797,N_2737);
nor U8818 (N_8818,N_2475,N_2664);
nor U8819 (N_8819,N_2540,N_402);
and U8820 (N_8820,N_4730,N_596);
nor U8821 (N_8821,N_516,N_3528);
and U8822 (N_8822,N_1771,N_4468);
and U8823 (N_8823,N_4215,N_3798);
and U8824 (N_8824,N_1032,N_3659);
or U8825 (N_8825,N_2828,N_2301);
nor U8826 (N_8826,N_689,N_3594);
nor U8827 (N_8827,N_3318,N_2551);
or U8828 (N_8828,N_2706,N_2564);
or U8829 (N_8829,N_4160,N_1325);
nor U8830 (N_8830,N_4367,N_877);
or U8831 (N_8831,N_254,N_2306);
or U8832 (N_8832,N_2861,N_3378);
nor U8833 (N_8833,N_442,N_2532);
nor U8834 (N_8834,N_4357,N_3184);
nor U8835 (N_8835,N_2266,N_420);
nor U8836 (N_8836,N_1799,N_2275);
xor U8837 (N_8837,N_1340,N_1258);
nand U8838 (N_8838,N_652,N_2078);
nand U8839 (N_8839,N_1618,N_3246);
and U8840 (N_8840,N_2667,N_2108);
nand U8841 (N_8841,N_2434,N_4433);
or U8842 (N_8842,N_2428,N_2626);
or U8843 (N_8843,N_1774,N_2823);
or U8844 (N_8844,N_3977,N_1116);
nor U8845 (N_8845,N_3882,N_2339);
nand U8846 (N_8846,N_1380,N_3826);
nand U8847 (N_8847,N_502,N_3112);
or U8848 (N_8848,N_2093,N_4798);
nor U8849 (N_8849,N_332,N_3167);
nand U8850 (N_8850,N_1591,N_612);
or U8851 (N_8851,N_3943,N_3576);
nand U8852 (N_8852,N_2706,N_216);
or U8853 (N_8853,N_604,N_4695);
nor U8854 (N_8854,N_1564,N_4185);
or U8855 (N_8855,N_4935,N_364);
and U8856 (N_8856,N_439,N_2024);
or U8857 (N_8857,N_1550,N_4292);
or U8858 (N_8858,N_4752,N_4542);
or U8859 (N_8859,N_2489,N_2418);
and U8860 (N_8860,N_889,N_1325);
nor U8861 (N_8861,N_3081,N_4743);
or U8862 (N_8862,N_4093,N_186);
and U8863 (N_8863,N_260,N_2125);
nand U8864 (N_8864,N_4569,N_1360);
or U8865 (N_8865,N_3830,N_696);
or U8866 (N_8866,N_1182,N_3612);
nand U8867 (N_8867,N_1869,N_4419);
nor U8868 (N_8868,N_326,N_756);
nor U8869 (N_8869,N_1182,N_2290);
and U8870 (N_8870,N_3647,N_286);
nand U8871 (N_8871,N_3688,N_4445);
nor U8872 (N_8872,N_4456,N_2065);
or U8873 (N_8873,N_4149,N_2830);
nand U8874 (N_8874,N_1772,N_376);
nor U8875 (N_8875,N_3094,N_4921);
nor U8876 (N_8876,N_4105,N_4414);
nand U8877 (N_8877,N_805,N_2112);
nand U8878 (N_8878,N_1998,N_4049);
and U8879 (N_8879,N_1274,N_1158);
nand U8880 (N_8880,N_1204,N_3320);
or U8881 (N_8881,N_4408,N_2364);
or U8882 (N_8882,N_4864,N_1934);
nand U8883 (N_8883,N_2552,N_755);
or U8884 (N_8884,N_387,N_1244);
nand U8885 (N_8885,N_2633,N_2175);
nand U8886 (N_8886,N_2652,N_2195);
and U8887 (N_8887,N_1450,N_1283);
and U8888 (N_8888,N_773,N_4998);
nand U8889 (N_8889,N_276,N_1477);
nand U8890 (N_8890,N_2758,N_1598);
or U8891 (N_8891,N_2473,N_1752);
nor U8892 (N_8892,N_24,N_725);
nand U8893 (N_8893,N_295,N_4652);
or U8894 (N_8894,N_206,N_1182);
nor U8895 (N_8895,N_1478,N_2147);
nand U8896 (N_8896,N_3280,N_3832);
nand U8897 (N_8897,N_1815,N_4286);
nor U8898 (N_8898,N_3579,N_3702);
and U8899 (N_8899,N_4784,N_1020);
nor U8900 (N_8900,N_4442,N_2175);
and U8901 (N_8901,N_3519,N_360);
or U8902 (N_8902,N_769,N_754);
and U8903 (N_8903,N_4228,N_2566);
nor U8904 (N_8904,N_2149,N_2463);
or U8905 (N_8905,N_4099,N_1153);
nand U8906 (N_8906,N_3,N_860);
or U8907 (N_8907,N_1315,N_2343);
nor U8908 (N_8908,N_4470,N_4304);
or U8909 (N_8909,N_2584,N_693);
nor U8910 (N_8910,N_872,N_2832);
and U8911 (N_8911,N_327,N_2598);
or U8912 (N_8912,N_4211,N_925);
nor U8913 (N_8913,N_1004,N_1809);
and U8914 (N_8914,N_1532,N_1741);
or U8915 (N_8915,N_3817,N_4123);
nor U8916 (N_8916,N_541,N_4530);
and U8917 (N_8917,N_1199,N_313);
or U8918 (N_8918,N_1722,N_4051);
nor U8919 (N_8919,N_2253,N_1904);
and U8920 (N_8920,N_3274,N_711);
or U8921 (N_8921,N_1028,N_1207);
nand U8922 (N_8922,N_2339,N_663);
nor U8923 (N_8923,N_1884,N_4998);
nand U8924 (N_8924,N_2427,N_4294);
nand U8925 (N_8925,N_3469,N_1317);
nor U8926 (N_8926,N_4095,N_2806);
and U8927 (N_8927,N_1347,N_4115);
nand U8928 (N_8928,N_3390,N_3628);
nand U8929 (N_8929,N_2596,N_3268);
or U8930 (N_8930,N_2182,N_400);
or U8931 (N_8931,N_1746,N_728);
nor U8932 (N_8932,N_1092,N_4402);
or U8933 (N_8933,N_1592,N_4991);
nand U8934 (N_8934,N_4493,N_1460);
nand U8935 (N_8935,N_3730,N_565);
or U8936 (N_8936,N_3618,N_556);
nand U8937 (N_8937,N_740,N_4019);
nand U8938 (N_8938,N_4942,N_2269);
nor U8939 (N_8939,N_949,N_3736);
nor U8940 (N_8940,N_977,N_4271);
nand U8941 (N_8941,N_4569,N_2287);
nor U8942 (N_8942,N_3782,N_4211);
nand U8943 (N_8943,N_3191,N_3691);
and U8944 (N_8944,N_3860,N_4019);
or U8945 (N_8945,N_3741,N_3820);
nor U8946 (N_8946,N_165,N_219);
and U8947 (N_8947,N_2839,N_4572);
and U8948 (N_8948,N_2774,N_3464);
and U8949 (N_8949,N_692,N_3918);
or U8950 (N_8950,N_596,N_61);
or U8951 (N_8951,N_4219,N_3608);
and U8952 (N_8952,N_1998,N_4632);
or U8953 (N_8953,N_277,N_1709);
nor U8954 (N_8954,N_3352,N_2301);
or U8955 (N_8955,N_61,N_2524);
nor U8956 (N_8956,N_2086,N_4305);
and U8957 (N_8957,N_2152,N_812);
nor U8958 (N_8958,N_1854,N_2340);
and U8959 (N_8959,N_4631,N_3650);
and U8960 (N_8960,N_3481,N_3001);
and U8961 (N_8961,N_1060,N_3687);
and U8962 (N_8962,N_4987,N_1023);
nor U8963 (N_8963,N_1674,N_902);
and U8964 (N_8964,N_4806,N_2950);
or U8965 (N_8965,N_4657,N_3442);
or U8966 (N_8966,N_399,N_873);
nor U8967 (N_8967,N_1844,N_238);
and U8968 (N_8968,N_4314,N_982);
nor U8969 (N_8969,N_4188,N_643);
or U8970 (N_8970,N_3765,N_3489);
or U8971 (N_8971,N_3175,N_1301);
nand U8972 (N_8972,N_2597,N_1271);
nand U8973 (N_8973,N_3411,N_1420);
and U8974 (N_8974,N_614,N_3728);
nor U8975 (N_8975,N_1666,N_1268);
nand U8976 (N_8976,N_3501,N_2970);
nand U8977 (N_8977,N_433,N_3308);
nor U8978 (N_8978,N_4984,N_2242);
and U8979 (N_8979,N_1442,N_4749);
nand U8980 (N_8980,N_4407,N_4309);
and U8981 (N_8981,N_1337,N_1881);
nor U8982 (N_8982,N_3519,N_4180);
nand U8983 (N_8983,N_3494,N_3688);
or U8984 (N_8984,N_1441,N_2644);
and U8985 (N_8985,N_3322,N_2366);
or U8986 (N_8986,N_2864,N_2664);
and U8987 (N_8987,N_1772,N_3909);
and U8988 (N_8988,N_3867,N_3017);
or U8989 (N_8989,N_1522,N_3734);
nor U8990 (N_8990,N_670,N_223);
nand U8991 (N_8991,N_1764,N_2322);
nand U8992 (N_8992,N_4281,N_1724);
or U8993 (N_8993,N_2747,N_82);
nand U8994 (N_8994,N_2472,N_514);
nor U8995 (N_8995,N_397,N_2704);
nor U8996 (N_8996,N_2403,N_937);
nor U8997 (N_8997,N_3758,N_4725);
nor U8998 (N_8998,N_3714,N_4079);
or U8999 (N_8999,N_4867,N_359);
or U9000 (N_9000,N_3908,N_3726);
and U9001 (N_9001,N_1963,N_4507);
nand U9002 (N_9002,N_930,N_2550);
nand U9003 (N_9003,N_4992,N_2136);
nand U9004 (N_9004,N_1022,N_1127);
and U9005 (N_9005,N_3382,N_1878);
or U9006 (N_9006,N_444,N_2564);
or U9007 (N_9007,N_4780,N_621);
nand U9008 (N_9008,N_1199,N_3623);
or U9009 (N_9009,N_2375,N_4399);
or U9010 (N_9010,N_4906,N_4693);
and U9011 (N_9011,N_1867,N_1948);
and U9012 (N_9012,N_3407,N_2939);
and U9013 (N_9013,N_3766,N_2561);
nor U9014 (N_9014,N_963,N_887);
and U9015 (N_9015,N_1270,N_742);
and U9016 (N_9016,N_3152,N_2059);
nand U9017 (N_9017,N_1235,N_2189);
nand U9018 (N_9018,N_2225,N_1865);
nand U9019 (N_9019,N_1285,N_2762);
and U9020 (N_9020,N_3349,N_4937);
nand U9021 (N_9021,N_1998,N_4260);
nor U9022 (N_9022,N_3649,N_4621);
nand U9023 (N_9023,N_813,N_1242);
and U9024 (N_9024,N_1093,N_3311);
nand U9025 (N_9025,N_1607,N_4179);
nand U9026 (N_9026,N_4926,N_910);
and U9027 (N_9027,N_2287,N_4760);
and U9028 (N_9028,N_3049,N_77);
xor U9029 (N_9029,N_3682,N_4309);
and U9030 (N_9030,N_2749,N_3516);
nor U9031 (N_9031,N_323,N_807);
and U9032 (N_9032,N_139,N_3386);
nor U9033 (N_9033,N_2703,N_1269);
nand U9034 (N_9034,N_3069,N_2441);
or U9035 (N_9035,N_3412,N_2429);
and U9036 (N_9036,N_2154,N_2056);
nand U9037 (N_9037,N_2230,N_551);
and U9038 (N_9038,N_4650,N_3702);
nand U9039 (N_9039,N_2192,N_1964);
or U9040 (N_9040,N_4961,N_4264);
and U9041 (N_9041,N_933,N_299);
or U9042 (N_9042,N_4680,N_1191);
and U9043 (N_9043,N_1074,N_2459);
nor U9044 (N_9044,N_3724,N_3088);
nand U9045 (N_9045,N_4496,N_601);
nand U9046 (N_9046,N_476,N_949);
and U9047 (N_9047,N_573,N_345);
or U9048 (N_9048,N_2318,N_3696);
nor U9049 (N_9049,N_4012,N_3698);
nor U9050 (N_9050,N_4707,N_117);
or U9051 (N_9051,N_3533,N_441);
or U9052 (N_9052,N_3559,N_70);
nor U9053 (N_9053,N_4709,N_1170);
and U9054 (N_9054,N_4244,N_1893);
nor U9055 (N_9055,N_4615,N_72);
and U9056 (N_9056,N_1372,N_1434);
nand U9057 (N_9057,N_3374,N_1086);
nand U9058 (N_9058,N_2045,N_3311);
or U9059 (N_9059,N_1156,N_3099);
and U9060 (N_9060,N_3338,N_4978);
nor U9061 (N_9061,N_2981,N_1634);
and U9062 (N_9062,N_3740,N_424);
or U9063 (N_9063,N_2074,N_3299);
or U9064 (N_9064,N_1271,N_500);
or U9065 (N_9065,N_2401,N_4992);
nand U9066 (N_9066,N_4231,N_2602);
nor U9067 (N_9067,N_3874,N_1700);
nand U9068 (N_9068,N_767,N_1610);
nand U9069 (N_9069,N_4764,N_3203);
nor U9070 (N_9070,N_1381,N_4753);
or U9071 (N_9071,N_530,N_4520);
and U9072 (N_9072,N_1057,N_324);
nand U9073 (N_9073,N_4023,N_4936);
or U9074 (N_9074,N_635,N_4225);
or U9075 (N_9075,N_3790,N_762);
and U9076 (N_9076,N_2598,N_1647);
nand U9077 (N_9077,N_1360,N_1546);
nand U9078 (N_9078,N_1403,N_585);
nor U9079 (N_9079,N_3702,N_4869);
nand U9080 (N_9080,N_3466,N_3933);
nor U9081 (N_9081,N_107,N_2983);
or U9082 (N_9082,N_3413,N_8);
and U9083 (N_9083,N_1579,N_3985);
and U9084 (N_9084,N_4401,N_452);
and U9085 (N_9085,N_2844,N_2935);
nand U9086 (N_9086,N_975,N_2511);
nor U9087 (N_9087,N_511,N_4797);
nand U9088 (N_9088,N_1931,N_4795);
nor U9089 (N_9089,N_206,N_2171);
nor U9090 (N_9090,N_2495,N_4295);
or U9091 (N_9091,N_3491,N_874);
or U9092 (N_9092,N_572,N_2800);
and U9093 (N_9093,N_193,N_1167);
nor U9094 (N_9094,N_4677,N_4312);
or U9095 (N_9095,N_2429,N_3280);
nand U9096 (N_9096,N_318,N_4784);
nor U9097 (N_9097,N_3656,N_3165);
and U9098 (N_9098,N_1362,N_3412);
nand U9099 (N_9099,N_4626,N_2869);
nand U9100 (N_9100,N_2168,N_4717);
nand U9101 (N_9101,N_3991,N_1220);
nor U9102 (N_9102,N_1060,N_1003);
nand U9103 (N_9103,N_3224,N_4023);
nand U9104 (N_9104,N_4076,N_869);
or U9105 (N_9105,N_497,N_2420);
nand U9106 (N_9106,N_525,N_2349);
nand U9107 (N_9107,N_4694,N_2487);
or U9108 (N_9108,N_291,N_1247);
nand U9109 (N_9109,N_748,N_1790);
nand U9110 (N_9110,N_1736,N_1318);
nor U9111 (N_9111,N_4533,N_1325);
nor U9112 (N_9112,N_2834,N_3510);
and U9113 (N_9113,N_2770,N_1777);
nor U9114 (N_9114,N_1191,N_100);
or U9115 (N_9115,N_2222,N_2794);
or U9116 (N_9116,N_2106,N_4086);
nor U9117 (N_9117,N_4875,N_1769);
and U9118 (N_9118,N_1465,N_2197);
nand U9119 (N_9119,N_524,N_4427);
and U9120 (N_9120,N_1825,N_3381);
nor U9121 (N_9121,N_1194,N_488);
and U9122 (N_9122,N_3304,N_838);
nor U9123 (N_9123,N_3491,N_2785);
and U9124 (N_9124,N_2577,N_3024);
and U9125 (N_9125,N_4943,N_2552);
and U9126 (N_9126,N_858,N_1526);
nor U9127 (N_9127,N_1214,N_1351);
and U9128 (N_9128,N_463,N_1476);
and U9129 (N_9129,N_2072,N_3735);
and U9130 (N_9130,N_3796,N_760);
and U9131 (N_9131,N_3935,N_3443);
nand U9132 (N_9132,N_4104,N_1940);
nand U9133 (N_9133,N_3378,N_27);
nand U9134 (N_9134,N_1559,N_100);
and U9135 (N_9135,N_3529,N_174);
nand U9136 (N_9136,N_1475,N_665);
or U9137 (N_9137,N_1346,N_2108);
nor U9138 (N_9138,N_3704,N_2941);
and U9139 (N_9139,N_1451,N_3581);
or U9140 (N_9140,N_2585,N_319);
nor U9141 (N_9141,N_1367,N_2488);
nor U9142 (N_9142,N_4725,N_571);
or U9143 (N_9143,N_1242,N_2783);
nor U9144 (N_9144,N_3403,N_2986);
or U9145 (N_9145,N_1333,N_2365);
nor U9146 (N_9146,N_4574,N_1678);
and U9147 (N_9147,N_2089,N_311);
nor U9148 (N_9148,N_1989,N_661);
and U9149 (N_9149,N_2247,N_826);
nor U9150 (N_9150,N_2890,N_2487);
nand U9151 (N_9151,N_1618,N_2635);
or U9152 (N_9152,N_1815,N_3566);
and U9153 (N_9153,N_3243,N_3201);
nor U9154 (N_9154,N_2556,N_4435);
and U9155 (N_9155,N_3627,N_586);
nand U9156 (N_9156,N_500,N_2458);
nor U9157 (N_9157,N_824,N_1658);
nand U9158 (N_9158,N_2566,N_4310);
or U9159 (N_9159,N_3516,N_474);
nand U9160 (N_9160,N_2752,N_3031);
nor U9161 (N_9161,N_1214,N_2352);
xnor U9162 (N_9162,N_781,N_4293);
and U9163 (N_9163,N_2446,N_1459);
nand U9164 (N_9164,N_1994,N_127);
and U9165 (N_9165,N_185,N_4228);
nand U9166 (N_9166,N_139,N_449);
and U9167 (N_9167,N_1104,N_1166);
nand U9168 (N_9168,N_3932,N_3724);
nand U9169 (N_9169,N_2478,N_3544);
nor U9170 (N_9170,N_3926,N_4397);
nor U9171 (N_9171,N_2775,N_580);
and U9172 (N_9172,N_2717,N_1754);
nor U9173 (N_9173,N_2503,N_4993);
nor U9174 (N_9174,N_3955,N_1402);
and U9175 (N_9175,N_3333,N_371);
or U9176 (N_9176,N_145,N_1859);
nand U9177 (N_9177,N_1500,N_1339);
nand U9178 (N_9178,N_729,N_1264);
nand U9179 (N_9179,N_364,N_1441);
or U9180 (N_9180,N_4516,N_2089);
nand U9181 (N_9181,N_846,N_517);
nor U9182 (N_9182,N_1032,N_1732);
nand U9183 (N_9183,N_702,N_2059);
or U9184 (N_9184,N_924,N_3900);
or U9185 (N_9185,N_746,N_1570);
nand U9186 (N_9186,N_216,N_1306);
or U9187 (N_9187,N_439,N_3424);
and U9188 (N_9188,N_1727,N_3292);
or U9189 (N_9189,N_3223,N_215);
nand U9190 (N_9190,N_2596,N_1934);
or U9191 (N_9191,N_303,N_3400);
or U9192 (N_9192,N_2199,N_3453);
and U9193 (N_9193,N_4235,N_4679);
or U9194 (N_9194,N_4798,N_4442);
and U9195 (N_9195,N_724,N_717);
and U9196 (N_9196,N_2166,N_3396);
nor U9197 (N_9197,N_1507,N_530);
nand U9198 (N_9198,N_4413,N_1473);
and U9199 (N_9199,N_2897,N_3114);
and U9200 (N_9200,N_3963,N_3148);
or U9201 (N_9201,N_4432,N_2825);
nand U9202 (N_9202,N_1890,N_1717);
nor U9203 (N_9203,N_25,N_2739);
nor U9204 (N_9204,N_2223,N_3159);
and U9205 (N_9205,N_2629,N_772);
nor U9206 (N_9206,N_3656,N_2754);
and U9207 (N_9207,N_2057,N_4224);
or U9208 (N_9208,N_245,N_2586);
nand U9209 (N_9209,N_3197,N_2313);
nand U9210 (N_9210,N_3983,N_692);
nor U9211 (N_9211,N_4037,N_1656);
or U9212 (N_9212,N_2857,N_4260);
nor U9213 (N_9213,N_902,N_245);
or U9214 (N_9214,N_4829,N_2202);
nand U9215 (N_9215,N_2908,N_2179);
nand U9216 (N_9216,N_2401,N_4525);
and U9217 (N_9217,N_3301,N_156);
and U9218 (N_9218,N_1415,N_2644);
nor U9219 (N_9219,N_3710,N_3600);
or U9220 (N_9220,N_782,N_2159);
and U9221 (N_9221,N_2192,N_2964);
or U9222 (N_9222,N_2933,N_3660);
xor U9223 (N_9223,N_707,N_4373);
and U9224 (N_9224,N_1572,N_4521);
or U9225 (N_9225,N_220,N_2787);
or U9226 (N_9226,N_3064,N_3811);
nor U9227 (N_9227,N_4227,N_4169);
or U9228 (N_9228,N_2922,N_4990);
or U9229 (N_9229,N_2598,N_588);
nor U9230 (N_9230,N_1690,N_1013);
or U9231 (N_9231,N_1964,N_871);
and U9232 (N_9232,N_14,N_4705);
and U9233 (N_9233,N_2911,N_11);
or U9234 (N_9234,N_1975,N_930);
or U9235 (N_9235,N_3973,N_3407);
nand U9236 (N_9236,N_3898,N_4577);
or U9237 (N_9237,N_4939,N_3881);
or U9238 (N_9238,N_2474,N_1060);
and U9239 (N_9239,N_3992,N_1395);
and U9240 (N_9240,N_51,N_3103);
nor U9241 (N_9241,N_2464,N_4527);
or U9242 (N_9242,N_1867,N_420);
nand U9243 (N_9243,N_645,N_275);
or U9244 (N_9244,N_3427,N_2786);
and U9245 (N_9245,N_4153,N_3210);
nand U9246 (N_9246,N_3652,N_889);
nor U9247 (N_9247,N_2639,N_62);
or U9248 (N_9248,N_2740,N_2119);
nor U9249 (N_9249,N_3751,N_1587);
nand U9250 (N_9250,N_4623,N_1885);
or U9251 (N_9251,N_2621,N_3600);
nor U9252 (N_9252,N_1991,N_4349);
xor U9253 (N_9253,N_780,N_4196);
nor U9254 (N_9254,N_4537,N_1897);
and U9255 (N_9255,N_2019,N_1507);
and U9256 (N_9256,N_1438,N_3236);
nand U9257 (N_9257,N_1836,N_1918);
and U9258 (N_9258,N_2681,N_2259);
nor U9259 (N_9259,N_566,N_2329);
nor U9260 (N_9260,N_4683,N_4696);
nand U9261 (N_9261,N_14,N_3283);
or U9262 (N_9262,N_2089,N_1227);
nor U9263 (N_9263,N_1563,N_1225);
nor U9264 (N_9264,N_1170,N_3748);
nand U9265 (N_9265,N_1394,N_2912);
nor U9266 (N_9266,N_602,N_4211);
nand U9267 (N_9267,N_3402,N_4060);
and U9268 (N_9268,N_3653,N_1020);
and U9269 (N_9269,N_154,N_1381);
nor U9270 (N_9270,N_3137,N_3273);
nor U9271 (N_9271,N_2462,N_16);
or U9272 (N_9272,N_4846,N_3071);
or U9273 (N_9273,N_440,N_4950);
and U9274 (N_9274,N_2853,N_3451);
xor U9275 (N_9275,N_1329,N_2121);
nand U9276 (N_9276,N_1081,N_2032);
nand U9277 (N_9277,N_1814,N_370);
and U9278 (N_9278,N_237,N_864);
and U9279 (N_9279,N_3473,N_760);
nor U9280 (N_9280,N_4663,N_3956);
and U9281 (N_9281,N_2655,N_4859);
nand U9282 (N_9282,N_82,N_1508);
nor U9283 (N_9283,N_3825,N_1402);
or U9284 (N_9284,N_2082,N_4595);
or U9285 (N_9285,N_529,N_2824);
and U9286 (N_9286,N_3386,N_1182);
nor U9287 (N_9287,N_3615,N_2854);
and U9288 (N_9288,N_1229,N_3111);
or U9289 (N_9289,N_1344,N_1842);
and U9290 (N_9290,N_908,N_2019);
nand U9291 (N_9291,N_4477,N_2494);
nand U9292 (N_9292,N_2957,N_4284);
nand U9293 (N_9293,N_470,N_3671);
nor U9294 (N_9294,N_2414,N_1325);
nor U9295 (N_9295,N_3822,N_2790);
nand U9296 (N_9296,N_1833,N_37);
nor U9297 (N_9297,N_2326,N_846);
and U9298 (N_9298,N_2921,N_4365);
nand U9299 (N_9299,N_4122,N_924);
and U9300 (N_9300,N_13,N_854);
nor U9301 (N_9301,N_3420,N_3518);
and U9302 (N_9302,N_3784,N_520);
or U9303 (N_9303,N_1451,N_3465);
or U9304 (N_9304,N_255,N_4985);
and U9305 (N_9305,N_846,N_3360);
or U9306 (N_9306,N_4729,N_3115);
or U9307 (N_9307,N_1092,N_232);
nand U9308 (N_9308,N_277,N_4672);
and U9309 (N_9309,N_1668,N_2533);
or U9310 (N_9310,N_2582,N_2074);
or U9311 (N_9311,N_1431,N_1736);
nand U9312 (N_9312,N_4373,N_3313);
nand U9313 (N_9313,N_3118,N_4450);
or U9314 (N_9314,N_3304,N_3016);
and U9315 (N_9315,N_2383,N_2463);
nand U9316 (N_9316,N_4413,N_4088);
and U9317 (N_9317,N_3274,N_3969);
nor U9318 (N_9318,N_1927,N_4217);
or U9319 (N_9319,N_2086,N_1696);
and U9320 (N_9320,N_1365,N_4986);
nor U9321 (N_9321,N_3719,N_1789);
nor U9322 (N_9322,N_4243,N_4723);
and U9323 (N_9323,N_2801,N_1201);
nor U9324 (N_9324,N_1047,N_1712);
and U9325 (N_9325,N_2733,N_1510);
and U9326 (N_9326,N_3527,N_44);
or U9327 (N_9327,N_4992,N_839);
nand U9328 (N_9328,N_4363,N_3895);
nand U9329 (N_9329,N_2607,N_703);
and U9330 (N_9330,N_1823,N_3129);
nor U9331 (N_9331,N_2803,N_4762);
nand U9332 (N_9332,N_4884,N_808);
nand U9333 (N_9333,N_4490,N_4599);
nor U9334 (N_9334,N_4843,N_3464);
and U9335 (N_9335,N_3354,N_4991);
nand U9336 (N_9336,N_2637,N_1853);
or U9337 (N_9337,N_1846,N_3812);
or U9338 (N_9338,N_3528,N_1217);
nand U9339 (N_9339,N_310,N_3512);
xor U9340 (N_9340,N_2542,N_2163);
nor U9341 (N_9341,N_1088,N_1755);
nand U9342 (N_9342,N_706,N_3920);
nor U9343 (N_9343,N_3546,N_1887);
and U9344 (N_9344,N_1903,N_2633);
or U9345 (N_9345,N_1579,N_2254);
nor U9346 (N_9346,N_2348,N_3759);
and U9347 (N_9347,N_1542,N_1029);
and U9348 (N_9348,N_4180,N_1222);
or U9349 (N_9349,N_3445,N_4281);
nor U9350 (N_9350,N_3947,N_1447);
or U9351 (N_9351,N_4214,N_2512);
nand U9352 (N_9352,N_3198,N_1854);
or U9353 (N_9353,N_729,N_1957);
or U9354 (N_9354,N_359,N_1918);
or U9355 (N_9355,N_510,N_1988);
or U9356 (N_9356,N_4681,N_4694);
nand U9357 (N_9357,N_611,N_362);
or U9358 (N_9358,N_2799,N_3);
nand U9359 (N_9359,N_3166,N_4151);
nor U9360 (N_9360,N_1604,N_2004);
nor U9361 (N_9361,N_2253,N_3546);
or U9362 (N_9362,N_83,N_3603);
or U9363 (N_9363,N_1273,N_399);
and U9364 (N_9364,N_4345,N_1144);
and U9365 (N_9365,N_4055,N_1118);
nor U9366 (N_9366,N_608,N_3285);
nor U9367 (N_9367,N_1608,N_3348);
nand U9368 (N_9368,N_1255,N_3805);
nor U9369 (N_9369,N_771,N_4217);
or U9370 (N_9370,N_3911,N_1514);
xnor U9371 (N_9371,N_1325,N_881);
nand U9372 (N_9372,N_4309,N_2907);
nand U9373 (N_9373,N_54,N_4559);
nand U9374 (N_9374,N_4840,N_337);
and U9375 (N_9375,N_647,N_172);
and U9376 (N_9376,N_2526,N_4419);
and U9377 (N_9377,N_3196,N_4264);
nand U9378 (N_9378,N_668,N_3492);
nor U9379 (N_9379,N_1101,N_3168);
nand U9380 (N_9380,N_1107,N_3313);
nand U9381 (N_9381,N_1043,N_1241);
nor U9382 (N_9382,N_3048,N_1139);
or U9383 (N_9383,N_3701,N_2757);
and U9384 (N_9384,N_4348,N_3558);
nor U9385 (N_9385,N_2234,N_1810);
or U9386 (N_9386,N_1256,N_4412);
and U9387 (N_9387,N_3116,N_14);
or U9388 (N_9388,N_272,N_4553);
nand U9389 (N_9389,N_3990,N_4826);
and U9390 (N_9390,N_3831,N_4686);
or U9391 (N_9391,N_2004,N_3283);
or U9392 (N_9392,N_4511,N_4028);
and U9393 (N_9393,N_2940,N_4332);
nand U9394 (N_9394,N_949,N_3050);
and U9395 (N_9395,N_4635,N_1192);
or U9396 (N_9396,N_4165,N_2645);
nor U9397 (N_9397,N_4426,N_4140);
and U9398 (N_9398,N_4211,N_2937);
or U9399 (N_9399,N_1643,N_1124);
nand U9400 (N_9400,N_2150,N_14);
nand U9401 (N_9401,N_1094,N_2391);
and U9402 (N_9402,N_2397,N_1697);
nand U9403 (N_9403,N_242,N_499);
and U9404 (N_9404,N_2603,N_4527);
nand U9405 (N_9405,N_4610,N_4059);
nor U9406 (N_9406,N_4344,N_195);
nand U9407 (N_9407,N_2645,N_4872);
or U9408 (N_9408,N_4436,N_3000);
nor U9409 (N_9409,N_2360,N_1824);
and U9410 (N_9410,N_3069,N_761);
nand U9411 (N_9411,N_4456,N_2660);
nor U9412 (N_9412,N_1781,N_2229);
and U9413 (N_9413,N_431,N_3536);
and U9414 (N_9414,N_776,N_2058);
or U9415 (N_9415,N_334,N_580);
nor U9416 (N_9416,N_190,N_2758);
nand U9417 (N_9417,N_4254,N_4451);
and U9418 (N_9418,N_3128,N_1133);
and U9419 (N_9419,N_731,N_4355);
and U9420 (N_9420,N_1907,N_1514);
or U9421 (N_9421,N_3449,N_1459);
and U9422 (N_9422,N_3921,N_997);
or U9423 (N_9423,N_1031,N_501);
and U9424 (N_9424,N_687,N_3881);
nor U9425 (N_9425,N_4500,N_665);
nand U9426 (N_9426,N_2250,N_4899);
or U9427 (N_9427,N_855,N_934);
nand U9428 (N_9428,N_1311,N_1928);
and U9429 (N_9429,N_685,N_645);
or U9430 (N_9430,N_2204,N_2669);
nor U9431 (N_9431,N_2186,N_683);
or U9432 (N_9432,N_309,N_3020);
and U9433 (N_9433,N_2144,N_4009);
and U9434 (N_9434,N_4113,N_2526);
or U9435 (N_9435,N_369,N_4856);
or U9436 (N_9436,N_4639,N_3304);
nor U9437 (N_9437,N_804,N_3651);
nor U9438 (N_9438,N_2610,N_460);
nor U9439 (N_9439,N_795,N_2769);
nor U9440 (N_9440,N_2265,N_1803);
nand U9441 (N_9441,N_3156,N_3030);
nand U9442 (N_9442,N_2618,N_4599);
nor U9443 (N_9443,N_2695,N_2630);
or U9444 (N_9444,N_4891,N_1978);
or U9445 (N_9445,N_1701,N_3175);
or U9446 (N_9446,N_4043,N_1421);
or U9447 (N_9447,N_958,N_2028);
nand U9448 (N_9448,N_4130,N_413);
nand U9449 (N_9449,N_1225,N_3271);
nand U9450 (N_9450,N_4600,N_4726);
and U9451 (N_9451,N_97,N_1815);
and U9452 (N_9452,N_1311,N_4625);
nor U9453 (N_9453,N_329,N_2686);
nand U9454 (N_9454,N_1354,N_4354);
nor U9455 (N_9455,N_3783,N_65);
nor U9456 (N_9456,N_4623,N_4922);
or U9457 (N_9457,N_647,N_897);
and U9458 (N_9458,N_2653,N_4213);
nor U9459 (N_9459,N_3859,N_4533);
nand U9460 (N_9460,N_100,N_857);
and U9461 (N_9461,N_3063,N_2364);
or U9462 (N_9462,N_1816,N_3119);
nand U9463 (N_9463,N_4030,N_2121);
or U9464 (N_9464,N_815,N_4801);
nor U9465 (N_9465,N_4628,N_3802);
or U9466 (N_9466,N_1687,N_4339);
nand U9467 (N_9467,N_1607,N_1810);
or U9468 (N_9468,N_3719,N_2021);
and U9469 (N_9469,N_4203,N_2037);
xor U9470 (N_9470,N_1369,N_2334);
nand U9471 (N_9471,N_3939,N_4008);
nand U9472 (N_9472,N_767,N_4702);
or U9473 (N_9473,N_4494,N_2877);
and U9474 (N_9474,N_3801,N_1213);
or U9475 (N_9475,N_3686,N_176);
or U9476 (N_9476,N_2669,N_4946);
nand U9477 (N_9477,N_2378,N_1877);
nand U9478 (N_9478,N_2716,N_674);
or U9479 (N_9479,N_1742,N_4024);
nor U9480 (N_9480,N_2335,N_856);
nand U9481 (N_9481,N_4720,N_3846);
or U9482 (N_9482,N_3904,N_52);
or U9483 (N_9483,N_1117,N_1597);
nor U9484 (N_9484,N_1367,N_4803);
or U9485 (N_9485,N_2543,N_3994);
nor U9486 (N_9486,N_3106,N_3800);
nor U9487 (N_9487,N_4991,N_527);
nand U9488 (N_9488,N_1015,N_2169);
xor U9489 (N_9489,N_4276,N_2555);
nand U9490 (N_9490,N_3560,N_3717);
or U9491 (N_9491,N_1205,N_3438);
nand U9492 (N_9492,N_2577,N_2607);
and U9493 (N_9493,N_545,N_746);
and U9494 (N_9494,N_4910,N_4510);
nand U9495 (N_9495,N_4129,N_3214);
nor U9496 (N_9496,N_2747,N_4451);
or U9497 (N_9497,N_228,N_2609);
and U9498 (N_9498,N_4725,N_3460);
and U9499 (N_9499,N_444,N_237);
nand U9500 (N_9500,N_2802,N_312);
or U9501 (N_9501,N_2138,N_1535);
and U9502 (N_9502,N_2999,N_3499);
and U9503 (N_9503,N_3260,N_4626);
nand U9504 (N_9504,N_30,N_25);
or U9505 (N_9505,N_1328,N_170);
or U9506 (N_9506,N_4463,N_4363);
nor U9507 (N_9507,N_1295,N_981);
and U9508 (N_9508,N_2782,N_4682);
nand U9509 (N_9509,N_2431,N_1194);
or U9510 (N_9510,N_4622,N_4774);
nor U9511 (N_9511,N_877,N_1080);
nor U9512 (N_9512,N_2545,N_1886);
and U9513 (N_9513,N_3548,N_2695);
and U9514 (N_9514,N_3091,N_1898);
and U9515 (N_9515,N_2369,N_311);
xnor U9516 (N_9516,N_4036,N_3642);
nand U9517 (N_9517,N_671,N_4900);
or U9518 (N_9518,N_2798,N_2799);
or U9519 (N_9519,N_1040,N_848);
nand U9520 (N_9520,N_3384,N_4458);
nand U9521 (N_9521,N_1239,N_3661);
nand U9522 (N_9522,N_3049,N_4269);
and U9523 (N_9523,N_160,N_3055);
and U9524 (N_9524,N_1766,N_2838);
or U9525 (N_9525,N_4220,N_3418);
nand U9526 (N_9526,N_3537,N_3335);
or U9527 (N_9527,N_317,N_1637);
or U9528 (N_9528,N_2806,N_535);
or U9529 (N_9529,N_2923,N_4584);
nand U9530 (N_9530,N_1086,N_616);
nor U9531 (N_9531,N_1495,N_2478);
or U9532 (N_9532,N_2197,N_1028);
or U9533 (N_9533,N_3642,N_2569);
nand U9534 (N_9534,N_226,N_2212);
nor U9535 (N_9535,N_4955,N_3103);
or U9536 (N_9536,N_1239,N_279);
nand U9537 (N_9537,N_4723,N_4194);
nand U9538 (N_9538,N_1179,N_901);
and U9539 (N_9539,N_1454,N_1746);
or U9540 (N_9540,N_3148,N_3576);
or U9541 (N_9541,N_4339,N_3302);
nand U9542 (N_9542,N_3581,N_2291);
or U9543 (N_9543,N_4204,N_3575);
and U9544 (N_9544,N_3648,N_1154);
nand U9545 (N_9545,N_1892,N_3403);
or U9546 (N_9546,N_998,N_3488);
nand U9547 (N_9547,N_2106,N_2529);
or U9548 (N_9548,N_4278,N_1158);
or U9549 (N_9549,N_1487,N_1687);
nor U9550 (N_9550,N_3028,N_1863);
or U9551 (N_9551,N_1685,N_1355);
nand U9552 (N_9552,N_3716,N_1690);
nand U9553 (N_9553,N_1619,N_1899);
and U9554 (N_9554,N_3919,N_4468);
nand U9555 (N_9555,N_2483,N_761);
nand U9556 (N_9556,N_3099,N_1814);
nor U9557 (N_9557,N_241,N_1385);
and U9558 (N_9558,N_1601,N_53);
nand U9559 (N_9559,N_113,N_585);
or U9560 (N_9560,N_442,N_1024);
nand U9561 (N_9561,N_2634,N_403);
or U9562 (N_9562,N_3513,N_1937);
or U9563 (N_9563,N_1249,N_1146);
or U9564 (N_9564,N_2449,N_4393);
nand U9565 (N_9565,N_3801,N_1224);
nand U9566 (N_9566,N_1944,N_3313);
or U9567 (N_9567,N_3856,N_2974);
or U9568 (N_9568,N_803,N_4770);
nor U9569 (N_9569,N_3707,N_3821);
and U9570 (N_9570,N_4482,N_1549);
and U9571 (N_9571,N_2594,N_2607);
nor U9572 (N_9572,N_758,N_4955);
nor U9573 (N_9573,N_1600,N_3588);
nor U9574 (N_9574,N_4417,N_1136);
or U9575 (N_9575,N_2050,N_367);
nand U9576 (N_9576,N_3183,N_2804);
and U9577 (N_9577,N_1573,N_4987);
or U9578 (N_9578,N_2257,N_129);
or U9579 (N_9579,N_1139,N_2582);
xnor U9580 (N_9580,N_2046,N_3642);
nor U9581 (N_9581,N_2169,N_429);
and U9582 (N_9582,N_6,N_4630);
and U9583 (N_9583,N_783,N_2281);
nand U9584 (N_9584,N_3688,N_1511);
nand U9585 (N_9585,N_2555,N_2962);
or U9586 (N_9586,N_2209,N_3876);
and U9587 (N_9587,N_1408,N_796);
and U9588 (N_9588,N_4847,N_1251);
nand U9589 (N_9589,N_4272,N_243);
nand U9590 (N_9590,N_121,N_403);
nor U9591 (N_9591,N_4363,N_1041);
and U9592 (N_9592,N_4601,N_1660);
nor U9593 (N_9593,N_4850,N_3362);
or U9594 (N_9594,N_595,N_2695);
and U9595 (N_9595,N_2152,N_384);
nor U9596 (N_9596,N_1624,N_4395);
or U9597 (N_9597,N_3632,N_3704);
nand U9598 (N_9598,N_4654,N_2339);
or U9599 (N_9599,N_1015,N_3886);
or U9600 (N_9600,N_1879,N_944);
or U9601 (N_9601,N_1964,N_1888);
and U9602 (N_9602,N_4740,N_1548);
and U9603 (N_9603,N_3639,N_2430);
or U9604 (N_9604,N_3220,N_4739);
or U9605 (N_9605,N_1361,N_3899);
nand U9606 (N_9606,N_3058,N_4469);
and U9607 (N_9607,N_2180,N_1093);
or U9608 (N_9608,N_993,N_4410);
nand U9609 (N_9609,N_284,N_4540);
or U9610 (N_9610,N_2326,N_3809);
and U9611 (N_9611,N_4389,N_3047);
nor U9612 (N_9612,N_3241,N_85);
or U9613 (N_9613,N_1059,N_1199);
and U9614 (N_9614,N_4957,N_1141);
and U9615 (N_9615,N_1057,N_4815);
or U9616 (N_9616,N_1457,N_77);
or U9617 (N_9617,N_428,N_4242);
and U9618 (N_9618,N_2692,N_359);
and U9619 (N_9619,N_2501,N_2040);
and U9620 (N_9620,N_2324,N_85);
nand U9621 (N_9621,N_795,N_2976);
or U9622 (N_9622,N_1386,N_2297);
and U9623 (N_9623,N_2306,N_1091);
nand U9624 (N_9624,N_1241,N_2456);
and U9625 (N_9625,N_1790,N_2738);
and U9626 (N_9626,N_4882,N_2629);
and U9627 (N_9627,N_2832,N_2891);
nor U9628 (N_9628,N_1221,N_3260);
or U9629 (N_9629,N_3019,N_1788);
nand U9630 (N_9630,N_821,N_2567);
nand U9631 (N_9631,N_1606,N_1441);
nor U9632 (N_9632,N_4767,N_1480);
nand U9633 (N_9633,N_2806,N_517);
and U9634 (N_9634,N_2705,N_4846);
xor U9635 (N_9635,N_4922,N_1392);
and U9636 (N_9636,N_4325,N_962);
nand U9637 (N_9637,N_3970,N_1804);
and U9638 (N_9638,N_2333,N_68);
nor U9639 (N_9639,N_51,N_3325);
and U9640 (N_9640,N_1302,N_1367);
nor U9641 (N_9641,N_1490,N_1304);
xnor U9642 (N_9642,N_4237,N_2401);
and U9643 (N_9643,N_3544,N_899);
nand U9644 (N_9644,N_3567,N_541);
and U9645 (N_9645,N_14,N_4491);
xor U9646 (N_9646,N_2403,N_1039);
nor U9647 (N_9647,N_3564,N_620);
nand U9648 (N_9648,N_170,N_34);
or U9649 (N_9649,N_4714,N_4993);
nand U9650 (N_9650,N_551,N_4328);
and U9651 (N_9651,N_4582,N_978);
nor U9652 (N_9652,N_1169,N_695);
or U9653 (N_9653,N_4371,N_1180);
or U9654 (N_9654,N_3003,N_3636);
or U9655 (N_9655,N_486,N_304);
or U9656 (N_9656,N_1280,N_1842);
nor U9657 (N_9657,N_707,N_341);
nor U9658 (N_9658,N_3553,N_1757);
nand U9659 (N_9659,N_2549,N_1692);
or U9660 (N_9660,N_2745,N_542);
xnor U9661 (N_9661,N_3436,N_1912);
and U9662 (N_9662,N_1332,N_4643);
and U9663 (N_9663,N_4315,N_808);
or U9664 (N_9664,N_2676,N_3898);
nor U9665 (N_9665,N_1846,N_1);
or U9666 (N_9666,N_904,N_1961);
and U9667 (N_9667,N_4963,N_40);
and U9668 (N_9668,N_4550,N_4056);
and U9669 (N_9669,N_3410,N_2546);
nor U9670 (N_9670,N_1046,N_2518);
nor U9671 (N_9671,N_4559,N_2873);
nor U9672 (N_9672,N_2665,N_4682);
or U9673 (N_9673,N_3059,N_1183);
nor U9674 (N_9674,N_4180,N_3253);
or U9675 (N_9675,N_2057,N_4495);
or U9676 (N_9676,N_1754,N_1449);
and U9677 (N_9677,N_4292,N_2697);
or U9678 (N_9678,N_2202,N_3712);
nor U9679 (N_9679,N_1355,N_1720);
or U9680 (N_9680,N_4193,N_2007);
or U9681 (N_9681,N_761,N_1020);
or U9682 (N_9682,N_1206,N_459);
nor U9683 (N_9683,N_84,N_397);
nor U9684 (N_9684,N_3707,N_506);
nand U9685 (N_9685,N_3248,N_84);
and U9686 (N_9686,N_4107,N_1793);
and U9687 (N_9687,N_3692,N_3622);
nand U9688 (N_9688,N_2989,N_2353);
and U9689 (N_9689,N_4913,N_1992);
nand U9690 (N_9690,N_3129,N_4562);
and U9691 (N_9691,N_4168,N_4470);
or U9692 (N_9692,N_3825,N_3965);
nor U9693 (N_9693,N_118,N_1644);
nor U9694 (N_9694,N_4598,N_1744);
or U9695 (N_9695,N_33,N_4548);
or U9696 (N_9696,N_1199,N_813);
nor U9697 (N_9697,N_637,N_1326);
nor U9698 (N_9698,N_2745,N_2250);
nor U9699 (N_9699,N_3894,N_1935);
nor U9700 (N_9700,N_383,N_1244);
or U9701 (N_9701,N_4852,N_554);
nor U9702 (N_9702,N_2871,N_4770);
or U9703 (N_9703,N_4481,N_4427);
nand U9704 (N_9704,N_102,N_4198);
nand U9705 (N_9705,N_3575,N_588);
nor U9706 (N_9706,N_1071,N_2754);
or U9707 (N_9707,N_2403,N_4313);
nand U9708 (N_9708,N_2593,N_4055);
and U9709 (N_9709,N_232,N_819);
or U9710 (N_9710,N_2072,N_4153);
nand U9711 (N_9711,N_2234,N_237);
nand U9712 (N_9712,N_2367,N_977);
or U9713 (N_9713,N_3490,N_3841);
nor U9714 (N_9714,N_2627,N_4570);
or U9715 (N_9715,N_2028,N_2742);
xor U9716 (N_9716,N_1448,N_1881);
nand U9717 (N_9717,N_369,N_2692);
and U9718 (N_9718,N_2554,N_1933);
and U9719 (N_9719,N_2292,N_4427);
or U9720 (N_9720,N_1756,N_3995);
nor U9721 (N_9721,N_1734,N_1622);
and U9722 (N_9722,N_1214,N_1292);
or U9723 (N_9723,N_381,N_2066);
nand U9724 (N_9724,N_971,N_1193);
and U9725 (N_9725,N_3504,N_1164);
nor U9726 (N_9726,N_4944,N_3023);
nor U9727 (N_9727,N_661,N_86);
nor U9728 (N_9728,N_380,N_2519);
nand U9729 (N_9729,N_601,N_73);
xor U9730 (N_9730,N_268,N_3672);
nor U9731 (N_9731,N_1907,N_2836);
or U9732 (N_9732,N_3585,N_3323);
and U9733 (N_9733,N_4688,N_3250);
nor U9734 (N_9734,N_1994,N_2358);
nand U9735 (N_9735,N_1217,N_1517);
nand U9736 (N_9736,N_4795,N_3799);
and U9737 (N_9737,N_4870,N_1584);
and U9738 (N_9738,N_2465,N_2410);
nand U9739 (N_9739,N_357,N_1838);
xnor U9740 (N_9740,N_4849,N_350);
nand U9741 (N_9741,N_776,N_4839);
nor U9742 (N_9742,N_4088,N_4368);
nand U9743 (N_9743,N_2185,N_3185);
nand U9744 (N_9744,N_1349,N_561);
and U9745 (N_9745,N_4416,N_3129);
nand U9746 (N_9746,N_1052,N_1077);
nor U9747 (N_9747,N_3319,N_4453);
and U9748 (N_9748,N_3617,N_1575);
and U9749 (N_9749,N_1305,N_1532);
nand U9750 (N_9750,N_3841,N_2190);
nand U9751 (N_9751,N_3330,N_3899);
nand U9752 (N_9752,N_2569,N_4625);
nand U9753 (N_9753,N_3847,N_1143);
nand U9754 (N_9754,N_3318,N_679);
and U9755 (N_9755,N_3822,N_3675);
and U9756 (N_9756,N_133,N_1143);
and U9757 (N_9757,N_2977,N_4951);
or U9758 (N_9758,N_239,N_384);
nand U9759 (N_9759,N_3259,N_2879);
nand U9760 (N_9760,N_1567,N_25);
and U9761 (N_9761,N_1522,N_207);
nand U9762 (N_9762,N_3379,N_4503);
nand U9763 (N_9763,N_1366,N_2987);
nand U9764 (N_9764,N_853,N_4424);
or U9765 (N_9765,N_1662,N_1764);
and U9766 (N_9766,N_2330,N_1972);
and U9767 (N_9767,N_204,N_1933);
nand U9768 (N_9768,N_3381,N_371);
nor U9769 (N_9769,N_4996,N_989);
or U9770 (N_9770,N_366,N_3161);
nand U9771 (N_9771,N_2022,N_216);
nor U9772 (N_9772,N_133,N_1997);
nor U9773 (N_9773,N_1332,N_3651);
and U9774 (N_9774,N_2598,N_4040);
or U9775 (N_9775,N_3032,N_4986);
nor U9776 (N_9776,N_2750,N_2695);
or U9777 (N_9777,N_4905,N_1996);
nor U9778 (N_9778,N_721,N_3108);
or U9779 (N_9779,N_2051,N_1932);
nand U9780 (N_9780,N_135,N_1240);
and U9781 (N_9781,N_1941,N_4905);
or U9782 (N_9782,N_4562,N_4585);
or U9783 (N_9783,N_4735,N_1362);
nor U9784 (N_9784,N_969,N_4514);
or U9785 (N_9785,N_4219,N_899);
nor U9786 (N_9786,N_3349,N_2414);
and U9787 (N_9787,N_2263,N_2455);
and U9788 (N_9788,N_4841,N_4147);
nand U9789 (N_9789,N_2056,N_942);
or U9790 (N_9790,N_1414,N_1349);
and U9791 (N_9791,N_1896,N_4181);
nand U9792 (N_9792,N_3849,N_4100);
nor U9793 (N_9793,N_2556,N_4745);
and U9794 (N_9794,N_178,N_3934);
and U9795 (N_9795,N_4287,N_621);
nor U9796 (N_9796,N_1221,N_4583);
and U9797 (N_9797,N_2332,N_3121);
nand U9798 (N_9798,N_460,N_2190);
and U9799 (N_9799,N_42,N_1467);
nor U9800 (N_9800,N_3503,N_1984);
or U9801 (N_9801,N_356,N_2354);
nor U9802 (N_9802,N_2380,N_419);
or U9803 (N_9803,N_1226,N_1455);
or U9804 (N_9804,N_2320,N_447);
and U9805 (N_9805,N_2550,N_960);
and U9806 (N_9806,N_4129,N_44);
nand U9807 (N_9807,N_582,N_4199);
nand U9808 (N_9808,N_1652,N_1744);
xnor U9809 (N_9809,N_4341,N_3954);
and U9810 (N_9810,N_1717,N_4795);
nor U9811 (N_9811,N_1361,N_1489);
and U9812 (N_9812,N_4811,N_629);
nor U9813 (N_9813,N_2826,N_4466);
or U9814 (N_9814,N_125,N_4656);
or U9815 (N_9815,N_712,N_2782);
or U9816 (N_9816,N_1203,N_4981);
and U9817 (N_9817,N_2755,N_2781);
nand U9818 (N_9818,N_717,N_4528);
nand U9819 (N_9819,N_1835,N_127);
and U9820 (N_9820,N_1552,N_3345);
and U9821 (N_9821,N_727,N_550);
or U9822 (N_9822,N_4173,N_650);
nor U9823 (N_9823,N_48,N_2678);
or U9824 (N_9824,N_4944,N_200);
and U9825 (N_9825,N_1863,N_4487);
and U9826 (N_9826,N_4466,N_3424);
and U9827 (N_9827,N_4637,N_3641);
or U9828 (N_9828,N_3904,N_2266);
and U9829 (N_9829,N_1064,N_2966);
nand U9830 (N_9830,N_446,N_474);
and U9831 (N_9831,N_1061,N_4813);
and U9832 (N_9832,N_665,N_539);
nand U9833 (N_9833,N_539,N_1920);
or U9834 (N_9834,N_2195,N_2073);
or U9835 (N_9835,N_4341,N_4633);
nand U9836 (N_9836,N_4789,N_4589);
and U9837 (N_9837,N_3718,N_4084);
nor U9838 (N_9838,N_2720,N_1152);
or U9839 (N_9839,N_430,N_1623);
nor U9840 (N_9840,N_4350,N_4021);
nand U9841 (N_9841,N_3943,N_3373);
or U9842 (N_9842,N_3681,N_3103);
and U9843 (N_9843,N_2776,N_2752);
nor U9844 (N_9844,N_2208,N_505);
and U9845 (N_9845,N_1428,N_3755);
nand U9846 (N_9846,N_2432,N_702);
or U9847 (N_9847,N_1572,N_599);
or U9848 (N_9848,N_2311,N_1452);
nand U9849 (N_9849,N_1793,N_953);
or U9850 (N_9850,N_1411,N_10);
nand U9851 (N_9851,N_3497,N_732);
nor U9852 (N_9852,N_2630,N_3729);
nand U9853 (N_9853,N_2040,N_3103);
nor U9854 (N_9854,N_2982,N_2487);
or U9855 (N_9855,N_1507,N_3990);
nand U9856 (N_9856,N_743,N_444);
and U9857 (N_9857,N_627,N_408);
or U9858 (N_9858,N_3112,N_3083);
nand U9859 (N_9859,N_3888,N_4351);
and U9860 (N_9860,N_3134,N_3084);
and U9861 (N_9861,N_2928,N_2554);
nand U9862 (N_9862,N_858,N_1196);
nor U9863 (N_9863,N_501,N_946);
nand U9864 (N_9864,N_622,N_3990);
nor U9865 (N_9865,N_877,N_3895);
nor U9866 (N_9866,N_3034,N_2248);
and U9867 (N_9867,N_4095,N_2492);
nor U9868 (N_9868,N_386,N_4597);
nand U9869 (N_9869,N_4668,N_4959);
or U9870 (N_9870,N_474,N_1808);
and U9871 (N_9871,N_541,N_3213);
and U9872 (N_9872,N_2391,N_2105);
or U9873 (N_9873,N_4091,N_3255);
nor U9874 (N_9874,N_3392,N_1538);
and U9875 (N_9875,N_3912,N_3373);
and U9876 (N_9876,N_2266,N_1816);
nand U9877 (N_9877,N_1876,N_3039);
and U9878 (N_9878,N_3578,N_2914);
or U9879 (N_9879,N_3559,N_1077);
and U9880 (N_9880,N_3244,N_678);
nor U9881 (N_9881,N_4529,N_1211);
or U9882 (N_9882,N_3085,N_3783);
nand U9883 (N_9883,N_4783,N_4499);
nor U9884 (N_9884,N_3137,N_852);
nand U9885 (N_9885,N_4234,N_831);
or U9886 (N_9886,N_2359,N_4854);
nand U9887 (N_9887,N_2493,N_2144);
nor U9888 (N_9888,N_3586,N_4964);
nor U9889 (N_9889,N_203,N_1693);
or U9890 (N_9890,N_3992,N_4560);
or U9891 (N_9891,N_2023,N_2908);
nor U9892 (N_9892,N_2365,N_1377);
and U9893 (N_9893,N_1780,N_2497);
and U9894 (N_9894,N_686,N_4888);
xor U9895 (N_9895,N_3100,N_3153);
and U9896 (N_9896,N_1536,N_3008);
nor U9897 (N_9897,N_3162,N_1116);
and U9898 (N_9898,N_4637,N_3116);
and U9899 (N_9899,N_2311,N_1808);
nand U9900 (N_9900,N_792,N_1572);
nand U9901 (N_9901,N_1454,N_1255);
or U9902 (N_9902,N_1312,N_3231);
nor U9903 (N_9903,N_1196,N_767);
and U9904 (N_9904,N_638,N_570);
nand U9905 (N_9905,N_4997,N_2582);
nor U9906 (N_9906,N_4452,N_1571);
nor U9907 (N_9907,N_1623,N_938);
nor U9908 (N_9908,N_1790,N_2972);
nor U9909 (N_9909,N_2221,N_1842);
xnor U9910 (N_9910,N_3029,N_3060);
or U9911 (N_9911,N_1420,N_4982);
and U9912 (N_9912,N_540,N_4552);
and U9913 (N_9913,N_4974,N_890);
nand U9914 (N_9914,N_678,N_2836);
and U9915 (N_9915,N_1566,N_4651);
nand U9916 (N_9916,N_1062,N_3798);
nand U9917 (N_9917,N_3667,N_560);
nand U9918 (N_9918,N_2468,N_2829);
and U9919 (N_9919,N_3963,N_3205);
and U9920 (N_9920,N_225,N_4986);
nand U9921 (N_9921,N_3180,N_4171);
or U9922 (N_9922,N_806,N_344);
nor U9923 (N_9923,N_352,N_3856);
and U9924 (N_9924,N_2568,N_2001);
and U9925 (N_9925,N_3515,N_4744);
nand U9926 (N_9926,N_831,N_2627);
or U9927 (N_9927,N_1649,N_1783);
or U9928 (N_9928,N_349,N_1896);
and U9929 (N_9929,N_3562,N_3831);
nor U9930 (N_9930,N_210,N_1404);
or U9931 (N_9931,N_2177,N_160);
and U9932 (N_9932,N_3837,N_3207);
nand U9933 (N_9933,N_3279,N_3117);
and U9934 (N_9934,N_4230,N_1324);
nand U9935 (N_9935,N_937,N_2589);
nand U9936 (N_9936,N_3546,N_8);
or U9937 (N_9937,N_2111,N_3819);
or U9938 (N_9938,N_4810,N_4669);
and U9939 (N_9939,N_3194,N_1236);
and U9940 (N_9940,N_387,N_2709);
and U9941 (N_9941,N_3830,N_4593);
nand U9942 (N_9942,N_1927,N_76);
nor U9943 (N_9943,N_2137,N_307);
nand U9944 (N_9944,N_2044,N_4377);
nand U9945 (N_9945,N_1643,N_4741);
and U9946 (N_9946,N_2911,N_1113);
nor U9947 (N_9947,N_1996,N_1766);
nor U9948 (N_9948,N_3564,N_2291);
nand U9949 (N_9949,N_130,N_1473);
nand U9950 (N_9950,N_3595,N_1314);
nand U9951 (N_9951,N_4664,N_706);
nand U9952 (N_9952,N_1303,N_410);
or U9953 (N_9953,N_4673,N_466);
or U9954 (N_9954,N_3460,N_169);
xor U9955 (N_9955,N_1487,N_1199);
nor U9956 (N_9956,N_3394,N_2378);
nand U9957 (N_9957,N_2312,N_3655);
or U9958 (N_9958,N_3290,N_1060);
nand U9959 (N_9959,N_430,N_1750);
nor U9960 (N_9960,N_3728,N_823);
or U9961 (N_9961,N_664,N_2274);
and U9962 (N_9962,N_3064,N_1846);
and U9963 (N_9963,N_3092,N_3918);
nor U9964 (N_9964,N_3384,N_4024);
or U9965 (N_9965,N_115,N_924);
and U9966 (N_9966,N_4795,N_3993);
or U9967 (N_9967,N_855,N_695);
and U9968 (N_9968,N_547,N_1360);
or U9969 (N_9969,N_3966,N_2924);
or U9970 (N_9970,N_829,N_4606);
nor U9971 (N_9971,N_2009,N_3660);
nor U9972 (N_9972,N_662,N_1166);
or U9973 (N_9973,N_793,N_4961);
or U9974 (N_9974,N_1108,N_3470);
or U9975 (N_9975,N_3603,N_1215);
and U9976 (N_9976,N_3577,N_1392);
nand U9977 (N_9977,N_4098,N_3979);
and U9978 (N_9978,N_1679,N_4800);
or U9979 (N_9979,N_2298,N_4282);
nor U9980 (N_9980,N_1241,N_3030);
and U9981 (N_9981,N_3207,N_4296);
and U9982 (N_9982,N_2410,N_4018);
or U9983 (N_9983,N_4866,N_2599);
nand U9984 (N_9984,N_2538,N_4392);
or U9985 (N_9985,N_4280,N_1769);
xnor U9986 (N_9986,N_380,N_588);
nand U9987 (N_9987,N_106,N_1971);
nand U9988 (N_9988,N_3545,N_2908);
and U9989 (N_9989,N_1464,N_4365);
and U9990 (N_9990,N_91,N_355);
nand U9991 (N_9991,N_2383,N_1371);
and U9992 (N_9992,N_1680,N_2166);
and U9993 (N_9993,N_2762,N_1620);
nor U9994 (N_9994,N_1741,N_1530);
or U9995 (N_9995,N_987,N_1516);
or U9996 (N_9996,N_3172,N_1881);
nand U9997 (N_9997,N_1126,N_2628);
nand U9998 (N_9998,N_1254,N_1745);
nand U9999 (N_9999,N_586,N_1635);
nor U10000 (N_10000,N_8776,N_7613);
nand U10001 (N_10001,N_7183,N_6828);
or U10002 (N_10002,N_7521,N_7588);
nor U10003 (N_10003,N_7676,N_9073);
and U10004 (N_10004,N_6583,N_6465);
or U10005 (N_10005,N_6692,N_7564);
nand U10006 (N_10006,N_9991,N_7773);
and U10007 (N_10007,N_8054,N_6187);
nand U10008 (N_10008,N_9317,N_9175);
and U10009 (N_10009,N_5822,N_6161);
or U10010 (N_10010,N_6594,N_6969);
nand U10011 (N_10011,N_6658,N_5545);
and U10012 (N_10012,N_9330,N_5236);
nand U10013 (N_10013,N_9208,N_5271);
nor U10014 (N_10014,N_7228,N_9614);
nor U10015 (N_10015,N_7808,N_6278);
or U10016 (N_10016,N_9830,N_6900);
nand U10017 (N_10017,N_6996,N_6769);
nor U10018 (N_10018,N_9191,N_8478);
and U10019 (N_10019,N_7212,N_9406);
or U10020 (N_10020,N_6163,N_8310);
nand U10021 (N_10021,N_5075,N_6604);
or U10022 (N_10022,N_5280,N_9782);
nand U10023 (N_10023,N_7900,N_5473);
or U10024 (N_10024,N_7140,N_5290);
nand U10025 (N_10025,N_6848,N_5849);
nor U10026 (N_10026,N_7738,N_7250);
nand U10027 (N_10027,N_9407,N_6506);
nor U10028 (N_10028,N_6273,N_9826);
nand U10029 (N_10029,N_7619,N_9138);
nand U10030 (N_10030,N_6007,N_7753);
nor U10031 (N_10031,N_6770,N_7560);
nor U10032 (N_10032,N_7308,N_7734);
or U10033 (N_10033,N_8167,N_6431);
or U10034 (N_10034,N_7710,N_7686);
nand U10035 (N_10035,N_5529,N_5159);
or U10036 (N_10036,N_7550,N_8994);
and U10037 (N_10037,N_8940,N_7713);
nor U10038 (N_10038,N_6182,N_7364);
nand U10039 (N_10039,N_5502,N_6002);
xnor U10040 (N_10040,N_9865,N_8085);
nand U10041 (N_10041,N_6829,N_9468);
nor U10042 (N_10042,N_5284,N_6267);
nand U10043 (N_10043,N_8065,N_8836);
nand U10044 (N_10044,N_5559,N_6740);
nand U10045 (N_10045,N_7598,N_5638);
and U10046 (N_10046,N_6189,N_8526);
or U10047 (N_10047,N_9464,N_8709);
nand U10048 (N_10048,N_8342,N_9291);
nor U10049 (N_10049,N_5828,N_7476);
or U10050 (N_10050,N_5999,N_8950);
nand U10051 (N_10051,N_5659,N_8520);
nand U10052 (N_10052,N_9557,N_7681);
nor U10053 (N_10053,N_8482,N_6176);
and U10054 (N_10054,N_7971,N_5338);
nor U10055 (N_10055,N_8751,N_8913);
or U10056 (N_10056,N_7406,N_5922);
nor U10057 (N_10057,N_7709,N_5371);
nand U10058 (N_10058,N_7347,N_8373);
or U10059 (N_10059,N_7336,N_7345);
and U10060 (N_10060,N_8487,N_8743);
nand U10061 (N_10061,N_9538,N_7885);
nand U10062 (N_10062,N_6058,N_5016);
or U10063 (N_10063,N_7931,N_6854);
or U10064 (N_10064,N_5213,N_7647);
nand U10065 (N_10065,N_9189,N_9900);
and U10066 (N_10066,N_7580,N_6018);
nor U10067 (N_10067,N_6714,N_8534);
nand U10068 (N_10068,N_6207,N_7174);
nand U10069 (N_10069,N_5851,N_5147);
and U10070 (N_10070,N_8860,N_8738);
nor U10071 (N_10071,N_6659,N_8975);
xor U10072 (N_10072,N_6721,N_8053);
nor U10073 (N_10073,N_9670,N_7634);
nand U10074 (N_10074,N_9853,N_9856);
or U10075 (N_10075,N_6496,N_8817);
nor U10076 (N_10076,N_5496,N_9397);
nor U10077 (N_10077,N_5649,N_8437);
xor U10078 (N_10078,N_7405,N_6832);
or U10079 (N_10079,N_7987,N_5970);
xor U10080 (N_10080,N_8544,N_8796);
nand U10081 (N_10081,N_5230,N_7799);
and U10082 (N_10082,N_5202,N_7671);
nand U10083 (N_10083,N_9551,N_8164);
nor U10084 (N_10084,N_6629,N_6749);
or U10085 (N_10085,N_9163,N_9558);
nand U10086 (N_10086,N_7302,N_7968);
nand U10087 (N_10087,N_7672,N_6849);
or U10088 (N_10088,N_7327,N_7126);
nor U10089 (N_10089,N_6787,N_5246);
or U10090 (N_10090,N_9320,N_5848);
nand U10091 (N_10091,N_6093,N_6766);
nor U10092 (N_10092,N_9343,N_9861);
and U10093 (N_10093,N_8171,N_6743);
and U10094 (N_10094,N_8283,N_6747);
nor U10095 (N_10095,N_6693,N_6455);
nand U10096 (N_10096,N_7068,N_5556);
or U10097 (N_10097,N_6222,N_5551);
nand U10098 (N_10098,N_6818,N_9592);
and U10099 (N_10099,N_9339,N_6399);
or U10100 (N_10100,N_9239,N_6905);
nor U10101 (N_10101,N_9076,N_5988);
nand U10102 (N_10102,N_9840,N_8648);
nand U10103 (N_10103,N_8925,N_7691);
and U10104 (N_10104,N_5198,N_8459);
or U10105 (N_10105,N_7537,N_8308);
and U10106 (N_10106,N_8550,N_6072);
nand U10107 (N_10107,N_9028,N_6188);
nand U10108 (N_10108,N_7760,N_5211);
nand U10109 (N_10109,N_5477,N_5486);
or U10110 (N_10110,N_5681,N_7571);
or U10111 (N_10111,N_9618,N_5466);
nand U10112 (N_10112,N_8402,N_7898);
nand U10113 (N_10113,N_8222,N_7323);
and U10114 (N_10114,N_6952,N_8151);
nand U10115 (N_10115,N_5569,N_5282);
nand U10116 (N_10116,N_6193,N_6197);
nor U10117 (N_10117,N_8233,N_6819);
and U10118 (N_10118,N_8503,N_6888);
nor U10119 (N_10119,N_8824,N_9103);
nor U10120 (N_10120,N_7304,N_8447);
and U10121 (N_10121,N_5878,N_5294);
and U10122 (N_10122,N_7023,N_6560);
nor U10123 (N_10123,N_7121,N_8168);
nand U10124 (N_10124,N_5967,N_7226);
and U10125 (N_10125,N_9367,N_6232);
or U10126 (N_10126,N_8299,N_7398);
nor U10127 (N_10127,N_7736,N_8440);
and U10128 (N_10128,N_7563,N_5724);
and U10129 (N_10129,N_8545,N_6263);
and U10130 (N_10130,N_6165,N_8837);
or U10131 (N_10131,N_6410,N_5357);
or U10132 (N_10132,N_9294,N_8352);
nand U10133 (N_10133,N_8135,N_5958);
xnor U10134 (N_10134,N_5074,N_7943);
or U10135 (N_10135,N_7331,N_9017);
nand U10136 (N_10136,N_8445,N_6785);
and U10137 (N_10137,N_7150,N_9411);
or U10138 (N_10138,N_6881,N_6094);
nand U10139 (N_10139,N_8006,N_6215);
and U10140 (N_10140,N_8987,N_8623);
nor U10141 (N_10141,N_9186,N_7587);
nand U10142 (N_10142,N_7101,N_9067);
nand U10143 (N_10143,N_8613,N_6964);
and U10144 (N_10144,N_7063,N_7219);
and U10145 (N_10145,N_5492,N_8281);
and U10146 (N_10146,N_8176,N_7396);
nor U10147 (N_10147,N_7813,N_9655);
nand U10148 (N_10148,N_6100,N_6809);
or U10149 (N_10149,N_5459,N_7471);
nor U10150 (N_10150,N_5188,N_7969);
nand U10151 (N_10151,N_9342,N_8013);
and U10152 (N_10152,N_7667,N_8527);
and U10153 (N_10153,N_8209,N_8026);
and U10154 (N_10154,N_9940,N_5021);
and U10155 (N_10155,N_5637,N_6739);
nor U10156 (N_10156,N_5445,N_5043);
nor U10157 (N_10157,N_9525,N_9431);
or U10158 (N_10158,N_5422,N_5648);
nor U10159 (N_10159,N_9135,N_8429);
nor U10160 (N_10160,N_7363,N_8384);
nand U10161 (N_10161,N_5312,N_6471);
nand U10162 (N_10162,N_8842,N_9668);
and U10163 (N_10163,N_5843,N_7169);
and U10164 (N_10164,N_5789,N_6039);
or U10165 (N_10165,N_6599,N_7459);
or U10166 (N_10166,N_7535,N_6154);
and U10167 (N_10167,N_9448,N_5864);
nor U10168 (N_10168,N_9494,N_6311);
or U10169 (N_10169,N_8884,N_9851);
and U10170 (N_10170,N_7849,N_6918);
and U10171 (N_10171,N_8242,N_8590);
nand U10172 (N_10172,N_6209,N_8676);
nand U10173 (N_10173,N_9504,N_7575);
xnor U10174 (N_10174,N_6283,N_8833);
or U10175 (N_10175,N_5114,N_7177);
or U10176 (N_10176,N_5933,N_8055);
or U10177 (N_10177,N_6525,N_5291);
nor U10178 (N_10178,N_9847,N_5417);
or U10179 (N_10179,N_8268,N_5152);
or U10180 (N_10180,N_8638,N_8827);
or U10181 (N_10181,N_9039,N_7367);
nor U10182 (N_10182,N_8543,N_8529);
or U10183 (N_10183,N_6711,N_5839);
or U10184 (N_10184,N_5436,N_8655);
or U10185 (N_10185,N_7907,N_8202);
or U10186 (N_10186,N_7292,N_8782);
nor U10187 (N_10187,N_7862,N_6902);
or U10188 (N_10188,N_7284,N_5019);
and U10189 (N_10189,N_5050,N_9071);
nand U10190 (N_10190,N_6345,N_6622);
or U10191 (N_10191,N_6571,N_8274);
nor U10192 (N_10192,N_9555,N_5966);
nor U10193 (N_10193,N_8442,N_7489);
nor U10194 (N_10194,N_5858,N_8012);
nor U10195 (N_10195,N_9562,N_9838);
nor U10196 (N_10196,N_5539,N_9619);
nor U10197 (N_10197,N_8536,N_6316);
nand U10198 (N_10198,N_7558,N_8811);
nand U10199 (N_10199,N_5158,N_6082);
or U10200 (N_10200,N_6020,N_7233);
xnor U10201 (N_10201,N_9285,N_7963);
nor U10202 (N_10202,N_7990,N_8554);
nand U10203 (N_10203,N_5454,N_8667);
nand U10204 (N_10204,N_7958,N_9395);
or U10205 (N_10205,N_7824,N_9387);
and U10206 (N_10206,N_5331,N_6166);
or U10207 (N_10207,N_8519,N_9211);
nand U10208 (N_10208,N_9055,N_6611);
or U10209 (N_10209,N_9245,N_7133);
nor U10210 (N_10210,N_8713,N_8084);
and U10211 (N_10211,N_6006,N_6130);
and U10212 (N_10212,N_6680,N_7790);
nor U10213 (N_10213,N_8309,N_6485);
or U10214 (N_10214,N_8294,N_9125);
and U10215 (N_10215,N_7225,N_9066);
and U10216 (N_10216,N_5034,N_7478);
nor U10217 (N_10217,N_8787,N_6035);
or U10218 (N_10218,N_9344,N_9750);
nand U10219 (N_10219,N_9476,N_9689);
and U10220 (N_10220,N_8301,N_7015);
nor U10221 (N_10221,N_6735,N_6127);
nand U10222 (N_10222,N_9503,N_8637);
and U10223 (N_10223,N_9000,N_6225);
or U10224 (N_10224,N_6073,N_7751);
nor U10225 (N_10225,N_8145,N_5541);
and U10226 (N_10226,N_8050,N_5823);
nor U10227 (N_10227,N_6871,N_7992);
or U10228 (N_10228,N_5164,N_8794);
and U10229 (N_10229,N_7814,N_8779);
nand U10230 (N_10230,N_7435,N_8612);
or U10231 (N_10231,N_6758,N_7545);
or U10232 (N_10232,N_7332,N_8835);
nor U10233 (N_10233,N_9430,N_8599);
nor U10234 (N_10234,N_8636,N_8383);
nor U10235 (N_10235,N_7793,N_7469);
or U10236 (N_10236,N_8472,N_6642);
and U10237 (N_10237,N_8314,N_8839);
nor U10238 (N_10238,N_8056,N_9418);
nor U10239 (N_10239,N_9014,N_6792);
nand U10240 (N_10240,N_8446,N_6268);
and U10241 (N_10241,N_6968,N_7611);
and U10242 (N_10242,N_5026,N_5562);
nand U10243 (N_10243,N_5469,N_9105);
nand U10244 (N_10244,N_5688,N_8593);
nand U10245 (N_10245,N_6904,N_7455);
nand U10246 (N_10246,N_6155,N_9134);
and U10247 (N_10247,N_6825,N_5209);
or U10248 (N_10248,N_7872,N_6446);
xor U10249 (N_10249,N_9799,N_9297);
or U10250 (N_10250,N_5444,N_6838);
nand U10251 (N_10251,N_5604,N_5695);
nor U10252 (N_10252,N_8219,N_9459);
nor U10253 (N_10253,N_8435,N_9057);
and U10254 (N_10254,N_9587,N_7220);
nand U10255 (N_10255,N_6863,N_6767);
and U10256 (N_10256,N_9903,N_7422);
and U10257 (N_10257,N_8724,N_6774);
nor U10258 (N_10258,N_5720,N_6103);
nor U10259 (N_10259,N_5163,N_6017);
nor U10260 (N_10260,N_6243,N_7871);
or U10261 (N_10261,N_5581,N_8589);
nor U10262 (N_10262,N_5673,N_8481);
xor U10263 (N_10263,N_5747,N_8237);
nor U10264 (N_10264,N_5571,N_8273);
nor U10265 (N_10265,N_7050,N_9905);
and U10266 (N_10266,N_9318,N_9258);
nand U10267 (N_10267,N_5093,N_6876);
or U10268 (N_10268,N_5153,N_9764);
and U10269 (N_10269,N_9739,N_6129);
nand U10270 (N_10270,N_5123,N_8546);
nor U10271 (N_10271,N_8806,N_9261);
or U10272 (N_10272,N_9930,N_8302);
and U10273 (N_10273,N_8074,N_5076);
nand U10274 (N_10274,N_8759,N_7848);
nand U10275 (N_10275,N_7244,N_8411);
nor U10276 (N_10276,N_9798,N_5238);
nor U10277 (N_10277,N_9954,N_7662);
and U10278 (N_10278,N_9207,N_8966);
and U10279 (N_10279,N_5596,N_7506);
or U10280 (N_10280,N_7029,N_8763);
and U10281 (N_10281,N_8998,N_9065);
nor U10282 (N_10282,N_9606,N_5352);
and U10283 (N_10283,N_9303,N_7493);
or U10284 (N_10284,N_8540,N_7446);
or U10285 (N_10285,N_7171,N_8270);
or U10286 (N_10286,N_8818,N_9353);
or U10287 (N_10287,N_7855,N_5262);
or U10288 (N_10288,N_7952,N_7920);
nand U10289 (N_10289,N_8017,N_9084);
and U10290 (N_10290,N_9621,N_9041);
nand U10291 (N_10291,N_8180,N_5712);
nand U10292 (N_10292,N_9398,N_8215);
nor U10293 (N_10293,N_5468,N_8316);
nand U10294 (N_10294,N_8325,N_7236);
and U10295 (N_10295,N_8409,N_8967);
nand U10296 (N_10296,N_6941,N_5614);
and U10297 (N_10297,N_9696,N_8029);
and U10298 (N_10298,N_9401,N_9915);
nand U10299 (N_10299,N_5548,N_5804);
and U10300 (N_10300,N_6198,N_6459);
nand U10301 (N_10301,N_5335,N_7106);
nor U10302 (N_10302,N_6857,N_6591);
nor U10303 (N_10303,N_5378,N_9686);
nand U10304 (N_10304,N_8256,N_8602);
or U10305 (N_10305,N_7770,N_7041);
nor U10306 (N_10306,N_7274,N_5139);
nor U10307 (N_10307,N_5689,N_8627);
and U10308 (N_10308,N_6710,N_8847);
and U10309 (N_10309,N_7949,N_5002);
or U10310 (N_10310,N_8394,N_6617);
or U10311 (N_10311,N_5913,N_8156);
nor U10312 (N_10312,N_5960,N_9193);
nand U10313 (N_10313,N_9901,N_9438);
and U10314 (N_10314,N_7644,N_8897);
nor U10315 (N_10315,N_6903,N_7179);
nor U10316 (N_10316,N_8891,N_8576);
and U10317 (N_10317,N_5762,N_5809);
or U10318 (N_10318,N_6240,N_9932);
nand U10319 (N_10319,N_5467,N_7004);
nor U10320 (N_10320,N_9335,N_9540);
and U10321 (N_10321,N_6022,N_5129);
and U10322 (N_10322,N_7276,N_9110);
nand U10323 (N_10323,N_5948,N_9796);
nor U10324 (N_10324,N_7679,N_6842);
nand U10325 (N_10325,N_8875,N_9391);
nor U10326 (N_10326,N_6099,N_7959);
or U10327 (N_10327,N_5326,N_5489);
nand U10328 (N_10328,N_6143,N_8434);
or U10329 (N_10329,N_7118,N_6448);
nor U10330 (N_10330,N_5721,N_5242);
nor U10331 (N_10331,N_7632,N_6047);
nor U10332 (N_10332,N_6490,N_9338);
or U10333 (N_10333,N_9854,N_8982);
or U10334 (N_10334,N_5623,N_6633);
xnor U10335 (N_10335,N_7136,N_9542);
nand U10336 (N_10336,N_5421,N_8805);
nand U10337 (N_10337,N_8114,N_7482);
nor U10338 (N_10338,N_6451,N_8977);
nand U10339 (N_10339,N_9528,N_7129);
and U10340 (N_10340,N_8714,N_5138);
nor U10341 (N_10341,N_5891,N_5815);
or U10342 (N_10342,N_9674,N_5782);
nand U10343 (N_10343,N_8014,N_8213);
nand U10344 (N_10344,N_7604,N_8821);
nor U10345 (N_10345,N_5430,N_5981);
or U10346 (N_10346,N_8804,N_5241);
or U10347 (N_10347,N_7241,N_8807);
nand U10348 (N_10348,N_7240,N_5844);
nand U10349 (N_10349,N_9229,N_7616);
or U10350 (N_10350,N_5535,N_7926);
nand U10351 (N_10351,N_7182,N_7636);
nand U10352 (N_10352,N_7562,N_6440);
and U10353 (N_10353,N_6912,N_5792);
nand U10354 (N_10354,N_9837,N_7551);
or U10355 (N_10355,N_5778,N_7904);
or U10356 (N_10356,N_6565,N_5363);
nand U10357 (N_10357,N_8036,N_5896);
nand U10358 (N_10358,N_8494,N_7116);
and U10359 (N_10359,N_7237,N_7071);
nand U10360 (N_10360,N_6419,N_7897);
and U10361 (N_10361,N_5013,N_9482);
nor U10362 (N_10362,N_9072,N_6219);
nor U10363 (N_10363,N_8082,N_7856);
or U10364 (N_10364,N_9658,N_7159);
and U10365 (N_10365,N_5217,N_5276);
nand U10366 (N_10366,N_7200,N_6044);
nand U10367 (N_10367,N_8669,N_5716);
or U10368 (N_10368,N_9451,N_8947);
nor U10369 (N_10369,N_8769,N_6028);
and U10370 (N_10370,N_9444,N_8427);
and U10371 (N_10371,N_5863,N_8185);
or U10372 (N_10372,N_9044,N_7700);
and U10373 (N_10373,N_8989,N_7067);
and U10374 (N_10374,N_5287,N_9310);
and U10375 (N_10375,N_7630,N_6349);
nand U10376 (N_10376,N_8922,N_7351);
nor U10377 (N_10377,N_6031,N_7498);
or U10378 (N_10378,N_7841,N_7497);
nand U10379 (N_10379,N_5068,N_5785);
or U10380 (N_10380,N_6773,N_6057);
nand U10381 (N_10381,N_5874,N_6036);
and U10382 (N_10382,N_5719,N_7196);
nor U10383 (N_10383,N_9436,N_7246);
nor U10384 (N_10384,N_8103,N_8284);
or U10385 (N_10385,N_5599,N_8957);
nor U10386 (N_10386,N_5432,N_7964);
nand U10387 (N_10387,N_7889,N_9777);
nor U10388 (N_10388,N_8814,N_9983);
and U10389 (N_10389,N_8236,N_9223);
nor U10390 (N_10390,N_9473,N_9973);
nand U10391 (N_10391,N_9855,N_7884);
nor U10392 (N_10392,N_7286,N_6985);
and U10393 (N_10393,N_7378,N_6407);
and U10394 (N_10394,N_9185,N_5984);
nor U10395 (N_10395,N_9230,N_9572);
nor U10396 (N_10396,N_5481,N_8094);
nand U10397 (N_10397,N_9969,N_8978);
or U10398 (N_10398,N_7853,N_8629);
nand U10399 (N_10399,N_5090,N_9765);
or U10400 (N_10400,N_8524,N_5343);
and U10401 (N_10401,N_9649,N_5140);
and U10402 (N_10402,N_9266,N_5300);
or U10403 (N_10403,N_6796,N_6625);
and U10404 (N_10404,N_5005,N_5146);
nand U10405 (N_10405,N_7317,N_7416);
nand U10406 (N_10406,N_9846,N_5664);
nor U10407 (N_10407,N_8376,N_6046);
nor U10408 (N_10408,N_7756,N_6323);
nand U10409 (N_10409,N_6548,N_5670);
nand U10410 (N_10410,N_7935,N_9726);
nor U10411 (N_10411,N_6503,N_5846);
nand U10412 (N_10412,N_6203,N_8490);
or U10413 (N_10413,N_6746,N_6977);
or U10414 (N_10414,N_8951,N_6001);
or U10415 (N_10415,N_6788,N_8568);
or U10416 (N_10416,N_8838,N_5166);
nor U10417 (N_10417,N_9348,N_8865);
nor U10418 (N_10418,N_6034,N_6489);
nand U10419 (N_10419,N_9937,N_5254);
nor U10420 (N_10420,N_6664,N_7701);
or U10421 (N_10421,N_8475,N_6672);
nand U10422 (N_10422,N_5675,N_9895);
and U10423 (N_10423,N_7420,N_7365);
or U10424 (N_10424,N_9491,N_8419);
or U10425 (N_10425,N_8730,N_8414);
nor U10426 (N_10426,N_8335,N_7725);
and U10427 (N_10427,N_8381,N_7507);
or U10428 (N_10428,N_7778,N_8461);
or U10429 (N_10429,N_6884,N_5910);
nor U10430 (N_10430,N_6145,N_6347);
nand U10431 (N_10431,N_9204,N_6689);
nor U10432 (N_10432,N_7253,N_9908);
nor U10433 (N_10433,N_9881,N_9989);
nor U10434 (N_10434,N_8406,N_6623);
and U10435 (N_10435,N_9472,N_6937);
and U10436 (N_10436,N_6694,N_9637);
nor U10437 (N_10437,N_8007,N_7127);
and U10438 (N_10438,N_9113,N_7873);
or U10439 (N_10439,N_6624,N_8953);
or U10440 (N_10440,N_5890,N_6174);
nand U10441 (N_10441,N_9456,N_5484);
nand U10442 (N_10442,N_8995,N_8668);
nor U10443 (N_10443,N_9870,N_9966);
or U10444 (N_10444,N_8143,N_6976);
xor U10445 (N_10445,N_7262,N_9646);
and U10446 (N_10446,N_5820,N_6606);
nor U10447 (N_10447,N_8869,N_9529);
and U10448 (N_10448,N_6110,N_7819);
nand U10449 (N_10449,N_8923,N_8748);
or U10450 (N_10450,N_7030,N_9087);
and U10451 (N_10451,N_8948,N_9679);
nor U10452 (N_10452,N_5205,N_9510);
or U10453 (N_10453,N_6194,N_5892);
or U10454 (N_10454,N_9508,N_5190);
or U10455 (N_10455,N_5808,N_5367);
or U10456 (N_10456,N_8772,N_6326);
or U10457 (N_10457,N_9030,N_5381);
nor U10458 (N_10458,N_5176,N_6290);
or U10459 (N_10459,N_9620,N_8578);
or U10460 (N_10460,N_9153,N_5185);
nand U10461 (N_10461,N_9527,N_7445);
nor U10462 (N_10462,N_9801,N_5014);
nor U10463 (N_10463,N_9887,N_7359);
nor U10464 (N_10464,N_9086,N_8770);
and U10465 (N_10465,N_8912,N_5046);
and U10466 (N_10466,N_7668,N_8898);
or U10467 (N_10467,N_9863,N_9467);
xnor U10468 (N_10468,N_5953,N_7750);
nand U10469 (N_10469,N_7340,N_6576);
nand U10470 (N_10470,N_9623,N_8893);
and U10471 (N_10471,N_8605,N_6896);
or U10472 (N_10472,N_9574,N_7014);
or U10473 (N_10473,N_9164,N_9250);
nand U10474 (N_10474,N_9374,N_5626);
nand U10475 (N_10475,N_8555,N_7865);
or U10476 (N_10476,N_5832,N_7798);
or U10477 (N_10477,N_6802,N_8452);
nand U10478 (N_10478,N_9075,N_9283);
or U10479 (N_10479,N_7031,N_6289);
or U10480 (N_10480,N_9483,N_5344);
or U10481 (N_10481,N_9060,N_9982);
nand U10482 (N_10482,N_9971,N_9036);
and U10483 (N_10483,N_7516,N_8186);
and U10484 (N_10484,N_6461,N_9329);
or U10485 (N_10485,N_9596,N_6195);
and U10486 (N_10486,N_8148,N_7462);
nor U10487 (N_10487,N_5992,N_6596);
nand U10488 (N_10488,N_5572,N_7732);
or U10489 (N_10489,N_9144,N_7056);
and U10490 (N_10490,N_8417,N_9156);
nand U10491 (N_10491,N_7826,N_5196);
nor U10492 (N_10492,N_9647,N_5817);
nand U10493 (N_10493,N_9427,N_6920);
nor U10494 (N_10494,N_7447,N_8361);
and U10495 (N_10495,N_7448,N_9909);
nand U10496 (N_10496,N_7419,N_5831);
nor U10497 (N_10497,N_8920,N_6220);
and U10498 (N_10498,N_7204,N_8644);
nand U10499 (N_10499,N_6978,N_5578);
or U10500 (N_10500,N_9298,N_8377);
or U10501 (N_10501,N_7037,N_8971);
and U10502 (N_10502,N_7361,N_6256);
nand U10503 (N_10503,N_5950,N_5234);
or U10504 (N_10504,N_8582,N_8707);
or U10505 (N_10505,N_5443,N_5684);
and U10506 (N_10506,N_8516,N_7170);
xor U10507 (N_10507,N_7527,N_5613);
and U10508 (N_10508,N_6432,N_8802);
nand U10509 (N_10509,N_9974,N_5298);
and U10510 (N_10510,N_5022,N_7615);
and U10511 (N_10511,N_5516,N_6481);
or U10512 (N_10512,N_5925,N_9154);
nor U10513 (N_10513,N_6467,N_7519);
nor U10514 (N_10514,N_8333,N_8771);
or U10515 (N_10515,N_8911,N_6634);
or U10516 (N_10516,N_7741,N_8130);
and U10517 (N_10517,N_7626,N_5265);
or U10518 (N_10518,N_5994,N_7869);
nand U10519 (N_10519,N_5324,N_6865);
and U10520 (N_10520,N_8501,N_8491);
and U10521 (N_10521,N_8689,N_9019);
nand U10522 (N_10522,N_6890,N_9565);
nor U10523 (N_10523,N_5244,N_8640);
or U10524 (N_10524,N_7484,N_6726);
and U10525 (N_10525,N_9956,N_5079);
nor U10526 (N_10526,N_6783,N_7186);
or U10527 (N_10527,N_9062,N_5836);
nor U10528 (N_10528,N_7603,N_8363);
or U10529 (N_10529,N_6898,N_5240);
and U10530 (N_10530,N_8557,N_8566);
or U10531 (N_10531,N_9997,N_7138);
and U10532 (N_10532,N_5373,N_5437);
nor U10533 (N_10533,N_6334,N_7021);
nand U10534 (N_10534,N_6635,N_7764);
nand U10535 (N_10535,N_7923,N_5212);
or U10536 (N_10536,N_9747,N_7088);
nand U10537 (N_10537,N_9366,N_8474);
nand U10538 (N_10538,N_8125,N_6641);
and U10539 (N_10539,N_6237,N_7428);
and U10540 (N_10540,N_7181,N_6423);
nor U10541 (N_10541,N_6539,N_5877);
and U10542 (N_10542,N_6435,N_8931);
or U10543 (N_10543,N_6752,N_6441);
and U10544 (N_10544,N_8182,N_8418);
nand U10545 (N_10545,N_8686,N_7830);
and U10546 (N_10546,N_5737,N_5397);
or U10547 (N_10547,N_5498,N_8705);
nor U10548 (N_10548,N_5744,N_6284);
nand U10549 (N_10549,N_9784,N_9912);
nand U10550 (N_10550,N_5306,N_5206);
nand U10551 (N_10551,N_7168,N_9002);
nor U10552 (N_10552,N_5342,N_5725);
nand U10553 (N_10553,N_8595,N_7621);
nand U10554 (N_10554,N_7628,N_8448);
and U10555 (N_10555,N_6914,N_7887);
or U10556 (N_10556,N_6652,N_6841);
or U10557 (N_10557,N_7032,N_8696);
nor U10558 (N_10558,N_7674,N_9094);
and U10559 (N_10559,N_7973,N_5311);
or U10560 (N_10560,N_6510,N_6135);
and U10561 (N_10561,N_6798,N_6056);
or U10562 (N_10562,N_9886,N_9669);
and U10563 (N_10563,N_7149,N_7944);
nand U10564 (N_10564,N_7514,N_8997);
and U10565 (N_10565,N_7569,N_8098);
nor U10566 (N_10566,N_5471,N_5134);
nor U10567 (N_10567,N_5813,N_5094);
nor U10568 (N_10568,N_8010,N_7999);
and U10569 (N_10569,N_7091,N_5488);
or U10570 (N_10570,N_9992,N_8463);
nand U10571 (N_10571,N_6088,N_8809);
nor U10572 (N_10572,N_7161,N_7036);
or U10573 (N_10573,N_6728,N_6229);
or U10574 (N_10574,N_5680,N_6425);
nor U10575 (N_10575,N_9560,N_9439);
or U10576 (N_10576,N_6897,N_7460);
and U10577 (N_10577,N_5930,N_5105);
and U10578 (N_10578,N_6156,N_6454);
nor U10579 (N_10579,N_9513,N_7916);
and U10580 (N_10580,N_5061,N_8153);
nand U10581 (N_10581,N_9936,N_5407);
and U10582 (N_10582,N_9820,N_9638);
and U10583 (N_10583,N_9766,N_9904);
nand U10584 (N_10584,N_9720,N_9729);
and U10585 (N_10585,N_7857,N_6913);
or U10586 (N_10586,N_7694,N_5587);
nand U10587 (N_10587,N_5947,N_5222);
nor U10588 (N_10588,N_9512,N_7151);
nand U10589 (N_10589,N_5893,N_6807);
nand U10590 (N_10590,N_5946,N_5682);
nor U10591 (N_10591,N_5310,N_8154);
or U10592 (N_10592,N_9770,N_5758);
xnor U10593 (N_10593,N_9640,N_6476);
or U10594 (N_10594,N_7677,N_8556);
or U10595 (N_10595,N_7976,N_7859);
or U10596 (N_10596,N_8639,N_6202);
and U10597 (N_10597,N_6866,N_5401);
nor U10598 (N_10598,N_6558,N_9493);
and U10599 (N_10599,N_8051,N_8832);
nand U10600 (N_10600,N_9024,N_6619);
nand U10601 (N_10601,N_7675,N_8736);
nor U10602 (N_10602,N_7062,N_5267);
or U10603 (N_10603,N_6361,N_7896);
nand U10604 (N_10604,N_9921,N_7242);
nand U10605 (N_10605,N_9441,N_7825);
nor U10606 (N_10606,N_5171,N_9927);
nor U10607 (N_10607,N_8173,N_9496);
or U10608 (N_10608,N_9414,N_8565);
nand U10609 (N_10609,N_9249,N_8458);
or U10610 (N_10610,N_7321,N_9146);
nand U10611 (N_10611,N_9688,N_6337);
xor U10612 (N_10612,N_9949,N_6621);
nand U10613 (N_10613,N_6816,N_5081);
nand U10614 (N_10614,N_7073,N_5431);
or U10615 (N_10615,N_8872,N_9745);
nor U10616 (N_10616,N_6131,N_9751);
or U10617 (N_10617,N_5642,N_9511);
or U10618 (N_10618,N_5207,N_6536);
nor U10619 (N_10619,N_9306,N_6882);
or U10620 (N_10620,N_6566,N_5483);
nand U10621 (N_10621,N_6943,N_9385);
nand U10622 (N_10622,N_9771,N_6847);
nor U10623 (N_10623,N_6869,N_8963);
nor U10624 (N_10624,N_9322,N_8601);
or U10625 (N_10625,N_8853,N_8290);
nor U10626 (N_10626,N_7297,N_6545);
nand U10627 (N_10627,N_6919,N_6703);
nand U10628 (N_10628,N_6452,N_9237);
nand U10629 (N_10629,N_7157,N_5534);
nand U10630 (N_10630,N_7265,N_7433);
nand U10631 (N_10631,N_8657,N_8773);
or U10632 (N_10632,N_6270,N_6860);
and U10633 (N_10633,N_6128,N_7354);
nor U10634 (N_10634,N_7468,N_9953);
nand U10635 (N_10635,N_9842,N_8856);
or U10636 (N_10636,N_7561,N_5656);
or U10637 (N_10637,N_7198,N_5531);
or U10638 (N_10638,N_8559,N_7761);
or U10639 (N_10639,N_7748,N_5755);
nand U10640 (N_10640,N_7704,N_5568);
nand U10641 (N_10641,N_6894,N_5962);
nor U10642 (N_10642,N_6813,N_6382);
and U10643 (N_10643,N_8144,N_7119);
nand U10644 (N_10644,N_7844,N_5221);
and U10645 (N_10645,N_9774,N_8132);
nand U10646 (N_10646,N_9651,N_6048);
and U10647 (N_10647,N_5441,N_6158);
nor U10648 (N_10648,N_6947,N_5606);
or U10649 (N_10649,N_8507,N_5769);
nor U10650 (N_10650,N_9682,N_7914);
or U10651 (N_10651,N_7651,N_8525);
nor U10652 (N_10652,N_5850,N_5628);
and U10653 (N_10653,N_9337,N_5091);
and U10654 (N_10654,N_9240,N_9505);
nor U10655 (N_10655,N_7235,N_7135);
nor U10656 (N_10656,N_7864,N_7957);
and U10657 (N_10657,N_8563,N_7554);
nand U10658 (N_10658,N_8579,N_6563);
nor U10659 (N_10659,N_6580,N_6445);
nor U10660 (N_10660,N_5155,N_9319);
nor U10661 (N_10661,N_6346,N_8685);
and U10662 (N_10662,N_7622,N_6385);
and U10663 (N_10663,N_7248,N_5971);
nor U10664 (N_10664,N_8798,N_7698);
and U10665 (N_10665,N_8577,N_8945);
nand U10666 (N_10666,N_5411,N_9762);
and U10667 (N_10667,N_7617,N_8005);
nand U10668 (N_10668,N_9914,N_6329);
or U10669 (N_10669,N_6845,N_7110);
nor U10670 (N_10670,N_6995,N_5500);
or U10671 (N_10671,N_5440,N_9563);
nand U10672 (N_10672,N_5997,N_5511);
and U10673 (N_10673,N_6991,N_5218);
and U10674 (N_10674,N_5837,N_6089);
or U10675 (N_10675,N_8471,N_7891);
nor U10676 (N_10676,N_8710,N_8537);
and U10677 (N_10677,N_8184,N_7444);
nor U10678 (N_10678,N_8788,N_8313);
nor U10679 (N_10679,N_5192,N_9461);
nand U10680 (N_10680,N_6214,N_7529);
or U10681 (N_10681,N_9216,N_7017);
and U10682 (N_10682,N_6938,N_6930);
and U10683 (N_10683,N_6105,N_5036);
nor U10684 (N_10684,N_9326,N_9735);
or U10685 (N_10685,N_7356,N_7152);
xor U10686 (N_10686,N_8254,N_8039);
nand U10687 (N_10687,N_7578,N_9964);
and U10688 (N_10688,N_6148,N_6660);
or U10689 (N_10689,N_9465,N_6970);
and U10690 (N_10690,N_6682,N_6861);
nand U10691 (N_10691,N_6921,N_8280);
and U10692 (N_10692,N_9034,N_5566);
or U10693 (N_10693,N_7103,N_9222);
and U10694 (N_10694,N_7531,N_8080);
nor U10695 (N_10695,N_7918,N_6872);
or U10696 (N_10696,N_8431,N_9405);
nand U10697 (N_10697,N_9161,N_8432);
and U10698 (N_10698,N_8206,N_7404);
or U10699 (N_10699,N_8066,N_6493);
and U10700 (N_10700,N_5619,N_6303);
or U10701 (N_10701,N_5003,N_9447);
and U10702 (N_10702,N_7839,N_9287);
or U10703 (N_10703,N_8999,N_8792);
and U10704 (N_10704,N_9043,N_8239);
or U10705 (N_10705,N_8514,N_6724);
nor U10706 (N_10706,N_8919,N_6404);
nand U10707 (N_10707,N_6950,N_9020);
and U10708 (N_10708,N_5726,N_7768);
nand U10709 (N_10709,N_9420,N_7387);
nand U10710 (N_10710,N_9781,N_9083);
or U10711 (N_10711,N_8868,N_6043);
and U10712 (N_10712,N_5314,N_5384);
and U10713 (N_10713,N_5025,N_5410);
nor U10714 (N_10714,N_5446,N_6644);
nand U10715 (N_10715,N_8894,N_8217);
and U10716 (N_10716,N_9008,N_7678);
nand U10717 (N_10717,N_7817,N_7965);
or U10718 (N_10718,N_7215,N_8161);
or U10719 (N_10719,N_7666,N_9892);
nor U10720 (N_10720,N_9470,N_5882);
and U10721 (N_10721,N_7010,N_7431);
and U10722 (N_10722,N_6379,N_8726);
nand U10723 (N_10723,N_7209,N_8739);
and U10724 (N_10724,N_6294,N_6000);
nand U10725 (N_10725,N_7641,N_7372);
nor U10726 (N_10726,N_5388,N_6277);
and U10727 (N_10727,N_9271,N_6893);
nor U10728 (N_10728,N_7495,N_9931);
and U10729 (N_10729,N_7130,N_9056);
nand U10730 (N_10730,N_8881,N_9290);
nand U10731 (N_10731,N_5657,N_8562);
nor U10732 (N_10732,N_6529,N_6377);
and U10733 (N_10733,N_6090,N_8349);
nor U10734 (N_10734,N_7477,N_7650);
or U10735 (N_10735,N_9705,N_7524);
or U10736 (N_10736,N_9289,N_5603);
and U10737 (N_10737,N_6469,N_6479);
nand U10738 (N_10738,N_7227,N_6915);
or U10739 (N_10739,N_6933,N_9443);
nor U10740 (N_10740,N_6052,N_9486);
or U10741 (N_10741,N_6456,N_6810);
and U10742 (N_10742,N_9497,N_5909);
or U10743 (N_10743,N_9951,N_6532);
or U10744 (N_10744,N_9730,N_8574);
and U10745 (N_10745,N_8397,N_6971);
and U10746 (N_10746,N_7095,N_6114);
or U10747 (N_10747,N_6534,N_5677);
nor U10748 (N_10748,N_7185,N_9526);
and U10749 (N_10749,N_7908,N_8768);
or U10750 (N_10750,N_7408,N_5773);
or U10751 (N_10751,N_5172,N_7867);
nor U10752 (N_10752,N_9716,N_9588);
nand U10753 (N_10753,N_6698,N_7858);
and U10754 (N_10754,N_5070,N_9981);
or U10755 (N_10755,N_7988,N_8296);
nand U10756 (N_10756,N_7513,N_7229);
or U10757 (N_10757,N_9754,N_5830);
or U10758 (N_10758,N_9760,N_6239);
nor U10759 (N_10759,N_9876,N_9742);
and U10760 (N_10760,N_6170,N_9013);
nand U10761 (N_10761,N_9147,N_6839);
or U10762 (N_10762,N_8015,N_6507);
nand U10763 (N_10763,N_8522,N_7530);
nor U10764 (N_10764,N_6782,N_5293);
or U10765 (N_10765,N_6180,N_7499);
and U10766 (N_10766,N_8060,N_8231);
nor U10767 (N_10767,N_5527,N_5433);
nor U10768 (N_10768,N_5279,N_8366);
nor U10769 (N_10769,N_5510,N_9174);
or U10770 (N_10770,N_9986,N_6965);
or U10771 (N_10771,N_5876,N_8831);
nor U10772 (N_10772,N_8253,N_5842);
nand U10773 (N_10773,N_7542,N_5513);
or U10774 (N_10774,N_7279,N_6702);
and U10775 (N_10775,N_8766,N_6852);
and U10776 (N_10776,N_7003,N_5739);
nand U10777 (N_10777,N_9365,N_5940);
and U10778 (N_10778,N_6380,N_6053);
nor U10779 (N_10779,N_8679,N_9758);
nand U10780 (N_10780,N_6958,N_5256);
nand U10781 (N_10781,N_7989,N_8140);
and U10782 (N_10782,N_9312,N_8939);
nor U10783 (N_10783,N_9814,N_6609);
nand U10784 (N_10784,N_8212,N_6620);
nand U10785 (N_10785,N_8407,N_6265);
or U10786 (N_10786,N_8552,N_6260);
nor U10787 (N_10787,N_8896,N_7600);
and U10788 (N_10788,N_6982,N_6486);
xnor U10789 (N_10789,N_8509,N_6508);
or U10790 (N_10790,N_7697,N_9740);
nor U10791 (N_10791,N_8495,N_5525);
or U10792 (N_10792,N_7609,N_9159);
and U10793 (N_10793,N_8965,N_9534);
and U10794 (N_10794,N_5136,N_8757);
and U10795 (N_10795,N_7137,N_5301);
nand U10796 (N_10796,N_6276,N_8393);
nand U10797 (N_10797,N_9979,N_7192);
nand U10798 (N_10798,N_7048,N_5715);
and U10799 (N_10799,N_7661,N_6827);
or U10800 (N_10800,N_8127,N_6926);
nand U10801 (N_10801,N_9732,N_9450);
or U10802 (N_10802,N_7925,N_5509);
or U10803 (N_10803,N_5683,N_9737);
nand U10804 (N_10804,N_5261,N_7070);
xnor U10805 (N_10805,N_7098,N_6556);
and U10806 (N_10806,N_9967,N_8070);
nor U10807 (N_10807,N_6515,N_5740);
nand U10808 (N_10808,N_9152,N_5391);
or U10809 (N_10809,N_6647,N_7188);
or U10810 (N_10810,N_8972,N_5520);
nor U10811 (N_10811,N_9101,N_5907);
and U10812 (N_10812,N_9819,N_5624);
and U10813 (N_10813,N_5973,N_8241);
nor U10814 (N_10814,N_9616,N_8147);
or U10815 (N_10815,N_8178,N_6434);
or U10816 (N_10816,N_5278,N_5029);
and U10817 (N_10817,N_9680,N_8041);
and U10818 (N_10818,N_8548,N_9656);
or U10819 (N_10819,N_8207,N_9040);
or U10820 (N_10820,N_6524,N_8528);
or U10821 (N_10821,N_9484,N_5149);
nand U10822 (N_10822,N_6674,N_5235);
xnor U10823 (N_10823,N_6453,N_6206);
nor U10824 (N_10824,N_8653,N_7703);
or U10825 (N_10825,N_7319,N_9049);
nand U10826 (N_10826,N_5540,N_9292);
nor U10827 (N_10827,N_9664,N_8892);
nand U10828 (N_10828,N_8672,N_8033);
and U10829 (N_10829,N_6874,N_8177);
and U10830 (N_10830,N_7536,N_6139);
nand U10831 (N_10831,N_5386,N_6756);
or U10832 (N_10832,N_9531,N_9453);
nor U10833 (N_10833,N_7288,N_8392);
and U10834 (N_10834,N_7089,N_6482);
nor U10835 (N_10835,N_7485,N_9933);
or U10836 (N_10836,N_5110,N_5330);
nand U10837 (N_10837,N_9054,N_5523);
and U10838 (N_10838,N_8293,N_6669);
nor U10839 (N_10839,N_5763,N_7458);
nand U10840 (N_10840,N_6643,N_9145);
or U10841 (N_10841,N_9278,N_5044);
and U10842 (N_10842,N_6318,N_6426);
nor U10843 (N_10843,N_8227,N_5887);
or U10844 (N_10844,N_9380,N_7932);
nand U10845 (N_10845,N_9607,N_6690);
nor U10846 (N_10846,N_8697,N_9082);
or U10847 (N_10847,N_7597,N_9323);
nand U10848 (N_10848,N_7252,N_5576);
nor U10849 (N_10849,N_8122,N_7163);
and U10850 (N_10850,N_8785,N_6447);
nand U10851 (N_10851,N_5042,N_7362);
and U10852 (N_10852,N_8046,N_5600);
or U10853 (N_10853,N_8251,N_6822);
nor U10854 (N_10854,N_6498,N_5366);
or U10855 (N_10855,N_7822,N_6648);
nand U10856 (N_10856,N_6060,N_8663);
nor U10857 (N_10857,N_8334,N_8974);
and U10858 (N_10858,N_7540,N_8307);
nand U10859 (N_10859,N_8425,N_7441);
nand U10860 (N_10860,N_7556,N_7967);
nand U10861 (N_10861,N_7072,N_7075);
nand U10862 (N_10862,N_7984,N_8203);
nor U10863 (N_10863,N_9115,N_9217);
or U10864 (N_10864,N_9099,N_7180);
or U10865 (N_10865,N_9723,N_7892);
or U10866 (N_10866,N_7719,N_8848);
and U10867 (N_10867,N_9202,N_8533);
nand U10868 (N_10868,N_8271,N_8312);
nor U10869 (N_10869,N_8128,N_7324);
nand U10870 (N_10870,N_6348,N_9603);
and U10871 (N_10871,N_6468,N_5435);
and U10872 (N_10872,N_9839,N_6923);
and U10873 (N_10873,N_9634,N_8479);
and U10874 (N_10874,N_6928,N_8071);
nor U10875 (N_10875,N_9288,N_7285);
or U10876 (N_10876,N_6147,N_8718);
or U10877 (N_10877,N_7049,N_5644);
or U10878 (N_10878,N_9996,N_8592);
xnor U10879 (N_10879,N_5237,N_7683);
and U10880 (N_10880,N_7566,N_8646);
nand U10881 (N_10881,N_9333,N_6394);
and U10882 (N_10882,N_9759,N_7721);
or U10883 (N_10883,N_6312,N_6662);
or U10884 (N_10884,N_8580,N_7707);
nand U10885 (N_10885,N_7909,N_5412);
nand U10886 (N_10886,N_9016,N_6497);
or U10887 (N_10887,N_9180,N_9350);
or U10888 (N_10888,N_7389,N_9466);
nor U10889 (N_10889,N_6330,N_9140);
or U10890 (N_10890,N_5771,N_8703);
nor U10891 (N_10891,N_7791,N_8077);
nor U10892 (N_10892,N_6172,N_8338);
or U10893 (N_10893,N_8901,N_5584);
nor U10894 (N_10894,N_6972,N_5383);
and U10895 (N_10895,N_7197,N_8133);
and U10896 (N_10896,N_5297,N_9753);
or U10897 (N_10897,N_7878,N_8091);
nand U10898 (N_10898,N_9373,N_6327);
nor U10899 (N_10899,N_9413,N_6014);
or U10900 (N_10900,N_9309,N_5069);
nand U10901 (N_10901,N_6697,N_5341);
and U10902 (N_10902,N_7974,N_7942);
nand U10903 (N_10903,N_9815,N_6901);
nor U10904 (N_10904,N_8364,N_6413);
or U10905 (N_10905,N_9661,N_5080);
nor U10906 (N_10906,N_9021,N_7099);
nor U10907 (N_10907,N_5952,N_7490);
and U10908 (N_10908,N_9006,N_9500);
and U10909 (N_10909,N_6679,N_8331);
nor U10910 (N_10910,N_5794,N_6929);
and U10911 (N_10911,N_7403,N_9896);
nand U10912 (N_10912,N_6012,N_9871);
and U10913 (N_10913,N_8249,N_6585);
and U10914 (N_10914,N_6781,N_9314);
nor U10915 (N_10915,N_6168,N_7449);
nand U10916 (N_10916,N_8908,N_6877);
and U10917 (N_10917,N_7218,N_5805);
nand U10918 (N_10918,N_9235,N_5037);
nand U10919 (N_10919,N_5004,N_5504);
nand U10920 (N_10920,N_6487,N_6613);
nor U10921 (N_10921,N_9582,N_5208);
nor U10922 (N_10922,N_9717,N_8606);
nor U10923 (N_10923,N_7728,N_6123);
or U10924 (N_10924,N_6024,N_7584);
nand U10925 (N_10925,N_8250,N_5018);
or U10926 (N_10926,N_7809,N_7705);
nor U10927 (N_10927,N_9399,N_9210);
and U10928 (N_10928,N_8341,N_8609);
and U10929 (N_10929,N_8700,N_8052);
nand U10930 (N_10930,N_8786,N_9813);
nor U10931 (N_10931,N_5563,N_7549);
and U10932 (N_10932,N_9190,N_5795);
nor U10933 (N_10933,N_9631,N_5008);
nor U10934 (N_10934,N_8008,N_5040);
or U10935 (N_10935,N_5434,N_9356);
and U10936 (N_10936,N_9962,N_9609);
nor U10937 (N_10937,N_7291,N_8918);
nor U10938 (N_10938,N_9721,N_9703);
nor U10939 (N_10939,N_5585,N_5506);
and U10940 (N_10940,N_8155,N_8024);
or U10941 (N_10941,N_7111,N_6603);
and U10942 (N_10942,N_8720,N_8174);
nor U10943 (N_10943,N_8157,N_8753);
and U10944 (N_10944,N_8887,N_5917);
or U10945 (N_10945,N_8022,N_7026);
nor U10946 (N_10946,N_7105,N_6688);
or U10947 (N_10947,N_6800,N_7802);
nand U10948 (N_10948,N_5601,N_9919);
nor U10949 (N_10949,N_9591,N_8829);
or U10950 (N_10950,N_5757,N_9736);
nand U10951 (N_10951,N_6526,N_7076);
nand U10952 (N_10952,N_9004,N_6814);
or U10953 (N_10953,N_6909,N_5055);
nand U10954 (N_10954,N_9693,N_7983);
nand U10955 (N_10955,N_6122,N_9509);
or U10956 (N_10956,N_8564,N_8422);
or U10957 (N_10957,N_9794,N_5425);
and U10958 (N_10958,N_6295,N_8188);
nor U10959 (N_10959,N_8412,N_6436);
nor U10960 (N_10960,N_6210,N_5708);
nand U10961 (N_10961,N_8863,N_8973);
or U10962 (N_10962,N_9127,N_8761);
nor U10963 (N_10963,N_8444,N_5418);
or U10964 (N_10964,N_8480,N_8867);
nor U10965 (N_10965,N_7147,N_9923);
nand U10966 (N_10966,N_6104,N_8614);
and U10967 (N_10967,N_7012,N_6175);
xor U10968 (N_10968,N_9942,N_6291);
nor U10969 (N_10969,N_6742,N_9786);
and U10970 (N_10970,N_7552,N_6070);
or U10971 (N_10971,N_6341,N_5098);
nand U10972 (N_10972,N_9543,N_8650);
and U10973 (N_10973,N_5372,N_7082);
nor U10974 (N_10974,N_5741,N_6981);
nand U10975 (N_10975,N_8882,N_5210);
nand U10976 (N_10976,N_5270,N_9570);
and U10977 (N_10977,N_8289,N_7505);
nor U10978 (N_10978,N_6398,N_6572);
and U10979 (N_10979,N_5693,N_9536);
nor U10980 (N_10980,N_8375,N_9088);
xnor U10981 (N_10981,N_8671,N_9061);
and U10982 (N_10982,N_5120,N_8190);
or U10983 (N_10983,N_7807,N_9789);
and U10984 (N_10984,N_5978,N_6338);
or U10985 (N_10985,N_7927,N_7199);
nand U10986 (N_10986,N_8141,N_6235);
nor U10987 (N_10987,N_7665,N_8252);
nor U10988 (N_10988,N_8722,N_8379);
and U10989 (N_10989,N_7480,N_7125);
nand U10990 (N_10990,N_6911,N_7762);
or U10991 (N_10991,N_9691,N_5824);
nand U10992 (N_10992,N_8129,N_5570);
nand U10993 (N_10993,N_6589,N_6424);
nand U10994 (N_10994,N_8961,N_6478);
and U10995 (N_10995,N_9275,N_6078);
and U10996 (N_10996,N_9827,N_7875);
nand U10997 (N_10997,N_7953,N_5796);
or U10998 (N_10998,N_6107,N_6450);
nor U10999 (N_10999,N_5888,N_5491);
and U11000 (N_11000,N_9346,N_5580);
or U11001 (N_11001,N_8658,N_5900);
nand U11002 (N_11002,N_6559,N_6948);
or U11003 (N_11003,N_7605,N_9257);
and U11004 (N_11004,N_9807,N_8876);
nor U11005 (N_11005,N_5296,N_6513);
and U11006 (N_11006,N_6120,N_5283);
nand U11007 (N_11007,N_7275,N_8484);
nand U11008 (N_11008,N_5508,N_7154);
nor U11009 (N_11009,N_8398,N_9198);
or U11010 (N_11010,N_7919,N_9652);
and U11011 (N_11011,N_5518,N_7415);
nor U11012 (N_11012,N_8899,N_7272);
nand U11013 (N_11013,N_7555,N_7623);
nand U11014 (N_11014,N_9699,N_7371);
or U11015 (N_11015,N_5223,N_7820);
or U11016 (N_11016,N_6150,N_6846);
or U11017 (N_11017,N_5260,N_8045);
or U11018 (N_11018,N_9943,N_8023);
or U11019 (N_11019,N_7020,N_8996);
and U11020 (N_11020,N_8674,N_7479);
or U11021 (N_11021,N_8142,N_5396);
or U11022 (N_11022,N_6027,N_8279);
nand U11023 (N_11023,N_7148,N_8087);
nand U11024 (N_11024,N_9728,N_9492);
or U11025 (N_11025,N_8021,N_6765);
or U11026 (N_11026,N_7466,N_6444);
nor U11027 (N_11027,N_5165,N_9518);
and U11028 (N_11028,N_7938,N_6065);
nor U11029 (N_11029,N_5655,N_5049);
and U11030 (N_11030,N_9768,N_8288);
nand U11031 (N_11031,N_6266,N_9628);
or U11032 (N_11032,N_7131,N_6274);
or U11033 (N_11033,N_9433,N_8354);
and U11034 (N_11034,N_5427,N_6908);
nand U11035 (N_11035,N_8618,N_9595);
nand U11036 (N_11036,N_5203,N_7723);
nor U11037 (N_11037,N_7876,N_8731);
nor U11038 (N_11038,N_9970,N_9090);
nor U11039 (N_11039,N_7108,N_5938);
or U11040 (N_11040,N_5183,N_9645);
nor U11041 (N_11041,N_5100,N_5975);
nand U11042 (N_11042,N_9719,N_7912);
and U11043 (N_11043,N_6892,N_5899);
or U11044 (N_11044,N_5866,N_5686);
nand U11045 (N_11045,N_9053,N_8581);
or U11046 (N_11046,N_7360,N_8789);
or U11047 (N_11047,N_5723,N_8265);
nand U11048 (N_11048,N_8264,N_5115);
and U11049 (N_11049,N_5197,N_9415);
nand U11050 (N_11050,N_5921,N_7109);
nor U11051 (N_11051,N_5275,N_5825);
or U11052 (N_11052,N_8877,N_8780);
or U11053 (N_11053,N_9868,N_9733);
nand U11054 (N_11054,N_6632,N_5672);
nor U11055 (N_11055,N_6661,N_7642);
or U11056 (N_11056,N_9256,N_6646);
or U11057 (N_11057,N_6883,N_7251);
or U11058 (N_11058,N_8930,N_7146);
or U11059 (N_11059,N_9449,N_8194);
nand U11060 (N_11060,N_8704,N_8727);
or U11061 (N_11061,N_5593,N_9128);
nand U11062 (N_11062,N_9829,N_9957);
or U11063 (N_11063,N_5886,N_6169);
and U11064 (N_11064,N_6557,N_7243);
and U11065 (N_11065,N_7541,N_6074);
or U11066 (N_11066,N_8043,N_7258);
or U11067 (N_11067,N_8047,N_8096);
nand U11068 (N_11068,N_9878,N_5728);
and U11069 (N_11069,N_6954,N_9778);
nand U11070 (N_11070,N_5592,N_5493);
or U11071 (N_11071,N_9547,N_8449);
nor U11072 (N_11072,N_7624,N_5787);
nor U11073 (N_11073,N_9233,N_5405);
or U11074 (N_11074,N_8767,N_8607);
nand U11075 (N_11075,N_9452,N_8652);
nand U11076 (N_11076,N_9775,N_8624);
nor U11077 (N_11077,N_6795,N_5920);
or U11078 (N_11078,N_6313,N_5116);
and U11079 (N_11079,N_8684,N_8196);
nand U11080 (N_11080,N_5699,N_9748);
or U11081 (N_11081,N_8958,N_9553);
xor U11082 (N_11082,N_5194,N_7888);
nor U11083 (N_11083,N_7586,N_9121);
xor U11084 (N_11084,N_7538,N_8214);
or U11085 (N_11085,N_9402,N_6768);
nor U11086 (N_11086,N_8990,N_5395);
nor U11087 (N_11087,N_8634,N_6736);
and U11088 (N_11088,N_8886,N_7599);
nand U11089 (N_11089,N_9063,N_5894);
nand U11090 (N_11090,N_7879,N_6124);
nor U11091 (N_11091,N_7934,N_7755);
nor U11092 (N_11092,N_6083,N_5860);
nor U11093 (N_11093,N_8390,N_9435);
or U11094 (N_11094,N_7504,N_7443);
xnor U11095 (N_11095,N_5322,N_6851);
and U11096 (N_11096,N_8750,N_8344);
or U11097 (N_11097,N_9769,N_7144);
or U11098 (N_11098,N_6732,N_6595);
and U11099 (N_11099,N_9752,N_8347);
and U11100 (N_11100,N_5536,N_9003);
or U11101 (N_11101,N_6520,N_7384);
xnor U11102 (N_11102,N_8849,N_5362);
nor U11103 (N_11103,N_7045,N_6830);
or U11104 (N_11104,N_5895,N_9648);
or U11105 (N_11105,N_8917,N_9522);
and U11106 (N_11106,N_8625,N_6961);
xnor U11107 (N_11107,N_5109,N_6258);
and U11108 (N_11108,N_9469,N_7758);
or U11109 (N_11109,N_5286,N_9234);
and U11110 (N_11110,N_8224,N_9695);
nor U11111 (N_11111,N_8924,N_5776);
nor U11112 (N_11112,N_6442,N_8277);
and U11113 (N_11113,N_6650,N_5327);
and U11114 (N_11114,N_5087,N_5419);
xnor U11115 (N_11115,N_6416,N_9636);
or U11116 (N_11116,N_5667,N_7461);
nand U11117 (N_11117,N_7838,N_7854);
nand U11118 (N_11118,N_7216,N_6867);
nand U11119 (N_11119,N_8691,N_8076);
nand U11120 (N_11120,N_7426,N_8306);
or U11121 (N_11121,N_9032,N_9363);
and U11122 (N_11122,N_6288,N_5052);
and U11123 (N_11123,N_9643,N_7173);
nor U11124 (N_11124,N_5393,N_7837);
or U11125 (N_11125,N_7543,N_9831);
or U11126 (N_11126,N_8521,N_7176);
nand U11127 (N_11127,N_6420,N_5024);
nand U11128 (N_11128,N_6910,N_5332);
or U11129 (N_11129,N_7720,N_5226);
nand U11130 (N_11130,N_9463,N_6402);
or U11131 (N_11131,N_5838,N_6411);
and U11132 (N_11132,N_8396,N_8245);
nor U11133 (N_11133,N_9157,N_9349);
nor U11134 (N_11134,N_6546,N_7692);
and U11135 (N_11135,N_5057,N_7850);
nand U11136 (N_11136,N_6255,N_8063);
and U11137 (N_11137,N_9790,N_5317);
nand U11138 (N_11138,N_5867,N_6328);
or U11139 (N_11139,N_6353,N_7335);
or U11140 (N_11140,N_6706,N_6627);
or U11141 (N_11141,N_7494,N_6614);
nor U11142 (N_11142,N_6167,N_9910);
nor U11143 (N_11143,N_9710,N_9843);
or U11144 (N_11144,N_9809,N_7391);
nor U11145 (N_11145,N_7905,N_6709);
nand U11146 (N_11146,N_7153,N_9307);
and U11147 (N_11147,N_5963,N_5112);
or U11148 (N_11148,N_6386,N_9673);
nor U11149 (N_11149,N_6133,N_7669);
nand U11150 (N_11150,N_8464,N_5915);
or U11151 (N_11151,N_5039,N_7264);
nor U11152 (N_11152,N_7774,N_5420);
or U11153 (N_11153,N_7684,N_8198);
or U11154 (N_11154,N_7155,N_8286);
and U11155 (N_11155,N_7509,N_5834);
nor U11156 (N_11156,N_9035,N_6899);
or U11157 (N_11157,N_7316,N_7158);
nand U11158 (N_11158,N_7257,N_6384);
nor U11159 (N_11159,N_8670,N_6843);
nand U11160 (N_11160,N_5974,N_6777);
and U11161 (N_11161,N_8617,N_9985);
or U11162 (N_11162,N_6505,N_9408);
or U11163 (N_11163,N_6010,N_8395);
nand U11164 (N_11164,N_7682,N_8985);
and U11165 (N_11165,N_7208,N_5505);
or U11166 (N_11166,N_9196,N_6457);
nor U11167 (N_11167,N_6250,N_6360);
or U11168 (N_11168,N_8598,N_7945);
or U11169 (N_11169,N_5713,N_7083);
nor U11170 (N_11170,N_8843,N_7840);
nand U11171 (N_11171,N_5941,N_7589);
nor U11172 (N_11172,N_6080,N_5390);
nor U11173 (N_11173,N_7084,N_8784);
and U11174 (N_11174,N_7320,N_8538);
nand U11175 (N_11175,N_7052,N_6655);
nand U11176 (N_11176,N_5189,N_7166);
and U11177 (N_11177,N_7994,N_5010);
nor U11178 (N_11178,N_8910,N_6759);
nand U11179 (N_11179,N_8195,N_6695);
or U11180 (N_11180,N_9273,N_5609);
or U11181 (N_11181,N_7440,N_5465);
nor U11182 (N_11182,N_6651,N_6562);
nand U11183 (N_11183,N_9852,N_8221);
nand U11184 (N_11184,N_8541,N_6475);
or U11185 (N_11185,N_8980,N_8935);
nand U11186 (N_11186,N_9007,N_8588);
nor U11187 (N_11187,N_9848,N_5552);
or U11188 (N_11188,N_9624,N_6403);
nand U11189 (N_11189,N_7381,N_5060);
or U11190 (N_11190,N_5702,N_8735);
nand U11191 (N_11191,N_6132,N_7039);
and U11192 (N_11192,N_5944,N_7517);
or U11193 (N_11193,N_6744,N_5652);
nor U11194 (N_11194,N_6537,N_9133);
nand U11195 (N_11195,N_6784,N_9129);
or U11196 (N_11196,N_5355,N_8031);
nor U11197 (N_11197,N_5485,N_7565);
nand U11198 (N_11198,N_9361,N_9875);
nand U11199 (N_11199,N_8621,N_7742);
or U11200 (N_11200,N_6665,N_5871);
or U11201 (N_11201,N_6144,N_5873);
nor U11202 (N_11202,N_9305,N_7903);
nor U11203 (N_11203,N_8929,N_5456);
or U11204 (N_11204,N_8104,N_7568);
nand U11205 (N_11205,N_7249,N_9767);
and U11206 (N_11206,N_5243,N_5986);
nand U11207 (N_11207,N_5045,N_9347);
nor U11208 (N_11208,N_7951,N_5687);
and U11209 (N_11209,N_6079,N_8888);
nor U11210 (N_11210,N_7341,N_8968);
nor U11211 (N_11211,N_8681,N_5065);
nand U11212 (N_11212,N_8883,N_7940);
nand U11213 (N_11213,N_6940,N_6296);
nor U11214 (N_11214,N_6106,N_9259);
nand U11215 (N_11215,N_7980,N_8259);
nand U11216 (N_11216,N_9918,N_5219);
and U11217 (N_11217,N_8687,N_9386);
nand U11218 (N_11218,N_9042,N_5937);
or U11219 (N_11219,N_8049,N_7266);
or U11220 (N_11220,N_9194,N_5071);
nand U11221 (N_11221,N_7344,N_5666);
and U11222 (N_11222,N_7401,N_7523);
nor U11223 (N_11223,N_8424,N_5375);
nand U11224 (N_11224,N_5062,N_6504);
or U11225 (N_11225,N_9605,N_5187);
or U11226 (N_11226,N_9219,N_7293);
and U11227 (N_11227,N_8774,N_5904);
nand U11228 (N_11228,N_6935,N_6984);
nor U11229 (N_11229,N_7438,N_8488);
and U11230 (N_11230,N_5735,N_6428);
nor U11231 (N_11231,N_9893,N_6406);
or U11232 (N_11232,N_8120,N_7207);
and U11233 (N_11233,N_9477,N_8126);
nand U11234 (N_11234,N_5376,N_6439);
nor U11235 (N_11235,N_7614,N_8423);
or U11236 (N_11236,N_7511,N_6032);
nor U11237 (N_11237,N_7966,N_9860);
nand U11238 (N_11238,N_8187,N_9205);
nand U11239 (N_11239,N_6371,N_5257);
and U11240 (N_11240,N_6004,N_8715);
nor U11241 (N_11241,N_7195,N_6564);
or U11242 (N_11242,N_8976,N_7977);
nand U11243 (N_11243,N_7629,N_5752);
nand U11244 (N_11244,N_5868,N_7307);
or U11245 (N_11245,N_9182,N_5951);
and U11246 (N_11246,N_6429,N_5608);
nand U11247 (N_11247,N_5954,N_9457);
nor U11248 (N_11248,N_8099,N_7310);
or U11249 (N_11249,N_6494,N_9328);
nand U11250 (N_11250,N_6684,N_9089);
and U11251 (N_11251,N_7047,N_8859);
nand U11252 (N_11252,N_7590,N_6671);
and U11253 (N_11253,N_5028,N_7863);
or U11254 (N_11254,N_7191,N_5854);
nand U11255 (N_11255,N_8558,N_8778);
nand U11256 (N_11256,N_9280,N_8421);
nand U11257 (N_11257,N_5325,N_8303);
nor U11258 (N_11258,N_9218,N_6325);
and U11259 (N_11259,N_8403,N_6750);
and U11260 (N_11260,N_8895,N_8586);
nand U11261 (N_11261,N_7979,N_5479);
and U11262 (N_11262,N_5965,N_9416);
or U11263 (N_11263,N_9499,N_9598);
nand U11264 (N_11264,N_5507,N_5464);
or U11265 (N_11265,N_5215,N_9537);
or U11266 (N_11266,N_7128,N_8258);
nand U11267 (N_11267,N_7290,N_7429);
xnor U11268 (N_11268,N_5522,N_8647);
or U11269 (N_11269,N_6111,N_8336);
nand U11270 (N_11270,N_7373,N_7267);
nand U11271 (N_11271,N_8615,N_5193);
and U11272 (N_11272,N_9890,N_9181);
or U11273 (N_11273,N_5746,N_7380);
or U11274 (N_11274,N_5957,N_5872);
and U11275 (N_11275,N_9800,N_5884);
or U11276 (N_11276,N_6817,N_5133);
nor U11277 (N_11277,N_6538,N_5277);
nor U11278 (N_11278,N_7502,N_6835);
nand U11279 (N_11279,N_6185,N_8587);
nor U11280 (N_11280,N_6856,N_9821);
nor U11281 (N_11281,N_5348,N_9168);
nand U11282 (N_11282,N_7018,N_5015);
and U11283 (N_11283,N_7906,N_5515);
nand U11284 (N_11284,N_7092,N_8721);
xnor U11285 (N_11285,N_5742,N_5012);
nand U11286 (N_11286,N_7792,N_9188);
or U11287 (N_11287,N_6764,N_5577);
nor U11288 (N_11288,N_9370,N_9126);
nor U11289 (N_11289,N_5788,N_8320);
and U11290 (N_11290,N_9779,N_6309);
nor U11291 (N_11291,N_6741,N_9541);
and U11292 (N_11292,N_5001,N_7722);
nand U11293 (N_11293,N_7114,N_6771);
nand U11294 (N_11294,N_9888,N_6389);
nor U11295 (N_11295,N_6939,N_5692);
nor U11296 (N_11296,N_5519,N_7368);
nor U11297 (N_11297,N_9849,N_5533);
nor U11298 (N_11298,N_6388,N_8660);
nor U11299 (N_11299,N_5108,N_9095);
or U11300 (N_11300,N_7436,N_7393);
and U11301 (N_11301,N_5901,N_6390);
nor U11302 (N_11302,N_9667,N_8729);
or U11303 (N_11303,N_5309,N_6369);
or U11304 (N_11304,N_6754,N_7592);
nor U11305 (N_11305,N_5379,N_6727);
nand U11306 (N_11306,N_5544,N_9485);
or U11307 (N_11307,N_7263,N_8042);
nor U11308 (N_11308,N_7087,N_5733);
nand U11309 (N_11309,N_8561,N_6725);
nor U11310 (N_11310,N_8716,N_7178);
and U11311 (N_11311,N_6805,N_8323);
nor U11312 (N_11312,N_7706,N_5784);
nor U11313 (N_11313,N_5073,N_9988);
nand U11314 (N_11314,N_5141,N_5557);
and U11315 (N_11315,N_7388,N_6653);
and U11316 (N_11316,N_7805,N_9641);
nor U11317 (N_11317,N_7221,N_7002);
nand U11318 (N_11318,N_6030,N_7743);
and U11319 (N_11319,N_8890,N_9850);
and U11320 (N_11320,N_9613,N_9351);
and U11321 (N_11321,N_9911,N_5463);
or U11322 (N_11322,N_9423,N_5748);
and U11323 (N_11323,N_7194,N_8986);
or U11324 (N_11324,N_8211,N_7740);
and U11325 (N_11325,N_5266,N_7933);
nand U11326 (N_11326,N_6957,N_9564);
nand U11327 (N_11327,N_7300,N_8800);
nor U11328 (N_11328,N_5161,N_8889);
or U11329 (N_11329,N_8368,N_8941);
or U11330 (N_11330,N_5200,N_5530);
or U11331 (N_11331,N_5339,N_6966);
nor U11332 (N_11332,N_9507,N_7390);
or U11333 (N_11333,N_7570,N_6066);
and U11334 (N_11334,N_8854,N_7417);
and U11335 (N_11335,N_9776,N_8297);
nor U11336 (N_11336,N_9738,N_6499);
and U11337 (N_11337,N_9015,N_6834);
nor U11338 (N_11338,N_7134,N_6535);
nor U11339 (N_11339,N_7834,N_6683);
nand U11340 (N_11340,N_8553,N_9990);
nor U11341 (N_11341,N_9355,N_5356);
or U11342 (N_11342,N_7473,N_9136);
nor U11343 (N_11343,N_8234,N_9544);
nand U11344 (N_11344,N_7077,N_8510);
nand U11345 (N_11345,N_6400,N_8717);
nor U11346 (N_11346,N_8962,N_7481);
or U11347 (N_11347,N_5054,N_6308);
or U11348 (N_11348,N_5945,N_5167);
nor U11349 (N_11349,N_7452,N_5928);
nand U11350 (N_11350,N_7789,N_5727);
nor U11351 (N_11351,N_7689,N_9209);
nand U11352 (N_11352,N_5857,N_5524);
and U11353 (N_11353,N_8542,N_7585);
and U11354 (N_11354,N_7787,N_9963);
or U11355 (N_11355,N_7394,N_9313);
nor U11356 (N_11356,N_5370,N_5059);
nand U11357 (N_11357,N_7450,N_5630);
nor U11358 (N_11358,N_7866,N_9176);
nand U11359 (N_11359,N_8508,N_5645);
nand U11360 (N_11360,N_8879,N_5889);
nand U11361 (N_11361,N_6373,N_8382);
or U11362 (N_11362,N_9010,N_7175);
and U11363 (N_11363,N_8035,N_5641);
and U11364 (N_11364,N_9045,N_6342);
and U11365 (N_11365,N_8369,N_9059);
and U11366 (N_11366,N_8956,N_8404);
nand U11367 (N_11367,N_9635,N_7796);
and U11368 (N_11368,N_5333,N_8111);
xnor U11369 (N_11369,N_8694,N_6626);
and U11370 (N_11370,N_7124,N_8530);
or U11371 (N_11371,N_9394,N_5816);
or U11372 (N_11372,N_8275,N_9251);
or U11373 (N_11373,N_8226,N_7211);
nor U11374 (N_11374,N_9808,N_5736);
and U11375 (N_11375,N_6973,N_8673);
nor U11376 (N_11376,N_8315,N_7601);
nor U11377 (N_11377,N_7357,N_5709);
or U11378 (N_11378,N_8208,N_8311);
or U11379 (N_11379,N_5555,N_5625);
and U11380 (N_11380,N_6547,N_8902);
nor U11381 (N_11381,N_5669,N_6408);
and U11382 (N_11382,N_5761,N_9960);
nor U11383 (N_11383,N_9662,N_6495);
nand U11384 (N_11384,N_8732,N_5354);
nand U11385 (N_11385,N_9697,N_5064);
and U11386 (N_11386,N_9573,N_6763);
or U11387 (N_11387,N_8492,N_6438);
nor U11388 (N_11388,N_8572,N_9657);
and U11389 (N_11389,N_5885,N_7217);
nor U11390 (N_11390,N_6636,N_6713);
or U11391 (N_11391,N_5442,N_5827);
or U11392 (N_11392,N_7009,N_6561);
or U11393 (N_11393,N_6477,N_9440);
or U11394 (N_11394,N_5903,N_6755);
nor U11395 (N_11395,N_6731,N_7635);
nor U11396 (N_11396,N_8531,N_9106);
and U11397 (N_11397,N_8937,N_5936);
or U11398 (N_11398,N_7733,N_5810);
nand U11399 (N_11399,N_7145,N_6618);
and U11400 (N_11400,N_5812,N_9480);
or U11401 (N_11401,N_7434,N_8600);
and U11402 (N_11402,N_7044,N_6162);
or U11403 (N_11403,N_6430,N_6821);
and U11404 (N_11404,N_6974,N_6569);
or U11405 (N_11405,N_7081,N_9978);
or U11406 (N_11406,N_8204,N_5020);
and U11407 (N_11407,N_9295,N_6196);
nand U11408 (N_11408,N_9149,N_6927);
or U11409 (N_11409,N_6136,N_7870);
or U11410 (N_11410,N_5328,N_6916);
nor U11411 (N_11411,N_9377,N_9877);
nor U11412 (N_11412,N_8191,N_9446);
or U11413 (N_11413,N_5546,N_8305);
or U11414 (N_11414,N_6275,N_5451);
nand U11415 (N_11415,N_5035,N_8356);
nor U11416 (N_11416,N_7515,N_9434);
nand U11417 (N_11417,N_7402,N_7812);
or U11418 (N_11418,N_9845,N_9025);
and U11419 (N_11419,N_9388,N_8632);
or U11420 (N_11420,N_6738,N_7456);
and U11421 (N_11421,N_6097,N_7961);
or U11422 (N_11422,N_6518,N_8822);
and U11423 (N_11423,N_6063,N_5048);
nor U11424 (N_11424,N_5121,N_5304);
nor U11425 (N_11425,N_5774,N_6831);
nand U11426 (N_11426,N_6137,N_9238);
nor U11427 (N_11427,N_7782,N_9676);
or U11428 (N_11428,N_5856,N_5658);
nor U11429 (N_11429,N_9299,N_6654);
or U11430 (N_11430,N_5906,N_5030);
and U11431 (N_11431,N_6737,N_5717);
nand U11432 (N_11432,N_7213,N_9944);
nand U11433 (N_11433,N_8943,N_7314);
and U11434 (N_11434,N_8959,N_9806);
and U11435 (N_11435,N_7289,N_5990);
and U11436 (N_11436,N_8218,N_7234);
or U11437 (N_11437,N_9340,N_7724);
nor U11438 (N_11438,N_5128,N_6712);
and U11439 (N_11439,N_5258,N_7526);
nand U11440 (N_11440,N_7423,N_8282);
or U11441 (N_11441,N_8246,N_9761);
or U11442 (N_11442,N_7268,N_9586);
or U11443 (N_11443,N_5631,N_9516);
nor U11444 (N_11444,N_9005,N_8630);
or U11445 (N_11445,N_6931,N_9873);
and U11446 (N_11446,N_9663,N_7895);
or U11447 (N_11447,N_9160,N_9336);
nand U11448 (N_11448,N_8367,N_7143);
nand U11449 (N_11449,N_5360,N_5359);
or U11450 (N_11450,N_9429,N_5033);
and U11451 (N_11451,N_8512,N_6945);
nor U11452 (N_11452,N_5765,N_5783);
nor U11453 (N_11453,N_8090,N_9756);
or U11454 (N_11454,N_8454,N_5495);
nand U11455 (N_11455,N_5582,N_9033);
or U11456 (N_11456,N_9672,N_5382);
nor U11457 (N_11457,N_9731,N_6081);
or U11458 (N_11458,N_9091,N_9487);
and U11459 (N_11459,N_8626,N_8551);
nor U11460 (N_11460,N_5084,N_6553);
or U11461 (N_11461,N_5912,N_8515);
or U11462 (N_11462,N_6241,N_5259);
nand U11463 (N_11463,N_7413,N_5247);
and U11464 (N_11464,N_7911,N_7379);
and U11465 (N_11465,N_9166,N_7086);
or U11466 (N_11466,N_9665,N_9100);
nand U11467 (N_11467,N_8240,N_7342);
and U11468 (N_11468,N_5989,N_6269);
xor U11469 (N_11469,N_6116,N_5780);
nand U11470 (N_11470,N_7189,N_6199);
nor U11471 (N_11471,N_9633,N_7534);
or U11472 (N_11472,N_7781,N_8926);
or U11473 (N_11473,N_7352,N_6708);
and U11474 (N_11474,N_7868,N_8758);
and U11475 (N_11475,N_6776,N_7167);
and U11476 (N_11476,N_9345,N_7810);
nor U11477 (N_11477,N_7797,N_8754);
or U11478 (N_11478,N_9262,N_6946);
or U11479 (N_11479,N_6108,N_5926);
or U11480 (N_11480,N_5679,N_9755);
and U11481 (N_11481,N_9549,N_7006);
and U11482 (N_11482,N_9352,N_7382);
or U11483 (N_11483,N_8645,N_9123);
and U11484 (N_11484,N_5605,N_5423);
or U11485 (N_11485,N_7727,N_6282);
and U11486 (N_11486,N_9360,N_5734);
nor U11487 (N_11487,N_8116,N_7193);
or U11488 (N_11488,N_5696,N_7085);
and U11489 (N_11489,N_7313,N_5478);
nor U11490 (N_11490,N_5101,N_6466);
nand U11491 (N_11491,N_7472,N_6443);
nand U11492 (N_11492,N_7139,N_8744);
or U11493 (N_11493,N_7271,N_8874);
nand U11494 (N_11494,N_9569,N_6994);
nor U11495 (N_11495,N_5879,N_9938);
and U11496 (N_11496,N_5151,N_8287);
nand U11497 (N_11497,N_7097,N_9037);
nor U11498 (N_11498,N_8575,N_6279);
and U11499 (N_11499,N_6335,N_7639);
nor U11500 (N_11500,N_5220,N_9364);
nand U11501 (N_11501,N_5416,N_6418);
or U11502 (N_11502,N_5067,N_7981);
nor U11503 (N_11503,N_9517,N_6942);
or U11504 (N_11504,N_5299,N_7815);
or U11505 (N_11505,N_8828,N_7744);
and U11506 (N_11506,N_7113,N_9857);
nand U11507 (N_11507,N_7654,N_9051);
or U11508 (N_11508,N_8905,N_5227);
or U11509 (N_11509,N_7747,N_8269);
nand U11510 (N_11510,N_5799,N_8992);
and U11511 (N_11511,N_8075,N_8456);
or U11512 (N_11512,N_7657,N_8346);
and U11513 (N_11513,N_9215,N_5852);
nor U11514 (N_11514,N_8433,N_9783);
and U11515 (N_11515,N_6396,N_8662);
nand U11516 (N_11516,N_5350,N_7583);
nor U11517 (N_11517,N_6298,N_7731);
nand U11518 (N_11518,N_8262,N_6050);
nand U11519 (N_11519,N_8276,N_7627);
and U11520 (N_11520,N_9248,N_8149);
or U11521 (N_11521,N_5455,N_8064);
or U11522 (N_11522,N_7828,N_6554);
nor U11523 (N_11523,N_7546,N_5798);
nand U11524 (N_11524,N_6987,N_8712);
nand U11525 (N_11525,N_6953,N_5319);
nand U11526 (N_11526,N_5408,N_9392);
nor U11527 (N_11527,N_5272,N_5880);
and U11528 (N_11528,N_5248,N_6975);
nor U11529 (N_11529,N_5629,N_6395);
nor U11530 (N_11530,N_5964,N_6956);
and U11531 (N_11531,N_7922,N_9872);
nor U11532 (N_11532,N_5898,N_6474);
nand U11533 (N_11533,N_6729,N_7399);
and U11534 (N_11534,N_5591,N_5826);
or U11535 (N_11535,N_5056,N_7548);
and U11536 (N_11536,N_7104,N_7637);
and U11537 (N_11537,N_7457,N_7115);
nand U11538 (N_11538,N_9376,N_8189);
and U11539 (N_11539,N_8952,N_6271);
and U11540 (N_11540,N_6791,N_6593);
or U11541 (N_11541,N_6949,N_9653);
nand U11542 (N_11542,N_6986,N_7022);
or U11543 (N_11543,N_6980,N_6932);
or U11544 (N_11544,N_8073,N_6201);
or U11545 (N_11545,N_5361,N_9179);
and U11546 (N_11546,N_8916,N_8871);
nor U11547 (N_11547,N_7432,N_7349);
and U11548 (N_11548,N_7205,N_7165);
xor U11549 (N_11549,N_6234,N_8808);
nand U11550 (N_11550,N_9530,N_9946);
and U11551 (N_11551,N_8944,N_6873);
and U11552 (N_11552,N_5553,N_8072);
nor U11553 (N_11553,N_9321,N_7064);
and U11554 (N_11554,N_6815,N_6285);
or U11555 (N_11555,N_5647,N_7061);
nand U11556 (N_11556,N_8719,N_8027);
and U11557 (N_11557,N_7369,N_8345);
and U11558 (N_11558,N_5385,N_8079);
or U11559 (N_11559,N_7687,N_6719);
nand U11560 (N_11560,N_7409,N_6668);
and U11561 (N_11561,N_7309,N_9524);
or U11562 (N_11562,N_7008,N_8870);
and U11563 (N_11563,N_5558,N_9520);
and U11564 (N_11564,N_8979,N_9812);
or U11565 (N_11565,N_5063,N_5460);
nand U11566 (N_11566,N_8124,N_5403);
nand U11567 (N_11567,N_5676,N_9187);
nand U11568 (N_11568,N_9421,N_6247);
nor U11569 (N_11569,N_9183,N_7921);
and U11570 (N_11570,N_7821,N_7055);
or U11571 (N_11571,N_8386,N_9027);
nor U11572 (N_11572,N_6287,N_5083);
or U11573 (N_11573,N_8934,N_6351);
or U11574 (N_11574,N_6336,N_7042);
and U11575 (N_11575,N_9727,N_7093);
nor U11576 (N_11576,N_7386,N_6357);
or U11577 (N_11577,N_7375,N_5394);
nor U11578 (N_11578,N_6244,N_8165);
or U11579 (N_11579,N_8711,N_7693);
nand U11580 (N_11580,N_6512,N_8820);
and U11581 (N_11581,N_9412,N_5621);
or U11582 (N_11582,N_6779,N_5521);
nand U11583 (N_11583,N_9109,N_8453);
nor U11584 (N_11584,N_9515,N_9018);
nand U11585 (N_11585,N_7929,N_6286);
and U11586 (N_11586,N_9575,N_5017);
nor U11587 (N_11587,N_5743,N_5191);
nand U11588 (N_11588,N_8089,N_7058);
nor U11589 (N_11589,N_5058,N_7325);
nand U11590 (N_11590,N_8083,N_8183);
nand U11591 (N_11591,N_7256,N_6944);
nand U11592 (N_11592,N_6315,N_5514);
nor U11593 (N_11593,N_9221,N_6427);
nor U11594 (N_11594,N_7827,N_7206);
nor U11595 (N_11595,N_6084,N_8597);
nand U11596 (N_11596,N_8266,N_8332);
and U11597 (N_11597,N_7295,N_8616);
and U11598 (N_11598,N_5424,N_9899);
nand U11599 (N_11599,N_9255,N_9437);
and U11600 (N_11600,N_8267,N_9601);
and U11601 (N_11601,N_8020,N_9502);
nand U11602 (N_11602,N_9122,N_7421);
and U11603 (N_11603,N_9561,N_9171);
nand U11604 (N_11604,N_7652,N_6245);
nand U11605 (N_11605,N_9184,N_6068);
nor U11606 (N_11606,N_7685,N_9884);
nand U11607 (N_11607,N_9859,N_6015);
or U11608 (N_11608,N_9177,N_7847);
and U11609 (N_11609,N_8247,N_7901);
or U11610 (N_11610,N_6322,N_8106);
nand U11611 (N_11611,N_8864,N_9993);
and U11612 (N_11612,N_9546,N_7303);
nand U11613 (N_11613,N_7803,N_9378);
nor U11614 (N_11614,N_5532,N_5821);
nor U11615 (N_11615,N_5565,N_6748);
nor U11616 (N_11616,N_6962,N_8439);
and U11617 (N_11617,N_9282,N_7670);
nor U11618 (N_11618,N_6091,N_9475);
or U11619 (N_11619,N_5598,N_5697);
and U11620 (N_11620,N_8136,N_8933);
and U11621 (N_11621,N_7337,N_6113);
nor U11622 (N_11622,N_6509,N_7057);
or U11623 (N_11623,N_9137,N_8225);
and U11624 (N_11624,N_5662,N_9968);
nand U11625 (N_11625,N_9488,N_6793);
and U11626 (N_11626,N_9615,N_7996);
and U11627 (N_11627,N_9012,N_5612);
nand U11628 (N_11628,N_5320,N_7296);
and U11629 (N_11629,N_8069,N_7278);
and U11630 (N_11630,N_9791,N_9879);
nand U11631 (N_11631,N_6840,N_7172);
nand U11632 (N_11632,N_8117,N_7033);
or U11633 (N_11633,N_5255,N_5934);
and U11634 (N_11634,N_9074,N_9718);
and U11635 (N_11635,N_9642,N_5998);
or U11636 (N_11636,N_5111,N_9112);
or U11637 (N_11637,N_9379,N_8927);
nor U11638 (N_11638,N_9471,N_7726);
nor U11639 (N_11639,N_5281,N_8583);
or U11640 (N_11640,N_5077,N_6226);
nand U11641 (N_11641,N_8119,N_6610);
and U11642 (N_11642,N_6602,N_6666);
or U11643 (N_11643,N_7520,N_7339);
and U11644 (N_11644,N_8585,N_6516);
nand U11645 (N_11645,N_6837,N_6700);
nand U11646 (N_11646,N_5650,N_6517);
or U11647 (N_11647,N_5574,N_9780);
or U11648 (N_11648,N_8199,N_5345);
nand U11649 (N_11649,N_7993,N_5169);
nand U11650 (N_11650,N_7411,N_5289);
or U11651 (N_11651,N_8608,N_8068);
nand U11652 (N_11652,N_6691,N_9995);
nor U11653 (N_11653,N_7054,N_8493);
or U11654 (N_11654,N_6533,N_5450);
nand U11655 (N_11655,N_6870,N_7986);
or U11656 (N_11656,N_7301,N_7735);
nor U11657 (N_11657,N_5174,N_7765);
and U11658 (N_11658,N_5620,N_5651);
nand U11659 (N_11659,N_7280,N_7572);
or U11660 (N_11660,N_5150,N_6363);
nand U11661 (N_11661,N_7508,N_9959);
and U11662 (N_11662,N_6358,N_6238);
and U11663 (N_11663,N_5818,N_7407);
or U11664 (N_11664,N_9506,N_7567);
nand U11665 (N_11665,N_5349,N_6029);
nor U11666 (N_11666,N_6592,N_8131);
and U11667 (N_11667,N_8298,N_9972);
nor U11668 (N_11668,N_6021,N_5583);
and U11669 (N_11669,N_9600,N_7776);
nor U11670 (N_11670,N_5622,N_8040);
and U11671 (N_11671,N_8483,N_8801);
nor U11672 (N_11672,N_6936,N_8248);
and U11673 (N_11673,N_5905,N_8216);
and U11674 (N_11674,N_7745,N_9132);
or U11675 (N_11675,N_9580,N_5092);
and U11676 (N_11676,N_6049,N_5085);
nand U11677 (N_11677,N_5847,N_7930);
or U11678 (N_11678,N_9117,N_5380);
or U11679 (N_11679,N_5336,N_8172);
nor U11680 (N_11680,N_8851,N_7633);
nor U11681 (N_11681,N_7027,N_8016);
nand U11682 (N_11682,N_6352,N_5916);
or U11683 (N_11683,N_9265,N_8228);
nor U11684 (N_11684,N_9410,N_9501);
or U11685 (N_11685,N_7645,N_8991);
nor U11686 (N_11686,N_8760,N_9763);
and U11687 (N_11687,N_8936,N_8067);
nand U11688 (N_11688,N_7080,N_8970);
nor U11689 (N_11689,N_5982,N_8137);
nand U11690 (N_11690,N_5347,N_7034);
nor U11691 (N_11691,N_8272,N_5767);
or U11692 (N_11692,N_6041,N_9304);
and U11693 (N_11693,N_9331,N_9227);
nand U11694 (N_11694,N_9029,N_9690);
and U11695 (N_11695,N_6685,N_6297);
nand U11696 (N_11696,N_7096,N_6778);
or U11697 (N_11697,N_7643,N_6649);
or U11698 (N_11698,N_9713,N_9228);
nand U11699 (N_11699,N_7486,N_5399);
nand U11700 (N_11700,N_6823,N_5731);
nor U11701 (N_11701,N_8371,N_8942);
nand U11702 (N_11702,N_6317,N_5201);
nand U11703 (N_11703,N_8677,N_6907);
and U11704 (N_11704,N_7245,N_7716);
or U11705 (N_11705,N_5616,N_7410);
nand U11706 (N_11706,N_8391,N_8350);
and U11707 (N_11707,N_5991,N_5881);
or U11708 (N_11708,N_7702,N_5461);
nor U11709 (N_11709,N_7001,N_9793);
nor U11710 (N_11710,N_6300,N_6038);
nand U11711 (N_11711,N_8355,N_9300);
or U11712 (N_11712,N_6696,N_9092);
or U11713 (N_11713,N_9519,N_7287);
or U11714 (N_11714,N_9481,N_6319);
nor U11715 (N_11715,N_5214,N_8292);
nand U11716 (N_11716,N_7451,N_6878);
and U11717 (N_11717,N_5224,N_9070);
nand U11718 (N_11718,N_5550,N_6421);
and U11719 (N_11719,N_7982,N_6631);
nor U11720 (N_11720,N_9617,N_5543);
and U11721 (N_11721,N_8166,N_9139);
and U11722 (N_11722,N_9243,N_8850);
nand U11723 (N_11723,N_6365,N_8095);
nand U11724 (N_11724,N_5738,N_7893);
xnor U11725 (N_11725,N_9001,N_7358);
nand U11726 (N_11726,N_7936,N_9825);
and U11727 (N_11727,N_8466,N_7831);
nand U11728 (N_11728,N_9267,N_8628);
nand U11729 (N_11729,N_8150,N_7845);
nand U11730 (N_11730,N_5177,N_7532);
or U11731 (N_11731,N_5011,N_9231);
nand U11732 (N_11732,N_7247,N_8635);
nand U11733 (N_11733,N_9785,N_6216);
nand U11734 (N_11734,N_8443,N_7730);
nor U11735 (N_11735,N_8358,N_9533);
nand U11736 (N_11736,N_5714,N_7496);
nor U11737 (N_11737,N_6433,N_5156);
nand U11738 (N_11738,N_9811,N_8468);
nor U11739 (N_11739,N_7804,N_7939);
or U11740 (N_11740,N_5476,N_5337);
or U11741 (N_11741,N_7201,N_9772);
xnor U11742 (N_11742,N_7612,N_7649);
nand U11743 (N_11743,N_9409,N_8500);
nor U11744 (N_11744,N_5770,N_6824);
nor U11745 (N_11745,N_6656,N_8799);
and U11746 (N_11746,N_6550,N_6864);
nand U11747 (N_11747,N_7069,N_9474);
nor U11748 (N_11748,N_8467,N_8319);
nand U11749 (N_11749,N_7607,N_5404);
or U11750 (N_11750,N_6364,N_8834);
and U11751 (N_11751,N_7059,N_9715);
or U11752 (N_11752,N_9926,N_8304);
and U11753 (N_11753,N_9131,N_7311);
and U11754 (N_11754,N_9822,N_6378);
nor U11755 (N_11755,N_8702,N_8059);
or U11756 (N_11756,N_8328,N_5448);
or U11757 (N_11757,N_8675,N_9214);
nand U11758 (N_11758,N_5811,N_7038);
nand U11759 (N_11759,N_5814,N_8981);
nor U11760 (N_11760,N_5547,N_6217);
or U11761 (N_11761,N_9545,N_9523);
and U11762 (N_11762,N_8357,N_9773);
and U11763 (N_11763,N_8830,N_5542);
and U11764 (N_11764,N_5549,N_9206);
nor U11765 (N_11765,N_7190,N_6790);
or U11766 (N_11766,N_6858,N_6179);
nand U11767 (N_11767,N_6775,N_9902);
and U11768 (N_11768,N_6314,N_6686);
nand U11769 (N_11769,N_8244,N_6142);
nand U11770 (N_11770,N_6797,N_7512);
and U11771 (N_11771,N_8436,N_9403);
nand U11772 (N_11772,N_6013,N_9612);
nor U11773 (N_11773,N_8642,N_7659);
nor U11774 (N_11774,N_5051,N_7123);
nand U11775 (N_11775,N_8088,N_9195);
or U11776 (N_11776,N_8938,N_6393);
xnor U11777 (N_11777,N_7377,N_8535);
nor U11778 (N_11778,N_9810,N_9594);
and U11779 (N_11779,N_9659,N_8993);
or U11780 (N_11780,N_8362,N_7312);
and U11781 (N_11781,N_6417,N_9281);
nand U11782 (N_11782,N_7772,N_8197);
nor U11783 (N_11783,N_8775,N_7203);
xor U11784 (N_11784,N_6344,N_9384);
nor U11785 (N_11785,N_7886,N_8416);
xnor U11786 (N_11786,N_9038,N_6705);
nand U11787 (N_11787,N_7960,N_5801);
nor U11788 (N_11788,N_5959,N_9802);
or U11789 (N_11789,N_9424,N_7525);
or U11790 (N_11790,N_8654,N_8108);
or U11791 (N_11791,N_8680,N_8037);
nand U11792 (N_11792,N_5143,N_6146);
and U11793 (N_11793,N_9080,N_7779);
nand U11794 (N_11794,N_8665,N_6415);
or U11795 (N_11795,N_5611,N_7656);
or U11796 (N_11796,N_9107,N_6368);
and U11797 (N_11797,N_5346,N_5996);
nor U11798 (N_11798,N_6673,N_5969);
nor U11799 (N_11799,N_7338,N_9173);
nor U11800 (N_11800,N_5671,N_8134);
or U11801 (N_11801,N_7890,N_5627);
nor U11802 (N_11802,N_7582,N_7852);
nor U11803 (N_11803,N_8742,N_5038);
or U11804 (N_11804,N_7299,N_6304);
nand U11805 (N_11805,N_9316,N_6745);
and U11806 (N_11806,N_6544,N_8960);
or U11807 (N_11807,N_6370,N_6121);
and U11808 (N_11808,N_5228,N_5602);
nor U11809 (N_11809,N_6675,N_6281);
and U11810 (N_11810,N_8949,N_9167);
nand U11811 (N_11811,N_9315,N_6437);
and U11812 (N_11812,N_9610,N_8683);
and U11813 (N_11813,N_5118,N_9660);
xor U11814 (N_11814,N_7574,N_6875);
and U11815 (N_11815,N_7392,N_8337);
nor U11816 (N_11816,N_7442,N_8983);
and U11817 (N_11817,N_5710,N_7019);
and U11818 (N_11818,N_7465,N_5803);
nor U11819 (N_11819,N_6879,N_9375);
or U11820 (N_11820,N_6062,N_7620);
nor U11821 (N_11821,N_9709,N_7117);
or U11822 (N_11822,N_9977,N_7282);
nand U11823 (N_11823,N_6458,N_5113);
nand U11824 (N_11824,N_8661,N_7273);
nand U11825 (N_11825,N_8643,N_7232);
nand U11826 (N_11826,N_7800,N_5939);
or U11827 (N_11827,N_6186,N_5122);
nand U11828 (N_11828,N_8852,N_6607);
nor U11829 (N_11829,N_7424,N_9263);
nand U11830 (N_11830,N_5269,N_5369);
and U11831 (N_11831,N_9604,N_9862);
nand U11832 (N_11832,N_7766,N_7843);
or U11833 (N_11833,N_6992,N_8353);
and U11834 (N_11834,N_7714,N_5095);
and U11835 (N_11835,N_5807,N_6401);
and U11836 (N_11836,N_8855,N_5142);
or U11837 (N_11837,N_9093,N_5184);
and U11838 (N_11838,N_9201,N_6473);
nand U11839 (N_11839,N_7991,N_7699);
nor U11840 (N_11840,N_6157,N_8793);
or U11841 (N_11841,N_8505,N_7164);
or U11842 (N_11842,N_9118,N_5517);
nand U11843 (N_11843,N_8101,N_5439);
or U11844 (N_11844,N_8430,N_5426);
or U11845 (N_11845,N_8360,N_5897);
nand U11846 (N_11846,N_7618,N_5745);
or U11847 (N_11847,N_8081,N_8300);
or U11848 (N_11848,N_6118,N_7270);
nor U11849 (N_11849,N_8746,N_5927);
and U11850 (N_11850,N_9241,N_6701);
or U11851 (N_11851,N_8062,N_5862);
or U11852 (N_11852,N_9625,N_9578);
or U11853 (N_11853,N_5305,N_7577);
nor U11854 (N_11854,N_9644,N_8928);
and U11855 (N_11855,N_8885,N_9489);
nor U11856 (N_11856,N_8641,N_7648);
nand U11857 (N_11857,N_9706,N_9270);
and U11858 (N_11858,N_8420,N_9702);
or U11859 (N_11859,N_5131,N_6354);
or U11860 (N_11860,N_5216,N_8946);
or U11861 (N_11861,N_5718,N_5759);
and U11862 (N_11862,N_5195,N_6246);
or U11863 (N_11863,N_9817,N_9141);
nand U11864 (N_11864,N_5908,N_5968);
nand U11865 (N_11865,N_9390,N_6257);
and U11866 (N_11866,N_8278,N_5023);
and U11867 (N_11867,N_5760,N_6757);
and U11868 (N_11868,N_5503,N_9422);
and U11869 (N_11869,N_6628,N_6772);
nand U11870 (N_11870,N_8984,N_9419);
xnor U11871 (N_11871,N_8243,N_9078);
and U11872 (N_11872,N_9889,N_6934);
and U11873 (N_11873,N_7606,N_8485);
nand U11874 (N_11874,N_8034,N_8330);
and U11875 (N_11875,N_6803,N_5232);
nor U11876 (N_11876,N_5835,N_5976);
nor U11877 (N_11877,N_6126,N_9692);
nand U11878 (N_11878,N_8038,N_5786);
or U11879 (N_11879,N_5653,N_8649);
and U11880 (N_11880,N_8438,N_6587);
nand U11881 (N_11881,N_5250,N_8465);
and U11882 (N_11882,N_5089,N_8666);
or U11883 (N_11883,N_8329,N_5251);
or U11884 (N_11884,N_8193,N_8019);
nand U11885 (N_11885,N_5983,N_5618);
and U11886 (N_11886,N_5179,N_7880);
or U11887 (N_11887,N_9948,N_8815);
nor U11888 (N_11888,N_8810,N_5268);
and U11889 (N_11889,N_8745,N_8610);
and U11890 (N_11890,N_5607,N_9236);
nor U11891 (N_11891,N_9987,N_9382);
and U11892 (N_11892,N_7763,N_5646);
or U11893 (N_11893,N_6292,N_5705);
and U11894 (N_11894,N_9332,N_5661);
and U11895 (N_11895,N_8497,N_7757);
or U11896 (N_11896,N_7518,N_5414);
nand U11897 (N_11897,N_8372,N_5617);
and U11898 (N_11898,N_5979,N_6310);
or U11899 (N_11899,N_9554,N_6960);
or U11900 (N_11900,N_7254,N_8783);
and U11901 (N_11901,N_8179,N_7437);
or U11902 (N_11902,N_5588,N_5855);
and U11903 (N_11903,N_5993,N_8032);
or U11904 (N_11904,N_7576,N_6574);
or U11905 (N_11905,N_5082,N_8915);
nor U11906 (N_11906,N_8932,N_5475);
or U11907 (N_11907,N_7334,N_5264);
nor U11908 (N_11908,N_6551,N_5711);
nor U11909 (N_11909,N_8539,N_8255);
and U11910 (N_11910,N_7653,N_6230);
or U11911 (N_11911,N_8523,N_5597);
nand U11912 (N_11912,N_5972,N_9311);
and U11913 (N_11913,N_6299,N_5302);
nor U11914 (N_11914,N_9260,N_5589);
nor U11915 (N_11915,N_9788,N_7995);
nand U11916 (N_11916,N_7946,N_6833);
nor U11917 (N_11917,N_7937,N_9077);
and U11918 (N_11918,N_7487,N_6678);
or U11919 (N_11919,N_6262,N_6171);
nand U11920 (N_11920,N_9929,N_5751);
nand U11921 (N_11921,N_8765,N_7142);
nor U11922 (N_11922,N_9749,N_5303);
nand U11923 (N_11923,N_8498,N_7016);
or U11924 (N_11924,N_6925,N_7547);
or U11925 (N_11925,N_9984,N_9671);
nand U11926 (N_11926,N_5288,N_9980);
and U11927 (N_11927,N_9539,N_9913);
and U11928 (N_11928,N_6192,N_7322);
nand U11929 (N_11929,N_6715,N_8620);
and U11930 (N_11930,N_9232,N_9804);
nand U11931 (N_11931,N_5000,N_8560);
nand U11932 (N_11932,N_6366,N_9023);
or U11933 (N_11933,N_7214,N_9906);
nor U11934 (N_11934,N_7100,N_8909);
and U11935 (N_11935,N_5595,N_9224);
or U11936 (N_11936,N_8025,N_6488);
xor U11937 (N_11937,N_6264,N_5487);
nand U11938 (N_11938,N_6638,N_7210);
nor U11939 (N_11939,N_6306,N_9711);
and U11940 (N_11940,N_7500,N_8181);
and U11941 (N_11941,N_5285,N_8428);
nor U11942 (N_11942,N_8698,N_9148);
and U11943 (N_11943,N_5924,N_5180);
nor U11944 (N_11944,N_7239,N_8112);
nor U11945 (N_11945,N_6076,N_5732);
or U11946 (N_11946,N_8682,N_9381);
and U11947 (N_11947,N_7985,N_8797);
nor U11948 (N_11948,N_8749,N_8570);
or U11949 (N_11949,N_7784,N_7269);
and U11950 (N_11950,N_8009,N_5663);
or U11951 (N_11951,N_8232,N_6630);
nand U11952 (N_11952,N_6573,N_7078);
and U11953 (N_11953,N_7956,N_5806);
nand U11954 (N_11954,N_6716,N_6998);
nor U11955 (N_11955,N_9264,N_5841);
nand U11956 (N_11956,N_7255,N_7501);
or U11957 (N_11957,N_5398,N_7040);
and U11958 (N_11958,N_7941,N_6173);
nor U11959 (N_11959,N_7544,N_6463);
and U11960 (N_11960,N_6789,N_9823);
or U11961 (N_11961,N_6259,N_6125);
nor U11962 (N_11962,N_7223,N_6811);
nor U11963 (N_11963,N_5729,N_6359);
and U11964 (N_11964,N_8169,N_6392);
nor U11965 (N_11965,N_7046,N_5144);
and U11966 (N_11966,N_6096,N_9894);
or U11967 (N_11967,N_7715,N_8410);
or U11968 (N_11968,N_8192,N_8906);
nand U11969 (N_11969,N_9225,N_5387);
nand U11970 (N_11970,N_6184,N_6071);
nand U11971 (N_11971,N_7439,N_5634);
nor U11972 (N_11972,N_8594,N_9576);
nand U11973 (N_11973,N_9426,N_8139);
nand U11974 (N_11974,N_7752,N_6887);
or U11975 (N_11975,N_9479,N_9058);
or U11976 (N_11976,N_7156,N_9400);
and U11977 (N_11977,N_7333,N_6412);
xor U11978 (N_11978,N_7608,N_9203);
nor U11979 (N_11979,N_5458,N_7355);
nand U11980 (N_11980,N_6374,N_5790);
or U11981 (N_11981,N_9445,N_5041);
nor U11982 (N_11982,N_8374,N_8486);
nor U11983 (N_11983,N_6734,N_6248);
nor U11984 (N_11984,N_6753,N_9212);
or U11985 (N_11985,N_7913,N_6794);
and U11986 (N_11986,N_6054,N_5462);
or U11987 (N_11987,N_5694,N_7769);
or U11988 (N_11988,N_6826,N_8160);
and U11989 (N_11989,N_7079,N_8504);
nand U11990 (N_11990,N_7746,N_5985);
nor U11991 (N_11991,N_8326,N_6733);
or U11992 (N_11992,N_6951,N_7202);
nor U11993 (N_11993,N_6579,N_7928);
and U11994 (N_11994,N_9050,N_6272);
or U11995 (N_11995,N_5124,N_8000);
nor U11996 (N_11996,N_9939,N_5955);
nor U11997 (N_11997,N_6492,N_8003);
or U11998 (N_11998,N_6372,N_6582);
nand U11999 (N_11999,N_6249,N_7718);
nor U12000 (N_12000,N_7491,N_6183);
nand U12001 (N_12001,N_6480,N_5902);
nor U12002 (N_12002,N_6997,N_9244);
nand U12003 (N_12003,N_7007,N_9832);
or U12004 (N_12004,N_5472,N_5853);
nand U12005 (N_12005,N_7998,N_5914);
nand U12006 (N_12006,N_7553,N_7281);
nand U12007 (N_12007,N_8469,N_9835);
nand U12008 (N_12008,N_5660,N_5590);
or U12009 (N_12009,N_5406,N_6608);
and U12010 (N_12010,N_9460,N_8001);
and U12011 (N_12011,N_6381,N_5072);
nor U12012 (N_12012,N_6151,N_8741);
and U12013 (N_12013,N_7712,N_7717);
or U12014 (N_12014,N_6521,N_7298);
or U12015 (N_12015,N_6301,N_5099);
nor U12016 (N_12016,N_6164,N_6577);
or U12017 (N_12017,N_7972,N_5665);
nand U12018 (N_12018,N_9478,N_9882);
nand U12019 (N_12019,N_8861,N_7522);
or U12020 (N_12020,N_6470,N_7187);
or U12021 (N_12021,N_6211,N_7860);
nand U12022 (N_12022,N_6552,N_9678);
and U12023 (N_12023,N_6581,N_9707);
nor U12024 (N_12024,N_5106,N_5107);
or U12025 (N_12025,N_6224,N_7024);
nand U12026 (N_12026,N_8163,N_6242);
or U12027 (N_12027,N_9242,N_5103);
or U12028 (N_12028,N_9666,N_5554);
nor U12029 (N_12029,N_7836,N_6307);
and U12030 (N_12030,N_6522,N_7533);
or U12031 (N_12031,N_7835,N_8777);
nor U12032 (N_12032,N_7184,N_9535);
or U12033 (N_12033,N_9632,N_7894);
nor U12034 (N_12034,N_9455,N_6227);
or U12035 (N_12035,N_9568,N_6152);
nor U12036 (N_12036,N_5980,N_5117);
nand U12037 (N_12037,N_7842,N_5160);
nand U12038 (N_12038,N_9584,N_9687);
nand U12039 (N_12039,N_5245,N_8747);
nand U12040 (N_12040,N_5567,N_5377);
nor U12041 (N_12041,N_5674,N_5935);
or U12042 (N_12042,N_8210,N_7094);
nor U12043 (N_12043,N_5119,N_5932);
and U12044 (N_12044,N_9744,N_5168);
nor U12045 (N_12045,N_5263,N_7780);
and U12046 (N_12046,N_8813,N_7801);
or U12047 (N_12047,N_6221,N_9357);
nand U12048 (N_12048,N_6836,N_6855);
nand U12049 (N_12049,N_6098,N_8791);
and U12050 (N_12050,N_7539,N_5032);
nor U12051 (N_12051,N_5364,N_8825);
nand U12052 (N_12052,N_8058,N_9417);
nor U12053 (N_12053,N_9925,N_7385);
and U12054 (N_12054,N_9022,N_6037);
or U12055 (N_12055,N_7767,N_9178);
or U12056 (N_12056,N_7483,N_5490);
and U12057 (N_12057,N_9694,N_7463);
and U12058 (N_12058,N_6812,N_9608);
nor U12059 (N_12059,N_8413,N_7581);
and U12060 (N_12060,N_8451,N_9172);
nand U12061 (N_12061,N_7492,N_9046);
and U12062 (N_12062,N_9792,N_6530);
and U12063 (N_12063,N_9945,N_9325);
and U12064 (N_12064,N_6615,N_5470);
nand U12065 (N_12065,N_5923,N_8002);
and U12066 (N_12066,N_8756,N_7596);
nor U12067 (N_12067,N_9683,N_7318);
nor U12068 (N_12068,N_8470,N_9583);
nand U12069 (N_12069,N_5006,N_7376);
nand U12070 (N_12070,N_8878,N_5753);
and U12071 (N_12071,N_6718,N_9490);
and U12072 (N_12072,N_9428,N_5704);
nand U12073 (N_12073,N_5334,N_6205);
or U12074 (N_12074,N_8152,N_9741);
nand U12075 (N_12075,N_6804,N_6055);
or U12076 (N_12076,N_5097,N_5685);
nor U12077 (N_12077,N_6367,N_5610);
or U12078 (N_12078,N_5573,N_6568);
and U12079 (N_12079,N_6808,N_7454);
and U12080 (N_12080,N_7120,N_7877);
or U12081 (N_12081,N_8229,N_9998);
and U12082 (N_12082,N_5253,N_6204);
nand U12083 (N_12083,N_6885,N_9787);
and U12084 (N_12084,N_7043,N_7528);
and U12085 (N_12085,N_9743,N_5764);
or U12086 (N_12086,N_9571,N_9272);
nand U12087 (N_12087,N_5707,N_6645);
nor U12088 (N_12088,N_8795,N_5698);
nor U12089 (N_12089,N_8327,N_6999);
nand U12090 (N_12090,N_8476,N_9795);
or U12091 (N_12091,N_6844,N_9577);
or U12092 (N_12092,N_7759,N_9858);
and U12093 (N_12093,N_7579,N_9891);
and U12094 (N_12094,N_7806,N_6799);
xnor U12095 (N_12095,N_7090,N_5329);
nand U12096 (N_12096,N_7414,N_5538);
nor U12097 (N_12097,N_6178,N_5777);
xor U12098 (N_12098,N_5754,N_5579);
and U12099 (N_12099,N_7353,N_7238);
nor U12100 (N_12100,N_6033,N_9327);
or U12101 (N_12101,N_7162,N_5009);
nor U12102 (N_12102,N_5374,N_9841);
and U12103 (N_12103,N_5501,N_9958);
nor U12104 (N_12104,N_5639,N_9192);
nor U12105 (N_12105,N_5918,N_6333);
and U12106 (N_12106,N_8230,N_5869);
and U12107 (N_12107,N_7948,N_8762);
and U12108 (N_12108,N_5170,N_5700);
nand U12109 (N_12109,N_9897,N_8078);
nand U12110 (N_12110,N_7832,N_6704);
and U12111 (N_12111,N_6600,N_9169);
nand U12112 (N_12112,N_7315,N_7729);
or U12113 (N_12113,N_6801,N_8840);
nor U12114 (N_12114,N_5772,N_5252);
and U12115 (N_12115,N_7074,N_7786);
nand U12116 (N_12116,N_8506,N_6141);
and U12117 (N_12117,N_9650,N_5643);
nor U12118 (N_12118,N_6095,N_9081);
or U12119 (N_12119,N_9626,N_5457);
and U12120 (N_12120,N_5615,N_5668);
or U12121 (N_12121,N_6730,N_6376);
and U12122 (N_12122,N_6391,N_6040);
and U12123 (N_12123,N_9934,N_6578);
and U12124 (N_12124,N_6191,N_7818);
nand U12125 (N_12125,N_8441,N_9143);
or U12126 (N_12126,N_5392,N_9372);
and U12127 (N_12127,N_6955,N_5066);
nand U12128 (N_12128,N_9009,N_7366);
nor U12129 (N_12129,N_8109,N_5499);
or U12130 (N_12130,N_7775,N_5865);
and U12131 (N_12131,N_6236,N_9253);
nand U12132 (N_12132,N_5127,N_5949);
and U12133 (N_12133,N_8591,N_9681);
and U12134 (N_12134,N_8816,N_5526);
or U12135 (N_12135,N_8567,N_8734);
and U12136 (N_12136,N_5703,N_9521);
nand U12137 (N_12137,N_8048,N_7785);
nor U12138 (N_12138,N_5706,N_7975);
nand U12139 (N_12139,N_9701,N_8633);
nand U12140 (N_12140,N_6075,N_7640);
or U12141 (N_12141,N_9200,N_7711);
nand U12142 (N_12142,N_7066,N_8348);
and U12143 (N_12143,N_8093,N_7846);
or U12144 (N_12144,N_7881,N_5126);
or U12145 (N_12145,N_9585,N_5819);
nand U12146 (N_12146,N_9698,N_8235);
and U12147 (N_12147,N_8790,N_7343);
or U12148 (N_12148,N_9654,N_8499);
and U12149 (N_12149,N_5861,N_7412);
nand U12150 (N_12150,N_9935,N_5691);
nand U12151 (N_12151,N_5560,N_6077);
nor U12152 (N_12152,N_8004,N_9151);
and U12153 (N_12153,N_9734,N_5182);
or U12154 (N_12154,N_6786,N_8584);
and U12155 (N_12155,N_6190,N_8365);
nor U12156 (N_12156,N_9268,N_5137);
nand U12157 (N_12157,N_5053,N_6003);
and U12158 (N_12158,N_7051,N_6859);
and U12159 (N_12159,N_6087,N_7000);
nand U12160 (N_12160,N_6850,N_6159);
or U12161 (N_12161,N_6362,N_6252);
or U12162 (N_12162,N_9116,N_6924);
nor U12163 (N_12163,N_9803,N_9630);
and U12164 (N_12164,N_9462,N_8728);
nand U12165 (N_12165,N_6025,N_9675);
and U12166 (N_12166,N_5995,N_7610);
or U12167 (N_12167,N_5756,N_6519);
or U12168 (N_12168,N_9566,N_7811);
nor U12169 (N_12169,N_5654,N_7224);
nor U12170 (N_12170,N_9142,N_9869);
and U12171 (N_12171,N_6223,N_7112);
nor U12172 (N_12172,N_6590,N_8028);
nor U12173 (N_12173,N_8200,N_7425);
or U12174 (N_12174,N_8450,N_6253);
and U12175 (N_12175,N_6092,N_5413);
nand U12176 (N_12176,N_9358,N_7053);
or U12177 (N_12177,N_9589,N_5162);
or U12178 (N_12178,N_5452,N_8699);
nor U12179 (N_12179,N_6051,N_7060);
nand U12180 (N_12180,N_5961,N_9597);
nor U12181 (N_12181,N_6387,N_6862);
or U12182 (N_12182,N_7260,N_8819);
or U12183 (N_12183,N_8399,N_6501);
nand U12184 (N_12184,N_5186,N_8113);
nor U12185 (N_12185,N_8969,N_9708);
or U12186 (N_12186,N_9880,N_5318);
or U12187 (N_12187,N_6414,N_9952);
or U12188 (N_12188,N_7453,N_6280);
nand U12189 (N_12189,N_8100,N_6117);
nand U12190 (N_12190,N_6115,N_5175);
or U12191 (N_12191,N_6597,N_5512);
nor U12192 (N_12192,N_9383,N_8263);
nor U12193 (N_12193,N_6906,N_5321);
xnor U12194 (N_12194,N_5409,N_5315);
or U12195 (N_12195,N_7160,N_8201);
nand U12196 (N_12196,N_8900,N_9757);
or U12197 (N_12197,N_9999,N_9556);
nand U12198 (N_12198,N_9119,N_7277);
and U12199 (N_12199,N_8688,N_5086);
and U12200 (N_12200,N_8123,N_5793);
nor U12201 (N_12201,N_8611,N_9828);
or U12202 (N_12202,N_5575,N_8725);
nand U12203 (N_12203,N_9302,N_7739);
or U12204 (N_12204,N_5402,N_7595);
nor U12205 (N_12205,N_9130,N_8803);
nand U12206 (N_12206,N_5494,N_9155);
and U12207 (N_12207,N_7829,N_8380);
nand U12208 (N_12208,N_5273,N_9454);
nor U12209 (N_12209,N_7559,N_5633);
nor U12210 (N_12210,N_7261,N_9269);
nor U12211 (N_12211,N_6584,N_6567);
and U12212 (N_12212,N_5307,N_9961);
or U12213 (N_12213,N_6963,N_6677);
nor U12214 (N_12214,N_6008,N_9629);
and U12215 (N_12215,N_6979,N_7430);
nor U12216 (N_12216,N_9170,N_6880);
nor U12217 (N_12217,N_6011,N_9550);
and U12218 (N_12218,N_6605,N_6138);
and U12219 (N_12219,N_8547,N_9627);
nor U12220 (N_12220,N_5148,N_6332);
and U12221 (N_12221,N_5047,N_6009);
nand U12222 (N_12222,N_8845,N_7690);
nand U12223 (N_12223,N_8285,N_9011);
nand U12224 (N_12224,N_6723,N_6531);
or U12225 (N_12225,N_6231,N_9498);
nand U12226 (N_12226,N_6153,N_8659);
or U12227 (N_12227,N_5365,N_8092);
nor U12228 (N_12228,N_8343,N_6375);
and U12229 (N_12229,N_6064,N_8359);
or U12230 (N_12230,N_6640,N_7326);
nand U12231 (N_12231,N_6305,N_8146);
and U12232 (N_12232,N_9301,N_8321);
or U12233 (N_12233,N_9097,N_5833);
nand U12234 (N_12234,N_9746,N_8690);
nand U12235 (N_12235,N_9712,N_8903);
or U12236 (N_12236,N_8317,N_5135);
nor U12237 (N_12237,N_9286,N_8238);
or U12238 (N_12238,N_7025,N_6397);
nand U12239 (N_12239,N_5750,N_6575);
or U12240 (N_12240,N_8086,N_9581);
nand U12241 (N_12241,N_7899,N_6462);
and U12242 (N_12242,N_6699,N_8517);
and U12243 (N_12243,N_6527,N_6422);
or U12244 (N_12244,N_5225,N_6598);
and U12245 (N_12245,N_6612,N_6409);
or U12246 (N_12246,N_8105,N_9371);
and U12247 (N_12247,N_8324,N_8532);
nor U12248 (N_12248,N_8260,N_7737);
or U12249 (N_12249,N_8904,N_5415);
or U12250 (N_12250,N_6570,N_6483);
nand U12251 (N_12251,N_7660,N_9362);
or U12252 (N_12252,N_6663,N_5791);
nand U12253 (N_12253,N_6676,N_6134);
nor U12254 (N_12254,N_7132,N_9928);
and U12255 (N_12255,N_9247,N_8604);
nand U12256 (N_12256,N_6806,N_8723);
nand U12257 (N_12257,N_5800,N_8388);
or U12258 (N_12258,N_6780,N_6541);
nor U12259 (N_12259,N_8781,N_8511);
and U12260 (N_12260,N_9816,N_5768);
or U12261 (N_12261,N_8907,N_8873);
nand U12262 (N_12262,N_7749,N_7673);
nor U12263 (N_12263,N_7474,N_6762);
and U12264 (N_12264,N_9396,N_6321);
and U12265 (N_12265,N_5125,N_7851);
or U12266 (N_12266,N_8914,N_5239);
nand U12267 (N_12267,N_7222,N_7370);
nor U12268 (N_12268,N_6200,N_5429);
nor U12269 (N_12269,N_5295,N_5157);
or U12270 (N_12270,N_6343,N_8477);
nand U12271 (N_12271,N_6959,N_9714);
or U12272 (N_12272,N_8387,N_8631);
or U12273 (N_12273,N_6549,N_7638);
nor U12274 (N_12274,N_9213,N_8513);
or U12275 (N_12275,N_6218,N_5447);
and U12276 (N_12276,N_8295,N_9341);
nand U12277 (N_12277,N_5749,N_8622);
and U12278 (N_12278,N_7788,N_5231);
nand U12279 (N_12279,N_7328,N_6637);
nand U12280 (N_12280,N_5870,N_8812);
or U12281 (N_12281,N_6502,N_9425);
nor U12282 (N_12282,N_5181,N_5353);
and U12283 (N_12283,N_6140,N_8030);
nor U12284 (N_12284,N_9197,N_6657);
and U12285 (N_12285,N_8011,N_5482);
or U12286 (N_12286,N_8862,N_8261);
and U12287 (N_12287,N_8121,N_5779);
nand U12288 (N_12288,N_5766,N_6460);
or U12289 (N_12289,N_9104,N_9246);
or U12290 (N_12290,N_7997,N_5929);
nand U12291 (N_12291,N_8656,N_8752);
or U12292 (N_12292,N_6853,N_6993);
nor U12293 (N_12293,N_9068,N_6989);
or U12294 (N_12294,N_6540,N_9069);
or U12295 (N_12295,N_8692,N_8706);
nand U12296 (N_12296,N_7631,N_5096);
and U12297 (N_12297,N_8518,N_7035);
and U12298 (N_12298,N_6005,N_6405);
nand U12299 (N_12299,N_8701,N_6681);
nand U12300 (N_12300,N_5249,N_9293);
nand U12301 (N_12301,N_8988,N_8408);
nor U12302 (N_12302,N_8205,N_9920);
and U12303 (N_12303,N_6639,N_8162);
or U12304 (N_12304,N_6181,N_5480);
or U12305 (N_12305,N_6355,N_6069);
or U12306 (N_12306,N_7065,N_9368);
or U12307 (N_12307,N_7329,N_9976);
and U12308 (N_12308,N_8596,N_6868);
and U12309 (N_12309,N_9296,N_5845);
nand U12310 (N_12310,N_6751,N_9048);
nor U12311 (N_12311,N_6233,N_6254);
or U12312 (N_12312,N_8678,N_5722);
nand U12313 (N_12313,N_8473,N_6542);
nor U12314 (N_12314,N_8138,N_9274);
nor U12315 (N_12315,N_9532,N_9797);
and U12316 (N_12316,N_6160,N_5078);
and U12317 (N_12317,N_9833,N_5316);
or U12318 (N_12318,N_5875,N_7470);
or U12319 (N_12319,N_7625,N_8571);
nor U12320 (N_12320,N_6302,N_8740);
and U12321 (N_12321,N_6339,N_6059);
and U12322 (N_12322,N_9079,N_6917);
nand U12323 (N_12323,N_5730,N_7011);
nand U12324 (N_12324,N_9404,N_9824);
and U12325 (N_12325,N_8223,N_8322);
and U12326 (N_12326,N_9898,N_8603);
and U12327 (N_12327,N_7330,N_9994);
or U12328 (N_12328,N_7557,N_7794);
or U12329 (N_12329,N_7696,N_6356);
nor U12330 (N_12330,N_9834,N_8880);
or U12331 (N_12331,N_9458,N_9611);
or U12332 (N_12332,N_8220,N_6500);
nor U12333 (N_12333,N_7777,N_5594);
nand U12334 (N_12334,N_5199,N_6464);
nand U12335 (N_12335,N_9047,N_9158);
or U12336 (N_12336,N_6109,N_9548);
nand U12337 (N_12337,N_9965,N_9354);
or U12338 (N_12338,N_7655,N_8826);
or U12339 (N_12339,N_9579,N_8405);
and U12340 (N_12340,N_6112,N_6616);
or U12341 (N_12341,N_9867,N_6324);
or U12342 (N_12342,N_5313,N_8664);
or U12343 (N_12343,N_5145,N_8502);
or U12344 (N_12344,N_6449,N_9599);
nor U12345 (N_12345,N_7594,N_5678);
and U12346 (N_12346,N_5102,N_8866);
and U12347 (N_12347,N_5323,N_6895);
nor U12348 (N_12348,N_5956,N_7475);
nor U12349 (N_12349,N_5635,N_8389);
nor U12350 (N_12350,N_8351,N_8858);
or U12351 (N_12351,N_8857,N_7573);
nor U12352 (N_12352,N_7005,N_8097);
nor U12353 (N_12353,N_8257,N_9252);
nor U12354 (N_12354,N_7230,N_9639);
nand U12355 (N_12355,N_9165,N_9102);
and U12356 (N_12356,N_7646,N_9941);
nand U12357 (N_12357,N_7346,N_7107);
nand U12358 (N_12358,N_9096,N_9874);
or U12359 (N_12359,N_5797,N_9593);
nor U12360 (N_12360,N_9864,N_9622);
and U12361 (N_12361,N_8764,N_6023);
nor U12362 (N_12362,N_6350,N_7902);
nand U12363 (N_12363,N_6717,N_6523);
nand U12364 (N_12364,N_9064,N_6045);
nor U12365 (N_12365,N_5690,N_9805);
and U12366 (N_12366,N_5178,N_7602);
nand U12367 (N_12367,N_8619,N_9722);
nor U12368 (N_12368,N_9052,N_7915);
or U12369 (N_12369,N_9590,N_5497);
nor U12370 (N_12370,N_5919,N_5781);
nor U12371 (N_12371,N_6016,N_6208);
or U12372 (N_12372,N_5292,N_5358);
nand U12373 (N_12373,N_9917,N_7467);
nor U12374 (N_12374,N_7658,N_8954);
and U12375 (N_12375,N_7771,N_7593);
nand U12376 (N_12376,N_5088,N_6967);
nor U12377 (N_12377,N_6213,N_5204);
or U12378 (N_12378,N_7464,N_8573);
or U12379 (N_12379,N_8489,N_9120);
or U12380 (N_12380,N_9924,N_5130);
and U12381 (N_12381,N_7917,N_5977);
nor U12382 (N_12382,N_5132,N_7795);
or U12383 (N_12383,N_6886,N_9284);
nand U12384 (N_12384,N_5636,N_7028);
and U12385 (N_12385,N_7141,N_8841);
and U12386 (N_12386,N_7861,N_6889);
xor U12387 (N_12387,N_9334,N_9226);
xnor U12388 (N_12388,N_7663,N_7374);
and U12389 (N_12389,N_9883,N_9907);
or U12390 (N_12390,N_6149,N_5537);
and U12391 (N_12391,N_6042,N_8755);
or U12392 (N_12392,N_8496,N_8569);
or U12393 (N_12393,N_8107,N_5561);
nor U12394 (N_12394,N_6086,N_9111);
nand U12395 (N_12395,N_5883,N_8118);
nand U12396 (N_12396,N_8175,N_5802);
nor U12397 (N_12397,N_8695,N_9836);
nand U12398 (N_12398,N_9818,N_8057);
or U12399 (N_12399,N_7259,N_9922);
or U12400 (N_12400,N_9724,N_6891);
or U12401 (N_12401,N_5308,N_5400);
and U12402 (N_12402,N_9567,N_5031);
or U12403 (N_12403,N_9514,N_5564);
nand U12404 (N_12404,N_6988,N_6514);
nor U12405 (N_12405,N_8651,N_7882);
and U12406 (N_12406,N_6102,N_9308);
or U12407 (N_12407,N_7874,N_6543);
nor U12408 (N_12408,N_9254,N_6588);
and U12409 (N_12409,N_6720,N_6101);
and U12410 (N_12410,N_6484,N_5453);
nor U12411 (N_12411,N_5389,N_7954);
and U12412 (N_12412,N_9114,N_6586);
and U12413 (N_12413,N_8457,N_5007);
or U12414 (N_12414,N_8844,N_7680);
nand U12415 (N_12415,N_9559,N_6820);
or U12416 (N_12416,N_7383,N_7294);
or U12417 (N_12417,N_9359,N_9098);
and U12418 (N_12418,N_9844,N_5701);
nor U12419 (N_12419,N_5775,N_9885);
nor U12420 (N_12420,N_8115,N_7910);
nor U12421 (N_12421,N_8159,N_8339);
nand U12422 (N_12422,N_6707,N_5632);
nor U12423 (N_12423,N_9389,N_8964);
nand U12424 (N_12424,N_8291,N_8415);
nand U12425 (N_12425,N_5274,N_9324);
and U12426 (N_12426,N_7962,N_9677);
or U12427 (N_12427,N_8549,N_7591);
and U12428 (N_12428,N_7816,N_6722);
nor U12429 (N_12429,N_6320,N_7348);
nand U12430 (N_12430,N_9602,N_9124);
or U12431 (N_12431,N_7510,N_5438);
and U12432 (N_12432,N_5829,N_8170);
nand U12433 (N_12433,N_6061,N_7664);
nand U12434 (N_12434,N_9947,N_8455);
nand U12435 (N_12435,N_6212,N_5154);
and U12436 (N_12436,N_9031,N_7503);
nand U12437 (N_12437,N_9220,N_9393);
nand U12438 (N_12438,N_6340,N_5840);
and U12439 (N_12439,N_5027,N_7688);
and U12440 (N_12440,N_8370,N_5474);
and U12441 (N_12441,N_8110,N_5987);
nand U12442 (N_12442,N_7833,N_8737);
nor U12443 (N_12443,N_9108,N_6293);
nand U12444 (N_12444,N_9685,N_5351);
nand U12445 (N_12445,N_6760,N_7231);
or U12446 (N_12446,N_7708,N_6261);
nand U12447 (N_12447,N_5233,N_8708);
and U12448 (N_12448,N_9276,N_5173);
or U12449 (N_12449,N_6670,N_7305);
nor U12450 (N_12450,N_9866,N_5586);
nand U12451 (N_12451,N_9277,N_6922);
nor U12452 (N_12452,N_8462,N_8102);
or U12453 (N_12453,N_6228,N_7400);
and U12454 (N_12454,N_6085,N_9085);
nand U12455 (N_12455,N_5528,N_7395);
and U12456 (N_12456,N_7947,N_7970);
and U12457 (N_12457,N_6026,N_7754);
or U12458 (N_12458,N_7783,N_8158);
or U12459 (N_12459,N_6761,N_7102);
nor U12460 (N_12460,N_7013,N_6019);
nand U12461 (N_12461,N_9552,N_5104);
nand U12462 (N_12462,N_8340,N_7418);
or U12463 (N_12463,N_8061,N_6251);
and U12464 (N_12464,N_9684,N_8401);
nand U12465 (N_12465,N_7397,N_6491);
or U12466 (N_12466,N_9700,N_9495);
nand U12467 (N_12467,N_9199,N_9725);
nor U12468 (N_12468,N_7978,N_6472);
or U12469 (N_12469,N_8460,N_5449);
or U12470 (N_12470,N_6511,N_9162);
nand U12471 (N_12471,N_6119,N_9950);
nor U12472 (N_12472,N_8400,N_9369);
nand U12473 (N_12473,N_9704,N_5368);
nand U12474 (N_12474,N_9150,N_5640);
or U12475 (N_12475,N_7955,N_8378);
and U12476 (N_12476,N_6177,N_7488);
nand U12477 (N_12477,N_8318,N_5340);
or U12478 (N_12478,N_7427,N_5428);
nor U12479 (N_12479,N_6555,N_9955);
nand U12480 (N_12480,N_7350,N_8044);
and U12481 (N_12481,N_6983,N_8693);
or U12482 (N_12482,N_8385,N_7283);
or U12483 (N_12483,N_5943,N_5931);
nor U12484 (N_12484,N_5229,N_8921);
and U12485 (N_12485,N_7823,N_6383);
nand U12486 (N_12486,N_9279,N_7950);
nand U12487 (N_12487,N_5859,N_8823);
nand U12488 (N_12488,N_9432,N_9442);
or U12489 (N_12489,N_8955,N_7306);
and U12490 (N_12490,N_9975,N_7924);
or U12491 (N_12491,N_6331,N_6990);
nand U12492 (N_12492,N_6067,N_7695);
and U12493 (N_12493,N_8846,N_6687);
or U12494 (N_12494,N_5911,N_7122);
and U12495 (N_12495,N_7883,N_6601);
or U12496 (N_12496,N_6667,N_9026);
nor U12497 (N_12497,N_8733,N_9916);
nor U12498 (N_12498,N_5942,N_8426);
nor U12499 (N_12499,N_8018,N_6528);
or U12500 (N_12500,N_8551,N_8109);
and U12501 (N_12501,N_6770,N_9117);
nand U12502 (N_12502,N_7182,N_8111);
nor U12503 (N_12503,N_5339,N_5111);
nand U12504 (N_12504,N_5587,N_9504);
nor U12505 (N_12505,N_8195,N_9474);
and U12506 (N_12506,N_8808,N_5831);
and U12507 (N_12507,N_5907,N_6109);
nand U12508 (N_12508,N_5624,N_7188);
nor U12509 (N_12509,N_5776,N_6631);
and U12510 (N_12510,N_6044,N_9283);
nand U12511 (N_12511,N_9728,N_9618);
nor U12512 (N_12512,N_6059,N_8065);
and U12513 (N_12513,N_9002,N_6379);
nand U12514 (N_12514,N_5862,N_5108);
and U12515 (N_12515,N_9478,N_5394);
nor U12516 (N_12516,N_6232,N_6414);
and U12517 (N_12517,N_6726,N_8742);
or U12518 (N_12518,N_7916,N_5488);
nor U12519 (N_12519,N_5071,N_9690);
and U12520 (N_12520,N_9999,N_6260);
nand U12521 (N_12521,N_5350,N_7741);
nand U12522 (N_12522,N_5381,N_8639);
or U12523 (N_12523,N_9210,N_9436);
or U12524 (N_12524,N_9888,N_7164);
or U12525 (N_12525,N_8631,N_6712);
nand U12526 (N_12526,N_9767,N_5309);
nor U12527 (N_12527,N_9801,N_9299);
or U12528 (N_12528,N_5924,N_8747);
nor U12529 (N_12529,N_6333,N_8249);
or U12530 (N_12530,N_6320,N_9410);
nor U12531 (N_12531,N_8063,N_7594);
and U12532 (N_12532,N_9975,N_5988);
or U12533 (N_12533,N_5980,N_5651);
nor U12534 (N_12534,N_6648,N_8813);
nand U12535 (N_12535,N_7531,N_6168);
nor U12536 (N_12536,N_9751,N_6480);
nor U12537 (N_12537,N_5123,N_9132);
nand U12538 (N_12538,N_6282,N_7798);
or U12539 (N_12539,N_6018,N_8061);
nand U12540 (N_12540,N_9647,N_8595);
and U12541 (N_12541,N_9195,N_9058);
nand U12542 (N_12542,N_9785,N_9658);
nor U12543 (N_12543,N_6433,N_8551);
nand U12544 (N_12544,N_5143,N_5259);
or U12545 (N_12545,N_7230,N_9758);
or U12546 (N_12546,N_7756,N_7795);
nand U12547 (N_12547,N_9781,N_6340);
and U12548 (N_12548,N_5227,N_6315);
and U12549 (N_12549,N_5965,N_5258);
or U12550 (N_12550,N_5919,N_9423);
nand U12551 (N_12551,N_9514,N_8309);
or U12552 (N_12552,N_7981,N_5821);
or U12553 (N_12553,N_8237,N_9843);
nand U12554 (N_12554,N_8961,N_9856);
nor U12555 (N_12555,N_8361,N_9350);
or U12556 (N_12556,N_6767,N_9542);
nor U12557 (N_12557,N_6603,N_8793);
nor U12558 (N_12558,N_5391,N_6715);
nand U12559 (N_12559,N_7119,N_9844);
nand U12560 (N_12560,N_6089,N_9714);
nor U12561 (N_12561,N_9182,N_9611);
or U12562 (N_12562,N_5395,N_5808);
or U12563 (N_12563,N_6786,N_9517);
or U12564 (N_12564,N_8802,N_7654);
nand U12565 (N_12565,N_5799,N_6875);
and U12566 (N_12566,N_9951,N_5662);
or U12567 (N_12567,N_6851,N_9113);
nor U12568 (N_12568,N_7699,N_7695);
nor U12569 (N_12569,N_5107,N_6519);
nor U12570 (N_12570,N_5054,N_8352);
or U12571 (N_12571,N_6008,N_5005);
nor U12572 (N_12572,N_5290,N_7879);
nor U12573 (N_12573,N_9783,N_5361);
nand U12574 (N_12574,N_6317,N_8013);
nand U12575 (N_12575,N_7636,N_7904);
or U12576 (N_12576,N_7858,N_8946);
nor U12577 (N_12577,N_9726,N_5381);
or U12578 (N_12578,N_5759,N_6826);
or U12579 (N_12579,N_8286,N_7185);
nor U12580 (N_12580,N_8894,N_6164);
nand U12581 (N_12581,N_5264,N_6057);
and U12582 (N_12582,N_6129,N_5409);
and U12583 (N_12583,N_5513,N_5245);
nor U12584 (N_12584,N_6432,N_8039);
or U12585 (N_12585,N_7083,N_5951);
and U12586 (N_12586,N_6817,N_9967);
nor U12587 (N_12587,N_6945,N_5121);
nand U12588 (N_12588,N_7642,N_6403);
nand U12589 (N_12589,N_5539,N_5786);
nor U12590 (N_12590,N_5367,N_5598);
or U12591 (N_12591,N_7440,N_5632);
and U12592 (N_12592,N_5875,N_8903);
and U12593 (N_12593,N_9068,N_9010);
and U12594 (N_12594,N_5500,N_8393);
nor U12595 (N_12595,N_5790,N_5327);
or U12596 (N_12596,N_8501,N_6991);
or U12597 (N_12597,N_5932,N_5249);
nand U12598 (N_12598,N_9084,N_5473);
nand U12599 (N_12599,N_5180,N_6403);
nand U12600 (N_12600,N_6610,N_9506);
nor U12601 (N_12601,N_7846,N_7245);
or U12602 (N_12602,N_8419,N_5626);
or U12603 (N_12603,N_7892,N_8099);
nand U12604 (N_12604,N_9477,N_8152);
nand U12605 (N_12605,N_6884,N_6660);
nand U12606 (N_12606,N_5112,N_7660);
or U12607 (N_12607,N_5704,N_5121);
nor U12608 (N_12608,N_6074,N_8085);
and U12609 (N_12609,N_7532,N_6931);
nand U12610 (N_12610,N_8919,N_7518);
nand U12611 (N_12611,N_9678,N_7771);
nor U12612 (N_12612,N_9427,N_8231);
or U12613 (N_12613,N_8661,N_6218);
or U12614 (N_12614,N_9752,N_8370);
nand U12615 (N_12615,N_7187,N_6647);
and U12616 (N_12616,N_5257,N_6224);
and U12617 (N_12617,N_7995,N_7856);
and U12618 (N_12618,N_5398,N_6191);
nor U12619 (N_12619,N_8235,N_8179);
and U12620 (N_12620,N_5114,N_6626);
nor U12621 (N_12621,N_8265,N_6134);
nor U12622 (N_12622,N_9521,N_9152);
nand U12623 (N_12623,N_9277,N_6200);
nand U12624 (N_12624,N_9946,N_8337);
and U12625 (N_12625,N_6385,N_6296);
nor U12626 (N_12626,N_5443,N_5127);
or U12627 (N_12627,N_5307,N_8286);
nand U12628 (N_12628,N_7341,N_9502);
nor U12629 (N_12629,N_8033,N_7318);
and U12630 (N_12630,N_8286,N_9033);
or U12631 (N_12631,N_5721,N_6643);
nor U12632 (N_12632,N_8295,N_9068);
nand U12633 (N_12633,N_9237,N_9563);
nor U12634 (N_12634,N_6228,N_5043);
or U12635 (N_12635,N_8964,N_7506);
or U12636 (N_12636,N_8829,N_5537);
or U12637 (N_12637,N_7843,N_8968);
nand U12638 (N_12638,N_7984,N_9257);
or U12639 (N_12639,N_8828,N_6717);
and U12640 (N_12640,N_6994,N_9960);
or U12641 (N_12641,N_5231,N_7291);
or U12642 (N_12642,N_9873,N_7671);
nand U12643 (N_12643,N_8126,N_7192);
or U12644 (N_12644,N_5792,N_9861);
and U12645 (N_12645,N_7806,N_5936);
nand U12646 (N_12646,N_6423,N_6113);
nand U12647 (N_12647,N_7638,N_7738);
nand U12648 (N_12648,N_6323,N_9841);
or U12649 (N_12649,N_6052,N_5248);
nand U12650 (N_12650,N_5004,N_7605);
or U12651 (N_12651,N_6663,N_6363);
nor U12652 (N_12652,N_6579,N_6059);
xor U12653 (N_12653,N_7657,N_9503);
nor U12654 (N_12654,N_6382,N_7914);
or U12655 (N_12655,N_8361,N_9623);
or U12656 (N_12656,N_7860,N_9665);
nor U12657 (N_12657,N_6823,N_8000);
nand U12658 (N_12658,N_9533,N_5763);
or U12659 (N_12659,N_6601,N_7681);
nand U12660 (N_12660,N_7202,N_7200);
nor U12661 (N_12661,N_8103,N_5817);
or U12662 (N_12662,N_9169,N_6020);
nand U12663 (N_12663,N_7343,N_8428);
nand U12664 (N_12664,N_8917,N_9130);
or U12665 (N_12665,N_9255,N_7327);
nand U12666 (N_12666,N_5154,N_5560);
and U12667 (N_12667,N_5309,N_5750);
nand U12668 (N_12668,N_9131,N_8664);
and U12669 (N_12669,N_6976,N_7850);
nor U12670 (N_12670,N_8757,N_5423);
and U12671 (N_12671,N_7202,N_6586);
and U12672 (N_12672,N_7106,N_8535);
and U12673 (N_12673,N_7337,N_5144);
nor U12674 (N_12674,N_7183,N_6124);
nor U12675 (N_12675,N_9736,N_5080);
or U12676 (N_12676,N_7160,N_8520);
nor U12677 (N_12677,N_5568,N_7595);
and U12678 (N_12678,N_8311,N_6526);
nand U12679 (N_12679,N_5415,N_7509);
or U12680 (N_12680,N_9257,N_8800);
nor U12681 (N_12681,N_7619,N_5607);
and U12682 (N_12682,N_7623,N_7989);
and U12683 (N_12683,N_5283,N_5425);
or U12684 (N_12684,N_5603,N_7019);
and U12685 (N_12685,N_6122,N_5195);
nand U12686 (N_12686,N_5749,N_7066);
or U12687 (N_12687,N_8385,N_8268);
or U12688 (N_12688,N_8866,N_5654);
or U12689 (N_12689,N_9215,N_5269);
nand U12690 (N_12690,N_8308,N_9851);
nand U12691 (N_12691,N_6109,N_7058);
nand U12692 (N_12692,N_7246,N_7985);
and U12693 (N_12693,N_9340,N_5023);
or U12694 (N_12694,N_5077,N_9060);
nor U12695 (N_12695,N_9992,N_6068);
xor U12696 (N_12696,N_8615,N_9994);
nand U12697 (N_12697,N_7741,N_7050);
and U12698 (N_12698,N_9163,N_9072);
and U12699 (N_12699,N_9884,N_5744);
and U12700 (N_12700,N_9472,N_6303);
nand U12701 (N_12701,N_6667,N_8306);
nor U12702 (N_12702,N_5263,N_6922);
nor U12703 (N_12703,N_6583,N_7375);
and U12704 (N_12704,N_8452,N_7446);
nor U12705 (N_12705,N_5619,N_6759);
and U12706 (N_12706,N_7201,N_5289);
or U12707 (N_12707,N_9498,N_5179);
nor U12708 (N_12708,N_7769,N_5234);
nor U12709 (N_12709,N_8293,N_7324);
nand U12710 (N_12710,N_6909,N_9012);
nand U12711 (N_12711,N_9041,N_9222);
and U12712 (N_12712,N_7886,N_7787);
or U12713 (N_12713,N_9311,N_6881);
and U12714 (N_12714,N_9422,N_7047);
and U12715 (N_12715,N_8651,N_9519);
and U12716 (N_12716,N_6301,N_6229);
and U12717 (N_12717,N_8815,N_6560);
nor U12718 (N_12718,N_7924,N_7988);
or U12719 (N_12719,N_8599,N_9179);
and U12720 (N_12720,N_8388,N_7078);
and U12721 (N_12721,N_8335,N_8893);
or U12722 (N_12722,N_8027,N_7764);
or U12723 (N_12723,N_6869,N_5035);
nor U12724 (N_12724,N_5590,N_6759);
or U12725 (N_12725,N_9381,N_8757);
or U12726 (N_12726,N_5026,N_6958);
or U12727 (N_12727,N_7027,N_5567);
or U12728 (N_12728,N_8568,N_6774);
nor U12729 (N_12729,N_8708,N_5606);
nand U12730 (N_12730,N_7308,N_8192);
and U12731 (N_12731,N_8636,N_9041);
nor U12732 (N_12732,N_8069,N_5459);
nor U12733 (N_12733,N_6257,N_6180);
nand U12734 (N_12734,N_8537,N_6962);
or U12735 (N_12735,N_9123,N_6239);
and U12736 (N_12736,N_6770,N_5800);
nor U12737 (N_12737,N_7578,N_8869);
nor U12738 (N_12738,N_7632,N_7562);
and U12739 (N_12739,N_5067,N_7086);
nand U12740 (N_12740,N_8684,N_7162);
and U12741 (N_12741,N_8961,N_6098);
nand U12742 (N_12742,N_9279,N_9228);
or U12743 (N_12743,N_5434,N_6848);
and U12744 (N_12744,N_9635,N_6471);
nand U12745 (N_12745,N_7148,N_5418);
xor U12746 (N_12746,N_9065,N_7779);
nand U12747 (N_12747,N_6468,N_7037);
or U12748 (N_12748,N_8160,N_5137);
and U12749 (N_12749,N_7199,N_6105);
nand U12750 (N_12750,N_6239,N_6103);
nor U12751 (N_12751,N_5026,N_7243);
nand U12752 (N_12752,N_8155,N_7020);
and U12753 (N_12753,N_8352,N_5477);
nor U12754 (N_12754,N_8420,N_9499);
or U12755 (N_12755,N_8679,N_8017);
or U12756 (N_12756,N_9544,N_9055);
nor U12757 (N_12757,N_5600,N_7083);
nand U12758 (N_12758,N_7301,N_7941);
or U12759 (N_12759,N_5088,N_7265);
and U12760 (N_12760,N_9913,N_9339);
or U12761 (N_12761,N_6218,N_6847);
nand U12762 (N_12762,N_7657,N_6547);
nor U12763 (N_12763,N_7725,N_8660);
and U12764 (N_12764,N_6244,N_7335);
or U12765 (N_12765,N_6293,N_8410);
or U12766 (N_12766,N_7544,N_6631);
and U12767 (N_12767,N_6560,N_6714);
nand U12768 (N_12768,N_9556,N_8597);
and U12769 (N_12769,N_9621,N_9422);
nand U12770 (N_12770,N_7746,N_6894);
nor U12771 (N_12771,N_7132,N_5174);
nor U12772 (N_12772,N_7238,N_5432);
nor U12773 (N_12773,N_5014,N_5254);
nor U12774 (N_12774,N_5919,N_8588);
nand U12775 (N_12775,N_9467,N_5954);
nand U12776 (N_12776,N_6941,N_8916);
and U12777 (N_12777,N_8279,N_6787);
nor U12778 (N_12778,N_7167,N_6511);
or U12779 (N_12779,N_8631,N_6659);
nand U12780 (N_12780,N_8416,N_5320);
nor U12781 (N_12781,N_9056,N_6438);
and U12782 (N_12782,N_8830,N_8502);
and U12783 (N_12783,N_9984,N_9639);
and U12784 (N_12784,N_7606,N_9586);
and U12785 (N_12785,N_5587,N_5131);
and U12786 (N_12786,N_9594,N_8617);
or U12787 (N_12787,N_9901,N_6708);
nand U12788 (N_12788,N_6243,N_8277);
or U12789 (N_12789,N_5626,N_9026);
and U12790 (N_12790,N_6854,N_9583);
and U12791 (N_12791,N_6143,N_7919);
nand U12792 (N_12792,N_6440,N_5805);
nor U12793 (N_12793,N_9458,N_7275);
or U12794 (N_12794,N_5154,N_9373);
nor U12795 (N_12795,N_5282,N_9264);
or U12796 (N_12796,N_7085,N_5848);
nand U12797 (N_12797,N_8183,N_7240);
nand U12798 (N_12798,N_6590,N_5714);
or U12799 (N_12799,N_7043,N_5480);
xor U12800 (N_12800,N_9741,N_9050);
or U12801 (N_12801,N_9831,N_8484);
and U12802 (N_12802,N_6031,N_9499);
and U12803 (N_12803,N_9573,N_6553);
and U12804 (N_12804,N_8189,N_7126);
and U12805 (N_12805,N_7071,N_5303);
and U12806 (N_12806,N_6151,N_5531);
nor U12807 (N_12807,N_7407,N_9540);
nand U12808 (N_12808,N_9851,N_5814);
or U12809 (N_12809,N_8690,N_8515);
nand U12810 (N_12810,N_9757,N_8385);
or U12811 (N_12811,N_5772,N_7200);
nor U12812 (N_12812,N_8462,N_6923);
nand U12813 (N_12813,N_6043,N_7512);
nor U12814 (N_12814,N_9550,N_5907);
and U12815 (N_12815,N_5104,N_5871);
and U12816 (N_12816,N_6589,N_9280);
nor U12817 (N_12817,N_9368,N_7411);
nor U12818 (N_12818,N_7490,N_8690);
nand U12819 (N_12819,N_8408,N_5671);
nor U12820 (N_12820,N_8676,N_8978);
or U12821 (N_12821,N_9001,N_8218);
nand U12822 (N_12822,N_8995,N_8999);
nor U12823 (N_12823,N_8357,N_8328);
or U12824 (N_12824,N_8181,N_8626);
nor U12825 (N_12825,N_6088,N_5660);
or U12826 (N_12826,N_8387,N_9295);
or U12827 (N_12827,N_5806,N_7557);
nor U12828 (N_12828,N_8940,N_7491);
nor U12829 (N_12829,N_9048,N_9330);
and U12830 (N_12830,N_8124,N_8982);
nor U12831 (N_12831,N_9107,N_6020);
nand U12832 (N_12832,N_7443,N_7834);
nor U12833 (N_12833,N_7473,N_5998);
and U12834 (N_12834,N_6331,N_7824);
nand U12835 (N_12835,N_6126,N_5634);
and U12836 (N_12836,N_7497,N_8293);
nand U12837 (N_12837,N_9698,N_6331);
and U12838 (N_12838,N_6365,N_8412);
or U12839 (N_12839,N_8935,N_7736);
and U12840 (N_12840,N_7126,N_5247);
nor U12841 (N_12841,N_6198,N_7539);
nand U12842 (N_12842,N_5822,N_5278);
and U12843 (N_12843,N_6294,N_5638);
nor U12844 (N_12844,N_5019,N_8213);
nor U12845 (N_12845,N_7224,N_8878);
or U12846 (N_12846,N_8719,N_6771);
or U12847 (N_12847,N_9588,N_7441);
or U12848 (N_12848,N_7582,N_9717);
nand U12849 (N_12849,N_5347,N_7146);
nor U12850 (N_12850,N_5631,N_7850);
nor U12851 (N_12851,N_8491,N_5941);
or U12852 (N_12852,N_7524,N_8242);
or U12853 (N_12853,N_5912,N_7364);
nand U12854 (N_12854,N_9510,N_6855);
or U12855 (N_12855,N_6256,N_5327);
nand U12856 (N_12856,N_8786,N_6987);
or U12857 (N_12857,N_9855,N_5367);
nor U12858 (N_12858,N_8794,N_9831);
and U12859 (N_12859,N_8874,N_6147);
nor U12860 (N_12860,N_5995,N_5678);
and U12861 (N_12861,N_8469,N_5591);
and U12862 (N_12862,N_8953,N_7152);
and U12863 (N_12863,N_8166,N_5971);
or U12864 (N_12864,N_5135,N_6542);
nor U12865 (N_12865,N_6846,N_9071);
nand U12866 (N_12866,N_7963,N_5263);
nand U12867 (N_12867,N_6512,N_8245);
and U12868 (N_12868,N_7631,N_7867);
or U12869 (N_12869,N_9853,N_7131);
nor U12870 (N_12870,N_6548,N_9951);
or U12871 (N_12871,N_6368,N_7268);
nor U12872 (N_12872,N_6738,N_5238);
or U12873 (N_12873,N_9512,N_9329);
and U12874 (N_12874,N_6655,N_6230);
nand U12875 (N_12875,N_8284,N_6457);
nor U12876 (N_12876,N_8610,N_5338);
or U12877 (N_12877,N_9645,N_9169);
nor U12878 (N_12878,N_5910,N_6071);
nand U12879 (N_12879,N_8422,N_5359);
nor U12880 (N_12880,N_9400,N_7653);
and U12881 (N_12881,N_5730,N_9723);
nand U12882 (N_12882,N_6704,N_8390);
and U12883 (N_12883,N_9907,N_7681);
and U12884 (N_12884,N_6753,N_7520);
and U12885 (N_12885,N_9423,N_8449);
or U12886 (N_12886,N_9951,N_8747);
or U12887 (N_12887,N_6300,N_9366);
nand U12888 (N_12888,N_8759,N_9262);
nor U12889 (N_12889,N_8583,N_9069);
nand U12890 (N_12890,N_7415,N_8411);
nand U12891 (N_12891,N_7428,N_5027);
and U12892 (N_12892,N_6387,N_7617);
or U12893 (N_12893,N_6220,N_7847);
and U12894 (N_12894,N_9559,N_9313);
or U12895 (N_12895,N_5166,N_5513);
nand U12896 (N_12896,N_8938,N_9799);
or U12897 (N_12897,N_5585,N_8556);
nor U12898 (N_12898,N_7226,N_5251);
and U12899 (N_12899,N_6874,N_9684);
and U12900 (N_12900,N_5747,N_9935);
nand U12901 (N_12901,N_9148,N_7715);
nor U12902 (N_12902,N_7174,N_8654);
nand U12903 (N_12903,N_7885,N_8770);
nand U12904 (N_12904,N_7083,N_7793);
nand U12905 (N_12905,N_5959,N_5642);
or U12906 (N_12906,N_5465,N_8931);
xor U12907 (N_12907,N_9779,N_7267);
and U12908 (N_12908,N_6397,N_5107);
or U12909 (N_12909,N_6254,N_6546);
nor U12910 (N_12910,N_7629,N_5906);
and U12911 (N_12911,N_6264,N_5421);
nor U12912 (N_12912,N_9499,N_6959);
nor U12913 (N_12913,N_6216,N_6731);
nand U12914 (N_12914,N_9006,N_8140);
or U12915 (N_12915,N_5085,N_9416);
nand U12916 (N_12916,N_6633,N_9819);
nor U12917 (N_12917,N_5341,N_6818);
nor U12918 (N_12918,N_8372,N_8782);
nor U12919 (N_12919,N_5306,N_6572);
nor U12920 (N_12920,N_6343,N_9544);
or U12921 (N_12921,N_9403,N_5435);
and U12922 (N_12922,N_7339,N_9601);
or U12923 (N_12923,N_8758,N_5480);
and U12924 (N_12924,N_6003,N_7011);
and U12925 (N_12925,N_9873,N_5495);
or U12926 (N_12926,N_7882,N_5821);
xnor U12927 (N_12927,N_9317,N_6713);
nor U12928 (N_12928,N_7858,N_5623);
nor U12929 (N_12929,N_7428,N_6119);
nor U12930 (N_12930,N_5318,N_7212);
nor U12931 (N_12931,N_7923,N_5884);
nor U12932 (N_12932,N_5891,N_7200);
and U12933 (N_12933,N_5473,N_7296);
or U12934 (N_12934,N_9709,N_7860);
nor U12935 (N_12935,N_5949,N_7669);
or U12936 (N_12936,N_6556,N_5043);
nor U12937 (N_12937,N_7060,N_5023);
or U12938 (N_12938,N_6942,N_6033);
or U12939 (N_12939,N_9089,N_6511);
and U12940 (N_12940,N_7489,N_7564);
nand U12941 (N_12941,N_7482,N_6672);
or U12942 (N_12942,N_9561,N_8862);
nand U12943 (N_12943,N_6092,N_5781);
and U12944 (N_12944,N_7759,N_5014);
and U12945 (N_12945,N_5326,N_7672);
nor U12946 (N_12946,N_6138,N_5899);
and U12947 (N_12947,N_5100,N_5737);
or U12948 (N_12948,N_5623,N_7326);
and U12949 (N_12949,N_6821,N_9598);
and U12950 (N_12950,N_7462,N_9096);
nand U12951 (N_12951,N_5771,N_5009);
nand U12952 (N_12952,N_6340,N_6959);
nand U12953 (N_12953,N_8653,N_5025);
or U12954 (N_12954,N_7543,N_9673);
nand U12955 (N_12955,N_6849,N_8375);
and U12956 (N_12956,N_9249,N_5450);
and U12957 (N_12957,N_5294,N_5678);
xnor U12958 (N_12958,N_5743,N_8739);
and U12959 (N_12959,N_9248,N_8836);
and U12960 (N_12960,N_9371,N_9171);
nor U12961 (N_12961,N_9801,N_9447);
and U12962 (N_12962,N_7394,N_9855);
and U12963 (N_12963,N_8441,N_8616);
nand U12964 (N_12964,N_5877,N_8841);
nor U12965 (N_12965,N_8610,N_9124);
nor U12966 (N_12966,N_8696,N_9968);
nor U12967 (N_12967,N_8940,N_9526);
nand U12968 (N_12968,N_6409,N_6258);
and U12969 (N_12969,N_7743,N_5589);
or U12970 (N_12970,N_6942,N_9175);
nor U12971 (N_12971,N_7293,N_7284);
nand U12972 (N_12972,N_9949,N_6655);
nor U12973 (N_12973,N_7559,N_7519);
nand U12974 (N_12974,N_7852,N_7958);
or U12975 (N_12975,N_7366,N_9821);
nor U12976 (N_12976,N_6340,N_8779);
or U12977 (N_12977,N_7681,N_7793);
nand U12978 (N_12978,N_9416,N_7836);
and U12979 (N_12979,N_9729,N_5579);
nand U12980 (N_12980,N_8359,N_6027);
nand U12981 (N_12981,N_9117,N_5664);
or U12982 (N_12982,N_7893,N_6610);
or U12983 (N_12983,N_5278,N_8228);
nand U12984 (N_12984,N_5556,N_5077);
and U12985 (N_12985,N_7477,N_9531);
and U12986 (N_12986,N_6654,N_9666);
or U12987 (N_12987,N_9721,N_7793);
or U12988 (N_12988,N_5172,N_9108);
nand U12989 (N_12989,N_6928,N_9929);
nand U12990 (N_12990,N_5627,N_8572);
and U12991 (N_12991,N_7602,N_8419);
or U12992 (N_12992,N_6986,N_7226);
nand U12993 (N_12993,N_9810,N_6890);
and U12994 (N_12994,N_6431,N_8259);
and U12995 (N_12995,N_7461,N_9531);
and U12996 (N_12996,N_7422,N_7832);
nand U12997 (N_12997,N_8079,N_7054);
nand U12998 (N_12998,N_5288,N_6476);
nor U12999 (N_12999,N_6890,N_7156);
xor U13000 (N_13000,N_9386,N_6303);
or U13001 (N_13001,N_6596,N_7858);
nand U13002 (N_13002,N_7080,N_6380);
nand U13003 (N_13003,N_5959,N_7775);
nor U13004 (N_13004,N_5840,N_7809);
and U13005 (N_13005,N_8927,N_8961);
nor U13006 (N_13006,N_9661,N_9101);
nand U13007 (N_13007,N_6184,N_9430);
nand U13008 (N_13008,N_7223,N_7063);
or U13009 (N_13009,N_7797,N_9471);
nor U13010 (N_13010,N_9408,N_9735);
nand U13011 (N_13011,N_6306,N_8810);
nor U13012 (N_13012,N_6941,N_6456);
and U13013 (N_13013,N_6719,N_9372);
nor U13014 (N_13014,N_7666,N_5245);
or U13015 (N_13015,N_6491,N_7578);
nor U13016 (N_13016,N_5471,N_7043);
nand U13017 (N_13017,N_7254,N_9666);
and U13018 (N_13018,N_7690,N_9770);
and U13019 (N_13019,N_5459,N_8618);
nor U13020 (N_13020,N_8306,N_5492);
nor U13021 (N_13021,N_9882,N_5758);
and U13022 (N_13022,N_7851,N_5330);
and U13023 (N_13023,N_6465,N_6958);
or U13024 (N_13024,N_5331,N_9294);
nand U13025 (N_13025,N_6063,N_5593);
nand U13026 (N_13026,N_7372,N_6663);
and U13027 (N_13027,N_9281,N_5234);
nand U13028 (N_13028,N_9318,N_7341);
nor U13029 (N_13029,N_7125,N_8734);
or U13030 (N_13030,N_9252,N_7680);
nor U13031 (N_13031,N_7098,N_6212);
and U13032 (N_13032,N_8563,N_7486);
or U13033 (N_13033,N_6807,N_6623);
nor U13034 (N_13034,N_5704,N_5881);
nor U13035 (N_13035,N_5381,N_7702);
nor U13036 (N_13036,N_6582,N_8514);
nor U13037 (N_13037,N_7430,N_6546);
or U13038 (N_13038,N_5705,N_8923);
and U13039 (N_13039,N_7013,N_7069);
nor U13040 (N_13040,N_5484,N_5925);
or U13041 (N_13041,N_5156,N_9000);
and U13042 (N_13042,N_6852,N_9833);
nor U13043 (N_13043,N_5746,N_5277);
and U13044 (N_13044,N_8353,N_9006);
nand U13045 (N_13045,N_7828,N_9885);
nor U13046 (N_13046,N_6323,N_8182);
or U13047 (N_13047,N_5545,N_7704);
or U13048 (N_13048,N_9754,N_5751);
or U13049 (N_13049,N_6934,N_8167);
or U13050 (N_13050,N_9452,N_9325);
or U13051 (N_13051,N_5946,N_6997);
or U13052 (N_13052,N_6138,N_8279);
and U13053 (N_13053,N_7930,N_5843);
nor U13054 (N_13054,N_9627,N_9950);
nand U13055 (N_13055,N_7160,N_5333);
nor U13056 (N_13056,N_7441,N_9344);
or U13057 (N_13057,N_6802,N_5678);
nand U13058 (N_13058,N_7672,N_9538);
nor U13059 (N_13059,N_9665,N_8647);
nor U13060 (N_13060,N_9194,N_6347);
nor U13061 (N_13061,N_8456,N_7038);
nand U13062 (N_13062,N_6458,N_6973);
and U13063 (N_13063,N_7866,N_6343);
nor U13064 (N_13064,N_9685,N_6409);
and U13065 (N_13065,N_8005,N_9663);
or U13066 (N_13066,N_7157,N_7261);
or U13067 (N_13067,N_8689,N_7153);
nor U13068 (N_13068,N_9186,N_5945);
nand U13069 (N_13069,N_9760,N_6781);
or U13070 (N_13070,N_6710,N_9781);
or U13071 (N_13071,N_6552,N_5424);
nor U13072 (N_13072,N_6089,N_8676);
or U13073 (N_13073,N_8955,N_8731);
and U13074 (N_13074,N_8264,N_6407);
or U13075 (N_13075,N_5510,N_7968);
nand U13076 (N_13076,N_6722,N_9853);
nor U13077 (N_13077,N_8961,N_7802);
nand U13078 (N_13078,N_8221,N_5144);
and U13079 (N_13079,N_6309,N_7942);
nor U13080 (N_13080,N_6417,N_6042);
nand U13081 (N_13081,N_6960,N_8173);
nor U13082 (N_13082,N_9548,N_7198);
nor U13083 (N_13083,N_5076,N_5764);
nand U13084 (N_13084,N_5569,N_7755);
nor U13085 (N_13085,N_9409,N_9266);
and U13086 (N_13086,N_6924,N_6327);
xor U13087 (N_13087,N_6475,N_7276);
or U13088 (N_13088,N_5055,N_8967);
or U13089 (N_13089,N_6779,N_6813);
or U13090 (N_13090,N_9464,N_6429);
nor U13091 (N_13091,N_5946,N_8595);
nor U13092 (N_13092,N_7752,N_6106);
nor U13093 (N_13093,N_6840,N_5434);
or U13094 (N_13094,N_6229,N_5342);
and U13095 (N_13095,N_8786,N_8183);
nor U13096 (N_13096,N_6707,N_6885);
and U13097 (N_13097,N_8477,N_5789);
nand U13098 (N_13098,N_5736,N_8203);
and U13099 (N_13099,N_7539,N_5351);
nand U13100 (N_13100,N_8044,N_5601);
nand U13101 (N_13101,N_8950,N_5720);
and U13102 (N_13102,N_7163,N_9456);
and U13103 (N_13103,N_8473,N_8375);
and U13104 (N_13104,N_6718,N_8054);
and U13105 (N_13105,N_9172,N_8211);
or U13106 (N_13106,N_8558,N_7728);
or U13107 (N_13107,N_5461,N_9189);
and U13108 (N_13108,N_8346,N_6652);
or U13109 (N_13109,N_5394,N_9582);
xor U13110 (N_13110,N_5315,N_8397);
or U13111 (N_13111,N_8732,N_5743);
or U13112 (N_13112,N_6537,N_8771);
and U13113 (N_13113,N_8225,N_7980);
nor U13114 (N_13114,N_8829,N_5287);
xnor U13115 (N_13115,N_8839,N_6761);
or U13116 (N_13116,N_8504,N_5824);
or U13117 (N_13117,N_8249,N_5308);
nand U13118 (N_13118,N_9297,N_8283);
nor U13119 (N_13119,N_8324,N_8255);
nand U13120 (N_13120,N_5817,N_6650);
nor U13121 (N_13121,N_5926,N_6903);
and U13122 (N_13122,N_6740,N_5452);
or U13123 (N_13123,N_6861,N_6357);
nand U13124 (N_13124,N_6128,N_8544);
nand U13125 (N_13125,N_5258,N_9333);
nor U13126 (N_13126,N_5392,N_5985);
or U13127 (N_13127,N_9264,N_5856);
and U13128 (N_13128,N_8850,N_8725);
nor U13129 (N_13129,N_5266,N_6164);
or U13130 (N_13130,N_6981,N_7893);
nor U13131 (N_13131,N_8860,N_7884);
nor U13132 (N_13132,N_7364,N_6021);
nor U13133 (N_13133,N_9511,N_5566);
or U13134 (N_13134,N_6532,N_7869);
nor U13135 (N_13135,N_7031,N_5793);
and U13136 (N_13136,N_5082,N_9889);
or U13137 (N_13137,N_6923,N_7456);
nor U13138 (N_13138,N_6411,N_8293);
nor U13139 (N_13139,N_8294,N_6313);
nor U13140 (N_13140,N_9428,N_9449);
nor U13141 (N_13141,N_9621,N_8109);
nor U13142 (N_13142,N_9993,N_5355);
or U13143 (N_13143,N_9869,N_9619);
nor U13144 (N_13144,N_8183,N_6015);
nor U13145 (N_13145,N_8587,N_7184);
and U13146 (N_13146,N_8431,N_9114);
or U13147 (N_13147,N_5612,N_9074);
nand U13148 (N_13148,N_8644,N_5160);
nand U13149 (N_13149,N_5512,N_9647);
and U13150 (N_13150,N_5271,N_5210);
and U13151 (N_13151,N_7142,N_8668);
and U13152 (N_13152,N_7983,N_6372);
and U13153 (N_13153,N_8461,N_6059);
nand U13154 (N_13154,N_7291,N_9586);
or U13155 (N_13155,N_7197,N_7920);
nor U13156 (N_13156,N_9967,N_5844);
or U13157 (N_13157,N_6181,N_9326);
or U13158 (N_13158,N_7139,N_9641);
or U13159 (N_13159,N_8313,N_8361);
nand U13160 (N_13160,N_9844,N_5690);
nand U13161 (N_13161,N_5162,N_7767);
nand U13162 (N_13162,N_6552,N_7969);
or U13163 (N_13163,N_6071,N_6338);
and U13164 (N_13164,N_7774,N_7721);
and U13165 (N_13165,N_8381,N_8538);
nor U13166 (N_13166,N_5180,N_8801);
and U13167 (N_13167,N_8977,N_6790);
nor U13168 (N_13168,N_8096,N_5562);
nor U13169 (N_13169,N_9520,N_9790);
and U13170 (N_13170,N_5740,N_5232);
xor U13171 (N_13171,N_8725,N_8874);
nand U13172 (N_13172,N_7197,N_8183);
nor U13173 (N_13173,N_9644,N_9501);
and U13174 (N_13174,N_6539,N_5327);
nor U13175 (N_13175,N_6255,N_7909);
xnor U13176 (N_13176,N_6321,N_7599);
nand U13177 (N_13177,N_7255,N_6341);
nand U13178 (N_13178,N_7493,N_7499);
nand U13179 (N_13179,N_6496,N_8926);
nand U13180 (N_13180,N_6158,N_8832);
nand U13181 (N_13181,N_6460,N_5719);
nor U13182 (N_13182,N_8946,N_9959);
or U13183 (N_13183,N_9705,N_8357);
nor U13184 (N_13184,N_7562,N_8659);
nor U13185 (N_13185,N_5223,N_6543);
or U13186 (N_13186,N_8025,N_9870);
nor U13187 (N_13187,N_5935,N_6676);
or U13188 (N_13188,N_8864,N_5253);
nor U13189 (N_13189,N_8353,N_5412);
nand U13190 (N_13190,N_9019,N_6622);
nor U13191 (N_13191,N_7820,N_6615);
nor U13192 (N_13192,N_8330,N_7758);
nand U13193 (N_13193,N_9141,N_5096);
nor U13194 (N_13194,N_5761,N_5955);
nor U13195 (N_13195,N_6855,N_9523);
nor U13196 (N_13196,N_7933,N_5689);
nor U13197 (N_13197,N_6174,N_9561);
and U13198 (N_13198,N_8607,N_9319);
or U13199 (N_13199,N_5757,N_5970);
and U13200 (N_13200,N_8871,N_7612);
nor U13201 (N_13201,N_5635,N_5785);
and U13202 (N_13202,N_8854,N_7931);
xnor U13203 (N_13203,N_9853,N_9700);
nor U13204 (N_13204,N_8320,N_6609);
nor U13205 (N_13205,N_7174,N_8468);
and U13206 (N_13206,N_5643,N_7268);
nand U13207 (N_13207,N_9262,N_8638);
nor U13208 (N_13208,N_8885,N_5247);
nand U13209 (N_13209,N_6456,N_9332);
nand U13210 (N_13210,N_9922,N_6047);
and U13211 (N_13211,N_6319,N_7985);
nor U13212 (N_13212,N_8415,N_5739);
nor U13213 (N_13213,N_8942,N_5943);
and U13214 (N_13214,N_8550,N_8345);
xnor U13215 (N_13215,N_9436,N_9996);
and U13216 (N_13216,N_5593,N_7702);
or U13217 (N_13217,N_5740,N_9366);
or U13218 (N_13218,N_5937,N_6842);
nand U13219 (N_13219,N_8737,N_7576);
nor U13220 (N_13220,N_9928,N_7628);
and U13221 (N_13221,N_8396,N_9333);
or U13222 (N_13222,N_8929,N_7662);
nand U13223 (N_13223,N_6575,N_8236);
nor U13224 (N_13224,N_7777,N_5226);
or U13225 (N_13225,N_7760,N_7837);
and U13226 (N_13226,N_5173,N_5032);
and U13227 (N_13227,N_8575,N_8652);
nor U13228 (N_13228,N_8021,N_9455);
xnor U13229 (N_13229,N_8485,N_6938);
and U13230 (N_13230,N_5320,N_9240);
or U13231 (N_13231,N_7382,N_7150);
and U13232 (N_13232,N_5000,N_6181);
nor U13233 (N_13233,N_9671,N_9972);
or U13234 (N_13234,N_8049,N_9120);
and U13235 (N_13235,N_6234,N_9688);
nor U13236 (N_13236,N_7229,N_7644);
or U13237 (N_13237,N_8080,N_8669);
nand U13238 (N_13238,N_6130,N_5626);
or U13239 (N_13239,N_8719,N_5263);
or U13240 (N_13240,N_9882,N_8322);
and U13241 (N_13241,N_5685,N_6033);
and U13242 (N_13242,N_5148,N_8816);
nand U13243 (N_13243,N_7228,N_6692);
and U13244 (N_13244,N_5690,N_9934);
nor U13245 (N_13245,N_8661,N_7163);
nand U13246 (N_13246,N_5532,N_9955);
nor U13247 (N_13247,N_5837,N_7336);
nor U13248 (N_13248,N_9114,N_9087);
nand U13249 (N_13249,N_6056,N_6777);
nand U13250 (N_13250,N_6791,N_5743);
nor U13251 (N_13251,N_9238,N_8836);
xor U13252 (N_13252,N_7833,N_9778);
nor U13253 (N_13253,N_8782,N_5163);
nand U13254 (N_13254,N_7761,N_9603);
nand U13255 (N_13255,N_6161,N_5889);
and U13256 (N_13256,N_5821,N_8215);
or U13257 (N_13257,N_8147,N_5626);
and U13258 (N_13258,N_8574,N_7080);
or U13259 (N_13259,N_7846,N_6777);
nor U13260 (N_13260,N_6477,N_6772);
nand U13261 (N_13261,N_8499,N_8069);
nor U13262 (N_13262,N_8695,N_9028);
and U13263 (N_13263,N_6405,N_6471);
nand U13264 (N_13264,N_7240,N_6004);
nand U13265 (N_13265,N_5345,N_9923);
and U13266 (N_13266,N_7901,N_7906);
nand U13267 (N_13267,N_9706,N_6236);
and U13268 (N_13268,N_8426,N_8709);
nor U13269 (N_13269,N_5496,N_6441);
and U13270 (N_13270,N_7465,N_7919);
nand U13271 (N_13271,N_8565,N_9628);
or U13272 (N_13272,N_8814,N_9785);
nand U13273 (N_13273,N_9897,N_5907);
or U13274 (N_13274,N_8964,N_8017);
nand U13275 (N_13275,N_8863,N_8707);
nand U13276 (N_13276,N_5138,N_5544);
nand U13277 (N_13277,N_5591,N_8044);
and U13278 (N_13278,N_7209,N_9935);
nor U13279 (N_13279,N_7820,N_8127);
nand U13280 (N_13280,N_7961,N_5125);
nand U13281 (N_13281,N_6157,N_9874);
and U13282 (N_13282,N_7636,N_6470);
nand U13283 (N_13283,N_6298,N_7281);
nand U13284 (N_13284,N_7486,N_9599);
and U13285 (N_13285,N_8630,N_6280);
or U13286 (N_13286,N_9215,N_8853);
or U13287 (N_13287,N_7833,N_5303);
or U13288 (N_13288,N_8763,N_9302);
or U13289 (N_13289,N_6586,N_6984);
or U13290 (N_13290,N_5209,N_7072);
or U13291 (N_13291,N_6929,N_6103);
or U13292 (N_13292,N_9031,N_6694);
nor U13293 (N_13293,N_5104,N_8650);
nand U13294 (N_13294,N_5064,N_7376);
and U13295 (N_13295,N_5618,N_7646);
and U13296 (N_13296,N_7121,N_7625);
nand U13297 (N_13297,N_5575,N_8362);
nand U13298 (N_13298,N_8789,N_8338);
nand U13299 (N_13299,N_5222,N_6680);
or U13300 (N_13300,N_6219,N_9593);
nor U13301 (N_13301,N_5357,N_9447);
and U13302 (N_13302,N_5356,N_5431);
and U13303 (N_13303,N_7401,N_6216);
and U13304 (N_13304,N_5557,N_9898);
nor U13305 (N_13305,N_5541,N_9040);
nor U13306 (N_13306,N_9484,N_7128);
and U13307 (N_13307,N_8590,N_7340);
and U13308 (N_13308,N_8542,N_8708);
or U13309 (N_13309,N_7996,N_8193);
nor U13310 (N_13310,N_5785,N_5538);
nand U13311 (N_13311,N_9699,N_6212);
nor U13312 (N_13312,N_6298,N_9775);
or U13313 (N_13313,N_6458,N_9783);
nand U13314 (N_13314,N_7886,N_7191);
and U13315 (N_13315,N_9975,N_9580);
and U13316 (N_13316,N_6329,N_5646);
nor U13317 (N_13317,N_7719,N_6609);
or U13318 (N_13318,N_9343,N_8713);
xnor U13319 (N_13319,N_8912,N_6996);
or U13320 (N_13320,N_7083,N_6865);
or U13321 (N_13321,N_7024,N_9799);
nand U13322 (N_13322,N_7786,N_5208);
nor U13323 (N_13323,N_8253,N_9267);
or U13324 (N_13324,N_9538,N_7990);
nor U13325 (N_13325,N_5653,N_7187);
and U13326 (N_13326,N_7228,N_7981);
and U13327 (N_13327,N_5942,N_6366);
nor U13328 (N_13328,N_9392,N_8494);
nand U13329 (N_13329,N_7948,N_5375);
and U13330 (N_13330,N_9820,N_9260);
xor U13331 (N_13331,N_9096,N_8896);
nor U13332 (N_13332,N_8883,N_5107);
nor U13333 (N_13333,N_6134,N_9177);
nor U13334 (N_13334,N_5168,N_9120);
nor U13335 (N_13335,N_6530,N_7076);
or U13336 (N_13336,N_8192,N_9135);
nor U13337 (N_13337,N_7446,N_6048);
nand U13338 (N_13338,N_6690,N_5713);
or U13339 (N_13339,N_9803,N_8978);
or U13340 (N_13340,N_9466,N_7001);
nand U13341 (N_13341,N_8358,N_9846);
nor U13342 (N_13342,N_7003,N_5602);
and U13343 (N_13343,N_9422,N_6372);
and U13344 (N_13344,N_5674,N_9813);
nand U13345 (N_13345,N_6259,N_8434);
or U13346 (N_13346,N_5601,N_5518);
nand U13347 (N_13347,N_8377,N_7092);
and U13348 (N_13348,N_5050,N_7822);
nor U13349 (N_13349,N_6182,N_7547);
and U13350 (N_13350,N_9659,N_5323);
and U13351 (N_13351,N_5236,N_5663);
nor U13352 (N_13352,N_9084,N_6866);
nor U13353 (N_13353,N_6762,N_8798);
nor U13354 (N_13354,N_7329,N_5718);
xor U13355 (N_13355,N_8097,N_5232);
nor U13356 (N_13356,N_7890,N_7018);
and U13357 (N_13357,N_9924,N_9883);
and U13358 (N_13358,N_9627,N_6909);
nor U13359 (N_13359,N_8150,N_7736);
or U13360 (N_13360,N_8221,N_8409);
or U13361 (N_13361,N_9053,N_6206);
and U13362 (N_13362,N_5244,N_7881);
nand U13363 (N_13363,N_5362,N_8758);
or U13364 (N_13364,N_6858,N_5652);
nand U13365 (N_13365,N_6152,N_6307);
or U13366 (N_13366,N_8509,N_8073);
nand U13367 (N_13367,N_7412,N_8261);
and U13368 (N_13368,N_8844,N_9700);
and U13369 (N_13369,N_7475,N_7436);
xor U13370 (N_13370,N_8041,N_7597);
or U13371 (N_13371,N_6772,N_8751);
nand U13372 (N_13372,N_6604,N_7387);
and U13373 (N_13373,N_7496,N_9260);
xnor U13374 (N_13374,N_6840,N_9991);
or U13375 (N_13375,N_6478,N_5196);
or U13376 (N_13376,N_9790,N_7590);
or U13377 (N_13377,N_9471,N_6507);
or U13378 (N_13378,N_5752,N_7660);
nor U13379 (N_13379,N_7093,N_8558);
nor U13380 (N_13380,N_8004,N_5265);
or U13381 (N_13381,N_8249,N_8082);
or U13382 (N_13382,N_5553,N_9737);
nor U13383 (N_13383,N_5807,N_6512);
nand U13384 (N_13384,N_8634,N_6241);
nor U13385 (N_13385,N_5969,N_9122);
and U13386 (N_13386,N_5139,N_8847);
or U13387 (N_13387,N_5817,N_9482);
or U13388 (N_13388,N_5436,N_8021);
xor U13389 (N_13389,N_9819,N_6951);
nor U13390 (N_13390,N_5068,N_8901);
nand U13391 (N_13391,N_8003,N_7105);
nor U13392 (N_13392,N_7378,N_8347);
nand U13393 (N_13393,N_6944,N_7925);
and U13394 (N_13394,N_6981,N_5242);
nand U13395 (N_13395,N_7461,N_6215);
nor U13396 (N_13396,N_9518,N_5873);
and U13397 (N_13397,N_6250,N_9223);
nor U13398 (N_13398,N_8848,N_8348);
or U13399 (N_13399,N_5106,N_7281);
or U13400 (N_13400,N_5917,N_7815);
nand U13401 (N_13401,N_6448,N_8567);
nor U13402 (N_13402,N_5190,N_7421);
nand U13403 (N_13403,N_7272,N_9180);
nor U13404 (N_13404,N_5038,N_9438);
and U13405 (N_13405,N_8785,N_5330);
and U13406 (N_13406,N_8641,N_8512);
or U13407 (N_13407,N_5832,N_5256);
nor U13408 (N_13408,N_9517,N_8278);
nor U13409 (N_13409,N_5016,N_9192);
or U13410 (N_13410,N_9764,N_6362);
nor U13411 (N_13411,N_7998,N_5420);
and U13412 (N_13412,N_7383,N_7240);
and U13413 (N_13413,N_6290,N_9167);
nand U13414 (N_13414,N_6976,N_6230);
nand U13415 (N_13415,N_5895,N_9253);
nor U13416 (N_13416,N_6416,N_5521);
nor U13417 (N_13417,N_8836,N_5393);
or U13418 (N_13418,N_5927,N_6774);
nor U13419 (N_13419,N_6537,N_6668);
and U13420 (N_13420,N_9298,N_9198);
nor U13421 (N_13421,N_8792,N_9995);
and U13422 (N_13422,N_6469,N_8523);
and U13423 (N_13423,N_5690,N_8204);
nor U13424 (N_13424,N_5270,N_6456);
nor U13425 (N_13425,N_5189,N_9895);
nand U13426 (N_13426,N_9381,N_7955);
and U13427 (N_13427,N_9455,N_8146);
and U13428 (N_13428,N_8154,N_5813);
and U13429 (N_13429,N_9602,N_7034);
nand U13430 (N_13430,N_6851,N_9452);
nand U13431 (N_13431,N_8852,N_5720);
nor U13432 (N_13432,N_8704,N_9929);
nor U13433 (N_13433,N_5731,N_7882);
and U13434 (N_13434,N_6846,N_9764);
and U13435 (N_13435,N_9907,N_8811);
nand U13436 (N_13436,N_6416,N_9069);
nor U13437 (N_13437,N_6418,N_5299);
nand U13438 (N_13438,N_7446,N_6724);
nor U13439 (N_13439,N_6419,N_9905);
xor U13440 (N_13440,N_6377,N_8344);
or U13441 (N_13441,N_5322,N_5791);
or U13442 (N_13442,N_6672,N_6918);
nor U13443 (N_13443,N_6797,N_5443);
and U13444 (N_13444,N_8298,N_8610);
nand U13445 (N_13445,N_5474,N_8248);
nor U13446 (N_13446,N_8840,N_8980);
or U13447 (N_13447,N_6645,N_6377);
nor U13448 (N_13448,N_8765,N_9304);
or U13449 (N_13449,N_6932,N_6007);
and U13450 (N_13450,N_6959,N_6057);
nor U13451 (N_13451,N_7043,N_6303);
or U13452 (N_13452,N_6302,N_5861);
nand U13453 (N_13453,N_5981,N_7821);
and U13454 (N_13454,N_5643,N_5234);
or U13455 (N_13455,N_6297,N_6565);
nor U13456 (N_13456,N_5857,N_7900);
or U13457 (N_13457,N_9305,N_5685);
or U13458 (N_13458,N_5008,N_7038);
and U13459 (N_13459,N_7372,N_5981);
or U13460 (N_13460,N_9846,N_5721);
nor U13461 (N_13461,N_5732,N_9489);
or U13462 (N_13462,N_7834,N_9965);
xor U13463 (N_13463,N_7347,N_5682);
nor U13464 (N_13464,N_8838,N_9939);
nand U13465 (N_13465,N_9010,N_9649);
or U13466 (N_13466,N_9216,N_9490);
nand U13467 (N_13467,N_8524,N_5810);
nand U13468 (N_13468,N_6598,N_9276);
nor U13469 (N_13469,N_6838,N_7576);
and U13470 (N_13470,N_8837,N_6248);
nor U13471 (N_13471,N_7491,N_6100);
nor U13472 (N_13472,N_7100,N_5494);
nand U13473 (N_13473,N_7704,N_9600);
or U13474 (N_13474,N_5122,N_7266);
and U13475 (N_13475,N_5554,N_9449);
or U13476 (N_13476,N_7450,N_6731);
nor U13477 (N_13477,N_8702,N_8435);
and U13478 (N_13478,N_6075,N_8084);
or U13479 (N_13479,N_6017,N_5723);
and U13480 (N_13480,N_9040,N_5649);
nor U13481 (N_13481,N_8041,N_7563);
nor U13482 (N_13482,N_5996,N_5419);
nand U13483 (N_13483,N_8021,N_6586);
and U13484 (N_13484,N_9154,N_7505);
nand U13485 (N_13485,N_7484,N_5236);
nor U13486 (N_13486,N_5746,N_7684);
and U13487 (N_13487,N_6661,N_9619);
xnor U13488 (N_13488,N_9089,N_9205);
nand U13489 (N_13489,N_6798,N_7693);
or U13490 (N_13490,N_7577,N_6140);
and U13491 (N_13491,N_6350,N_6688);
nor U13492 (N_13492,N_8392,N_6829);
nor U13493 (N_13493,N_7314,N_9072);
xnor U13494 (N_13494,N_7553,N_7355);
or U13495 (N_13495,N_7012,N_7603);
and U13496 (N_13496,N_6594,N_7733);
nor U13497 (N_13497,N_8075,N_7054);
nand U13498 (N_13498,N_6476,N_7906);
and U13499 (N_13499,N_9614,N_6372);
xnor U13500 (N_13500,N_7335,N_5384);
or U13501 (N_13501,N_8460,N_9927);
or U13502 (N_13502,N_7806,N_8198);
nand U13503 (N_13503,N_7480,N_9711);
or U13504 (N_13504,N_6301,N_5522);
nand U13505 (N_13505,N_5569,N_8971);
or U13506 (N_13506,N_8302,N_7183);
nand U13507 (N_13507,N_6163,N_5305);
and U13508 (N_13508,N_8232,N_7794);
or U13509 (N_13509,N_6434,N_5986);
and U13510 (N_13510,N_9564,N_5793);
nor U13511 (N_13511,N_5493,N_5982);
nand U13512 (N_13512,N_9555,N_7530);
and U13513 (N_13513,N_7927,N_8412);
nor U13514 (N_13514,N_5921,N_8149);
or U13515 (N_13515,N_9738,N_8102);
and U13516 (N_13516,N_5401,N_9811);
and U13517 (N_13517,N_5189,N_8337);
nand U13518 (N_13518,N_5515,N_8824);
or U13519 (N_13519,N_5175,N_7830);
or U13520 (N_13520,N_7688,N_5917);
nor U13521 (N_13521,N_9631,N_9637);
or U13522 (N_13522,N_6327,N_8532);
or U13523 (N_13523,N_8363,N_8312);
and U13524 (N_13524,N_7297,N_6285);
nand U13525 (N_13525,N_5313,N_7027);
nand U13526 (N_13526,N_7659,N_6623);
and U13527 (N_13527,N_8672,N_5114);
nor U13528 (N_13528,N_5742,N_8206);
nand U13529 (N_13529,N_9310,N_6719);
nor U13530 (N_13530,N_9194,N_8726);
nor U13531 (N_13531,N_7988,N_7286);
and U13532 (N_13532,N_7155,N_8329);
and U13533 (N_13533,N_5750,N_5080);
or U13534 (N_13534,N_7607,N_5472);
nand U13535 (N_13535,N_7622,N_7257);
nand U13536 (N_13536,N_5679,N_9975);
nand U13537 (N_13537,N_9247,N_9353);
and U13538 (N_13538,N_6031,N_6967);
nor U13539 (N_13539,N_6217,N_8249);
nand U13540 (N_13540,N_5922,N_6407);
or U13541 (N_13541,N_8468,N_8671);
nor U13542 (N_13542,N_8510,N_8741);
or U13543 (N_13543,N_6958,N_8260);
and U13544 (N_13544,N_9757,N_7828);
and U13545 (N_13545,N_7550,N_7655);
and U13546 (N_13546,N_7877,N_9194);
nor U13547 (N_13547,N_6493,N_8441);
nor U13548 (N_13548,N_6945,N_5764);
nand U13549 (N_13549,N_7049,N_8663);
or U13550 (N_13550,N_5094,N_7854);
nand U13551 (N_13551,N_9295,N_5113);
nand U13552 (N_13552,N_9286,N_7334);
or U13553 (N_13553,N_9517,N_7051);
and U13554 (N_13554,N_8424,N_5904);
or U13555 (N_13555,N_5770,N_9507);
or U13556 (N_13556,N_5233,N_7470);
nand U13557 (N_13557,N_7833,N_5233);
nor U13558 (N_13558,N_9207,N_6750);
and U13559 (N_13559,N_5479,N_5647);
or U13560 (N_13560,N_6570,N_5708);
and U13561 (N_13561,N_5610,N_8288);
nand U13562 (N_13562,N_9291,N_9615);
and U13563 (N_13563,N_7979,N_5167);
nand U13564 (N_13564,N_8522,N_7238);
nor U13565 (N_13565,N_6622,N_9565);
and U13566 (N_13566,N_5210,N_7229);
nand U13567 (N_13567,N_6469,N_5122);
nand U13568 (N_13568,N_7141,N_8239);
and U13569 (N_13569,N_9782,N_9122);
nand U13570 (N_13570,N_8330,N_5438);
nor U13571 (N_13571,N_8869,N_7209);
nand U13572 (N_13572,N_5582,N_5020);
nand U13573 (N_13573,N_7653,N_7911);
and U13574 (N_13574,N_8278,N_6222);
nand U13575 (N_13575,N_6704,N_5646);
or U13576 (N_13576,N_7269,N_9063);
or U13577 (N_13577,N_7795,N_7668);
nand U13578 (N_13578,N_8096,N_7107);
nor U13579 (N_13579,N_5741,N_9377);
nand U13580 (N_13580,N_8955,N_5003);
nand U13581 (N_13581,N_7705,N_9029);
nand U13582 (N_13582,N_8110,N_9739);
nor U13583 (N_13583,N_6858,N_7481);
nand U13584 (N_13584,N_7676,N_5010);
and U13585 (N_13585,N_9671,N_8666);
nand U13586 (N_13586,N_7428,N_5969);
nor U13587 (N_13587,N_7002,N_7786);
and U13588 (N_13588,N_7778,N_8714);
nand U13589 (N_13589,N_5627,N_5148);
nor U13590 (N_13590,N_7660,N_8610);
or U13591 (N_13591,N_8759,N_9097);
or U13592 (N_13592,N_6054,N_7371);
nand U13593 (N_13593,N_5970,N_7664);
nand U13594 (N_13594,N_5360,N_7720);
nand U13595 (N_13595,N_7753,N_5114);
nand U13596 (N_13596,N_8082,N_6894);
nand U13597 (N_13597,N_5771,N_8395);
or U13598 (N_13598,N_9707,N_8305);
and U13599 (N_13599,N_5888,N_5089);
nor U13600 (N_13600,N_5541,N_9645);
and U13601 (N_13601,N_5753,N_5860);
nor U13602 (N_13602,N_5962,N_5970);
nor U13603 (N_13603,N_9942,N_9390);
or U13604 (N_13604,N_5959,N_7627);
or U13605 (N_13605,N_7259,N_7820);
nand U13606 (N_13606,N_9165,N_5999);
xor U13607 (N_13607,N_8018,N_7731);
nor U13608 (N_13608,N_9410,N_5398);
nor U13609 (N_13609,N_6224,N_5628);
xnor U13610 (N_13610,N_6624,N_5550);
and U13611 (N_13611,N_5225,N_7493);
or U13612 (N_13612,N_9762,N_5584);
or U13613 (N_13613,N_8359,N_6632);
and U13614 (N_13614,N_7649,N_8749);
or U13615 (N_13615,N_9486,N_8257);
nand U13616 (N_13616,N_6807,N_6904);
or U13617 (N_13617,N_8833,N_9645);
nand U13618 (N_13618,N_8664,N_9394);
and U13619 (N_13619,N_7337,N_8630);
and U13620 (N_13620,N_5953,N_9238);
and U13621 (N_13621,N_9245,N_5836);
nand U13622 (N_13622,N_6661,N_6404);
and U13623 (N_13623,N_6730,N_6266);
nor U13624 (N_13624,N_7626,N_5697);
or U13625 (N_13625,N_5643,N_9216);
or U13626 (N_13626,N_6114,N_6367);
or U13627 (N_13627,N_9682,N_7117);
and U13628 (N_13628,N_9538,N_9158);
nand U13629 (N_13629,N_9394,N_7607);
nor U13630 (N_13630,N_7189,N_7386);
nand U13631 (N_13631,N_7275,N_9207);
nand U13632 (N_13632,N_5936,N_8974);
and U13633 (N_13633,N_6427,N_9081);
nor U13634 (N_13634,N_8606,N_6175);
and U13635 (N_13635,N_7077,N_8936);
and U13636 (N_13636,N_6701,N_6672);
nor U13637 (N_13637,N_5431,N_7264);
or U13638 (N_13638,N_6391,N_8991);
and U13639 (N_13639,N_7768,N_8332);
nand U13640 (N_13640,N_6070,N_7619);
or U13641 (N_13641,N_8192,N_7846);
and U13642 (N_13642,N_6291,N_6633);
nor U13643 (N_13643,N_8924,N_8693);
nor U13644 (N_13644,N_5567,N_9237);
or U13645 (N_13645,N_8738,N_5027);
nor U13646 (N_13646,N_5094,N_7962);
or U13647 (N_13647,N_9400,N_6319);
nand U13648 (N_13648,N_8197,N_6147);
nor U13649 (N_13649,N_6720,N_8060);
or U13650 (N_13650,N_9409,N_9105);
or U13651 (N_13651,N_8799,N_9078);
nor U13652 (N_13652,N_5924,N_9624);
and U13653 (N_13653,N_9004,N_6836);
or U13654 (N_13654,N_7755,N_5502);
or U13655 (N_13655,N_6138,N_7310);
nor U13656 (N_13656,N_5367,N_7600);
or U13657 (N_13657,N_8041,N_6141);
or U13658 (N_13658,N_6813,N_9895);
or U13659 (N_13659,N_6288,N_9236);
nor U13660 (N_13660,N_7515,N_6259);
or U13661 (N_13661,N_6424,N_8449);
and U13662 (N_13662,N_7703,N_7976);
nor U13663 (N_13663,N_7913,N_7058);
or U13664 (N_13664,N_6311,N_5648);
and U13665 (N_13665,N_8636,N_7254);
nor U13666 (N_13666,N_5235,N_8564);
and U13667 (N_13667,N_6632,N_5816);
and U13668 (N_13668,N_8786,N_5641);
nand U13669 (N_13669,N_5324,N_7216);
nand U13670 (N_13670,N_5139,N_7826);
and U13671 (N_13671,N_7551,N_9259);
and U13672 (N_13672,N_7236,N_8012);
or U13673 (N_13673,N_9189,N_7549);
nor U13674 (N_13674,N_7188,N_5964);
or U13675 (N_13675,N_5282,N_8864);
nor U13676 (N_13676,N_9232,N_5859);
nor U13677 (N_13677,N_5575,N_9785);
nand U13678 (N_13678,N_6702,N_7031);
and U13679 (N_13679,N_5492,N_5034);
or U13680 (N_13680,N_5488,N_9839);
and U13681 (N_13681,N_8943,N_7296);
nor U13682 (N_13682,N_5328,N_7436);
nand U13683 (N_13683,N_9829,N_7094);
nor U13684 (N_13684,N_9304,N_8335);
nor U13685 (N_13685,N_5614,N_9599);
and U13686 (N_13686,N_7166,N_5790);
nand U13687 (N_13687,N_9298,N_5246);
nor U13688 (N_13688,N_9576,N_9751);
and U13689 (N_13689,N_6384,N_9516);
or U13690 (N_13690,N_8653,N_6495);
nor U13691 (N_13691,N_6569,N_7372);
and U13692 (N_13692,N_8344,N_6696);
or U13693 (N_13693,N_8024,N_8147);
and U13694 (N_13694,N_9458,N_9533);
nor U13695 (N_13695,N_5472,N_6183);
or U13696 (N_13696,N_5359,N_7013);
nor U13697 (N_13697,N_8616,N_6562);
or U13698 (N_13698,N_9283,N_7486);
nand U13699 (N_13699,N_5222,N_7703);
or U13700 (N_13700,N_6817,N_6854);
or U13701 (N_13701,N_8813,N_5777);
nand U13702 (N_13702,N_9933,N_7134);
or U13703 (N_13703,N_6442,N_6405);
and U13704 (N_13704,N_7992,N_7101);
nor U13705 (N_13705,N_5902,N_5074);
and U13706 (N_13706,N_8266,N_5515);
or U13707 (N_13707,N_5732,N_7148);
nand U13708 (N_13708,N_8035,N_8730);
or U13709 (N_13709,N_7847,N_6526);
nor U13710 (N_13710,N_6528,N_8458);
nand U13711 (N_13711,N_7462,N_6602);
nand U13712 (N_13712,N_7852,N_7084);
nand U13713 (N_13713,N_9692,N_7030);
nand U13714 (N_13714,N_9549,N_7415);
nor U13715 (N_13715,N_7282,N_7453);
and U13716 (N_13716,N_8662,N_6110);
nand U13717 (N_13717,N_8427,N_8337);
nand U13718 (N_13718,N_7957,N_5894);
and U13719 (N_13719,N_6686,N_8437);
or U13720 (N_13720,N_5218,N_5894);
nor U13721 (N_13721,N_5732,N_5232);
nor U13722 (N_13722,N_5987,N_5907);
or U13723 (N_13723,N_8433,N_5583);
nor U13724 (N_13724,N_8081,N_6174);
nand U13725 (N_13725,N_9429,N_6634);
and U13726 (N_13726,N_7619,N_6160);
and U13727 (N_13727,N_6928,N_7224);
nand U13728 (N_13728,N_9109,N_5699);
or U13729 (N_13729,N_9148,N_6341);
nand U13730 (N_13730,N_5976,N_5561);
nor U13731 (N_13731,N_7918,N_6996);
and U13732 (N_13732,N_6712,N_7353);
or U13733 (N_13733,N_6970,N_5663);
nand U13734 (N_13734,N_6390,N_5979);
nand U13735 (N_13735,N_8111,N_7338);
or U13736 (N_13736,N_7798,N_7568);
xor U13737 (N_13737,N_8898,N_7467);
and U13738 (N_13738,N_8015,N_5334);
nor U13739 (N_13739,N_8176,N_5063);
and U13740 (N_13740,N_6523,N_8776);
nand U13741 (N_13741,N_6799,N_9682);
nand U13742 (N_13742,N_8890,N_5954);
nor U13743 (N_13743,N_5322,N_9249);
or U13744 (N_13744,N_8841,N_8189);
or U13745 (N_13745,N_5692,N_5686);
and U13746 (N_13746,N_5055,N_8075);
or U13747 (N_13747,N_7267,N_5593);
nor U13748 (N_13748,N_8230,N_5676);
nand U13749 (N_13749,N_5610,N_9123);
and U13750 (N_13750,N_6605,N_5700);
or U13751 (N_13751,N_5591,N_6108);
nand U13752 (N_13752,N_6606,N_9348);
or U13753 (N_13753,N_7345,N_6093);
and U13754 (N_13754,N_8821,N_6506);
and U13755 (N_13755,N_9749,N_8646);
nand U13756 (N_13756,N_8197,N_8876);
or U13757 (N_13757,N_5735,N_7053);
nor U13758 (N_13758,N_9422,N_7485);
and U13759 (N_13759,N_7379,N_5588);
nand U13760 (N_13760,N_7653,N_7309);
nor U13761 (N_13761,N_9705,N_9161);
nor U13762 (N_13762,N_9659,N_8659);
and U13763 (N_13763,N_9175,N_8577);
nand U13764 (N_13764,N_8642,N_6641);
nor U13765 (N_13765,N_6101,N_9901);
nor U13766 (N_13766,N_8270,N_5694);
nor U13767 (N_13767,N_7124,N_7187);
nand U13768 (N_13768,N_5452,N_8575);
or U13769 (N_13769,N_6063,N_5022);
nand U13770 (N_13770,N_5414,N_8325);
and U13771 (N_13771,N_8691,N_5275);
nand U13772 (N_13772,N_7709,N_8318);
or U13773 (N_13773,N_6961,N_9345);
nand U13774 (N_13774,N_5735,N_6093);
nand U13775 (N_13775,N_5212,N_5412);
or U13776 (N_13776,N_5979,N_6313);
nand U13777 (N_13777,N_7947,N_7681);
nand U13778 (N_13778,N_7988,N_7803);
nor U13779 (N_13779,N_5015,N_6653);
or U13780 (N_13780,N_8545,N_6874);
and U13781 (N_13781,N_6814,N_7626);
or U13782 (N_13782,N_6488,N_5005);
and U13783 (N_13783,N_9626,N_6237);
and U13784 (N_13784,N_8116,N_9491);
and U13785 (N_13785,N_8795,N_7196);
nor U13786 (N_13786,N_8279,N_7988);
and U13787 (N_13787,N_7756,N_5140);
nand U13788 (N_13788,N_6140,N_6739);
nand U13789 (N_13789,N_8389,N_7999);
or U13790 (N_13790,N_6056,N_7520);
or U13791 (N_13791,N_7429,N_7212);
nand U13792 (N_13792,N_6551,N_5081);
nor U13793 (N_13793,N_5725,N_7909);
or U13794 (N_13794,N_8518,N_6085);
nor U13795 (N_13795,N_6928,N_7557);
or U13796 (N_13796,N_6457,N_5808);
and U13797 (N_13797,N_8503,N_6123);
or U13798 (N_13798,N_9262,N_6299);
nor U13799 (N_13799,N_5325,N_6944);
nor U13800 (N_13800,N_5464,N_6115);
and U13801 (N_13801,N_9413,N_6572);
and U13802 (N_13802,N_6511,N_6327);
nand U13803 (N_13803,N_8165,N_6181);
nand U13804 (N_13804,N_8766,N_7783);
nor U13805 (N_13805,N_6199,N_8877);
or U13806 (N_13806,N_5734,N_5228);
nor U13807 (N_13807,N_5446,N_6890);
nor U13808 (N_13808,N_8997,N_5319);
and U13809 (N_13809,N_6832,N_7798);
or U13810 (N_13810,N_8217,N_7620);
nor U13811 (N_13811,N_6328,N_9640);
nor U13812 (N_13812,N_9651,N_5666);
and U13813 (N_13813,N_8097,N_7629);
or U13814 (N_13814,N_6763,N_7998);
nand U13815 (N_13815,N_9123,N_8779);
nand U13816 (N_13816,N_9227,N_7656);
nand U13817 (N_13817,N_5209,N_9073);
and U13818 (N_13818,N_8257,N_7693);
and U13819 (N_13819,N_5607,N_9739);
nand U13820 (N_13820,N_5628,N_5698);
or U13821 (N_13821,N_6916,N_9718);
nor U13822 (N_13822,N_5311,N_9201);
and U13823 (N_13823,N_7036,N_9933);
nor U13824 (N_13824,N_6764,N_5801);
and U13825 (N_13825,N_8173,N_7333);
nor U13826 (N_13826,N_9649,N_9044);
and U13827 (N_13827,N_6552,N_8075);
and U13828 (N_13828,N_8179,N_5096);
and U13829 (N_13829,N_7603,N_9498);
nand U13830 (N_13830,N_9313,N_7666);
and U13831 (N_13831,N_9245,N_7087);
or U13832 (N_13832,N_7438,N_8768);
or U13833 (N_13833,N_9400,N_9158);
nand U13834 (N_13834,N_8434,N_6804);
nor U13835 (N_13835,N_5641,N_5803);
nand U13836 (N_13836,N_5530,N_6362);
nand U13837 (N_13837,N_6978,N_6003);
nand U13838 (N_13838,N_7602,N_6093);
and U13839 (N_13839,N_6306,N_6716);
nor U13840 (N_13840,N_5450,N_7693);
or U13841 (N_13841,N_8262,N_6920);
nand U13842 (N_13842,N_9068,N_9829);
nor U13843 (N_13843,N_7120,N_6659);
and U13844 (N_13844,N_6319,N_6312);
or U13845 (N_13845,N_7824,N_5216);
nor U13846 (N_13846,N_6077,N_8178);
and U13847 (N_13847,N_6697,N_8571);
nand U13848 (N_13848,N_5424,N_7892);
nand U13849 (N_13849,N_9115,N_7893);
nor U13850 (N_13850,N_6380,N_6244);
or U13851 (N_13851,N_5835,N_9903);
nand U13852 (N_13852,N_8234,N_5625);
nand U13853 (N_13853,N_7810,N_5767);
or U13854 (N_13854,N_9915,N_7311);
and U13855 (N_13855,N_6452,N_8869);
nand U13856 (N_13856,N_8565,N_6536);
and U13857 (N_13857,N_7273,N_5785);
nor U13858 (N_13858,N_8706,N_8789);
or U13859 (N_13859,N_6967,N_8942);
nor U13860 (N_13860,N_7557,N_6471);
or U13861 (N_13861,N_7140,N_7511);
or U13862 (N_13862,N_6099,N_7347);
nor U13863 (N_13863,N_5735,N_8988);
and U13864 (N_13864,N_8509,N_9804);
or U13865 (N_13865,N_7143,N_8953);
and U13866 (N_13866,N_9488,N_7096);
nor U13867 (N_13867,N_7330,N_6987);
or U13868 (N_13868,N_7866,N_6367);
or U13869 (N_13869,N_5392,N_8410);
or U13870 (N_13870,N_6328,N_7067);
xnor U13871 (N_13871,N_7029,N_5179);
nand U13872 (N_13872,N_9469,N_6426);
and U13873 (N_13873,N_6588,N_7801);
or U13874 (N_13874,N_6980,N_7826);
nor U13875 (N_13875,N_8134,N_9850);
nor U13876 (N_13876,N_6360,N_9076);
nand U13877 (N_13877,N_6953,N_6898);
nor U13878 (N_13878,N_6709,N_7757);
nand U13879 (N_13879,N_7875,N_5964);
nor U13880 (N_13880,N_6840,N_6909);
and U13881 (N_13881,N_6351,N_7091);
or U13882 (N_13882,N_7498,N_9127);
nand U13883 (N_13883,N_9213,N_7458);
or U13884 (N_13884,N_7899,N_6110);
nand U13885 (N_13885,N_7091,N_8944);
and U13886 (N_13886,N_6560,N_5036);
nor U13887 (N_13887,N_8231,N_5022);
nand U13888 (N_13888,N_7053,N_8579);
nand U13889 (N_13889,N_6396,N_7276);
or U13890 (N_13890,N_9138,N_7957);
and U13891 (N_13891,N_8045,N_5357);
and U13892 (N_13892,N_8763,N_5168);
nand U13893 (N_13893,N_5101,N_8170);
and U13894 (N_13894,N_7765,N_8712);
and U13895 (N_13895,N_7630,N_5235);
and U13896 (N_13896,N_6908,N_5611);
nor U13897 (N_13897,N_7465,N_9111);
or U13898 (N_13898,N_5894,N_5917);
nor U13899 (N_13899,N_6761,N_8266);
nor U13900 (N_13900,N_9731,N_6876);
nor U13901 (N_13901,N_7982,N_8261);
or U13902 (N_13902,N_6836,N_9463);
nor U13903 (N_13903,N_5584,N_6087);
or U13904 (N_13904,N_7618,N_7148);
nor U13905 (N_13905,N_9430,N_6988);
or U13906 (N_13906,N_8310,N_5396);
and U13907 (N_13907,N_6953,N_8320);
nor U13908 (N_13908,N_6709,N_5954);
nor U13909 (N_13909,N_9783,N_6264);
and U13910 (N_13910,N_5542,N_9126);
and U13911 (N_13911,N_7250,N_5974);
nand U13912 (N_13912,N_9673,N_5153);
nand U13913 (N_13913,N_5387,N_8400);
nand U13914 (N_13914,N_8286,N_8383);
nor U13915 (N_13915,N_5601,N_5042);
or U13916 (N_13916,N_7985,N_9498);
nor U13917 (N_13917,N_8656,N_8374);
or U13918 (N_13918,N_9744,N_6803);
or U13919 (N_13919,N_8535,N_9784);
or U13920 (N_13920,N_6256,N_6866);
or U13921 (N_13921,N_7272,N_7244);
or U13922 (N_13922,N_9177,N_7583);
and U13923 (N_13923,N_8457,N_7112);
nor U13924 (N_13924,N_6904,N_6654);
or U13925 (N_13925,N_7690,N_5710);
or U13926 (N_13926,N_7801,N_5293);
or U13927 (N_13927,N_9204,N_5965);
and U13928 (N_13928,N_6463,N_8700);
and U13929 (N_13929,N_8722,N_5035);
and U13930 (N_13930,N_8007,N_7050);
and U13931 (N_13931,N_5358,N_5962);
and U13932 (N_13932,N_9912,N_5672);
and U13933 (N_13933,N_6055,N_8622);
nor U13934 (N_13934,N_5547,N_7781);
xor U13935 (N_13935,N_5957,N_6631);
nand U13936 (N_13936,N_8882,N_9282);
nor U13937 (N_13937,N_8861,N_9047);
or U13938 (N_13938,N_5710,N_9558);
nand U13939 (N_13939,N_9029,N_6231);
nand U13940 (N_13940,N_8970,N_6967);
nor U13941 (N_13941,N_7816,N_9956);
nor U13942 (N_13942,N_8931,N_5584);
nor U13943 (N_13943,N_7314,N_8060);
or U13944 (N_13944,N_8443,N_9294);
nand U13945 (N_13945,N_5154,N_5376);
and U13946 (N_13946,N_9041,N_9660);
and U13947 (N_13947,N_9556,N_6242);
nor U13948 (N_13948,N_8323,N_6301);
or U13949 (N_13949,N_9988,N_6230);
nor U13950 (N_13950,N_6200,N_8559);
or U13951 (N_13951,N_8796,N_5754);
xor U13952 (N_13952,N_7850,N_9515);
nor U13953 (N_13953,N_7996,N_8664);
nand U13954 (N_13954,N_8488,N_5465);
and U13955 (N_13955,N_9574,N_9588);
and U13956 (N_13956,N_7023,N_8716);
nand U13957 (N_13957,N_5254,N_6621);
and U13958 (N_13958,N_7714,N_5825);
nand U13959 (N_13959,N_9129,N_8098);
or U13960 (N_13960,N_8173,N_5772);
or U13961 (N_13961,N_5969,N_5156);
or U13962 (N_13962,N_8119,N_5512);
nand U13963 (N_13963,N_7541,N_8178);
and U13964 (N_13964,N_6672,N_6256);
and U13965 (N_13965,N_8292,N_5846);
nand U13966 (N_13966,N_8990,N_7209);
or U13967 (N_13967,N_6010,N_7824);
and U13968 (N_13968,N_7353,N_7134);
or U13969 (N_13969,N_9325,N_6658);
or U13970 (N_13970,N_7050,N_7209);
xnor U13971 (N_13971,N_7257,N_5347);
nand U13972 (N_13972,N_8575,N_9869);
and U13973 (N_13973,N_6105,N_5657);
or U13974 (N_13974,N_8890,N_7440);
and U13975 (N_13975,N_7398,N_8314);
or U13976 (N_13976,N_8553,N_6827);
and U13977 (N_13977,N_8871,N_5394);
nor U13978 (N_13978,N_7314,N_8380);
and U13979 (N_13979,N_9953,N_6680);
nand U13980 (N_13980,N_9103,N_6357);
nand U13981 (N_13981,N_9810,N_7012);
nor U13982 (N_13982,N_6114,N_8890);
or U13983 (N_13983,N_9908,N_7598);
or U13984 (N_13984,N_5379,N_7100);
or U13985 (N_13985,N_5704,N_9120);
nand U13986 (N_13986,N_8480,N_5100);
and U13987 (N_13987,N_5758,N_8748);
nand U13988 (N_13988,N_8235,N_8964);
nand U13989 (N_13989,N_7114,N_9035);
or U13990 (N_13990,N_8997,N_9160);
nor U13991 (N_13991,N_5462,N_7561);
or U13992 (N_13992,N_6743,N_5104);
nor U13993 (N_13993,N_9851,N_7727);
nand U13994 (N_13994,N_8556,N_9316);
and U13995 (N_13995,N_9320,N_8525);
nor U13996 (N_13996,N_5767,N_7147);
and U13997 (N_13997,N_9872,N_7151);
nor U13998 (N_13998,N_8791,N_8960);
nor U13999 (N_13999,N_6435,N_9160);
or U14000 (N_14000,N_6774,N_9143);
or U14001 (N_14001,N_7067,N_9821);
nor U14002 (N_14002,N_9068,N_7910);
and U14003 (N_14003,N_9421,N_8836);
nor U14004 (N_14004,N_9144,N_8072);
or U14005 (N_14005,N_7926,N_8993);
and U14006 (N_14006,N_8692,N_7107);
nor U14007 (N_14007,N_8681,N_9840);
and U14008 (N_14008,N_5902,N_9385);
nand U14009 (N_14009,N_5186,N_6386);
nand U14010 (N_14010,N_5822,N_8440);
or U14011 (N_14011,N_9962,N_6765);
and U14012 (N_14012,N_9513,N_6662);
or U14013 (N_14013,N_6665,N_9532);
and U14014 (N_14014,N_5306,N_7438);
nor U14015 (N_14015,N_9908,N_7263);
or U14016 (N_14016,N_6062,N_9845);
nand U14017 (N_14017,N_9845,N_8583);
nor U14018 (N_14018,N_8270,N_8568);
or U14019 (N_14019,N_6287,N_7316);
xor U14020 (N_14020,N_9817,N_8787);
nor U14021 (N_14021,N_5413,N_5806);
nand U14022 (N_14022,N_5595,N_9808);
or U14023 (N_14023,N_8925,N_7492);
and U14024 (N_14024,N_6524,N_7268);
or U14025 (N_14025,N_5937,N_8693);
nor U14026 (N_14026,N_9778,N_8824);
nor U14027 (N_14027,N_5663,N_5824);
or U14028 (N_14028,N_7593,N_7582);
nand U14029 (N_14029,N_8391,N_7966);
or U14030 (N_14030,N_8700,N_8261);
or U14031 (N_14031,N_8595,N_5525);
or U14032 (N_14032,N_8852,N_5281);
and U14033 (N_14033,N_7958,N_8245);
nor U14034 (N_14034,N_9078,N_5079);
nor U14035 (N_14035,N_7753,N_8601);
nor U14036 (N_14036,N_9529,N_8904);
or U14037 (N_14037,N_7755,N_6770);
nand U14038 (N_14038,N_5245,N_5438);
nor U14039 (N_14039,N_8262,N_7168);
nor U14040 (N_14040,N_9499,N_9968);
nor U14041 (N_14041,N_8888,N_5397);
and U14042 (N_14042,N_7335,N_9839);
or U14043 (N_14043,N_5390,N_8638);
nor U14044 (N_14044,N_6727,N_5743);
nor U14045 (N_14045,N_8500,N_5026);
nand U14046 (N_14046,N_5033,N_8310);
or U14047 (N_14047,N_8927,N_6472);
and U14048 (N_14048,N_8279,N_9256);
and U14049 (N_14049,N_9327,N_6921);
nand U14050 (N_14050,N_8369,N_9006);
xor U14051 (N_14051,N_6651,N_7463);
nand U14052 (N_14052,N_6720,N_6232);
or U14053 (N_14053,N_7812,N_9967);
nor U14054 (N_14054,N_8468,N_9689);
nor U14055 (N_14055,N_5711,N_8959);
nor U14056 (N_14056,N_7842,N_9019);
or U14057 (N_14057,N_5265,N_7100);
nor U14058 (N_14058,N_9559,N_7250);
or U14059 (N_14059,N_6837,N_8185);
and U14060 (N_14060,N_8438,N_7708);
or U14061 (N_14061,N_9660,N_7325);
and U14062 (N_14062,N_8629,N_9858);
and U14063 (N_14063,N_7918,N_8156);
nor U14064 (N_14064,N_6568,N_7597);
nand U14065 (N_14065,N_5008,N_7303);
or U14066 (N_14066,N_8920,N_8881);
nor U14067 (N_14067,N_8524,N_7224);
or U14068 (N_14068,N_9633,N_8509);
nand U14069 (N_14069,N_7384,N_7573);
or U14070 (N_14070,N_5995,N_7382);
nand U14071 (N_14071,N_6044,N_7269);
nand U14072 (N_14072,N_5658,N_5199);
or U14073 (N_14073,N_7027,N_5116);
nor U14074 (N_14074,N_8672,N_7866);
nand U14075 (N_14075,N_9747,N_7950);
nor U14076 (N_14076,N_8523,N_6927);
nand U14077 (N_14077,N_6355,N_8919);
or U14078 (N_14078,N_7801,N_9190);
and U14079 (N_14079,N_7609,N_6677);
nor U14080 (N_14080,N_6529,N_8701);
or U14081 (N_14081,N_8620,N_7224);
nand U14082 (N_14082,N_9769,N_7251);
or U14083 (N_14083,N_7496,N_7543);
nor U14084 (N_14084,N_5939,N_6720);
xor U14085 (N_14085,N_8867,N_8105);
nor U14086 (N_14086,N_6031,N_9455);
nor U14087 (N_14087,N_7187,N_8304);
nand U14088 (N_14088,N_5378,N_5307);
nor U14089 (N_14089,N_9798,N_7317);
nand U14090 (N_14090,N_5217,N_6968);
nor U14091 (N_14091,N_7308,N_9519);
or U14092 (N_14092,N_9770,N_9544);
nor U14093 (N_14093,N_5869,N_6973);
or U14094 (N_14094,N_6692,N_9013);
nor U14095 (N_14095,N_5111,N_5881);
nor U14096 (N_14096,N_6066,N_8566);
nor U14097 (N_14097,N_8147,N_6970);
and U14098 (N_14098,N_9755,N_9559);
nor U14099 (N_14099,N_5911,N_8840);
and U14100 (N_14100,N_9232,N_6702);
nor U14101 (N_14101,N_6394,N_9980);
and U14102 (N_14102,N_6269,N_6120);
nand U14103 (N_14103,N_6457,N_7106);
or U14104 (N_14104,N_8954,N_6601);
and U14105 (N_14105,N_5808,N_7824);
nor U14106 (N_14106,N_8665,N_6290);
and U14107 (N_14107,N_5445,N_9133);
nor U14108 (N_14108,N_9879,N_9562);
and U14109 (N_14109,N_7579,N_8474);
nor U14110 (N_14110,N_9411,N_7930);
nor U14111 (N_14111,N_8690,N_8651);
and U14112 (N_14112,N_6655,N_9555);
nand U14113 (N_14113,N_6114,N_5726);
nor U14114 (N_14114,N_7674,N_5721);
nor U14115 (N_14115,N_7134,N_6002);
or U14116 (N_14116,N_9376,N_8770);
and U14117 (N_14117,N_5294,N_6979);
nand U14118 (N_14118,N_7025,N_9265);
or U14119 (N_14119,N_5853,N_5891);
and U14120 (N_14120,N_8832,N_6879);
nor U14121 (N_14121,N_9651,N_6115);
or U14122 (N_14122,N_9506,N_8979);
nor U14123 (N_14123,N_7423,N_5515);
or U14124 (N_14124,N_9608,N_5170);
nor U14125 (N_14125,N_5605,N_9346);
nand U14126 (N_14126,N_7168,N_9881);
nand U14127 (N_14127,N_7432,N_7490);
or U14128 (N_14128,N_6435,N_8664);
nand U14129 (N_14129,N_7896,N_5511);
nand U14130 (N_14130,N_7402,N_6553);
and U14131 (N_14131,N_5868,N_7659);
nand U14132 (N_14132,N_6294,N_9631);
nor U14133 (N_14133,N_7638,N_6637);
and U14134 (N_14134,N_6881,N_6955);
nor U14135 (N_14135,N_5553,N_5749);
nand U14136 (N_14136,N_7831,N_9000);
or U14137 (N_14137,N_5334,N_6505);
nor U14138 (N_14138,N_8775,N_9758);
nand U14139 (N_14139,N_5185,N_7372);
nor U14140 (N_14140,N_5077,N_9647);
and U14141 (N_14141,N_6732,N_6805);
nand U14142 (N_14142,N_8128,N_5563);
or U14143 (N_14143,N_7561,N_5953);
or U14144 (N_14144,N_8882,N_6116);
nor U14145 (N_14145,N_5205,N_8050);
or U14146 (N_14146,N_5625,N_9565);
nor U14147 (N_14147,N_8028,N_9975);
nor U14148 (N_14148,N_5969,N_9681);
nor U14149 (N_14149,N_7512,N_8503);
nor U14150 (N_14150,N_8734,N_8026);
nand U14151 (N_14151,N_9806,N_9646);
and U14152 (N_14152,N_7029,N_8867);
nand U14153 (N_14153,N_9187,N_6107);
or U14154 (N_14154,N_7159,N_5055);
or U14155 (N_14155,N_8601,N_9735);
nand U14156 (N_14156,N_6716,N_9996);
nand U14157 (N_14157,N_5754,N_9730);
nor U14158 (N_14158,N_6469,N_8362);
or U14159 (N_14159,N_6254,N_6953);
nand U14160 (N_14160,N_7601,N_9414);
or U14161 (N_14161,N_6050,N_5796);
or U14162 (N_14162,N_5754,N_5343);
and U14163 (N_14163,N_7057,N_6080);
nand U14164 (N_14164,N_9010,N_8856);
and U14165 (N_14165,N_8849,N_6825);
or U14166 (N_14166,N_5773,N_7436);
nand U14167 (N_14167,N_7219,N_9997);
and U14168 (N_14168,N_6240,N_8915);
nand U14169 (N_14169,N_7534,N_9360);
nor U14170 (N_14170,N_6182,N_5935);
nor U14171 (N_14171,N_8223,N_6325);
or U14172 (N_14172,N_9561,N_6888);
or U14173 (N_14173,N_5571,N_5490);
and U14174 (N_14174,N_7695,N_7206);
and U14175 (N_14175,N_8083,N_6063);
nor U14176 (N_14176,N_8271,N_6210);
nor U14177 (N_14177,N_7274,N_6903);
nand U14178 (N_14178,N_5558,N_5850);
and U14179 (N_14179,N_6485,N_7151);
or U14180 (N_14180,N_8826,N_5345);
and U14181 (N_14181,N_5131,N_5238);
or U14182 (N_14182,N_7482,N_5461);
or U14183 (N_14183,N_5160,N_6740);
or U14184 (N_14184,N_9081,N_7630);
nor U14185 (N_14185,N_5488,N_9500);
or U14186 (N_14186,N_7810,N_6692);
nand U14187 (N_14187,N_8557,N_7924);
nor U14188 (N_14188,N_5192,N_6299);
nand U14189 (N_14189,N_8358,N_6587);
and U14190 (N_14190,N_7696,N_5762);
or U14191 (N_14191,N_9343,N_6936);
and U14192 (N_14192,N_9656,N_7712);
and U14193 (N_14193,N_8968,N_6079);
nand U14194 (N_14194,N_6922,N_7076);
xor U14195 (N_14195,N_8994,N_6663);
nand U14196 (N_14196,N_7681,N_9013);
or U14197 (N_14197,N_8964,N_9563);
nor U14198 (N_14198,N_8302,N_6085);
or U14199 (N_14199,N_6627,N_7188);
or U14200 (N_14200,N_7329,N_7913);
or U14201 (N_14201,N_8417,N_5454);
or U14202 (N_14202,N_8896,N_6265);
nor U14203 (N_14203,N_5617,N_5494);
nor U14204 (N_14204,N_9974,N_7049);
or U14205 (N_14205,N_9038,N_6035);
and U14206 (N_14206,N_8783,N_9436);
nand U14207 (N_14207,N_9748,N_5886);
and U14208 (N_14208,N_9091,N_7639);
nand U14209 (N_14209,N_5894,N_6016);
nor U14210 (N_14210,N_7850,N_7573);
and U14211 (N_14211,N_9553,N_9436);
nand U14212 (N_14212,N_5065,N_9666);
or U14213 (N_14213,N_5684,N_5570);
or U14214 (N_14214,N_7887,N_9721);
or U14215 (N_14215,N_5009,N_9952);
and U14216 (N_14216,N_5270,N_8280);
nor U14217 (N_14217,N_5436,N_7343);
nand U14218 (N_14218,N_7279,N_9097);
xnor U14219 (N_14219,N_5057,N_7749);
nand U14220 (N_14220,N_8176,N_7666);
or U14221 (N_14221,N_9805,N_6384);
and U14222 (N_14222,N_7807,N_8734);
nand U14223 (N_14223,N_9447,N_9778);
and U14224 (N_14224,N_8597,N_7917);
nand U14225 (N_14225,N_5869,N_7452);
or U14226 (N_14226,N_5994,N_9455);
nand U14227 (N_14227,N_8979,N_9336);
nand U14228 (N_14228,N_8664,N_8610);
nand U14229 (N_14229,N_8364,N_8067);
nor U14230 (N_14230,N_8334,N_9210);
or U14231 (N_14231,N_8088,N_7875);
and U14232 (N_14232,N_8604,N_6903);
and U14233 (N_14233,N_6365,N_9299);
nor U14234 (N_14234,N_6632,N_6001);
and U14235 (N_14235,N_6426,N_6882);
nand U14236 (N_14236,N_7353,N_8536);
or U14237 (N_14237,N_8744,N_6554);
or U14238 (N_14238,N_5752,N_9929);
or U14239 (N_14239,N_7172,N_9258);
nor U14240 (N_14240,N_7269,N_9970);
nand U14241 (N_14241,N_6128,N_9906);
nand U14242 (N_14242,N_5843,N_9397);
and U14243 (N_14243,N_5888,N_9183);
nor U14244 (N_14244,N_9950,N_8705);
or U14245 (N_14245,N_6470,N_9485);
and U14246 (N_14246,N_6829,N_7466);
nand U14247 (N_14247,N_8030,N_5279);
and U14248 (N_14248,N_9191,N_6098);
nor U14249 (N_14249,N_6217,N_5563);
and U14250 (N_14250,N_5251,N_6670);
or U14251 (N_14251,N_5681,N_7367);
and U14252 (N_14252,N_5806,N_7171);
or U14253 (N_14253,N_8013,N_7643);
and U14254 (N_14254,N_8295,N_6748);
nor U14255 (N_14255,N_6413,N_8814);
or U14256 (N_14256,N_9666,N_6142);
nor U14257 (N_14257,N_8562,N_9751);
or U14258 (N_14258,N_7517,N_8960);
and U14259 (N_14259,N_8853,N_6228);
nor U14260 (N_14260,N_5254,N_9980);
and U14261 (N_14261,N_6220,N_9875);
or U14262 (N_14262,N_9696,N_7503);
nor U14263 (N_14263,N_9365,N_7728);
nand U14264 (N_14264,N_6481,N_9673);
nor U14265 (N_14265,N_6122,N_5584);
nand U14266 (N_14266,N_8568,N_7637);
and U14267 (N_14267,N_5619,N_8433);
nand U14268 (N_14268,N_6036,N_5583);
or U14269 (N_14269,N_5727,N_7918);
or U14270 (N_14270,N_7849,N_9297);
nor U14271 (N_14271,N_6067,N_9643);
or U14272 (N_14272,N_7795,N_6990);
nand U14273 (N_14273,N_6303,N_6220);
nor U14274 (N_14274,N_8794,N_8337);
nor U14275 (N_14275,N_7921,N_9784);
and U14276 (N_14276,N_9018,N_8440);
nand U14277 (N_14277,N_7844,N_6624);
nor U14278 (N_14278,N_6092,N_6150);
nor U14279 (N_14279,N_9141,N_5342);
nor U14280 (N_14280,N_5225,N_5714);
or U14281 (N_14281,N_9704,N_8301);
and U14282 (N_14282,N_5525,N_5364);
nand U14283 (N_14283,N_5347,N_6037);
nor U14284 (N_14284,N_9092,N_6047);
and U14285 (N_14285,N_7511,N_7184);
and U14286 (N_14286,N_7785,N_8138);
or U14287 (N_14287,N_8223,N_8604);
or U14288 (N_14288,N_8857,N_5564);
nand U14289 (N_14289,N_5577,N_9872);
or U14290 (N_14290,N_6773,N_9223);
nor U14291 (N_14291,N_5817,N_7483);
nand U14292 (N_14292,N_5231,N_5518);
and U14293 (N_14293,N_9603,N_5185);
and U14294 (N_14294,N_5588,N_8648);
nand U14295 (N_14295,N_5177,N_5557);
nand U14296 (N_14296,N_9494,N_9631);
nand U14297 (N_14297,N_7471,N_6321);
nand U14298 (N_14298,N_8926,N_5508);
nor U14299 (N_14299,N_8804,N_9307);
or U14300 (N_14300,N_5694,N_7317);
or U14301 (N_14301,N_8627,N_9640);
or U14302 (N_14302,N_7719,N_7797);
nand U14303 (N_14303,N_8855,N_9444);
nor U14304 (N_14304,N_6872,N_6562);
nor U14305 (N_14305,N_8771,N_8914);
nor U14306 (N_14306,N_5776,N_6446);
nand U14307 (N_14307,N_6601,N_8852);
xnor U14308 (N_14308,N_5475,N_8660);
or U14309 (N_14309,N_7423,N_7090);
nor U14310 (N_14310,N_7575,N_5893);
nor U14311 (N_14311,N_6383,N_5487);
or U14312 (N_14312,N_7417,N_8816);
and U14313 (N_14313,N_6750,N_6295);
and U14314 (N_14314,N_8375,N_6503);
nor U14315 (N_14315,N_6633,N_5122);
nor U14316 (N_14316,N_5980,N_6789);
and U14317 (N_14317,N_5097,N_5630);
or U14318 (N_14318,N_7165,N_8675);
nand U14319 (N_14319,N_7206,N_6242);
nor U14320 (N_14320,N_6031,N_5694);
nand U14321 (N_14321,N_7173,N_6246);
or U14322 (N_14322,N_5030,N_5050);
and U14323 (N_14323,N_5890,N_6833);
nand U14324 (N_14324,N_8835,N_9152);
or U14325 (N_14325,N_7578,N_7406);
and U14326 (N_14326,N_9878,N_8079);
nand U14327 (N_14327,N_7694,N_5200);
nand U14328 (N_14328,N_9174,N_9198);
nand U14329 (N_14329,N_6481,N_5133);
nand U14330 (N_14330,N_8159,N_9359);
and U14331 (N_14331,N_6670,N_5867);
nand U14332 (N_14332,N_5320,N_9955);
and U14333 (N_14333,N_8065,N_7179);
nor U14334 (N_14334,N_7383,N_6442);
or U14335 (N_14335,N_8980,N_9734);
nor U14336 (N_14336,N_5135,N_5862);
nor U14337 (N_14337,N_6626,N_6890);
and U14338 (N_14338,N_7395,N_6771);
or U14339 (N_14339,N_6574,N_6192);
and U14340 (N_14340,N_7003,N_6578);
nand U14341 (N_14341,N_7013,N_8804);
nand U14342 (N_14342,N_5493,N_8860);
nand U14343 (N_14343,N_7929,N_5477);
nor U14344 (N_14344,N_9626,N_9055);
and U14345 (N_14345,N_5768,N_8671);
nand U14346 (N_14346,N_9272,N_9443);
or U14347 (N_14347,N_7118,N_6461);
nor U14348 (N_14348,N_5056,N_7448);
and U14349 (N_14349,N_6860,N_9830);
or U14350 (N_14350,N_9605,N_6462);
and U14351 (N_14351,N_5880,N_9211);
nand U14352 (N_14352,N_5593,N_9640);
nor U14353 (N_14353,N_7643,N_7739);
and U14354 (N_14354,N_5094,N_8304);
and U14355 (N_14355,N_5191,N_6420);
or U14356 (N_14356,N_9216,N_7122);
nor U14357 (N_14357,N_6045,N_6161);
nand U14358 (N_14358,N_5829,N_6847);
and U14359 (N_14359,N_6767,N_5659);
and U14360 (N_14360,N_8792,N_9943);
nand U14361 (N_14361,N_8890,N_8010);
and U14362 (N_14362,N_5264,N_5002);
nor U14363 (N_14363,N_7983,N_5762);
nor U14364 (N_14364,N_6167,N_6251);
or U14365 (N_14365,N_8515,N_6808);
and U14366 (N_14366,N_5436,N_8771);
nand U14367 (N_14367,N_8210,N_5437);
nand U14368 (N_14368,N_7719,N_8413);
and U14369 (N_14369,N_7508,N_6194);
nor U14370 (N_14370,N_6268,N_7311);
and U14371 (N_14371,N_9574,N_8707);
nand U14372 (N_14372,N_5865,N_5266);
or U14373 (N_14373,N_7237,N_8669);
nor U14374 (N_14374,N_9871,N_7401);
nor U14375 (N_14375,N_9635,N_8564);
or U14376 (N_14376,N_9430,N_6566);
nor U14377 (N_14377,N_7860,N_5402);
or U14378 (N_14378,N_8063,N_5108);
nor U14379 (N_14379,N_8470,N_6110);
nor U14380 (N_14380,N_5257,N_6383);
and U14381 (N_14381,N_8577,N_6608);
and U14382 (N_14382,N_9464,N_5520);
nand U14383 (N_14383,N_8149,N_6240);
nand U14384 (N_14384,N_9462,N_6213);
or U14385 (N_14385,N_8294,N_9973);
or U14386 (N_14386,N_9279,N_9602);
or U14387 (N_14387,N_7574,N_8060);
nor U14388 (N_14388,N_9384,N_9317);
nand U14389 (N_14389,N_7221,N_8673);
nor U14390 (N_14390,N_6372,N_7811);
nand U14391 (N_14391,N_7417,N_9723);
and U14392 (N_14392,N_7143,N_9660);
nor U14393 (N_14393,N_5043,N_7540);
nand U14394 (N_14394,N_8716,N_8154);
and U14395 (N_14395,N_9452,N_9987);
or U14396 (N_14396,N_6523,N_8211);
nor U14397 (N_14397,N_6929,N_9541);
or U14398 (N_14398,N_8319,N_6367);
or U14399 (N_14399,N_6722,N_6430);
nand U14400 (N_14400,N_9354,N_6957);
or U14401 (N_14401,N_6030,N_7475);
or U14402 (N_14402,N_7514,N_9390);
nand U14403 (N_14403,N_7969,N_5306);
nand U14404 (N_14404,N_5276,N_5960);
nor U14405 (N_14405,N_7434,N_6592);
and U14406 (N_14406,N_5490,N_6831);
and U14407 (N_14407,N_8215,N_5348);
or U14408 (N_14408,N_5658,N_6809);
nand U14409 (N_14409,N_7736,N_6111);
nand U14410 (N_14410,N_8939,N_5559);
or U14411 (N_14411,N_5947,N_9391);
and U14412 (N_14412,N_6439,N_9793);
and U14413 (N_14413,N_5120,N_5591);
or U14414 (N_14414,N_7294,N_8060);
nand U14415 (N_14415,N_5609,N_7180);
and U14416 (N_14416,N_9461,N_8903);
or U14417 (N_14417,N_7184,N_7898);
nor U14418 (N_14418,N_7259,N_7994);
and U14419 (N_14419,N_8550,N_9598);
nand U14420 (N_14420,N_7611,N_9676);
and U14421 (N_14421,N_8852,N_5736);
and U14422 (N_14422,N_5134,N_5723);
nand U14423 (N_14423,N_5832,N_5200);
nor U14424 (N_14424,N_5896,N_7901);
or U14425 (N_14425,N_5784,N_8971);
nor U14426 (N_14426,N_8682,N_6807);
or U14427 (N_14427,N_8202,N_8249);
nand U14428 (N_14428,N_9200,N_7468);
nor U14429 (N_14429,N_6454,N_9922);
or U14430 (N_14430,N_9097,N_9271);
xnor U14431 (N_14431,N_7076,N_6186);
nor U14432 (N_14432,N_9358,N_5342);
nand U14433 (N_14433,N_6362,N_6277);
and U14434 (N_14434,N_6647,N_5686);
nor U14435 (N_14435,N_5747,N_6729);
or U14436 (N_14436,N_5579,N_6783);
nor U14437 (N_14437,N_6077,N_8765);
and U14438 (N_14438,N_7835,N_5701);
or U14439 (N_14439,N_5685,N_9133);
nand U14440 (N_14440,N_6018,N_7381);
and U14441 (N_14441,N_8120,N_7617);
or U14442 (N_14442,N_8724,N_7342);
nand U14443 (N_14443,N_9015,N_7098);
and U14444 (N_14444,N_6003,N_5695);
and U14445 (N_14445,N_6454,N_9183);
nor U14446 (N_14446,N_6526,N_9350);
nand U14447 (N_14447,N_9075,N_5760);
or U14448 (N_14448,N_7215,N_5406);
nand U14449 (N_14449,N_5898,N_7841);
nor U14450 (N_14450,N_8324,N_7418);
or U14451 (N_14451,N_8856,N_6465);
nand U14452 (N_14452,N_8235,N_7080);
nand U14453 (N_14453,N_8845,N_8868);
nand U14454 (N_14454,N_6403,N_5467);
or U14455 (N_14455,N_7582,N_7496);
and U14456 (N_14456,N_7452,N_9989);
nor U14457 (N_14457,N_7238,N_9305);
nand U14458 (N_14458,N_6343,N_6250);
and U14459 (N_14459,N_5941,N_7130);
nand U14460 (N_14460,N_7749,N_7020);
or U14461 (N_14461,N_9949,N_6455);
and U14462 (N_14462,N_9186,N_8698);
and U14463 (N_14463,N_6788,N_8379);
nand U14464 (N_14464,N_5149,N_7282);
or U14465 (N_14465,N_9415,N_5735);
nand U14466 (N_14466,N_6578,N_7250);
or U14467 (N_14467,N_6267,N_5371);
and U14468 (N_14468,N_5687,N_6927);
nand U14469 (N_14469,N_6553,N_9036);
nand U14470 (N_14470,N_8951,N_5213);
and U14471 (N_14471,N_9898,N_5229);
nor U14472 (N_14472,N_8086,N_8713);
xnor U14473 (N_14473,N_6746,N_5333);
nor U14474 (N_14474,N_7346,N_7234);
or U14475 (N_14475,N_9415,N_9856);
nand U14476 (N_14476,N_7055,N_8899);
and U14477 (N_14477,N_9002,N_8317);
or U14478 (N_14478,N_6095,N_5632);
nor U14479 (N_14479,N_6016,N_5200);
or U14480 (N_14480,N_5971,N_5986);
and U14481 (N_14481,N_7449,N_8389);
or U14482 (N_14482,N_9190,N_8090);
and U14483 (N_14483,N_9609,N_8325);
or U14484 (N_14484,N_8258,N_9434);
nand U14485 (N_14485,N_7822,N_8978);
nand U14486 (N_14486,N_8864,N_6577);
nand U14487 (N_14487,N_5759,N_9430);
and U14488 (N_14488,N_9199,N_6967);
and U14489 (N_14489,N_8459,N_7129);
or U14490 (N_14490,N_9709,N_9794);
nor U14491 (N_14491,N_6354,N_6875);
nor U14492 (N_14492,N_5889,N_8438);
and U14493 (N_14493,N_7709,N_5809);
or U14494 (N_14494,N_5806,N_9877);
or U14495 (N_14495,N_8015,N_5392);
or U14496 (N_14496,N_5003,N_8370);
or U14497 (N_14497,N_5141,N_5007);
nand U14498 (N_14498,N_8106,N_9610);
and U14499 (N_14499,N_8917,N_9981);
or U14500 (N_14500,N_5330,N_9803);
and U14501 (N_14501,N_6996,N_9227);
nor U14502 (N_14502,N_9240,N_6263);
or U14503 (N_14503,N_7935,N_7489);
nand U14504 (N_14504,N_9823,N_7935);
nand U14505 (N_14505,N_7789,N_9340);
nand U14506 (N_14506,N_8743,N_5712);
nor U14507 (N_14507,N_6211,N_9973);
or U14508 (N_14508,N_6087,N_8068);
nand U14509 (N_14509,N_8533,N_6387);
and U14510 (N_14510,N_7536,N_5006);
and U14511 (N_14511,N_5994,N_5601);
or U14512 (N_14512,N_6403,N_6331);
nor U14513 (N_14513,N_8495,N_8681);
or U14514 (N_14514,N_8108,N_6436);
and U14515 (N_14515,N_6431,N_9502);
and U14516 (N_14516,N_7682,N_8144);
or U14517 (N_14517,N_5671,N_6786);
nor U14518 (N_14518,N_9183,N_5810);
nand U14519 (N_14519,N_6624,N_9558);
nor U14520 (N_14520,N_8820,N_8869);
nor U14521 (N_14521,N_7515,N_6779);
or U14522 (N_14522,N_6631,N_6739);
or U14523 (N_14523,N_8191,N_9764);
or U14524 (N_14524,N_8999,N_6181);
and U14525 (N_14525,N_9434,N_6789);
and U14526 (N_14526,N_6884,N_6372);
nor U14527 (N_14527,N_5747,N_6044);
or U14528 (N_14528,N_8190,N_7441);
or U14529 (N_14529,N_7734,N_7045);
nor U14530 (N_14530,N_9942,N_9408);
or U14531 (N_14531,N_5745,N_6433);
nor U14532 (N_14532,N_6949,N_5428);
nand U14533 (N_14533,N_9418,N_8237);
nand U14534 (N_14534,N_7227,N_5990);
or U14535 (N_14535,N_9226,N_6107);
and U14536 (N_14536,N_7231,N_6111);
or U14537 (N_14537,N_7351,N_6209);
nor U14538 (N_14538,N_6012,N_8128);
nor U14539 (N_14539,N_8342,N_6028);
and U14540 (N_14540,N_6103,N_9540);
and U14541 (N_14541,N_7355,N_9188);
or U14542 (N_14542,N_5793,N_9910);
nand U14543 (N_14543,N_8421,N_5027);
nand U14544 (N_14544,N_8773,N_6726);
and U14545 (N_14545,N_9932,N_5052);
or U14546 (N_14546,N_9561,N_8610);
nor U14547 (N_14547,N_8741,N_8176);
nor U14548 (N_14548,N_7807,N_6998);
nor U14549 (N_14549,N_8183,N_5208);
and U14550 (N_14550,N_7791,N_5780);
or U14551 (N_14551,N_5433,N_8504);
nand U14552 (N_14552,N_7894,N_9961);
nor U14553 (N_14553,N_5326,N_7160);
nand U14554 (N_14554,N_8500,N_6192);
nand U14555 (N_14555,N_8690,N_9906);
or U14556 (N_14556,N_7806,N_7695);
nor U14557 (N_14557,N_6635,N_6230);
and U14558 (N_14558,N_6934,N_7416);
nor U14559 (N_14559,N_8923,N_7890);
nand U14560 (N_14560,N_8018,N_9668);
nor U14561 (N_14561,N_5217,N_8734);
and U14562 (N_14562,N_9496,N_5093);
nor U14563 (N_14563,N_5309,N_9919);
or U14564 (N_14564,N_8606,N_5581);
nand U14565 (N_14565,N_6446,N_9624);
or U14566 (N_14566,N_7541,N_9095);
or U14567 (N_14567,N_7979,N_7630);
nand U14568 (N_14568,N_6869,N_8221);
and U14569 (N_14569,N_8721,N_7423);
nand U14570 (N_14570,N_9928,N_6718);
and U14571 (N_14571,N_7435,N_9891);
and U14572 (N_14572,N_9646,N_8907);
or U14573 (N_14573,N_7471,N_7535);
nand U14574 (N_14574,N_9122,N_8115);
nand U14575 (N_14575,N_5101,N_7896);
nand U14576 (N_14576,N_9674,N_8046);
or U14577 (N_14577,N_8701,N_9302);
nand U14578 (N_14578,N_7444,N_9548);
and U14579 (N_14579,N_7349,N_9301);
or U14580 (N_14580,N_9353,N_6819);
nand U14581 (N_14581,N_7813,N_8875);
or U14582 (N_14582,N_9398,N_8698);
or U14583 (N_14583,N_9371,N_9573);
or U14584 (N_14584,N_8367,N_7683);
nor U14585 (N_14585,N_6798,N_9633);
nand U14586 (N_14586,N_7082,N_9516);
nor U14587 (N_14587,N_9871,N_6613);
or U14588 (N_14588,N_8134,N_8084);
nand U14589 (N_14589,N_6717,N_5109);
or U14590 (N_14590,N_9842,N_5941);
or U14591 (N_14591,N_7360,N_8454);
and U14592 (N_14592,N_9648,N_9892);
nand U14593 (N_14593,N_7883,N_9237);
nor U14594 (N_14594,N_8481,N_9523);
nor U14595 (N_14595,N_7448,N_8829);
nand U14596 (N_14596,N_9689,N_9260);
and U14597 (N_14597,N_8867,N_9120);
and U14598 (N_14598,N_8662,N_5810);
nor U14599 (N_14599,N_6969,N_9317);
nand U14600 (N_14600,N_9969,N_5743);
and U14601 (N_14601,N_5621,N_9953);
nor U14602 (N_14602,N_9864,N_7773);
or U14603 (N_14603,N_7871,N_5873);
and U14604 (N_14604,N_6441,N_5480);
and U14605 (N_14605,N_8181,N_8658);
or U14606 (N_14606,N_7314,N_8159);
and U14607 (N_14607,N_8700,N_5659);
and U14608 (N_14608,N_6354,N_9578);
and U14609 (N_14609,N_5894,N_6890);
nand U14610 (N_14610,N_6955,N_5219);
nand U14611 (N_14611,N_9371,N_9315);
nor U14612 (N_14612,N_6019,N_5144);
nand U14613 (N_14613,N_8515,N_9934);
nand U14614 (N_14614,N_7563,N_9491);
nor U14615 (N_14615,N_9332,N_6699);
nand U14616 (N_14616,N_6236,N_7605);
nor U14617 (N_14617,N_7728,N_7133);
nor U14618 (N_14618,N_6143,N_5979);
nand U14619 (N_14619,N_8368,N_8743);
or U14620 (N_14620,N_8183,N_7507);
or U14621 (N_14621,N_7159,N_7828);
nand U14622 (N_14622,N_6325,N_7590);
nor U14623 (N_14623,N_5876,N_7444);
or U14624 (N_14624,N_5431,N_9346);
or U14625 (N_14625,N_9033,N_5376);
nor U14626 (N_14626,N_6190,N_6841);
or U14627 (N_14627,N_5034,N_7644);
nor U14628 (N_14628,N_8740,N_6492);
and U14629 (N_14629,N_5776,N_9885);
nand U14630 (N_14630,N_7376,N_9827);
and U14631 (N_14631,N_7656,N_7305);
or U14632 (N_14632,N_8125,N_8758);
or U14633 (N_14633,N_6779,N_8540);
nor U14634 (N_14634,N_9828,N_8066);
and U14635 (N_14635,N_7670,N_6437);
nor U14636 (N_14636,N_9702,N_6701);
nor U14637 (N_14637,N_5750,N_6166);
or U14638 (N_14638,N_7595,N_6589);
or U14639 (N_14639,N_9589,N_7247);
nor U14640 (N_14640,N_8474,N_8523);
nor U14641 (N_14641,N_5241,N_8927);
and U14642 (N_14642,N_7461,N_6595);
nand U14643 (N_14643,N_9520,N_9830);
or U14644 (N_14644,N_6948,N_9451);
or U14645 (N_14645,N_8581,N_8996);
nand U14646 (N_14646,N_5609,N_7375);
and U14647 (N_14647,N_9033,N_8566);
nand U14648 (N_14648,N_7993,N_9968);
nor U14649 (N_14649,N_6798,N_7854);
or U14650 (N_14650,N_5787,N_7662);
and U14651 (N_14651,N_6299,N_8725);
and U14652 (N_14652,N_6975,N_8836);
nor U14653 (N_14653,N_9376,N_6443);
nand U14654 (N_14654,N_6904,N_7408);
or U14655 (N_14655,N_8851,N_6215);
and U14656 (N_14656,N_9427,N_5084);
nand U14657 (N_14657,N_9710,N_6982);
and U14658 (N_14658,N_5104,N_5922);
and U14659 (N_14659,N_9011,N_8360);
nand U14660 (N_14660,N_5238,N_6689);
and U14661 (N_14661,N_8115,N_6770);
nand U14662 (N_14662,N_5128,N_8702);
and U14663 (N_14663,N_9550,N_8143);
nand U14664 (N_14664,N_6082,N_6106);
nand U14665 (N_14665,N_7781,N_6184);
or U14666 (N_14666,N_5567,N_8947);
or U14667 (N_14667,N_7310,N_8863);
nor U14668 (N_14668,N_5631,N_5286);
nor U14669 (N_14669,N_5906,N_5686);
nor U14670 (N_14670,N_9397,N_6457);
nor U14671 (N_14671,N_6014,N_9919);
nor U14672 (N_14672,N_5353,N_7421);
and U14673 (N_14673,N_5726,N_5043);
nand U14674 (N_14674,N_8035,N_6376);
nand U14675 (N_14675,N_5045,N_7707);
nor U14676 (N_14676,N_7193,N_7441);
or U14677 (N_14677,N_9326,N_7801);
nor U14678 (N_14678,N_9673,N_8041);
nand U14679 (N_14679,N_9201,N_9890);
nand U14680 (N_14680,N_8146,N_7601);
nor U14681 (N_14681,N_6388,N_9216);
and U14682 (N_14682,N_5038,N_6238);
nor U14683 (N_14683,N_7516,N_6872);
nand U14684 (N_14684,N_7373,N_5907);
nand U14685 (N_14685,N_8120,N_9480);
nand U14686 (N_14686,N_7078,N_8459);
or U14687 (N_14687,N_7316,N_7751);
and U14688 (N_14688,N_7968,N_5941);
nor U14689 (N_14689,N_5726,N_7275);
or U14690 (N_14690,N_6597,N_7767);
nor U14691 (N_14691,N_7290,N_7545);
nand U14692 (N_14692,N_8310,N_9378);
nor U14693 (N_14693,N_5376,N_9786);
nor U14694 (N_14694,N_6248,N_5366);
nand U14695 (N_14695,N_9975,N_7268);
nand U14696 (N_14696,N_6538,N_8233);
xor U14697 (N_14697,N_8472,N_9566);
or U14698 (N_14698,N_6577,N_6658);
and U14699 (N_14699,N_6481,N_6273);
nand U14700 (N_14700,N_8173,N_8163);
nor U14701 (N_14701,N_6741,N_9614);
or U14702 (N_14702,N_6773,N_7739);
nor U14703 (N_14703,N_7667,N_7116);
nand U14704 (N_14704,N_9316,N_6861);
or U14705 (N_14705,N_7345,N_7672);
and U14706 (N_14706,N_7690,N_7099);
or U14707 (N_14707,N_6420,N_8410);
nor U14708 (N_14708,N_6126,N_5599);
nor U14709 (N_14709,N_6951,N_7160);
or U14710 (N_14710,N_5811,N_6281);
and U14711 (N_14711,N_8564,N_8534);
nor U14712 (N_14712,N_9776,N_8749);
and U14713 (N_14713,N_8185,N_5040);
nor U14714 (N_14714,N_8793,N_6042);
nand U14715 (N_14715,N_7175,N_8523);
and U14716 (N_14716,N_6252,N_7366);
nor U14717 (N_14717,N_8324,N_9990);
or U14718 (N_14718,N_5366,N_9713);
nand U14719 (N_14719,N_8791,N_7488);
and U14720 (N_14720,N_7558,N_9860);
nor U14721 (N_14721,N_6068,N_7109);
nand U14722 (N_14722,N_5884,N_5324);
nor U14723 (N_14723,N_9206,N_6726);
nand U14724 (N_14724,N_7334,N_8889);
or U14725 (N_14725,N_7714,N_9074);
or U14726 (N_14726,N_6561,N_5046);
nor U14727 (N_14727,N_6025,N_9163);
or U14728 (N_14728,N_9002,N_6298);
and U14729 (N_14729,N_9466,N_5579);
or U14730 (N_14730,N_5408,N_6111);
nand U14731 (N_14731,N_9011,N_6892);
and U14732 (N_14732,N_8869,N_7697);
nor U14733 (N_14733,N_9456,N_9751);
nor U14734 (N_14734,N_8699,N_6739);
nand U14735 (N_14735,N_6945,N_5628);
or U14736 (N_14736,N_6568,N_7772);
or U14737 (N_14737,N_9289,N_7651);
nand U14738 (N_14738,N_8482,N_8121);
nand U14739 (N_14739,N_7928,N_5536);
nand U14740 (N_14740,N_6631,N_7964);
or U14741 (N_14741,N_5589,N_5333);
nand U14742 (N_14742,N_7808,N_9889);
and U14743 (N_14743,N_5022,N_5674);
and U14744 (N_14744,N_5597,N_5675);
nor U14745 (N_14745,N_8700,N_7716);
nor U14746 (N_14746,N_8765,N_7715);
and U14747 (N_14747,N_8024,N_7612);
or U14748 (N_14748,N_9848,N_5163);
or U14749 (N_14749,N_8127,N_9458);
xnor U14750 (N_14750,N_8931,N_6339);
nor U14751 (N_14751,N_8272,N_6283);
or U14752 (N_14752,N_7668,N_9893);
and U14753 (N_14753,N_9713,N_6323);
xnor U14754 (N_14754,N_5324,N_5521);
and U14755 (N_14755,N_6258,N_9005);
or U14756 (N_14756,N_9074,N_8005);
nor U14757 (N_14757,N_8539,N_6742);
nor U14758 (N_14758,N_7792,N_8078);
and U14759 (N_14759,N_9490,N_9144);
nand U14760 (N_14760,N_9599,N_7167);
and U14761 (N_14761,N_9832,N_9777);
nand U14762 (N_14762,N_8958,N_6395);
nand U14763 (N_14763,N_6429,N_8245);
and U14764 (N_14764,N_5270,N_7033);
nor U14765 (N_14765,N_9703,N_7292);
or U14766 (N_14766,N_6137,N_9556);
and U14767 (N_14767,N_8426,N_6288);
and U14768 (N_14768,N_8807,N_6931);
nand U14769 (N_14769,N_8264,N_5256);
and U14770 (N_14770,N_6452,N_9550);
or U14771 (N_14771,N_5007,N_6709);
nor U14772 (N_14772,N_6019,N_6252);
nand U14773 (N_14773,N_8313,N_7496);
nand U14774 (N_14774,N_7845,N_6184);
or U14775 (N_14775,N_5924,N_5826);
nand U14776 (N_14776,N_7630,N_7555);
nor U14777 (N_14777,N_6336,N_9842);
and U14778 (N_14778,N_9345,N_5666);
nand U14779 (N_14779,N_6535,N_7922);
or U14780 (N_14780,N_9339,N_7282);
nand U14781 (N_14781,N_8664,N_7810);
nor U14782 (N_14782,N_5374,N_7970);
or U14783 (N_14783,N_9279,N_6098);
nand U14784 (N_14784,N_6043,N_8386);
nand U14785 (N_14785,N_8949,N_7999);
and U14786 (N_14786,N_8783,N_6494);
or U14787 (N_14787,N_6639,N_6951);
and U14788 (N_14788,N_7330,N_8037);
nor U14789 (N_14789,N_6155,N_8729);
nand U14790 (N_14790,N_5725,N_6432);
nand U14791 (N_14791,N_9563,N_7840);
nor U14792 (N_14792,N_6167,N_5235);
or U14793 (N_14793,N_8944,N_9696);
or U14794 (N_14794,N_7506,N_8836);
nand U14795 (N_14795,N_8694,N_7324);
or U14796 (N_14796,N_9380,N_6264);
nor U14797 (N_14797,N_6024,N_5314);
or U14798 (N_14798,N_9618,N_7016);
or U14799 (N_14799,N_9699,N_8590);
nand U14800 (N_14800,N_6600,N_7586);
or U14801 (N_14801,N_5139,N_7917);
and U14802 (N_14802,N_5137,N_6296);
or U14803 (N_14803,N_6235,N_8601);
and U14804 (N_14804,N_7395,N_9375);
and U14805 (N_14805,N_9345,N_9515);
nor U14806 (N_14806,N_9048,N_8356);
nor U14807 (N_14807,N_9768,N_6849);
nand U14808 (N_14808,N_8984,N_5937);
nor U14809 (N_14809,N_5391,N_5101);
or U14810 (N_14810,N_7673,N_6394);
and U14811 (N_14811,N_6035,N_6604);
nand U14812 (N_14812,N_6278,N_5058);
nand U14813 (N_14813,N_8873,N_9355);
nor U14814 (N_14814,N_7626,N_8894);
nand U14815 (N_14815,N_8347,N_5870);
or U14816 (N_14816,N_7658,N_7912);
and U14817 (N_14817,N_8225,N_9880);
and U14818 (N_14818,N_7998,N_6792);
and U14819 (N_14819,N_9299,N_7752);
nor U14820 (N_14820,N_7363,N_7285);
nand U14821 (N_14821,N_5841,N_6047);
nand U14822 (N_14822,N_5741,N_8032);
nand U14823 (N_14823,N_7464,N_7959);
nor U14824 (N_14824,N_6060,N_6306);
nor U14825 (N_14825,N_7660,N_7610);
and U14826 (N_14826,N_9441,N_5928);
or U14827 (N_14827,N_8727,N_7889);
nor U14828 (N_14828,N_8941,N_7962);
or U14829 (N_14829,N_5122,N_8166);
and U14830 (N_14830,N_7817,N_6220);
and U14831 (N_14831,N_7690,N_6035);
nor U14832 (N_14832,N_7628,N_5469);
or U14833 (N_14833,N_5294,N_5924);
and U14834 (N_14834,N_8195,N_9434);
and U14835 (N_14835,N_8117,N_9510);
or U14836 (N_14836,N_5482,N_6258);
nor U14837 (N_14837,N_5219,N_7617);
nand U14838 (N_14838,N_5914,N_5155);
or U14839 (N_14839,N_6106,N_5700);
nor U14840 (N_14840,N_8563,N_8371);
and U14841 (N_14841,N_9885,N_7022);
and U14842 (N_14842,N_7767,N_6419);
nor U14843 (N_14843,N_6750,N_8236);
and U14844 (N_14844,N_7727,N_8605);
or U14845 (N_14845,N_5743,N_7057);
nor U14846 (N_14846,N_8630,N_9449);
nor U14847 (N_14847,N_8357,N_7581);
and U14848 (N_14848,N_8710,N_6326);
nand U14849 (N_14849,N_6964,N_6805);
and U14850 (N_14850,N_8680,N_6870);
nand U14851 (N_14851,N_6187,N_5369);
nand U14852 (N_14852,N_9633,N_8237);
nand U14853 (N_14853,N_7674,N_5176);
and U14854 (N_14854,N_8306,N_9407);
nand U14855 (N_14855,N_8220,N_5711);
or U14856 (N_14856,N_8363,N_7680);
nor U14857 (N_14857,N_6820,N_6560);
nand U14858 (N_14858,N_9276,N_5293);
nand U14859 (N_14859,N_5556,N_6210);
nor U14860 (N_14860,N_9660,N_9631);
or U14861 (N_14861,N_8657,N_6830);
or U14862 (N_14862,N_9131,N_5953);
or U14863 (N_14863,N_7231,N_7173);
nand U14864 (N_14864,N_5358,N_8858);
nor U14865 (N_14865,N_6818,N_8693);
or U14866 (N_14866,N_7336,N_8730);
nand U14867 (N_14867,N_7593,N_7776);
nor U14868 (N_14868,N_9162,N_5075);
or U14869 (N_14869,N_5001,N_5632);
and U14870 (N_14870,N_8596,N_5612);
and U14871 (N_14871,N_7946,N_8797);
nor U14872 (N_14872,N_8583,N_8867);
nor U14873 (N_14873,N_7394,N_9735);
nand U14874 (N_14874,N_7990,N_5518);
nor U14875 (N_14875,N_7401,N_9575);
or U14876 (N_14876,N_9587,N_5740);
and U14877 (N_14877,N_9527,N_8420);
nand U14878 (N_14878,N_5115,N_5487);
nor U14879 (N_14879,N_9077,N_6045);
nand U14880 (N_14880,N_5458,N_8425);
or U14881 (N_14881,N_7852,N_6946);
or U14882 (N_14882,N_6423,N_5959);
or U14883 (N_14883,N_8339,N_5922);
nand U14884 (N_14884,N_9421,N_8976);
or U14885 (N_14885,N_8533,N_7678);
and U14886 (N_14886,N_9419,N_9792);
and U14887 (N_14887,N_8841,N_5732);
nor U14888 (N_14888,N_8686,N_6083);
nand U14889 (N_14889,N_6783,N_8459);
nand U14890 (N_14890,N_5704,N_6121);
xor U14891 (N_14891,N_6643,N_5826);
or U14892 (N_14892,N_5862,N_7683);
or U14893 (N_14893,N_5746,N_9177);
nand U14894 (N_14894,N_5950,N_8909);
and U14895 (N_14895,N_6367,N_8482);
and U14896 (N_14896,N_9107,N_8361);
and U14897 (N_14897,N_8950,N_6259);
nand U14898 (N_14898,N_7317,N_5033);
nand U14899 (N_14899,N_6552,N_8657);
nand U14900 (N_14900,N_8250,N_7038);
nand U14901 (N_14901,N_9141,N_5836);
nor U14902 (N_14902,N_8538,N_5538);
nand U14903 (N_14903,N_6191,N_5848);
and U14904 (N_14904,N_9755,N_9811);
or U14905 (N_14905,N_6434,N_9036);
nand U14906 (N_14906,N_6036,N_7282);
or U14907 (N_14907,N_7634,N_7544);
nand U14908 (N_14908,N_8583,N_5434);
or U14909 (N_14909,N_8692,N_8702);
nand U14910 (N_14910,N_7922,N_6219);
and U14911 (N_14911,N_8089,N_6978);
nand U14912 (N_14912,N_7488,N_6661);
and U14913 (N_14913,N_9636,N_6931);
nor U14914 (N_14914,N_6023,N_9150);
or U14915 (N_14915,N_5758,N_9564);
and U14916 (N_14916,N_9377,N_8780);
or U14917 (N_14917,N_9931,N_8995);
nor U14918 (N_14918,N_7325,N_6106);
and U14919 (N_14919,N_9882,N_9008);
and U14920 (N_14920,N_6652,N_9706);
and U14921 (N_14921,N_5924,N_7191);
nand U14922 (N_14922,N_8162,N_7275);
nor U14923 (N_14923,N_6220,N_7837);
nor U14924 (N_14924,N_5403,N_7840);
or U14925 (N_14925,N_7517,N_5450);
nor U14926 (N_14926,N_5599,N_6896);
nand U14927 (N_14927,N_8987,N_9965);
nand U14928 (N_14928,N_5883,N_7239);
nor U14929 (N_14929,N_9821,N_6500);
nand U14930 (N_14930,N_8336,N_6858);
or U14931 (N_14931,N_6696,N_9778);
and U14932 (N_14932,N_9210,N_9901);
or U14933 (N_14933,N_5040,N_5876);
nor U14934 (N_14934,N_5911,N_7773);
xor U14935 (N_14935,N_5062,N_5104);
nand U14936 (N_14936,N_7488,N_9062);
or U14937 (N_14937,N_9880,N_5520);
nor U14938 (N_14938,N_5932,N_8525);
nor U14939 (N_14939,N_9788,N_7531);
or U14940 (N_14940,N_7538,N_9527);
nand U14941 (N_14941,N_5153,N_6139);
nor U14942 (N_14942,N_5329,N_8077);
nand U14943 (N_14943,N_8040,N_5222);
and U14944 (N_14944,N_9035,N_8392);
and U14945 (N_14945,N_9398,N_6709);
or U14946 (N_14946,N_9217,N_9939);
or U14947 (N_14947,N_7420,N_6530);
nor U14948 (N_14948,N_7752,N_5510);
and U14949 (N_14949,N_9731,N_5016);
and U14950 (N_14950,N_9604,N_7892);
or U14951 (N_14951,N_8745,N_9218);
or U14952 (N_14952,N_8058,N_6600);
nand U14953 (N_14953,N_8915,N_7389);
or U14954 (N_14954,N_5100,N_5284);
nand U14955 (N_14955,N_7630,N_9937);
or U14956 (N_14956,N_5638,N_6725);
nor U14957 (N_14957,N_8359,N_7267);
nor U14958 (N_14958,N_8742,N_7749);
and U14959 (N_14959,N_6705,N_5636);
or U14960 (N_14960,N_9627,N_9363);
or U14961 (N_14961,N_6346,N_8330);
nand U14962 (N_14962,N_6269,N_5286);
or U14963 (N_14963,N_6936,N_6543);
nand U14964 (N_14964,N_5652,N_6835);
nor U14965 (N_14965,N_9265,N_5762);
and U14966 (N_14966,N_5314,N_6882);
and U14967 (N_14967,N_5720,N_8533);
and U14968 (N_14968,N_9239,N_7689);
or U14969 (N_14969,N_7000,N_8267);
nand U14970 (N_14970,N_7844,N_8017);
nand U14971 (N_14971,N_9882,N_5495);
or U14972 (N_14972,N_6822,N_8258);
or U14973 (N_14973,N_5236,N_8993);
or U14974 (N_14974,N_7872,N_5875);
nand U14975 (N_14975,N_5825,N_9648);
nand U14976 (N_14976,N_8064,N_6673);
and U14977 (N_14977,N_9456,N_9023);
nor U14978 (N_14978,N_6389,N_5383);
and U14979 (N_14979,N_8343,N_7433);
or U14980 (N_14980,N_9996,N_7683);
or U14981 (N_14981,N_8708,N_9633);
nand U14982 (N_14982,N_5224,N_8891);
and U14983 (N_14983,N_9715,N_5860);
nand U14984 (N_14984,N_5959,N_9224);
and U14985 (N_14985,N_9374,N_9355);
or U14986 (N_14986,N_9924,N_9510);
nor U14987 (N_14987,N_7430,N_5537);
and U14988 (N_14988,N_6280,N_7939);
nor U14989 (N_14989,N_7255,N_7900);
nand U14990 (N_14990,N_9443,N_5405);
nor U14991 (N_14991,N_8389,N_8185);
or U14992 (N_14992,N_5638,N_8973);
or U14993 (N_14993,N_6990,N_9658);
nand U14994 (N_14994,N_9138,N_6174);
nor U14995 (N_14995,N_7472,N_6860);
or U14996 (N_14996,N_6624,N_7769);
xnor U14997 (N_14997,N_6342,N_7233);
nand U14998 (N_14998,N_9125,N_9614);
nor U14999 (N_14999,N_7458,N_6964);
nor U15000 (N_15000,N_11921,N_12466);
and U15001 (N_15001,N_13698,N_14022);
and U15002 (N_15002,N_11286,N_11375);
nor U15003 (N_15003,N_11260,N_12828);
and U15004 (N_15004,N_13091,N_13900);
nand U15005 (N_15005,N_12240,N_12589);
nor U15006 (N_15006,N_13283,N_14618);
and U15007 (N_15007,N_10816,N_14107);
nor U15008 (N_15008,N_10478,N_12030);
nand U15009 (N_15009,N_12621,N_14904);
nand U15010 (N_15010,N_11185,N_10272);
and U15011 (N_15011,N_11846,N_12208);
and U15012 (N_15012,N_10602,N_10205);
and U15013 (N_15013,N_14450,N_11961);
and U15014 (N_15014,N_13986,N_14795);
nor U15015 (N_15015,N_12900,N_14941);
or U15016 (N_15016,N_10723,N_14512);
nor U15017 (N_15017,N_14222,N_12756);
and U15018 (N_15018,N_10435,N_13401);
and U15019 (N_15019,N_11712,N_13046);
and U15020 (N_15020,N_11917,N_12242);
and U15021 (N_15021,N_10082,N_10563);
or U15022 (N_15022,N_12041,N_14766);
nor U15023 (N_15023,N_14288,N_11928);
nand U15024 (N_15024,N_14625,N_10818);
and U15025 (N_15025,N_12063,N_13076);
or U15026 (N_15026,N_14835,N_10288);
nor U15027 (N_15027,N_14575,N_13786);
or U15028 (N_15028,N_14370,N_14111);
or U15029 (N_15029,N_14953,N_12293);
nor U15030 (N_15030,N_13133,N_14465);
or U15031 (N_15031,N_14602,N_13482);
or U15032 (N_15032,N_11896,N_14734);
or U15033 (N_15033,N_14106,N_10040);
and U15034 (N_15034,N_14898,N_10778);
or U15035 (N_15035,N_14113,N_14736);
or U15036 (N_15036,N_12543,N_14627);
nand U15037 (N_15037,N_13866,N_10540);
nand U15038 (N_15038,N_10860,N_12630);
and U15039 (N_15039,N_11445,N_11674);
and U15040 (N_15040,N_10611,N_12893);
or U15041 (N_15041,N_13135,N_11740);
and U15042 (N_15042,N_14387,N_13831);
and U15043 (N_15043,N_10826,N_11782);
or U15044 (N_15044,N_12953,N_12952);
and U15045 (N_15045,N_12949,N_10008);
nor U15046 (N_15046,N_13129,N_14037);
or U15047 (N_15047,N_13600,N_14571);
nand U15048 (N_15048,N_13883,N_13782);
or U15049 (N_15049,N_14368,N_13053);
nand U15050 (N_15050,N_11687,N_10653);
nand U15051 (N_15051,N_10733,N_10779);
nor U15052 (N_15052,N_14403,N_11758);
nand U15053 (N_15053,N_11125,N_11654);
nand U15054 (N_15054,N_13180,N_12812);
and U15055 (N_15055,N_13483,N_13325);
or U15056 (N_15056,N_12838,N_13776);
and U15057 (N_15057,N_13275,N_13265);
nand U15058 (N_15058,N_10041,N_13909);
nand U15059 (N_15059,N_13708,N_12593);
nand U15060 (N_15060,N_13722,N_14710);
nand U15061 (N_15061,N_13902,N_10195);
nor U15062 (N_15062,N_13707,N_11717);
and U15063 (N_15063,N_12750,N_14500);
and U15064 (N_15064,N_10992,N_10843);
nand U15065 (N_15065,N_10949,N_10343);
and U15066 (N_15066,N_11090,N_14066);
nor U15067 (N_15067,N_14744,N_10169);
nand U15068 (N_15068,N_12707,N_10242);
nand U15069 (N_15069,N_10572,N_14347);
or U15070 (N_15070,N_13243,N_10708);
and U15071 (N_15071,N_13004,N_13832);
and U15072 (N_15072,N_11535,N_13457);
or U15073 (N_15073,N_10409,N_14281);
or U15074 (N_15074,N_12633,N_13285);
or U15075 (N_15075,N_14899,N_12637);
nor U15076 (N_15076,N_11910,N_11924);
nor U15077 (N_15077,N_11297,N_12212);
nand U15078 (N_15078,N_12183,N_10077);
nand U15079 (N_15079,N_13274,N_13881);
and U15080 (N_15080,N_13514,N_10419);
or U15081 (N_15081,N_14349,N_11888);
nand U15082 (N_15082,N_11123,N_11413);
nor U15083 (N_15083,N_11056,N_12358);
nand U15084 (N_15084,N_11424,N_14934);
and U15085 (N_15085,N_13822,N_12825);
and U15086 (N_15086,N_11834,N_12808);
nand U15087 (N_15087,N_13979,N_13005);
nor U15088 (N_15088,N_12917,N_12930);
nor U15089 (N_15089,N_12165,N_14345);
nor U15090 (N_15090,N_14320,N_11513);
nand U15091 (N_15091,N_13587,N_13977);
nor U15092 (N_15092,N_12380,N_11680);
nor U15093 (N_15093,N_13565,N_10799);
or U15094 (N_15094,N_12347,N_11761);
nand U15095 (N_15095,N_10166,N_10386);
nor U15096 (N_15096,N_12537,N_12145);
nor U15097 (N_15097,N_11985,N_13888);
and U15098 (N_15098,N_13801,N_13235);
nor U15099 (N_15099,N_13984,N_12426);
nand U15100 (N_15100,N_14930,N_10857);
nor U15101 (N_15101,N_11038,N_13259);
nand U15102 (N_15102,N_14140,N_11007);
nand U15103 (N_15103,N_11823,N_12547);
or U15104 (N_15104,N_13719,N_10274);
and U15105 (N_15105,N_10156,N_10050);
and U15106 (N_15106,N_11875,N_12153);
and U15107 (N_15107,N_12156,N_10861);
nor U15108 (N_15108,N_11841,N_11762);
or U15109 (N_15109,N_12104,N_12186);
nand U15110 (N_15110,N_10675,N_10269);
nand U15111 (N_15111,N_12856,N_14585);
nand U15112 (N_15112,N_13706,N_14606);
and U15113 (N_15113,N_10113,N_12939);
and U15114 (N_15114,N_12877,N_10475);
and U15115 (N_15115,N_11509,N_12790);
or U15116 (N_15116,N_13659,N_10796);
or U15117 (N_15117,N_14142,N_11974);
or U15118 (N_15118,N_13586,N_14435);
or U15119 (N_15119,N_11374,N_10890);
or U15120 (N_15120,N_12540,N_11963);
nand U15121 (N_15121,N_14876,N_13501);
and U15122 (N_15122,N_11996,N_11763);
and U15123 (N_15123,N_13637,N_11912);
and U15124 (N_15124,N_11227,N_13924);
nand U15125 (N_15125,N_11266,N_11950);
or U15126 (N_15126,N_14259,N_14467);
and U15127 (N_15127,N_14544,N_11043);
nor U15128 (N_15128,N_10640,N_12205);
and U15129 (N_15129,N_12309,N_12913);
nor U15130 (N_15130,N_14681,N_11771);
nand U15131 (N_15131,N_13442,N_13226);
or U15132 (N_15132,N_12399,N_14346);
and U15133 (N_15133,N_11534,N_14531);
nor U15134 (N_15134,N_12978,N_11252);
nor U15135 (N_15135,N_11991,N_10736);
and U15136 (N_15136,N_11719,N_10815);
or U15137 (N_15137,N_12495,N_11517);
nand U15138 (N_15138,N_12308,N_14129);
nor U15139 (N_15139,N_12510,N_10732);
or U15140 (N_15140,N_14502,N_13804);
or U15141 (N_15141,N_10183,N_14595);
and U15142 (N_15142,N_13910,N_10445);
xor U15143 (N_15143,N_14741,N_12757);
or U15144 (N_15144,N_13111,N_14237);
nand U15145 (N_15145,N_12775,N_10026);
and U15146 (N_15146,N_14514,N_10937);
nand U15147 (N_15147,N_11546,N_12470);
xor U15148 (N_15148,N_13648,N_11222);
and U15149 (N_15149,N_14203,N_11666);
nand U15150 (N_15150,N_12502,N_14511);
and U15151 (N_15151,N_10748,N_13069);
or U15152 (N_15152,N_12754,N_10609);
nand U15153 (N_15153,N_10509,N_10657);
nor U15154 (N_15154,N_12420,N_10803);
nand U15155 (N_15155,N_10024,N_12749);
nand U15156 (N_15156,N_12962,N_11840);
or U15157 (N_15157,N_11436,N_13421);
and U15158 (N_15158,N_13360,N_12159);
xnor U15159 (N_15159,N_12627,N_10381);
nand U15160 (N_15160,N_10241,N_11965);
and U15161 (N_15161,N_13165,N_12146);
and U15162 (N_15162,N_14838,N_14060);
nor U15163 (N_15163,N_14378,N_14718);
nor U15164 (N_15164,N_12103,N_11756);
or U15165 (N_15165,N_12769,N_12517);
nor U15166 (N_15166,N_14683,N_11272);
nor U15167 (N_15167,N_13519,N_14960);
nor U15168 (N_15168,N_11933,N_12742);
nor U15169 (N_15169,N_12954,N_11549);
or U15170 (N_15170,N_14938,N_13836);
and U15171 (N_15171,N_10498,N_13830);
or U15172 (N_15172,N_12849,N_12360);
and U15173 (N_15173,N_13149,N_14495);
nand U15174 (N_15174,N_14994,N_12709);
or U15175 (N_15175,N_12227,N_14810);
and U15176 (N_15176,N_13625,N_10063);
nor U15177 (N_15177,N_11315,N_10384);
and U15178 (N_15178,N_13879,N_12260);
nor U15179 (N_15179,N_12112,N_11214);
nor U15180 (N_15180,N_13552,N_14555);
nand U15181 (N_15181,N_13415,N_10821);
and U15182 (N_15182,N_10016,N_13153);
or U15183 (N_15183,N_10883,N_11516);
nor U15184 (N_15184,N_10994,N_12759);
nor U15185 (N_15185,N_12291,N_11200);
or U15186 (N_15186,N_11156,N_13969);
and U15187 (N_15187,N_14025,N_12128);
nor U15188 (N_15188,N_12278,N_14947);
nand U15189 (N_15189,N_11064,N_14784);
nand U15190 (N_15190,N_11778,N_12752);
and U15191 (N_15191,N_10112,N_10713);
nand U15192 (N_15192,N_11023,N_13861);
nor U15193 (N_15193,N_12125,N_11229);
or U15194 (N_15194,N_13343,N_12698);
nor U15195 (N_15195,N_11789,N_10940);
and U15196 (N_15196,N_12343,N_14139);
or U15197 (N_15197,N_11372,N_10226);
nand U15198 (N_15198,N_11481,N_11028);
or U15199 (N_15199,N_14217,N_14959);
nor U15200 (N_15200,N_14956,N_14305);
xnor U15201 (N_15201,N_14837,N_10373);
nand U15202 (N_15202,N_13263,N_10812);
nor U15203 (N_15203,N_11948,N_13895);
nor U15204 (N_15204,N_12014,N_10967);
or U15205 (N_15205,N_12109,N_14707);
nand U15206 (N_15206,N_14522,N_11897);
and U15207 (N_15207,N_12081,N_10094);
or U15208 (N_15208,N_14038,N_13264);
nand U15209 (N_15209,N_12765,N_13916);
or U15210 (N_15210,N_12615,N_11166);
or U15211 (N_15211,N_14570,N_14358);
nor U15212 (N_15212,N_13915,N_14191);
nor U15213 (N_15213,N_14123,N_11442);
nor U15214 (N_15214,N_11766,N_10551);
nor U15215 (N_15215,N_14887,N_10366);
and U15216 (N_15216,N_13276,N_11721);
nor U15217 (N_15217,N_11063,N_13777);
nor U15218 (N_15218,N_13917,N_11514);
and U15219 (N_15219,N_11569,N_14819);
nand U15220 (N_15220,N_11865,N_13997);
nor U15221 (N_15221,N_12976,N_10402);
nor U15222 (N_15222,N_10989,N_11678);
or U15223 (N_15223,N_13225,N_10938);
and U15224 (N_15224,N_13674,N_12704);
nand U15225 (N_15225,N_11695,N_11464);
and U15226 (N_15226,N_14829,N_11004);
and U15227 (N_15227,N_14210,N_11280);
and U15228 (N_15228,N_10814,N_11640);
or U15229 (N_15229,N_12028,N_13035);
nor U15230 (N_15230,N_10827,N_13184);
or U15231 (N_15231,N_14893,N_13377);
nor U15232 (N_15232,N_13738,N_11314);
and U15233 (N_15233,N_14176,N_13368);
and U15234 (N_15234,N_11988,N_13268);
nand U15235 (N_15235,N_13006,N_10762);
nand U15236 (N_15236,N_11303,N_10404);
nor U15237 (N_15237,N_12942,N_14411);
or U15238 (N_15238,N_14015,N_14613);
and U15239 (N_15239,N_14189,N_10273);
nor U15240 (N_15240,N_12780,N_11368);
or U15241 (N_15241,N_14473,N_12904);
and U15242 (N_15242,N_11002,N_14270);
nor U15243 (N_15243,N_11136,N_14386);
nand U15244 (N_15244,N_14763,N_11418);
and U15245 (N_15245,N_12440,N_11845);
or U15246 (N_15246,N_12029,N_10870);
nand U15247 (N_15247,N_13124,N_11816);
nand U15248 (N_15248,N_13667,N_12070);
or U15249 (N_15249,N_13538,N_14033);
or U15250 (N_15250,N_12150,N_13658);
xnor U15251 (N_15251,N_10214,N_13548);
nor U15252 (N_15252,N_12268,N_10131);
nand U15253 (N_15253,N_11079,N_14916);
nor U15254 (N_15254,N_10872,N_12501);
and U15255 (N_15255,N_14642,N_13468);
and U15256 (N_15256,N_12441,N_13178);
nand U15257 (N_15257,N_10283,N_14536);
nand U15258 (N_15258,N_14634,N_12503);
and U15259 (N_15259,N_12496,N_10412);
nor U15260 (N_15260,N_13663,N_13399);
and U15261 (N_15261,N_12386,N_13778);
or U15262 (N_15262,N_10891,N_14289);
or U15263 (N_15263,N_13281,N_10901);
nand U15264 (N_15264,N_12715,N_12901);
or U15265 (N_15265,N_10904,N_11600);
and U15266 (N_15266,N_14223,N_11207);
nand U15267 (N_15267,N_11751,N_12580);
and U15268 (N_15268,N_10126,N_12875);
xor U15269 (N_15269,N_13718,N_14126);
and U15270 (N_15270,N_12694,N_12654);
and U15271 (N_15271,N_12179,N_11025);
nor U15272 (N_15272,N_12985,N_12349);
nand U15273 (N_15273,N_12894,N_14943);
nor U15274 (N_15274,N_11074,N_13388);
or U15275 (N_15275,N_13595,N_14405);
nor U15276 (N_15276,N_14484,N_14909);
nor U15277 (N_15277,N_12974,N_11582);
or U15278 (N_15278,N_10852,N_13349);
or U15279 (N_15279,N_10962,N_12273);
nor U15280 (N_15280,N_11860,N_11001);
nand U15281 (N_15281,N_13452,N_12193);
nand U15282 (N_15282,N_12243,N_14709);
nor U15283 (N_15283,N_13928,N_14933);
nor U15284 (N_15284,N_14644,N_10232);
nor U15285 (N_15285,N_14727,N_13607);
or U15286 (N_15286,N_10911,N_14521);
and U15287 (N_15287,N_11389,N_12906);
nand U15288 (N_15288,N_14871,N_13002);
nand U15289 (N_15289,N_14961,N_13673);
and U15290 (N_15290,N_14005,N_11645);
or U15291 (N_15291,N_11706,N_14043);
and U15292 (N_15292,N_13988,N_13704);
or U15293 (N_15293,N_12181,N_10106);
nand U15294 (N_15294,N_14751,N_13267);
or U15295 (N_15295,N_10141,N_12903);
and U15296 (N_15296,N_13952,N_13375);
nor U15297 (N_15297,N_10934,N_13992);
or U15298 (N_15298,N_11512,N_14458);
or U15299 (N_15299,N_13875,N_10281);
nor U15300 (N_15300,N_10154,N_12883);
nand U15301 (N_15301,N_10292,N_11739);
or U15302 (N_15302,N_12272,N_13340);
or U15303 (N_15303,N_13374,N_11365);
nor U15304 (N_15304,N_12591,N_11699);
and U15305 (N_15305,N_13887,N_12523);
or U15306 (N_15306,N_12254,N_13182);
nand U15307 (N_15307,N_14132,N_12073);
or U15308 (N_15308,N_10933,N_14291);
or U15309 (N_15309,N_13838,N_10715);
nor U15310 (N_15310,N_12132,N_14851);
and U15311 (N_15311,N_13662,N_10033);
nand U15312 (N_15312,N_13039,N_13392);
nand U15313 (N_15313,N_11279,N_13232);
nor U15314 (N_15314,N_11657,N_12782);
nand U15315 (N_15315,N_10158,N_13271);
nand U15316 (N_15316,N_13258,N_14050);
and U15317 (N_15317,N_14350,N_11998);
nor U15318 (N_15318,N_14753,N_13333);
or U15319 (N_15319,N_10757,N_14483);
nor U15320 (N_15320,N_12133,N_12803);
or U15321 (N_15321,N_12472,N_14457);
or U15322 (N_15322,N_11526,N_10727);
nand U15323 (N_15323,N_10314,N_12642);
nor U15324 (N_15324,N_14410,N_14393);
and U15325 (N_15325,N_11573,N_13899);
or U15326 (N_15326,N_10278,N_14341);
or U15327 (N_15327,N_11482,N_13371);
nand U15328 (N_15328,N_10341,N_10134);
nand U15329 (N_15329,N_13459,N_13562);
nand U15330 (N_15330,N_10544,N_13622);
nand U15331 (N_15331,N_12732,N_14992);
nand U15332 (N_15332,N_13498,N_11217);
nor U15333 (N_15333,N_14556,N_13545);
and U15334 (N_15334,N_14508,N_12527);
or U15335 (N_15335,N_12880,N_14926);
nand U15336 (N_15336,N_14286,N_13451);
or U15337 (N_15337,N_10262,N_13199);
nand U15338 (N_15338,N_10930,N_14371);
or U15339 (N_15339,N_14218,N_13985);
nor U15340 (N_15340,N_11926,N_11343);
xnor U15341 (N_15341,N_11632,N_11670);
nand U15342 (N_15342,N_11171,N_11127);
and U15343 (N_15343,N_11115,N_12407);
or U15344 (N_15344,N_11119,N_11357);
and U15345 (N_15345,N_11664,N_12442);
or U15346 (N_15346,N_11525,N_10577);
nand U15347 (N_15347,N_12197,N_13508);
or U15348 (N_15348,N_12361,N_14152);
and U15349 (N_15349,N_10078,N_10036);
nand U15350 (N_15350,N_10575,N_14392);
nor U15351 (N_15351,N_14799,N_12219);
and U15352 (N_15352,N_11018,N_10880);
and U15353 (N_15353,N_10634,N_14955);
or U15354 (N_15354,N_10737,N_11745);
nor U15355 (N_15355,N_11275,N_14175);
nand U15356 (N_15356,N_13387,N_11929);
and U15357 (N_15357,N_12173,N_14932);
and U15358 (N_15358,N_12912,N_11407);
and U15359 (N_15359,N_11385,N_14180);
nor U15360 (N_15360,N_14099,N_13958);
nand U15361 (N_15361,N_11801,N_10403);
or U15362 (N_15362,N_13774,N_12310);
nor U15363 (N_15363,N_10344,N_14630);
or U15364 (N_15364,N_13589,N_10615);
nor U15365 (N_15365,N_11285,N_14576);
and U15366 (N_15366,N_13594,N_12480);
and U15367 (N_15367,N_11749,N_11396);
nand U15368 (N_15368,N_12872,N_12712);
and U15369 (N_15369,N_10886,N_13829);
nor U15370 (N_15370,N_10758,N_13533);
nor U15371 (N_15371,N_10467,N_14390);
nand U15372 (N_15372,N_12252,N_12682);
or U15373 (N_15373,N_14888,N_13125);
or U15374 (N_15374,N_13300,N_13351);
nor U15375 (N_15375,N_11259,N_13769);
nand U15376 (N_15376,N_13834,N_14779);
nand U15377 (N_15377,N_13029,N_13438);
nand U15378 (N_15378,N_11711,N_14702);
and U15379 (N_15379,N_12220,N_13982);
nor U15380 (N_15380,N_13554,N_14389);
or U15381 (N_15381,N_13183,N_13148);
and U15382 (N_15382,N_11530,N_14588);
nand U15383 (N_15383,N_11468,N_11827);
or U15384 (N_15384,N_10393,N_11052);
nand U15385 (N_15385,N_12071,N_12788);
or U15386 (N_15386,N_13689,N_12600);
nand U15387 (N_15387,N_13932,N_13746);
nand U15388 (N_15388,N_11510,N_13294);
nor U15389 (N_15389,N_14265,N_11918);
nor U15390 (N_15390,N_10510,N_11121);
nand U15391 (N_15391,N_10355,N_12973);
nand U15392 (N_15392,N_12218,N_11324);
or U15393 (N_15393,N_13756,N_14115);
or U15394 (N_15394,N_11548,N_13079);
nand U15395 (N_15395,N_10869,N_13494);
nand U15396 (N_15396,N_14342,N_10309);
or U15397 (N_15397,N_10461,N_10349);
or U15398 (N_15398,N_11784,N_11972);
and U15399 (N_15399,N_12533,N_13121);
or U15400 (N_15400,N_11946,N_13332);
nor U15401 (N_15401,N_13592,N_14914);
or U15402 (N_15402,N_13207,N_10623);
nand U15403 (N_15403,N_10415,N_12332);
or U15404 (N_15404,N_11172,N_12889);
or U15405 (N_15405,N_14680,N_14839);
nor U15406 (N_15406,N_11159,N_10781);
or U15407 (N_15407,N_13669,N_13423);
nand U15408 (N_15408,N_12324,N_13015);
nor U15409 (N_15409,N_12024,N_13266);
or U15410 (N_15410,N_14031,N_10382);
nand U15411 (N_15411,N_10842,N_11820);
nor U15412 (N_15412,N_11300,N_11165);
xnor U15413 (N_15413,N_10444,N_13356);
or U15414 (N_15414,N_10661,N_13302);
and U15415 (N_15415,N_13870,N_11147);
nor U15416 (N_15416,N_10110,N_10836);
and U15417 (N_15417,N_10570,N_14832);
and U15418 (N_15418,N_11192,N_13461);
nand U15419 (N_15419,N_10523,N_14145);
nand U15420 (N_15420,N_13602,N_10353);
and U15421 (N_15421,N_12649,N_10754);
nand U15422 (N_15422,N_14742,N_14296);
or U15423 (N_15423,N_10636,N_10589);
or U15424 (N_15424,N_14809,N_12123);
nand U15425 (N_15425,N_10954,N_12982);
and U15426 (N_15426,N_12055,N_14052);
nand U15427 (N_15427,N_14474,N_11561);
nor U15428 (N_15428,N_13237,N_14657);
or U15429 (N_15429,N_10390,N_14211);
or U15430 (N_15430,N_13931,N_11892);
nor U15431 (N_15431,N_12626,N_14748);
or U15432 (N_15432,N_14164,N_11175);
or U15433 (N_15433,N_14523,N_11455);
and U15434 (N_15434,N_10742,N_14737);
nand U15435 (N_15435,N_13835,N_12101);
nor U15436 (N_15436,N_12816,N_12972);
and U15437 (N_15437,N_12222,N_13536);
nand U15438 (N_15438,N_10271,N_10053);
nor U15439 (N_15439,N_10357,N_10706);
or U15440 (N_15440,N_10248,N_12546);
or U15441 (N_15441,N_12459,N_13289);
or U15442 (N_15442,N_11915,N_10721);
or U15443 (N_15443,N_14660,N_11096);
nand U15444 (N_15444,N_14794,N_12172);
and U15445 (N_15445,N_10287,N_14905);
nor U15446 (N_15446,N_12512,N_11939);
nor U15447 (N_15447,N_13167,N_11454);
and U15448 (N_15448,N_12054,N_10527);
xnor U15449 (N_15449,N_12735,N_13677);
or U15450 (N_15450,N_10442,N_14714);
or U15451 (N_15451,N_12049,N_10590);
nand U15452 (N_15452,N_10389,N_12666);
and U15453 (N_15453,N_14398,N_10520);
or U15454 (N_15454,N_11738,N_11938);
and U15455 (N_15455,N_12673,N_10494);
nor U15456 (N_15456,N_12261,N_12207);
nor U15457 (N_15457,N_14421,N_10607);
or U15458 (N_15458,N_12943,N_12933);
or U15459 (N_15459,N_10437,N_13551);
and U15460 (N_15460,N_10569,N_11731);
or U15461 (N_15461,N_12991,N_12538);
nor U15462 (N_15462,N_10299,N_10541);
nor U15463 (N_15463,N_13036,N_11497);
xor U15464 (N_15464,N_13209,N_10761);
nand U15465 (N_15465,N_10454,N_10969);
nand U15466 (N_15466,N_11358,N_14747);
or U15467 (N_15467,N_14783,N_10327);
and U15468 (N_15468,N_14407,N_14501);
nand U15469 (N_15469,N_12603,N_14250);
and U15470 (N_15470,N_12967,N_13695);
and U15471 (N_15471,N_12795,N_14815);
and U15472 (N_15472,N_11021,N_14105);
and U15473 (N_15473,N_14979,N_14706);
or U15474 (N_15474,N_14833,N_13112);
nand U15475 (N_15475,N_14638,N_11579);
and U15476 (N_15476,N_13028,N_11869);
and U15477 (N_15477,N_13903,N_13889);
and U15478 (N_15478,N_14920,N_14340);
nand U15479 (N_15479,N_12623,N_10682);
xnor U15480 (N_15480,N_11142,N_14593);
or U15481 (N_15481,N_11451,N_13848);
nand U15482 (N_15482,N_14429,N_13606);
and U15483 (N_15483,N_13130,N_13311);
and U15484 (N_15484,N_13873,N_11710);
nor U15485 (N_15485,N_10542,N_14449);
nand U15486 (N_15486,N_13190,N_13480);
or U15487 (N_15487,N_14771,N_10557);
or U15488 (N_15488,N_10217,N_12570);
nor U15489 (N_15489,N_14789,N_14154);
xnor U15490 (N_15490,N_14054,N_11319);
and U15491 (N_15491,N_13676,N_10695);
and U15492 (N_15492,N_12339,N_11764);
nor U15493 (N_15493,N_14061,N_10958);
nor U15494 (N_15494,N_13713,N_11646);
nand U15495 (N_15495,N_11157,N_12114);
and U15496 (N_15496,N_14738,N_13413);
nand U15497 (N_15497,N_10545,N_10512);
and U15498 (N_15498,N_11086,N_13488);
or U15499 (N_15499,N_14122,N_13393);
nor U15500 (N_15500,N_14455,N_12850);
or U15501 (N_15501,N_10772,N_11466);
or U15502 (N_15502,N_12705,N_12006);
and U15503 (N_15503,N_12667,N_11610);
and U15504 (N_15504,N_14664,N_11124);
and U15505 (N_15505,N_13974,N_13813);
nand U15506 (N_15506,N_13110,N_13327);
and U15507 (N_15507,N_14408,N_12595);
nor U15508 (N_15508,N_11291,N_12005);
or U15509 (N_15509,N_13402,N_11073);
and U15510 (N_15510,N_12628,N_10745);
and U15511 (N_15511,N_14042,N_13994);
nand U15512 (N_15512,N_14791,N_13161);
or U15513 (N_15513,N_10800,N_13995);
nand U15514 (N_15514,N_11715,N_10650);
nand U15515 (N_15515,N_13664,N_12734);
or U15516 (N_15516,N_14055,N_10418);
or U15517 (N_15517,N_13138,N_11603);
nand U15518 (N_15518,N_10229,N_10369);
or U15519 (N_15519,N_13410,N_14759);
nand U15520 (N_15520,N_13042,N_14667);
nor U15521 (N_15521,N_10658,N_11379);
or U15522 (N_15522,N_11053,N_14353);
and U15523 (N_15523,N_12988,N_12706);
and U15524 (N_15524,N_12955,N_11070);
or U15525 (N_15525,N_11274,N_10767);
and U15526 (N_15526,N_14552,N_13050);
nand U15527 (N_15527,N_13038,N_10674);
or U15528 (N_15528,N_14619,N_12562);
or U15529 (N_15529,N_11893,N_13196);
or U15530 (N_15530,N_14177,N_13559);
or U15531 (N_15531,N_11164,N_12490);
nand U15532 (N_15532,N_13789,N_10775);
nor U15533 (N_15533,N_13828,N_11293);
xor U15534 (N_15534,N_12017,N_13636);
or U15535 (N_15535,N_10250,N_14277);
nor U15536 (N_15536,N_11168,N_14978);
nand U15537 (N_15537,N_11443,N_13239);
nand U15538 (N_15538,N_11339,N_13730);
nand U15539 (N_15539,N_13605,N_12120);
or U15540 (N_15540,N_10491,N_11855);
and U15541 (N_15541,N_11467,N_12866);
and U15542 (N_15542,N_11634,N_10651);
and U15543 (N_15543,N_12516,N_12200);
nor U15544 (N_15544,N_14873,N_11110);
nand U15545 (N_15545,N_10124,N_11877);
nor U15546 (N_15546,N_13071,N_10605);
nand U15547 (N_15547,N_12577,N_10019);
nand U15548 (N_15548,N_12393,N_10452);
nand U15549 (N_15549,N_11256,N_10211);
nor U15550 (N_15550,N_13181,N_14146);
and U15551 (N_15551,N_12660,N_11474);
or U15552 (N_15552,N_10447,N_11619);
and U15553 (N_15553,N_13792,N_12052);
nand U15554 (N_15554,N_14257,N_10638);
or U15555 (N_15555,N_13502,N_11889);
or U15556 (N_15556,N_14973,N_13741);
or U15557 (N_15557,N_12842,N_14194);
nor U15558 (N_15558,N_12373,N_11984);
or U15559 (N_15559,N_11470,N_14863);
nand U15560 (N_15560,N_13198,N_11230);
and U15561 (N_15561,N_10871,N_11606);
and U15562 (N_15562,N_10300,N_12053);
xor U15563 (N_15563,N_14862,N_12082);
or U15564 (N_15564,N_14225,N_12390);
and U15565 (N_15565,N_12369,N_13395);
and U15566 (N_15566,N_10873,N_10506);
and U15567 (N_15567,N_11105,N_12202);
nor U15568 (N_15568,N_11898,N_10251);
nor U15569 (N_15569,N_13642,N_10522);
or U15570 (N_15570,N_13416,N_12829);
nand U15571 (N_15571,N_12773,N_12266);
nand U15572 (N_15572,N_12995,N_12381);
nand U15573 (N_15573,N_12095,N_12733);
nand U15574 (N_15574,N_12851,N_10279);
or U15575 (N_15575,N_10079,N_13493);
or U15576 (N_15576,N_11832,N_13440);
xnor U15577 (N_15577,N_14968,N_10606);
and U15578 (N_15578,N_12141,N_10738);
nand U15579 (N_15579,N_13630,N_12198);
nor U15580 (N_15580,N_12986,N_10173);
and U15581 (N_15581,N_11085,N_10218);
xor U15582 (N_15582,N_12237,N_10788);
and U15583 (N_15583,N_11099,N_14083);
and U15584 (N_15584,N_11432,N_13847);
xnor U15585 (N_15585,N_10237,N_11189);
or U15586 (N_15586,N_14462,N_11033);
nor U15587 (N_15587,N_10068,N_14275);
or U15588 (N_15588,N_13603,N_10099);
nand U15589 (N_15589,N_10848,N_11042);
nor U15590 (N_15590,N_10986,N_14755);
nand U15591 (N_15591,N_10717,N_13011);
or U15592 (N_15592,N_10867,N_13874);
and U15593 (N_15593,N_10030,N_12225);
nor U15594 (N_15594,N_10247,N_11927);
and U15595 (N_15595,N_10428,N_14509);
and U15596 (N_15596,N_13060,N_12508);
and U15597 (N_15597,N_13965,N_13597);
xnor U15598 (N_15598,N_14253,N_11387);
nand U15599 (N_15599,N_13967,N_12271);
nor U15600 (N_15600,N_11973,N_11197);
or U15601 (N_15601,N_11744,N_12344);
nor U15602 (N_15602,N_14962,N_13099);
nor U15603 (N_15603,N_10604,N_13208);
nand U15604 (N_15604,N_12463,N_14285);
or U15605 (N_15605,N_10220,N_11296);
and U15606 (N_15606,N_13615,N_14775);
or U15607 (N_15607,N_14482,N_10175);
nand U15608 (N_15608,N_10120,N_12462);
or U15609 (N_15609,N_11703,N_13886);
and U15610 (N_15610,N_12807,N_13734);
or U15611 (N_15611,N_12044,N_11696);
nor U15612 (N_15612,N_14732,N_11377);
or U15613 (N_15613,N_14604,N_12236);
nand U15614 (N_15614,N_11457,N_14461);
or U15615 (N_15615,N_14633,N_11819);
nor U15616 (N_15616,N_14214,N_14656);
nor U15617 (N_15617,N_12563,N_14293);
nand U15618 (N_15618,N_14685,N_12837);
or U15619 (N_15619,N_11627,N_10177);
nand U15620 (N_15620,N_11618,N_13938);
nor U15621 (N_15621,N_12238,N_14437);
or U15622 (N_15622,N_12922,N_11876);
nand U15623 (N_15623,N_12003,N_13305);
or U15624 (N_15624,N_11523,N_10324);
nor U15625 (N_15625,N_14963,N_14911);
nor U15626 (N_15626,N_11777,N_11810);
nor U15627 (N_15627,N_14244,N_12191);
or U15628 (N_15628,N_14078,N_13684);
or U15629 (N_15629,N_11900,N_12571);
and U15630 (N_15630,N_12650,N_11013);
or U15631 (N_15631,N_11848,N_12576);
nor U15632 (N_15632,N_10993,N_11490);
nor U15633 (N_15633,N_11630,N_14767);
nor U15634 (N_15634,N_11944,N_11177);
or U15635 (N_15635,N_11748,N_12194);
and U15636 (N_15636,N_11886,N_11909);
nand U15637 (N_15637,N_11773,N_11511);
or U15638 (N_15638,N_10664,N_11397);
or U15639 (N_15639,N_14002,N_14489);
or U15640 (N_15640,N_14205,N_14640);
and U15641 (N_15641,N_13222,N_12387);
and U15642 (N_15642,N_10942,N_14252);
nor U15643 (N_15643,N_14772,N_10996);
nand U15644 (N_15644,N_12249,N_13693);
or U15645 (N_15645,N_12318,N_13223);
or U15646 (N_15646,N_10011,N_10647);
nand U15647 (N_15647,N_11458,N_10104);
nor U15648 (N_15648,N_13282,N_10002);
and U15649 (N_15649,N_11193,N_10420);
or U15650 (N_15650,N_14527,N_14884);
and U15651 (N_15651,N_14670,N_14266);
and U15652 (N_15652,N_12451,N_13162);
and U15653 (N_15653,N_10219,N_14469);
nand U15654 (N_15654,N_11383,N_14331);
nor U15655 (N_15655,N_12468,N_13582);
and U15656 (N_15656,N_12348,N_13211);
and U15657 (N_15657,N_11936,N_10552);
or U15658 (N_15658,N_14750,N_10155);
and U15659 (N_15659,N_13398,N_13323);
or U15660 (N_15660,N_11048,N_10817);
and U15661 (N_15661,N_10770,N_11791);
and U15662 (N_15662,N_12535,N_14196);
nor U15663 (N_15663,N_10466,N_11287);
nand U15664 (N_15664,N_11224,N_11465);
nor U15665 (N_15665,N_10319,N_14517);
and U15666 (N_15666,N_12004,N_14404);
or U15667 (N_15667,N_11066,N_12713);
nor U15668 (N_15668,N_11952,N_13299);
nor U15669 (N_15669,N_13082,N_14843);
or U15670 (N_15670,N_13897,N_14985);
nor U15671 (N_15671,N_11725,N_12859);
nand U15672 (N_15672,N_11806,N_12007);
nor U15673 (N_15673,N_13935,N_12811);
nand U15674 (N_15674,N_13660,N_11679);
nand U15675 (N_15675,N_14024,N_11329);
nand U15676 (N_15676,N_12087,N_13681);
and U15677 (N_15677,N_12211,N_13064);
and U15678 (N_15678,N_11187,N_14616);
and U15679 (N_15679,N_10691,N_14650);
nor U15680 (N_15680,N_12277,N_14261);
and U15681 (N_15681,N_13960,N_14768);
nor U15682 (N_15682,N_12443,N_13301);
or U15683 (N_15683,N_12931,N_12886);
nand U15684 (N_15684,N_10123,N_12121);
nand U15685 (N_15685,N_12264,N_13627);
nor U15686 (N_15686,N_11447,N_13250);
or U15687 (N_15687,N_14415,N_11624);
or U15688 (N_15688,N_14859,N_12089);
and U15689 (N_15689,N_13815,N_14141);
nor U15690 (N_15690,N_12918,N_13728);
nand U15691 (N_15691,N_12902,N_14974);
and U15692 (N_15692,N_10303,N_12263);
nor U15693 (N_15693,N_13943,N_14151);
and U15694 (N_15694,N_14114,N_12558);
or U15695 (N_15695,N_13114,N_11577);
and U15696 (N_15696,N_11084,N_14589);
and U15697 (N_15697,N_13269,N_14677);
or U15698 (N_15698,N_12356,N_13429);
or U15699 (N_15699,N_11498,N_14069);
nand U15700 (N_15700,N_13346,N_10618);
or U15701 (N_15701,N_12336,N_13077);
nor U15702 (N_15702,N_13455,N_11599);
nor U15703 (N_15703,N_12355,N_14841);
xor U15704 (N_15704,N_12341,N_11206);
nor U15705 (N_15705,N_12970,N_10593);
and U15706 (N_15706,N_12086,N_11010);
nand U15707 (N_15707,N_12406,N_13764);
nor U15708 (N_15708,N_13688,N_14023);
or U15709 (N_15709,N_10153,N_10525);
nor U15710 (N_15710,N_13370,N_14749);
nor U15711 (N_15711,N_12365,N_13260);
and U15712 (N_15712,N_12979,N_10162);
or U15713 (N_15713,N_11149,N_14695);
or U15714 (N_15714,N_14188,N_12556);
and U15715 (N_15715,N_11796,N_12739);
nand U15716 (N_15716,N_14027,N_14842);
nor U15717 (N_15717,N_12680,N_12408);
and U15718 (N_15718,N_14858,N_10685);
or U15719 (N_15719,N_11659,N_12478);
and U15720 (N_15720,N_13795,N_10896);
nor U15721 (N_15721,N_10686,N_10773);
or U15722 (N_15722,N_10567,N_12761);
nand U15723 (N_15723,N_13680,N_11661);
nor U15724 (N_15724,N_13939,N_10286);
xnor U15725 (N_15725,N_14162,N_12098);
nor U15726 (N_15726,N_11461,N_13843);
and U15727 (N_15727,N_13896,N_14922);
nor U15728 (N_15728,N_13231,N_12090);
or U15729 (N_15729,N_10795,N_12575);
nand U15730 (N_15730,N_12199,N_13107);
or U15731 (N_15731,N_11393,N_14519);
nor U15732 (N_15732,N_11245,N_14659);
and U15733 (N_15733,N_10297,N_12963);
and U15734 (N_15734,N_10206,N_14688);
nor U15735 (N_15735,N_14335,N_13251);
and U15736 (N_15736,N_11993,N_14073);
nand U15737 (N_15737,N_11281,N_14605);
nor U15738 (N_15738,N_11433,N_10953);
or U15739 (N_15739,N_11566,N_11960);
nor U15740 (N_15740,N_13692,N_14471);
or U15741 (N_15741,N_10550,N_12932);
or U15742 (N_15742,N_10808,N_12945);
and U15743 (N_15743,N_11062,N_11551);
nand U15744 (N_15744,N_10961,N_10760);
nor U15745 (N_15745,N_10932,N_11268);
and U15746 (N_15746,N_10365,N_10021);
or U15747 (N_15747,N_13650,N_10417);
and U15748 (N_15748,N_12681,N_12882);
nor U15749 (N_15749,N_11024,N_10917);
and U15750 (N_15750,N_12460,N_13414);
nand U15751 (N_15751,N_11203,N_13543);
nand U15752 (N_15752,N_11653,N_14464);
nand U15753 (N_15753,N_10627,N_13770);
nand U15754 (N_15754,N_14103,N_11570);
nand U15755 (N_15755,N_14216,N_13812);
nor U15756 (N_15756,N_13462,N_13626);
nor U15757 (N_15757,N_14937,N_13557);
and U15758 (N_15758,N_10581,N_13160);
nor U15759 (N_15759,N_11437,N_10925);
or U15760 (N_15760,N_13316,N_11223);
and U15761 (N_15761,N_14121,N_10321);
nand U15762 (N_15762,N_11765,N_10599);
or U15763 (N_15763,N_10087,N_13661);
and U15764 (N_15764,N_13027,N_11003);
or U15765 (N_15765,N_10908,N_11883);
xnor U15766 (N_15766,N_10802,N_11029);
nand U15767 (N_15767,N_14491,N_11908);
nand U15768 (N_15768,N_11117,N_12997);
nor U15769 (N_15769,N_10375,N_10356);
or U15770 (N_15770,N_12002,N_14966);
nand U15771 (N_15771,N_13228,N_12176);
and U15772 (N_15772,N_10794,N_14672);
nor U15773 (N_15773,N_12398,N_11977);
nand U15774 (N_15774,N_13255,N_11327);
nand U15775 (N_15775,N_11854,N_12521);
and U15776 (N_15776,N_14090,N_14396);
nand U15777 (N_15777,N_10774,N_10703);
nand U15778 (N_15778,N_11026,N_12566);
nor U15779 (N_15779,N_14255,N_11290);
or U15780 (N_15780,N_14541,N_12169);
or U15781 (N_15781,N_11698,N_10924);
nor U15782 (N_15782,N_12895,N_14730);
and U15783 (N_15783,N_12987,N_12204);
and U15784 (N_15784,N_10174,N_13021);
and U15785 (N_15785,N_14820,N_10060);
and U15786 (N_15786,N_13070,N_10844);
nor U15787 (N_15787,N_11065,N_14039);
or U15788 (N_15788,N_10731,N_13860);
nor U15789 (N_15789,N_14631,N_10587);
and U15790 (N_15790,N_13752,N_14875);
and U15791 (N_15791,N_13858,N_13563);
and U15792 (N_15792,N_11675,N_14561);
and U15793 (N_15793,N_14192,N_12640);
and U15794 (N_15794,N_11522,N_11395);
or U15795 (N_15795,N_13212,N_11528);
or U15796 (N_15796,N_14564,N_13458);
xor U15797 (N_15797,N_11492,N_10429);
or U15798 (N_15798,N_14646,N_10603);
and U15799 (N_15799,N_13702,N_14545);
or U15800 (N_15800,N_12154,N_14021);
or U15801 (N_15801,N_12822,N_14227);
nand U15802 (N_15802,N_13631,N_13588);
and U15803 (N_15803,N_12937,N_10085);
or U15804 (N_15804,N_13220,N_11403);
nand U15805 (N_15805,N_12035,N_14085);
nor U15806 (N_15806,N_13697,N_13106);
and U15807 (N_15807,N_11656,N_13878);
and U15808 (N_15808,N_12136,N_11781);
nand U15809 (N_15809,N_11682,N_14850);
nand U15810 (N_15810,N_10700,N_14171);
nor U15811 (N_15811,N_14276,N_13257);
or U15812 (N_15812,N_13516,N_12653);
nor U15813 (N_15813,N_14365,N_14826);
nor U15814 (N_15814,N_11753,N_10920);
or U15815 (N_15815,N_11058,N_11401);
nor U15816 (N_15816,N_12166,N_10228);
nand U15817 (N_15817,N_13532,N_14704);
nand U15818 (N_15818,N_11178,N_14120);
or U15819 (N_15819,N_14553,N_10728);
or U15820 (N_15820,N_12482,N_14239);
and U15821 (N_15821,N_14836,N_10784);
or U15822 (N_15822,N_13751,N_10425);
nand U15823 (N_15823,N_12096,N_11239);
and U15824 (N_15824,N_12209,N_12094);
or U15825 (N_15825,N_12221,N_12382);
and U15826 (N_15826,N_12815,N_10828);
nor U15827 (N_15827,N_12311,N_12662);
and U15828 (N_15828,N_14422,N_13185);
nor U15829 (N_15829,N_11945,N_10900);
or U15830 (N_15830,N_12776,N_10439);
nor U15831 (N_15831,N_10484,N_10170);
nor U15832 (N_15832,N_13634,N_12697);
and U15833 (N_15833,N_14828,N_14299);
nor U15834 (N_15834,N_14917,N_13014);
nand U15835 (N_15835,N_11643,N_14765);
nand U15836 (N_15836,N_13108,N_11539);
or U15837 (N_15837,N_14550,N_13530);
or U15838 (N_15838,N_13526,N_12609);
and U15839 (N_15839,N_11697,N_12180);
and U15840 (N_15840,N_13580,N_12910);
or U15841 (N_15841,N_10449,N_12896);
nand U15842 (N_15842,N_10061,N_10455);
nand U15843 (N_15843,N_14549,N_13816);
nor U15844 (N_15844,N_13010,N_13134);
nand U15845 (N_15845,N_10705,N_13657);
or U15846 (N_15846,N_10586,N_13337);
and U15847 (N_15847,N_14929,N_13022);
and U15848 (N_15848,N_12119,N_10460);
and U15849 (N_15849,N_13033,N_13863);
nor U15850 (N_15850,N_10031,N_13304);
and U15851 (N_15851,N_10140,N_13740);
nor U15852 (N_15852,N_11158,N_10160);
nand U15853 (N_15853,N_13179,N_13590);
nor U15854 (N_15854,N_13845,N_10505);
nand U15855 (N_15855,N_11507,N_13705);
nor U15856 (N_15856,N_13334,N_13609);
nand U15857 (N_15857,N_12488,N_14481);
nand U15858 (N_15858,N_13639,N_13041);
or U15859 (N_15859,N_11613,N_12471);
or U15860 (N_15860,N_12530,N_14769);
and U15861 (N_15861,N_10948,N_14610);
or U15862 (N_15862,N_13313,N_11616);
and U15863 (N_15863,N_14391,N_14629);
nor U15864 (N_15864,N_11212,N_12647);
nor U15865 (N_15865,N_10834,N_10838);
nand U15866 (N_15866,N_11337,N_11684);
or U15867 (N_15867,N_11746,N_11439);
nor U15868 (N_15868,N_14100,N_12884);
nand U15869 (N_15869,N_14662,N_12612);
or U15870 (N_15870,N_11732,N_11760);
or U15871 (N_15871,N_12477,N_10032);
nor U15872 (N_15872,N_10697,N_10810);
or U15873 (N_15873,N_14233,N_12057);
or U15874 (N_15874,N_12607,N_12817);
or U15875 (N_15875,N_10334,N_13244);
nor U15876 (N_15876,N_12461,N_12852);
or U15877 (N_15877,N_12022,N_10579);
nor U15878 (N_15878,N_10006,N_10988);
and U15879 (N_15879,N_12826,N_13724);
nor U15880 (N_15880,N_13403,N_12313);
nor U15881 (N_15881,N_14125,N_13147);
and U15882 (N_15882,N_14439,N_10335);
nor U15883 (N_15883,N_13572,N_10252);
or U15884 (N_15884,N_13534,N_10304);
nand U15885 (N_15885,N_11790,N_13427);
and U15886 (N_15886,N_10496,N_14725);
and U15887 (N_15887,N_10362,N_10102);
nor U15888 (N_15888,N_14310,N_14375);
and U15889 (N_15889,N_13120,N_13044);
nor U15890 (N_15890,N_13143,N_11132);
or U15891 (N_15891,N_10724,N_11051);
nor U15892 (N_15892,N_12203,N_11567);
and U15893 (N_15893,N_13556,N_10866);
nor U15894 (N_15894,N_13826,N_11752);
and U15895 (N_15895,N_10979,N_14294);
and U15896 (N_15896,N_12947,N_11364);
and U15897 (N_15897,N_14444,N_11243);
and U15898 (N_15898,N_12847,N_10644);
or U15899 (N_15899,N_14016,N_13000);
xnor U15900 (N_15900,N_10811,N_11793);
and U15901 (N_15901,N_12269,N_12280);
nand U15902 (N_15902,N_10312,N_14967);
nor U15903 (N_15903,N_10296,N_12143);
or U15904 (N_15904,N_10943,N_10038);
nor U15905 (N_15905,N_11797,N_14942);
or U15906 (N_15906,N_14452,N_14857);
nor U15907 (N_15907,N_11262,N_12267);
and U15908 (N_15908,N_14206,N_10469);
nand U15909 (N_15909,N_10837,N_14713);
nor U15910 (N_15910,N_14611,N_14432);
nand U15911 (N_15911,N_14183,N_10884);
nor U15912 (N_15912,N_14267,N_10822);
nor U15913 (N_15913,N_11334,N_11444);
nand U15914 (N_15914,N_14328,N_14118);
and U15915 (N_15915,N_12525,N_10673);
nand U15916 (N_15916,N_13528,N_10559);
and U15917 (N_15917,N_10188,N_10877);
and U15918 (N_15918,N_13061,N_10865);
and U15919 (N_15919,N_11173,N_12130);
nand U15920 (N_15920,N_11094,N_11638);
nor U15921 (N_15921,N_13051,N_12663);
or U15922 (N_15922,N_10885,N_11662);
nand U15923 (N_15923,N_12582,N_14940);
nand U15924 (N_15924,N_12989,N_14409);
or U15925 (N_15925,N_11162,N_12685);
and U15926 (N_15926,N_14944,N_13062);
nand U15927 (N_15927,N_13785,N_13570);
nand U15928 (N_15928,N_14885,N_10655);
or U15929 (N_15929,N_14156,N_10597);
nand U15930 (N_15930,N_12684,N_12670);
nor U15931 (N_15931,N_11311,N_11017);
or U15932 (N_15932,N_14246,N_12042);
nor U15933 (N_15933,N_11122,N_10531);
nand U15934 (N_15934,N_10340,N_10332);
or U15935 (N_15935,N_11022,N_12127);
and U15936 (N_15936,N_10221,N_14716);
and U15937 (N_15937,N_10069,N_11294);
and U15938 (N_15938,N_10001,N_14568);
or U15939 (N_15939,N_12544,N_12897);
nand U15940 (N_15940,N_13779,N_14665);
nor U15941 (N_15941,N_12135,N_13781);
nand U15942 (N_15942,N_12905,N_12492);
or U15943 (N_15943,N_13849,N_11815);
and U15944 (N_15944,N_11336,N_12235);
nand U15945 (N_15945,N_11160,N_10022);
and U15946 (N_15946,N_10368,N_14480);
and U15947 (N_15947,N_12333,N_12585);
nor U15948 (N_15948,N_10255,N_10020);
nand U15949 (N_15949,N_12748,N_12140);
nand U15950 (N_15950,N_13319,N_10687);
or U15951 (N_15951,N_12964,N_11078);
nand U15952 (N_15952,N_14312,N_12514);
and U15953 (N_15953,N_11644,N_13247);
nand U15954 (N_15954,N_11037,N_11864);
or U15955 (N_15955,N_12342,N_13744);
and U15956 (N_15956,N_13396,N_13049);
or U15957 (N_15957,N_12403,N_13799);
nand U15958 (N_15958,N_10625,N_11263);
and U15959 (N_15959,N_13083,N_13983);
or U15960 (N_15960,N_11333,N_11821);
nor U15961 (N_15961,N_14890,N_11859);
or U15962 (N_15962,N_13944,N_11805);
nand U15963 (N_15963,N_13380,N_13170);
or U15964 (N_15964,N_10472,N_14931);
or U15965 (N_15965,N_12518,N_11012);
xnor U15966 (N_15966,N_12170,N_14431);
nand U15967 (N_15967,N_14058,N_14112);
xor U15968 (N_15968,N_11087,N_11414);
and U15969 (N_15969,N_14300,N_14572);
nand U15970 (N_15970,N_13460,N_10698);
and U15971 (N_15971,N_10632,N_10755);
or U15972 (N_15972,N_12710,N_13105);
nor U15973 (N_15973,N_12553,N_10184);
and U15974 (N_15974,N_10642,N_14032);
nor U15975 (N_15975,N_14013,N_12483);
and U15976 (N_15976,N_12522,N_11195);
nor U15977 (N_15977,N_12561,N_12999);
nor U15978 (N_15978,N_14321,N_12325);
and U15979 (N_15979,N_13772,N_11835);
and U15980 (N_15980,N_10400,N_10763);
nor U15981 (N_15981,N_11380,N_11292);
and U15982 (N_15982,N_12118,N_14179);
nor U15983 (N_15983,N_11210,N_10122);
nor U15984 (N_15984,N_10186,N_14104);
nor U15985 (N_15985,N_11080,N_12487);
or U15986 (N_15986,N_14699,N_12032);
and U15987 (N_15987,N_14700,N_10118);
nor U15988 (N_15988,N_11126,N_12787);
and U15989 (N_15989,N_10018,N_13175);
nand U15990 (N_15990,N_14258,N_12857);
nand U15991 (N_15991,N_13252,N_11935);
nand U15992 (N_15992,N_12890,N_12439);
nor U15993 (N_15993,N_14134,N_13731);
nor U15994 (N_15994,N_10610,N_13287);
nor U15995 (N_15995,N_14694,N_14195);
xnor U15996 (N_15996,N_14130,N_12911);
or U15997 (N_15997,N_12813,N_12213);
and U15998 (N_15998,N_11989,N_10128);
nor U15999 (N_15999,N_14803,N_10430);
and U16000 (N_16000,N_11435,N_13621);
or U16001 (N_16001,N_12519,N_13474);
nand U16002 (N_16002,N_11689,N_11720);
and U16003 (N_16003,N_12216,N_12453);
nor U16004 (N_16004,N_14554,N_14578);
or U16005 (N_16005,N_12397,N_13906);
and U16006 (N_16006,N_13098,N_10316);
and U16007 (N_16007,N_12051,N_13090);
nand U16008 (N_16008,N_11852,N_13709);
and U16009 (N_16009,N_10725,N_14507);
nand U16010 (N_16010,N_11504,N_11787);
or U16011 (N_16011,N_13871,N_11800);
or U16012 (N_16012,N_12671,N_11344);
and U16013 (N_16013,N_11571,N_13394);
and U16014 (N_16014,N_13644,N_10083);
and U16015 (N_16015,N_14327,N_10555);
nand U16016 (N_16016,N_12944,N_13101);
nor U16017 (N_16017,N_14679,N_11968);
or U16018 (N_16018,N_12074,N_13810);
nor U16019 (N_16019,N_11345,N_12745);
nand U16020 (N_16020,N_11000,N_11556);
nand U16021 (N_16021,N_14989,N_11250);
nor U16022 (N_16022,N_11308,N_12046);
or U16023 (N_16023,N_13635,N_12551);
nor U16024 (N_16024,N_10176,N_11404);
and U16025 (N_16025,N_12447,N_13197);
nand U16026 (N_16026,N_13918,N_12618);
nand U16027 (N_16027,N_12298,N_11242);
nand U16028 (N_16028,N_10726,N_10538);
nor U16029 (N_16029,N_13714,N_13547);
nand U16030 (N_16030,N_11098,N_14065);
nor U16031 (N_16031,N_11853,N_12744);
and U16032 (N_16032,N_13656,N_10092);
nand U16033 (N_16033,N_12655,N_12534);
or U16034 (N_16034,N_11194,N_12796);
or U16035 (N_16035,N_14770,N_10566);
nand U16036 (N_16036,N_14546,N_14138);
nand U16037 (N_16037,N_14423,N_13716);
and U16038 (N_16038,N_12606,N_14454);
xor U16039 (N_16039,N_11649,N_12012);
and U16040 (N_16040,N_14598,N_13694);
nand U16041 (N_16041,N_14226,N_13964);
nand U16042 (N_16042,N_11718,N_14172);
nor U16043 (N_16043,N_13241,N_14814);
nand U16044 (N_16044,N_10582,N_12389);
nand U16045 (N_16045,N_10633,N_14456);
and U16046 (N_16046,N_10216,N_11349);
or U16047 (N_16047,N_11647,N_11601);
and U16048 (N_16048,N_12763,N_13016);
or U16049 (N_16049,N_12839,N_10630);
and U16050 (N_16050,N_13477,N_10839);
and U16051 (N_16051,N_12564,N_11997);
nand U16052 (N_16052,N_11681,N_14459);
nor U16053 (N_16053,N_14790,N_11479);
or U16054 (N_16054,N_14822,N_10488);
nand U16055 (N_16055,N_12672,N_11419);
and U16056 (N_16056,N_12476,N_12424);
or U16057 (N_16057,N_10246,N_11446);
nor U16058 (N_16058,N_13550,N_14505);
and U16059 (N_16059,N_13814,N_11373);
nor U16060 (N_16060,N_13978,N_11352);
nand U16061 (N_16061,N_13476,N_14918);
or U16062 (N_16062,N_12465,N_12863);
nor U16063 (N_16063,N_10285,N_13620);
nor U16064 (N_16064,N_10831,N_11356);
or U16065 (N_16065,N_14158,N_12296);
and U16066 (N_16066,N_14362,N_10909);
and U16067 (N_16067,N_10151,N_13940);
nor U16068 (N_16068,N_11005,N_14207);
or U16069 (N_16069,N_10264,N_13761);
nand U16070 (N_16070,N_13654,N_12401);
nand U16071 (N_16071,N_13723,N_12645);
or U16072 (N_16072,N_12421,N_14720);
and U16073 (N_16073,N_12688,N_10769);
nor U16074 (N_16074,N_10797,N_11919);
nor U16075 (N_16075,N_14580,N_11148);
nor U16076 (N_16076,N_10619,N_14202);
nand U16077 (N_16077,N_11323,N_13486);
or U16078 (N_16078,N_10508,N_11775);
and U16079 (N_16079,N_13113,N_11077);
nor U16080 (N_16080,N_10612,N_11906);
and U16081 (N_16081,N_11476,N_10945);
and U16082 (N_16082,N_13649,N_13102);
or U16083 (N_16083,N_13397,N_14951);
nor U16084 (N_16084,N_11705,N_12692);
nand U16085 (N_16085,N_12085,N_14721);
and U16086 (N_16086,N_14238,N_14204);
or U16087 (N_16087,N_13382,N_13126);
or U16088 (N_16088,N_11956,N_13956);
and U16089 (N_16089,N_12804,N_14557);
and U16090 (N_16090,N_12678,N_10676);
or U16091 (N_16091,N_13720,N_13229);
or U16092 (N_16092,N_13385,N_11836);
and U16093 (N_16093,N_11736,N_12444);
nor U16094 (N_16094,N_11742,N_11428);
or U16095 (N_16095,N_10266,N_12108);
nand U16096 (N_16096,N_14143,N_13298);
and U16097 (N_16097,N_10193,N_10315);
nand U16098 (N_16098,N_13523,N_11267);
nand U16099 (N_16099,N_14048,N_10464);
nand U16100 (N_16100,N_14271,N_13768);
and U16101 (N_16101,N_11264,N_10624);
and U16102 (N_16102,N_12020,N_13216);
or U16103 (N_16103,N_11179,N_12728);
nand U16104 (N_16104,N_14671,N_12644);
and U16105 (N_16105,N_10983,N_10681);
and U16106 (N_16106,N_13509,N_14476);
and U16107 (N_16107,N_11390,N_14852);
nor U16108 (N_16108,N_12479,N_13202);
or U16109 (N_16109,N_11772,N_12624);
or U16110 (N_16110,N_14303,N_11359);
nand U16111 (N_16111,N_14283,N_10470);
and U16112 (N_16112,N_10549,N_14668);
or U16113 (N_16113,N_12505,N_12372);
nand U16114 (N_16114,N_11532,N_13678);
nand U16115 (N_16115,N_13643,N_12772);
and U16116 (N_16116,N_10458,N_13524);
nor U16117 (N_16117,N_12724,N_14017);
or U16118 (N_16118,N_12774,N_14723);
nand U16119 (N_16119,N_12305,N_11722);
or U16120 (N_16120,N_10507,N_13624);
nor U16121 (N_16121,N_12996,N_11278);
xor U16122 (N_16122,N_12965,N_13372);
nor U16123 (N_16123,N_13297,N_12862);
nor U16124 (N_16124,N_11449,N_11502);
or U16125 (N_16125,N_12786,N_10013);
nand U16126 (N_16126,N_10704,N_10854);
nor U16127 (N_16127,N_10202,N_14881);
nand U16128 (N_16128,N_13171,N_12411);
nand U16129 (N_16129,N_14361,N_11691);
and U16130 (N_16130,N_11955,N_11369);
and U16131 (N_16131,N_11215,N_12276);
nand U16132 (N_16132,N_10829,N_10646);
nor U16133 (N_16133,N_13855,N_11181);
or U16134 (N_16134,N_11020,N_10875);
or U16135 (N_16135,N_10028,N_12321);
nand U16136 (N_16136,N_14357,N_14907);
or U16137 (N_16137,N_14532,N_14487);
nor U16138 (N_16138,N_10503,N_13092);
nor U16139 (N_16139,N_10722,N_11868);
and U16140 (N_16140,N_10119,N_12975);
nor U16141 (N_16141,N_10929,N_14844);
and U16142 (N_16142,N_13145,N_14682);
and U16143 (N_16143,N_14297,N_11174);
and U16144 (N_16144,N_13430,N_13217);
nand U16145 (N_16145,N_13807,N_14883);
or U16146 (N_16146,N_10719,N_14717);
nor U16147 (N_16147,N_10238,N_14201);
nor U16148 (N_16148,N_10114,N_11994);
or U16149 (N_16149,N_11964,N_10516);
nand U16150 (N_16150,N_10233,N_13640);
nor U16151 (N_16151,N_12840,N_10388);
nor U16152 (N_16152,N_12379,N_12080);
and U16153 (N_16153,N_12693,N_13696);
or U16154 (N_16154,N_10121,N_13616);
nand U16155 (N_16155,N_10422,N_14174);
or U16156 (N_16156,N_11325,N_10426);
or U16157 (N_16157,N_12604,N_12789);
xor U16158 (N_16158,N_11034,N_10326);
or U16159 (N_16159,N_14900,N_13152);
and U16160 (N_16160,N_12025,N_12148);
nand U16161 (N_16161,N_12229,N_14026);
or U16162 (N_16162,N_14029,N_10256);
nor U16163 (N_16163,N_13564,N_13358);
nor U16164 (N_16164,N_13177,N_13966);
or U16165 (N_16165,N_14761,N_12846);
nor U16166 (N_16166,N_14463,N_12797);
or U16167 (N_16167,N_13336,N_11008);
nor U16168 (N_16168,N_12524,N_13953);
and U16169 (N_16169,N_10172,N_13844);
or U16170 (N_16170,N_13204,N_13839);
and U16171 (N_16171,N_14330,N_13484);
nand U16172 (N_16172,N_14997,N_10096);
or U16173 (N_16173,N_10284,N_13186);
nor U16174 (N_16174,N_13389,N_11055);
nand U16175 (N_16175,N_11591,N_13700);
nand U16176 (N_16176,N_13759,N_14800);
nor U16177 (N_16177,N_14394,N_12100);
nand U16178 (N_16178,N_10935,N_11335);
nand U16179 (N_16179,N_13651,N_10057);
and U16180 (N_16180,N_13465,N_11218);
nor U16181 (N_16181,N_12329,N_11188);
nand U16182 (N_16182,N_12665,N_11694);
nand U16183 (N_16183,N_14674,N_12446);
or U16184 (N_16184,N_11733,N_11254);
nand U16185 (N_16185,N_10098,N_14443);
nand U16186 (N_16186,N_10350,N_14302);
or U16187 (N_16187,N_10595,N_10666);
or U16188 (N_16188,N_12746,N_14381);
nor U16189 (N_16189,N_14046,N_11231);
nor U16190 (N_16190,N_14208,N_13767);
and U16191 (N_16191,N_12040,N_12306);
or U16192 (N_16192,N_14044,N_12738);
or U16193 (N_16193,N_13025,N_14127);
and U16194 (N_16194,N_13058,N_14870);
nand U16195 (N_16195,N_11995,N_12686);
and U16196 (N_16196,N_13496,N_11615);
or U16197 (N_16197,N_14565,N_14260);
nor U16198 (N_16198,N_12569,N_14057);
or U16199 (N_16199,N_10142,N_11594);
or U16200 (N_16200,N_12634,N_10502);
nand U16201 (N_16201,N_14998,N_14355);
and U16202 (N_16202,N_10305,N_14701);
nand U16203 (N_16203,N_14077,N_12779);
or U16204 (N_16204,N_13762,N_12432);
and U16205 (N_16205,N_13613,N_13577);
nor U16206 (N_16206,N_11220,N_10480);
and U16207 (N_16207,N_11818,N_13633);
and U16208 (N_16208,N_12422,N_14697);
and U16209 (N_16209,N_14936,N_11521);
nand U16210 (N_16210,N_11152,N_10116);
or U16211 (N_16211,N_12892,N_13775);
and U16212 (N_16212,N_10434,N_12865);
nor U16213 (N_16213,N_12458,N_14209);
and U16214 (N_16214,N_12506,N_11044);
nor U16215 (N_16215,N_14693,N_12299);
or U16216 (N_16216,N_11575,N_14860);
or U16217 (N_16217,N_10997,N_14678);
or U16218 (N_16218,N_14592,N_14692);
nand U16219 (N_16219,N_11190,N_14247);
and U16220 (N_16220,N_14867,N_10894);
nand U16221 (N_16221,N_10354,N_14243);
and U16222 (N_16222,N_14864,N_13409);
nor U16223 (N_16223,N_11312,N_14777);
and U16224 (N_16224,N_12450,N_10825);
nor U16225 (N_16225,N_13352,N_12928);
or U16226 (N_16226,N_14488,N_13732);
and U16227 (N_16227,N_10711,N_14470);
or U16228 (N_16228,N_10450,N_12499);
nand U16229 (N_16229,N_14466,N_10367);
and U16230 (N_16230,N_12723,N_11161);
nor U16231 (N_16231,N_10459,N_10960);
nor U16232 (N_16232,N_12171,N_13701);
nor U16233 (N_16233,N_12383,N_12434);
and U16234 (N_16234,N_14343,N_10200);
nand U16235 (N_16235,N_12635,N_13927);
nor U16236 (N_16236,N_10753,N_10906);
and U16237 (N_16237,N_14957,N_11366);
nor U16238 (N_16238,N_10337,N_13448);
and U16239 (N_16239,N_11992,N_13094);
nand U16240 (N_16240,N_13853,N_14560);
or U16241 (N_16241,N_13441,N_10091);
nor U16242 (N_16242,N_11685,N_12881);
nand U16243 (N_16243,N_12334,N_12255);
xnor U16244 (N_16244,N_13386,N_12168);
nor U16245 (N_16245,N_10637,N_10793);
nor U16246 (N_16246,N_12920,N_13331);
nand U16247 (N_16247,N_10530,N_12743);
nand U16248 (N_16248,N_14645,N_13194);
nand U16249 (N_16249,N_10298,N_14324);
xor U16250 (N_16250,N_13140,N_14804);
and U16251 (N_16251,N_10995,N_14280);
and U16252 (N_16252,N_13363,N_11138);
and U16253 (N_16253,N_12137,N_10876);
nand U16254 (N_16254,N_12289,N_13020);
and U16255 (N_16255,N_12536,N_10376);
or U16256 (N_16256,N_12353,N_14366);
or U16257 (N_16257,N_14150,N_11081);
or U16258 (N_16258,N_10922,N_11131);
and U16259 (N_16259,N_10840,N_10379);
and U16260 (N_16260,N_13350,N_13963);
and U16261 (N_16261,N_11982,N_10878);
or U16262 (N_16262,N_12256,N_11269);
nand U16263 (N_16263,N_14011,N_14691);
and U16264 (N_16264,N_14586,N_14792);
nor U16265 (N_16265,N_13315,N_12337);
nor U16266 (N_16266,N_11540,N_10980);
or U16267 (N_16267,N_10338,N_11743);
and U16268 (N_16268,N_13710,N_14818);
or U16269 (N_16269,N_13236,N_13215);
and U16270 (N_16270,N_12449,N_11707);
nand U16271 (N_16271,N_14318,N_13950);
nor U16272 (N_16272,N_12037,N_13946);
or U16273 (N_16273,N_13851,N_14801);
or U16274 (N_16274,N_11108,N_10080);
nand U16275 (N_16275,N_13975,N_14587);
nor U16276 (N_16276,N_12016,N_14854);
nor U16277 (N_16277,N_12320,N_14098);
nand U16278 (N_16278,N_10819,N_13200);
nor U16279 (N_16279,N_13426,N_13715);
nand U16280 (N_16280,N_12766,N_10045);
nor U16281 (N_16281,N_13652,N_10766);
nand U16282 (N_16282,N_12303,N_13818);
nor U16283 (N_16283,N_11822,N_14921);
nand U16284 (N_16284,N_10660,N_12674);
and U16285 (N_16285,N_11894,N_14584);
nor U16286 (N_16286,N_14397,N_10571);
nand U16287 (N_16287,N_10801,N_14062);
or U16288 (N_16288,N_11604,N_10267);
nand U16289 (N_16289,N_10065,N_13671);
nand U16290 (N_16290,N_13808,N_10260);
or U16291 (N_16291,N_14551,N_14735);
and U16292 (N_16292,N_10125,N_13475);
or U16293 (N_16293,N_11704,N_12088);
nor U16294 (N_16294,N_10361,N_14230);
nand U16295 (N_16295,N_10813,N_13998);
and U16296 (N_16296,N_11729,N_11714);
or U16297 (N_16297,N_13447,N_12270);
nor U16298 (N_16298,N_10405,N_14581);
nor U16299 (N_16299,N_11102,N_12396);
or U16300 (N_16300,N_11109,N_13433);
nand U16301 (N_16301,N_13470,N_13852);
nand U16302 (N_16302,N_11626,N_12454);
or U16303 (N_16303,N_11780,N_13436);
or U16304 (N_16304,N_13366,N_12885);
and U16305 (N_16305,N_11462,N_10027);
and U16306 (N_16306,N_13568,N_11113);
and U16307 (N_16307,N_10790,N_13471);
nand U16308 (N_16308,N_10859,N_13893);
nor U16309 (N_16309,N_13993,N_13317);
nor U16310 (N_16310,N_13518,N_12423);
nand U16311 (N_16311,N_10477,N_10963);
nor U16312 (N_16312,N_14426,N_14632);
or U16313 (N_16313,N_11842,N_13877);
and U16314 (N_16314,N_10012,N_11786);
or U16315 (N_16315,N_10947,N_13925);
and U16316 (N_16316,N_14533,N_13001);
nor U16317 (N_16317,N_11506,N_12110);
and U16318 (N_16318,N_14856,N_11039);
and U16319 (N_16319,N_11340,N_12821);
or U16320 (N_16320,N_11093,N_13872);
nand U16321 (N_16321,N_12214,N_13566);
nand U16322 (N_16322,N_12568,N_10493);
and U16323 (N_16323,N_10111,N_14441);
and U16324 (N_16324,N_13400,N_11376);
nor U16325 (N_16325,N_11271,N_10659);
nor U16326 (N_16326,N_10014,N_10129);
nand U16327 (N_16327,N_11592,N_14658);
or U16328 (N_16328,N_11089,N_14478);
nand U16329 (N_16329,N_14304,N_10858);
or U16330 (N_16330,N_10497,N_14248);
and U16331 (N_16331,N_10783,N_14754);
and U16332 (N_16332,N_12675,N_11830);
nor U16333 (N_16333,N_14637,N_10187);
and U16334 (N_16334,N_11655,N_11204);
or U16335 (N_16335,N_11755,N_14648);
nor U16336 (N_16336,N_13286,N_10201);
nor U16337 (N_16337,N_12656,N_13802);
or U16338 (N_16338,N_10209,N_12284);
or U16339 (N_16339,N_11406,N_11460);
nand U16340 (N_16340,N_14880,N_13345);
nand U16341 (N_16341,N_12664,N_14855);
nor U16342 (N_16342,N_13742,N_14924);
nor U16343 (N_16343,N_14919,N_11941);
or U16344 (N_16344,N_11837,N_14124);
nor U16345 (N_16345,N_13527,N_14170);
xor U16346 (N_16346,N_12151,N_10529);
and U16347 (N_16347,N_12574,N_11112);
nand U16348 (N_16348,N_12992,N_14879);
or U16349 (N_16349,N_12631,N_14607);
or U16350 (N_16350,N_11240,N_12658);
and U16351 (N_16351,N_12455,N_12830);
nand U16352 (N_16352,N_12304,N_12331);
nand U16353 (N_16353,N_11885,N_14866);
nor U16354 (N_16354,N_11241,N_11554);
nor U16355 (N_16355,N_14952,N_14364);
and U16356 (N_16356,N_14006,N_10628);
or U16357 (N_16357,N_11354,N_12404);
or U16358 (N_16358,N_10990,N_13013);
nor U16359 (N_16359,N_13907,N_14673);
or U16360 (N_16360,N_10798,N_11234);
nor U16361 (N_16361,N_13892,N_13037);
nor U16362 (N_16362,N_10694,N_11151);
and U16363 (N_16363,N_14352,N_14109);
nor U16364 (N_16364,N_10465,N_12064);
and U16365 (N_16365,N_12158,N_14075);
and U16366 (N_16366,N_11346,N_13882);
xnor U16367 (N_16367,N_11809,N_13084);
or U16368 (N_16368,N_11332,N_11903);
or U16369 (N_16369,N_12275,N_11030);
nor U16370 (N_16370,N_12250,N_11833);
nand U16371 (N_16371,N_11082,N_12590);
nand U16372 (N_16372,N_14601,N_11301);
and U16373 (N_16373,N_10049,N_13806);
nor U16374 (N_16374,N_10734,N_10163);
and U16375 (N_16375,N_14007,N_11041);
and U16376 (N_16376,N_10835,N_14185);
nand U16377 (N_16377,N_14802,N_14781);
and U16378 (N_16378,N_13619,N_12783);
nand U16379 (N_16379,N_13466,N_13798);
nand U16380 (N_16380,N_10923,N_13913);
nand U16381 (N_16381,N_13169,N_10351);
nor U16382 (N_16382,N_10329,N_14696);
or U16383 (N_16383,N_11676,N_14597);
nor U16384 (N_16384,N_13672,N_13233);
and U16385 (N_16385,N_11104,N_12914);
nand U16386 (N_16386,N_14894,N_13074);
nor U16387 (N_16387,N_13824,N_11560);
nand U16388 (N_16388,N_10856,N_13962);
nor U16389 (N_16389,N_13856,N_14599);
nor U16390 (N_16390,N_10179,N_10669);
nor U16391 (N_16391,N_10042,N_14834);
and U16392 (N_16392,N_13373,N_12257);
nand U16393 (N_16393,N_13408,N_10010);
nand U16394 (N_16394,N_11137,N_12539);
and U16395 (N_16395,N_12916,N_14910);
nand U16396 (N_16396,N_10075,N_10991);
nor U16397 (N_16397,N_14436,N_12239);
nand U16398 (N_16398,N_13078,N_10276);
nand U16399 (N_16399,N_12960,N_11186);
and U16400 (N_16400,N_10342,N_13837);
and U16401 (N_16401,N_13141,N_12129);
nand U16402 (N_16402,N_12683,N_14051);
nand U16403 (N_16403,N_14708,N_10574);
nand U16404 (N_16404,N_10359,N_12695);
nand U16405 (N_16405,N_11633,N_11459);
nor U16406 (N_16406,N_13491,N_12941);
or U16407 (N_16407,N_13246,N_10936);
and U16408 (N_16408,N_10423,N_14325);
nand U16409 (N_16409,N_12493,N_14388);
nor U16410 (N_16410,N_14830,N_11341);
and U16411 (N_16411,N_12034,N_11580);
and U16412 (N_16412,N_10850,N_11471);
nor U16413 (N_16413,N_13894,N_10643);
nor U16414 (N_16414,N_13093,N_14376);
nand U16415 (N_16415,N_10970,N_14084);
or U16416 (N_16416,N_12245,N_14372);
and U16417 (N_16417,N_10198,N_13320);
nor U16418 (N_16418,N_13628,N_14928);
nand U16419 (N_16419,N_14198,N_11057);
and U16420 (N_16420,N_11728,N_14983);
or U16421 (N_16421,N_11839,N_12990);
nor U16422 (N_16422,N_13214,N_12810);
nand U16423 (N_16423,N_10974,N_14492);
or U16424 (N_16424,N_10749,N_11605);
or U16425 (N_16425,N_12259,N_12115);
nand U16426 (N_16426,N_13142,N_13342);
xnor U16427 (N_16427,N_14144,N_12282);
nor U16428 (N_16428,N_11440,N_10089);
or U16429 (N_16429,N_10641,N_10482);
and U16430 (N_16430,N_12107,N_11727);
and U16431 (N_16431,N_13144,N_13923);
nor U16432 (N_16432,N_12874,N_12391);
nand U16433 (N_16433,N_10684,N_13412);
and U16434 (N_16434,N_11975,N_12001);
or U16435 (N_16435,N_14460,N_11792);
and U16436 (N_16436,N_10138,N_14472);
nor U16437 (N_16437,N_13210,N_11947);
or U16438 (N_16438,N_12286,N_12613);
or U16439 (N_16439,N_11183,N_11503);
or U16440 (N_16440,N_14724,N_10712);
and U16441 (N_16441,N_14891,N_10268);
nor U16442 (N_16442,N_11402,N_14273);
nand U16443 (N_16443,N_10699,N_13206);
or U16444 (N_16444,N_12233,N_11672);
nand U16445 (N_16445,N_13278,N_13017);
or U16446 (N_16446,N_10622,N_10568);
and U16447 (N_16447,N_10951,N_13771);
and U16448 (N_16448,N_10317,N_12625);
nor U16449 (N_16449,N_14234,N_14774);
and U16450 (N_16450,N_11590,N_14136);
nand U16451 (N_16451,N_12346,N_11351);
or U16452 (N_16452,N_14344,N_11987);
nand U16453 (N_16453,N_11016,N_13087);
nand U16454 (N_16454,N_14817,N_14231);
nor U16455 (N_16455,N_14169,N_11226);
nand U16456 (N_16456,N_14301,N_11475);
nor U16457 (N_16457,N_10387,N_10515);
nand U16458 (N_16458,N_13936,N_13357);
and U16459 (N_16459,N_13089,N_13670);
and U16460 (N_16460,N_11499,N_10109);
and U16461 (N_16461,N_12909,N_12691);
nor U16462 (N_16462,N_12661,N_10413);
nand U16463 (N_16463,N_11426,N_13085);
and U16464 (N_16464,N_10000,N_11636);
nand U16465 (N_16465,N_14072,N_10310);
or U16466 (N_16466,N_10481,N_11990);
and U16467 (N_16467,N_10108,N_12617);
nor U16468 (N_16468,N_11309,N_12307);
nor U16469 (N_16469,N_11452,N_11191);
nand U16470 (N_16470,N_10048,N_10560);
nor U16471 (N_16471,N_13760,N_11083);
or U16472 (N_16472,N_11608,N_13213);
or U16473 (N_16473,N_12702,N_13819);
nor U16474 (N_16474,N_11759,N_14166);
nand U16475 (N_16475,N_14418,N_11091);
and U16476 (N_16476,N_12971,N_13503);
nor U16477 (N_16477,N_13520,N_10629);
nand U16478 (N_16478,N_12781,N_14520);
nand U16479 (N_16479,N_11529,N_12915);
and U16480 (N_16480,N_11586,N_10414);
nor U16481 (N_16481,N_10671,N_11130);
nand U16482 (N_16482,N_10702,N_14382);
or U16483 (N_16483,N_11584,N_12919);
nand U16484 (N_16484,N_11472,N_11027);
and U16485 (N_16485,N_12091,N_13840);
nor U16486 (N_16486,N_14882,N_13166);
nand U16487 (N_16487,N_13691,N_10576);
nor U16488 (N_16488,N_11363,N_13348);
nand U16489 (N_16489,N_14846,N_12368);
nand U16490 (N_16490,N_11411,N_14993);
nor U16491 (N_16491,N_12228,N_11949);
and U16492 (N_16492,N_11572,N_12155);
nand U16493 (N_16493,N_14187,N_13122);
or U16494 (N_16494,N_10107,N_14413);
or U16495 (N_16495,N_14133,N_13219);
and U16496 (N_16496,N_13638,N_14163);
and U16497 (N_16497,N_12418,N_13495);
nor U16498 (N_16498,N_11154,N_14018);
or U16499 (N_16499,N_11544,N_10752);
nor U16500 (N_16500,N_11228,N_13584);
or U16501 (N_16501,N_12414,N_11920);
nand U16502 (N_16502,N_10968,N_13783);
nand U16503 (N_16503,N_13240,N_12162);
nor U16504 (N_16504,N_14232,N_11969);
and U16505 (N_16505,N_12554,N_14315);
nand U16506 (N_16506,N_10254,N_14128);
and U16507 (N_16507,N_10971,N_11932);
or U16508 (N_16508,N_11911,N_11768);
xnor U16509 (N_16509,N_11542,N_13168);
or U16510 (N_16510,N_14108,N_12870);
nand U16511 (N_16511,N_10159,N_13193);
nand U16512 (N_16512,N_13367,N_13987);
or U16513 (N_16513,N_11563,N_14518);
or U16514 (N_16514,N_12491,N_12144);
and U16515 (N_16515,N_10391,N_10765);
nand U16516 (N_16516,N_14036,N_14782);
or U16517 (N_16517,N_14314,N_14402);
nor U16518 (N_16518,N_12283,N_11270);
or U16519 (N_16519,N_11803,N_12977);
or U16520 (N_16520,N_13703,N_10981);
or U16521 (N_16521,N_11494,N_13529);
nand U16522 (N_16522,N_14181,N_13056);
or U16523 (N_16523,N_10191,N_11866);
nand U16524 (N_16524,N_11448,N_11660);
or U16525 (N_16525,N_13561,N_13230);
and U16526 (N_16526,N_11248,N_13757);
nor U16527 (N_16527,N_12452,N_11533);
or U16528 (N_16528,N_12799,N_12565);
nor U16529 (N_16529,N_13312,N_13727);
and U16530 (N_16530,N_10833,N_13857);
nand U16531 (N_16531,N_12936,N_11754);
or U16532 (N_16532,N_14279,N_11957);
or U16533 (N_16533,N_13151,N_11916);
nand U16534 (N_16534,N_13736,N_14684);
or U16535 (N_16535,N_14184,N_10656);
nand U16536 (N_16536,N_13322,N_12584);
or U16537 (N_16537,N_12818,N_14612);
nand U16538 (N_16538,N_12714,N_11802);
nor U16539 (N_16539,N_10670,N_10034);
nor U16540 (N_16540,N_11798,N_10072);
and U16541 (N_16541,N_11258,N_11617);
or U16542 (N_16542,N_14086,N_12545);
or U16543 (N_16543,N_10225,N_10345);
and U16544 (N_16544,N_14912,N_10689);
nand U16545 (N_16545,N_13617,N_10243);
nor U16546 (N_16546,N_11794,N_12437);
or U16547 (N_16547,N_14228,N_12801);
and U16548 (N_16548,N_12182,N_10397);
nor U16549 (N_16549,N_14805,N_14628);
or U16550 (N_16550,N_14797,N_10171);
nand U16551 (N_16551,N_11305,N_12363);
nand U16552 (N_16552,N_10433,N_11904);
nor U16553 (N_16553,N_13072,N_13941);
and U16554 (N_16554,N_13481,N_13825);
or U16555 (N_16555,N_10787,N_13439);
nand U16556 (N_16556,N_14594,N_13890);
nor U16557 (N_16557,N_11399,N_14096);
or U16558 (N_16558,N_12940,N_12588);
or U16559 (N_16559,N_12583,N_10785);
nand U16560 (N_16560,N_10978,N_14153);
nand U16561 (N_16561,N_10168,N_14263);
and U16562 (N_16562,N_10208,N_14135);
and U16563 (N_16563,N_12167,N_10720);
and U16564 (N_16564,N_13227,N_13355);
or U16565 (N_16565,N_13238,N_12160);
and U16566 (N_16566,N_11238,N_12961);
or U16567 (N_16567,N_11692,N_14513);
nand U16568 (N_16568,N_10290,N_10534);
and U16569 (N_16569,N_13687,N_13192);
and U16570 (N_16570,N_13338,N_10474);
nor U16571 (N_16571,N_14626,N_12921);
and U16572 (N_16572,N_10683,N_11651);
nand U16573 (N_16573,N_14719,N_13745);
nor U16574 (N_16574,N_11856,N_13306);
or U16575 (N_16575,N_13254,N_11493);
and U16576 (N_16576,N_14406,N_10227);
nand U16577 (N_16577,N_13195,N_13809);
and U16578 (N_16578,N_11469,N_10062);
nor U16579 (N_16579,N_11251,N_10044);
and U16580 (N_16580,N_10371,N_11384);
nor U16581 (N_16581,N_12687,N_14147);
or U16582 (N_16582,N_11641,N_13292);
nor U16583 (N_16583,N_14726,N_13359);
or U16584 (N_16584,N_12068,N_12009);
nand U16585 (N_16585,N_11700,N_10897);
nor U16586 (N_16586,N_13065,N_13914);
nand U16587 (N_16587,N_11581,N_10144);
xor U16588 (N_16588,N_11814,N_12117);
and U16589 (N_16589,N_10431,N_12226);
nor U16590 (N_16590,N_12668,N_12509);
or U16591 (N_16591,N_13443,N_11631);
and U16592 (N_16592,N_13846,N_10476);
or U16593 (N_16593,N_11669,N_14034);
nand U16594 (N_16594,N_10401,N_10236);
and U16595 (N_16595,N_10517,N_14675);
nor U16596 (N_16596,N_11114,N_13949);
nand U16597 (N_16597,N_11683,N_11902);
nand U16598 (N_16598,N_12716,N_14949);
and U16599 (N_16599,N_10245,N_12473);
and U16600 (N_16600,N_13256,N_10791);
nor U16601 (N_16601,N_14946,N_13364);
nor U16602 (N_16602,N_12195,N_10846);
or U16603 (N_16603,N_13632,N_14268);
nand U16604 (N_16604,N_12793,N_14272);
or U16605 (N_16605,N_14865,N_10383);
or U16606 (N_16606,N_14262,N_10194);
and U16607 (N_16607,N_11235,N_10614);
and U16608 (N_16608,N_10678,N_11249);
nand U16609 (N_16609,N_11543,N_12597);
and U16610 (N_16610,N_12113,N_12043);
nand U16611 (N_16611,N_10578,N_13666);
or U16612 (N_16612,N_10853,N_11184);
and U16613 (N_16613,N_14240,N_13596);
nand U16614 (N_16614,N_12425,N_12105);
nand U16615 (N_16615,N_10086,N_11006);
and U16616 (N_16616,N_10764,N_14635);
nand U16617 (N_16617,N_13717,N_10580);
and U16618 (N_16618,N_14609,N_13303);
nor U16619 (N_16619,N_10149,N_11167);
nand U16620 (N_16620,N_12069,N_13136);
or U16621 (N_16621,N_10984,N_14004);
and U16622 (N_16622,N_12770,N_14030);
nor U16623 (N_16623,N_10394,N_10741);
nand U16624 (N_16624,N_13104,N_14224);
or U16625 (N_16625,N_14760,N_14245);
nand U16626 (N_16626,N_13748,N_13116);
and U16627 (N_16627,N_12541,N_11688);
and U16628 (N_16628,N_13811,N_14787);
nand U16629 (N_16629,N_12721,N_14600);
or U16630 (N_16630,N_10436,N_10223);
and U16631 (N_16631,N_14939,N_10845);
and U16632 (N_16632,N_14477,N_14117);
nor U16633 (N_16633,N_10302,N_11673);
nand U16634 (N_16634,N_12066,N_12287);
nand U16635 (N_16635,N_14903,N_14845);
or U16636 (N_16636,N_11980,N_14019);
and U16637 (N_16637,N_11872,N_14427);
and U16638 (N_16638,N_14193,N_11076);
and U16639 (N_16639,N_12247,N_12834);
nor U16640 (N_16640,N_11838,N_10820);
nor U16641 (N_16641,N_12178,N_10490);
nor U16642 (N_16642,N_13335,N_12281);
nor U16643 (N_16643,N_10537,N_11219);
nand U16644 (N_16644,N_10157,N_13539);
or U16645 (N_16645,N_14639,N_10448);
and U16646 (N_16646,N_12887,N_14490);
xor U16647 (N_16647,N_11118,N_14537);
or U16648 (N_16648,N_14326,N_12819);
or U16649 (N_16649,N_11518,N_12072);
nor U16650 (N_16650,N_13555,N_11547);
nand U16651 (N_16651,N_14510,N_10003);
or U16652 (N_16652,N_11774,N_12097);
or U16653 (N_16653,N_12557,N_12038);
and U16654 (N_16654,N_10263,N_13378);
nor U16655 (N_16655,N_14313,N_12013);
or U16656 (N_16656,N_10039,N_10239);
nand U16657 (N_16657,N_10081,N_13086);
or U16658 (N_16658,N_10976,N_14306);
and U16659 (N_16659,N_12433,N_11937);
or U16660 (N_16660,N_13749,N_13904);
and U16661 (N_16661,N_12611,N_12703);
nand U16662 (N_16662,N_10931,N_11014);
or U16663 (N_16663,N_14582,N_10771);
nand U16664 (N_16664,N_14831,N_12456);
and U16665 (N_16665,N_11813,N_10396);
nand U16666 (N_16666,N_12065,N_10029);
nand U16667 (N_16667,N_14621,N_10807);
and U16668 (N_16668,N_13307,N_12351);
nor U16669 (N_16669,N_12258,N_10667);
nor U16670 (N_16670,N_10224,N_10489);
nand U16671 (N_16671,N_11648,N_11891);
nor U16672 (N_16672,N_11307,N_12378);
nand U16673 (N_16673,N_14624,N_13608);
nand U16674 (N_16674,N_13711,N_12362);
nand U16675 (N_16675,N_12994,N_10585);
nor U16676 (N_16676,N_11289,N_11558);
and U16677 (N_16677,N_11671,N_10213);
or U16678 (N_16678,N_10150,N_12019);
nand U16679 (N_16679,N_11930,N_11953);
nor U16680 (N_16680,N_13841,N_14796);
or U16681 (N_16681,N_14711,N_14311);
nand U16682 (N_16682,N_14740,N_11614);
nand U16683 (N_16683,N_10416,N_12048);
nand U16684 (N_16684,N_12983,N_10921);
nor U16685 (N_16685,N_14076,N_11019);
and U16686 (N_16686,N_14762,N_13788);
nand U16687 (N_16687,N_10514,N_13279);
or U16688 (N_16688,N_12142,N_11485);
or U16689 (N_16689,N_14976,N_14840);
nor U16690 (N_16690,N_12833,N_14282);
nor U16691 (N_16691,N_12292,N_14028);
and U16692 (N_16692,N_10662,N_10881);
or U16693 (N_16693,N_12241,N_13525);
and U16694 (N_16694,N_13054,N_10964);
nor U16695 (N_16695,N_13059,N_14686);
nor U16696 (N_16696,N_14095,N_11463);
nor U16697 (N_16697,N_10410,N_11966);
nor U16698 (N_16698,N_13513,N_12594);
and U16699 (N_16699,N_11611,N_10377);
and U16700 (N_16700,N_14401,N_10654);
or U16701 (N_16701,N_10910,N_13954);
or U16702 (N_16702,N_10046,N_10893);
or U16703 (N_16703,N_10318,N_12364);
nand U16704 (N_16704,N_11450,N_14416);
nand U16705 (N_16705,N_10750,N_10583);
or U16706 (N_16706,N_12075,N_11741);
nand U16707 (N_16707,N_14971,N_14093);
or U16708 (N_16708,N_12317,N_11981);
nand U16709 (N_16709,N_14497,N_14566);
nand U16710 (N_16710,N_10902,N_11129);
or U16711 (N_16711,N_10665,N_12083);
or U16712 (N_16712,N_14161,N_12124);
nor U16713 (N_16713,N_13601,N_11409);
or U16714 (N_16714,N_11488,N_13347);
nand U16715 (N_16715,N_12767,N_14579);
or U16716 (N_16716,N_12598,N_10548);
nand U16717 (N_16717,N_10780,N_11635);
and U16718 (N_16718,N_12428,N_10499);
nand U16719 (N_16719,N_10235,N_11735);
or U16720 (N_16720,N_10805,N_11922);
nor U16721 (N_16721,N_11843,N_14356);
and U16722 (N_16722,N_11306,N_12384);
or U16723 (N_16723,N_12177,N_12785);
and U16724 (N_16724,N_13793,N_13034);
or U16725 (N_16725,N_12045,N_10913);
or U16726 (N_16726,N_10584,N_12078);
and U16727 (N_16727,N_14102,N_11907);
and U16728 (N_16728,N_13739,N_14651);
nand U16729 (N_16729,N_11412,N_12301);
nor U16730 (N_16730,N_11623,N_12026);
or U16731 (N_16731,N_13500,N_10406);
nor U16732 (N_16732,N_10768,N_10103);
and U16733 (N_16733,N_12802,N_11976);
nor U16734 (N_16734,N_12102,N_14446);
and U16735 (N_16735,N_12529,N_10047);
nor U16736 (N_16736,N_11831,N_12326);
or U16737 (N_16737,N_11829,N_13869);
nor U16738 (N_16738,N_10743,N_11347);
nor U16739 (N_16739,N_13623,N_11478);
nor U16740 (N_16740,N_14442,N_10895);
or U16741 (N_16741,N_10015,N_13544);
and U16742 (N_16742,N_12314,N_13489);
or U16743 (N_16743,N_11205,N_13743);
nor U16744 (N_16744,N_13942,N_13467);
nor U16745 (N_16745,N_13437,N_11316);
or U16746 (N_16746,N_13645,N_14958);
nor U16747 (N_16747,N_11519,N_10443);
nor U16748 (N_16748,N_13173,N_12188);
and U16749 (N_16749,N_13612,N_14996);
nand U16750 (N_16750,N_12737,N_11031);
nand U16751 (N_16751,N_14614,N_12800);
and U16752 (N_16752,N_10130,N_10374);
and U16753 (N_16753,N_11890,N_13420);
nor U16754 (N_16754,N_14950,N_13976);
or U16755 (N_16755,N_13540,N_11621);
or U16756 (N_16756,N_13510,N_11310);
nor U16757 (N_16757,N_10101,N_13405);
nor U16758 (N_16758,N_10730,N_11708);
nand U16759 (N_16759,N_12350,N_13542);
and U16760 (N_16760,N_13407,N_10485);
nand U16761 (N_16761,N_12106,N_13492);
and U16762 (N_16762,N_14116,N_14131);
and U16763 (N_16763,N_12959,N_10364);
and U16764 (N_16764,N_12388,N_13293);
and U16765 (N_16765,N_12578,N_12898);
or U16766 (N_16766,N_13766,N_12302);
nor U16767 (N_16767,N_12676,N_13558);
nand U16768 (N_16768,N_10847,N_13862);
nor U16769 (N_16769,N_10133,N_10916);
and U16770 (N_16770,N_10352,N_11817);
and U16771 (N_16771,N_12504,N_13919);
nand U16772 (N_16772,N_12371,N_11201);
or U16773 (N_16773,N_13948,N_10879);
nor U16774 (N_16774,N_14982,N_12950);
and U16775 (N_16775,N_14813,N_11862);
nand U16776 (N_16776,N_10258,N_10998);
and U16777 (N_16777,N_14889,N_10649);
nand U16778 (N_16778,N_11180,N_14892);
and U16779 (N_16779,N_11198,N_12555);
nand U16780 (N_16780,N_14999,N_10064);
nor U16781 (N_16781,N_13750,N_11767);
or U16782 (N_16782,N_14923,N_12060);
nor U16783 (N_16783,N_13411,N_11011);
and U16784 (N_16784,N_14807,N_11565);
or U16785 (N_16785,N_13773,N_11578);
nand U16786 (N_16786,N_14155,N_14419);
or U16787 (N_16787,N_11564,N_10291);
nor U16788 (N_16788,N_11103,N_12295);
nand U16789 (N_16789,N_11625,N_12844);
nand U16790 (N_16790,N_10270,N_14874);
nor U16791 (N_16791,N_11779,N_13354);
or U16792 (N_16792,N_10668,N_11596);
and U16793 (N_16793,N_12099,N_14515);
or U16794 (N_16794,N_12659,N_10347);
or U16795 (N_16795,N_10441,N_12929);
nor U16796 (N_16796,N_13787,N_10192);
nor U16797 (N_16797,N_13791,N_12848);
or U16798 (N_16798,N_13531,N_14219);
nor U16799 (N_16799,N_11557,N_11330);
and U16800 (N_16800,N_13154,N_12620);
or U16801 (N_16801,N_11326,N_11967);
nand U16802 (N_16802,N_12845,N_12552);
or U16803 (N_16803,N_12722,N_14986);
nor U16804 (N_16804,N_12192,N_13868);
and U16805 (N_16805,N_14063,N_11508);
or U16806 (N_16806,N_11520,N_14091);
or U16807 (N_16807,N_11107,N_11795);
and U16808 (N_16808,N_14608,N_14827);
xor U16809 (N_16809,N_12507,N_13721);
or U16810 (N_16810,N_14590,N_10740);
and U16811 (N_16811,N_13567,N_10282);
nand U16812 (N_16812,N_14798,N_13218);
nand U16813 (N_16813,N_13449,N_13585);
nor U16814 (N_16814,N_10626,N_11049);
nand U16815 (N_16815,N_12322,N_12573);
nand U16816 (N_16816,N_12669,N_13068);
nand U16817 (N_16817,N_10320,N_11505);
nand U16818 (N_16818,N_10982,N_10204);
nor U16819 (N_16819,N_14945,N_12050);
and U16820 (N_16820,N_14948,N_13945);
and U16821 (N_16821,N_14757,N_13203);
nand U16822 (N_16822,N_11734,N_13490);
or U16823 (N_16823,N_13934,N_10735);
nor U16824 (N_16824,N_10863,N_10608);
nor U16825 (N_16825,N_14424,N_11895);
nor U16826 (N_16826,N_10639,N_14384);
and U16827 (N_16827,N_11870,N_12528);
or U16828 (N_16828,N_14548,N_14251);
nand U16829 (N_16829,N_11225,N_10074);
or U16830 (N_16830,N_14010,N_14620);
and U16831 (N_16831,N_10399,N_11211);
nor U16832 (N_16832,N_10486,N_12147);
nor U16833 (N_16833,N_12438,N_11331);
nand U16834 (N_16834,N_11500,N_11237);
nand U16835 (N_16835,N_10136,N_12843);
nor U16836 (N_16836,N_10898,N_12059);
nand U16837 (N_16837,N_10463,N_12806);
and U16838 (N_16838,N_14539,N_10518);
nand U16839 (N_16839,N_12592,N_10792);
nand U16840 (N_16840,N_11527,N_10398);
and U16841 (N_16841,N_10056,N_14977);
nand U16842 (N_16842,N_14712,N_12409);
nand U16843 (N_16843,N_11668,N_11587);
or U16844 (N_16844,N_14788,N_11170);
and U16845 (N_16845,N_12567,N_14168);
and U16846 (N_16846,N_10446,N_11106);
or U16847 (N_16847,N_14199,N_11060);
and U16848 (N_16848,N_10438,N_14728);
or U16849 (N_16849,N_13827,N_12357);
or U16850 (N_16850,N_13679,N_11553);
or U16851 (N_16851,N_13618,N_12189);
and U16852 (N_16852,N_12500,N_11050);
nor U16853 (N_16853,N_13284,N_10333);
and U16854 (N_16854,N_13277,N_10210);
xnor U16855 (N_16855,N_11361,N_11940);
nor U16856 (N_16856,N_12741,N_13464);
nor U16857 (N_16857,N_14535,N_12814);
nor U16858 (N_16858,N_12711,N_10946);
nand U16859 (N_16859,N_11713,N_12395);
nand U16860 (N_16860,N_13499,N_10181);
or U16861 (N_16861,N_12548,N_13604);
or U16862 (N_16862,N_11213,N_14808);
and U16863 (N_16863,N_12494,N_13968);
nor U16864 (N_16864,N_10959,N_13131);
nand U16865 (N_16865,N_13445,N_12616);
or U16866 (N_16866,N_14400,N_14895);
or U16867 (N_16867,N_10513,N_12858);
nand U16868 (N_16868,N_14351,N_14534);
or U16869 (N_16869,N_10234,N_10759);
nor U16870 (N_16870,N_11568,N_12926);
nand U16871 (N_16871,N_13150,N_12542);
or U16872 (N_16872,N_14925,N_10167);
or U16873 (N_16873,N_13097,N_14448);
nor U16874 (N_16874,N_14908,N_13270);
nor U16875 (N_16875,N_14498,N_12327);
xnor U16876 (N_16876,N_12526,N_13249);
or U16877 (N_16877,N_11541,N_12475);
and U16878 (N_16878,N_14746,N_11360);
nor U16879 (N_16879,N_13189,N_12116);
or U16880 (N_16880,N_11983,N_14160);
nor U16881 (N_16881,N_11163,N_10212);
nand U16882 (N_16882,N_12036,N_12768);
nand U16883 (N_16883,N_13521,N_10147);
nor U16884 (N_16884,N_10620,N_11321);
nand U16885 (N_16885,N_14053,N_14825);
or U16886 (N_16886,N_12718,N_13981);
nand U16887 (N_16887,N_13996,N_14793);
nor U16888 (N_16888,N_10546,N_10556);
nand U16889 (N_16889,N_10370,N_13823);
and U16890 (N_16890,N_10492,N_10950);
nor U16891 (N_16891,N_14001,N_14070);
and U16892 (N_16892,N_11394,N_12957);
or U16893 (N_16893,N_10621,N_14786);
and U16894 (N_16894,N_14110,N_10746);
xor U16895 (N_16895,N_14009,N_10451);
and U16896 (N_16896,N_12485,N_14338);
xnor U16897 (N_16897,N_14990,N_14148);
nand U16898 (N_16898,N_13898,N_10471);
and U16899 (N_16899,N_13817,N_11667);
or U16900 (N_16900,N_12935,N_10143);
nor U16901 (N_16901,N_10888,N_13419);
and U16902 (N_16902,N_13579,N_10230);
nor U16903 (N_16903,N_14558,N_12513);
and U16904 (N_16904,N_13047,N_13080);
nor U16905 (N_16905,N_10776,N_10592);
or U16906 (N_16906,N_14984,N_13641);
and U16907 (N_16907,N_12764,N_10966);
and U16908 (N_16908,N_11299,N_13063);
nor U16909 (N_16909,N_12300,N_10955);
nand U16910 (N_16910,N_11690,N_11477);
nand U16911 (N_16911,N_14690,N_12376);
and U16912 (N_16912,N_14676,N_12998);
or U16913 (N_16913,N_14165,N_11923);
nor U16914 (N_16914,N_10164,N_12725);
nor U16915 (N_16915,N_13344,N_12196);
and U16916 (N_16916,N_11261,N_13262);
and U16917 (N_16917,N_13737,N_13574);
xnor U16918 (N_16918,N_10648,N_10231);
nor U16919 (N_16919,N_14256,N_11597);
or U16920 (N_16920,N_12290,N_13201);
nand U16921 (N_16921,N_12747,N_11850);
or U16922 (N_16922,N_13753,N_10090);
nand U16923 (N_16923,N_10944,N_12489);
and U16924 (N_16924,N_11295,N_11847);
nand U16925 (N_16925,N_11144,N_13973);
nor U16926 (N_16926,N_13755,N_13989);
or U16927 (N_16927,N_10189,N_14322);
or U16928 (N_16928,N_12934,N_10672);
or U16929 (N_16929,N_10701,N_11799);
nand U16930 (N_16930,N_11092,N_11723);
and U16931 (N_16931,N_10892,N_10716);
or U16932 (N_16932,N_11128,N_11515);
nor U16933 (N_16933,N_11054,N_13726);
or U16934 (N_16934,N_11233,N_13123);
xor U16935 (N_16935,N_11288,N_14067);
or U16936 (N_16936,N_10598,N_14395);
nand U16937 (N_16937,N_13003,N_10501);
or U16938 (N_16938,N_14159,N_13991);
nand U16939 (N_16939,N_11143,N_14975);
nand U16940 (N_16940,N_11392,N_12279);
nor U16941 (N_16941,N_13132,N_11342);
or U16942 (N_16942,N_11371,N_13505);
and U16943 (N_16943,N_13158,N_10185);
or U16944 (N_16944,N_12392,N_13339);
and U16945 (N_16945,N_10025,N_12729);
nor U16946 (N_16946,N_11867,N_11496);
or U16947 (N_16947,N_14445,N_13790);
nor U16948 (N_16948,N_14778,N_13431);
nor U16949 (N_16949,N_13156,N_11236);
and U16950 (N_16950,N_12285,N_14064);
and U16951 (N_16951,N_13578,N_12431);
or U16952 (N_16952,N_12246,N_10088);
or U16953 (N_16953,N_13052,N_14902);
nand U16954 (N_16954,N_12312,N_11857);
and U16955 (N_16955,N_12262,N_11302);
or U16956 (N_16956,N_11979,N_10985);
or U16957 (N_16957,N_12511,N_11537);
and U16958 (N_16958,N_10453,N_12531);
nand U16959 (N_16959,N_13362,N_13758);
nand U16960 (N_16960,N_14698,N_14569);
or U16961 (N_16961,N_11962,N_13404);
or U16962 (N_16962,N_13234,N_13794);
nor U16963 (N_16963,N_11067,N_11209);
or U16964 (N_16964,N_14333,N_14323);
or U16965 (N_16965,N_14643,N_10182);
or U16966 (N_16966,N_13921,N_12288);
nor U16967 (N_16967,N_12076,N_10887);
nand U16968 (N_16968,N_11427,N_14559);
and U16969 (N_16969,N_10055,N_11150);
and U16970 (N_16970,N_12736,N_12824);
nand U16971 (N_16971,N_11978,N_13971);
and U16972 (N_16972,N_13381,N_12629);
and U16973 (N_16973,N_10907,N_10965);
and U16974 (N_16974,N_14970,N_14235);
nand U16975 (N_16975,N_11199,N_12415);
xnor U16976 (N_16976,N_12359,N_10440);
nand U16977 (N_16977,N_10710,N_10165);
and U16978 (N_16978,N_13920,N_10095);
or U16979 (N_16979,N_14615,N_14241);
nand U16980 (N_16980,N_11265,N_12836);
nor U16981 (N_16981,N_14317,N_12033);
nand U16982 (N_16982,N_12354,N_13280);
nand U16983 (N_16983,N_11097,N_11826);
nor U16984 (N_16984,N_11318,N_11970);
nand U16985 (N_16985,N_13163,N_13859);
and U16986 (N_16986,N_11612,N_11040);
and U16987 (N_16987,N_11284,N_10424);
nor U16988 (N_16988,N_11607,N_13675);
and U16989 (N_16989,N_14705,N_12021);
nand U16990 (N_16990,N_10117,N_14074);
or U16991 (N_16991,N_12217,N_11276);
and U16992 (N_16992,N_11958,N_13406);
and U16993 (N_16993,N_14739,N_12690);
and U16994 (N_16994,N_13456,N_12457);
xor U16995 (N_16995,N_14583,N_12297);
or U16996 (N_16996,N_13780,N_11045);
and U16997 (N_16997,N_12740,N_10468);
or U16998 (N_16998,N_11429,N_11531);
nor U16999 (N_16999,N_12402,N_13560);
nor U17000 (N_17000,N_11255,N_11884);
and U17001 (N_17001,N_10054,N_14878);
or U17002 (N_17002,N_12265,N_11438);
and U17003 (N_17003,N_13030,N_11120);
or U17004 (N_17004,N_13833,N_10139);
or U17005 (N_17005,N_11686,N_13803);
nor U17006 (N_17006,N_12027,N_12187);
and U17007 (N_17007,N_10331,N_10693);
or U17008 (N_17008,N_10037,N_12869);
or U17009 (N_17009,N_11153,N_10222);
and U17010 (N_17010,N_12520,N_11808);
or U17011 (N_17011,N_13842,N_12366);
or U17012 (N_17012,N_11348,N_11650);
and U17013 (N_17013,N_13088,N_12469);
xor U17014 (N_17014,N_11253,N_11381);
nor U17015 (N_17015,N_11702,N_10306);
or U17016 (N_17016,N_10190,N_13535);
and U17017 (N_17017,N_14731,N_12646);
and U17018 (N_17018,N_10207,N_10280);
nand U17019 (N_17019,N_10385,N_14089);
nand U17020 (N_17020,N_12855,N_11202);
nor U17021 (N_17021,N_12201,N_13784);
and U17022 (N_17022,N_10782,N_14906);
and U17023 (N_17023,N_11304,N_14617);
or U17024 (N_17024,N_11486,N_11887);
and U17025 (N_17025,N_14506,N_11046);
nand U17026 (N_17026,N_14337,N_10408);
or U17027 (N_17027,N_14524,N_10526);
and U17028 (N_17028,N_12924,N_14215);
nor U17029 (N_17029,N_11216,N_10004);
nand U17030 (N_17030,N_11501,N_11776);
or U17031 (N_17031,N_14045,N_13007);
and U17032 (N_17032,N_14689,N_13733);
nor U17033 (N_17033,N_12416,N_13417);
nor U17034 (N_17034,N_14773,N_12549);
and U17035 (N_17035,N_10524,N_10536);
nand U17036 (N_17036,N_11047,N_11208);
nand U17037 (N_17037,N_10677,N_10058);
nand U17038 (N_17038,N_13454,N_10322);
or U17039 (N_17039,N_10680,N_10178);
nand U17040 (N_17040,N_11737,N_12760);
nor U17041 (N_17041,N_11328,N_12231);
or U17042 (N_17042,N_14399,N_13690);
or U17043 (N_17043,N_11487,N_10849);
nand U17044 (N_17044,N_14284,N_14412);
or U17045 (N_17045,N_14059,N_13308);
and U17046 (N_17046,N_12614,N_13067);
nand U17047 (N_17047,N_11881,N_13376);
nor U17048 (N_17048,N_14525,N_13850);
and U17049 (N_17049,N_14373,N_13506);
nor U17050 (N_17050,N_11410,N_12484);
nand U17051 (N_17051,N_12835,N_13805);
or U17052 (N_17052,N_13683,N_12184);
and U17053 (N_17053,N_11658,N_12223);
and U17054 (N_17054,N_14901,N_13653);
and U17055 (N_17055,N_12031,N_11620);
or U17056 (N_17056,N_12111,N_14236);
nor U17057 (N_17057,N_13128,N_11273);
nand U17058 (N_17058,N_11140,N_10928);
and U17059 (N_17059,N_12092,N_12352);
nand U17060 (N_17060,N_14927,N_10115);
or U17061 (N_17061,N_13424,N_12794);
and U17062 (N_17062,N_14980,N_10987);
or U17063 (N_17063,N_11757,N_10874);
nand U17064 (N_17064,N_10395,N_12798);
or U17065 (N_17065,N_14420,N_13747);
or U17066 (N_17066,N_14020,N_11901);
and U17067 (N_17067,N_12925,N_14516);
nor U17068 (N_17068,N_10889,N_10973);
nor U17069 (N_17069,N_12464,N_13867);
nand U17070 (N_17070,N_14092,N_11355);
and U17071 (N_17071,N_13453,N_10532);
nor U17072 (N_17072,N_10927,N_14503);
nand U17073 (N_17073,N_10739,N_14149);
and U17074 (N_17074,N_12430,N_10148);
and U17075 (N_17075,N_10127,N_12445);
nor U17076 (N_17076,N_12367,N_13951);
and U17077 (N_17077,N_11282,N_13800);
nor U17078 (N_17078,N_11257,N_12927);
and U17079 (N_17079,N_10718,N_13242);
or U17080 (N_17080,N_14641,N_10588);
nand U17081 (N_17081,N_11422,N_13328);
nor U17082 (N_17082,N_13478,N_12436);
or U17083 (N_17083,N_10161,N_14047);
or U17084 (N_17084,N_14935,N_13599);
nor U17085 (N_17085,N_13224,N_11934);
and U17086 (N_17086,N_14972,N_13324);
nor U17087 (N_17087,N_13912,N_12730);
nand U17088 (N_17088,N_13341,N_10307);
and U17089 (N_17089,N_11595,N_11844);
or U17090 (N_17090,N_10862,N_12230);
nand U17091 (N_17091,N_10690,N_14654);
and U17092 (N_17092,N_14360,N_11423);
nand U17093 (N_17093,N_13008,N_10203);
nor U17094 (N_17094,N_10473,N_13908);
nand U17095 (N_17095,N_13040,N_12771);
nand U17096 (N_17096,N_12638,N_13391);
nand U17097 (N_17097,N_12602,N_10616);
and U17098 (N_17098,N_12908,N_10809);
or U17099 (N_17099,N_13865,N_13383);
and U17100 (N_17100,N_13955,N_12232);
nand U17101 (N_17101,N_11931,N_11701);
nand U17102 (N_17102,N_14012,N_14178);
nand U17103 (N_17103,N_12315,N_10330);
nand U17104 (N_17104,N_13487,N_11473);
nor U17105 (N_17105,N_12899,N_14451);
or U17106 (N_17106,N_14080,N_10145);
and U17107 (N_17107,N_11873,N_13820);
or U17108 (N_17108,N_14715,N_14806);
nand U17109 (N_17109,N_12878,N_12605);
nor U17110 (N_17110,N_12412,N_14332);
or U17111 (N_17111,N_10346,N_11882);
nor U17112 (N_17112,N_12677,N_12174);
or U17113 (N_17113,N_10707,N_12435);
or U17114 (N_17114,N_11538,N_14591);
nor U17115 (N_17115,N_10093,N_14666);
nand U17116 (N_17116,N_10744,N_13326);
or U17117 (N_17117,N_11182,N_10483);
or U17118 (N_17118,N_14119,N_13164);
nor U17119 (N_17119,N_12868,N_12946);
and U17120 (N_17120,N_14097,N_13479);
and U17121 (N_17121,N_13291,N_12727);
and U17122 (N_17122,N_10097,N_14729);
and U17123 (N_17123,N_11747,N_14896);
or U17124 (N_17124,N_13712,N_10975);
nand U17125 (N_17125,N_10977,N_13361);
or U17126 (N_17126,N_10999,N_11555);
or U17127 (N_17127,N_13422,N_14577);
nor U17128 (N_17128,N_11609,N_10427);
nand U17129 (N_17129,N_14574,N_14812);
or U17130 (N_17130,N_10009,N_13290);
and U17131 (N_17131,N_13933,N_13507);
nor U17132 (N_17132,N_12888,N_13469);
nand U17133 (N_17133,N_13137,N_13763);
nor U17134 (N_17134,N_11133,N_14661);
xor U17135 (N_17135,N_11111,N_11726);
nor U17136 (N_17136,N_13066,N_13174);
and U17137 (N_17137,N_14821,N_13115);
nand U17138 (N_17138,N_11350,N_10903);
or U17139 (N_17139,N_10328,N_14897);
nor U17140 (N_17140,N_14428,N_12873);
or U17141 (N_17141,N_13365,N_14307);
nand U17142 (N_17142,N_12234,N_11313);
nor U17143 (N_17143,N_13668,N_11628);
nor U17144 (N_17144,N_14687,N_11388);
or U17145 (N_17145,N_12015,N_14652);
nor U17146 (N_17146,N_14528,N_14988);
and U17147 (N_17147,N_13019,N_12777);
and U17148 (N_17148,N_14496,N_10152);
nor U17149 (N_17149,N_10539,N_14853);
or U17150 (N_17150,N_11009,N_12316);
nor U17151 (N_17151,N_13961,N_10882);
nor U17152 (N_17152,N_12067,N_13930);
or U17153 (N_17153,N_13043,N_14776);
and U17154 (N_17154,N_12784,N_11959);
nor U17155 (N_17155,N_10275,N_13610);
nand U17156 (N_17156,N_11602,N_11622);
or U17157 (N_17157,N_13321,N_14056);
nand U17158 (N_17158,N_11559,N_11637);
or U17159 (N_17159,N_13444,N_12093);
or U17160 (N_17160,N_10613,N_10696);
and U17161 (N_17161,N_13117,N_13012);
or U17162 (N_17162,N_14264,N_14379);
and U17163 (N_17163,N_12891,N_12405);
nor U17164 (N_17164,N_12958,N_14254);
and U17165 (N_17165,N_13884,N_13435);
nor U17166 (N_17166,N_14295,N_12701);
nor U17167 (N_17167,N_14529,N_13073);
nand U17168 (N_17168,N_13591,N_14987);
and U17169 (N_17169,N_13473,N_12134);
nand U17170 (N_17170,N_12719,N_12679);
and U17171 (N_17171,N_12651,N_11524);
nand U17172 (N_17172,N_12079,N_12827);
nor U17173 (N_17173,N_14623,N_12966);
or U17174 (N_17174,N_12861,N_12061);
nand U17175 (N_17175,N_12131,N_13318);
or U17176 (N_17176,N_14316,N_13032);
or U17177 (N_17177,N_11480,N_13187);
nor U17178 (N_17178,N_12056,N_12340);
xor U17179 (N_17179,N_10456,N_14964);
or U17180 (N_17180,N_13957,N_14499);
nor U17181 (N_17181,N_13310,N_12632);
and U17182 (N_17182,N_11386,N_11134);
and U17183 (N_17183,N_14220,N_13155);
nor U17184 (N_17184,N_13754,N_12008);
nor U17185 (N_17185,N_12345,N_10411);
nor U17186 (N_17186,N_12385,N_12319);
or U17187 (N_17187,N_12610,N_14383);
nand U17188 (N_17188,N_12791,N_13023);
and U17189 (N_17189,N_12248,N_12394);
xor U17190 (N_17190,N_13288,N_11899);
nor U17191 (N_17191,N_10663,N_14369);
nand U17192 (N_17192,N_12210,N_12550);
nand U17193 (N_17193,N_10553,N_11585);
nand U17194 (N_17194,N_10023,N_11155);
and U17195 (N_17195,N_11824,N_10392);
and U17196 (N_17196,N_14752,N_12185);
nor U17197 (N_17197,N_10363,N_12696);
nor U17198 (N_17198,N_10912,N_12374);
nand U17199 (N_17199,N_12854,N_10804);
or U17200 (N_17200,N_11430,N_11986);
nor U17201 (N_17201,N_11417,N_10952);
or U17202 (N_17202,N_11863,N_14636);
or U17203 (N_17203,N_14008,N_13512);
or U17204 (N_17204,N_14433,N_12823);
nand U17205 (N_17205,N_12860,N_14756);
nor U17206 (N_17206,N_14082,N_14334);
nand U17207 (N_17207,N_12010,N_12058);
and U17208 (N_17208,N_11785,N_13024);
nand U17209 (N_17209,N_14094,N_11434);
and U17210 (N_17210,N_10253,N_12328);
nand U17211 (N_17211,N_11072,N_10939);
nor U17212 (N_17212,N_10421,N_12152);
or U17213 (N_17213,N_13901,N_11545);
or U17214 (N_17214,N_13972,N_12587);
and U17215 (N_17215,N_10591,N_10059);
and U17216 (N_17216,N_12579,N_14329);
nand U17217 (N_17217,N_13055,N_11677);
nand U17218 (N_17218,N_12157,N_13330);
nor U17219 (N_17219,N_12018,N_11942);
and U17220 (N_17220,N_11788,N_14849);
nand U17221 (N_17221,N_13821,N_12599);
nor U17222 (N_17222,N_10479,N_14758);
nand U17223 (N_17223,N_14229,N_14969);
and U17224 (N_17224,N_12948,N_14290);
or U17225 (N_17225,N_10504,N_11905);
nor U17226 (N_17226,N_11807,N_12938);
and U17227 (N_17227,N_11420,N_13517);
or U17228 (N_17228,N_12608,N_10957);
nor U17229 (N_17229,N_10105,N_10919);
nand U17230 (N_17230,N_13096,N_14212);
xnor U17231 (N_17231,N_13522,N_13057);
nor U17232 (N_17232,N_12481,N_14811);
or U17233 (N_17233,N_11075,N_13497);
nand U17234 (N_17234,N_12417,N_12375);
or U17235 (N_17235,N_10257,N_11035);
or U17236 (N_17236,N_13450,N_10301);
nor U17237 (N_17237,N_10197,N_11317);
nor U17238 (N_17238,N_13665,N_13296);
nor U17239 (N_17239,N_10554,N_11415);
nand U17240 (N_17240,N_13425,N_13583);
nor U17241 (N_17241,N_12400,N_12841);
and U17242 (N_17242,N_14173,N_13314);
or U17243 (N_17243,N_10100,N_13109);
nand U17244 (N_17244,N_12330,N_14380);
nand U17245 (N_17245,N_14743,N_10652);
nor U17246 (N_17246,N_12980,N_10339);
nand U17247 (N_17247,N_14995,N_14348);
or U17248 (N_17248,N_10543,N_10511);
nand U17249 (N_17249,N_13418,N_12755);
nor U17250 (N_17250,N_13463,N_13329);
and U17251 (N_17251,N_12689,N_10823);
or U17252 (N_17252,N_10528,N_12700);
and U17253 (N_17253,N_14824,N_14363);
nor U17254 (N_17254,N_14954,N_11730);
and U17255 (N_17255,N_12601,N_10348);
or U17256 (N_17256,N_11724,N_13546);
or U17257 (N_17257,N_13432,N_13081);
or U17258 (N_17258,N_12429,N_14530);
nor U17259 (N_17259,N_13553,N_10679);
nand U17260 (N_17260,N_14981,N_11769);
nand U17261 (N_17261,N_14653,N_10070);
nand U17262 (N_17262,N_11576,N_10864);
nor U17263 (N_17263,N_10709,N_13864);
nor U17264 (N_17264,N_14040,N_10336);
nand U17265 (N_17265,N_11101,N_14186);
nand U17266 (N_17266,N_13127,N_13854);
nand U17267 (N_17267,N_10372,N_10519);
nor U17268 (N_17268,N_11593,N_12419);
or U17269 (N_17269,N_11176,N_11382);
or U17270 (N_17270,N_14035,N_13146);
or U17271 (N_17271,N_10941,N_11431);
or U17272 (N_17272,N_14493,N_12758);
nor U17273 (N_17273,N_11032,N_13253);
nor U17274 (N_17274,N_14068,N_10786);
nand U17275 (N_17275,N_14504,N_11095);
nor U17276 (N_17276,N_10914,N_12497);
or U17277 (N_17277,N_11750,N_10432);
nor U17278 (N_17278,N_10824,N_14430);
and U17279 (N_17279,N_11408,N_11999);
nand U17280 (N_17280,N_14547,N_12805);
nor U17281 (N_17281,N_10457,N_14197);
or U17282 (N_17282,N_10521,N_12751);
and U17283 (N_17283,N_14213,N_13205);
nand U17284 (N_17284,N_11146,N_14596);
nand U17285 (N_17285,N_11061,N_11244);
nor U17286 (N_17286,N_14339,N_11878);
and U17287 (N_17287,N_14003,N_13048);
nand U17288 (N_17288,N_13159,N_12370);
or U17289 (N_17289,N_14733,N_14417);
and U17290 (N_17290,N_14308,N_12648);
and U17291 (N_17291,N_13646,N_13796);
and U17292 (N_17292,N_11145,N_10323);
or U17293 (N_17293,N_13765,N_14354);
nor U17294 (N_17294,N_12122,N_14847);
or U17295 (N_17295,N_10535,N_10565);
nor U17296 (N_17296,N_14816,N_11247);
nor U17297 (N_17297,N_12572,N_11951);
nor U17298 (N_17298,N_11652,N_13511);
or U17299 (N_17299,N_10600,N_14647);
or U17300 (N_17300,N_14157,N_13885);
nor U17301 (N_17301,N_14071,N_13018);
nor U17302 (N_17302,N_11141,N_13273);
and U17303 (N_17303,N_11416,N_10007);
nor U17304 (N_17304,N_11370,N_14722);
or U17305 (N_17305,N_14526,N_14374);
or U17306 (N_17306,N_11583,N_14453);
nor U17307 (N_17307,N_12253,N_11298);
nand U17308 (N_17308,N_12410,N_14475);
nand U17309 (N_17309,N_11943,N_11849);
nand U17310 (N_17310,N_13031,N_14872);
or U17311 (N_17311,N_12832,N_12427);
nand U17312 (N_17312,N_10601,N_10146);
nand U17313 (N_17313,N_11812,N_10071);
nor U17314 (N_17314,N_14087,N_13593);
and U17315 (N_17315,N_11858,N_10841);
nand U17316 (N_17316,N_11536,N_13119);
and U17317 (N_17317,N_11874,N_13937);
or U17318 (N_17318,N_14336,N_12879);
nand U17319 (N_17319,N_10199,N_11491);
or U17320 (N_17320,N_11804,N_13472);
nand U17321 (N_17321,N_10249,N_10596);
and U17322 (N_17322,N_12413,N_13434);
or U17323 (N_17323,N_13880,N_10751);
or U17324 (N_17324,N_14563,N_10084);
nand U17325 (N_17325,N_11552,N_14655);
or U17326 (N_17326,N_12993,N_13959);
nand U17327 (N_17327,N_14780,N_10076);
nand U17328 (N_17328,N_13176,N_12969);
nand U17329 (N_17329,N_14249,N_10294);
nor U17330 (N_17330,N_12726,N_14991);
or U17331 (N_17331,N_14000,N_10196);
nor U17332 (N_17332,N_14764,N_11828);
nor U17333 (N_17333,N_13515,N_12871);
or U17334 (N_17334,N_14877,N_11483);
nand U17335 (N_17335,N_10067,N_11391);
and U17336 (N_17336,N_14414,N_11879);
or U17337 (N_17337,N_14479,N_10132);
nor U17338 (N_17338,N_11954,N_11036);
nor U17339 (N_17339,N_13157,N_11914);
or U17340 (N_17340,N_12474,N_14081);
nor U17341 (N_17341,N_14367,N_10244);
and U17342 (N_17342,N_14603,N_13891);
and U17343 (N_17343,N_10261,N_11825);
nor U17344 (N_17344,N_11405,N_14182);
nand U17345 (N_17345,N_13100,N_10806);
and U17346 (N_17346,N_11221,N_12149);
or U17347 (N_17347,N_10380,N_12515);
or U17348 (N_17348,N_12708,N_11665);
or U17349 (N_17349,N_11484,N_13390);
or U17350 (N_17350,N_11322,N_12323);
nor U17351 (N_17351,N_12164,N_13221);
or U17352 (N_17352,N_11069,N_12831);
nor U17353 (N_17353,N_10311,N_13118);
or U17354 (N_17354,N_14309,N_14965);
and U17355 (N_17355,N_13103,N_14359);
or U17356 (N_17356,N_14221,N_12639);
nand U17357 (N_17357,N_12175,N_10495);
nand U17358 (N_17358,N_11693,N_12622);
and U17359 (N_17359,N_12907,N_14785);
or U17360 (N_17360,N_14269,N_13682);
and U17361 (N_17361,N_13549,N_13685);
nand U17362 (N_17362,N_13699,N_11421);
nor U17363 (N_17363,N_13614,N_10277);
and U17364 (N_17364,N_10360,N_11338);
nor U17365 (N_17365,N_12641,N_12023);
nor U17366 (N_17366,N_12047,N_10358);
and U17367 (N_17367,N_11495,N_11015);
nor U17368 (N_17368,N_14434,N_13353);
and U17369 (N_17369,N_10135,N_10956);
and U17370 (N_17370,N_14913,N_14848);
nand U17371 (N_17371,N_14562,N_13384);
or U17372 (N_17372,N_11196,N_10573);
or U17373 (N_17373,N_10729,N_10215);
nor U17374 (N_17374,N_14703,N_13999);
and U17375 (N_17375,N_10378,N_13261);
or U17376 (N_17376,N_13905,N_12619);
or U17377 (N_17377,N_12062,N_10855);
nor U17378 (N_17378,N_13735,N_10289);
nand U17379 (N_17379,N_14573,N_11574);
or U17380 (N_17380,N_12968,N_11398);
nand U17381 (N_17381,N_10635,N_14101);
nand U17382 (N_17382,N_14292,N_10035);
xor U17383 (N_17383,N_11362,N_14868);
nor U17384 (N_17384,N_14088,N_12876);
and U17385 (N_17385,N_11232,N_14377);
and U17386 (N_17386,N_12984,N_14869);
nor U17387 (N_17387,N_11456,N_13729);
and U17388 (N_17388,N_13970,N_12206);
or U17389 (N_17389,N_12596,N_11663);
nand U17390 (N_17390,N_12956,N_11400);
nand U17391 (N_17391,N_12084,N_14274);
nand U17392 (N_17392,N_14014,N_10562);
or U17393 (N_17393,N_11088,N_12077);
and U17394 (N_17394,N_14494,N_10915);
nand U17395 (N_17395,N_10051,N_12448);
or U17396 (N_17396,N_11642,N_14319);
nor U17397 (N_17397,N_12762,N_14287);
or U17398 (N_17398,N_13655,N_10747);
or U17399 (N_17399,N_12190,N_14622);
and U17400 (N_17400,N_13576,N_10688);
and U17401 (N_17401,N_13571,N_12294);
nand U17402 (N_17402,N_13245,N_12699);
or U17403 (N_17403,N_10617,N_13379);
and U17404 (N_17404,N_10899,N_13537);
nor U17405 (N_17405,N_13929,N_14438);
and U17406 (N_17406,N_10308,N_14079);
or U17407 (N_17407,N_10851,N_10137);
or U17408 (N_17408,N_11246,N_14298);
or U17409 (N_17409,N_11639,N_12338);
or U17410 (N_17410,N_14425,N_12498);
nor U17411 (N_17411,N_14540,N_14538);
or U17412 (N_17412,N_10830,N_12251);
or U17413 (N_17413,N_13980,N_12792);
nor U17414 (N_17414,N_12717,N_12981);
nor U17415 (N_17415,N_10293,N_11320);
nand U17416 (N_17416,N_12486,N_10240);
nand U17417 (N_17417,N_14447,N_11925);
and U17418 (N_17418,N_13188,N_14861);
nor U17419 (N_17419,N_10017,N_14485);
xnor U17420 (N_17420,N_10564,N_11100);
nor U17421 (N_17421,N_10756,N_12138);
nor U17422 (N_17422,N_11871,N_10052);
xor U17423 (N_17423,N_14278,N_13686);
nand U17424 (N_17424,N_13026,N_12560);
or U17425 (N_17425,N_13922,N_10533);
and U17426 (N_17426,N_10631,N_10926);
and U17427 (N_17427,N_14486,N_13629);
nand U17428 (N_17428,N_12853,N_13990);
xor U17429 (N_17429,N_12867,N_13191);
and U17430 (N_17430,N_13485,N_13139);
and U17431 (N_17431,N_12039,N_10558);
and U17432 (N_17432,N_14663,N_14200);
and U17433 (N_17433,N_13581,N_12720);
nand U17434 (N_17434,N_12244,N_11811);
nor U17435 (N_17435,N_11169,N_11425);
and U17436 (N_17436,N_12581,N_10645);
or U17437 (N_17437,N_12377,N_14543);
nand U17438 (N_17438,N_10325,N_13009);
nor U17439 (N_17439,N_11598,N_11709);
nand U17440 (N_17440,N_12274,N_14915);
and U17441 (N_17441,N_11851,N_14385);
or U17442 (N_17442,N_14049,N_10692);
xor U17443 (N_17443,N_12467,N_11562);
and U17444 (N_17444,N_12820,N_10295);
nor U17445 (N_17445,N_13172,N_11783);
nand U17446 (N_17446,N_12643,N_13075);
or U17447 (N_17447,N_14567,N_12731);
nand U17448 (N_17448,N_12532,N_13647);
or U17449 (N_17449,N_11059,N_10905);
nand U17450 (N_17450,N_14669,N_12139);
nor U17451 (N_17451,N_11135,N_11353);
or U17452 (N_17452,N_11367,N_12126);
nor U17453 (N_17453,N_12215,N_10462);
or U17454 (N_17454,N_14468,N_12923);
and U17455 (N_17455,N_11489,N_14137);
and U17456 (N_17456,N_13369,N_10073);
nand U17457 (N_17457,N_13611,N_10265);
nor U17458 (N_17458,N_11139,N_13295);
nand U17459 (N_17459,N_12163,N_11971);
and U17460 (N_17460,N_10005,N_11629);
nand U17461 (N_17461,N_10407,N_11550);
nand U17462 (N_17462,N_11283,N_10500);
or U17463 (N_17463,N_13095,N_12000);
or U17464 (N_17464,N_10066,N_13446);
or U17465 (N_17465,N_12586,N_11068);
nor U17466 (N_17466,N_11453,N_14167);
and U17467 (N_17467,N_10487,N_10043);
and U17468 (N_17468,N_13428,N_14823);
nand U17469 (N_17469,N_11913,N_13575);
nand U17470 (N_17470,N_11880,N_10594);
and U17471 (N_17471,N_11770,N_13573);
or U17472 (N_17472,N_13598,N_13926);
nor U17473 (N_17473,N_13725,N_14041);
and U17474 (N_17474,N_14190,N_11071);
and U17475 (N_17475,N_12161,N_14649);
or U17476 (N_17476,N_10777,N_12864);
nand U17477 (N_17477,N_10918,N_10714);
and U17478 (N_17478,N_12636,N_10547);
nand U17479 (N_17479,N_14542,N_10561);
or U17480 (N_17480,N_12951,N_12657);
xnor U17481 (N_17481,N_13911,N_10868);
nor U17482 (N_17482,N_11716,N_14242);
nand U17483 (N_17483,N_14440,N_11441);
or U17484 (N_17484,N_13947,N_12652);
or U17485 (N_17485,N_10972,N_13045);
or U17486 (N_17486,N_11277,N_11589);
nand U17487 (N_17487,N_11116,N_11588);
and U17488 (N_17488,N_13569,N_12224);
nor U17489 (N_17489,N_13504,N_11861);
nor U17490 (N_17490,N_13309,N_13797);
nand U17491 (N_17491,N_12809,N_10832);
and U17492 (N_17492,N_13876,N_14886);
xnor U17493 (N_17493,N_13248,N_14745);
nand U17494 (N_17494,N_13541,N_10180);
nor U17495 (N_17495,N_13272,N_10259);
nor U17496 (N_17496,N_12559,N_10789);
or U17497 (N_17497,N_11378,N_12753);
and U17498 (N_17498,N_12335,N_10313);
and U17499 (N_17499,N_12778,N_12011);
and U17500 (N_17500,N_14048,N_12113);
or U17501 (N_17501,N_10467,N_14255);
nand U17502 (N_17502,N_10677,N_14741);
nand U17503 (N_17503,N_13714,N_10822);
and U17504 (N_17504,N_13808,N_11748);
nor U17505 (N_17505,N_13425,N_12739);
or U17506 (N_17506,N_13248,N_12961);
and U17507 (N_17507,N_13532,N_11154);
or U17508 (N_17508,N_14238,N_10668);
and U17509 (N_17509,N_11889,N_10074);
or U17510 (N_17510,N_12072,N_13018);
nor U17511 (N_17511,N_12526,N_10979);
and U17512 (N_17512,N_12510,N_14828);
nand U17513 (N_17513,N_11164,N_11165);
and U17514 (N_17514,N_14227,N_14507);
nand U17515 (N_17515,N_11608,N_14391);
nand U17516 (N_17516,N_14474,N_14684);
nor U17517 (N_17517,N_14631,N_13929);
nand U17518 (N_17518,N_10862,N_11711);
nand U17519 (N_17519,N_10100,N_10011);
or U17520 (N_17520,N_10639,N_14558);
and U17521 (N_17521,N_11241,N_12387);
or U17522 (N_17522,N_14845,N_10610);
or U17523 (N_17523,N_14679,N_13910);
nor U17524 (N_17524,N_10670,N_13096);
nor U17525 (N_17525,N_13312,N_12402);
and U17526 (N_17526,N_14916,N_14016);
nor U17527 (N_17527,N_11073,N_10437);
and U17528 (N_17528,N_11786,N_12911);
and U17529 (N_17529,N_11237,N_12679);
or U17530 (N_17530,N_14098,N_14333);
and U17531 (N_17531,N_10767,N_12827);
nand U17532 (N_17532,N_13720,N_10743);
or U17533 (N_17533,N_11800,N_10052);
and U17534 (N_17534,N_12792,N_12197);
nand U17535 (N_17535,N_12822,N_13280);
or U17536 (N_17536,N_11449,N_12515);
or U17537 (N_17537,N_12813,N_10647);
nor U17538 (N_17538,N_10678,N_14955);
nor U17539 (N_17539,N_11703,N_10931);
and U17540 (N_17540,N_11360,N_10691);
nor U17541 (N_17541,N_12822,N_11814);
nor U17542 (N_17542,N_11906,N_13641);
or U17543 (N_17543,N_14684,N_11601);
or U17544 (N_17544,N_14909,N_14847);
nand U17545 (N_17545,N_13520,N_12209);
and U17546 (N_17546,N_12712,N_13996);
nand U17547 (N_17547,N_11439,N_12006);
nand U17548 (N_17548,N_13704,N_13987);
nor U17549 (N_17549,N_12387,N_10520);
nand U17550 (N_17550,N_14125,N_12664);
nand U17551 (N_17551,N_12628,N_13085);
nand U17552 (N_17552,N_12329,N_14539);
nor U17553 (N_17553,N_14257,N_12850);
and U17554 (N_17554,N_11853,N_10170);
and U17555 (N_17555,N_11585,N_14252);
or U17556 (N_17556,N_14636,N_11278);
nor U17557 (N_17557,N_14172,N_14435);
nand U17558 (N_17558,N_14721,N_13643);
nor U17559 (N_17559,N_10820,N_14017);
nor U17560 (N_17560,N_11518,N_14360);
and U17561 (N_17561,N_14678,N_14021);
nand U17562 (N_17562,N_11751,N_12479);
and U17563 (N_17563,N_13739,N_10387);
nand U17564 (N_17564,N_13223,N_13316);
nand U17565 (N_17565,N_11703,N_11146);
nor U17566 (N_17566,N_10510,N_12551);
or U17567 (N_17567,N_10617,N_10831);
nand U17568 (N_17568,N_11497,N_14749);
nor U17569 (N_17569,N_11609,N_10051);
nor U17570 (N_17570,N_13974,N_13501);
and U17571 (N_17571,N_11074,N_14666);
or U17572 (N_17572,N_14259,N_12335);
nand U17573 (N_17573,N_11070,N_14870);
nand U17574 (N_17574,N_11085,N_10414);
or U17575 (N_17575,N_10644,N_11425);
nand U17576 (N_17576,N_12603,N_14843);
or U17577 (N_17577,N_12559,N_11937);
nand U17578 (N_17578,N_11971,N_12973);
and U17579 (N_17579,N_11560,N_12375);
xnor U17580 (N_17580,N_13954,N_14944);
and U17581 (N_17581,N_10752,N_10196);
nor U17582 (N_17582,N_11691,N_12213);
nor U17583 (N_17583,N_12842,N_10125);
nor U17584 (N_17584,N_13457,N_10805);
and U17585 (N_17585,N_10533,N_11123);
and U17586 (N_17586,N_10984,N_10278);
or U17587 (N_17587,N_11577,N_11104);
nor U17588 (N_17588,N_14992,N_10862);
or U17589 (N_17589,N_12430,N_10104);
nand U17590 (N_17590,N_14912,N_14062);
nand U17591 (N_17591,N_11211,N_14369);
nand U17592 (N_17592,N_11562,N_13980);
and U17593 (N_17593,N_13590,N_10336);
nor U17594 (N_17594,N_13394,N_14717);
and U17595 (N_17595,N_14949,N_12306);
or U17596 (N_17596,N_12551,N_13171);
and U17597 (N_17597,N_10440,N_12610);
nor U17598 (N_17598,N_12956,N_13739);
nand U17599 (N_17599,N_14007,N_14162);
nand U17600 (N_17600,N_14948,N_12047);
nor U17601 (N_17601,N_13220,N_11162);
or U17602 (N_17602,N_12218,N_10484);
and U17603 (N_17603,N_13032,N_10339);
nor U17604 (N_17604,N_10906,N_14159);
or U17605 (N_17605,N_14103,N_13227);
or U17606 (N_17606,N_10873,N_13476);
nor U17607 (N_17607,N_10673,N_13927);
or U17608 (N_17608,N_11517,N_10776);
nor U17609 (N_17609,N_14747,N_10004);
or U17610 (N_17610,N_10384,N_11760);
and U17611 (N_17611,N_10409,N_11314);
nor U17612 (N_17612,N_13855,N_10648);
xnor U17613 (N_17613,N_10460,N_11709);
or U17614 (N_17614,N_10821,N_13635);
and U17615 (N_17615,N_12957,N_10875);
and U17616 (N_17616,N_14156,N_10259);
and U17617 (N_17617,N_13186,N_14830);
nor U17618 (N_17618,N_12509,N_13642);
xor U17619 (N_17619,N_12990,N_12108);
or U17620 (N_17620,N_11334,N_12339);
nand U17621 (N_17621,N_10037,N_12308);
or U17622 (N_17622,N_11808,N_14115);
nand U17623 (N_17623,N_12327,N_10925);
nand U17624 (N_17624,N_14927,N_12137);
and U17625 (N_17625,N_11119,N_10494);
or U17626 (N_17626,N_14850,N_14676);
and U17627 (N_17627,N_10217,N_10716);
nand U17628 (N_17628,N_13852,N_10576);
nor U17629 (N_17629,N_14122,N_11838);
or U17630 (N_17630,N_13245,N_13662);
nand U17631 (N_17631,N_13970,N_12329);
nor U17632 (N_17632,N_13354,N_10634);
or U17633 (N_17633,N_14696,N_13202);
nand U17634 (N_17634,N_13601,N_14242);
or U17635 (N_17635,N_13852,N_13129);
or U17636 (N_17636,N_12469,N_14806);
nor U17637 (N_17637,N_11881,N_10398);
nor U17638 (N_17638,N_10649,N_11104);
or U17639 (N_17639,N_11426,N_12744);
nand U17640 (N_17640,N_13640,N_10565);
nand U17641 (N_17641,N_12017,N_13894);
nor U17642 (N_17642,N_12608,N_12640);
nand U17643 (N_17643,N_14533,N_10758);
nor U17644 (N_17644,N_13841,N_11514);
nand U17645 (N_17645,N_10704,N_14951);
or U17646 (N_17646,N_11896,N_14369);
nand U17647 (N_17647,N_10512,N_11428);
nand U17648 (N_17648,N_13708,N_14730);
nand U17649 (N_17649,N_13449,N_10125);
nor U17650 (N_17650,N_11917,N_10637);
nand U17651 (N_17651,N_11156,N_10965);
and U17652 (N_17652,N_11935,N_12641);
and U17653 (N_17653,N_11131,N_12007);
or U17654 (N_17654,N_11743,N_14423);
and U17655 (N_17655,N_11306,N_13300);
and U17656 (N_17656,N_13068,N_11457);
or U17657 (N_17657,N_11446,N_12756);
nor U17658 (N_17658,N_12133,N_14325);
and U17659 (N_17659,N_10468,N_10678);
and U17660 (N_17660,N_13466,N_14499);
or U17661 (N_17661,N_14737,N_13139);
and U17662 (N_17662,N_12761,N_10007);
and U17663 (N_17663,N_11696,N_10318);
or U17664 (N_17664,N_13840,N_12387);
and U17665 (N_17665,N_10021,N_12911);
nand U17666 (N_17666,N_11638,N_13567);
nand U17667 (N_17667,N_10451,N_10780);
nand U17668 (N_17668,N_11846,N_13477);
or U17669 (N_17669,N_13804,N_12812);
nor U17670 (N_17670,N_11034,N_12980);
nor U17671 (N_17671,N_10785,N_11139);
nand U17672 (N_17672,N_11057,N_11501);
nand U17673 (N_17673,N_10587,N_11061);
nor U17674 (N_17674,N_10576,N_11426);
and U17675 (N_17675,N_11573,N_11398);
nand U17676 (N_17676,N_11812,N_13401);
nand U17677 (N_17677,N_12835,N_12177);
nor U17678 (N_17678,N_14543,N_14851);
and U17679 (N_17679,N_10832,N_11739);
and U17680 (N_17680,N_12299,N_11430);
nor U17681 (N_17681,N_10637,N_10006);
and U17682 (N_17682,N_12094,N_11322);
or U17683 (N_17683,N_11726,N_12672);
and U17684 (N_17684,N_12809,N_14831);
or U17685 (N_17685,N_12444,N_12227);
nor U17686 (N_17686,N_13174,N_12144);
and U17687 (N_17687,N_13974,N_10987);
or U17688 (N_17688,N_10318,N_13791);
nor U17689 (N_17689,N_11911,N_14289);
nor U17690 (N_17690,N_14574,N_11320);
and U17691 (N_17691,N_12088,N_14004);
and U17692 (N_17692,N_13503,N_13288);
nand U17693 (N_17693,N_10216,N_11671);
and U17694 (N_17694,N_10929,N_10642);
and U17695 (N_17695,N_14044,N_10390);
nand U17696 (N_17696,N_12931,N_12093);
nor U17697 (N_17697,N_11800,N_13271);
nand U17698 (N_17698,N_14635,N_11383);
or U17699 (N_17699,N_10778,N_14842);
nand U17700 (N_17700,N_14513,N_12229);
and U17701 (N_17701,N_13534,N_12821);
nor U17702 (N_17702,N_10679,N_13482);
and U17703 (N_17703,N_13217,N_10280);
or U17704 (N_17704,N_14829,N_11778);
nand U17705 (N_17705,N_11527,N_13651);
nor U17706 (N_17706,N_11677,N_13819);
nand U17707 (N_17707,N_13115,N_10954);
nor U17708 (N_17708,N_13306,N_13770);
nor U17709 (N_17709,N_11715,N_10398);
and U17710 (N_17710,N_13780,N_10605);
nor U17711 (N_17711,N_13538,N_10602);
nor U17712 (N_17712,N_11963,N_11935);
nor U17713 (N_17713,N_11539,N_11848);
or U17714 (N_17714,N_11948,N_11392);
or U17715 (N_17715,N_12455,N_10877);
or U17716 (N_17716,N_12416,N_13216);
nand U17717 (N_17717,N_13845,N_13512);
or U17718 (N_17718,N_12005,N_11667);
nor U17719 (N_17719,N_14899,N_14476);
nand U17720 (N_17720,N_12031,N_12579);
and U17721 (N_17721,N_12545,N_11884);
nand U17722 (N_17722,N_11398,N_11289);
nor U17723 (N_17723,N_12690,N_13569);
nand U17724 (N_17724,N_14158,N_10854);
nand U17725 (N_17725,N_11016,N_10325);
and U17726 (N_17726,N_11856,N_12168);
nand U17727 (N_17727,N_11251,N_14410);
nand U17728 (N_17728,N_14355,N_11174);
and U17729 (N_17729,N_11767,N_12037);
or U17730 (N_17730,N_11954,N_11352);
nand U17731 (N_17731,N_10768,N_14749);
or U17732 (N_17732,N_10115,N_11146);
nor U17733 (N_17733,N_13447,N_12384);
or U17734 (N_17734,N_12620,N_13706);
nor U17735 (N_17735,N_13619,N_10918);
and U17736 (N_17736,N_13804,N_14980);
nor U17737 (N_17737,N_11621,N_11588);
nand U17738 (N_17738,N_10229,N_10613);
nand U17739 (N_17739,N_12406,N_10568);
and U17740 (N_17740,N_14121,N_14412);
nand U17741 (N_17741,N_14628,N_11305);
or U17742 (N_17742,N_11560,N_11695);
and U17743 (N_17743,N_12186,N_10544);
nand U17744 (N_17744,N_12780,N_12331);
nand U17745 (N_17745,N_13447,N_14200);
nor U17746 (N_17746,N_14292,N_13463);
nor U17747 (N_17747,N_14218,N_12485);
nand U17748 (N_17748,N_11546,N_12209);
or U17749 (N_17749,N_12806,N_10882);
nand U17750 (N_17750,N_13592,N_12252);
and U17751 (N_17751,N_13285,N_13194);
nand U17752 (N_17752,N_11164,N_11480);
nand U17753 (N_17753,N_10513,N_13296);
or U17754 (N_17754,N_12707,N_10848);
nand U17755 (N_17755,N_14471,N_13073);
and U17756 (N_17756,N_14115,N_14984);
or U17757 (N_17757,N_12097,N_14982);
and U17758 (N_17758,N_14242,N_10439);
nand U17759 (N_17759,N_12417,N_12204);
nor U17760 (N_17760,N_11687,N_14958);
nor U17761 (N_17761,N_10143,N_12875);
nand U17762 (N_17762,N_13435,N_10648);
or U17763 (N_17763,N_12619,N_13766);
nor U17764 (N_17764,N_14078,N_13979);
and U17765 (N_17765,N_13169,N_11567);
nor U17766 (N_17766,N_14457,N_12848);
or U17767 (N_17767,N_14843,N_13255);
and U17768 (N_17768,N_14520,N_10225);
nor U17769 (N_17769,N_14208,N_10320);
nand U17770 (N_17770,N_10794,N_11596);
nand U17771 (N_17771,N_10010,N_12707);
nor U17772 (N_17772,N_14606,N_13587);
nor U17773 (N_17773,N_12766,N_13167);
nor U17774 (N_17774,N_14065,N_10892);
nand U17775 (N_17775,N_10857,N_13618);
and U17776 (N_17776,N_13214,N_14584);
or U17777 (N_17777,N_12563,N_14428);
nand U17778 (N_17778,N_12247,N_14849);
nand U17779 (N_17779,N_12866,N_13575);
nor U17780 (N_17780,N_14675,N_13397);
and U17781 (N_17781,N_10378,N_10557);
and U17782 (N_17782,N_14204,N_14451);
nor U17783 (N_17783,N_13829,N_10635);
or U17784 (N_17784,N_11865,N_12989);
or U17785 (N_17785,N_14313,N_13488);
or U17786 (N_17786,N_13917,N_14235);
nor U17787 (N_17787,N_12827,N_13531);
nand U17788 (N_17788,N_11400,N_10585);
and U17789 (N_17789,N_10387,N_13369);
nand U17790 (N_17790,N_10006,N_13191);
nor U17791 (N_17791,N_13187,N_11479);
nor U17792 (N_17792,N_14437,N_11540);
nand U17793 (N_17793,N_14817,N_14462);
nor U17794 (N_17794,N_11174,N_13043);
nor U17795 (N_17795,N_11652,N_11804);
nand U17796 (N_17796,N_14551,N_11574);
nor U17797 (N_17797,N_10715,N_14403);
nor U17798 (N_17798,N_10416,N_10527);
nor U17799 (N_17799,N_14426,N_11842);
nand U17800 (N_17800,N_11778,N_11790);
and U17801 (N_17801,N_13423,N_12623);
and U17802 (N_17802,N_14507,N_10655);
and U17803 (N_17803,N_13417,N_10230);
nor U17804 (N_17804,N_11399,N_11209);
nand U17805 (N_17805,N_10037,N_12890);
nor U17806 (N_17806,N_14361,N_12749);
or U17807 (N_17807,N_13659,N_12361);
xnor U17808 (N_17808,N_13732,N_11075);
and U17809 (N_17809,N_12821,N_13700);
nand U17810 (N_17810,N_11074,N_14152);
or U17811 (N_17811,N_13339,N_14684);
nor U17812 (N_17812,N_10621,N_13271);
nand U17813 (N_17813,N_10077,N_13540);
and U17814 (N_17814,N_11642,N_14261);
nand U17815 (N_17815,N_10684,N_10664);
nand U17816 (N_17816,N_11140,N_14102);
and U17817 (N_17817,N_14892,N_11053);
nand U17818 (N_17818,N_13466,N_12550);
nor U17819 (N_17819,N_14975,N_10059);
and U17820 (N_17820,N_14091,N_14155);
nand U17821 (N_17821,N_10126,N_14056);
nor U17822 (N_17822,N_11765,N_14842);
or U17823 (N_17823,N_12109,N_10207);
or U17824 (N_17824,N_13489,N_10314);
nand U17825 (N_17825,N_11327,N_13664);
or U17826 (N_17826,N_10888,N_14821);
or U17827 (N_17827,N_13472,N_11400);
nor U17828 (N_17828,N_12928,N_11569);
nand U17829 (N_17829,N_13108,N_12626);
nand U17830 (N_17830,N_13233,N_11695);
nor U17831 (N_17831,N_11512,N_10920);
and U17832 (N_17832,N_14075,N_12316);
nand U17833 (N_17833,N_14953,N_13259);
or U17834 (N_17834,N_14995,N_11488);
and U17835 (N_17835,N_10487,N_14121);
and U17836 (N_17836,N_12326,N_13222);
nor U17837 (N_17837,N_12819,N_14123);
and U17838 (N_17838,N_13739,N_12862);
nor U17839 (N_17839,N_11756,N_12639);
and U17840 (N_17840,N_14207,N_11137);
or U17841 (N_17841,N_13019,N_12604);
nor U17842 (N_17842,N_12386,N_13906);
nor U17843 (N_17843,N_11869,N_14366);
nor U17844 (N_17844,N_11830,N_14718);
nor U17845 (N_17845,N_11138,N_14864);
and U17846 (N_17846,N_10460,N_11430);
nor U17847 (N_17847,N_12037,N_10428);
nand U17848 (N_17848,N_13967,N_11800);
or U17849 (N_17849,N_14969,N_11593);
or U17850 (N_17850,N_10282,N_11985);
and U17851 (N_17851,N_14359,N_14595);
and U17852 (N_17852,N_13138,N_10393);
nor U17853 (N_17853,N_12886,N_11186);
and U17854 (N_17854,N_12757,N_12117);
nor U17855 (N_17855,N_13936,N_13424);
nor U17856 (N_17856,N_12327,N_12855);
nor U17857 (N_17857,N_13529,N_11107);
or U17858 (N_17858,N_14853,N_13470);
or U17859 (N_17859,N_13702,N_14458);
nor U17860 (N_17860,N_10758,N_14746);
and U17861 (N_17861,N_14453,N_14920);
or U17862 (N_17862,N_13027,N_10656);
or U17863 (N_17863,N_12332,N_10589);
and U17864 (N_17864,N_14244,N_11250);
nor U17865 (N_17865,N_12298,N_12680);
and U17866 (N_17866,N_13648,N_14263);
or U17867 (N_17867,N_10082,N_13877);
or U17868 (N_17868,N_11131,N_14815);
nand U17869 (N_17869,N_10675,N_14989);
nand U17870 (N_17870,N_11055,N_12457);
nand U17871 (N_17871,N_14375,N_12299);
nor U17872 (N_17872,N_10125,N_10694);
or U17873 (N_17873,N_14944,N_11892);
and U17874 (N_17874,N_14674,N_14466);
or U17875 (N_17875,N_11814,N_14225);
nand U17876 (N_17876,N_14638,N_11713);
nor U17877 (N_17877,N_13843,N_10448);
nand U17878 (N_17878,N_11547,N_11982);
nand U17879 (N_17879,N_14998,N_10217);
nor U17880 (N_17880,N_14018,N_10913);
nand U17881 (N_17881,N_10377,N_13045);
nand U17882 (N_17882,N_11429,N_14911);
and U17883 (N_17883,N_11042,N_14873);
nand U17884 (N_17884,N_11067,N_11472);
and U17885 (N_17885,N_13773,N_11406);
nand U17886 (N_17886,N_13758,N_14756);
or U17887 (N_17887,N_13029,N_12883);
nor U17888 (N_17888,N_10289,N_13246);
nor U17889 (N_17889,N_14618,N_11299);
nand U17890 (N_17890,N_14904,N_11685);
nor U17891 (N_17891,N_11331,N_10211);
or U17892 (N_17892,N_13094,N_12491);
and U17893 (N_17893,N_10161,N_12545);
nand U17894 (N_17894,N_13543,N_11702);
nand U17895 (N_17895,N_10790,N_10542);
or U17896 (N_17896,N_11861,N_13905);
nor U17897 (N_17897,N_10167,N_13562);
and U17898 (N_17898,N_13343,N_14062);
or U17899 (N_17899,N_13935,N_11708);
nor U17900 (N_17900,N_11204,N_11571);
nand U17901 (N_17901,N_10848,N_14318);
nand U17902 (N_17902,N_10429,N_13707);
nor U17903 (N_17903,N_13301,N_13995);
nand U17904 (N_17904,N_11714,N_14805);
nand U17905 (N_17905,N_12617,N_10778);
and U17906 (N_17906,N_12544,N_12466);
nor U17907 (N_17907,N_13460,N_12474);
nor U17908 (N_17908,N_12465,N_14253);
nor U17909 (N_17909,N_11013,N_14457);
or U17910 (N_17910,N_14511,N_11236);
or U17911 (N_17911,N_10118,N_12375);
or U17912 (N_17912,N_14550,N_14884);
or U17913 (N_17913,N_10958,N_11410);
nand U17914 (N_17914,N_14880,N_14959);
nand U17915 (N_17915,N_12557,N_12516);
and U17916 (N_17916,N_13849,N_12937);
nor U17917 (N_17917,N_14101,N_13768);
nor U17918 (N_17918,N_13922,N_14488);
and U17919 (N_17919,N_12470,N_14885);
and U17920 (N_17920,N_12428,N_11843);
nor U17921 (N_17921,N_14491,N_12747);
nor U17922 (N_17922,N_13649,N_10390);
or U17923 (N_17923,N_11264,N_12415);
nand U17924 (N_17924,N_11598,N_12908);
and U17925 (N_17925,N_14097,N_10500);
nand U17926 (N_17926,N_12042,N_10616);
and U17927 (N_17927,N_13098,N_12102);
and U17928 (N_17928,N_11845,N_10503);
nand U17929 (N_17929,N_11098,N_11179);
nor U17930 (N_17930,N_12230,N_12042);
and U17931 (N_17931,N_12546,N_13754);
and U17932 (N_17932,N_13457,N_14823);
nand U17933 (N_17933,N_10703,N_12914);
and U17934 (N_17934,N_13432,N_11871);
nand U17935 (N_17935,N_13224,N_13385);
and U17936 (N_17936,N_13884,N_10866);
or U17937 (N_17937,N_13020,N_13903);
nor U17938 (N_17938,N_13283,N_14171);
nor U17939 (N_17939,N_11442,N_10802);
nand U17940 (N_17940,N_11229,N_14049);
nand U17941 (N_17941,N_11393,N_12097);
and U17942 (N_17942,N_11060,N_12536);
nand U17943 (N_17943,N_12633,N_11399);
or U17944 (N_17944,N_12176,N_11949);
and U17945 (N_17945,N_12815,N_11722);
and U17946 (N_17946,N_11376,N_13132);
or U17947 (N_17947,N_14694,N_14850);
nand U17948 (N_17948,N_12255,N_10745);
nor U17949 (N_17949,N_11965,N_10677);
nand U17950 (N_17950,N_10392,N_10463);
nand U17951 (N_17951,N_11596,N_11845);
nor U17952 (N_17952,N_14125,N_14429);
or U17953 (N_17953,N_11508,N_12508);
or U17954 (N_17954,N_14138,N_14806);
or U17955 (N_17955,N_14214,N_11322);
and U17956 (N_17956,N_10818,N_13054);
or U17957 (N_17957,N_12082,N_14135);
nand U17958 (N_17958,N_10414,N_13256);
and U17959 (N_17959,N_13661,N_12446);
or U17960 (N_17960,N_11063,N_12252);
nor U17961 (N_17961,N_12381,N_12939);
or U17962 (N_17962,N_13479,N_12986);
or U17963 (N_17963,N_14439,N_12619);
nor U17964 (N_17964,N_11420,N_10266);
and U17965 (N_17965,N_13910,N_13705);
nand U17966 (N_17966,N_12223,N_10914);
and U17967 (N_17967,N_13328,N_14725);
nor U17968 (N_17968,N_11167,N_10930);
nand U17969 (N_17969,N_10848,N_10129);
nor U17970 (N_17970,N_12776,N_14580);
or U17971 (N_17971,N_13968,N_12557);
or U17972 (N_17972,N_10030,N_10126);
nor U17973 (N_17973,N_13245,N_11533);
xnor U17974 (N_17974,N_14196,N_14857);
nor U17975 (N_17975,N_14196,N_10299);
and U17976 (N_17976,N_13171,N_11446);
nand U17977 (N_17977,N_11463,N_10335);
nand U17978 (N_17978,N_14772,N_12685);
or U17979 (N_17979,N_11195,N_13089);
nand U17980 (N_17980,N_12244,N_10714);
nand U17981 (N_17981,N_13426,N_14297);
nand U17982 (N_17982,N_13048,N_12414);
nand U17983 (N_17983,N_11448,N_12789);
nor U17984 (N_17984,N_11660,N_10435);
nand U17985 (N_17985,N_14697,N_14035);
or U17986 (N_17986,N_10362,N_13004);
and U17987 (N_17987,N_14139,N_14579);
nor U17988 (N_17988,N_12458,N_11019);
xnor U17989 (N_17989,N_12607,N_14154);
nand U17990 (N_17990,N_14626,N_14244);
and U17991 (N_17991,N_14941,N_10406);
and U17992 (N_17992,N_13195,N_14189);
nor U17993 (N_17993,N_14457,N_10673);
nand U17994 (N_17994,N_14454,N_10593);
and U17995 (N_17995,N_12448,N_12430);
nor U17996 (N_17996,N_12116,N_12200);
and U17997 (N_17997,N_12846,N_12948);
and U17998 (N_17998,N_14911,N_11613);
nor U17999 (N_17999,N_12265,N_12225);
and U18000 (N_18000,N_14999,N_14053);
or U18001 (N_18001,N_12375,N_11673);
nor U18002 (N_18002,N_14546,N_13377);
nand U18003 (N_18003,N_10345,N_13466);
or U18004 (N_18004,N_11664,N_10518);
and U18005 (N_18005,N_12114,N_14886);
and U18006 (N_18006,N_12682,N_11406);
nor U18007 (N_18007,N_12183,N_12391);
and U18008 (N_18008,N_12689,N_13817);
and U18009 (N_18009,N_12889,N_14126);
nor U18010 (N_18010,N_12312,N_12035);
nand U18011 (N_18011,N_12466,N_13193);
nand U18012 (N_18012,N_12269,N_11826);
nor U18013 (N_18013,N_14045,N_12259);
and U18014 (N_18014,N_10950,N_10029);
nor U18015 (N_18015,N_14826,N_14137);
nor U18016 (N_18016,N_13595,N_14326);
nor U18017 (N_18017,N_13174,N_14974);
or U18018 (N_18018,N_10358,N_10366);
and U18019 (N_18019,N_12180,N_12746);
and U18020 (N_18020,N_11357,N_11033);
or U18021 (N_18021,N_12815,N_14498);
nand U18022 (N_18022,N_13414,N_14706);
nor U18023 (N_18023,N_12456,N_14626);
and U18024 (N_18024,N_12971,N_14567);
nor U18025 (N_18025,N_13125,N_11221);
and U18026 (N_18026,N_12446,N_14753);
nor U18027 (N_18027,N_11361,N_13320);
or U18028 (N_18028,N_11606,N_14504);
nand U18029 (N_18029,N_11859,N_14985);
and U18030 (N_18030,N_11338,N_10363);
nor U18031 (N_18031,N_14313,N_14401);
and U18032 (N_18032,N_11569,N_11698);
and U18033 (N_18033,N_14292,N_10107);
nand U18034 (N_18034,N_14573,N_10529);
nor U18035 (N_18035,N_10551,N_10160);
nand U18036 (N_18036,N_14911,N_10574);
and U18037 (N_18037,N_13555,N_14322);
or U18038 (N_18038,N_11802,N_11277);
and U18039 (N_18039,N_12257,N_14473);
or U18040 (N_18040,N_11440,N_12700);
or U18041 (N_18041,N_11527,N_10439);
or U18042 (N_18042,N_12747,N_10408);
and U18043 (N_18043,N_13162,N_11031);
nor U18044 (N_18044,N_12754,N_10060);
nor U18045 (N_18045,N_11830,N_14916);
or U18046 (N_18046,N_11745,N_12562);
nor U18047 (N_18047,N_10432,N_10235);
nor U18048 (N_18048,N_12323,N_13628);
and U18049 (N_18049,N_12329,N_14008);
or U18050 (N_18050,N_14344,N_13182);
or U18051 (N_18051,N_13893,N_13990);
or U18052 (N_18052,N_14790,N_10816);
nor U18053 (N_18053,N_11970,N_14206);
nand U18054 (N_18054,N_11550,N_14919);
or U18055 (N_18055,N_10996,N_13269);
nor U18056 (N_18056,N_10403,N_11945);
nor U18057 (N_18057,N_12950,N_14703);
and U18058 (N_18058,N_11560,N_12918);
and U18059 (N_18059,N_14586,N_11393);
nand U18060 (N_18060,N_10279,N_13914);
and U18061 (N_18061,N_11508,N_12954);
nor U18062 (N_18062,N_11971,N_13064);
or U18063 (N_18063,N_13075,N_10502);
or U18064 (N_18064,N_14585,N_13581);
and U18065 (N_18065,N_14300,N_13999);
or U18066 (N_18066,N_14074,N_12181);
nor U18067 (N_18067,N_12839,N_13954);
nand U18068 (N_18068,N_13429,N_11182);
nand U18069 (N_18069,N_12682,N_14217);
nand U18070 (N_18070,N_10096,N_11286);
nor U18071 (N_18071,N_10950,N_12288);
and U18072 (N_18072,N_12517,N_13338);
and U18073 (N_18073,N_11279,N_12215);
nand U18074 (N_18074,N_14691,N_14567);
nand U18075 (N_18075,N_11786,N_12190);
nor U18076 (N_18076,N_12535,N_10658);
and U18077 (N_18077,N_10119,N_13421);
or U18078 (N_18078,N_14078,N_13234);
nor U18079 (N_18079,N_12380,N_11517);
nand U18080 (N_18080,N_11897,N_10695);
nand U18081 (N_18081,N_11772,N_14339);
nor U18082 (N_18082,N_10070,N_13521);
nand U18083 (N_18083,N_11770,N_10452);
nand U18084 (N_18084,N_10546,N_10865);
nor U18085 (N_18085,N_11762,N_12540);
nand U18086 (N_18086,N_13678,N_13412);
xor U18087 (N_18087,N_13767,N_12429);
and U18088 (N_18088,N_12816,N_11566);
nor U18089 (N_18089,N_12245,N_10152);
nand U18090 (N_18090,N_12298,N_10335);
nor U18091 (N_18091,N_13084,N_12345);
or U18092 (N_18092,N_10966,N_11951);
and U18093 (N_18093,N_10263,N_13944);
and U18094 (N_18094,N_13559,N_14217);
and U18095 (N_18095,N_10110,N_12682);
or U18096 (N_18096,N_10798,N_10545);
nor U18097 (N_18097,N_13650,N_12801);
or U18098 (N_18098,N_11643,N_11186);
and U18099 (N_18099,N_13379,N_13046);
and U18100 (N_18100,N_13994,N_11767);
nor U18101 (N_18101,N_10303,N_10203);
or U18102 (N_18102,N_11303,N_12888);
nand U18103 (N_18103,N_14878,N_14389);
nor U18104 (N_18104,N_11375,N_10203);
nand U18105 (N_18105,N_11759,N_10693);
nand U18106 (N_18106,N_11948,N_12173);
nand U18107 (N_18107,N_13466,N_10853);
and U18108 (N_18108,N_14537,N_11694);
and U18109 (N_18109,N_13902,N_14689);
or U18110 (N_18110,N_13337,N_13344);
nor U18111 (N_18111,N_10884,N_12145);
and U18112 (N_18112,N_10129,N_14627);
nand U18113 (N_18113,N_13502,N_10586);
nor U18114 (N_18114,N_14650,N_14731);
or U18115 (N_18115,N_11713,N_12512);
or U18116 (N_18116,N_10659,N_14118);
nor U18117 (N_18117,N_11896,N_12209);
or U18118 (N_18118,N_11144,N_14485);
nor U18119 (N_18119,N_11704,N_10990);
nand U18120 (N_18120,N_12748,N_14757);
nor U18121 (N_18121,N_11226,N_12722);
and U18122 (N_18122,N_13920,N_10784);
nand U18123 (N_18123,N_11596,N_10076);
or U18124 (N_18124,N_13878,N_12575);
nand U18125 (N_18125,N_11272,N_13900);
nor U18126 (N_18126,N_11022,N_10092);
and U18127 (N_18127,N_13364,N_10241);
or U18128 (N_18128,N_13750,N_11286);
or U18129 (N_18129,N_10921,N_10073);
and U18130 (N_18130,N_14302,N_12265);
and U18131 (N_18131,N_10553,N_13566);
nor U18132 (N_18132,N_11750,N_14144);
nand U18133 (N_18133,N_12616,N_10596);
nor U18134 (N_18134,N_13436,N_11588);
or U18135 (N_18135,N_12775,N_10153);
nor U18136 (N_18136,N_11080,N_10358);
or U18137 (N_18137,N_11014,N_11885);
or U18138 (N_18138,N_13344,N_13305);
and U18139 (N_18139,N_10372,N_14973);
nand U18140 (N_18140,N_13110,N_12894);
and U18141 (N_18141,N_13739,N_11056);
nor U18142 (N_18142,N_14698,N_12072);
and U18143 (N_18143,N_10746,N_14070);
nand U18144 (N_18144,N_13062,N_14471);
or U18145 (N_18145,N_14502,N_13329);
nand U18146 (N_18146,N_13863,N_11162);
and U18147 (N_18147,N_12315,N_10141);
nor U18148 (N_18148,N_11210,N_12413);
nand U18149 (N_18149,N_11262,N_14721);
and U18150 (N_18150,N_12761,N_12843);
and U18151 (N_18151,N_11043,N_13411);
and U18152 (N_18152,N_11601,N_14394);
or U18153 (N_18153,N_12891,N_11827);
nand U18154 (N_18154,N_11479,N_13804);
or U18155 (N_18155,N_11376,N_10052);
nand U18156 (N_18156,N_11414,N_14088);
nand U18157 (N_18157,N_13587,N_10520);
or U18158 (N_18158,N_14241,N_13263);
nand U18159 (N_18159,N_13254,N_10609);
or U18160 (N_18160,N_10024,N_11405);
nor U18161 (N_18161,N_12778,N_14348);
nand U18162 (N_18162,N_12497,N_11193);
nor U18163 (N_18163,N_10515,N_12509);
nor U18164 (N_18164,N_11723,N_10888);
nor U18165 (N_18165,N_11414,N_14924);
nand U18166 (N_18166,N_14774,N_14443);
or U18167 (N_18167,N_11859,N_10256);
and U18168 (N_18168,N_14641,N_13211);
and U18169 (N_18169,N_12180,N_13063);
or U18170 (N_18170,N_12084,N_12613);
nand U18171 (N_18171,N_13581,N_12126);
nand U18172 (N_18172,N_12405,N_14081);
and U18173 (N_18173,N_12668,N_11393);
and U18174 (N_18174,N_10108,N_13712);
or U18175 (N_18175,N_10514,N_14968);
and U18176 (N_18176,N_11327,N_12889);
or U18177 (N_18177,N_12327,N_14153);
nor U18178 (N_18178,N_11810,N_10620);
or U18179 (N_18179,N_14900,N_10221);
nor U18180 (N_18180,N_10655,N_13523);
and U18181 (N_18181,N_13822,N_11332);
nand U18182 (N_18182,N_10824,N_14792);
and U18183 (N_18183,N_13959,N_13723);
nand U18184 (N_18184,N_13962,N_14405);
nor U18185 (N_18185,N_12597,N_10402);
and U18186 (N_18186,N_14497,N_13337);
nand U18187 (N_18187,N_13950,N_14471);
and U18188 (N_18188,N_13624,N_10848);
or U18189 (N_18189,N_10533,N_10986);
nor U18190 (N_18190,N_13107,N_12288);
and U18191 (N_18191,N_11078,N_14205);
and U18192 (N_18192,N_10366,N_10651);
or U18193 (N_18193,N_14997,N_11695);
nand U18194 (N_18194,N_10314,N_13125);
nand U18195 (N_18195,N_12589,N_14972);
nand U18196 (N_18196,N_10199,N_12897);
nor U18197 (N_18197,N_10570,N_10417);
or U18198 (N_18198,N_14216,N_14564);
nand U18199 (N_18199,N_14679,N_10488);
or U18200 (N_18200,N_10562,N_13706);
nor U18201 (N_18201,N_12058,N_14953);
nor U18202 (N_18202,N_13256,N_13370);
nor U18203 (N_18203,N_11317,N_10216);
or U18204 (N_18204,N_11670,N_14256);
nand U18205 (N_18205,N_13653,N_12357);
nor U18206 (N_18206,N_13168,N_10282);
xor U18207 (N_18207,N_11168,N_11065);
or U18208 (N_18208,N_11235,N_10044);
nand U18209 (N_18209,N_13323,N_11285);
or U18210 (N_18210,N_13537,N_13761);
and U18211 (N_18211,N_11258,N_11361);
and U18212 (N_18212,N_14810,N_10427);
or U18213 (N_18213,N_14492,N_10610);
and U18214 (N_18214,N_11448,N_12900);
nand U18215 (N_18215,N_13277,N_11562);
nand U18216 (N_18216,N_12485,N_13416);
and U18217 (N_18217,N_13095,N_14091);
or U18218 (N_18218,N_10321,N_11418);
or U18219 (N_18219,N_12087,N_10435);
nor U18220 (N_18220,N_14809,N_14721);
nor U18221 (N_18221,N_14218,N_10559);
nor U18222 (N_18222,N_13603,N_14610);
nand U18223 (N_18223,N_12397,N_12863);
nand U18224 (N_18224,N_14344,N_10312);
nand U18225 (N_18225,N_14362,N_13910);
nand U18226 (N_18226,N_13110,N_14924);
and U18227 (N_18227,N_10192,N_12794);
nor U18228 (N_18228,N_12166,N_14345);
xor U18229 (N_18229,N_14513,N_12052);
or U18230 (N_18230,N_13428,N_11522);
nand U18231 (N_18231,N_14761,N_13310);
nand U18232 (N_18232,N_13981,N_12402);
nand U18233 (N_18233,N_13928,N_12852);
and U18234 (N_18234,N_11323,N_11777);
nor U18235 (N_18235,N_14074,N_11026);
or U18236 (N_18236,N_14985,N_10792);
and U18237 (N_18237,N_10158,N_14042);
nor U18238 (N_18238,N_12589,N_13826);
nor U18239 (N_18239,N_14642,N_13379);
nand U18240 (N_18240,N_10917,N_11874);
nand U18241 (N_18241,N_14080,N_11785);
and U18242 (N_18242,N_11672,N_14692);
nand U18243 (N_18243,N_10392,N_11508);
or U18244 (N_18244,N_12453,N_10308);
nand U18245 (N_18245,N_14546,N_12134);
nand U18246 (N_18246,N_14016,N_12613);
nand U18247 (N_18247,N_14621,N_10809);
and U18248 (N_18248,N_14579,N_11876);
or U18249 (N_18249,N_12360,N_14252);
nor U18250 (N_18250,N_12121,N_11395);
nand U18251 (N_18251,N_11746,N_12083);
nand U18252 (N_18252,N_11225,N_13168);
or U18253 (N_18253,N_12365,N_11103);
nor U18254 (N_18254,N_10610,N_11599);
and U18255 (N_18255,N_12464,N_12814);
nand U18256 (N_18256,N_10542,N_14624);
and U18257 (N_18257,N_10497,N_13110);
nor U18258 (N_18258,N_12559,N_11106);
and U18259 (N_18259,N_13824,N_13021);
and U18260 (N_18260,N_12808,N_12587);
nor U18261 (N_18261,N_14772,N_10302);
nand U18262 (N_18262,N_13055,N_11202);
nand U18263 (N_18263,N_14256,N_13059);
or U18264 (N_18264,N_13719,N_14887);
and U18265 (N_18265,N_11436,N_12565);
nand U18266 (N_18266,N_12189,N_10723);
and U18267 (N_18267,N_12749,N_12244);
nand U18268 (N_18268,N_14603,N_12562);
nand U18269 (N_18269,N_14851,N_10886);
and U18270 (N_18270,N_11730,N_10994);
nand U18271 (N_18271,N_14867,N_14311);
or U18272 (N_18272,N_13833,N_14294);
or U18273 (N_18273,N_10512,N_10764);
nor U18274 (N_18274,N_13544,N_10705);
nand U18275 (N_18275,N_11719,N_11779);
or U18276 (N_18276,N_10654,N_11066);
and U18277 (N_18277,N_10785,N_13207);
and U18278 (N_18278,N_11932,N_12779);
and U18279 (N_18279,N_10288,N_14999);
nand U18280 (N_18280,N_13757,N_12451);
nand U18281 (N_18281,N_10159,N_13285);
or U18282 (N_18282,N_14173,N_11456);
or U18283 (N_18283,N_13652,N_13421);
and U18284 (N_18284,N_12175,N_12034);
nand U18285 (N_18285,N_13459,N_14551);
or U18286 (N_18286,N_12172,N_14044);
nand U18287 (N_18287,N_14711,N_10193);
nand U18288 (N_18288,N_10081,N_10488);
or U18289 (N_18289,N_11056,N_12947);
and U18290 (N_18290,N_11339,N_14528);
and U18291 (N_18291,N_10994,N_12096);
nand U18292 (N_18292,N_10110,N_13797);
nor U18293 (N_18293,N_10982,N_12150);
nor U18294 (N_18294,N_11140,N_14406);
nand U18295 (N_18295,N_11286,N_10086);
and U18296 (N_18296,N_12330,N_12778);
nand U18297 (N_18297,N_13359,N_11671);
nand U18298 (N_18298,N_12773,N_11280);
nor U18299 (N_18299,N_11683,N_10999);
or U18300 (N_18300,N_13553,N_13550);
nor U18301 (N_18301,N_13649,N_11036);
nand U18302 (N_18302,N_10147,N_12550);
nor U18303 (N_18303,N_12889,N_14828);
or U18304 (N_18304,N_14888,N_10430);
or U18305 (N_18305,N_14911,N_11792);
nor U18306 (N_18306,N_12540,N_12521);
nor U18307 (N_18307,N_10883,N_11136);
or U18308 (N_18308,N_13277,N_14316);
nand U18309 (N_18309,N_13995,N_11364);
and U18310 (N_18310,N_11254,N_14881);
nor U18311 (N_18311,N_11092,N_13704);
or U18312 (N_18312,N_13932,N_10113);
and U18313 (N_18313,N_14163,N_11650);
nor U18314 (N_18314,N_13959,N_14878);
and U18315 (N_18315,N_12722,N_14777);
nand U18316 (N_18316,N_11303,N_10326);
and U18317 (N_18317,N_12781,N_14068);
nand U18318 (N_18318,N_10732,N_12764);
and U18319 (N_18319,N_14708,N_10323);
and U18320 (N_18320,N_10359,N_12517);
nand U18321 (N_18321,N_12179,N_14875);
nand U18322 (N_18322,N_13211,N_10473);
or U18323 (N_18323,N_14829,N_14965);
or U18324 (N_18324,N_12943,N_11869);
nand U18325 (N_18325,N_14947,N_13465);
or U18326 (N_18326,N_14083,N_10303);
and U18327 (N_18327,N_12209,N_14882);
nor U18328 (N_18328,N_11845,N_11847);
nand U18329 (N_18329,N_13515,N_10474);
or U18330 (N_18330,N_13686,N_11573);
or U18331 (N_18331,N_12710,N_14561);
and U18332 (N_18332,N_11079,N_14260);
nor U18333 (N_18333,N_14734,N_11723);
nand U18334 (N_18334,N_13032,N_10191);
and U18335 (N_18335,N_14087,N_13984);
and U18336 (N_18336,N_10068,N_10771);
nand U18337 (N_18337,N_12072,N_11408);
or U18338 (N_18338,N_12861,N_13437);
or U18339 (N_18339,N_10395,N_13627);
nand U18340 (N_18340,N_14852,N_13928);
or U18341 (N_18341,N_11106,N_12951);
nand U18342 (N_18342,N_14453,N_13347);
nor U18343 (N_18343,N_11015,N_14467);
and U18344 (N_18344,N_14705,N_14618);
and U18345 (N_18345,N_11263,N_13551);
nor U18346 (N_18346,N_13655,N_12005);
nor U18347 (N_18347,N_11092,N_14741);
and U18348 (N_18348,N_12760,N_10039);
nand U18349 (N_18349,N_11725,N_14260);
nand U18350 (N_18350,N_10147,N_14521);
or U18351 (N_18351,N_10794,N_14331);
nand U18352 (N_18352,N_10954,N_14621);
nor U18353 (N_18353,N_11184,N_13041);
nor U18354 (N_18354,N_11892,N_10334);
and U18355 (N_18355,N_10470,N_12554);
nand U18356 (N_18356,N_12232,N_11838);
and U18357 (N_18357,N_14093,N_10607);
and U18358 (N_18358,N_12594,N_10481);
nor U18359 (N_18359,N_13940,N_12273);
nor U18360 (N_18360,N_14206,N_14093);
or U18361 (N_18361,N_11414,N_10597);
or U18362 (N_18362,N_12942,N_14977);
nor U18363 (N_18363,N_11141,N_12394);
nand U18364 (N_18364,N_10472,N_13744);
nand U18365 (N_18365,N_12909,N_14865);
nand U18366 (N_18366,N_10713,N_10939);
and U18367 (N_18367,N_11926,N_10190);
and U18368 (N_18368,N_11281,N_11596);
or U18369 (N_18369,N_12908,N_11233);
and U18370 (N_18370,N_10886,N_12768);
nor U18371 (N_18371,N_11063,N_12004);
nor U18372 (N_18372,N_11911,N_13278);
or U18373 (N_18373,N_10536,N_13546);
or U18374 (N_18374,N_14614,N_12715);
and U18375 (N_18375,N_10181,N_14753);
and U18376 (N_18376,N_10116,N_13271);
or U18377 (N_18377,N_10755,N_11747);
nor U18378 (N_18378,N_12789,N_14927);
and U18379 (N_18379,N_13629,N_10686);
or U18380 (N_18380,N_12269,N_13741);
or U18381 (N_18381,N_12297,N_11440);
nand U18382 (N_18382,N_11803,N_12128);
and U18383 (N_18383,N_11095,N_11739);
nand U18384 (N_18384,N_11186,N_13522);
nor U18385 (N_18385,N_13248,N_11507);
or U18386 (N_18386,N_14603,N_14763);
and U18387 (N_18387,N_14659,N_10063);
xnor U18388 (N_18388,N_14681,N_11545);
or U18389 (N_18389,N_12889,N_14306);
nor U18390 (N_18390,N_10228,N_10483);
nand U18391 (N_18391,N_11906,N_12211);
xnor U18392 (N_18392,N_11131,N_10770);
and U18393 (N_18393,N_13066,N_13117);
nand U18394 (N_18394,N_11791,N_11204);
nor U18395 (N_18395,N_11044,N_10539);
or U18396 (N_18396,N_10376,N_10135);
and U18397 (N_18397,N_13983,N_12142);
and U18398 (N_18398,N_12057,N_14488);
nand U18399 (N_18399,N_14485,N_12635);
or U18400 (N_18400,N_13143,N_10187);
or U18401 (N_18401,N_14304,N_14791);
nand U18402 (N_18402,N_12804,N_11865);
or U18403 (N_18403,N_10838,N_11680);
xor U18404 (N_18404,N_14146,N_14502);
xnor U18405 (N_18405,N_14306,N_12139);
nand U18406 (N_18406,N_14869,N_12886);
or U18407 (N_18407,N_12989,N_10330);
and U18408 (N_18408,N_10887,N_11515);
or U18409 (N_18409,N_14764,N_14251);
xnor U18410 (N_18410,N_14926,N_14097);
nor U18411 (N_18411,N_10220,N_14661);
or U18412 (N_18412,N_12925,N_13474);
and U18413 (N_18413,N_14189,N_10116);
and U18414 (N_18414,N_13559,N_13057);
nand U18415 (N_18415,N_14287,N_13587);
nor U18416 (N_18416,N_11772,N_10298);
nand U18417 (N_18417,N_14205,N_11070);
and U18418 (N_18418,N_12407,N_13539);
or U18419 (N_18419,N_13397,N_12915);
or U18420 (N_18420,N_12584,N_14769);
and U18421 (N_18421,N_11165,N_11503);
nor U18422 (N_18422,N_10827,N_11351);
nand U18423 (N_18423,N_12437,N_10412);
and U18424 (N_18424,N_10114,N_10573);
nor U18425 (N_18425,N_13907,N_10135);
and U18426 (N_18426,N_13442,N_10445);
or U18427 (N_18427,N_13993,N_11921);
and U18428 (N_18428,N_14370,N_14237);
and U18429 (N_18429,N_11815,N_14419);
and U18430 (N_18430,N_10921,N_13733);
or U18431 (N_18431,N_11637,N_10643);
nand U18432 (N_18432,N_14666,N_11485);
or U18433 (N_18433,N_10282,N_13133);
or U18434 (N_18434,N_11613,N_11304);
nor U18435 (N_18435,N_12478,N_12805);
nand U18436 (N_18436,N_14969,N_14298);
nor U18437 (N_18437,N_11594,N_13436);
and U18438 (N_18438,N_10466,N_11263);
nand U18439 (N_18439,N_12118,N_14086);
and U18440 (N_18440,N_12996,N_11139);
nand U18441 (N_18441,N_14429,N_14257);
nand U18442 (N_18442,N_11444,N_13578);
or U18443 (N_18443,N_13065,N_14639);
nand U18444 (N_18444,N_12834,N_13195);
and U18445 (N_18445,N_14546,N_10245);
nand U18446 (N_18446,N_11255,N_11249);
and U18447 (N_18447,N_10376,N_14855);
nor U18448 (N_18448,N_14374,N_12789);
or U18449 (N_18449,N_14155,N_13151);
nor U18450 (N_18450,N_14409,N_12293);
or U18451 (N_18451,N_13789,N_13060);
nor U18452 (N_18452,N_10095,N_13651);
nor U18453 (N_18453,N_13597,N_12246);
and U18454 (N_18454,N_14146,N_13237);
nor U18455 (N_18455,N_14391,N_14003);
nor U18456 (N_18456,N_12469,N_11419);
nand U18457 (N_18457,N_10292,N_14561);
nor U18458 (N_18458,N_11518,N_10480);
and U18459 (N_18459,N_11147,N_13235);
nor U18460 (N_18460,N_12285,N_14489);
nor U18461 (N_18461,N_11923,N_10459);
or U18462 (N_18462,N_14542,N_12976);
nand U18463 (N_18463,N_14278,N_10486);
nand U18464 (N_18464,N_11159,N_11061);
or U18465 (N_18465,N_10613,N_13812);
or U18466 (N_18466,N_12597,N_13534);
nor U18467 (N_18467,N_12406,N_12668);
and U18468 (N_18468,N_11351,N_13800);
and U18469 (N_18469,N_10205,N_12608);
or U18470 (N_18470,N_13700,N_12390);
nor U18471 (N_18471,N_14035,N_12656);
or U18472 (N_18472,N_12946,N_12638);
nor U18473 (N_18473,N_12057,N_13245);
or U18474 (N_18474,N_11926,N_14883);
or U18475 (N_18475,N_11793,N_14684);
nor U18476 (N_18476,N_10290,N_13285);
or U18477 (N_18477,N_14196,N_14023);
nand U18478 (N_18478,N_13314,N_10271);
and U18479 (N_18479,N_10129,N_11774);
and U18480 (N_18480,N_10795,N_12648);
or U18481 (N_18481,N_12245,N_10459);
and U18482 (N_18482,N_10552,N_14365);
or U18483 (N_18483,N_14472,N_12532);
xnor U18484 (N_18484,N_10247,N_11252);
and U18485 (N_18485,N_14845,N_14201);
and U18486 (N_18486,N_11747,N_13382);
nand U18487 (N_18487,N_10442,N_13153);
nor U18488 (N_18488,N_12783,N_11438);
or U18489 (N_18489,N_12444,N_12635);
nor U18490 (N_18490,N_11135,N_14709);
nor U18491 (N_18491,N_14411,N_10227);
and U18492 (N_18492,N_11104,N_11703);
nand U18493 (N_18493,N_12539,N_13795);
or U18494 (N_18494,N_12605,N_12345);
nand U18495 (N_18495,N_13134,N_10295);
nand U18496 (N_18496,N_12650,N_14301);
nor U18497 (N_18497,N_11636,N_13645);
nor U18498 (N_18498,N_13780,N_10014);
nor U18499 (N_18499,N_11826,N_11421);
nand U18500 (N_18500,N_14521,N_13994);
or U18501 (N_18501,N_13908,N_11464);
nor U18502 (N_18502,N_13481,N_11562);
and U18503 (N_18503,N_11193,N_14249);
and U18504 (N_18504,N_10927,N_11109);
nor U18505 (N_18505,N_14125,N_10545);
nor U18506 (N_18506,N_12544,N_10144);
and U18507 (N_18507,N_11937,N_14913);
or U18508 (N_18508,N_14525,N_12701);
or U18509 (N_18509,N_14933,N_11037);
nand U18510 (N_18510,N_13882,N_11119);
nand U18511 (N_18511,N_12949,N_11651);
nand U18512 (N_18512,N_12572,N_13650);
or U18513 (N_18513,N_10155,N_12360);
and U18514 (N_18514,N_10135,N_10276);
nor U18515 (N_18515,N_12153,N_14034);
nand U18516 (N_18516,N_10707,N_12312);
nor U18517 (N_18517,N_12199,N_11497);
or U18518 (N_18518,N_11512,N_14437);
or U18519 (N_18519,N_11501,N_10045);
or U18520 (N_18520,N_14054,N_13394);
and U18521 (N_18521,N_13513,N_11215);
nor U18522 (N_18522,N_12663,N_10679);
or U18523 (N_18523,N_10857,N_12841);
nand U18524 (N_18524,N_14638,N_14490);
nor U18525 (N_18525,N_14336,N_11357);
nand U18526 (N_18526,N_13240,N_12931);
or U18527 (N_18527,N_11371,N_10958);
or U18528 (N_18528,N_10843,N_13242);
nor U18529 (N_18529,N_11313,N_12963);
and U18530 (N_18530,N_13354,N_14851);
nor U18531 (N_18531,N_12691,N_12150);
xor U18532 (N_18532,N_11567,N_10311);
nor U18533 (N_18533,N_10074,N_11958);
or U18534 (N_18534,N_10554,N_14049);
nand U18535 (N_18535,N_10204,N_12017);
nor U18536 (N_18536,N_11703,N_11565);
or U18537 (N_18537,N_11578,N_13710);
and U18538 (N_18538,N_14298,N_12989);
or U18539 (N_18539,N_11792,N_10924);
nand U18540 (N_18540,N_12695,N_11136);
nor U18541 (N_18541,N_12140,N_14249);
or U18542 (N_18542,N_12955,N_11799);
nor U18543 (N_18543,N_14309,N_11124);
or U18544 (N_18544,N_11592,N_11736);
nor U18545 (N_18545,N_11368,N_12999);
nor U18546 (N_18546,N_12985,N_13721);
and U18547 (N_18547,N_13671,N_14392);
nor U18548 (N_18548,N_11426,N_13768);
or U18549 (N_18549,N_14993,N_12181);
and U18550 (N_18550,N_13957,N_13741);
and U18551 (N_18551,N_10668,N_12562);
nand U18552 (N_18552,N_11141,N_10984);
nand U18553 (N_18553,N_11648,N_13372);
or U18554 (N_18554,N_13268,N_13299);
nor U18555 (N_18555,N_11844,N_13735);
and U18556 (N_18556,N_13740,N_11113);
and U18557 (N_18557,N_11946,N_13323);
nor U18558 (N_18558,N_11223,N_10459);
nor U18559 (N_18559,N_10936,N_10307);
nand U18560 (N_18560,N_14212,N_12299);
or U18561 (N_18561,N_12820,N_12082);
or U18562 (N_18562,N_11635,N_14070);
nor U18563 (N_18563,N_12095,N_13586);
nor U18564 (N_18564,N_13898,N_11106);
and U18565 (N_18565,N_10324,N_12372);
or U18566 (N_18566,N_13549,N_14288);
or U18567 (N_18567,N_14302,N_12050);
nor U18568 (N_18568,N_11044,N_10451);
nand U18569 (N_18569,N_13762,N_11784);
and U18570 (N_18570,N_13685,N_13959);
nor U18571 (N_18571,N_11011,N_12733);
nor U18572 (N_18572,N_13939,N_14441);
nor U18573 (N_18573,N_10172,N_12827);
and U18574 (N_18574,N_10800,N_13061);
and U18575 (N_18575,N_10644,N_13868);
nand U18576 (N_18576,N_11173,N_13144);
nand U18577 (N_18577,N_12889,N_11959);
nor U18578 (N_18578,N_14345,N_11511);
and U18579 (N_18579,N_12909,N_11722);
or U18580 (N_18580,N_14571,N_14106);
nand U18581 (N_18581,N_10218,N_10422);
nand U18582 (N_18582,N_11028,N_12912);
and U18583 (N_18583,N_13194,N_14938);
and U18584 (N_18584,N_14679,N_13518);
nor U18585 (N_18585,N_11047,N_12167);
nand U18586 (N_18586,N_10223,N_11442);
nand U18587 (N_18587,N_11890,N_10978);
or U18588 (N_18588,N_14118,N_11061);
nor U18589 (N_18589,N_14830,N_13830);
or U18590 (N_18590,N_13290,N_14782);
and U18591 (N_18591,N_13139,N_14206);
or U18592 (N_18592,N_11687,N_13930);
nand U18593 (N_18593,N_13755,N_12401);
or U18594 (N_18594,N_11241,N_14342);
nand U18595 (N_18595,N_11470,N_11720);
nand U18596 (N_18596,N_11653,N_14993);
or U18597 (N_18597,N_11518,N_13717);
or U18598 (N_18598,N_13059,N_11743);
nand U18599 (N_18599,N_13879,N_10625);
or U18600 (N_18600,N_12002,N_12509);
nor U18601 (N_18601,N_14029,N_13854);
and U18602 (N_18602,N_10573,N_12310);
or U18603 (N_18603,N_12172,N_11868);
nor U18604 (N_18604,N_10040,N_11598);
xor U18605 (N_18605,N_13409,N_11593);
nor U18606 (N_18606,N_12728,N_12142);
or U18607 (N_18607,N_11704,N_13458);
and U18608 (N_18608,N_13980,N_12598);
or U18609 (N_18609,N_12733,N_12816);
nor U18610 (N_18610,N_14853,N_13428);
nor U18611 (N_18611,N_14882,N_14139);
nor U18612 (N_18612,N_11471,N_14309);
nor U18613 (N_18613,N_14230,N_11512);
nand U18614 (N_18614,N_11715,N_13170);
nand U18615 (N_18615,N_11628,N_13303);
nor U18616 (N_18616,N_14534,N_11093);
or U18617 (N_18617,N_10546,N_12037);
nor U18618 (N_18618,N_12581,N_12689);
nand U18619 (N_18619,N_10428,N_14181);
and U18620 (N_18620,N_12366,N_11105);
nor U18621 (N_18621,N_14879,N_10655);
nand U18622 (N_18622,N_11546,N_13888);
and U18623 (N_18623,N_13503,N_11900);
nor U18624 (N_18624,N_13570,N_12663);
nand U18625 (N_18625,N_14599,N_13868);
or U18626 (N_18626,N_13334,N_10508);
nor U18627 (N_18627,N_13211,N_11507);
nor U18628 (N_18628,N_10869,N_14353);
or U18629 (N_18629,N_11832,N_11452);
nor U18630 (N_18630,N_13257,N_12065);
nor U18631 (N_18631,N_12349,N_14793);
or U18632 (N_18632,N_11526,N_11233);
and U18633 (N_18633,N_13825,N_10140);
or U18634 (N_18634,N_10923,N_10126);
and U18635 (N_18635,N_10513,N_10580);
and U18636 (N_18636,N_14410,N_13234);
or U18637 (N_18637,N_11179,N_11485);
or U18638 (N_18638,N_12635,N_14073);
or U18639 (N_18639,N_12403,N_13432);
or U18640 (N_18640,N_13049,N_14519);
nand U18641 (N_18641,N_13909,N_10185);
or U18642 (N_18642,N_12300,N_12445);
nand U18643 (N_18643,N_13316,N_14598);
nor U18644 (N_18644,N_10125,N_14233);
nor U18645 (N_18645,N_14521,N_11677);
or U18646 (N_18646,N_11212,N_11667);
nor U18647 (N_18647,N_14672,N_10265);
and U18648 (N_18648,N_13788,N_11075);
or U18649 (N_18649,N_11821,N_11647);
and U18650 (N_18650,N_13962,N_10410);
nor U18651 (N_18651,N_14934,N_11275);
nor U18652 (N_18652,N_10613,N_14807);
or U18653 (N_18653,N_13074,N_11068);
nor U18654 (N_18654,N_11590,N_12124);
or U18655 (N_18655,N_13184,N_14561);
nor U18656 (N_18656,N_11408,N_11395);
nor U18657 (N_18657,N_11119,N_10311);
nand U18658 (N_18658,N_13005,N_11614);
nand U18659 (N_18659,N_11541,N_13283);
or U18660 (N_18660,N_12128,N_11831);
or U18661 (N_18661,N_13150,N_13905);
nand U18662 (N_18662,N_14921,N_13770);
nor U18663 (N_18663,N_14411,N_10616);
and U18664 (N_18664,N_12713,N_11682);
nor U18665 (N_18665,N_14050,N_11582);
and U18666 (N_18666,N_12239,N_11820);
and U18667 (N_18667,N_13468,N_11468);
or U18668 (N_18668,N_14478,N_11537);
and U18669 (N_18669,N_12012,N_12011);
nor U18670 (N_18670,N_13745,N_13422);
or U18671 (N_18671,N_14535,N_14250);
nor U18672 (N_18672,N_14465,N_12123);
nand U18673 (N_18673,N_12548,N_11575);
nor U18674 (N_18674,N_12610,N_12989);
nand U18675 (N_18675,N_14111,N_12255);
xor U18676 (N_18676,N_12558,N_13819);
or U18677 (N_18677,N_10007,N_11633);
and U18678 (N_18678,N_12687,N_14993);
and U18679 (N_18679,N_14465,N_10587);
nand U18680 (N_18680,N_10795,N_13655);
xnor U18681 (N_18681,N_12122,N_14078);
nor U18682 (N_18682,N_11395,N_13747);
nand U18683 (N_18683,N_10636,N_12428);
or U18684 (N_18684,N_11443,N_14795);
or U18685 (N_18685,N_12507,N_12655);
nor U18686 (N_18686,N_10445,N_14470);
and U18687 (N_18687,N_11061,N_13333);
nor U18688 (N_18688,N_11567,N_12018);
nor U18689 (N_18689,N_14233,N_12544);
and U18690 (N_18690,N_10978,N_10291);
nor U18691 (N_18691,N_11801,N_10532);
and U18692 (N_18692,N_13462,N_10223);
nand U18693 (N_18693,N_13863,N_11550);
and U18694 (N_18694,N_10730,N_10788);
nor U18695 (N_18695,N_12901,N_11211);
nor U18696 (N_18696,N_14261,N_13686);
or U18697 (N_18697,N_11522,N_14886);
nor U18698 (N_18698,N_12139,N_11486);
nand U18699 (N_18699,N_11284,N_13217);
and U18700 (N_18700,N_12010,N_10795);
and U18701 (N_18701,N_10227,N_10927);
and U18702 (N_18702,N_13420,N_13981);
or U18703 (N_18703,N_12843,N_12393);
or U18704 (N_18704,N_13572,N_11140);
and U18705 (N_18705,N_13630,N_13803);
or U18706 (N_18706,N_13865,N_14590);
nand U18707 (N_18707,N_13291,N_10316);
nand U18708 (N_18708,N_10938,N_14151);
or U18709 (N_18709,N_12504,N_12757);
or U18710 (N_18710,N_11095,N_12305);
and U18711 (N_18711,N_14669,N_10890);
nor U18712 (N_18712,N_12267,N_13531);
nor U18713 (N_18713,N_14948,N_13974);
nor U18714 (N_18714,N_10560,N_10107);
nand U18715 (N_18715,N_14455,N_12762);
nand U18716 (N_18716,N_12986,N_13523);
nand U18717 (N_18717,N_12990,N_11120);
or U18718 (N_18718,N_10283,N_14756);
nand U18719 (N_18719,N_12773,N_12003);
or U18720 (N_18720,N_13607,N_12730);
or U18721 (N_18721,N_14445,N_13851);
nand U18722 (N_18722,N_11424,N_11601);
or U18723 (N_18723,N_12055,N_10880);
nand U18724 (N_18724,N_12071,N_12353);
nor U18725 (N_18725,N_13516,N_10181);
nand U18726 (N_18726,N_11795,N_13409);
nor U18727 (N_18727,N_12061,N_10636);
nor U18728 (N_18728,N_10127,N_11385);
nand U18729 (N_18729,N_14320,N_12097);
or U18730 (N_18730,N_10560,N_13098);
nor U18731 (N_18731,N_12098,N_12161);
xor U18732 (N_18732,N_11603,N_14732);
or U18733 (N_18733,N_14083,N_14629);
nand U18734 (N_18734,N_10892,N_11060);
and U18735 (N_18735,N_11783,N_10951);
and U18736 (N_18736,N_10451,N_14493);
and U18737 (N_18737,N_10747,N_11220);
and U18738 (N_18738,N_12546,N_12138);
nor U18739 (N_18739,N_11523,N_12544);
or U18740 (N_18740,N_11093,N_10863);
nor U18741 (N_18741,N_14915,N_11319);
nand U18742 (N_18742,N_14511,N_14192);
or U18743 (N_18743,N_14629,N_12306);
or U18744 (N_18744,N_11360,N_14578);
nor U18745 (N_18745,N_12998,N_11467);
or U18746 (N_18746,N_12742,N_14240);
xor U18747 (N_18747,N_11163,N_13222);
nand U18748 (N_18748,N_13160,N_13449);
nand U18749 (N_18749,N_13268,N_11360);
nand U18750 (N_18750,N_13344,N_12161);
or U18751 (N_18751,N_10028,N_12789);
nor U18752 (N_18752,N_14740,N_14567);
or U18753 (N_18753,N_11907,N_12689);
nor U18754 (N_18754,N_14422,N_10360);
nand U18755 (N_18755,N_14340,N_12246);
and U18756 (N_18756,N_11504,N_14907);
xor U18757 (N_18757,N_11764,N_11489);
nor U18758 (N_18758,N_13703,N_14084);
and U18759 (N_18759,N_13492,N_10517);
and U18760 (N_18760,N_12199,N_11247);
nand U18761 (N_18761,N_14976,N_13574);
nand U18762 (N_18762,N_13730,N_11292);
or U18763 (N_18763,N_14350,N_14410);
or U18764 (N_18764,N_13210,N_11712);
nand U18765 (N_18765,N_14846,N_13764);
nand U18766 (N_18766,N_14120,N_10364);
nand U18767 (N_18767,N_13071,N_14172);
and U18768 (N_18768,N_12698,N_14307);
nor U18769 (N_18769,N_11166,N_14748);
nor U18770 (N_18770,N_13515,N_10299);
and U18771 (N_18771,N_10917,N_12441);
and U18772 (N_18772,N_11940,N_13098);
nand U18773 (N_18773,N_10652,N_10481);
nand U18774 (N_18774,N_12148,N_12595);
nand U18775 (N_18775,N_14856,N_12624);
nand U18776 (N_18776,N_10017,N_11380);
nand U18777 (N_18777,N_14093,N_10858);
nor U18778 (N_18778,N_14572,N_10078);
nor U18779 (N_18779,N_11943,N_14015);
and U18780 (N_18780,N_10566,N_12386);
nand U18781 (N_18781,N_13038,N_10235);
nand U18782 (N_18782,N_10768,N_12009);
or U18783 (N_18783,N_14641,N_14752);
nand U18784 (N_18784,N_10568,N_10758);
or U18785 (N_18785,N_14085,N_12213);
and U18786 (N_18786,N_14157,N_10205);
and U18787 (N_18787,N_10144,N_10989);
nand U18788 (N_18788,N_13090,N_10619);
nor U18789 (N_18789,N_10904,N_13005);
nor U18790 (N_18790,N_13481,N_13111);
or U18791 (N_18791,N_14662,N_12243);
nand U18792 (N_18792,N_14767,N_11286);
nand U18793 (N_18793,N_13934,N_12265);
nor U18794 (N_18794,N_11194,N_13173);
and U18795 (N_18795,N_11050,N_14600);
nor U18796 (N_18796,N_13606,N_12355);
and U18797 (N_18797,N_14715,N_12473);
nor U18798 (N_18798,N_11906,N_10900);
or U18799 (N_18799,N_11394,N_13154);
or U18800 (N_18800,N_10492,N_14272);
or U18801 (N_18801,N_14552,N_14980);
nand U18802 (N_18802,N_11597,N_13533);
or U18803 (N_18803,N_12964,N_11547);
or U18804 (N_18804,N_13213,N_10175);
or U18805 (N_18805,N_12114,N_10044);
nor U18806 (N_18806,N_13250,N_13589);
and U18807 (N_18807,N_11598,N_12382);
and U18808 (N_18808,N_12758,N_10247);
nand U18809 (N_18809,N_10383,N_12859);
or U18810 (N_18810,N_12269,N_14760);
or U18811 (N_18811,N_13570,N_14374);
nor U18812 (N_18812,N_14926,N_11716);
nor U18813 (N_18813,N_13131,N_13158);
nand U18814 (N_18814,N_10907,N_10824);
or U18815 (N_18815,N_12017,N_13834);
nand U18816 (N_18816,N_12535,N_10631);
and U18817 (N_18817,N_11628,N_10721);
and U18818 (N_18818,N_12388,N_12517);
and U18819 (N_18819,N_11760,N_13411);
or U18820 (N_18820,N_11853,N_11329);
or U18821 (N_18821,N_12086,N_14194);
nand U18822 (N_18822,N_10682,N_10423);
nand U18823 (N_18823,N_13958,N_14468);
and U18824 (N_18824,N_11971,N_13460);
or U18825 (N_18825,N_12149,N_10963);
nor U18826 (N_18826,N_14752,N_11921);
and U18827 (N_18827,N_11639,N_10265);
or U18828 (N_18828,N_14571,N_10614);
and U18829 (N_18829,N_12904,N_11523);
or U18830 (N_18830,N_12650,N_10323);
or U18831 (N_18831,N_10574,N_13887);
or U18832 (N_18832,N_14386,N_14493);
and U18833 (N_18833,N_11300,N_13765);
nor U18834 (N_18834,N_13696,N_14163);
nor U18835 (N_18835,N_11182,N_14642);
and U18836 (N_18836,N_13010,N_14387);
nand U18837 (N_18837,N_11312,N_12930);
and U18838 (N_18838,N_14788,N_11054);
nor U18839 (N_18839,N_10987,N_11360);
nand U18840 (N_18840,N_11715,N_14911);
and U18841 (N_18841,N_13530,N_14211);
or U18842 (N_18842,N_13460,N_14337);
nor U18843 (N_18843,N_13496,N_12381);
or U18844 (N_18844,N_10336,N_10910);
and U18845 (N_18845,N_12203,N_11309);
nor U18846 (N_18846,N_11038,N_14970);
nor U18847 (N_18847,N_11138,N_13862);
nand U18848 (N_18848,N_10658,N_11514);
nor U18849 (N_18849,N_12125,N_14934);
and U18850 (N_18850,N_13306,N_10865);
or U18851 (N_18851,N_14522,N_12106);
nor U18852 (N_18852,N_12340,N_14501);
nor U18853 (N_18853,N_12329,N_12764);
nor U18854 (N_18854,N_10221,N_10504);
nor U18855 (N_18855,N_10009,N_11523);
or U18856 (N_18856,N_14618,N_13163);
nor U18857 (N_18857,N_10801,N_11242);
nand U18858 (N_18858,N_10179,N_10785);
nand U18859 (N_18859,N_10302,N_13724);
nor U18860 (N_18860,N_12603,N_11517);
nor U18861 (N_18861,N_11879,N_10035);
and U18862 (N_18862,N_10013,N_11412);
or U18863 (N_18863,N_13978,N_11374);
nand U18864 (N_18864,N_11110,N_12205);
or U18865 (N_18865,N_10067,N_10991);
or U18866 (N_18866,N_14287,N_13506);
or U18867 (N_18867,N_10085,N_12585);
nor U18868 (N_18868,N_10130,N_13643);
or U18869 (N_18869,N_12869,N_14509);
or U18870 (N_18870,N_13928,N_11283);
nand U18871 (N_18871,N_11368,N_10791);
or U18872 (N_18872,N_12960,N_10203);
nand U18873 (N_18873,N_14290,N_13792);
nand U18874 (N_18874,N_12770,N_14062);
or U18875 (N_18875,N_13023,N_10066);
or U18876 (N_18876,N_13546,N_14341);
nand U18877 (N_18877,N_12651,N_13438);
nor U18878 (N_18878,N_10945,N_10174);
and U18879 (N_18879,N_10802,N_11539);
nand U18880 (N_18880,N_13150,N_10205);
nand U18881 (N_18881,N_13650,N_13166);
nor U18882 (N_18882,N_12275,N_12461);
nor U18883 (N_18883,N_13806,N_14395);
or U18884 (N_18884,N_14769,N_12429);
or U18885 (N_18885,N_11315,N_10798);
or U18886 (N_18886,N_10231,N_13568);
or U18887 (N_18887,N_13687,N_12455);
nor U18888 (N_18888,N_13369,N_10468);
or U18889 (N_18889,N_12232,N_11661);
or U18890 (N_18890,N_12908,N_13903);
or U18891 (N_18891,N_13878,N_14982);
nand U18892 (N_18892,N_11937,N_13785);
nor U18893 (N_18893,N_11636,N_10700);
nor U18894 (N_18894,N_14129,N_12483);
or U18895 (N_18895,N_10747,N_12522);
or U18896 (N_18896,N_13309,N_11823);
or U18897 (N_18897,N_10972,N_14232);
nor U18898 (N_18898,N_13200,N_14137);
nand U18899 (N_18899,N_13806,N_12507);
and U18900 (N_18900,N_13584,N_10850);
or U18901 (N_18901,N_13496,N_14639);
nor U18902 (N_18902,N_13764,N_12499);
and U18903 (N_18903,N_11399,N_12492);
nand U18904 (N_18904,N_13194,N_11547);
nand U18905 (N_18905,N_11105,N_10585);
nand U18906 (N_18906,N_11669,N_14921);
and U18907 (N_18907,N_11473,N_12943);
and U18908 (N_18908,N_13138,N_10982);
and U18909 (N_18909,N_13567,N_14718);
or U18910 (N_18910,N_11554,N_10318);
nor U18911 (N_18911,N_13031,N_11105);
nor U18912 (N_18912,N_13203,N_10477);
nor U18913 (N_18913,N_13538,N_12365);
nand U18914 (N_18914,N_11400,N_11826);
nand U18915 (N_18915,N_12085,N_13666);
or U18916 (N_18916,N_12508,N_13411);
and U18917 (N_18917,N_11076,N_11469);
and U18918 (N_18918,N_10392,N_10705);
or U18919 (N_18919,N_11645,N_14713);
nor U18920 (N_18920,N_12507,N_11380);
nand U18921 (N_18921,N_13061,N_13529);
nand U18922 (N_18922,N_14810,N_11280);
and U18923 (N_18923,N_14339,N_10348);
nand U18924 (N_18924,N_13295,N_14811);
or U18925 (N_18925,N_11767,N_10899);
and U18926 (N_18926,N_14974,N_10775);
and U18927 (N_18927,N_11584,N_13076);
and U18928 (N_18928,N_10227,N_12640);
nor U18929 (N_18929,N_11872,N_13216);
and U18930 (N_18930,N_11273,N_10648);
nand U18931 (N_18931,N_12662,N_14770);
nand U18932 (N_18932,N_11641,N_14749);
nor U18933 (N_18933,N_10955,N_12813);
and U18934 (N_18934,N_12392,N_12705);
nor U18935 (N_18935,N_10218,N_12936);
and U18936 (N_18936,N_14995,N_11963);
or U18937 (N_18937,N_11018,N_14025);
or U18938 (N_18938,N_10305,N_12923);
nand U18939 (N_18939,N_11268,N_11276);
nand U18940 (N_18940,N_11680,N_12748);
or U18941 (N_18941,N_12222,N_11995);
nand U18942 (N_18942,N_12697,N_11560);
nand U18943 (N_18943,N_12995,N_10571);
xor U18944 (N_18944,N_11115,N_12301);
nor U18945 (N_18945,N_10618,N_10757);
or U18946 (N_18946,N_14209,N_14177);
nand U18947 (N_18947,N_13797,N_14055);
nor U18948 (N_18948,N_11867,N_12142);
nand U18949 (N_18949,N_11656,N_13632);
and U18950 (N_18950,N_13781,N_12531);
nor U18951 (N_18951,N_10314,N_12135);
nor U18952 (N_18952,N_14931,N_11124);
or U18953 (N_18953,N_14259,N_10107);
or U18954 (N_18954,N_14505,N_13274);
nor U18955 (N_18955,N_13496,N_12024);
or U18956 (N_18956,N_13587,N_13687);
or U18957 (N_18957,N_12302,N_12682);
or U18958 (N_18958,N_10630,N_13641);
or U18959 (N_18959,N_12774,N_14929);
nor U18960 (N_18960,N_13496,N_13644);
and U18961 (N_18961,N_11958,N_13088);
and U18962 (N_18962,N_11996,N_14769);
nand U18963 (N_18963,N_11467,N_12381);
and U18964 (N_18964,N_13035,N_13322);
nor U18965 (N_18965,N_13868,N_12880);
and U18966 (N_18966,N_13710,N_14324);
and U18967 (N_18967,N_13277,N_13010);
and U18968 (N_18968,N_13698,N_13814);
nand U18969 (N_18969,N_11193,N_12930);
xor U18970 (N_18970,N_13354,N_10185);
or U18971 (N_18971,N_14189,N_13931);
nor U18972 (N_18972,N_12625,N_14371);
nand U18973 (N_18973,N_12018,N_13574);
and U18974 (N_18974,N_14034,N_10664);
or U18975 (N_18975,N_13328,N_11318);
or U18976 (N_18976,N_11975,N_12445);
or U18977 (N_18977,N_13456,N_12299);
or U18978 (N_18978,N_11728,N_12487);
nor U18979 (N_18979,N_11949,N_13929);
nor U18980 (N_18980,N_12997,N_10200);
or U18981 (N_18981,N_12335,N_11790);
nor U18982 (N_18982,N_14264,N_12775);
or U18983 (N_18983,N_14948,N_11688);
or U18984 (N_18984,N_14586,N_10269);
nor U18985 (N_18985,N_10811,N_14983);
or U18986 (N_18986,N_12570,N_14652);
nand U18987 (N_18987,N_13029,N_12091);
nand U18988 (N_18988,N_11511,N_14780);
nand U18989 (N_18989,N_11445,N_12235);
nand U18990 (N_18990,N_10216,N_13003);
nand U18991 (N_18991,N_13731,N_10439);
nor U18992 (N_18992,N_11140,N_14057);
or U18993 (N_18993,N_14576,N_14921);
xor U18994 (N_18994,N_10534,N_14677);
nor U18995 (N_18995,N_10687,N_11218);
and U18996 (N_18996,N_13579,N_14559);
and U18997 (N_18997,N_13580,N_12653);
nor U18998 (N_18998,N_10610,N_14170);
or U18999 (N_18999,N_10604,N_10686);
nor U19000 (N_19000,N_12942,N_13219);
nor U19001 (N_19001,N_13932,N_14330);
and U19002 (N_19002,N_10023,N_11906);
nand U19003 (N_19003,N_14191,N_12821);
nor U19004 (N_19004,N_13754,N_11052);
or U19005 (N_19005,N_11304,N_10554);
and U19006 (N_19006,N_13503,N_12271);
nand U19007 (N_19007,N_14119,N_10951);
nand U19008 (N_19008,N_12150,N_14829);
or U19009 (N_19009,N_11775,N_12517);
or U19010 (N_19010,N_14070,N_10024);
nand U19011 (N_19011,N_13955,N_10855);
and U19012 (N_19012,N_12674,N_12663);
nor U19013 (N_19013,N_14776,N_14838);
and U19014 (N_19014,N_12521,N_14293);
nor U19015 (N_19015,N_11157,N_14015);
or U19016 (N_19016,N_11598,N_13505);
and U19017 (N_19017,N_13508,N_10100);
nor U19018 (N_19018,N_12981,N_14487);
and U19019 (N_19019,N_14383,N_11808);
or U19020 (N_19020,N_10543,N_11806);
nor U19021 (N_19021,N_10783,N_12785);
nand U19022 (N_19022,N_14081,N_14934);
or U19023 (N_19023,N_11225,N_13878);
nor U19024 (N_19024,N_11288,N_13260);
or U19025 (N_19025,N_13307,N_14517);
or U19026 (N_19026,N_13828,N_12169);
nor U19027 (N_19027,N_11127,N_12083);
nor U19028 (N_19028,N_14614,N_10930);
or U19029 (N_19029,N_11623,N_13705);
and U19030 (N_19030,N_11321,N_14281);
and U19031 (N_19031,N_10714,N_14697);
nand U19032 (N_19032,N_13933,N_13656);
nand U19033 (N_19033,N_11884,N_10955);
and U19034 (N_19034,N_14137,N_14838);
or U19035 (N_19035,N_11589,N_13556);
nand U19036 (N_19036,N_13641,N_11726);
nor U19037 (N_19037,N_14942,N_13410);
and U19038 (N_19038,N_12527,N_13027);
and U19039 (N_19039,N_14049,N_13162);
or U19040 (N_19040,N_12727,N_11063);
or U19041 (N_19041,N_11515,N_12034);
nor U19042 (N_19042,N_14133,N_13513);
nand U19043 (N_19043,N_14330,N_13571);
nand U19044 (N_19044,N_13609,N_13730);
and U19045 (N_19045,N_10695,N_12513);
and U19046 (N_19046,N_13197,N_12155);
nor U19047 (N_19047,N_10637,N_14818);
or U19048 (N_19048,N_10044,N_12825);
and U19049 (N_19049,N_11887,N_11738);
or U19050 (N_19050,N_10153,N_11641);
xnor U19051 (N_19051,N_11621,N_11836);
nand U19052 (N_19052,N_11162,N_10158);
or U19053 (N_19053,N_10120,N_13432);
nand U19054 (N_19054,N_10980,N_11625);
nor U19055 (N_19055,N_13785,N_11784);
nand U19056 (N_19056,N_11864,N_12162);
nand U19057 (N_19057,N_11810,N_13694);
nand U19058 (N_19058,N_14698,N_12935);
nor U19059 (N_19059,N_14546,N_14095);
or U19060 (N_19060,N_13077,N_12589);
nor U19061 (N_19061,N_11258,N_10723);
nor U19062 (N_19062,N_12085,N_10097);
or U19063 (N_19063,N_13339,N_12338);
and U19064 (N_19064,N_14362,N_11554);
nand U19065 (N_19065,N_11844,N_13409);
and U19066 (N_19066,N_14042,N_11086);
nand U19067 (N_19067,N_10916,N_12388);
nor U19068 (N_19068,N_13341,N_11355);
nor U19069 (N_19069,N_10408,N_13473);
and U19070 (N_19070,N_11293,N_11487);
or U19071 (N_19071,N_14099,N_11276);
and U19072 (N_19072,N_12235,N_14163);
nand U19073 (N_19073,N_10372,N_12039);
nor U19074 (N_19074,N_11931,N_14756);
nand U19075 (N_19075,N_13242,N_13974);
nand U19076 (N_19076,N_10584,N_10008);
or U19077 (N_19077,N_14422,N_12919);
nor U19078 (N_19078,N_12078,N_12065);
nand U19079 (N_19079,N_13702,N_13712);
nand U19080 (N_19080,N_14203,N_11083);
nand U19081 (N_19081,N_12507,N_11729);
or U19082 (N_19082,N_12929,N_12388);
nor U19083 (N_19083,N_11650,N_10482);
or U19084 (N_19084,N_11708,N_13053);
nor U19085 (N_19085,N_12117,N_10200);
nor U19086 (N_19086,N_13610,N_14347);
nand U19087 (N_19087,N_13939,N_10585);
or U19088 (N_19088,N_12871,N_14198);
nor U19089 (N_19089,N_12193,N_14306);
or U19090 (N_19090,N_13206,N_13986);
nor U19091 (N_19091,N_10888,N_11437);
nor U19092 (N_19092,N_10719,N_10723);
and U19093 (N_19093,N_12472,N_12180);
nor U19094 (N_19094,N_12871,N_14547);
or U19095 (N_19095,N_12888,N_11311);
or U19096 (N_19096,N_10511,N_14252);
or U19097 (N_19097,N_12338,N_10122);
nor U19098 (N_19098,N_11940,N_12468);
nand U19099 (N_19099,N_10287,N_14885);
nand U19100 (N_19100,N_12565,N_14899);
or U19101 (N_19101,N_11725,N_12800);
or U19102 (N_19102,N_14185,N_13536);
nor U19103 (N_19103,N_12857,N_10490);
and U19104 (N_19104,N_14819,N_10183);
nand U19105 (N_19105,N_11988,N_10404);
or U19106 (N_19106,N_14986,N_13832);
and U19107 (N_19107,N_12023,N_13129);
and U19108 (N_19108,N_11733,N_14310);
nand U19109 (N_19109,N_10175,N_12703);
nand U19110 (N_19110,N_13950,N_13798);
and U19111 (N_19111,N_14483,N_12700);
or U19112 (N_19112,N_12113,N_14504);
or U19113 (N_19113,N_10781,N_14992);
and U19114 (N_19114,N_11201,N_11241);
nand U19115 (N_19115,N_11473,N_12996);
and U19116 (N_19116,N_14549,N_10049);
and U19117 (N_19117,N_12855,N_14807);
nand U19118 (N_19118,N_14715,N_10987);
or U19119 (N_19119,N_11299,N_13505);
nor U19120 (N_19120,N_13155,N_13867);
nand U19121 (N_19121,N_11280,N_14449);
or U19122 (N_19122,N_14993,N_13979);
or U19123 (N_19123,N_10800,N_12335);
and U19124 (N_19124,N_10628,N_11042);
nand U19125 (N_19125,N_14762,N_10751);
and U19126 (N_19126,N_11261,N_12950);
nor U19127 (N_19127,N_10368,N_12061);
or U19128 (N_19128,N_13244,N_14063);
and U19129 (N_19129,N_10404,N_11727);
and U19130 (N_19130,N_10511,N_10277);
nor U19131 (N_19131,N_11588,N_11682);
nand U19132 (N_19132,N_13263,N_13638);
nand U19133 (N_19133,N_13961,N_13798);
xor U19134 (N_19134,N_14820,N_14689);
nor U19135 (N_19135,N_10099,N_13981);
and U19136 (N_19136,N_14504,N_10355);
nor U19137 (N_19137,N_12512,N_10243);
or U19138 (N_19138,N_11265,N_12837);
and U19139 (N_19139,N_13610,N_12456);
and U19140 (N_19140,N_11972,N_13501);
nor U19141 (N_19141,N_10263,N_13305);
nor U19142 (N_19142,N_13134,N_12176);
nor U19143 (N_19143,N_11331,N_12410);
and U19144 (N_19144,N_13754,N_14137);
or U19145 (N_19145,N_13305,N_10435);
nor U19146 (N_19146,N_12785,N_10189);
nor U19147 (N_19147,N_14728,N_11121);
nand U19148 (N_19148,N_14814,N_12150);
nand U19149 (N_19149,N_13256,N_14503);
nor U19150 (N_19150,N_11242,N_14374);
nor U19151 (N_19151,N_11552,N_12047);
nand U19152 (N_19152,N_10349,N_10537);
and U19153 (N_19153,N_11560,N_10669);
or U19154 (N_19154,N_13264,N_11812);
nand U19155 (N_19155,N_14904,N_12414);
and U19156 (N_19156,N_13885,N_12262);
and U19157 (N_19157,N_14014,N_13726);
and U19158 (N_19158,N_13919,N_13467);
or U19159 (N_19159,N_12256,N_11004);
or U19160 (N_19160,N_11062,N_11801);
nor U19161 (N_19161,N_11065,N_12666);
or U19162 (N_19162,N_14287,N_14899);
and U19163 (N_19163,N_13181,N_10605);
nand U19164 (N_19164,N_14998,N_10345);
or U19165 (N_19165,N_13418,N_11450);
nand U19166 (N_19166,N_14016,N_14967);
or U19167 (N_19167,N_10074,N_14859);
and U19168 (N_19168,N_12586,N_10832);
nand U19169 (N_19169,N_14006,N_13862);
nor U19170 (N_19170,N_12131,N_12845);
or U19171 (N_19171,N_10183,N_14750);
and U19172 (N_19172,N_12987,N_13009);
and U19173 (N_19173,N_14504,N_12422);
nor U19174 (N_19174,N_10023,N_11755);
nand U19175 (N_19175,N_13347,N_10032);
or U19176 (N_19176,N_12706,N_14499);
nand U19177 (N_19177,N_12644,N_12204);
and U19178 (N_19178,N_12626,N_11983);
or U19179 (N_19179,N_10975,N_11186);
and U19180 (N_19180,N_14686,N_13861);
nor U19181 (N_19181,N_10568,N_10711);
and U19182 (N_19182,N_11001,N_12977);
and U19183 (N_19183,N_12818,N_10107);
or U19184 (N_19184,N_13098,N_12132);
nand U19185 (N_19185,N_10528,N_13903);
and U19186 (N_19186,N_13332,N_12901);
and U19187 (N_19187,N_13149,N_10102);
nand U19188 (N_19188,N_10940,N_14075);
and U19189 (N_19189,N_13544,N_12256);
and U19190 (N_19190,N_13198,N_12999);
nor U19191 (N_19191,N_12547,N_10112);
or U19192 (N_19192,N_13901,N_13538);
or U19193 (N_19193,N_14757,N_14133);
and U19194 (N_19194,N_14571,N_11868);
nand U19195 (N_19195,N_12155,N_10352);
or U19196 (N_19196,N_11547,N_13599);
and U19197 (N_19197,N_10748,N_11548);
and U19198 (N_19198,N_10357,N_14489);
nor U19199 (N_19199,N_11897,N_14984);
and U19200 (N_19200,N_12679,N_14711);
and U19201 (N_19201,N_14138,N_11458);
and U19202 (N_19202,N_10205,N_13448);
and U19203 (N_19203,N_12443,N_14009);
nor U19204 (N_19204,N_14225,N_10075);
and U19205 (N_19205,N_13592,N_12041);
or U19206 (N_19206,N_14007,N_13025);
nand U19207 (N_19207,N_12051,N_12541);
or U19208 (N_19208,N_14648,N_14968);
and U19209 (N_19209,N_14345,N_14721);
nand U19210 (N_19210,N_12372,N_11945);
nand U19211 (N_19211,N_14364,N_12214);
nand U19212 (N_19212,N_12317,N_11558);
or U19213 (N_19213,N_11267,N_10173);
and U19214 (N_19214,N_11564,N_13759);
and U19215 (N_19215,N_11329,N_13144);
xnor U19216 (N_19216,N_12318,N_10776);
nor U19217 (N_19217,N_12085,N_12555);
nand U19218 (N_19218,N_13198,N_14652);
nor U19219 (N_19219,N_10458,N_10050);
and U19220 (N_19220,N_10565,N_13717);
and U19221 (N_19221,N_14702,N_12095);
nand U19222 (N_19222,N_11070,N_10096);
or U19223 (N_19223,N_12920,N_13920);
nor U19224 (N_19224,N_13451,N_11913);
and U19225 (N_19225,N_10452,N_10434);
nor U19226 (N_19226,N_10870,N_11611);
nand U19227 (N_19227,N_13054,N_12207);
nand U19228 (N_19228,N_12189,N_10746);
and U19229 (N_19229,N_12980,N_14482);
and U19230 (N_19230,N_14181,N_10586);
nor U19231 (N_19231,N_13091,N_10765);
nand U19232 (N_19232,N_13085,N_13344);
nor U19233 (N_19233,N_10504,N_11152);
and U19234 (N_19234,N_14286,N_12753);
nand U19235 (N_19235,N_14984,N_10964);
and U19236 (N_19236,N_11569,N_11575);
nor U19237 (N_19237,N_10417,N_13652);
nand U19238 (N_19238,N_11615,N_12686);
nand U19239 (N_19239,N_11841,N_10549);
and U19240 (N_19240,N_13969,N_13151);
and U19241 (N_19241,N_13511,N_11935);
nor U19242 (N_19242,N_12058,N_12408);
nand U19243 (N_19243,N_12709,N_11695);
nor U19244 (N_19244,N_11509,N_14065);
or U19245 (N_19245,N_14157,N_12310);
nor U19246 (N_19246,N_13994,N_11621);
nand U19247 (N_19247,N_12958,N_13802);
and U19248 (N_19248,N_11101,N_10717);
nor U19249 (N_19249,N_10413,N_13634);
or U19250 (N_19250,N_13891,N_11360);
nor U19251 (N_19251,N_13226,N_13643);
nor U19252 (N_19252,N_10403,N_10471);
or U19253 (N_19253,N_12414,N_11599);
or U19254 (N_19254,N_14446,N_10772);
nor U19255 (N_19255,N_11119,N_10110);
nand U19256 (N_19256,N_13838,N_10600);
and U19257 (N_19257,N_13007,N_12226);
nand U19258 (N_19258,N_10928,N_11655);
xnor U19259 (N_19259,N_14352,N_10589);
nand U19260 (N_19260,N_10493,N_10114);
and U19261 (N_19261,N_13605,N_10197);
and U19262 (N_19262,N_13929,N_14565);
nor U19263 (N_19263,N_11656,N_12533);
nor U19264 (N_19264,N_10146,N_13801);
nor U19265 (N_19265,N_10269,N_11669);
nor U19266 (N_19266,N_10477,N_12065);
or U19267 (N_19267,N_12626,N_12091);
and U19268 (N_19268,N_13838,N_14998);
and U19269 (N_19269,N_12675,N_13755);
nor U19270 (N_19270,N_11520,N_10508);
nand U19271 (N_19271,N_12261,N_12629);
nand U19272 (N_19272,N_11070,N_10994);
nor U19273 (N_19273,N_12397,N_14840);
and U19274 (N_19274,N_10809,N_10093);
or U19275 (N_19275,N_14773,N_13003);
nor U19276 (N_19276,N_10265,N_10735);
and U19277 (N_19277,N_14101,N_13083);
nand U19278 (N_19278,N_10545,N_13838);
or U19279 (N_19279,N_12111,N_14491);
nand U19280 (N_19280,N_14185,N_13365);
or U19281 (N_19281,N_10327,N_13059);
or U19282 (N_19282,N_11043,N_11040);
nor U19283 (N_19283,N_12352,N_11218);
and U19284 (N_19284,N_11957,N_13672);
nor U19285 (N_19285,N_10539,N_13018);
nand U19286 (N_19286,N_13162,N_12379);
or U19287 (N_19287,N_14231,N_12057);
or U19288 (N_19288,N_13348,N_10375);
nor U19289 (N_19289,N_10274,N_11481);
nor U19290 (N_19290,N_10120,N_13878);
nand U19291 (N_19291,N_10624,N_11517);
or U19292 (N_19292,N_10865,N_11044);
and U19293 (N_19293,N_12799,N_11529);
and U19294 (N_19294,N_14828,N_10631);
nor U19295 (N_19295,N_12641,N_14588);
and U19296 (N_19296,N_14329,N_14437);
nor U19297 (N_19297,N_13216,N_10089);
nor U19298 (N_19298,N_11206,N_13980);
nand U19299 (N_19299,N_12219,N_10706);
nand U19300 (N_19300,N_10016,N_13839);
or U19301 (N_19301,N_13004,N_12886);
nor U19302 (N_19302,N_14500,N_14108);
and U19303 (N_19303,N_14497,N_10009);
or U19304 (N_19304,N_11105,N_13811);
or U19305 (N_19305,N_13194,N_12054);
nor U19306 (N_19306,N_14191,N_14703);
and U19307 (N_19307,N_12530,N_14611);
or U19308 (N_19308,N_14417,N_12509);
and U19309 (N_19309,N_11334,N_14448);
and U19310 (N_19310,N_14310,N_11889);
and U19311 (N_19311,N_10342,N_14066);
nand U19312 (N_19312,N_13980,N_10642);
and U19313 (N_19313,N_10362,N_13683);
nand U19314 (N_19314,N_14170,N_11525);
nand U19315 (N_19315,N_12561,N_12594);
or U19316 (N_19316,N_11358,N_12188);
or U19317 (N_19317,N_12960,N_10314);
nand U19318 (N_19318,N_13317,N_12705);
nand U19319 (N_19319,N_14102,N_13322);
and U19320 (N_19320,N_11527,N_13306);
and U19321 (N_19321,N_14394,N_12500);
nand U19322 (N_19322,N_10796,N_14214);
nand U19323 (N_19323,N_12272,N_12675);
nand U19324 (N_19324,N_11956,N_10823);
nor U19325 (N_19325,N_13342,N_11169);
or U19326 (N_19326,N_14321,N_14735);
nand U19327 (N_19327,N_11552,N_12599);
nor U19328 (N_19328,N_12729,N_13428);
nor U19329 (N_19329,N_12047,N_10931);
or U19330 (N_19330,N_10683,N_10672);
nand U19331 (N_19331,N_14084,N_10073);
xnor U19332 (N_19332,N_13144,N_12518);
nand U19333 (N_19333,N_11279,N_11338);
xor U19334 (N_19334,N_12028,N_10161);
or U19335 (N_19335,N_12358,N_12956);
nand U19336 (N_19336,N_11659,N_12553);
nor U19337 (N_19337,N_13205,N_12882);
or U19338 (N_19338,N_13577,N_12464);
nand U19339 (N_19339,N_14440,N_14828);
nor U19340 (N_19340,N_13694,N_12297);
nor U19341 (N_19341,N_10596,N_14745);
nor U19342 (N_19342,N_10090,N_11879);
and U19343 (N_19343,N_11322,N_13435);
or U19344 (N_19344,N_10536,N_14262);
and U19345 (N_19345,N_10697,N_12377);
nor U19346 (N_19346,N_12471,N_14505);
xor U19347 (N_19347,N_10088,N_12485);
and U19348 (N_19348,N_11051,N_12772);
or U19349 (N_19349,N_14741,N_12831);
or U19350 (N_19350,N_12338,N_14886);
and U19351 (N_19351,N_14868,N_11617);
and U19352 (N_19352,N_13440,N_11160);
and U19353 (N_19353,N_10248,N_10886);
nand U19354 (N_19354,N_14442,N_12227);
and U19355 (N_19355,N_11242,N_14800);
nor U19356 (N_19356,N_12032,N_14928);
nor U19357 (N_19357,N_10538,N_13978);
nand U19358 (N_19358,N_11496,N_12680);
nand U19359 (N_19359,N_11792,N_11748);
or U19360 (N_19360,N_11259,N_14780);
nor U19361 (N_19361,N_12408,N_12593);
nor U19362 (N_19362,N_12360,N_14107);
nand U19363 (N_19363,N_11208,N_13237);
nor U19364 (N_19364,N_10829,N_11704);
or U19365 (N_19365,N_11932,N_14213);
nor U19366 (N_19366,N_11398,N_12835);
nor U19367 (N_19367,N_12819,N_10759);
nand U19368 (N_19368,N_11629,N_13814);
and U19369 (N_19369,N_11845,N_10721);
or U19370 (N_19370,N_11069,N_12409);
and U19371 (N_19371,N_11978,N_13733);
or U19372 (N_19372,N_10346,N_13060);
nand U19373 (N_19373,N_13578,N_14347);
and U19374 (N_19374,N_12343,N_13308);
nor U19375 (N_19375,N_11531,N_11326);
nand U19376 (N_19376,N_14346,N_14221);
nor U19377 (N_19377,N_11554,N_10145);
and U19378 (N_19378,N_10276,N_12060);
nand U19379 (N_19379,N_13380,N_10043);
and U19380 (N_19380,N_14600,N_11851);
and U19381 (N_19381,N_13739,N_12331);
nor U19382 (N_19382,N_13914,N_13288);
or U19383 (N_19383,N_11722,N_12596);
or U19384 (N_19384,N_14975,N_13831);
and U19385 (N_19385,N_10035,N_12973);
nor U19386 (N_19386,N_11622,N_10449);
nand U19387 (N_19387,N_14108,N_13823);
nand U19388 (N_19388,N_13533,N_12487);
and U19389 (N_19389,N_12739,N_14027);
and U19390 (N_19390,N_13711,N_12005);
nand U19391 (N_19391,N_14888,N_10966);
or U19392 (N_19392,N_12049,N_13982);
nor U19393 (N_19393,N_13709,N_10917);
nand U19394 (N_19394,N_13148,N_13537);
nor U19395 (N_19395,N_14396,N_12104);
nand U19396 (N_19396,N_10376,N_10397);
nand U19397 (N_19397,N_13362,N_14480);
and U19398 (N_19398,N_11911,N_12731);
nor U19399 (N_19399,N_10167,N_11300);
or U19400 (N_19400,N_13843,N_14202);
nor U19401 (N_19401,N_11212,N_13667);
and U19402 (N_19402,N_14560,N_11589);
or U19403 (N_19403,N_13598,N_14641);
nand U19404 (N_19404,N_14289,N_10107);
or U19405 (N_19405,N_12696,N_10654);
or U19406 (N_19406,N_10459,N_11926);
or U19407 (N_19407,N_14297,N_10273);
and U19408 (N_19408,N_13787,N_10726);
or U19409 (N_19409,N_14302,N_12286);
and U19410 (N_19410,N_12627,N_11663);
and U19411 (N_19411,N_11359,N_14265);
nand U19412 (N_19412,N_13680,N_14509);
or U19413 (N_19413,N_13094,N_13251);
xnor U19414 (N_19414,N_10323,N_14216);
nand U19415 (N_19415,N_11006,N_11603);
or U19416 (N_19416,N_13493,N_14975);
nor U19417 (N_19417,N_14544,N_14863);
nor U19418 (N_19418,N_12091,N_14320);
nor U19419 (N_19419,N_11295,N_11433);
nand U19420 (N_19420,N_13744,N_12363);
or U19421 (N_19421,N_13847,N_14924);
and U19422 (N_19422,N_14164,N_10330);
and U19423 (N_19423,N_11115,N_14301);
nor U19424 (N_19424,N_10703,N_14818);
nor U19425 (N_19425,N_12682,N_14724);
nand U19426 (N_19426,N_11944,N_13209);
nand U19427 (N_19427,N_13586,N_11571);
nor U19428 (N_19428,N_14174,N_14223);
nor U19429 (N_19429,N_11592,N_11104);
nand U19430 (N_19430,N_12424,N_14931);
or U19431 (N_19431,N_12266,N_11426);
or U19432 (N_19432,N_12986,N_11377);
and U19433 (N_19433,N_14920,N_12090);
or U19434 (N_19434,N_13166,N_11631);
and U19435 (N_19435,N_12146,N_14702);
xor U19436 (N_19436,N_10276,N_11473);
and U19437 (N_19437,N_13278,N_10638);
or U19438 (N_19438,N_13376,N_11569);
nor U19439 (N_19439,N_12555,N_11537);
nor U19440 (N_19440,N_12626,N_12606);
nand U19441 (N_19441,N_10926,N_14691);
nand U19442 (N_19442,N_14048,N_12059);
nand U19443 (N_19443,N_14840,N_14718);
or U19444 (N_19444,N_14417,N_14588);
nor U19445 (N_19445,N_11311,N_11268);
nand U19446 (N_19446,N_14472,N_14469);
and U19447 (N_19447,N_10487,N_13206);
nand U19448 (N_19448,N_14706,N_13382);
nor U19449 (N_19449,N_13494,N_14004);
or U19450 (N_19450,N_13420,N_11599);
nand U19451 (N_19451,N_13343,N_14130);
nand U19452 (N_19452,N_13870,N_10051);
and U19453 (N_19453,N_12668,N_10036);
and U19454 (N_19454,N_11279,N_11802);
xor U19455 (N_19455,N_11615,N_13964);
nor U19456 (N_19456,N_10360,N_13963);
and U19457 (N_19457,N_12946,N_11775);
or U19458 (N_19458,N_11644,N_10885);
or U19459 (N_19459,N_10422,N_14902);
nand U19460 (N_19460,N_14399,N_10110);
nor U19461 (N_19461,N_12813,N_14504);
and U19462 (N_19462,N_10083,N_13671);
or U19463 (N_19463,N_11362,N_12207);
or U19464 (N_19464,N_12765,N_10626);
or U19465 (N_19465,N_11763,N_13751);
and U19466 (N_19466,N_12915,N_10029);
nand U19467 (N_19467,N_13190,N_13358);
nand U19468 (N_19468,N_11811,N_13518);
and U19469 (N_19469,N_14328,N_14371);
or U19470 (N_19470,N_13207,N_13165);
nand U19471 (N_19471,N_10755,N_12087);
nand U19472 (N_19472,N_10685,N_12315);
or U19473 (N_19473,N_14694,N_11171);
or U19474 (N_19474,N_11319,N_12088);
nor U19475 (N_19475,N_10907,N_13538);
and U19476 (N_19476,N_12188,N_14809);
or U19477 (N_19477,N_12291,N_11099);
or U19478 (N_19478,N_13260,N_14333);
nand U19479 (N_19479,N_12046,N_11094);
nand U19480 (N_19480,N_12445,N_14826);
nand U19481 (N_19481,N_11767,N_11029);
or U19482 (N_19482,N_10732,N_14323);
or U19483 (N_19483,N_14028,N_10292);
or U19484 (N_19484,N_10744,N_12755);
nand U19485 (N_19485,N_12113,N_14199);
or U19486 (N_19486,N_11263,N_10274);
nor U19487 (N_19487,N_13595,N_10491);
nand U19488 (N_19488,N_14644,N_10275);
and U19489 (N_19489,N_10782,N_13153);
and U19490 (N_19490,N_13383,N_11660);
nand U19491 (N_19491,N_13287,N_13840);
or U19492 (N_19492,N_11634,N_12676);
nand U19493 (N_19493,N_13931,N_11971);
nor U19494 (N_19494,N_14050,N_12577);
nand U19495 (N_19495,N_13674,N_14967);
and U19496 (N_19496,N_13184,N_12120);
and U19497 (N_19497,N_14387,N_10623);
and U19498 (N_19498,N_12634,N_12454);
nor U19499 (N_19499,N_14920,N_12271);
and U19500 (N_19500,N_10242,N_10286);
and U19501 (N_19501,N_10178,N_10356);
nand U19502 (N_19502,N_14108,N_14898);
or U19503 (N_19503,N_11377,N_10674);
and U19504 (N_19504,N_10857,N_13393);
nor U19505 (N_19505,N_13139,N_10539);
nor U19506 (N_19506,N_11292,N_12994);
or U19507 (N_19507,N_11601,N_11505);
and U19508 (N_19508,N_12893,N_11757);
or U19509 (N_19509,N_10203,N_12477);
and U19510 (N_19510,N_14112,N_11628);
and U19511 (N_19511,N_11029,N_12585);
and U19512 (N_19512,N_13249,N_14611);
or U19513 (N_19513,N_11271,N_13236);
or U19514 (N_19514,N_13183,N_14181);
nor U19515 (N_19515,N_13388,N_11325);
or U19516 (N_19516,N_10202,N_12966);
and U19517 (N_19517,N_13606,N_10611);
nor U19518 (N_19518,N_13917,N_12476);
or U19519 (N_19519,N_11974,N_10055);
nand U19520 (N_19520,N_11932,N_10479);
nor U19521 (N_19521,N_12981,N_12088);
nor U19522 (N_19522,N_11057,N_10801);
or U19523 (N_19523,N_10052,N_12086);
nor U19524 (N_19524,N_10933,N_10614);
nand U19525 (N_19525,N_11537,N_13060);
nand U19526 (N_19526,N_14480,N_14796);
nor U19527 (N_19527,N_10726,N_13318);
and U19528 (N_19528,N_13770,N_14498);
or U19529 (N_19529,N_12484,N_11741);
or U19530 (N_19530,N_13674,N_11897);
nand U19531 (N_19531,N_11192,N_10682);
nor U19532 (N_19532,N_10740,N_11649);
nand U19533 (N_19533,N_12478,N_13268);
nor U19534 (N_19534,N_12947,N_12757);
or U19535 (N_19535,N_14861,N_10743);
nand U19536 (N_19536,N_11197,N_13635);
nor U19537 (N_19537,N_14203,N_13862);
nand U19538 (N_19538,N_11531,N_13804);
and U19539 (N_19539,N_11285,N_12780);
and U19540 (N_19540,N_11437,N_11551);
and U19541 (N_19541,N_12740,N_14212);
nor U19542 (N_19542,N_10403,N_13756);
or U19543 (N_19543,N_12690,N_14775);
nor U19544 (N_19544,N_14271,N_14951);
and U19545 (N_19545,N_10673,N_11793);
and U19546 (N_19546,N_10400,N_11775);
and U19547 (N_19547,N_12783,N_14532);
or U19548 (N_19548,N_12252,N_13614);
nor U19549 (N_19549,N_11309,N_11339);
and U19550 (N_19550,N_13798,N_12924);
nor U19551 (N_19551,N_14649,N_10219);
nand U19552 (N_19552,N_12395,N_12212);
nand U19553 (N_19553,N_14916,N_11514);
nor U19554 (N_19554,N_13427,N_12853);
and U19555 (N_19555,N_10760,N_10732);
nand U19556 (N_19556,N_13419,N_14561);
nand U19557 (N_19557,N_11261,N_12202);
or U19558 (N_19558,N_10854,N_10091);
nor U19559 (N_19559,N_14404,N_14068);
or U19560 (N_19560,N_11482,N_12875);
and U19561 (N_19561,N_13017,N_12831);
nand U19562 (N_19562,N_13826,N_14740);
or U19563 (N_19563,N_13048,N_11421);
nand U19564 (N_19564,N_11052,N_11699);
or U19565 (N_19565,N_10713,N_11848);
nand U19566 (N_19566,N_13562,N_11011);
and U19567 (N_19567,N_10949,N_14618);
nand U19568 (N_19568,N_11546,N_10795);
nand U19569 (N_19569,N_12477,N_10089);
or U19570 (N_19570,N_11907,N_11924);
and U19571 (N_19571,N_14568,N_14613);
nand U19572 (N_19572,N_11786,N_10446);
and U19573 (N_19573,N_10226,N_11852);
and U19574 (N_19574,N_11043,N_12701);
or U19575 (N_19575,N_12293,N_13333);
nor U19576 (N_19576,N_10965,N_12970);
and U19577 (N_19577,N_13568,N_11980);
or U19578 (N_19578,N_13294,N_13827);
nor U19579 (N_19579,N_12214,N_11584);
or U19580 (N_19580,N_12152,N_11327);
or U19581 (N_19581,N_13425,N_14090);
nor U19582 (N_19582,N_11244,N_12549);
and U19583 (N_19583,N_10914,N_14747);
and U19584 (N_19584,N_14570,N_13512);
nand U19585 (N_19585,N_10428,N_13208);
nand U19586 (N_19586,N_10841,N_12058);
and U19587 (N_19587,N_11780,N_12923);
or U19588 (N_19588,N_14553,N_13932);
and U19589 (N_19589,N_12422,N_14668);
or U19590 (N_19590,N_12228,N_11406);
and U19591 (N_19591,N_12787,N_14263);
nor U19592 (N_19592,N_14011,N_14812);
or U19593 (N_19593,N_11556,N_12857);
or U19594 (N_19594,N_12432,N_12528);
or U19595 (N_19595,N_10876,N_14352);
nand U19596 (N_19596,N_10160,N_12329);
nor U19597 (N_19597,N_13293,N_12731);
nor U19598 (N_19598,N_10237,N_12493);
nor U19599 (N_19599,N_12701,N_10182);
or U19600 (N_19600,N_13211,N_14763);
or U19601 (N_19601,N_10417,N_12131);
and U19602 (N_19602,N_13354,N_13474);
nor U19603 (N_19603,N_12522,N_13144);
or U19604 (N_19604,N_14330,N_10056);
nor U19605 (N_19605,N_13871,N_12679);
or U19606 (N_19606,N_12704,N_14949);
xnor U19607 (N_19607,N_14661,N_13059);
nor U19608 (N_19608,N_14636,N_11430);
nand U19609 (N_19609,N_10683,N_13584);
nor U19610 (N_19610,N_12638,N_13493);
nor U19611 (N_19611,N_12243,N_13139);
nor U19612 (N_19612,N_13316,N_12287);
or U19613 (N_19613,N_10366,N_13249);
nor U19614 (N_19614,N_14164,N_11114);
or U19615 (N_19615,N_14171,N_14443);
nor U19616 (N_19616,N_13264,N_12457);
and U19617 (N_19617,N_11296,N_10724);
and U19618 (N_19618,N_12962,N_14690);
or U19619 (N_19619,N_13531,N_11563);
and U19620 (N_19620,N_10061,N_10943);
nor U19621 (N_19621,N_10020,N_13760);
and U19622 (N_19622,N_10597,N_12952);
or U19623 (N_19623,N_13161,N_11474);
and U19624 (N_19624,N_11195,N_12961);
or U19625 (N_19625,N_13629,N_13497);
and U19626 (N_19626,N_14509,N_11940);
and U19627 (N_19627,N_11522,N_11932);
or U19628 (N_19628,N_10229,N_14682);
and U19629 (N_19629,N_12226,N_14216);
and U19630 (N_19630,N_14232,N_13129);
or U19631 (N_19631,N_12939,N_11253);
nand U19632 (N_19632,N_14602,N_12927);
nor U19633 (N_19633,N_14074,N_12941);
nor U19634 (N_19634,N_14330,N_10642);
and U19635 (N_19635,N_10257,N_14389);
nor U19636 (N_19636,N_13525,N_11949);
and U19637 (N_19637,N_13546,N_12444);
nor U19638 (N_19638,N_12726,N_13181);
and U19639 (N_19639,N_12800,N_12497);
nor U19640 (N_19640,N_10854,N_13494);
or U19641 (N_19641,N_12590,N_11886);
nand U19642 (N_19642,N_11403,N_10832);
nor U19643 (N_19643,N_12323,N_14919);
and U19644 (N_19644,N_14652,N_12429);
or U19645 (N_19645,N_10778,N_14708);
nor U19646 (N_19646,N_11883,N_11216);
and U19647 (N_19647,N_10484,N_12872);
and U19648 (N_19648,N_13147,N_14857);
nand U19649 (N_19649,N_10599,N_10050);
nand U19650 (N_19650,N_12809,N_14660);
nor U19651 (N_19651,N_14370,N_14211);
nand U19652 (N_19652,N_14878,N_13858);
nand U19653 (N_19653,N_11543,N_12423);
nand U19654 (N_19654,N_14753,N_13058);
and U19655 (N_19655,N_14155,N_14348);
nor U19656 (N_19656,N_10681,N_12076);
nor U19657 (N_19657,N_12696,N_13615);
or U19658 (N_19658,N_13356,N_14129);
nand U19659 (N_19659,N_13356,N_10278);
nor U19660 (N_19660,N_11412,N_12756);
nand U19661 (N_19661,N_10861,N_10146);
and U19662 (N_19662,N_14005,N_14870);
nor U19663 (N_19663,N_10819,N_14221);
or U19664 (N_19664,N_13389,N_14232);
and U19665 (N_19665,N_10770,N_11934);
and U19666 (N_19666,N_14373,N_11511);
nand U19667 (N_19667,N_10450,N_11521);
or U19668 (N_19668,N_13898,N_13901);
nor U19669 (N_19669,N_11231,N_13894);
nand U19670 (N_19670,N_13583,N_13348);
and U19671 (N_19671,N_12126,N_10444);
nand U19672 (N_19672,N_14979,N_10462);
nand U19673 (N_19673,N_14967,N_10526);
nor U19674 (N_19674,N_10979,N_14446);
nand U19675 (N_19675,N_14417,N_12519);
nor U19676 (N_19676,N_14379,N_13378);
xnor U19677 (N_19677,N_12257,N_14641);
nor U19678 (N_19678,N_14751,N_10965);
nor U19679 (N_19679,N_12310,N_14990);
xor U19680 (N_19680,N_11814,N_11609);
and U19681 (N_19681,N_14129,N_12265);
or U19682 (N_19682,N_10874,N_14123);
nor U19683 (N_19683,N_13515,N_10004);
nor U19684 (N_19684,N_12489,N_11396);
or U19685 (N_19685,N_10830,N_10846);
nand U19686 (N_19686,N_14009,N_11842);
and U19687 (N_19687,N_12426,N_14570);
or U19688 (N_19688,N_10357,N_12794);
and U19689 (N_19689,N_14278,N_12083);
nor U19690 (N_19690,N_12222,N_13462);
nand U19691 (N_19691,N_13269,N_11749);
and U19692 (N_19692,N_14175,N_10937);
nor U19693 (N_19693,N_11012,N_11842);
xnor U19694 (N_19694,N_13286,N_11451);
and U19695 (N_19695,N_14974,N_10728);
nand U19696 (N_19696,N_12977,N_12798);
nor U19697 (N_19697,N_13922,N_11724);
nand U19698 (N_19698,N_10729,N_10402);
nor U19699 (N_19699,N_11364,N_12270);
nor U19700 (N_19700,N_11172,N_14220);
nand U19701 (N_19701,N_10303,N_11077);
or U19702 (N_19702,N_13539,N_10640);
and U19703 (N_19703,N_13781,N_11394);
or U19704 (N_19704,N_11890,N_13735);
nor U19705 (N_19705,N_10121,N_14875);
or U19706 (N_19706,N_12104,N_13208);
nand U19707 (N_19707,N_12705,N_12474);
and U19708 (N_19708,N_11843,N_10835);
xor U19709 (N_19709,N_14042,N_11782);
nand U19710 (N_19710,N_12064,N_13802);
and U19711 (N_19711,N_10401,N_13124);
and U19712 (N_19712,N_10733,N_14888);
or U19713 (N_19713,N_13995,N_11671);
nor U19714 (N_19714,N_11829,N_10643);
or U19715 (N_19715,N_13118,N_13403);
nor U19716 (N_19716,N_13599,N_11252);
nand U19717 (N_19717,N_10765,N_11290);
or U19718 (N_19718,N_13373,N_11341);
nand U19719 (N_19719,N_12976,N_11929);
xor U19720 (N_19720,N_14094,N_10036);
nor U19721 (N_19721,N_11734,N_10998);
nor U19722 (N_19722,N_11768,N_10111);
nand U19723 (N_19723,N_14683,N_12197);
nand U19724 (N_19724,N_10288,N_11190);
nand U19725 (N_19725,N_12879,N_10533);
and U19726 (N_19726,N_12194,N_14053);
nand U19727 (N_19727,N_13165,N_11092);
nor U19728 (N_19728,N_14614,N_14412);
and U19729 (N_19729,N_11977,N_13193);
or U19730 (N_19730,N_14913,N_11229);
and U19731 (N_19731,N_12607,N_11452);
xnor U19732 (N_19732,N_14599,N_14564);
nor U19733 (N_19733,N_11309,N_13618);
or U19734 (N_19734,N_12576,N_12828);
and U19735 (N_19735,N_12521,N_11013);
and U19736 (N_19736,N_10835,N_10435);
or U19737 (N_19737,N_14778,N_10380);
or U19738 (N_19738,N_13388,N_14537);
and U19739 (N_19739,N_13897,N_14067);
nor U19740 (N_19740,N_10821,N_13836);
nor U19741 (N_19741,N_11037,N_12566);
or U19742 (N_19742,N_13566,N_11669);
nor U19743 (N_19743,N_13646,N_14062);
and U19744 (N_19744,N_13840,N_11855);
and U19745 (N_19745,N_12458,N_10435);
nand U19746 (N_19746,N_10702,N_14818);
and U19747 (N_19747,N_10068,N_13962);
and U19748 (N_19748,N_11414,N_12563);
nor U19749 (N_19749,N_10584,N_14488);
nor U19750 (N_19750,N_13671,N_12899);
nor U19751 (N_19751,N_11137,N_11647);
or U19752 (N_19752,N_11514,N_14386);
and U19753 (N_19753,N_11680,N_10141);
and U19754 (N_19754,N_11765,N_11696);
nor U19755 (N_19755,N_13373,N_12314);
xnor U19756 (N_19756,N_12572,N_12179);
or U19757 (N_19757,N_14571,N_14537);
nor U19758 (N_19758,N_10441,N_13385);
or U19759 (N_19759,N_11626,N_11892);
nand U19760 (N_19760,N_10990,N_12098);
or U19761 (N_19761,N_10793,N_11787);
or U19762 (N_19762,N_12268,N_14478);
and U19763 (N_19763,N_10117,N_12082);
nand U19764 (N_19764,N_13894,N_11999);
or U19765 (N_19765,N_14053,N_11467);
nor U19766 (N_19766,N_13128,N_11465);
nor U19767 (N_19767,N_11166,N_12800);
nor U19768 (N_19768,N_13988,N_13128);
nor U19769 (N_19769,N_14740,N_10784);
nand U19770 (N_19770,N_13331,N_14709);
or U19771 (N_19771,N_12584,N_13883);
nand U19772 (N_19772,N_14181,N_12160);
or U19773 (N_19773,N_14116,N_14710);
and U19774 (N_19774,N_14299,N_10822);
xnor U19775 (N_19775,N_11296,N_10463);
or U19776 (N_19776,N_12367,N_10536);
nand U19777 (N_19777,N_10813,N_10066);
or U19778 (N_19778,N_10955,N_14352);
nand U19779 (N_19779,N_10252,N_13987);
nand U19780 (N_19780,N_12825,N_13596);
and U19781 (N_19781,N_12541,N_13431);
nor U19782 (N_19782,N_11472,N_14347);
or U19783 (N_19783,N_14350,N_13504);
nor U19784 (N_19784,N_11528,N_11782);
and U19785 (N_19785,N_11792,N_14938);
nand U19786 (N_19786,N_11277,N_14367);
or U19787 (N_19787,N_10535,N_14236);
nor U19788 (N_19788,N_12438,N_12369);
and U19789 (N_19789,N_14370,N_10039);
and U19790 (N_19790,N_10897,N_10506);
nor U19791 (N_19791,N_12392,N_13241);
or U19792 (N_19792,N_12877,N_12274);
nor U19793 (N_19793,N_10707,N_10299);
nor U19794 (N_19794,N_12014,N_10244);
xor U19795 (N_19795,N_12318,N_10473);
or U19796 (N_19796,N_14380,N_10691);
and U19797 (N_19797,N_13233,N_13720);
and U19798 (N_19798,N_14499,N_12365);
or U19799 (N_19799,N_12109,N_14351);
nand U19800 (N_19800,N_12290,N_13728);
nor U19801 (N_19801,N_13967,N_14931);
nor U19802 (N_19802,N_13898,N_14261);
and U19803 (N_19803,N_12831,N_13375);
nor U19804 (N_19804,N_11754,N_13858);
nor U19805 (N_19805,N_12684,N_14538);
nor U19806 (N_19806,N_11975,N_13312);
and U19807 (N_19807,N_12178,N_12413);
nand U19808 (N_19808,N_10029,N_11356);
and U19809 (N_19809,N_10866,N_12224);
nand U19810 (N_19810,N_12740,N_10432);
nor U19811 (N_19811,N_10948,N_12700);
or U19812 (N_19812,N_12887,N_14152);
nand U19813 (N_19813,N_11704,N_11489);
or U19814 (N_19814,N_14171,N_14782);
nor U19815 (N_19815,N_12005,N_13150);
nand U19816 (N_19816,N_12867,N_12379);
nand U19817 (N_19817,N_14301,N_13831);
and U19818 (N_19818,N_13273,N_11787);
nor U19819 (N_19819,N_12866,N_11873);
nand U19820 (N_19820,N_10417,N_10733);
nor U19821 (N_19821,N_11159,N_10720);
or U19822 (N_19822,N_13805,N_13258);
nand U19823 (N_19823,N_13094,N_11413);
or U19824 (N_19824,N_14504,N_14007);
nor U19825 (N_19825,N_10809,N_12936);
or U19826 (N_19826,N_11081,N_13480);
nor U19827 (N_19827,N_11139,N_14905);
or U19828 (N_19828,N_10918,N_12232);
nand U19829 (N_19829,N_10569,N_13508);
and U19830 (N_19830,N_12492,N_12975);
or U19831 (N_19831,N_13144,N_10663);
and U19832 (N_19832,N_10751,N_11433);
nand U19833 (N_19833,N_11162,N_10566);
and U19834 (N_19834,N_13511,N_12262);
and U19835 (N_19835,N_10444,N_12897);
nor U19836 (N_19836,N_10877,N_13194);
and U19837 (N_19837,N_12589,N_12651);
and U19838 (N_19838,N_12550,N_12289);
nand U19839 (N_19839,N_10241,N_14441);
nor U19840 (N_19840,N_13547,N_14042);
nor U19841 (N_19841,N_11774,N_14062);
or U19842 (N_19842,N_12117,N_14413);
or U19843 (N_19843,N_14218,N_13643);
nand U19844 (N_19844,N_11948,N_12678);
nor U19845 (N_19845,N_13993,N_12144);
nand U19846 (N_19846,N_13617,N_10406);
and U19847 (N_19847,N_10175,N_14942);
nand U19848 (N_19848,N_13579,N_10971);
nand U19849 (N_19849,N_13799,N_11959);
nor U19850 (N_19850,N_14774,N_14449);
and U19851 (N_19851,N_13443,N_14273);
nand U19852 (N_19852,N_12421,N_13811);
xor U19853 (N_19853,N_14217,N_12103);
or U19854 (N_19854,N_12718,N_14509);
and U19855 (N_19855,N_10180,N_10476);
and U19856 (N_19856,N_11175,N_12731);
or U19857 (N_19857,N_14108,N_12572);
or U19858 (N_19858,N_13640,N_11759);
nor U19859 (N_19859,N_10677,N_12385);
and U19860 (N_19860,N_12025,N_14593);
or U19861 (N_19861,N_14302,N_11606);
or U19862 (N_19862,N_12363,N_10719);
or U19863 (N_19863,N_13162,N_12169);
nor U19864 (N_19864,N_10551,N_11119);
and U19865 (N_19865,N_11345,N_10055);
and U19866 (N_19866,N_10061,N_14852);
and U19867 (N_19867,N_14978,N_14299);
nor U19868 (N_19868,N_14547,N_14404);
nand U19869 (N_19869,N_13244,N_11908);
nor U19870 (N_19870,N_14173,N_11116);
and U19871 (N_19871,N_11892,N_14209);
or U19872 (N_19872,N_11800,N_14333);
and U19873 (N_19873,N_11593,N_11928);
nor U19874 (N_19874,N_11329,N_13303);
nor U19875 (N_19875,N_12096,N_10024);
or U19876 (N_19876,N_12387,N_14334);
and U19877 (N_19877,N_13724,N_14817);
nand U19878 (N_19878,N_13772,N_11971);
or U19879 (N_19879,N_14748,N_12368);
or U19880 (N_19880,N_12569,N_14993);
and U19881 (N_19881,N_10156,N_12281);
nor U19882 (N_19882,N_10183,N_13530);
nor U19883 (N_19883,N_11886,N_11291);
nand U19884 (N_19884,N_12420,N_12990);
nand U19885 (N_19885,N_14719,N_10379);
nor U19886 (N_19886,N_13920,N_13590);
nand U19887 (N_19887,N_14323,N_13670);
nor U19888 (N_19888,N_14153,N_12715);
and U19889 (N_19889,N_11960,N_13190);
nand U19890 (N_19890,N_14887,N_12143);
or U19891 (N_19891,N_12908,N_13956);
and U19892 (N_19892,N_13156,N_14504);
nand U19893 (N_19893,N_11246,N_10893);
nor U19894 (N_19894,N_14612,N_14301);
nor U19895 (N_19895,N_13873,N_13013);
nand U19896 (N_19896,N_12940,N_13586);
and U19897 (N_19897,N_11057,N_10501);
and U19898 (N_19898,N_10637,N_10063);
and U19899 (N_19899,N_13864,N_12546);
or U19900 (N_19900,N_10541,N_13884);
and U19901 (N_19901,N_12472,N_12543);
and U19902 (N_19902,N_12615,N_12096);
nand U19903 (N_19903,N_14563,N_10769);
nand U19904 (N_19904,N_14963,N_11811);
nand U19905 (N_19905,N_11361,N_13104);
or U19906 (N_19906,N_14724,N_11447);
and U19907 (N_19907,N_13277,N_13806);
nand U19908 (N_19908,N_14943,N_11860);
nand U19909 (N_19909,N_14069,N_10448);
or U19910 (N_19910,N_13225,N_11555);
nand U19911 (N_19911,N_11163,N_14736);
or U19912 (N_19912,N_12005,N_13389);
nand U19913 (N_19913,N_10812,N_10799);
nand U19914 (N_19914,N_13879,N_11774);
and U19915 (N_19915,N_11331,N_12148);
or U19916 (N_19916,N_13519,N_14572);
or U19917 (N_19917,N_12902,N_12397);
and U19918 (N_19918,N_14094,N_14677);
or U19919 (N_19919,N_10359,N_10509);
or U19920 (N_19920,N_11395,N_13654);
or U19921 (N_19921,N_10987,N_10269);
nor U19922 (N_19922,N_14705,N_14961);
or U19923 (N_19923,N_11695,N_14237);
and U19924 (N_19924,N_10550,N_13146);
nand U19925 (N_19925,N_14616,N_12283);
nand U19926 (N_19926,N_14465,N_10160);
and U19927 (N_19927,N_11510,N_13565);
nand U19928 (N_19928,N_10121,N_12068);
and U19929 (N_19929,N_11197,N_12470);
nor U19930 (N_19930,N_11976,N_14614);
and U19931 (N_19931,N_13752,N_10908);
nor U19932 (N_19932,N_11920,N_14719);
nor U19933 (N_19933,N_14002,N_11513);
nand U19934 (N_19934,N_12786,N_14714);
nand U19935 (N_19935,N_12971,N_12868);
and U19936 (N_19936,N_11750,N_14816);
and U19937 (N_19937,N_14432,N_11460);
nand U19938 (N_19938,N_14495,N_12417);
nor U19939 (N_19939,N_11243,N_12041);
nor U19940 (N_19940,N_10719,N_13632);
nand U19941 (N_19941,N_13827,N_11656);
or U19942 (N_19942,N_10496,N_12309);
or U19943 (N_19943,N_14225,N_14918);
or U19944 (N_19944,N_13116,N_12033);
nor U19945 (N_19945,N_12901,N_10281);
and U19946 (N_19946,N_10088,N_11763);
and U19947 (N_19947,N_10177,N_13825);
and U19948 (N_19948,N_14308,N_11560);
or U19949 (N_19949,N_14366,N_12266);
or U19950 (N_19950,N_12943,N_10101);
and U19951 (N_19951,N_11874,N_10823);
and U19952 (N_19952,N_12940,N_14233);
nor U19953 (N_19953,N_13928,N_13276);
nand U19954 (N_19954,N_14697,N_14671);
or U19955 (N_19955,N_12276,N_10829);
or U19956 (N_19956,N_12074,N_11125);
nor U19957 (N_19957,N_13680,N_11253);
or U19958 (N_19958,N_13773,N_14396);
nand U19959 (N_19959,N_14301,N_10519);
nand U19960 (N_19960,N_14191,N_13686);
or U19961 (N_19961,N_10544,N_14032);
nand U19962 (N_19962,N_14958,N_11099);
or U19963 (N_19963,N_12812,N_12271);
and U19964 (N_19964,N_14158,N_10045);
and U19965 (N_19965,N_11793,N_11412);
nor U19966 (N_19966,N_10297,N_14510);
and U19967 (N_19967,N_14012,N_14263);
nor U19968 (N_19968,N_13105,N_14840);
nor U19969 (N_19969,N_13458,N_12739);
nor U19970 (N_19970,N_10447,N_13451);
nand U19971 (N_19971,N_14683,N_11229);
nor U19972 (N_19972,N_11270,N_13188);
and U19973 (N_19973,N_14286,N_14177);
or U19974 (N_19974,N_12023,N_13603);
and U19975 (N_19975,N_13799,N_11214);
nand U19976 (N_19976,N_11769,N_10979);
nor U19977 (N_19977,N_13836,N_10303);
and U19978 (N_19978,N_10194,N_14043);
nand U19979 (N_19979,N_13270,N_13030);
nor U19980 (N_19980,N_11110,N_11175);
or U19981 (N_19981,N_13156,N_11955);
nand U19982 (N_19982,N_10248,N_12404);
and U19983 (N_19983,N_12461,N_14895);
nor U19984 (N_19984,N_12531,N_12336);
nand U19985 (N_19985,N_11273,N_11667);
nor U19986 (N_19986,N_14304,N_10218);
nand U19987 (N_19987,N_13053,N_14094);
xor U19988 (N_19988,N_13009,N_13337);
nand U19989 (N_19989,N_12285,N_10019);
and U19990 (N_19990,N_11381,N_13804);
nor U19991 (N_19991,N_11171,N_12217);
and U19992 (N_19992,N_10093,N_11293);
nand U19993 (N_19993,N_14415,N_11808);
and U19994 (N_19994,N_10407,N_11649);
nand U19995 (N_19995,N_14254,N_14984);
and U19996 (N_19996,N_13273,N_14944);
nand U19997 (N_19997,N_13372,N_13361);
and U19998 (N_19998,N_13180,N_11063);
and U19999 (N_19999,N_12373,N_14744);
or UO_0 (O_0,N_16068,N_15123);
nand UO_1 (O_1,N_16123,N_17774);
and UO_2 (O_2,N_19561,N_18496);
nor UO_3 (O_3,N_17385,N_18592);
nand UO_4 (O_4,N_15838,N_19708);
or UO_5 (O_5,N_15917,N_19462);
and UO_6 (O_6,N_18628,N_19446);
or UO_7 (O_7,N_17225,N_15555);
or UO_8 (O_8,N_16987,N_19823);
nand UO_9 (O_9,N_19623,N_16568);
nand UO_10 (O_10,N_15837,N_15736);
nand UO_11 (O_11,N_17358,N_16795);
nand UO_12 (O_12,N_17512,N_15598);
nor UO_13 (O_13,N_15044,N_15621);
and UO_14 (O_14,N_18549,N_15546);
and UO_15 (O_15,N_19893,N_17172);
nand UO_16 (O_16,N_18754,N_15386);
or UO_17 (O_17,N_15881,N_19532);
and UO_18 (O_18,N_16133,N_16562);
and UO_19 (O_19,N_17231,N_17042);
or UO_20 (O_20,N_19171,N_16408);
and UO_21 (O_21,N_18387,N_19923);
nand UO_22 (O_22,N_17612,N_15325);
nand UO_23 (O_23,N_19678,N_19688);
nor UO_24 (O_24,N_19494,N_17443);
nand UO_25 (O_25,N_15474,N_15094);
and UO_26 (O_26,N_15814,N_15345);
nand UO_27 (O_27,N_19890,N_17088);
or UO_28 (O_28,N_19151,N_15657);
and UO_29 (O_29,N_16625,N_16648);
nor UO_30 (O_30,N_16375,N_18283);
nand UO_31 (O_31,N_15296,N_15456);
nand UO_32 (O_32,N_19711,N_15284);
or UO_33 (O_33,N_15161,N_15676);
or UO_34 (O_34,N_19249,N_19858);
nor UO_35 (O_35,N_16790,N_16907);
or UO_36 (O_36,N_15844,N_18260);
and UO_37 (O_37,N_19056,N_16362);
or UO_38 (O_38,N_16727,N_19605);
nor UO_39 (O_39,N_15693,N_19182);
nand UO_40 (O_40,N_19727,N_16631);
and UO_41 (O_41,N_16360,N_19029);
nand UO_42 (O_42,N_18012,N_17335);
nor UO_43 (O_43,N_16837,N_18282);
and UO_44 (O_44,N_16298,N_15246);
and UO_45 (O_45,N_19503,N_19864);
and UO_46 (O_46,N_18824,N_16311);
and UO_47 (O_47,N_18925,N_17145);
and UO_48 (O_48,N_19598,N_16176);
nor UO_49 (O_49,N_16682,N_19633);
nand UO_50 (O_50,N_16555,N_19108);
nor UO_51 (O_51,N_15504,N_17921);
nor UO_52 (O_52,N_17851,N_18704);
and UO_53 (O_53,N_18511,N_18054);
nor UO_54 (O_54,N_15453,N_16368);
nand UO_55 (O_55,N_17028,N_19048);
and UO_56 (O_56,N_16300,N_17157);
nand UO_57 (O_57,N_17895,N_15348);
nor UO_58 (O_58,N_15304,N_17303);
nor UO_59 (O_59,N_15472,N_15965);
and UO_60 (O_60,N_15997,N_15822);
or UO_61 (O_61,N_18993,N_18093);
nor UO_62 (O_62,N_15212,N_16819);
nand UO_63 (O_63,N_15600,N_15198);
nand UO_64 (O_64,N_18558,N_17782);
nand UO_65 (O_65,N_18077,N_18867);
nor UO_66 (O_66,N_17486,N_16764);
or UO_67 (O_67,N_16023,N_15203);
nand UO_68 (O_68,N_17993,N_18419);
nor UO_69 (O_69,N_19081,N_17841);
or UO_70 (O_70,N_18882,N_16499);
nor UO_71 (O_71,N_19447,N_16855);
nor UO_72 (O_72,N_19519,N_15960);
xor UO_73 (O_73,N_15433,N_17577);
nor UO_74 (O_74,N_18380,N_16827);
and UO_75 (O_75,N_16915,N_16219);
and UO_76 (O_76,N_15383,N_18618);
or UO_77 (O_77,N_17757,N_18295);
and UO_78 (O_78,N_17448,N_17215);
nor UO_79 (O_79,N_15556,N_15860);
or UO_80 (O_80,N_19964,N_15309);
nor UO_81 (O_81,N_17917,N_16378);
or UO_82 (O_82,N_19386,N_17123);
or UO_83 (O_83,N_17384,N_17827);
or UO_84 (O_84,N_17437,N_15595);
nand UO_85 (O_85,N_15671,N_19536);
nand UO_86 (O_86,N_18251,N_17656);
nor UO_87 (O_87,N_18021,N_15479);
nand UO_88 (O_88,N_17425,N_18798);
and UO_89 (O_89,N_19988,N_16725);
nand UO_90 (O_90,N_18846,N_15624);
nand UO_91 (O_91,N_17732,N_19908);
and UO_92 (O_92,N_15627,N_18414);
or UO_93 (O_93,N_17901,N_19839);
nand UO_94 (O_94,N_15957,N_15031);
and UO_95 (O_95,N_18017,N_18660);
or UO_96 (O_96,N_15353,N_16352);
nand UO_97 (O_97,N_17666,N_16692);
nor UO_98 (O_98,N_19847,N_19990);
and UO_99 (O_99,N_19251,N_15443);
nand UO_100 (O_100,N_15679,N_18930);
nor UO_101 (O_101,N_19981,N_16472);
nand UO_102 (O_102,N_19947,N_18536);
or UO_103 (O_103,N_17083,N_15717);
or UO_104 (O_104,N_18743,N_17814);
nand UO_105 (O_105,N_18935,N_17012);
and UO_106 (O_106,N_18574,N_15232);
and UO_107 (O_107,N_15154,N_18098);
and UO_108 (O_108,N_16025,N_15109);
or UO_109 (O_109,N_18449,N_17371);
nand UO_110 (O_110,N_19467,N_18774);
nand UO_111 (O_111,N_15520,N_15145);
nor UO_112 (O_112,N_16044,N_16397);
nor UO_113 (O_113,N_16338,N_18421);
or UO_114 (O_114,N_19816,N_19911);
and UO_115 (O_115,N_16815,N_16245);
and UO_116 (O_116,N_15097,N_19828);
nor UO_117 (O_117,N_16047,N_17957);
nor UO_118 (O_118,N_17558,N_18318);
and UO_119 (O_119,N_17529,N_15892);
nand UO_120 (O_120,N_16112,N_17220);
nor UO_121 (O_121,N_17079,N_16026);
and UO_122 (O_122,N_19231,N_16657);
xor UO_123 (O_123,N_16564,N_18290);
nand UO_124 (O_124,N_17155,N_16593);
or UO_125 (O_125,N_19228,N_16763);
nor UO_126 (O_126,N_17379,N_17580);
or UO_127 (O_127,N_16936,N_19229);
or UO_128 (O_128,N_19872,N_18241);
nor UO_129 (O_129,N_18783,N_18550);
nand UO_130 (O_130,N_19498,N_18719);
nor UO_131 (O_131,N_19651,N_18941);
and UO_132 (O_132,N_15698,N_16822);
and UO_133 (O_133,N_17680,N_19546);
and UO_134 (O_134,N_17572,N_17600);
nand UO_135 (O_135,N_18502,N_19366);
or UO_136 (O_136,N_16921,N_18084);
nor UO_137 (O_137,N_18636,N_15082);
nand UO_138 (O_138,N_19009,N_16859);
or UO_139 (O_139,N_17941,N_18028);
and UO_140 (O_140,N_17234,N_18321);
and UO_141 (O_141,N_16152,N_17184);
nand UO_142 (O_142,N_16367,N_19523);
and UO_143 (O_143,N_18067,N_16899);
and UO_144 (O_144,N_15707,N_17620);
nor UO_145 (O_145,N_16970,N_18631);
nor UO_146 (O_146,N_15511,N_19756);
and UO_147 (O_147,N_15491,N_16503);
or UO_148 (O_148,N_18906,N_17775);
nand UO_149 (O_149,N_15942,N_17866);
nand UO_150 (O_150,N_17690,N_16779);
nor UO_151 (O_151,N_16677,N_17206);
nor UO_152 (O_152,N_19132,N_16228);
xor UO_153 (O_153,N_16869,N_18855);
nor UO_154 (O_154,N_16542,N_16616);
nand UO_155 (O_155,N_19738,N_15642);
nand UO_156 (O_156,N_19423,N_19272);
or UO_157 (O_157,N_15823,N_17167);
nand UO_158 (O_158,N_15393,N_17203);
or UO_159 (O_159,N_19513,N_15066);
and UO_160 (O_160,N_19206,N_16086);
or UO_161 (O_161,N_16350,N_17763);
nor UO_162 (O_162,N_18126,N_18371);
and UO_163 (O_163,N_15124,N_15761);
and UO_164 (O_164,N_17561,N_18864);
nor UO_165 (O_165,N_19754,N_16414);
or UO_166 (O_166,N_17034,N_16178);
and UO_167 (O_167,N_16106,N_19359);
nand UO_168 (O_168,N_19715,N_19665);
and UO_169 (O_169,N_19175,N_16642);
nand UO_170 (O_170,N_15974,N_17038);
and UO_171 (O_171,N_16076,N_16359);
and UO_172 (O_172,N_15062,N_19010);
and UO_173 (O_173,N_16247,N_15078);
and UO_174 (O_174,N_17254,N_18398);
nor UO_175 (O_175,N_15297,N_19892);
nand UO_176 (O_176,N_19552,N_19607);
or UO_177 (O_177,N_19232,N_15128);
and UO_178 (O_178,N_15253,N_15160);
or UO_179 (O_179,N_16536,N_18812);
nor UO_180 (O_180,N_19028,N_15603);
nand UO_181 (O_181,N_18438,N_15730);
and UO_182 (O_182,N_16759,N_17228);
or UO_183 (O_183,N_16002,N_17191);
nand UO_184 (O_184,N_17696,N_18689);
or UO_185 (O_185,N_18988,N_16433);
nand UO_186 (O_186,N_15057,N_18199);
and UO_187 (O_187,N_18471,N_17352);
nor UO_188 (O_188,N_17129,N_16250);
or UO_189 (O_189,N_19138,N_18327);
and UO_190 (O_190,N_16190,N_15139);
and UO_191 (O_191,N_17938,N_17699);
and UO_192 (O_192,N_17534,N_16212);
nand UO_193 (O_193,N_16854,N_19619);
nor UO_194 (O_194,N_15011,N_18816);
or UO_195 (O_195,N_17216,N_16128);
and UO_196 (O_196,N_17758,N_17170);
or UO_197 (O_197,N_15898,N_17090);
nor UO_198 (O_198,N_19578,N_17240);
nand UO_199 (O_199,N_17647,N_16556);
and UO_200 (O_200,N_19308,N_18477);
or UO_201 (O_201,N_18141,N_15702);
nand UO_202 (O_202,N_19874,N_17826);
nor UO_203 (O_203,N_15508,N_16448);
and UO_204 (O_204,N_16345,N_15445);
or UO_205 (O_205,N_18480,N_19174);
or UO_206 (O_206,N_18825,N_17188);
and UO_207 (O_207,N_18364,N_18587);
nand UO_208 (O_208,N_17608,N_19710);
or UO_209 (O_209,N_18270,N_16947);
and UO_210 (O_210,N_18742,N_18157);
nand UO_211 (O_211,N_18722,N_17973);
or UO_212 (O_212,N_19415,N_16806);
and UO_213 (O_213,N_19608,N_19095);
nor UO_214 (O_214,N_16811,N_17196);
nor UO_215 (O_215,N_18542,N_16391);
or UO_216 (O_216,N_17791,N_15442);
and UO_217 (O_217,N_19969,N_15537);
or UO_218 (O_218,N_18728,N_17786);
nor UO_219 (O_219,N_15426,N_15695);
or UO_220 (O_220,N_17771,N_19723);
nand UO_221 (O_221,N_16505,N_17421);
nor UO_222 (O_222,N_16817,N_19783);
or UO_223 (O_223,N_15735,N_18795);
nor UO_224 (O_224,N_15008,N_15867);
or UO_225 (O_225,N_17644,N_16363);
and UO_226 (O_226,N_19420,N_17236);
nand UO_227 (O_227,N_16195,N_15009);
and UO_228 (O_228,N_16485,N_15899);
nand UO_229 (O_229,N_16193,N_19504);
or UO_230 (O_230,N_19920,N_17544);
nor UO_231 (O_231,N_17549,N_16316);
nor UO_232 (O_232,N_15397,N_19841);
or UO_233 (O_233,N_15184,N_19378);
nand UO_234 (O_234,N_18853,N_15054);
and UO_235 (O_235,N_16614,N_17970);
nor UO_236 (O_236,N_16846,N_17643);
or UO_237 (O_237,N_19904,N_19616);
or UO_238 (O_238,N_18443,N_19334);
nor UO_239 (O_239,N_19398,N_15968);
and UO_240 (O_240,N_18643,N_17756);
nand UO_241 (O_241,N_17395,N_18350);
and UO_242 (O_242,N_18200,N_18514);
nand UO_243 (O_243,N_15638,N_17397);
nor UO_244 (O_244,N_19838,N_19840);
nand UO_245 (O_245,N_18959,N_18595);
and UO_246 (O_246,N_15843,N_16005);
nor UO_247 (O_247,N_15204,N_16490);
and UO_248 (O_248,N_15694,N_18810);
nor UO_249 (O_249,N_16781,N_15469);
nor UO_250 (O_250,N_16425,N_18073);
nand UO_251 (O_251,N_16634,N_17165);
nand UO_252 (O_252,N_18361,N_18366);
nand UO_253 (O_253,N_18437,N_17905);
or UO_254 (O_254,N_18478,N_15873);
and UO_255 (O_255,N_15356,N_18917);
and UO_256 (O_256,N_15220,N_19256);
or UO_257 (O_257,N_16778,N_19945);
nand UO_258 (O_258,N_16856,N_17072);
nand UO_259 (O_259,N_18580,N_19648);
and UO_260 (O_260,N_18777,N_15288);
nor UO_261 (O_261,N_15940,N_18405);
and UO_262 (O_262,N_15678,N_18519);
and UO_263 (O_263,N_16398,N_16435);
or UO_264 (O_264,N_19127,N_16624);
nand UO_265 (O_265,N_15135,N_19271);
nand UO_266 (O_266,N_18138,N_18064);
and UO_267 (O_267,N_18927,N_16723);
and UO_268 (O_268,N_16515,N_18785);
and UO_269 (O_269,N_18258,N_18145);
nor UO_270 (O_270,N_19167,N_17609);
nor UO_271 (O_271,N_17710,N_19338);
or UO_272 (O_272,N_18139,N_16407);
nand UO_273 (O_273,N_16701,N_19163);
or UO_274 (O_274,N_17306,N_19038);
and UO_275 (O_275,N_16775,N_19291);
nand UO_276 (O_276,N_15579,N_17502);
or UO_277 (O_277,N_18828,N_15774);
and UO_278 (O_278,N_17844,N_15853);
nor UO_279 (O_279,N_18302,N_15835);
or UO_280 (O_280,N_16691,N_16931);
nand UO_281 (O_281,N_16438,N_15883);
or UO_282 (O_282,N_15271,N_17117);
nand UO_283 (O_283,N_15489,N_15709);
and UO_284 (O_284,N_17366,N_16709);
or UO_285 (O_285,N_16920,N_17825);
nor UO_286 (O_286,N_16347,N_16379);
nor UO_287 (O_287,N_15257,N_17388);
nor UO_288 (O_288,N_17845,N_16153);
or UO_289 (O_289,N_19321,N_19744);
nor UO_290 (O_290,N_18717,N_15497);
nor UO_291 (O_291,N_18630,N_19012);
nor UO_292 (O_292,N_19413,N_18588);
and UO_293 (O_293,N_19758,N_19070);
nand UO_294 (O_294,N_17013,N_16999);
and UO_295 (O_295,N_19582,N_15685);
nand UO_296 (O_296,N_19279,N_16813);
or UO_297 (O_297,N_17725,N_19343);
or UO_298 (O_298,N_16538,N_16240);
nor UO_299 (O_299,N_15112,N_15742);
nor UO_300 (O_300,N_15850,N_15071);
or UO_301 (O_301,N_16405,N_17007);
or UO_302 (O_302,N_16879,N_17682);
and UO_303 (O_303,N_15310,N_16617);
nand UO_304 (O_304,N_15586,N_16157);
and UO_305 (O_305,N_17991,N_19897);
nand UO_306 (O_306,N_16891,N_18512);
or UO_307 (O_307,N_18726,N_15982);
and UO_308 (O_308,N_15434,N_15366);
and UO_309 (O_309,N_15306,N_16985);
and UO_310 (O_310,N_18344,N_15795);
or UO_311 (O_311,N_17711,N_15408);
nand UO_312 (O_312,N_19703,N_19815);
and UO_313 (O_313,N_19778,N_15248);
or UO_314 (O_314,N_15983,N_19869);
and UO_315 (O_315,N_18695,N_18184);
nor UO_316 (O_316,N_17359,N_16188);
nand UO_317 (O_317,N_15688,N_19062);
nor UO_318 (O_318,N_18040,N_16605);
or UO_319 (O_319,N_15049,N_15745);
nor UO_320 (O_320,N_16623,N_16808);
nor UO_321 (O_321,N_17438,N_16635);
nand UO_322 (O_322,N_17390,N_19496);
or UO_323 (O_323,N_17653,N_19912);
or UO_324 (O_324,N_19829,N_15074);
and UO_325 (O_325,N_17361,N_19166);
or UO_326 (O_326,N_16863,N_15151);
nor UO_327 (O_327,N_19800,N_18349);
and UO_328 (O_328,N_18818,N_15649);
nor UO_329 (O_329,N_16475,N_15592);
or UO_330 (O_330,N_18446,N_15557);
nand UO_331 (O_331,N_17717,N_19773);
and UO_332 (O_332,N_17838,N_15105);
and UO_333 (O_333,N_16473,N_16736);
nor UO_334 (O_334,N_18222,N_15585);
nand UO_335 (O_335,N_16599,N_15374);
or UO_336 (O_336,N_16658,N_17927);
nand UO_337 (O_337,N_17551,N_18155);
nand UO_338 (O_338,N_18649,N_17280);
or UO_339 (O_339,N_16698,N_18950);
nor UO_340 (O_340,N_16753,N_17279);
nand UO_341 (O_341,N_19719,N_19385);
nor UO_342 (O_342,N_19451,N_15714);
or UO_343 (O_343,N_19159,N_19377);
and UO_344 (O_344,N_18790,N_16258);
or UO_345 (O_345,N_17916,N_17897);
or UO_346 (O_346,N_18577,N_19919);
or UO_347 (O_347,N_17963,N_18460);
and UO_348 (O_348,N_15089,N_15133);
or UO_349 (O_349,N_16847,N_17598);
nand UO_350 (O_350,N_19674,N_18658);
or UO_351 (O_351,N_19954,N_19025);
and UO_352 (O_352,N_15087,N_17484);
or UO_353 (O_353,N_17546,N_16539);
or UO_354 (O_354,N_15068,N_18887);
nor UO_355 (O_355,N_16576,N_18195);
nor UO_356 (O_356,N_15267,N_17355);
nand UO_357 (O_357,N_17799,N_17198);
nand UO_358 (O_358,N_19922,N_17103);
nor UO_359 (O_359,N_15211,N_19131);
nand UO_360 (O_360,N_18926,N_18936);
nand UO_361 (O_361,N_17487,N_17144);
nor UO_362 (O_362,N_17902,N_17573);
or UO_363 (O_363,N_18500,N_19208);
or UO_364 (O_364,N_17089,N_16321);
nor UO_365 (O_365,N_16954,N_18412);
or UO_366 (O_366,N_19495,N_19746);
and UO_367 (O_367,N_18890,N_15549);
nand UO_368 (O_368,N_19520,N_16961);
nand UO_369 (O_369,N_16988,N_18561);
nor UO_370 (O_370,N_19280,N_17816);
nor UO_371 (O_371,N_15575,N_19512);
nand UO_372 (O_372,N_19573,N_19772);
or UO_373 (O_373,N_17006,N_18188);
or UO_374 (O_374,N_16618,N_15423);
or UO_375 (O_375,N_17942,N_19960);
and UO_376 (O_376,N_19417,N_16085);
nand UO_377 (O_377,N_18038,N_17033);
and UO_378 (O_378,N_16209,N_19455);
and UO_379 (O_379,N_17019,N_17979);
nor UO_380 (O_380,N_19088,N_19568);
nand UO_381 (O_381,N_16637,N_18978);
or UO_382 (O_382,N_16489,N_18505);
nand UO_383 (O_383,N_16877,N_16783);
or UO_384 (O_384,N_19917,N_17187);
or UO_385 (O_385,N_17798,N_18434);
nor UO_386 (O_386,N_15941,N_18980);
and UO_387 (O_387,N_18457,N_16826);
or UO_388 (O_388,N_17663,N_16802);
or UO_389 (O_389,N_18183,N_19528);
nand UO_390 (O_390,N_19460,N_15395);
nand UO_391 (O_391,N_15692,N_18730);
or UO_392 (O_392,N_18305,N_16122);
and UO_393 (O_393,N_15530,N_15780);
and UO_394 (O_394,N_19325,N_17108);
or UO_395 (O_395,N_19690,N_18900);
or UO_396 (O_396,N_15744,N_16421);
or UO_397 (O_397,N_15849,N_17417);
nand UO_398 (O_398,N_16067,N_17273);
nand UO_399 (O_399,N_16010,N_18019);
and UO_400 (O_400,N_16261,N_17436);
nor UO_401 (O_401,N_17550,N_19720);
or UO_402 (O_402,N_19946,N_15322);
nand UO_403 (O_403,N_17407,N_16332);
and UO_404 (O_404,N_15137,N_17192);
nand UO_405 (O_405,N_19312,N_18875);
nor UO_406 (O_406,N_18203,N_17064);
and UO_407 (O_407,N_19937,N_15975);
nand UO_408 (O_408,N_19364,N_18897);
and UO_409 (O_409,N_17541,N_17607);
and UO_410 (O_410,N_19968,N_18032);
nand UO_411 (O_411,N_15483,N_17208);
and UO_412 (O_412,N_18607,N_16716);
nor UO_413 (O_413,N_17300,N_17347);
nand UO_414 (O_414,N_17101,N_19692);
or UO_415 (O_415,N_16744,N_18007);
or UO_416 (O_416,N_19384,N_16581);
and UO_417 (O_417,N_17634,N_19372);
and UO_418 (O_418,N_18947,N_17059);
or UO_419 (O_419,N_17937,N_17950);
nor UO_420 (O_420,N_17483,N_16787);
nor UO_421 (O_421,N_19168,N_18298);
and UO_422 (O_422,N_16487,N_15613);
and UO_423 (O_423,N_15513,N_16038);
and UO_424 (O_424,N_16833,N_17376);
or UO_425 (O_425,N_16700,N_15132);
nor UO_426 (O_426,N_15093,N_16339);
and UO_427 (O_427,N_17207,N_17336);
nand UO_428 (O_428,N_15858,N_17285);
nand UO_429 (O_429,N_19843,N_16181);
nor UO_430 (O_430,N_16979,N_17780);
nand UO_431 (O_431,N_16655,N_19531);
nor UO_432 (O_432,N_19331,N_17375);
nor UO_433 (O_433,N_17183,N_18583);
nand UO_434 (O_434,N_19775,N_15070);
nand UO_435 (O_435,N_17724,N_16860);
or UO_436 (O_436,N_19534,N_18527);
and UO_437 (O_437,N_15228,N_16455);
nor UO_438 (O_438,N_18310,N_17731);
and UO_439 (O_439,N_16197,N_16317);
nor UO_440 (O_440,N_19313,N_19296);
and UO_441 (O_441,N_15162,N_17314);
and UO_442 (O_442,N_16051,N_17507);
nand UO_443 (O_443,N_19706,N_19091);
nand UO_444 (O_444,N_19476,N_16675);
and UO_445 (O_445,N_16201,N_19030);
nand UO_446 (O_446,N_19885,N_17383);
nor UO_447 (O_447,N_19612,N_18787);
nor UO_448 (O_448,N_19553,N_17433);
or UO_449 (O_449,N_19871,N_18657);
or UO_450 (O_450,N_19555,N_17186);
and UO_451 (O_451,N_19222,N_15373);
or UO_452 (O_452,N_17247,N_18154);
nor UO_453 (O_453,N_17290,N_18422);
nor UO_454 (O_454,N_16517,N_15174);
and UO_455 (O_455,N_17224,N_19736);
and UO_456 (O_456,N_19647,N_18212);
and UO_457 (O_457,N_17233,N_16294);
nand UO_458 (O_458,N_16647,N_15864);
nand UO_459 (O_459,N_16450,N_16114);
nand UO_460 (O_460,N_17065,N_16057);
or UO_461 (O_461,N_17565,N_19146);
or UO_462 (O_462,N_16230,N_17147);
and UO_463 (O_463,N_18360,N_16602);
nor UO_464 (O_464,N_17069,N_19907);
nand UO_465 (O_465,N_15784,N_18150);
and UO_466 (O_466,N_16745,N_15358);
nor UO_467 (O_467,N_16981,N_16966);
or UO_468 (O_468,N_18644,N_17521);
nor UO_469 (O_469,N_18475,N_19486);
and UO_470 (O_470,N_18257,N_15757);
nand UO_471 (O_471,N_15043,N_17381);
or UO_472 (O_472,N_17779,N_16402);
and UO_473 (O_473,N_15428,N_16075);
nor UO_474 (O_474,N_19258,N_15039);
nor UO_475 (O_475,N_15064,N_15811);
nor UO_476 (O_476,N_18602,N_18441);
nand UO_477 (O_477,N_15216,N_17043);
and UO_478 (O_478,N_17880,N_15399);
nor UO_479 (O_479,N_18319,N_16020);
and UO_480 (O_480,N_16284,N_18322);
or UO_481 (O_481,N_16477,N_19630);
or UO_482 (O_482,N_19626,N_19787);
nand UO_483 (O_483,N_17091,N_18807);
and UO_484 (O_484,N_15376,N_19564);
and UO_485 (O_485,N_16458,N_15010);
nor UO_486 (O_486,N_16340,N_17316);
and UO_487 (O_487,N_18665,N_15003);
nor UO_488 (O_488,N_17560,N_18079);
nand UO_489 (O_489,N_16953,N_15498);
nor UO_490 (O_490,N_15460,N_18884);
or UO_491 (O_491,N_15545,N_16563);
or UO_492 (O_492,N_17781,N_15805);
and UO_493 (O_493,N_15697,N_16441);
nand UO_494 (O_494,N_18244,N_17721);
nor UO_495 (O_495,N_19395,N_19197);
or UO_496 (O_496,N_17299,N_15169);
nand UO_497 (O_497,N_18370,N_17804);
nor UO_498 (O_498,N_17085,N_18202);
nor UO_499 (O_499,N_15930,N_15462);
or UO_500 (O_500,N_18140,N_17773);
nor UO_501 (O_501,N_15650,N_18768);
and UO_502 (O_502,N_15653,N_19218);
or UO_503 (O_503,N_16356,N_17641);
or UO_504 (O_504,N_16027,N_16690);
nand UO_505 (O_505,N_16537,N_19219);
nand UO_506 (O_506,N_17931,N_17002);
and UO_507 (O_507,N_16208,N_16079);
or UO_508 (O_508,N_18381,N_15193);
nor UO_509 (O_509,N_18530,N_18840);
and UO_510 (O_510,N_17618,N_17327);
or UO_511 (O_511,N_19382,N_19429);
or UO_512 (O_512,N_15027,N_15173);
nor UO_513 (O_513,N_16858,N_18292);
nor UO_514 (O_514,N_17199,N_18190);
nor UO_515 (O_515,N_16192,N_15086);
nor UO_516 (O_516,N_15851,N_16509);
nor UO_517 (O_517,N_18492,N_17205);
and UO_518 (O_518,N_19204,N_15894);
nand UO_519 (O_519,N_19935,N_15943);
or UO_520 (O_520,N_15775,N_19924);
nand UO_521 (O_521,N_18969,N_15833);
nand UO_522 (O_522,N_16922,N_16371);
nand UO_523 (O_523,N_19664,N_19567);
or UO_524 (O_524,N_16520,N_15791);
nor UO_525 (O_525,N_19147,N_17239);
nand UO_526 (O_526,N_17967,N_15308);
or UO_527 (O_527,N_16622,N_18096);
and UO_528 (O_528,N_18357,N_19562);
nor UO_529 (O_529,N_18097,N_17989);
and UO_530 (O_530,N_19047,N_19414);
nand UO_531 (O_531,N_17025,N_15007);
or UO_532 (O_532,N_15401,N_19779);
or UO_533 (O_533,N_17073,N_17867);
and UO_534 (O_534,N_19879,N_17542);
and UO_535 (O_535,N_18430,N_16793);
or UO_536 (O_536,N_18033,N_19604);
nor UO_537 (O_537,N_19263,N_16059);
nand UO_538 (O_538,N_16031,N_18559);
or UO_539 (O_539,N_16333,N_16377);
and UO_540 (O_540,N_18876,N_15130);
or UO_541 (O_541,N_16540,N_15562);
or UO_542 (O_542,N_15492,N_15413);
nor UO_543 (O_543,N_18573,N_17708);
or UO_544 (O_544,N_16668,N_18481);
and UO_545 (O_545,N_18235,N_18210);
and UO_546 (O_546,N_18613,N_15721);
nand UO_547 (O_547,N_15655,N_15646);
nand UO_548 (O_548,N_15282,N_19794);
nand UO_549 (O_549,N_18211,N_15716);
nor UO_550 (O_550,N_19973,N_15236);
nand UO_551 (O_551,N_18132,N_16324);
nor UO_552 (O_552,N_19215,N_19225);
or UO_553 (O_553,N_17513,N_15990);
or UO_554 (O_554,N_17175,N_15857);
nand UO_555 (O_555,N_15380,N_16275);
nand UO_556 (O_556,N_15118,N_17338);
or UO_557 (O_557,N_17664,N_18656);
and UO_558 (O_558,N_17720,N_19276);
nor UO_559 (O_559,N_18453,N_18997);
nor UO_560 (O_560,N_18690,N_18025);
nand UO_561 (O_561,N_17538,N_16268);
or UO_562 (O_562,N_19090,N_15647);
or UO_563 (O_563,N_19315,N_19732);
nand UO_564 (O_564,N_19658,N_15452);
nor UO_565 (O_565,N_15280,N_16717);
or UO_566 (O_566,N_16444,N_15724);
and UO_567 (O_567,N_15015,N_18506);
or UO_568 (O_568,N_15708,N_15321);
xor UO_569 (O_569,N_15063,N_15856);
nor UO_570 (O_570,N_17559,N_15327);
and UO_571 (O_571,N_19896,N_18130);
nor UO_572 (O_572,N_19461,N_19100);
nand UO_573 (O_573,N_15909,N_16158);
and UO_574 (O_574,N_19301,N_19199);
and UO_575 (O_575,N_19269,N_17744);
nand UO_576 (O_576,N_16018,N_17980);
and UO_577 (O_577,N_17142,N_17982);
and UO_578 (O_578,N_16882,N_16480);
nand UO_579 (O_579,N_16773,N_16103);
and UO_580 (O_580,N_17463,N_19653);
nand UO_581 (O_581,N_15351,N_18499);
or UO_582 (O_582,N_18539,N_16632);
nor UO_583 (O_583,N_15448,N_15379);
and UO_584 (O_584,N_19404,N_19442);
or UO_585 (O_585,N_16428,N_18720);
nand UO_586 (O_586,N_17959,N_15584);
nand UO_587 (O_587,N_17116,N_16434);
nor UO_588 (O_588,N_18484,N_18232);
nand UO_589 (O_589,N_17289,N_17587);
nand UO_590 (O_590,N_18031,N_17334);
or UO_591 (O_591,N_17194,N_19238);
and UO_592 (O_592,N_15146,N_16714);
or UO_593 (O_593,N_16273,N_16955);
and UO_594 (O_594,N_17621,N_19196);
or UO_595 (O_595,N_18013,N_18023);
nand UO_596 (O_596,N_19143,N_18958);
nand UO_597 (O_597,N_17344,N_17493);
xnor UO_598 (O_598,N_19071,N_18648);
nand UO_599 (O_599,N_19548,N_16403);
nor UO_600 (O_600,N_16728,N_15252);
nand UO_601 (O_601,N_19971,N_18646);
or UO_602 (O_602,N_17702,N_15636);
or UO_603 (O_603,N_17122,N_17026);
nor UO_604 (O_604,N_19045,N_19942);
nor UO_605 (O_605,N_19928,N_19195);
or UO_606 (O_606,N_18131,N_18326);
nor UO_607 (O_607,N_15040,N_18348);
nand UO_608 (O_608,N_17987,N_16236);
or UO_609 (O_609,N_17996,N_16529);
or UO_610 (O_610,N_17353,N_16665);
and UO_611 (O_611,N_17671,N_16415);
nor UO_612 (O_612,N_16547,N_16383);
and UO_613 (O_613,N_18336,N_17251);
or UO_614 (O_614,N_18470,N_15770);
or UO_615 (O_615,N_15669,N_17934);
nor UO_616 (O_616,N_18329,N_16182);
nand UO_617 (O_617,N_19116,N_17741);
xnor UO_618 (O_618,N_16831,N_15108);
nand UO_619 (O_619,N_17354,N_16670);
or UO_620 (O_620,N_19286,N_17946);
nor UO_621 (O_621,N_17315,N_18147);
and UO_622 (O_622,N_17181,N_19551);
and UO_623 (O_623,N_16949,N_16770);
nor UO_624 (O_624,N_16767,N_19165);
nand UO_625 (O_625,N_17249,N_16227);
nand UO_626 (O_626,N_16975,N_19424);
or UO_627 (O_627,N_17442,N_18061);
and UO_628 (O_628,N_17282,N_16263);
or UO_629 (O_629,N_15432,N_19625);
or UO_630 (O_630,N_17174,N_16260);
or UO_631 (O_631,N_18307,N_19054);
and UO_632 (O_632,N_15659,N_16307);
or UO_633 (O_633,N_19187,N_16366);
nand UO_634 (O_634,N_17179,N_18273);
or UO_635 (O_635,N_17037,N_17270);
or UO_636 (O_636,N_15266,N_17268);
nor UO_637 (O_637,N_16829,N_17488);
nor UO_638 (O_638,N_15768,N_19832);
or UO_639 (O_639,N_15680,N_16501);
nor UO_640 (O_640,N_16436,N_18827);
nor UO_641 (O_641,N_16894,N_18036);
nand UO_642 (O_642,N_15166,N_19522);
nand UO_643 (O_643,N_17557,N_18538);
nand UO_644 (O_644,N_17326,N_19376);
and UO_645 (O_645,N_19844,N_18564);
xnor UO_646 (O_646,N_17755,N_17195);
nor UO_647 (O_647,N_15470,N_19852);
or UO_648 (O_648,N_15229,N_19011);
nand UO_649 (O_649,N_17466,N_18885);
and UO_650 (O_650,N_19729,N_17855);
and UO_651 (O_651,N_17005,N_19768);
and UO_652 (O_652,N_18008,N_17302);
nand UO_653 (O_653,N_18953,N_18928);
and UO_654 (O_654,N_15620,N_17795);
nand UO_655 (O_655,N_18761,N_18046);
or UO_656 (O_656,N_19324,N_15859);
and UO_657 (O_657,N_16121,N_17614);
nor UO_658 (O_658,N_17377,N_18233);
and UO_659 (O_659,N_16012,N_16823);
or UO_660 (O_660,N_18035,N_18390);
or UO_661 (O_661,N_17943,N_18863);
nand UO_662 (O_662,N_15467,N_19481);
nand UO_663 (O_663,N_17271,N_18584);
or UO_664 (O_664,N_16288,N_16610);
and UO_665 (O_665,N_17015,N_17528);
or UO_666 (O_666,N_18526,N_18240);
and UO_667 (O_667,N_19705,N_19584);
nor UO_668 (O_668,N_18214,N_19214);
nor UO_669 (O_669,N_18889,N_15163);
and UO_670 (O_670,N_17579,N_19408);
nor UO_671 (O_671,N_19643,N_18975);
nand UO_672 (O_672,N_16934,N_17923);
and UO_673 (O_673,N_15258,N_15606);
or UO_674 (O_674,N_15444,N_15360);
nor UO_675 (O_675,N_19614,N_18468);
and UO_676 (O_676,N_16334,N_18727);
nor UO_677 (O_677,N_15152,N_18923);
nand UO_678 (O_678,N_19371,N_15301);
or UO_679 (O_679,N_18714,N_17440);
and UO_680 (O_680,N_19975,N_17903);
nor UO_681 (O_681,N_17962,N_16429);
nor UO_682 (O_682,N_15269,N_16636);
or UO_683 (O_683,N_18284,N_16748);
nor UO_684 (O_684,N_16619,N_19212);
and UO_685 (O_685,N_19484,N_18776);
and UO_686 (O_686,N_15989,N_18766);
or UO_687 (O_687,N_18440,N_17633);
nand UO_688 (O_688,N_15713,N_17001);
nor UO_689 (O_689,N_19743,N_17113);
nand UO_690 (O_690,N_15848,N_16303);
or UO_691 (O_691,N_18169,N_19638);
nand UO_692 (O_692,N_19760,N_16382);
nor UO_693 (O_693,N_15904,N_19103);
nor UO_694 (O_694,N_17482,N_17748);
or UO_695 (O_695,N_16596,N_19289);
or UO_696 (O_696,N_18281,N_16980);
or UO_697 (O_697,N_16948,N_19121);
nor UO_698 (O_698,N_17777,N_19040);
nand UO_699 (O_699,N_16687,N_15703);
nor UO_700 (O_700,N_17317,N_17833);
and UO_701 (O_701,N_19808,N_17834);
nor UO_702 (O_702,N_18095,N_17066);
nor UO_703 (O_703,N_17691,N_19083);
or UO_704 (O_704,N_18151,N_17429);
nand UO_705 (O_705,N_15148,N_19391);
and UO_706 (O_706,N_18103,N_19035);
and UO_707 (O_707,N_18059,N_19862);
or UO_708 (O_708,N_19621,N_19317);
or UO_709 (O_709,N_17591,N_17688);
and UO_710 (O_710,N_15018,N_16638);
or UO_711 (O_711,N_16565,N_17133);
nand UO_712 (O_712,N_19644,N_15938);
nor UO_713 (O_713,N_17622,N_18769);
nor UO_714 (O_714,N_19016,N_16290);
nor UO_715 (O_715,N_16828,N_17023);
and UO_716 (O_716,N_19431,N_17998);
and UO_717 (O_717,N_19903,N_18943);
or UO_718 (O_718,N_17457,N_16226);
and UO_719 (O_719,N_16234,N_17652);
or UO_720 (O_720,N_19668,N_19518);
nand UO_721 (O_721,N_16579,N_17555);
or UO_722 (O_722,N_16006,N_17372);
nor UO_723 (O_723,N_17854,N_15392);
nor UO_724 (O_724,N_19834,N_16296);
and UO_725 (O_725,N_17599,N_17726);
or UO_726 (O_726,N_18178,N_15390);
nand UO_727 (O_727,N_15095,N_16984);
nor UO_728 (O_728,N_19043,N_15727);
and UO_729 (O_729,N_16958,N_19769);
nor UO_730 (O_730,N_17859,N_16078);
xor UO_731 (O_731,N_19535,N_16460);
nor UO_732 (O_732,N_19819,N_18065);
nor UO_733 (O_733,N_16865,N_15519);
nand UO_734 (O_734,N_19766,N_16818);
nand UO_735 (O_735,N_19170,N_19683);
nor UO_736 (O_736,N_17891,N_19039);
xnor UO_737 (O_737,N_16660,N_16496);
and UO_738 (O_738,N_18495,N_15218);
or UO_739 (O_739,N_17399,N_19405);
nand UO_740 (O_740,N_19060,N_16091);
nor UO_741 (O_741,N_17713,N_19194);
nand UO_742 (O_742,N_15461,N_19477);
nand UO_743 (O_743,N_18068,N_16730);
or UO_744 (O_744,N_18523,N_16761);
xnor UO_745 (O_745,N_19142,N_16544);
nor UO_746 (O_746,N_18105,N_17197);
nand UO_747 (O_747,N_18991,N_19005);
nand UO_748 (O_748,N_19403,N_19473);
or UO_749 (O_749,N_15357,N_17070);
nand UO_750 (O_750,N_15431,N_18697);
or UO_751 (O_751,N_18731,N_18010);
nor UO_752 (O_752,N_16216,N_18683);
and UO_753 (O_753,N_17000,N_18528);
or UO_754 (O_754,N_17027,N_19655);
nor UO_755 (O_755,N_17067,N_17693);
nand UO_756 (O_756,N_18784,N_17667);
nor UO_757 (O_757,N_17461,N_16174);
nor UO_758 (O_758,N_16591,N_15645);
nand UO_759 (O_759,N_19939,N_17102);
and UO_760 (O_760,N_18881,N_17229);
and UO_761 (O_761,N_18316,N_17926);
or UO_762 (O_762,N_19902,N_16679);
nand UO_763 (O_763,N_17050,N_17956);
or UO_764 (O_764,N_17835,N_19441);
and UO_765 (O_765,N_17506,N_16643);
or UO_766 (O_766,N_15171,N_19262);
or UO_767 (O_767,N_15182,N_17792);
and UO_768 (O_768,N_19330,N_16420);
nand UO_769 (O_769,N_15091,N_15457);
nor UO_770 (O_770,N_17968,N_17110);
or UO_771 (O_771,N_17893,N_15013);
or UO_772 (O_772,N_15237,N_19824);
or UO_773 (O_773,N_19645,N_19537);
nor UO_774 (O_774,N_16328,N_15701);
nand UO_775 (O_775,N_19474,N_16447);
or UO_776 (O_776,N_18677,N_19192);
or UO_777 (O_777,N_18149,N_18226);
and UO_778 (O_778,N_15424,N_18426);
or UO_779 (O_779,N_16184,N_18762);
and UO_780 (O_780,N_19119,N_17508);
xnor UO_781 (O_781,N_17177,N_19875);
nand UO_782 (O_782,N_15531,N_15739);
or UO_783 (O_783,N_18356,N_16718);
or UO_784 (O_784,N_15202,N_15318);
nor UO_785 (O_785,N_15048,N_15566);
or UO_786 (O_786,N_19026,N_17135);
nor UO_787 (O_787,N_19014,N_16302);
nand UO_788 (O_788,N_18119,N_18859);
and UO_789 (O_789,N_15891,N_16521);
nand UO_790 (O_790,N_16257,N_16686);
and UO_791 (O_791,N_18277,N_16992);
and UO_792 (O_792,N_18267,N_16160);
or UO_793 (O_793,N_19191,N_16080);
and UO_794 (O_794,N_16785,N_19041);
or UO_795 (O_795,N_19906,N_15014);
and UO_796 (O_796,N_15937,N_18767);
nor UO_797 (O_797,N_19997,N_19412);
nor UO_798 (O_798,N_19448,N_18562);
and UO_799 (O_799,N_18009,N_15060);
nor UO_800 (O_800,N_19790,N_19635);
nor UO_801 (O_801,N_18858,N_18806);
and UO_802 (O_802,N_17533,N_17811);
nor UO_803 (O_803,N_15931,N_15954);
and UO_804 (O_804,N_18817,N_18027);
and UO_805 (O_805,N_19671,N_19949);
nand UO_806 (O_806,N_17351,N_16862);
nor UO_807 (O_807,N_17759,N_15352);
nor UO_808 (O_808,N_18368,N_17734);
nor UO_809 (O_809,N_19346,N_18729);
or UO_810 (O_810,N_18042,N_15876);
or UO_811 (O_811,N_16265,N_19126);
or UO_812 (O_812,N_15217,N_18990);
nor UO_813 (O_813,N_19470,N_18317);
and UO_814 (O_814,N_16930,N_16645);
nand UO_815 (O_815,N_15346,N_18243);
nand UO_816 (O_816,N_15734,N_19101);
nand UO_817 (O_817,N_17003,N_15387);
nor UO_818 (O_818,N_17350,N_16912);
and UO_819 (O_819,N_18553,N_17460);
and UO_820 (O_820,N_17099,N_17589);
or UO_821 (O_821,N_18451,N_16030);
or UO_822 (O_822,N_16974,N_18454);
and UO_823 (O_823,N_15025,N_17242);
nor UO_824 (O_824,N_16967,N_17817);
nor UO_825 (O_825,N_16532,N_17221);
nor UO_826 (O_826,N_16941,N_16697);
and UO_827 (O_827,N_19594,N_17953);
nor UO_828 (O_828,N_17178,N_17619);
nand UO_829 (O_829,N_17768,N_17872);
or UO_830 (O_830,N_16801,N_19627);
and UO_831 (O_831,N_17272,N_16279);
and UO_832 (O_832,N_18192,N_16782);
nor UO_833 (O_833,N_17427,N_19193);
nand UO_834 (O_834,N_18075,N_17411);
nor UO_835 (O_835,N_19268,N_17878);
and UO_836 (O_836,N_16327,N_18486);
or UO_837 (O_837,N_17406,N_17753);
nand UO_838 (O_838,N_15820,N_15882);
and UO_839 (O_839,N_19777,N_17564);
or UO_840 (O_840,N_19440,N_18782);
nand UO_841 (O_841,N_15998,N_15440);
xnor UO_842 (O_842,N_17097,N_17788);
or UO_843 (O_843,N_19863,N_15633);
and UO_844 (O_844,N_18122,N_17646);
nand UO_845 (O_845,N_17430,N_16722);
or UO_846 (O_846,N_17503,N_16558);
or UO_847 (O_847,N_16577,N_18913);
nand UO_848 (O_848,N_17909,N_18312);
xnor UO_849 (O_849,N_18399,N_15754);
or UO_850 (O_850,N_18117,N_16150);
or UO_851 (O_851,N_15749,N_16463);
nor UO_852 (O_852,N_17930,N_15072);
nor UO_853 (O_853,N_18672,N_18967);
or UO_854 (O_854,N_16644,N_15959);
nor UO_855 (O_855,N_19135,N_18862);
and UO_856 (O_856,N_18497,N_15992);
or UO_857 (O_857,N_19066,N_17389);
and UO_858 (O_858,N_18972,N_16163);
and UO_859 (O_859,N_16445,N_17039);
nand UO_860 (O_860,N_15999,N_18420);
nand UO_861 (O_861,N_18604,N_18715);
or UO_862 (O_862,N_17449,N_15559);
nand UO_863 (O_863,N_18070,N_19064);
and UO_864 (O_864,N_16752,N_17983);
nand UO_865 (O_865,N_16418,N_18764);
or UO_866 (O_866,N_19433,N_16081);
or UO_867 (O_867,N_17246,N_15629);
nand UO_868 (O_868,N_18288,N_19725);
or UO_869 (O_869,N_19245,N_15824);
nor UO_870 (O_870,N_18285,N_16097);
nor UO_871 (O_871,N_16661,N_19401);
nand UO_872 (O_872,N_18759,N_17030);
nand UO_873 (O_873,N_19958,N_15543);
nor UO_874 (O_874,N_18271,N_18334);
and UO_875 (O_875,N_15170,N_18246);
and UO_876 (O_876,N_18166,N_19713);
nor UO_877 (O_877,N_15654,N_15101);
and UO_878 (O_878,N_18191,N_15662);
nand UO_879 (O_879,N_15710,N_15855);
nand UO_880 (O_880,N_17819,N_15933);
nor UO_881 (O_881,N_18205,N_18699);
or UO_882 (O_882,N_17243,N_18264);
nor UO_883 (O_883,N_16353,N_18537);
and UO_884 (O_884,N_18984,N_18351);
or UO_885 (O_885,N_15815,N_19322);
nor UO_886 (O_886,N_16168,N_17202);
nor UO_887 (O_887,N_19125,N_18170);
nand UO_888 (O_888,N_18503,N_19139);
and UO_889 (O_889,N_19201,N_19905);
and UO_890 (O_890,N_17828,N_17797);
nand UO_891 (O_891,N_15962,N_19517);
nand UO_892 (O_892,N_16629,N_15270);
and UO_893 (O_893,N_17789,N_18994);
or UO_894 (O_894,N_19541,N_18745);
nor UO_895 (O_895,N_16694,N_15286);
nand UO_896 (O_896,N_16180,N_15747);
or UO_897 (O_897,N_16065,N_19615);
nor UO_898 (O_898,N_17913,N_15958);
and UO_899 (O_899,N_17997,N_18324);
nand UO_900 (O_900,N_15922,N_15578);
nand UO_901 (O_901,N_16125,N_17412);
nand UO_902 (O_902,N_19243,N_16118);
nand UO_903 (O_903,N_19110,N_19347);
or UO_904 (O_904,N_19735,N_15502);
nor UO_905 (O_905,N_17166,N_18554);
and UO_906 (O_906,N_17341,N_16009);
or UO_907 (O_907,N_16842,N_18161);
nor UO_908 (O_908,N_17261,N_16419);
or UO_909 (O_909,N_15699,N_18823);
nand UO_910 (O_910,N_18746,N_17523);
or UO_911 (O_911,N_16749,N_16492);
and UO_912 (O_912,N_19021,N_15782);
and UO_913 (O_913,N_18375,N_16437);
and UO_914 (O_914,N_18163,N_17180);
and UO_915 (O_915,N_15996,N_17974);
nor UO_916 (O_916,N_16630,N_18219);
nand UO_917 (O_917,N_15821,N_16171);
and UO_918 (O_918,N_19999,N_18700);
or UO_919 (O_919,N_19427,N_18877);
and UO_920 (O_920,N_17813,N_16483);
and UO_921 (O_921,N_16968,N_19857);
and UO_922 (O_922,N_16486,N_19082);
nor UO_923 (O_923,N_16867,N_15312);
nor UO_924 (O_924,N_17296,N_19294);
xnor UO_925 (O_925,N_17343,N_17583);
nand UO_926 (O_926,N_16325,N_15471);
and UO_927 (O_927,N_18546,N_19153);
nor UO_928 (O_928,N_15935,N_19295);
nor UO_929 (O_929,N_15667,N_18407);
or UO_930 (O_930,N_19560,N_17394);
nand UO_931 (O_931,N_19487,N_16839);
nor UO_932 (O_932,N_19886,N_18622);
or UO_933 (O_933,N_18171,N_15781);
xnor UO_934 (O_934,N_17276,N_19734);
xor UO_935 (O_935,N_17704,N_19203);
nor UO_936 (O_936,N_19008,N_17911);
xor UO_937 (O_937,N_18933,N_18829);
nand UO_938 (O_938,N_18099,N_19689);
nor UO_939 (O_939,N_15675,N_19499);
and UO_940 (O_940,N_17985,N_16220);
nor UO_941 (O_941,N_19854,N_17951);
or UO_942 (O_942,N_16788,N_19966);
nand UO_943 (O_943,N_16107,N_17515);
and UO_944 (O_944,N_18090,N_19622);
or UO_945 (O_945,N_19927,N_18392);
or UO_946 (O_946,N_16913,N_16707);
nor UO_947 (O_947,N_15888,N_19557);
nor UO_948 (O_948,N_15597,N_18841);
nor UO_949 (O_949,N_15487,N_18029);
or UO_950 (O_950,N_15278,N_15004);
nand UO_951 (O_951,N_15370,N_18118);
or UO_952 (O_952,N_19634,N_16516);
nand UO_953 (O_953,N_19093,N_15382);
nand UO_954 (O_954,N_16207,N_15901);
and UO_955 (O_955,N_17679,N_19400);
nor UO_956 (O_956,N_18932,N_15567);
and UO_957 (O_957,N_16684,N_15664);
nand UO_958 (O_958,N_19781,N_19807);
nor UO_959 (O_959,N_16306,N_15328);
nor UO_960 (O_960,N_18651,N_19620);
and UO_961 (O_961,N_18898,N_18662);
or UO_962 (O_962,N_16470,N_15179);
and UO_963 (O_963,N_18087,N_18914);
or UO_964 (O_964,N_17651,N_19748);
nand UO_965 (O_965,N_17029,N_18916);
and UO_966 (O_966,N_17669,N_18534);
nand UO_967 (O_967,N_15993,N_19453);
and UO_968 (O_968,N_17772,N_16890);
or UO_969 (O_969,N_15799,N_19704);
nor UO_970 (O_970,N_15381,N_18245);
or UO_971 (O_971,N_18760,N_18679);
nor UO_972 (O_972,N_16140,N_18049);
and UO_973 (O_973,N_15515,N_15181);
nand UO_974 (O_974,N_16270,N_17382);
nor UO_975 (O_975,N_16462,N_17603);
or UO_976 (O_976,N_17104,N_18710);
nand UO_977 (O_977,N_18891,N_18655);
and UO_978 (O_978,N_16908,N_17747);
and UO_979 (O_979,N_17853,N_19438);
and UO_980 (O_980,N_17124,N_19592);
nor UO_981 (O_981,N_18741,N_16997);
nand UO_982 (O_982,N_17237,N_19712);
nand UO_983 (O_983,N_17868,N_18752);
nor UO_984 (O_984,N_19747,N_18705);
nand UO_985 (O_985,N_15540,N_17736);
or UO_986 (O_986,N_17976,N_17400);
and UO_987 (O_987,N_16597,N_16482);
nor UO_988 (O_988,N_19456,N_15496);
nand UO_989 (O_989,N_19696,N_17151);
nand UO_990 (O_990,N_16500,N_16530);
nand UO_991 (O_991,N_18789,N_16843);
nand UO_992 (O_992,N_18548,N_16659);
or UO_993 (O_993,N_15807,N_18272);
nand UO_994 (O_994,N_15085,N_16586);
nor UO_995 (O_995,N_18433,N_17365);
or UO_996 (O_996,N_16161,N_17310);
or UO_997 (O_997,N_17462,N_18747);
nand UO_998 (O_998,N_17320,N_17024);
nand UO_999 (O_999,N_19866,N_16395);
or UO_1000 (O_1000,N_17783,N_19351);
or UO_1001 (O_1001,N_15035,N_15334);
or UO_1002 (O_1002,N_16286,N_16897);
nor UO_1003 (O_1003,N_15019,N_18179);
or UO_1004 (O_1004,N_17936,N_17562);
and UO_1005 (O_1005,N_16127,N_18134);
nand UO_1006 (O_1006,N_19918,N_18173);
xnor UO_1007 (O_1007,N_18543,N_15485);
and UO_1008 (O_1008,N_15924,N_19435);
nor UO_1009 (O_1009,N_18055,N_16177);
or UO_1010 (O_1010,N_15178,N_19235);
or UO_1011 (O_1011,N_15611,N_16351);
and UO_1012 (O_1012,N_15869,N_19112);
and UO_1013 (O_1013,N_16554,N_15340);
nand UO_1014 (O_1014,N_17743,N_17552);
nor UO_1015 (O_1015,N_17661,N_16364);
and UO_1016 (O_1016,N_15187,N_18629);
nor UO_1017 (O_1017,N_19387,N_18268);
or UO_1018 (O_1018,N_17801,N_19240);
nor UO_1019 (O_1019,N_16070,N_16004);
xnor UO_1020 (O_1020,N_15751,N_18685);
nand UO_1021 (O_1021,N_18389,N_16821);
or UO_1022 (O_1022,N_18424,N_19606);
or UO_1023 (O_1023,N_15758,N_18347);
and UO_1024 (O_1024,N_15759,N_17908);
or UO_1025 (O_1025,N_17475,N_19850);
nand UO_1026 (O_1026,N_15878,N_15053);
nor UO_1027 (O_1027,N_17918,N_16525);
or UO_1028 (O_1028,N_19253,N_18069);
and UO_1029 (O_1029,N_15787,N_15136);
nand UO_1030 (O_1030,N_17342,N_17687);
nor UO_1031 (O_1031,N_15719,N_19996);
nand UO_1032 (O_1032,N_16903,N_19285);
nand UO_1033 (O_1033,N_18555,N_19457);
nor UO_1034 (O_1034,N_19061,N_19445);
nand UO_1035 (O_1035,N_17537,N_18403);
and UO_1036 (O_1036,N_17277,N_18071);
or UO_1037 (O_1037,N_16589,N_15865);
nor UO_1038 (O_1038,N_15001,N_17323);
nand UO_1039 (O_1039,N_19335,N_17063);
or UO_1040 (O_1040,N_15347,N_16287);
nand UO_1041 (O_1041,N_15594,N_15354);
and UO_1042 (O_1042,N_19216,N_16361);
and UO_1043 (O_1043,N_16357,N_15326);
nor UO_1044 (O_1044,N_19884,N_19998);
or UO_1045 (O_1045,N_16794,N_15665);
nand UO_1046 (O_1046,N_16765,N_16066);
nor UO_1047 (O_1047,N_16295,N_17636);
nor UO_1048 (O_1048,N_15866,N_15871);
and UO_1049 (O_1049,N_19654,N_15126);
nand UO_1050 (O_1050,N_17729,N_19042);
and UO_1051 (O_1051,N_18968,N_16136);
and UO_1052 (O_1052,N_18472,N_18755);
and UO_1053 (O_1053,N_18483,N_18831);
nand UO_1054 (O_1054,N_16454,N_18142);
and UO_1055 (O_1055,N_19057,N_19628);
nor UO_1056 (O_1056,N_15687,N_17120);
nand UO_1057 (O_1057,N_19023,N_16491);
or UO_1058 (O_1058,N_15803,N_16896);
nor UO_1059 (O_1059,N_15656,N_17136);
nand UO_1060 (O_1060,N_18597,N_17929);
nor UO_1061 (O_1061,N_19444,N_15264);
nand UO_1062 (O_1062,N_17535,N_16381);
nand UO_1063 (O_1063,N_17418,N_15818);
nand UO_1064 (O_1064,N_19977,N_18091);
nand UO_1065 (O_1065,N_15544,N_18603);
nand UO_1066 (O_1066,N_19299,N_18127);
and UO_1067 (O_1067,N_18606,N_16995);
nor UO_1068 (O_1068,N_16109,N_16570);
and UO_1069 (O_1069,N_19730,N_15092);
xor UO_1070 (O_1070,N_19277,N_16706);
nor UO_1071 (O_1071,N_18739,N_16758);
nand UO_1072 (O_1072,N_18507,N_15733);
or UO_1073 (O_1073,N_19416,N_16633);
or UO_1074 (O_1074,N_18888,N_18227);
nand UO_1075 (O_1075,N_17865,N_19891);
nor UO_1076 (O_1076,N_17410,N_19300);
nand UO_1077 (O_1077,N_17393,N_15829);
and UO_1078 (O_1078,N_17718,N_19640);
and UO_1079 (O_1079,N_19610,N_15979);
nand UO_1080 (O_1080,N_18167,N_19855);
nand UO_1081 (O_1081,N_16702,N_16355);
nand UO_1082 (O_1082,N_17241,N_17848);
nor UO_1083 (O_1083,N_16225,N_17932);
or UO_1084 (O_1084,N_18225,N_16870);
nor UO_1085 (O_1085,N_17380,N_15532);
nand UO_1086 (O_1086,N_15652,N_18144);
nor UO_1087 (O_1087,N_16432,N_17749);
nor UO_1088 (O_1088,N_19802,N_16598);
or UO_1089 (O_1089,N_15069,N_16810);
and UO_1090 (O_1090,N_16015,N_17501);
and UO_1091 (O_1091,N_16202,N_15500);
nand UO_1092 (O_1092,N_19795,N_17309);
or UO_1093 (O_1093,N_15507,N_15885);
nand UO_1094 (O_1094,N_19586,N_19629);
and UO_1095 (O_1095,N_16143,N_18335);
nand UO_1096 (O_1096,N_19859,N_17152);
or UO_1097 (O_1097,N_18688,N_18153);
nand UO_1098 (O_1098,N_19363,N_16943);
nor UO_1099 (O_1099,N_19354,N_17036);
and UO_1100 (O_1100,N_17949,N_16812);
and UO_1101 (O_1101,N_19609,N_19213);
nand UO_1102 (O_1102,N_16342,N_16919);
nor UO_1103 (O_1103,N_18003,N_17875);
nand UO_1104 (O_1104,N_19089,N_15765);
and UO_1105 (O_1105,N_15831,N_17750);
or UO_1106 (O_1106,N_15243,N_18886);
or UO_1107 (O_1107,N_17790,N_15666);
and UO_1108 (O_1108,N_16889,N_17047);
and UO_1109 (O_1109,N_17307,N_18359);
and UO_1110 (O_1110,N_15365,N_17944);
nor UO_1111 (O_1111,N_16571,N_18609);
nor UO_1112 (O_1112,N_15190,N_17298);
nand UO_1113 (O_1113,N_17362,N_18137);
and UO_1114 (O_1114,N_18265,N_17201);
or UO_1115 (O_1115,N_18601,N_19452);
nand UO_1116 (O_1116,N_19459,N_16768);
and UO_1117 (O_1117,N_16550,N_19682);
nor UO_1118 (O_1118,N_18280,N_18664);
nand UO_1119 (O_1119,N_17516,N_15637);
nor UO_1120 (O_1120,N_16746,N_17297);
or UO_1121 (O_1121,N_19207,N_18666);
nor UO_1122 (O_1122,N_16762,N_16159);
or UO_1123 (O_1123,N_18308,N_17527);
or UO_1124 (O_1124,N_17032,N_19901);
nand UO_1125 (O_1125,N_19292,N_19880);
nor UO_1126 (O_1126,N_18086,N_17517);
or UO_1127 (O_1127,N_18228,N_19278);
and UO_1128 (O_1128,N_16994,N_19264);
nor UO_1129 (O_1129,N_18946,N_19646);
nand UO_1130 (O_1130,N_17485,N_17659);
nand UO_1131 (O_1131,N_19031,N_18957);
nor UO_1132 (O_1132,N_18425,N_16669);
or UO_1133 (O_1133,N_15406,N_16726);
nor UO_1134 (O_1134,N_19926,N_17785);
nor UO_1135 (O_1135,N_19739,N_18937);
or UO_1136 (O_1136,N_15167,N_17928);
and UO_1137 (O_1137,N_15711,N_19959);
and UO_1138 (O_1138,N_16089,N_19162);
nor UO_1139 (O_1139,N_16732,N_18712);
xor UO_1140 (O_1140,N_19352,N_17824);
nor UO_1141 (O_1141,N_19764,N_16663);
or UO_1142 (O_1142,N_17329,N_19114);
or UO_1143 (O_1143,N_15548,N_19987);
and UO_1144 (O_1144,N_19497,N_18439);
and UO_1145 (O_1145,N_17008,N_16792);
nor UO_1146 (O_1146,N_18463,N_16543);
or UO_1147 (O_1147,N_18608,N_19842);
nand UO_1148 (O_1148,N_17345,N_15828);
and UO_1149 (O_1149,N_15976,N_15192);
or UO_1150 (O_1150,N_17995,N_18895);
or UO_1151 (O_1151,N_17645,N_19767);
nor UO_1152 (O_1152,N_15934,N_15320);
or UO_1153 (O_1153,N_18156,N_18100);
and UO_1154 (O_1154,N_16147,N_15221);
or UO_1155 (O_1155,N_18541,N_18148);
and UO_1156 (O_1156,N_19524,N_16343);
or UO_1157 (O_1157,N_17049,N_18751);
and UO_1158 (O_1158,N_17093,N_19003);
nand UO_1159 (O_1159,N_15614,N_17404);
nor UO_1160 (O_1160,N_18868,N_15225);
nor UO_1161 (O_1161,N_19128,N_16251);
nor UO_1162 (O_1162,N_18707,N_18455);
nor UO_1163 (O_1163,N_16620,N_15168);
nand UO_1164 (O_1164,N_17637,N_16963);
nor UO_1165 (O_1165,N_19379,N_19550);
nand UO_1166 (O_1166,N_17140,N_19934);
nor UO_1167 (O_1167,N_15547,N_18820);
and UO_1168 (O_1168,N_17248,N_18814);
or UO_1169 (O_1169,N_19618,N_18848);
or UO_1170 (O_1170,N_17899,N_16453);
nand UO_1171 (O_1171,N_18902,N_17616);
or UO_1172 (O_1172,N_16132,N_19617);
or UO_1173 (O_1173,N_19480,N_17189);
and UO_1174 (O_1174,N_16053,N_18104);
nand UO_1175 (O_1175,N_17518,N_18493);
xor UO_1176 (O_1176,N_16393,N_16459);
and UO_1177 (O_1177,N_15804,N_18802);
or UO_1178 (O_1178,N_15493,N_17971);
nor UO_1179 (O_1179,N_16399,N_15533);
and UO_1180 (O_1180,N_17709,N_15926);
or UO_1181 (O_1181,N_15466,N_15362);
nor UO_1182 (O_1182,N_18152,N_15250);
or UO_1183 (O_1183,N_17578,N_18566);
nand UO_1184 (O_1184,N_18718,N_17889);
nor UO_1185 (O_1185,N_15553,N_15536);
nor UO_1186 (O_1186,N_15315,N_17526);
or UO_1187 (O_1187,N_17053,N_19983);
or UO_1188 (O_1188,N_19613,N_18488);
nand UO_1189 (O_1189,N_15122,N_17211);
nor UO_1190 (O_1190,N_19716,N_18879);
nand UO_1191 (O_1191,N_18525,N_17111);
or UO_1192 (O_1192,N_15601,N_19188);
and UO_1193 (O_1193,N_15020,N_18873);
nand UO_1194 (O_1194,N_18343,N_18015);
nand UO_1195 (O_1195,N_18638,N_15577);
and UO_1196 (O_1196,N_19699,N_19701);
and UO_1197 (O_1197,N_15032,N_15914);
nand UO_1198 (O_1198,N_17947,N_15631);
and UO_1199 (O_1199,N_15651,N_16742);
nor UO_1200 (O_1200,N_16451,N_17294);
and UO_1201 (O_1201,N_17628,N_15574);
or UO_1202 (O_1202,N_19817,N_16535);
nor UO_1203 (O_1203,N_19933,N_16750);
or UO_1204 (O_1204,N_17060,N_18860);
nor UO_1205 (O_1205,N_17869,N_19309);
and UO_1206 (O_1206,N_17451,N_16553);
nor UO_1207 (O_1207,N_18465,N_19227);
nand UO_1208 (O_1208,N_19603,N_19172);
or UO_1209 (O_1209,N_17984,N_18338);
nand UO_1210 (O_1210,N_15210,N_15140);
nor UO_1211 (O_1211,N_16695,N_17857);
and UO_1212 (O_1212,N_18633,N_17398);
and UO_1213 (O_1213,N_17455,N_15180);
or UO_1214 (O_1214,N_17126,N_18082);
or UO_1215 (O_1215,N_18018,N_19798);
or UO_1216 (O_1216,N_17794,N_15839);
or UO_1217 (O_1217,N_17048,N_17256);
nand UO_1218 (O_1218,N_15558,N_15746);
or UO_1219 (O_1219,N_17472,N_15125);
nand UO_1220 (O_1220,N_15542,N_15969);
nor UO_1221 (O_1221,N_15030,N_18300);
nor UO_1222 (O_1222,N_18473,N_17585);
nor UO_1223 (O_1223,N_18661,N_18293);
nor UO_1224 (O_1224,N_15840,N_18189);
nand UO_1225 (O_1225,N_18215,N_19233);
nor UO_1226 (O_1226,N_16776,N_16777);
nor UO_1227 (O_1227,N_17776,N_17348);
nor UO_1228 (O_1228,N_15593,N_15036);
or UO_1229 (O_1229,N_18158,N_16498);
nor UO_1230 (O_1230,N_15668,N_15417);
nand UO_1231 (O_1231,N_18586,N_17009);
nand UO_1232 (O_1232,N_15260,N_15690);
or UO_1233 (O_1233,N_17582,N_19956);
or UO_1234 (O_1234,N_18899,N_15435);
and UO_1235 (O_1235,N_15475,N_17751);
and UO_1236 (O_1236,N_19239,N_17958);
nor UO_1237 (O_1237,N_18620,N_17479);
or UO_1238 (O_1238,N_19761,N_18081);
and UO_1239 (O_1239,N_18596,N_17793);
nor UO_1240 (O_1240,N_16126,N_16204);
nand UO_1241 (O_1241,N_15403,N_17884);
nand UO_1242 (O_1242,N_17808,N_17662);
nor UO_1243 (O_1243,N_16796,N_18107);
nor UO_1244 (O_1244,N_15342,N_16254);
nor UO_1245 (O_1245,N_15771,N_16071);
nand UO_1246 (O_1246,N_15201,N_17305);
nand UO_1247 (O_1247,N_15812,N_17745);
nor UO_1248 (O_1248,N_19198,N_19851);
and UO_1249 (O_1249,N_19976,N_18627);
or UO_1250 (O_1250,N_15576,N_17182);
nor UO_1251 (O_1251,N_15550,N_16942);
nor UO_1252 (O_1252,N_17163,N_18623);
nor UO_1253 (O_1253,N_19493,N_19458);
and UO_1254 (O_1254,N_15663,N_16108);
and UO_1255 (O_1255,N_19836,N_17130);
and UO_1256 (O_1256,N_15259,N_19148);
or UO_1257 (O_1257,N_17235,N_18247);
and UO_1258 (O_1258,N_18164,N_18501);
or UO_1259 (O_1259,N_15464,N_16165);
nor UO_1260 (O_1260,N_18462,N_16809);
nand UO_1261 (O_1261,N_18365,N_17031);
nor UO_1262 (O_1262,N_19096,N_19122);
or UO_1263 (O_1263,N_16430,N_18815);
and UO_1264 (O_1264,N_19450,N_18788);
nand UO_1265 (O_1265,N_15769,N_19259);
nor UO_1266 (O_1266,N_18918,N_16604);
nand UO_1267 (O_1267,N_16264,N_15421);
and UO_1268 (O_1268,N_18218,N_19202);
nand UO_1269 (O_1269,N_17548,N_17888);
nor UO_1270 (O_1270,N_16918,N_15404);
or UO_1271 (O_1271,N_18072,N_19731);
xor UO_1272 (O_1272,N_18617,N_16583);
and UO_1273 (O_1273,N_15641,N_18524);
nand UO_1274 (O_1274,N_15047,N_15065);
nor UO_1275 (O_1275,N_17975,N_15349);
and UO_1276 (O_1276,N_15422,N_19179);
or UO_1277 (O_1277,N_16478,N_15908);
and UO_1278 (O_1278,N_15681,N_19681);
nor UO_1279 (O_1279,N_19304,N_16214);
nand UO_1280 (O_1280,N_19830,N_15149);
nand UO_1281 (O_1281,N_15893,N_17990);
or UO_1282 (O_1282,N_17554,N_17171);
xor UO_1283 (O_1283,N_19718,N_15729);
nor UO_1284 (O_1284,N_18965,N_17283);
and UO_1285 (O_1285,N_16200,N_18625);
nor UO_1286 (O_1286,N_17452,N_17858);
nand UO_1287 (O_1287,N_15023,N_18352);
nand UO_1288 (O_1288,N_17004,N_17232);
nand UO_1289 (O_1289,N_17862,N_16740);
nor UO_1290 (O_1290,N_15915,N_16093);
and UO_1291 (O_1291,N_19793,N_15391);
nand UO_1292 (O_1292,N_18799,N_17581);
nand UO_1293 (O_1293,N_16205,N_17952);
nand UO_1294 (O_1294,N_17020,N_15478);
or UO_1295 (O_1295,N_19580,N_16113);
nor UO_1296 (O_1296,N_16548,N_18386);
nand UO_1297 (O_1297,N_15596,N_17553);
and UO_1298 (O_1298,N_15317,N_17017);
nand UO_1299 (O_1299,N_17575,N_16139);
or UO_1300 (O_1300,N_17245,N_16838);
or UO_1301 (O_1301,N_17977,N_19642);
and UO_1302 (O_1302,N_15977,N_18115);
nand UO_1303 (O_1303,N_16341,N_16804);
nor UO_1304 (O_1304,N_15861,N_15777);
nor UO_1305 (O_1305,N_18469,N_15042);
nor UO_1306 (O_1306,N_15446,N_17569);
and UO_1307 (O_1307,N_16715,N_19468);
nor UO_1308 (O_1308,N_15956,N_17041);
and UO_1309 (O_1309,N_19342,N_15131);
and UO_1310 (O_1310,N_16416,N_16533);
nor UO_1311 (O_1311,N_15115,N_15337);
nor UO_1312 (O_1312,N_19695,N_15623);
nand UO_1313 (O_1313,N_16194,N_17766);
or UO_1314 (O_1314,N_16853,N_16055);
nor UO_1315 (O_1315,N_16210,N_16729);
and UO_1316 (O_1316,N_16310,N_16417);
and UO_1317 (O_1317,N_19013,N_17076);
or UO_1318 (O_1318,N_16090,N_15505);
or UO_1319 (O_1319,N_15872,N_15599);
nand UO_1320 (O_1320,N_15234,N_19319);
or UO_1321 (O_1321,N_18182,N_19388);
nand UO_1322 (O_1322,N_18669,N_16021);
nand UO_1323 (O_1323,N_15449,N_15056);
nand UO_1324 (O_1324,N_17605,N_15902);
and UO_1325 (O_1325,N_16766,N_17396);
nand UO_1326 (O_1326,N_17337,N_15388);
or UO_1327 (O_1327,N_17806,N_17127);
nand UO_1328 (O_1328,N_16130,N_18223);
or UO_1329 (O_1329,N_16269,N_15028);
or UO_1330 (O_1330,N_16213,N_19034);
nor UO_1331 (O_1331,N_15241,N_17058);
and UO_1332 (O_1332,N_17476,N_17778);
and UO_1333 (O_1333,N_18921,N_17689);
and UO_1334 (O_1334,N_17369,N_16925);
and UO_1335 (O_1335,N_15794,N_17121);
or UO_1336 (O_1336,N_15465,N_15329);
and UO_1337 (O_1337,N_17056,N_15458);
nor UO_1338 (O_1338,N_19307,N_18445);
and UO_1339 (O_1339,N_18289,N_15274);
nand UO_1340 (O_1340,N_17100,N_16155);
xnor UO_1341 (O_1341,N_18578,N_16681);
nand UO_1342 (O_1342,N_18522,N_18231);
and UO_1343 (O_1343,N_15240,N_18482);
nand UO_1344 (O_1344,N_16052,N_17374);
nand UO_1345 (O_1345,N_19157,N_15541);
and UO_1346 (O_1346,N_18129,N_18735);
nor UO_1347 (O_1347,N_15918,N_16246);
and UO_1348 (O_1348,N_15106,N_18680);
nand UO_1349 (O_1349,N_15052,N_16039);
or UO_1350 (O_1350,N_15970,N_17966);
or UO_1351 (O_1351,N_19514,N_18404);
or UO_1352 (O_1352,N_19751,N_16534);
nand UO_1353 (O_1353,N_15763,N_16845);
or UO_1354 (O_1354,N_16461,N_15339);
nand UO_1355 (O_1355,N_15238,N_19302);
or UO_1356 (O_1356,N_15359,N_16964);
and UO_1357 (O_1357,N_18384,N_18050);
or UO_1358 (O_1358,N_18942,N_15144);
and UO_1359 (O_1359,N_17595,N_18970);
and UO_1360 (O_1360,N_19978,N_16276);
and UO_1361 (O_1361,N_19230,N_17471);
and UO_1362 (O_1362,N_18269,N_18805);
nand UO_1363 (O_1363,N_17413,N_16048);
nand UO_1364 (O_1364,N_15772,N_18266);
and UO_1365 (O_1365,N_17871,N_15117);
and UO_1366 (O_1366,N_18363,N_15400);
or UO_1367 (O_1367,N_19326,N_19814);
xor UO_1368 (O_1368,N_15696,N_19515);
and UO_1369 (O_1369,N_19693,N_16998);
or UO_1370 (O_1370,N_16373,N_18314);
xor UO_1371 (O_1371,N_18605,N_17293);
and UO_1372 (O_1372,N_15067,N_15798);
and UO_1373 (O_1373,N_17873,N_19001);
and UO_1374 (O_1374,N_18600,N_15110);
and UO_1375 (O_1375,N_16467,N_17807);
nor UO_1376 (O_1376,N_15034,N_19936);
and UO_1377 (O_1377,N_17322,N_15523);
nand UO_1378 (O_1378,N_15529,N_16386);
or UO_1379 (O_1379,N_15022,N_16282);
nor UO_1380 (O_1380,N_19835,N_19052);
nand UO_1381 (O_1381,N_15364,N_16468);
and UO_1382 (O_1382,N_17464,N_18678);
nand UO_1383 (O_1383,N_16678,N_15175);
nand UO_1384 (O_1384,N_16154,N_15205);
or UO_1385 (O_1385,N_19492,N_17615);
and UO_1386 (O_1386,N_19432,N_16875);
and UO_1387 (O_1387,N_17217,N_15224);
nor UO_1388 (O_1388,N_19092,N_18749);
and UO_1389 (O_1389,N_17061,N_19805);
or UO_1390 (O_1390,N_15394,N_15551);
or UO_1391 (O_1391,N_17764,N_19853);
or UO_1392 (O_1392,N_15164,N_19714);
nor UO_1393 (O_1393,N_15737,N_17278);
and UO_1394 (O_1394,N_19281,N_17077);
nand UO_1395 (O_1395,N_19019,N_19017);
nor UO_1396 (O_1396,N_15459,N_15055);
and UO_1397 (O_1397,N_19115,N_16082);
nand UO_1398 (O_1398,N_16346,N_17253);
or UO_1399 (O_1399,N_17459,N_18174);
or UO_1400 (O_1400,N_19931,N_19587);
nor UO_1401 (O_1401,N_15589,N_16387);
nand UO_1402 (O_1402,N_16627,N_17604);
or UO_1403 (O_1403,N_19144,N_19952);
and UO_1404 (O_1404,N_18962,N_15874);
nor UO_1405 (O_1405,N_16584,N_17912);
nor UO_1406 (O_1406,N_16510,N_17156);
xnor UO_1407 (O_1407,N_17499,N_18920);
or UO_1408 (O_1408,N_19986,N_18076);
nand UO_1409 (O_1409,N_17169,N_16131);
nand UO_1410 (O_1410,N_16406,N_16117);
and UO_1411 (O_1411,N_15870,N_16927);
nand UO_1412 (O_1412,N_18239,N_18989);
and UO_1413 (O_1413,N_19257,N_16336);
nor UO_1414 (O_1414,N_16074,N_17469);
or UO_1415 (O_1415,N_19305,N_17668);
or UO_1416 (O_1416,N_19357,N_19984);
or UO_1417 (O_1417,N_18136,N_17505);
nand UO_1418 (O_1418,N_18976,N_18581);
nor UO_1419 (O_1419,N_19339,N_19593);
and UO_1420 (O_1420,N_17588,N_16484);
nand UO_1421 (O_1421,N_17439,N_19337);
nand UO_1422 (O_1422,N_19883,N_18221);
nand UO_1423 (O_1423,N_17761,N_17522);
nor UO_1424 (O_1424,N_17556,N_15527);
and UO_1425 (O_1425,N_18893,N_17707);
nand UO_1426 (O_1426,N_17992,N_16242);
and UO_1427 (O_1427,N_16374,N_15779);
and UO_1428 (O_1428,N_15494,N_18843);
nor UO_1429 (O_1429,N_19821,N_15948);
nand UO_1430 (O_1430,N_15953,N_15830);
nand UO_1431 (O_1431,N_15568,N_16173);
and UO_1432 (O_1432,N_17874,N_16522);
nor UO_1433 (O_1433,N_16289,N_17052);
and UO_1434 (O_1434,N_18301,N_15437);
nor UO_1435 (O_1435,N_17877,N_18060);
nand UO_1436 (O_1436,N_17654,N_15425);
nor UO_1437 (O_1437,N_15635,N_19428);
nand UO_1438 (O_1438,N_15686,N_15565);
nand UO_1439 (O_1439,N_18954,N_15295);
nand UO_1440 (O_1440,N_17597,N_19670);
nand UO_1441 (O_1441,N_18811,N_19811);
or UO_1442 (O_1442,N_16119,N_19590);
or UO_1443 (O_1443,N_18845,N_15764);
or UO_1444 (O_1444,N_18753,N_18966);
and UO_1445 (O_1445,N_16394,N_17706);
nor UO_1446 (O_1446,N_17264,N_17504);
and UO_1447 (O_1447,N_19837,N_19680);
nor UO_1448 (O_1448,N_17630,N_17883);
or UO_1449 (O_1449,N_16380,N_15099);
and UO_1450 (O_1450,N_17770,N_19637);
and UO_1451 (O_1451,N_15265,N_15096);
nand UO_1452 (O_1452,N_15877,N_18772);
or UO_1453 (O_1453,N_19006,N_18504);
nor UO_1454 (O_1454,N_15341,N_15418);
nand UO_1455 (O_1455,N_18444,N_17715);
nand UO_1456 (O_1456,N_15255,N_18778);
and UO_1457 (O_1457,N_15021,N_16549);
nand UO_1458 (O_1458,N_17649,N_19248);
nor UO_1459 (O_1459,N_16905,N_18193);
or UO_1460 (O_1460,N_18821,N_18971);
nand UO_1461 (O_1461,N_17655,N_17635);
nor UO_1462 (O_1462,N_15554,N_19549);
or UO_1463 (O_1463,N_19136,N_16923);
or UO_1464 (O_1464,N_19007,N_15338);
nor UO_1465 (O_1465,N_18177,N_16945);
or UO_1466 (O_1466,N_19265,N_17514);
nor UO_1467 (O_1467,N_16944,N_15420);
nor UO_1468 (O_1468,N_16965,N_17164);
and UO_1469 (O_1469,N_15223,N_16222);
and UO_1470 (O_1470,N_19303,N_15880);
nand UO_1471 (O_1471,N_17863,N_19267);
and UO_1472 (O_1472,N_17885,N_19466);
nor UO_1473 (O_1473,N_18383,N_15972);
nor UO_1474 (O_1474,N_17284,N_16069);
nand UO_1475 (O_1475,N_17238,N_17596);
or UO_1476 (O_1476,N_16218,N_15330);
nor UO_1477 (O_1477,N_19018,N_19963);
nor UO_1478 (O_1478,N_18044,N_16683);
nand UO_1479 (O_1479,N_16886,N_18869);
or UO_1480 (O_1480,N_18242,N_17658);
and UO_1481 (O_1481,N_16224,N_15427);
nand UO_1482 (O_1482,N_19649,N_19974);
and UO_1483 (O_1483,N_17965,N_18533);
and UO_1484 (O_1484,N_18956,N_19502);
nand UO_1485 (O_1485,N_15037,N_19659);
xnor UO_1486 (O_1486,N_17258,N_18306);
nor UO_1487 (O_1487,N_15628,N_15712);
nand UO_1488 (O_1488,N_15632,N_16392);
or UO_1489 (O_1489,N_18532,N_18196);
nor UO_1490 (O_1490,N_17567,N_17409);
and UO_1491 (O_1491,N_16162,N_18448);
and UO_1492 (O_1492,N_16573,N_19574);
or UO_1493 (O_1493,N_17568,N_16323);
nor UO_1494 (O_1494,N_16906,N_17910);
nor UO_1495 (O_1495,N_15378,N_18634);
and UO_1496 (O_1496,N_18593,N_17422);
nand UO_1497 (O_1497,N_15402,N_19941);
nor UO_1498 (O_1498,N_19806,N_16884);
nand UO_1499 (O_1499,N_19827,N_16880);
nor UO_1500 (O_1500,N_16412,N_18194);
nand UO_1501 (O_1501,N_17160,N_16621);
xnor UO_1502 (O_1502,N_16151,N_16092);
nor UO_1503 (O_1503,N_19506,N_19154);
nand UO_1504 (O_1504,N_18973,N_17574);
or UO_1505 (O_1505,N_15564,N_18797);
nand UO_1506 (O_1506,N_16000,N_19993);
nor UO_1507 (O_1507,N_18000,N_15369);
nor UO_1508 (O_1508,N_17760,N_17405);
nand UO_1509 (O_1509,N_15153,N_16996);
nor UO_1510 (O_1510,N_19944,N_16301);
or UO_1511 (O_1511,N_16959,N_18694);
nand UO_1512 (O_1512,N_19085,N_16280);
or UO_1513 (O_1513,N_16524,N_17458);
nor UO_1514 (O_1514,N_18983,N_16786);
nor UO_1515 (O_1515,N_16518,N_19055);
and UO_1516 (O_1516,N_16559,N_15800);
and UO_1517 (O_1517,N_16594,N_15582);
and UO_1518 (O_1518,N_15396,N_16101);
nand UO_1519 (O_1519,N_16731,N_19209);
and UO_1520 (O_1520,N_19350,N_19050);
and UO_1521 (O_1521,N_19375,N_15524);
nand UO_1522 (O_1522,N_15966,N_17318);
nor UO_1523 (O_1523,N_15017,N_17159);
nand UO_1524 (O_1524,N_16654,N_18094);
or UO_1525 (O_1525,N_16235,N_16384);
nand UO_1526 (O_1526,N_16741,N_15482);
and UO_1527 (O_1527,N_19036,N_19033);
or UO_1528 (O_1528,N_17520,N_15923);
or UO_1529 (O_1529,N_17252,N_16541);
xor UO_1530 (O_1530,N_19980,N_15098);
nand UO_1531 (O_1531,N_17672,N_17601);
nor UO_1532 (O_1532,N_18053,N_16456);
and UO_1533 (O_1533,N_17260,N_19694);
nand UO_1534 (O_1534,N_17904,N_17403);
nand UO_1535 (O_1535,N_17378,N_17094);
nor UO_1536 (O_1536,N_15024,N_19176);
nor UO_1537 (O_1537,N_18865,N_19916);
nor UO_1538 (O_1538,N_18692,N_19728);
nand UO_1539 (O_1539,N_16186,N_15046);
nand UO_1540 (O_1540,N_19511,N_16582);
or UO_1541 (O_1541,N_15756,N_16309);
or UO_1542 (O_1542,N_17387,N_17473);
and UO_1543 (O_1543,N_16211,N_16376);
and UO_1544 (O_1544,N_16427,N_19234);
or UO_1545 (O_1545,N_16871,N_18124);
nand UO_1546 (O_1546,N_17681,N_18332);
and UO_1547 (O_1547,N_15677,N_17510);
nand UO_1548 (O_1548,N_16248,N_15986);
nand UO_1549 (O_1549,N_19686,N_18474);
nor UO_1550 (O_1550,N_19180,N_15363);
nor UO_1551 (O_1551,N_16885,N_16986);
and UO_1552 (O_1552,N_15429,N_17849);
or UO_1553 (O_1553,N_16791,N_17695);
nor UO_1554 (O_1554,N_15743,N_15073);
nand UO_1555 (O_1555,N_16574,N_16956);
or UO_1556 (O_1556,N_15213,N_17489);
nand UO_1557 (O_1557,N_17295,N_16557);
and UO_1558 (O_1558,N_15033,N_16196);
nand UO_1559 (O_1559,N_16993,N_17900);
and UO_1560 (O_1560,N_18197,N_19273);
nand UO_1561 (O_1561,N_16215,N_15890);
nand UO_1562 (O_1562,N_19559,N_17370);
or UO_1563 (O_1563,N_16552,N_18614);
or UO_1564 (O_1564,N_16183,N_16299);
nor UO_1565 (O_1565,N_16146,N_16603);
or UO_1566 (O_1566,N_19488,N_18520);
nand UO_1567 (O_1567,N_19992,N_16312);
or UO_1568 (O_1568,N_15268,N_19776);
nor UO_1569 (O_1569,N_18663,N_15331);
nand UO_1570 (O_1570,N_16527,N_19069);
and UO_1571 (O_1571,N_16674,N_15660);
nor UO_1572 (O_1572,N_16064,N_15911);
nor UO_1573 (O_1573,N_19910,N_18299);
nor UO_1574 (O_1574,N_16724,N_16929);
nor UO_1575 (O_1575,N_18571,N_15889);
nor UO_1576 (O_1576,N_19733,N_17856);
or UO_1577 (O_1577,N_19707,N_15913);
nor UO_1578 (O_1578,N_17754,N_18723);
and UO_1579 (O_1579,N_16977,N_17566);
nand UO_1580 (O_1580,N_17540,N_15026);
and UO_1581 (O_1581,N_15910,N_16626);
and UO_1582 (O_1582,N_16805,N_17602);
or UO_1583 (O_1583,N_18508,N_17924);
nand UO_1584 (O_1584,N_19469,N_16024);
and UO_1585 (O_1585,N_16840,N_19876);
or UO_1586 (O_1586,N_15410,N_19463);
nor UO_1587 (O_1587,N_19226,N_16909);
or UO_1588 (O_1588,N_18125,N_18250);
nand UO_1589 (O_1589,N_18995,N_16096);
nor UO_1590 (O_1590,N_19846,N_17685);
or UO_1591 (O_1591,N_19073,N_19938);
nor UO_1592 (O_1592,N_17266,N_18088);
and UO_1593 (O_1593,N_16232,N_15375);
and UO_1594 (O_1594,N_16699,N_19569);
or UO_1595 (O_1595,N_19205,N_15191);
nor UO_1596 (O_1596,N_15616,N_18297);
and UO_1597 (O_1597,N_16848,N_19482);
and UO_1598 (O_1598,N_16098,N_16972);
nand UO_1599 (O_1599,N_15495,N_19530);
nand UO_1600 (O_1600,N_16600,N_16580);
or UO_1601 (O_1601,N_15102,N_16016);
or UO_1602 (O_1602,N_18259,N_19742);
nor UO_1603 (O_1603,N_16874,N_18599);
and UO_1604 (O_1604,N_18744,N_15038);
nand UO_1605 (O_1605,N_18803,N_15522);
nor UO_1606 (O_1606,N_17739,N_18102);
nor UO_1607 (O_1607,N_17920,N_15521);
nand UO_1608 (O_1608,N_18979,N_19652);
nand UO_1609 (O_1609,N_19032,N_16850);
nor UO_1610 (O_1610,N_17274,N_15868);
and UO_1611 (O_1611,N_18476,N_16471);
and UO_1612 (O_1612,N_17638,N_18572);
or UO_1613 (O_1613,N_16703,N_16673);
nor UO_1614 (O_1614,N_15061,N_16901);
and UO_1615 (O_1615,N_15610,N_15058);
nand UO_1616 (O_1616,N_16297,N_16951);
or UO_1617 (O_1617,N_18830,N_19000);
and UO_1618 (O_1618,N_16575,N_18786);
nor UO_1619 (O_1619,N_19595,N_15372);
nand UO_1620 (O_1620,N_19380,N_19717);
nor UO_1621 (O_1621,N_17146,N_19369);
or UO_1622 (O_1622,N_17700,N_17740);
nor UO_1623 (O_1623,N_19283,N_15196);
or UO_1624 (O_1624,N_19950,N_18585);
or UO_1625 (O_1625,N_16926,N_19636);
nand UO_1626 (O_1626,N_15287,N_18388);
nand UO_1627 (O_1627,N_18461,N_16976);
nand UO_1628 (O_1628,N_18491,N_15797);
and UO_1629 (O_1629,N_15760,N_15704);
nand UO_1630 (O_1630,N_18836,N_18883);
nand UO_1631 (O_1631,N_17705,N_18263);
or UO_1632 (O_1632,N_17200,N_18952);
or UO_1633 (O_1633,N_19507,N_19575);
and UO_1634 (O_1634,N_16797,N_17986);
and UO_1635 (O_1635,N_15762,N_16037);
nor UO_1636 (O_1636,N_19223,N_16060);
nor UO_1637 (O_1637,N_18331,N_16832);
or UO_1638 (O_1638,N_16370,N_16738);
and UO_1639 (O_1639,N_15343,N_16708);
nand UO_1640 (O_1640,N_16935,N_18034);
nor UO_1641 (O_1641,N_16233,N_17960);
or UO_1642 (O_1642,N_17919,N_18116);
nand UO_1643 (O_1643,N_16737,N_15790);
nand UO_1644 (O_1644,N_19002,N_18234);
or UO_1645 (O_1645,N_16523,N_16861);
and UO_1646 (O_1646,N_15896,N_18905);
nor UO_1647 (O_1647,N_19994,N_19471);
or UO_1648 (O_1648,N_16652,N_18341);
nand UO_1649 (O_1649,N_18939,N_17969);
nand UO_1650 (O_1650,N_15509,N_19120);
nor UO_1651 (O_1651,N_16531,N_17401);
and UO_1652 (O_1652,N_19698,N_17226);
nor UO_1653 (O_1653,N_16138,N_17981);
nand UO_1654 (O_1654,N_18748,N_19672);
or UO_1655 (O_1655,N_16110,N_15188);
nor UO_1656 (O_1656,N_19913,N_15415);
or UO_1657 (O_1657,N_19687,N_15963);
or UO_1658 (O_1658,N_17112,N_19130);
and UO_1659 (O_1659,N_18892,N_17617);
or UO_1660 (O_1660,N_16253,N_19788);
or UO_1661 (O_1661,N_19373,N_16073);
nor UO_1662 (O_1662,N_18442,N_15634);
nand UO_1663 (O_1663,N_15189,N_16609);
nor UO_1664 (O_1664,N_19804,N_18320);
and UO_1665 (O_1665,N_17881,N_18992);
nand UO_1666 (O_1666,N_16595,N_18675);
nor UO_1667 (O_1667,N_15503,N_18372);
or UO_1668 (O_1668,N_15256,N_15226);
nor UO_1669 (O_1669,N_15583,N_17727);
nand UO_1670 (O_1670,N_19323,N_19105);
nand UO_1671 (O_1671,N_17765,N_15477);
nand UO_1672 (O_1672,N_19895,N_19673);
or UO_1673 (O_1673,N_18909,N_18485);
nand UO_1674 (O_1674,N_17627,N_15846);
nand UO_1675 (O_1675,N_19650,N_19812);
nor UO_1676 (O_1676,N_19774,N_18758);
and UO_1677 (O_1677,N_17701,N_15141);
and UO_1678 (O_1678,N_16029,N_17332);
and UO_1679 (O_1679,N_17408,N_16413);
nand UO_1680 (O_1680,N_18668,N_19856);
nand UO_1681 (O_1681,N_19979,N_19909);
or UO_1682 (O_1682,N_15944,N_17373);
nor UO_1683 (O_1683,N_17496,N_19782);
nor UO_1684 (O_1684,N_16189,N_15481);
and UO_1685 (O_1685,N_16513,N_18951);
and UO_1686 (O_1686,N_18521,N_16104);
nand UO_1687 (O_1687,N_18850,N_19173);
or UO_1688 (O_1688,N_19430,N_16369);
nand UO_1689 (O_1689,N_16191,N_19164);
nor UO_1690 (O_1690,N_16238,N_16145);
nand UO_1691 (O_1691,N_17346,N_18834);
or UO_1692 (O_1692,N_17509,N_16292);
nor UO_1693 (O_1693,N_17349,N_17288);
and UO_1694 (O_1694,N_18423,N_18409);
and UO_1695 (O_1695,N_17114,N_19293);
nand UO_1696 (O_1696,N_19344,N_19410);
and UO_1697 (O_1697,N_17218,N_15921);
nand UO_1698 (O_1698,N_16957,N_15673);
and UO_1699 (O_1699,N_18535,N_19244);
nand UO_1700 (O_1700,N_19539,N_19237);
or UO_1701 (O_1701,N_19022,N_16710);
nor UO_1702 (O_1702,N_19318,N_15104);
nor UO_1703 (O_1703,N_15514,N_18206);
and UO_1704 (O_1704,N_18896,N_18369);
nand UO_1705 (O_1705,N_16172,N_15207);
and UO_1706 (O_1706,N_19024,N_16239);
or UO_1707 (O_1707,N_19189,N_17787);
or UO_1708 (O_1708,N_18589,N_15640);
nand UO_1709 (O_1709,N_15159,N_17592);
nor UO_1710 (O_1710,N_18985,N_18133);
and UO_1711 (O_1711,N_16318,N_19868);
nand UO_1712 (O_1712,N_17168,N_18490);
nor UO_1713 (O_1713,N_18880,N_15316);
nand UO_1714 (O_1714,N_17478,N_15895);
and UO_1715 (O_1715,N_15081,N_17018);
nand UO_1716 (O_1716,N_19789,N_19087);
xor UO_1717 (O_1717,N_16267,N_16940);
nor UO_1718 (O_1718,N_17150,N_19422);
or UO_1719 (O_1719,N_19113,N_16688);
and UO_1720 (O_1720,N_15276,N_16003);
or UO_1721 (O_1721,N_19765,N_19601);
or UO_1722 (O_1722,N_17068,N_17470);
and UO_1723 (O_1723,N_17821,N_15955);
nor UO_1724 (O_1724,N_17275,N_19183);
or UO_1725 (O_1725,N_19399,N_15506);
nand UO_1726 (O_1726,N_16685,N_17392);
and UO_1727 (O_1727,N_18854,N_17531);
and UO_1728 (O_1728,N_19368,N_19786);
or UO_1729 (O_1729,N_17831,N_15119);
nand UO_1730 (O_1730,N_19780,N_18237);
xor UO_1731 (O_1731,N_15121,N_19771);
nor UO_1732 (O_1732,N_17474,N_17864);
nand UO_1733 (O_1733,N_16693,N_18591);
nor UO_1734 (O_1734,N_19740,N_16313);
and UO_1735 (O_1735,N_16335,N_17728);
or UO_1736 (O_1736,N_18216,N_17840);
nand UO_1737 (O_1737,N_17368,N_18693);
nand UO_1738 (O_1738,N_17843,N_18001);
or UO_1739 (O_1739,N_19152,N_17269);
nor UO_1740 (O_1740,N_15247,N_16902);
or UO_1741 (O_1741,N_15605,N_16560);
and UO_1742 (O_1742,N_16950,N_18517);
or UO_1743 (O_1743,N_18220,N_19702);
and UO_1744 (O_1744,N_15741,N_18101);
and UO_1745 (O_1745,N_15808,N_18974);
and UO_1746 (O_1746,N_17330,N_17767);
nand UO_1747 (O_1747,N_17733,N_17805);
nor UO_1748 (O_1748,N_15630,N_19079);
and UO_1749 (O_1749,N_17762,N_19266);
nand UO_1750 (O_1750,N_17988,N_15819);
nand UO_1751 (O_1751,N_19051,N_19306);
or UO_1752 (O_1752,N_15886,N_16007);
nand UO_1753 (O_1753,N_17154,N_17084);
or UO_1754 (O_1754,N_16888,N_18108);
nand UO_1755 (O_1755,N_16754,N_15517);
or UO_1756 (O_1756,N_19921,N_16816);
or UO_1757 (O_1757,N_19861,N_15368);
and UO_1758 (O_1758,N_15919,N_18408);
xor UO_1759 (O_1759,N_15526,N_16271);
and UO_1760 (O_1760,N_16982,N_18304);
nor UO_1761 (O_1761,N_19270,N_18557);
nand UO_1762 (O_1762,N_19261,N_18198);
nor UO_1763 (O_1763,N_16479,N_19989);
nand UO_1764 (O_1764,N_17571,N_16390);
and UO_1765 (O_1765,N_17312,N_18106);
nor UO_1766 (O_1766,N_19250,N_16612);
nand UO_1767 (O_1767,N_15971,N_15570);
nand UO_1768 (O_1768,N_16465,N_17610);
xnor UO_1769 (O_1769,N_15407,N_18047);
nor UO_1770 (O_1770,N_16969,N_19406);
nand UO_1771 (O_1771,N_19392,N_18342);
or UO_1772 (O_1772,N_15766,N_19065);
or UO_1773 (O_1773,N_15964,N_17677);
and UO_1774 (O_1774,N_18915,N_17525);
nand UO_1775 (O_1775,N_18498,N_16008);
and UO_1776 (O_1776,N_19867,N_17139);
nand UO_1777 (O_1777,N_15604,N_17096);
or UO_1778 (O_1778,N_15332,N_15409);
and UO_1779 (O_1779,N_19316,N_15242);
and UO_1780 (O_1780,N_16917,N_17014);
and UO_1781 (O_1781,N_16611,N_17468);
nor UO_1782 (O_1782,N_19374,N_19004);
nand UO_1783 (O_1783,N_18907,N_16244);
and UO_1784 (O_1784,N_17648,N_19491);
nor UO_1785 (O_1785,N_17081,N_15076);
nor UO_1786 (O_1786,N_18396,N_15499);
or UO_1787 (O_1787,N_17162,N_17287);
and UO_1788 (O_1788,N_19877,N_15617);
nor UO_1789 (O_1789,N_19078,N_19169);
and UO_1790 (O_1790,N_18417,N_19677);
nor UO_1791 (O_1791,N_17935,N_17678);
nor UO_1792 (O_1792,N_19156,N_15313);
nor UO_1793 (O_1793,N_17490,N_16322);
or UO_1794 (O_1794,N_15927,N_19362);
nor UO_1795 (O_1795,N_15817,N_15834);
nand UO_1796 (O_1796,N_18135,N_19370);
or UO_1797 (O_1797,N_18866,N_17498);
or UO_1798 (O_1798,N_18180,N_18945);
or UO_1799 (O_1799,N_18590,N_15715);
or UO_1800 (O_1800,N_16720,N_15981);
and UO_1801 (O_1801,N_15648,N_17313);
nand UO_1802 (O_1802,N_16148,N_17074);
and UO_1803 (O_1803,N_17331,N_18837);
nand UO_1804 (O_1804,N_16916,N_18275);
nand UO_1805 (O_1805,N_16167,N_18458);
nand UO_1806 (O_1806,N_19465,N_17454);
nor UO_1807 (O_1807,N_16606,N_15920);
or UO_1808 (O_1808,N_17402,N_15832);
nor UO_1809 (O_1809,N_15706,N_18402);
nor UO_1810 (O_1810,N_15773,N_16072);
and UO_1811 (O_1811,N_17328,N_19540);
nor UO_1812 (O_1812,N_18006,N_18870);
and UO_1813 (O_1813,N_17815,N_19571);
xor UO_1814 (O_1814,N_18619,N_16175);
nand UO_1815 (O_1815,N_15080,N_16308);
nand UO_1816 (O_1816,N_18998,N_17158);
or UO_1817 (O_1817,N_15324,N_15622);
and UO_1818 (O_1818,N_17830,N_19955);
nand UO_1819 (O_1819,N_19124,N_18856);
or UO_1820 (O_1820,N_18737,N_19770);
and UO_1821 (O_1821,N_16932,N_15206);
and UO_1822 (O_1822,N_15113,N_19217);
nand UO_1823 (O_1823,N_19327,N_15371);
nor UO_1824 (O_1824,N_15887,N_17613);
nor UO_1825 (O_1825,N_15946,N_15767);
or UO_1826 (O_1826,N_17870,N_15293);
or UO_1827 (O_1827,N_19137,N_19809);
or UO_1828 (O_1828,N_17925,N_17898);
nand UO_1829 (O_1829,N_19210,N_18172);
nand UO_1830 (O_1830,N_16231,N_19985);
or UO_1831 (O_1831,N_18849,N_19353);
or UO_1832 (O_1832,N_18919,N_15012);
nor UO_1833 (O_1833,N_15984,N_17119);
nand UO_1834 (O_1834,N_19563,N_16504);
nor UO_1835 (O_1835,N_16400,N_18640);
nor UO_1836 (O_1836,N_18416,N_16640);
nand UO_1837 (O_1837,N_15314,N_19818);
and UO_1838 (O_1838,N_17259,N_19418);
and UO_1839 (O_1839,N_15438,N_19389);
nor UO_1840 (O_1840,N_16442,N_16747);
or UO_1841 (O_1841,N_16423,N_18376);
nand UO_1842 (O_1842,N_17367,N_19849);
nor UO_1843 (O_1843,N_17945,N_15111);
and UO_1844 (O_1844,N_15016,N_18757);
or UO_1845 (O_1845,N_18254,N_19290);
or UO_1846 (O_1846,N_15689,N_15658);
or UO_1847 (O_1847,N_19865,N_18711);
nor UO_1848 (O_1848,N_17584,N_19887);
nand UO_1849 (O_1849,N_16262,N_19358);
and UO_1850 (O_1850,N_16680,N_16449);
or UO_1851 (O_1851,N_16315,N_18835);
or UO_1852 (O_1852,N_16043,N_18563);
nand UO_1853 (O_1853,N_17210,N_15802);
nor UO_1854 (O_1854,N_19588,N_16229);
and UO_1855 (O_1855,N_15796,N_15209);
and UO_1856 (O_1856,N_18871,N_15841);
nor UO_1857 (O_1857,N_16431,N_19246);
nand UO_1858 (O_1858,N_18256,N_18703);
and UO_1859 (O_1859,N_17415,N_16035);
nor UO_1860 (O_1860,N_15473,N_16135);
and UO_1861 (O_1861,N_15588,N_17752);
nand UO_1862 (O_1862,N_17057,N_15740);
nand UO_1863 (O_1863,N_19898,N_17022);
nor UO_1864 (O_1864,N_16664,N_17660);
xnor UO_1865 (O_1865,N_19542,N_19951);
and UO_1866 (O_1866,N_18213,N_18545);
or UO_1867 (O_1867,N_15900,N_18547);
or UO_1868 (O_1868,N_18670,N_17846);
or UO_1869 (O_1869,N_18315,N_18901);
or UO_1870 (O_1870,N_17624,N_19508);
nand UO_1871 (O_1871,N_16551,N_15227);
nand UO_1872 (O_1872,N_18276,N_19583);
nor UO_1873 (O_1873,N_15303,N_19178);
or UO_1874 (O_1874,N_15273,N_16613);
and UO_1875 (O_1875,N_16820,N_19419);
or UO_1876 (O_1876,N_18513,N_17570);
nor UO_1877 (O_1877,N_15361,N_15518);
nor UO_1878 (O_1878,N_17594,N_16266);
or UO_1879 (O_1879,N_15142,N_18986);
or UO_1880 (O_1880,N_15783,N_19763);
nor UO_1881 (O_1881,N_15776,N_15006);
nor UO_1882 (O_1882,N_16983,N_16772);
nand UO_1883 (O_1883,N_15333,N_17955);
or UO_1884 (O_1884,N_17650,N_17391);
nor UO_1885 (O_1885,N_16170,N_15300);
or UO_1886 (O_1886,N_15552,N_19046);
nand UO_1887 (O_1887,N_17227,N_18447);
and UO_1888 (O_1888,N_16526,N_16034);
or UO_1889 (O_1889,N_15615,N_19753);
or UO_1890 (O_1890,N_15090,N_19675);
nor UO_1891 (O_1891,N_15991,N_18641);
and UO_1892 (O_1892,N_18908,N_16798);
nand UO_1893 (O_1893,N_18560,N_16156);
or UO_1894 (O_1894,N_19067,N_15994);
and UO_1895 (O_1895,N_15305,N_16488);
or UO_1896 (O_1896,N_19409,N_16084);
nor UO_1897 (O_1897,N_18765,N_18903);
nand UO_1898 (O_1898,N_19873,N_16641);
nor UO_1899 (O_1899,N_15279,N_19275);
and UO_1900 (O_1900,N_17011,N_19355);
nor UO_1901 (O_1901,N_16354,N_19483);
or UO_1902 (O_1902,N_17742,N_17586);
nand UO_1903 (O_1903,N_18687,N_17062);
and UO_1904 (O_1904,N_18847,N_19084);
and UO_1905 (O_1905,N_18011,N_18796);
or UO_1906 (O_1906,N_16978,N_19063);
and UO_1907 (O_1907,N_17697,N_16166);
or UO_1908 (O_1908,N_18083,N_17860);
nand UO_1909 (O_1909,N_15134,N_15277);
or UO_1910 (O_1910,N_16990,N_17086);
nand UO_1911 (O_1911,N_15084,N_16898);
and UO_1912 (O_1912,N_15261,N_17321);
or UO_1913 (O_1913,N_18929,N_18894);
nand UO_1914 (O_1914,N_19242,N_19589);
nand UO_1915 (O_1915,N_19407,N_15929);
nand UO_1916 (O_1916,N_15501,N_17796);
xnor UO_1917 (O_1917,N_18291,N_19075);
and UO_1918 (O_1918,N_15752,N_15644);
and UO_1919 (O_1919,N_16734,N_18624);
and UO_1920 (O_1920,N_17109,N_18411);
nor UO_1921 (O_1921,N_18510,N_18652);
or UO_1922 (O_1922,N_17447,N_17632);
xor UO_1923 (O_1923,N_18791,N_18981);
and UO_1924 (O_1924,N_15539,N_18940);
xor UO_1925 (O_1925,N_16041,N_18842);
nand UO_1926 (O_1926,N_16223,N_18391);
nand UO_1927 (O_1927,N_15945,N_17185);
nand UO_1928 (O_1928,N_19426,N_15450);
or UO_1929 (O_1929,N_15826,N_19411);
nor UO_1930 (O_1930,N_19076,N_19962);
nor UO_1931 (O_1931,N_19211,N_17098);
or UO_1932 (O_1932,N_18089,N_18516);
nor UO_1933 (O_1933,N_18819,N_15691);
nand UO_1934 (O_1934,N_17539,N_15625);
nand UO_1935 (O_1935,N_19117,N_17735);
or UO_1936 (O_1936,N_18230,N_16241);
nand UO_1937 (O_1937,N_18579,N_19597);
xnor UO_1938 (O_1938,N_17623,N_19611);
and UO_1939 (O_1939,N_18039,N_18551);
nor UO_1940 (O_1940,N_18397,N_15245);
nor UO_1941 (O_1941,N_16824,N_16876);
nand UO_1942 (O_1942,N_18217,N_18294);
and UO_1943 (O_1943,N_17657,N_18176);
nand UO_1944 (O_1944,N_16671,N_17933);
or UO_1945 (O_1945,N_19252,N_17149);
or UO_1946 (O_1946,N_15002,N_15718);
or UO_1947 (O_1947,N_19341,N_18681);
or UO_1948 (O_1948,N_18186,N_17223);
or UO_1949 (O_1949,N_15863,N_17948);
nor UO_1950 (O_1950,N_18713,N_15335);
or UO_1951 (O_1951,N_16319,N_19361);
or UO_1952 (O_1952,N_16780,N_16836);
nor UO_1953 (O_1953,N_19554,N_15619);
nor UO_1954 (O_1954,N_17176,N_16825);
and UO_1955 (O_1955,N_17092,N_18393);
or UO_1956 (O_1956,N_18732,N_19332);
and UO_1957 (O_1957,N_19058,N_19068);
nor UO_1958 (O_1958,N_18175,N_18452);
nor UO_1959 (O_1959,N_16099,N_15319);
or UO_1960 (O_1960,N_17882,N_15789);
nand UO_1961 (O_1961,N_17894,N_18781);
or UO_1962 (O_1962,N_15785,N_15298);
nand UO_1963 (O_1963,N_16495,N_19479);
nand UO_1964 (O_1964,N_18642,N_15158);
or UO_1965 (O_1965,N_16291,N_15683);
and UO_1966 (O_1966,N_17832,N_17543);
or UO_1967 (O_1967,N_16063,N_18395);
or UO_1968 (O_1968,N_16962,N_15726);
or UO_1969 (O_1969,N_17173,N_19190);
or UO_1970 (O_1970,N_18671,N_18676);
nor UO_1971 (O_1971,N_18394,N_16615);
or UO_1972 (O_1972,N_16646,N_18701);
or UO_1973 (O_1973,N_19037,N_16019);
or UO_1974 (O_1974,N_15454,N_18401);
or UO_1975 (O_1975,N_19356,N_17500);
nand UO_1976 (O_1976,N_18724,N_16866);
nor UO_1977 (O_1977,N_19221,N_15903);
nor UO_1978 (O_1978,N_15916,N_18353);
or UO_1979 (O_1979,N_15419,N_15172);
nor UO_1980 (O_1980,N_19915,N_15949);
nand UO_1981 (O_1981,N_19282,N_18698);
nand UO_1982 (O_1982,N_17087,N_17994);
nand UO_1983 (O_1983,N_19044,N_17631);
nor UO_1984 (O_1984,N_15480,N_15103);
and UO_1985 (O_1985,N_16711,N_18832);
nor UO_1986 (O_1986,N_18659,N_18456);
nor UO_1987 (O_1987,N_17915,N_19929);
and UO_1988 (O_1988,N_19888,N_18066);
or UO_1989 (O_1989,N_17675,N_16784);
or UO_1990 (O_1990,N_19801,N_16061);
and UO_1991 (O_1991,N_18540,N_18159);
and UO_1992 (O_1992,N_18653,N_16348);
and UO_1993 (O_1993,N_17075,N_15385);
or UO_1994 (O_1994,N_17265,N_15925);
and UO_1995 (O_1995,N_18333,N_16272);
nand UO_1996 (O_1996,N_18770,N_15244);
or UO_1997 (O_1997,N_18208,N_19241);
or UO_1998 (O_1998,N_15412,N_15289);
and UO_1999 (O_1999,N_19538,N_19543);
nor UO_2000 (O_2000,N_19402,N_18436);
or UO_2001 (O_2001,N_18598,N_16087);
and UO_2002 (O_2002,N_15836,N_18635);
nand UO_2003 (O_2003,N_16022,N_19957);
nor UO_2004 (O_2004,N_16443,N_18080);
or UO_2005 (O_2005,N_15672,N_19894);
nand UO_2006 (O_2006,N_19724,N_19421);
nand UO_2007 (O_2007,N_19820,N_19472);
or UO_2008 (O_2008,N_17876,N_18328);
nor UO_2009 (O_2009,N_16102,N_15197);
nand UO_2010 (O_2010,N_17153,N_17105);
nor UO_2011 (O_2011,N_18809,N_17886);
or UO_2012 (O_2012,N_16651,N_15302);
or UO_2013 (O_2013,N_16141,N_19596);
nand UO_2014 (O_2014,N_16857,N_16056);
nor UO_2015 (O_2015,N_19098,N_19485);
xnor UO_2016 (O_2016,N_19641,N_18910);
nor UO_2017 (O_2017,N_19544,N_18934);
nor UO_2018 (O_2018,N_17722,N_15000);
nand UO_2019 (O_2019,N_15608,N_17714);
and UO_2020 (O_2020,N_17497,N_16446);
or UO_2021 (O_2021,N_18385,N_19397);
nor UO_2022 (O_2022,N_17267,N_18645);
nor UO_2023 (O_2023,N_16757,N_16739);
nor UO_2024 (O_2024,N_18330,N_17892);
or UO_2025 (O_2025,N_15129,N_17626);
or UO_2026 (O_2026,N_16424,N_15235);
xnor UO_2027 (O_2027,N_15254,N_19762);
nand UO_2028 (O_2028,N_18691,N_15239);
nor UO_2029 (O_2029,N_19982,N_18738);
and UO_2030 (O_2030,N_17434,N_15441);
or UO_2031 (O_2031,N_15609,N_15249);
xor UO_2032 (O_2032,N_17115,N_17907);
or UO_2033 (O_2033,N_18309,N_18063);
or UO_2034 (O_2034,N_18255,N_19247);
nand UO_2035 (O_2035,N_19149,N_17530);
or UO_2036 (O_2036,N_19490,N_19661);
or UO_2037 (O_2037,N_18702,N_17456);
nand UO_2038 (O_2038,N_15961,N_18002);
or UO_2039 (O_2039,N_19970,N_17939);
and UO_2040 (O_2040,N_16799,N_16502);
nor UO_2041 (O_2041,N_18209,N_19185);
nor UO_2042 (O_2042,N_15750,N_19750);
and UO_2043 (O_2043,N_16439,N_19521);
xnor UO_2044 (O_2044,N_16198,N_15005);
or UO_2045 (O_2045,N_17890,N_16834);
or UO_2046 (O_2046,N_15639,N_19991);
and UO_2047 (O_2047,N_16179,N_19632);
nor UO_2048 (O_2048,N_19527,N_16662);
and UO_2049 (O_2049,N_15563,N_19943);
nand UO_2050 (O_2050,N_15723,N_18674);
nand UO_2051 (O_2051,N_17703,N_17495);
and UO_2052 (O_2052,N_16566,N_15906);
and UO_2053 (O_2053,N_17078,N_16713);
nor UO_2054 (O_2054,N_16206,N_16404);
or UO_2055 (O_2055,N_18109,N_18912);
and UO_2056 (O_2056,N_16546,N_19501);
and UO_2057 (O_2057,N_19900,N_15626);
nor UO_2058 (O_2058,N_19639,N_16274);
or UO_2059 (O_2059,N_17852,N_18058);
nor UO_2060 (O_2060,N_16105,N_18400);
nand UO_2061 (O_2061,N_17445,N_15307);
nor UO_2062 (O_2062,N_15107,N_19097);
and UO_2063 (O_2063,N_18518,N_16388);
or UO_2064 (O_2064,N_16033,N_15561);
nor UO_2065 (O_2065,N_16628,N_17214);
and UO_2066 (O_2066,N_15405,N_15936);
nor UO_2067 (O_2067,N_19667,N_17692);
nor UO_2068 (O_2068,N_15114,N_18311);
nor UO_2069 (O_2069,N_15806,N_17250);
and UO_2070 (O_2070,N_19333,N_15643);
and UO_2071 (O_2071,N_19669,N_18367);
and UO_2072 (O_2072,N_18725,N_17213);
and UO_2073 (O_2073,N_15075,N_15200);
nor UO_2074 (O_2074,N_18878,N_18682);
or UO_2075 (O_2075,N_17132,N_18611);
nor UO_2076 (O_2076,N_17532,N_17961);
nand UO_2077 (O_2077,N_18278,N_16474);
and UO_2078 (O_2078,N_17850,N_18780);
or UO_2079 (O_2079,N_18261,N_16578);
and UO_2080 (O_2080,N_15150,N_19826);
or UO_2081 (O_2081,N_15231,N_16011);
and UO_2082 (O_2082,N_17193,N_19889);
nor UO_2083 (O_2083,N_19080,N_16164);
nand UO_2084 (O_2084,N_15932,N_17291);
and UO_2085 (O_2085,N_18851,N_15602);
nand UO_2086 (O_2086,N_15512,N_15587);
nor UO_2087 (O_2087,N_19109,N_17446);
nor UO_2088 (O_2088,N_16124,N_16385);
nor UO_2089 (O_2089,N_17684,N_18804);
nor UO_2090 (O_2090,N_15607,N_19123);
nand UO_2091 (O_2091,N_19393,N_19311);
nor UO_2092 (O_2092,N_15436,N_17450);
and UO_2093 (O_2093,N_19565,N_19107);
nor UO_2094 (O_2094,N_17940,N_18051);
nand UO_2095 (O_2095,N_15398,N_19570);
nor UO_2096 (O_2096,N_17810,N_15816);
nand UO_2097 (O_2097,N_15311,N_17593);
nand UO_2098 (O_2098,N_19831,N_19579);
nand UO_2099 (O_2099,N_16255,N_18262);
nand UO_2100 (O_2100,N_15251,N_18556);
nand UO_2101 (O_2101,N_17818,N_19140);
and UO_2102 (O_2102,N_16077,N_15120);
or UO_2103 (O_2103,N_15510,N_16800);
and UO_2104 (O_2104,N_16396,N_15827);
or UO_2105 (O_2105,N_18296,N_18224);
nor UO_2106 (O_2106,N_16883,N_16493);
nand UO_2107 (O_2107,N_16221,N_19141);
and UO_2108 (O_2108,N_15281,N_19015);
or UO_2109 (O_2109,N_16511,N_19914);
nor UO_2110 (O_2110,N_15050,N_16733);
or UO_2111 (O_2111,N_17839,N_16991);
nand UO_2112 (O_2112,N_15155,N_18026);
or UO_2113 (O_2113,N_17639,N_17016);
and UO_2114 (O_2114,N_15705,N_18464);
or UO_2115 (O_2115,N_15219,N_15350);
nand UO_2116 (O_2116,N_18716,N_17324);
nand UO_2117 (O_2117,N_19489,N_19129);
nor UO_2118 (O_2118,N_18987,N_18078);
or UO_2119 (O_2119,N_17045,N_19464);
or UO_2120 (O_2120,N_16137,N_16569);
or UO_2121 (O_2121,N_19310,N_16401);
and UO_2122 (O_2122,N_16952,N_16751);
nand UO_2123 (O_2123,N_16656,N_18092);
nand UO_2124 (O_2124,N_16088,N_19478);
xnor UO_2125 (O_2125,N_19860,N_17686);
nand UO_2126 (O_2126,N_15905,N_19186);
and UO_2127 (O_2127,N_18043,N_18429);
nor UO_2128 (O_2128,N_18286,N_15275);
or UO_2129 (O_2129,N_18861,N_18570);
nor UO_2130 (O_2130,N_16771,N_18740);
nand UO_2131 (O_2131,N_18632,N_16365);
or UO_2132 (O_2132,N_17611,N_19833);
or UO_2133 (O_2133,N_16062,N_18568);
nor UO_2134 (O_2134,N_17673,N_19086);
nor UO_2135 (O_2135,N_15845,N_19700);
and UO_2136 (O_2136,N_19881,N_16928);
or UO_2137 (O_2137,N_17698,N_17255);
or UO_2138 (O_2138,N_16389,N_19576);
nor UO_2139 (O_2139,N_19726,N_17746);
nor UO_2140 (O_2140,N_17244,N_17212);
nor UO_2141 (O_2141,N_18252,N_16014);
or UO_2142 (O_2142,N_19749,N_17304);
and UO_2143 (O_2143,N_19602,N_18313);
nand UO_2144 (O_2144,N_17143,N_17629);
or UO_2145 (O_2145,N_17999,N_17545);
nor UO_2146 (O_2146,N_15214,N_15186);
nand UO_2147 (O_2147,N_19509,N_19556);
nand UO_2148 (O_2148,N_16507,N_15292);
or UO_2149 (O_2149,N_16281,N_15988);
nand UO_2150 (O_2150,N_15674,N_17257);
nor UO_2151 (O_2151,N_15980,N_15879);
and UO_2152 (O_2152,N_19822,N_16830);
or UO_2153 (O_2153,N_15538,N_17491);
or UO_2154 (O_2154,N_18358,N_16094);
nand UO_2155 (O_2155,N_15875,N_17784);
nor UO_2156 (O_2156,N_17964,N_18165);
nand UO_2157 (O_2157,N_15077,N_19160);
nor UO_2158 (O_2158,N_15285,N_17847);
nor UO_2159 (O_2159,N_15344,N_17125);
or UO_2160 (O_2160,N_15290,N_18612);
and UO_2161 (O_2161,N_19099,N_18110);
nor UO_2162 (O_2162,N_18354,N_16900);
or UO_2163 (O_2163,N_15810,N_18874);
nor UO_2164 (O_2164,N_18249,N_15967);
and UO_2165 (O_2165,N_15455,N_19150);
or UO_2166 (O_2166,N_18734,N_18872);
nand UO_2167 (O_2167,N_16144,N_16314);
nor UO_2168 (O_2168,N_17694,N_16519);
nand UO_2169 (O_2169,N_16667,N_16001);
or UO_2170 (O_2170,N_15590,N_16835);
nand UO_2171 (O_2171,N_19737,N_17441);
nor UO_2172 (O_2172,N_18373,N_16587);
and UO_2173 (O_2173,N_18673,N_15847);
xnor UO_2174 (O_2174,N_16512,N_19425);
xnor UO_2175 (O_2175,N_17809,N_17222);
and UO_2176 (O_2176,N_17887,N_17161);
nor UO_2177 (O_2177,N_17524,N_15852);
and UO_2178 (O_2178,N_15801,N_16705);
and UO_2179 (O_2179,N_17311,N_18977);
nand UO_2180 (O_2180,N_18779,N_16481);
nor UO_2181 (O_2181,N_16508,N_17356);
nor UO_2182 (O_2182,N_18552,N_16914);
and UO_2183 (O_2183,N_16639,N_15283);
or UO_2184 (O_2184,N_15199,N_19396);
or UO_2185 (O_2185,N_17822,N_17082);
nand UO_2186 (O_2186,N_18052,N_17128);
nand UO_2187 (O_2187,N_15439,N_18489);
nor UO_2188 (O_2188,N_16049,N_15778);
and UO_2189 (O_2189,N_17642,N_17137);
and UO_2190 (O_2190,N_15842,N_16814);
nand UO_2191 (O_2191,N_19394,N_19390);
or UO_2192 (O_2192,N_19449,N_18014);
and UO_2193 (O_2193,N_18567,N_17054);
nor UO_2194 (O_2194,N_16601,N_15792);
or UO_2195 (O_2195,N_18236,N_16946);
nor UO_2196 (O_2196,N_18639,N_18709);
or UO_2197 (O_2197,N_18948,N_19722);
nor UO_2198 (O_2198,N_16217,N_16422);
nor UO_2199 (O_2199,N_15912,N_15661);
nand UO_2200 (O_2200,N_17106,N_15738);
or UO_2201 (O_2201,N_19381,N_16046);
or UO_2202 (O_2202,N_16924,N_16650);
or UO_2203 (O_2203,N_19020,N_17138);
xnor UO_2204 (O_2204,N_18826,N_15100);
nand UO_2205 (O_2205,N_15722,N_15195);
xnor UO_2206 (O_2206,N_19752,N_16285);
nand UO_2207 (O_2207,N_18793,N_16017);
nor UO_2208 (O_2208,N_19118,N_15262);
nand UO_2209 (O_2209,N_15486,N_18248);
and UO_2210 (O_2210,N_15215,N_17606);
nor UO_2211 (O_2211,N_18610,N_16756);
and UO_2212 (O_2212,N_15447,N_18187);
nor UO_2213 (O_2213,N_19220,N_17141);
and UO_2214 (O_2214,N_19545,N_18024);
or UO_2215 (O_2215,N_15825,N_19784);
or UO_2216 (O_2216,N_19932,N_16672);
or UO_2217 (O_2217,N_18432,N_18355);
and UO_2218 (O_2218,N_16134,N_16409);
and UO_2219 (O_2219,N_19074,N_19791);
or UO_2220 (O_2220,N_15995,N_16410);
nand UO_2221 (O_2221,N_18428,N_19656);
and UO_2222 (O_2222,N_18162,N_19439);
nand UO_2223 (O_2223,N_18924,N_17209);
nand UO_2224 (O_2224,N_19360,N_19158);
and UO_2225 (O_2225,N_16358,N_18016);
and UO_2226 (O_2226,N_19328,N_17420);
nand UO_2227 (O_2227,N_16696,N_18838);
nor UO_2228 (O_2228,N_17386,N_19236);
or UO_2229 (O_2229,N_15525,N_15862);
and UO_2230 (O_2230,N_15476,N_18822);
and UO_2231 (O_2231,N_18792,N_16868);
nor UO_2232 (O_2232,N_19345,N_19948);
nand UO_2233 (O_2233,N_18181,N_17021);
nand UO_2234 (O_2234,N_15230,N_16278);
nand UO_2235 (O_2235,N_18771,N_18004);
or UO_2236 (O_2236,N_18345,N_17820);
or UO_2237 (O_2237,N_16040,N_18431);
and UO_2238 (O_2238,N_19679,N_18686);
or UO_2239 (O_2239,N_16588,N_17428);
and UO_2240 (O_2240,N_18030,N_18406);
and UO_2241 (O_2241,N_16372,N_16203);
nor UO_2242 (O_2242,N_17453,N_15907);
nand UO_2243 (O_2243,N_17879,N_15484);
or UO_2244 (O_2244,N_18057,N_16572);
nand UO_2245 (O_2245,N_17432,N_15488);
nand UO_2246 (O_2246,N_19155,N_15950);
nand UO_2247 (O_2247,N_19437,N_16933);
and UO_2248 (O_2248,N_18467,N_19287);
or UO_2249 (O_2249,N_17301,N_15463);
nor UO_2250 (O_2250,N_19925,N_18808);
and UO_2251 (O_2251,N_18852,N_18487);
nor UO_2252 (O_2252,N_15928,N_18185);
nand UO_2253 (O_2253,N_18146,N_16497);
or UO_2254 (O_2254,N_16440,N_15618);
nor UO_2255 (O_2255,N_17481,N_19529);
nor UO_2256 (O_2256,N_18427,N_16249);
or UO_2257 (O_2257,N_18575,N_15384);
nor UO_2258 (O_2258,N_16760,N_17922);
nand UO_2259 (O_2259,N_16585,N_16528);
nor UO_2260 (O_2260,N_15177,N_18056);
nor UO_2261 (O_2261,N_17492,N_16590);
and UO_2262 (O_2262,N_16083,N_16608);
nand UO_2263 (O_2263,N_19547,N_19899);
or UO_2264 (O_2264,N_15952,N_19572);
and UO_2265 (O_2265,N_16887,N_17107);
and UO_2266 (O_2266,N_19745,N_18794);
nor UO_2267 (O_2267,N_16426,N_16971);
nor UO_2268 (O_2268,N_15291,N_19224);
nor UO_2269 (O_2269,N_17737,N_18274);
and UO_2270 (O_2270,N_16803,N_18253);
nand UO_2271 (O_2271,N_19255,N_18374);
or UO_2272 (O_2272,N_16852,N_17536);
nor UO_2273 (O_2273,N_17800,N_19741);
or UO_2274 (O_2274,N_19053,N_19657);
and UO_2275 (O_2275,N_15138,N_19930);
and UO_2276 (O_2276,N_18621,N_15272);
and UO_2277 (O_2277,N_15147,N_18569);
nand UO_2278 (O_2278,N_15183,N_15083);
and UO_2279 (O_2279,N_15079,N_16464);
or UO_2280 (O_2280,N_15813,N_15323);
nor UO_2281 (O_2281,N_18931,N_18123);
nand UO_2282 (O_2282,N_17972,N_19785);
nand UO_2283 (O_2283,N_18121,N_16844);
nor UO_2284 (O_2284,N_18479,N_17426);
nor UO_2285 (O_2285,N_16494,N_18763);
or UO_2286 (O_2286,N_15786,N_19365);
nor UO_2287 (O_2287,N_16743,N_15157);
and UO_2288 (O_2288,N_15854,N_16036);
and UO_2289 (O_2289,N_17339,N_15728);
or UO_2290 (O_2290,N_16807,N_19434);
nand UO_2291 (O_2291,N_16938,N_15573);
nor UO_2292 (O_2292,N_18857,N_17423);
nor UO_2293 (O_2293,N_18833,N_15299);
nor UO_2294 (O_2294,N_19882,N_18647);
nor UO_2295 (O_2295,N_18706,N_18616);
or UO_2296 (O_2296,N_15793,N_18450);
and UO_2297 (O_2297,N_18637,N_19666);
nand UO_2298 (O_2298,N_17325,N_16304);
and UO_2299 (O_2299,N_18565,N_19577);
or UO_2300 (O_2300,N_19533,N_16607);
nand UO_2301 (O_2301,N_18410,N_16028);
and UO_2302 (O_2302,N_16095,N_18062);
nand UO_2303 (O_2303,N_16349,N_16042);
nand UO_2304 (O_2304,N_18168,N_15897);
or UO_2305 (O_2305,N_16032,N_15753);
and UO_2306 (O_2306,N_18801,N_19585);
and UO_2307 (O_2307,N_16960,N_19663);
nand UO_2308 (O_2308,N_15569,N_15294);
and UO_2309 (O_2309,N_19940,N_15788);
nor UO_2310 (O_2310,N_17286,N_19443);
and UO_2311 (O_2311,N_16989,N_18160);
nor UO_2312 (O_2312,N_18287,N_19383);
nor UO_2313 (O_2313,N_16476,N_19111);
nand UO_2314 (O_2314,N_19329,N_16045);
or UO_2315 (O_2315,N_19367,N_18325);
or UO_2316 (O_2316,N_19755,N_18041);
or UO_2317 (O_2317,N_17480,N_16689);
and UO_2318 (O_2318,N_15670,N_16466);
and UO_2319 (O_2319,N_19965,N_19516);
or UO_2320 (O_2320,N_18813,N_17055);
or UO_2321 (O_2321,N_15194,N_15127);
or UO_2322 (O_2322,N_17292,N_17010);
nand UO_2323 (O_2323,N_18340,N_16142);
or UO_2324 (O_2324,N_15411,N_17134);
nor UO_2325 (O_2325,N_18750,N_17071);
and UO_2326 (O_2326,N_17738,N_16666);
and UO_2327 (O_2327,N_19797,N_18982);
nand UO_2328 (O_2328,N_17230,N_15947);
and UO_2329 (O_2329,N_16293,N_19161);
and UO_2330 (O_2330,N_19260,N_17861);
nor UO_2331 (O_2331,N_17444,N_15978);
nor UO_2332 (O_2332,N_17842,N_17978);
and UO_2333 (O_2333,N_18415,N_16187);
nand UO_2334 (O_2334,N_18020,N_18362);
nand UO_2335 (O_2335,N_18435,N_16305);
nand UO_2336 (O_2336,N_18684,N_18773);
nand UO_2337 (O_2337,N_18238,N_18708);
nand UO_2338 (O_2338,N_19591,N_19184);
and UO_2339 (O_2339,N_18594,N_19177);
nand UO_2340 (O_2340,N_17435,N_16149);
and UO_2341 (O_2341,N_16054,N_16904);
nor UO_2342 (O_2342,N_16892,N_19340);
nand UO_2343 (O_2343,N_18733,N_18626);
or UO_2344 (O_2344,N_16769,N_17723);
nor UO_2345 (O_2345,N_17769,N_19810);
and UO_2346 (O_2346,N_16120,N_16185);
and UO_2347 (O_2347,N_17837,N_16864);
and UO_2348 (O_2348,N_18085,N_19475);
nor UO_2349 (O_2349,N_18494,N_19104);
nand UO_2350 (O_2350,N_19953,N_15045);
or UO_2351 (O_2351,N_19254,N_15682);
nand UO_2352 (O_2352,N_19077,N_17640);
nor UO_2353 (O_2353,N_17040,N_17802);
and UO_2354 (O_2354,N_16567,N_17547);
nand UO_2355 (O_2355,N_17080,N_15580);
nor UO_2356 (O_2356,N_16704,N_15468);
or UO_2357 (O_2357,N_15725,N_16895);
nor UO_2358 (O_2358,N_16676,N_17340);
and UO_2359 (O_2359,N_18922,N_17674);
and UO_2360 (O_2360,N_15156,N_17319);
or UO_2361 (O_2361,N_17670,N_17364);
or UO_2362 (O_2362,N_19660,N_19697);
and UO_2363 (O_2363,N_16100,N_15528);
and UO_2364 (O_2364,N_16514,N_17576);
or UO_2365 (O_2365,N_17051,N_19624);
or UO_2366 (O_2366,N_17148,N_15732);
nand UO_2367 (O_2367,N_15684,N_17914);
nand UO_2368 (O_2368,N_17416,N_19757);
or UO_2369 (O_2369,N_18378,N_17511);
or UO_2370 (O_2370,N_19759,N_18418);
or UO_2371 (O_2371,N_16506,N_18844);
nor UO_2372 (O_2372,N_19288,N_18582);
or UO_2373 (O_2373,N_17414,N_15041);
or UO_2374 (O_2374,N_16411,N_19094);
and UO_2375 (O_2375,N_15416,N_19878);
nand UO_2376 (O_2376,N_17044,N_18339);
and UO_2377 (O_2377,N_15233,N_19796);
nand UO_2378 (O_2378,N_19436,N_16237);
nor UO_2379 (O_2379,N_16721,N_15222);
nor UO_2380 (O_2380,N_18938,N_15535);
nor UO_2381 (O_2381,N_15560,N_17035);
nor UO_2382 (O_2382,N_18303,N_16199);
nand UO_2383 (O_2383,N_16256,N_17519);
or UO_2384 (O_2384,N_15700,N_17467);
nand UO_2385 (O_2385,N_18459,N_16050);
nor UO_2386 (O_2386,N_19600,N_15748);
nor UO_2387 (O_2387,N_16735,N_19072);
nand UO_2388 (O_2388,N_18207,N_18839);
nand UO_2389 (O_2389,N_17906,N_19972);
and UO_2390 (O_2390,N_16452,N_19803);
or UO_2391 (O_2391,N_15336,N_16330);
nor UO_2392 (O_2392,N_17431,N_17219);
nand UO_2393 (O_2393,N_19825,N_19059);
nand UO_2394 (O_2394,N_18615,N_16849);
or UO_2395 (O_2395,N_18346,N_19848);
or UO_2396 (O_2396,N_16129,N_19320);
and UO_2397 (O_2397,N_19106,N_18022);
and UO_2398 (O_2398,N_15263,N_19558);
and UO_2399 (O_2399,N_19349,N_17263);
nand UO_2400 (O_2400,N_19684,N_16331);
nand UO_2401 (O_2401,N_19500,N_16277);
or UO_2402 (O_2402,N_16259,N_18037);
or UO_2403 (O_2403,N_16329,N_18377);
and UO_2404 (O_2404,N_16283,N_17095);
and UO_2405 (O_2405,N_15414,N_19721);
nor UO_2406 (O_2406,N_15377,N_19870);
and UO_2407 (O_2407,N_18949,N_16013);
and UO_2408 (O_2408,N_16719,N_18963);
nor UO_2409 (O_2409,N_17419,N_15059);
nand UO_2410 (O_2410,N_17118,N_17836);
nor UO_2411 (O_2411,N_17360,N_15165);
and UO_2412 (O_2412,N_18382,N_15731);
nor UO_2413 (O_2413,N_19298,N_18229);
and UO_2414 (O_2414,N_18961,N_16592);
or UO_2415 (O_2415,N_17477,N_18736);
nor UO_2416 (O_2416,N_16973,N_18279);
nand UO_2417 (O_2417,N_15516,N_17262);
nor UO_2418 (O_2418,N_15355,N_17829);
and UO_2419 (O_2419,N_17954,N_16469);
and UO_2420 (O_2420,N_15029,N_19510);
nand UO_2421 (O_2421,N_17204,N_16910);
and UO_2422 (O_2422,N_17730,N_16326);
or UO_2423 (O_2423,N_17712,N_16116);
nor UO_2424 (O_2424,N_16851,N_15755);
nor UO_2425 (O_2425,N_19631,N_18721);
and UO_2426 (O_2426,N_17676,N_17281);
or UO_2427 (O_2427,N_17357,N_15208);
nand UO_2428 (O_2428,N_15809,N_15185);
or UO_2429 (O_2429,N_19676,N_18964);
or UO_2430 (O_2430,N_18143,N_15985);
or UO_2431 (O_2431,N_19845,N_16115);
nor UO_2432 (O_2432,N_16169,N_17625);
or UO_2433 (O_2433,N_18509,N_17683);
and UO_2434 (O_2434,N_17665,N_15939);
nand UO_2435 (O_2435,N_16893,N_15051);
nand UO_2436 (O_2436,N_15116,N_19274);
nand UO_2437 (O_2437,N_19967,N_19145);
or UO_2438 (O_2438,N_17424,N_15571);
nor UO_2439 (O_2439,N_19599,N_18667);
nand UO_2440 (O_2440,N_16337,N_18911);
or UO_2441 (O_2441,N_19566,N_15490);
nand UO_2442 (O_2442,N_19454,N_19134);
nand UO_2443 (O_2443,N_16937,N_17803);
nand UO_2444 (O_2444,N_15591,N_18696);
and UO_2445 (O_2445,N_15973,N_18654);
nor UO_2446 (O_2446,N_19961,N_18005);
or UO_2447 (O_2447,N_16872,N_15884);
nand UO_2448 (O_2448,N_17363,N_18204);
or UO_2449 (O_2449,N_17046,N_16111);
nor UO_2450 (O_2450,N_15367,N_15176);
nor UO_2451 (O_2451,N_18515,N_19685);
or UO_2452 (O_2452,N_15534,N_18111);
or UO_2453 (O_2453,N_17131,N_17308);
or UO_2454 (O_2454,N_15430,N_18323);
nor UO_2455 (O_2455,N_18201,N_15987);
nand UO_2456 (O_2456,N_18074,N_16873);
or UO_2457 (O_2457,N_18800,N_17333);
nor UO_2458 (O_2458,N_17823,N_15581);
and UO_2459 (O_2459,N_17563,N_17812);
and UO_2460 (O_2460,N_19792,N_19181);
and UO_2461 (O_2461,N_17465,N_19200);
nor UO_2462 (O_2462,N_18413,N_18960);
and UO_2463 (O_2463,N_16243,N_19297);
or UO_2464 (O_2464,N_16712,N_19314);
and UO_2465 (O_2465,N_19581,N_19348);
nor UO_2466 (O_2466,N_19525,N_16841);
and UO_2467 (O_2467,N_15451,N_16774);
and UO_2468 (O_2468,N_18120,N_19526);
and UO_2469 (O_2469,N_15572,N_18112);
nand UO_2470 (O_2470,N_19662,N_16561);
nand UO_2471 (O_2471,N_18048,N_19133);
nand UO_2472 (O_2472,N_16545,N_18337);
nand UO_2473 (O_2473,N_17494,N_18128);
and UO_2474 (O_2474,N_16878,N_18529);
nand UO_2475 (O_2475,N_16457,N_19505);
nor UO_2476 (O_2476,N_18904,N_17716);
xor UO_2477 (O_2477,N_15389,N_19102);
and UO_2478 (O_2478,N_16789,N_16939);
and UO_2479 (O_2479,N_19691,N_18114);
or UO_2480 (O_2480,N_16755,N_19799);
and UO_2481 (O_2481,N_15951,N_17590);
nor UO_2482 (O_2482,N_15088,N_15612);
nand UO_2483 (O_2483,N_18775,N_16320);
and UO_2484 (O_2484,N_15720,N_18531);
and UO_2485 (O_2485,N_17719,N_17896);
or UO_2486 (O_2486,N_17190,N_16653);
nand UO_2487 (O_2487,N_18955,N_16911);
nor UO_2488 (O_2488,N_18944,N_15143);
and UO_2489 (O_2489,N_19995,N_19049);
or UO_2490 (O_2490,N_16252,N_19709);
or UO_2491 (O_2491,N_18379,N_18996);
nand UO_2492 (O_2492,N_16881,N_16649);
nor UO_2493 (O_2493,N_18113,N_19336);
and UO_2494 (O_2494,N_16058,N_18999);
nor UO_2495 (O_2495,N_19813,N_18650);
or UO_2496 (O_2496,N_18544,N_18756);
or UO_2497 (O_2497,N_16344,N_18045);
nor UO_2498 (O_2498,N_19027,N_18466);
nor UO_2499 (O_2499,N_19284,N_18576);
endmodule