module basic_1000_10000_1500_50_levels_10xor_1(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999;
xnor U0 (N_0,In_760,In_612);
and U1 (N_1,In_295,In_347);
nor U2 (N_2,In_616,In_134);
or U3 (N_3,In_31,In_702);
xnor U4 (N_4,In_706,In_653);
or U5 (N_5,In_609,In_438);
or U6 (N_6,In_276,In_499);
nor U7 (N_7,In_819,In_376);
or U8 (N_8,In_326,In_696);
and U9 (N_9,In_593,In_88);
nand U10 (N_10,In_373,In_838);
nand U11 (N_11,In_816,In_130);
nor U12 (N_12,In_607,In_308);
nand U13 (N_13,In_492,In_414);
nor U14 (N_14,In_305,In_666);
and U15 (N_15,In_747,In_831);
or U16 (N_16,In_823,In_493);
xor U17 (N_17,In_287,In_721);
nor U18 (N_18,In_193,In_79);
or U19 (N_19,In_942,In_695);
and U20 (N_20,In_58,In_476);
nor U21 (N_21,In_210,In_804);
nand U22 (N_22,In_788,In_313);
xnor U23 (N_23,In_230,In_726);
and U24 (N_24,In_524,In_146);
or U25 (N_25,In_681,In_581);
nand U26 (N_26,In_453,In_885);
xor U27 (N_27,In_328,In_754);
or U28 (N_28,In_163,In_660);
and U29 (N_29,In_259,In_181);
nor U30 (N_30,In_899,In_14);
or U31 (N_31,In_461,In_446);
xor U32 (N_32,In_997,In_97);
xor U33 (N_33,In_106,In_893);
nand U34 (N_34,In_472,In_950);
nand U35 (N_35,In_491,In_474);
nor U36 (N_36,In_393,In_201);
and U37 (N_37,In_458,In_693);
and U38 (N_38,In_68,In_521);
xor U39 (N_39,In_519,In_473);
and U40 (N_40,In_451,In_84);
xor U41 (N_41,In_735,In_741);
or U42 (N_42,In_686,In_140);
nor U43 (N_43,In_963,In_535);
nor U44 (N_44,In_711,In_80);
and U45 (N_45,In_656,In_209);
nand U46 (N_46,In_763,In_150);
nand U47 (N_47,In_759,In_452);
or U48 (N_48,In_707,In_9);
or U49 (N_49,In_918,In_18);
and U50 (N_50,In_24,In_489);
or U51 (N_51,In_306,In_20);
or U52 (N_52,In_176,In_537);
or U53 (N_53,In_590,In_868);
nand U54 (N_54,In_188,In_319);
and U55 (N_55,In_157,In_538);
xor U56 (N_56,In_278,In_813);
nand U57 (N_57,In_239,In_636);
and U58 (N_58,In_516,In_737);
or U59 (N_59,In_664,In_575);
xor U60 (N_60,In_485,In_620);
or U61 (N_61,In_121,In_301);
nand U62 (N_62,In_40,In_783);
or U63 (N_63,In_951,In_113);
xor U64 (N_64,In_90,In_646);
nand U65 (N_65,In_290,In_345);
nor U66 (N_66,In_947,In_95);
and U67 (N_67,In_3,In_714);
or U68 (N_68,In_954,In_606);
or U69 (N_69,In_513,In_862);
and U70 (N_70,In_882,In_333);
or U71 (N_71,In_829,In_17);
nor U72 (N_72,In_404,In_228);
and U73 (N_73,In_247,In_559);
or U74 (N_74,In_423,In_520);
or U75 (N_75,In_204,In_526);
and U76 (N_76,In_49,In_381);
xnor U77 (N_77,In_975,In_149);
nor U78 (N_78,In_124,In_43);
or U79 (N_79,In_943,In_488);
or U80 (N_80,In_985,In_625);
or U81 (N_81,In_350,In_628);
and U82 (N_82,In_256,In_967);
nand U83 (N_83,In_322,In_314);
nor U84 (N_84,In_364,In_530);
xor U85 (N_85,In_263,In_57);
nor U86 (N_86,In_953,In_850);
and U87 (N_87,In_379,In_733);
nand U88 (N_88,In_812,In_502);
or U89 (N_89,In_802,In_396);
nor U90 (N_90,In_361,In_743);
xnor U91 (N_91,In_403,In_839);
nor U92 (N_92,In_861,In_155);
and U93 (N_93,In_425,In_131);
nor U94 (N_94,In_969,In_260);
or U95 (N_95,In_731,In_938);
and U96 (N_96,In_728,In_678);
xnor U97 (N_97,In_591,In_10);
or U98 (N_98,In_2,In_346);
xnor U99 (N_99,In_349,In_481);
nand U100 (N_100,In_398,In_486);
nor U101 (N_101,In_145,In_320);
nor U102 (N_102,In_37,In_872);
or U103 (N_103,In_164,In_633);
and U104 (N_104,In_991,In_303);
nand U105 (N_105,In_649,In_337);
or U106 (N_106,In_53,In_236);
and U107 (N_107,In_579,In_470);
nor U108 (N_108,In_156,In_500);
xor U109 (N_109,In_927,In_198);
or U110 (N_110,In_42,In_920);
xor U111 (N_111,In_915,In_577);
or U112 (N_112,In_852,In_223);
and U113 (N_113,In_662,In_237);
or U114 (N_114,In_922,In_51);
and U115 (N_115,In_116,In_832);
or U116 (N_116,In_898,In_460);
xor U117 (N_117,In_801,In_264);
nor U118 (N_118,In_830,In_439);
nand U119 (N_119,In_744,In_761);
xnor U120 (N_120,In_317,In_98);
and U121 (N_121,In_610,In_136);
nand U122 (N_122,In_548,In_187);
xnor U123 (N_123,In_677,In_386);
nor U124 (N_124,In_498,In_454);
xnor U125 (N_125,In_907,In_689);
nand U126 (N_126,In_336,In_279);
and U127 (N_127,In_652,In_160);
or U128 (N_128,In_367,In_244);
or U129 (N_129,In_261,In_117);
nor U130 (N_130,In_22,In_304);
nor U131 (N_131,In_369,In_529);
nand U132 (N_132,In_478,In_874);
and U133 (N_133,In_151,In_688);
or U134 (N_134,In_494,In_400);
nand U135 (N_135,In_437,In_974);
and U136 (N_136,In_856,In_551);
nor U137 (N_137,In_430,In_341);
and U138 (N_138,In_307,In_252);
or U139 (N_139,In_762,In_30);
nand U140 (N_140,In_23,In_324);
nand U141 (N_141,In_642,In_72);
nand U142 (N_142,In_700,In_509);
and U143 (N_143,In_573,In_148);
or U144 (N_144,In_45,In_385);
and U145 (N_145,In_343,In_528);
nand U146 (N_146,In_335,In_890);
nor U147 (N_147,In_797,In_576);
or U148 (N_148,In_701,In_296);
or U149 (N_149,In_709,In_312);
or U150 (N_150,In_175,In_374);
nor U151 (N_151,In_420,In_195);
nand U152 (N_152,In_266,In_826);
xor U153 (N_153,In_558,In_986);
nand U154 (N_154,In_318,In_869);
xnor U155 (N_155,In_909,In_756);
or U156 (N_156,In_771,In_299);
and U157 (N_157,In_128,In_183);
and U158 (N_158,In_758,In_571);
xnor U159 (N_159,In_232,In_705);
nor U160 (N_160,In_178,In_387);
or U161 (N_161,In_723,In_253);
nor U162 (N_162,In_370,In_545);
nand U163 (N_163,In_574,In_680);
and U164 (N_164,In_397,In_311);
and U165 (N_165,In_41,In_618);
xor U166 (N_166,In_123,In_732);
and U167 (N_167,In_557,In_196);
xnor U168 (N_168,In_354,In_879);
or U169 (N_169,In_778,In_93);
or U170 (N_170,In_162,In_29);
and U171 (N_171,In_566,In_358);
and U172 (N_172,In_791,In_837);
and U173 (N_173,In_101,In_89);
and U174 (N_174,In_300,In_977);
xor U175 (N_175,In_685,In_836);
or U176 (N_176,In_125,In_623);
and U177 (N_177,In_392,In_621);
nor U178 (N_178,In_543,In_399);
nand U179 (N_179,In_217,In_380);
nor U180 (N_180,In_940,In_456);
nand U181 (N_181,In_627,In_988);
xnor U182 (N_182,In_939,In_592);
or U183 (N_183,In_382,In_608);
or U184 (N_184,In_567,In_817);
nand U185 (N_185,In_442,In_600);
nand U186 (N_186,In_613,In_746);
nor U187 (N_187,In_448,In_959);
nor U188 (N_188,In_161,In_325);
xor U189 (N_189,In_233,In_866);
nand U190 (N_190,In_835,In_365);
xor U191 (N_191,In_873,In_497);
nor U192 (N_192,In_539,In_824);
and U193 (N_193,In_888,In_171);
xor U194 (N_194,In_235,In_34);
nor U195 (N_195,In_434,In_903);
nor U196 (N_196,In_805,In_841);
and U197 (N_197,In_806,In_378);
nor U198 (N_198,In_993,In_703);
nor U199 (N_199,In_546,In_968);
xnor U200 (N_200,N_174,In_562);
xor U201 (N_201,N_163,In_415);
nand U202 (N_202,In_135,In_902);
xnor U203 (N_203,N_54,In_989);
nor U204 (N_204,In_471,In_202);
nand U205 (N_205,N_92,In_26);
xnor U206 (N_206,N_2,In_243);
nand U207 (N_207,In_821,In_441);
or U208 (N_208,In_203,In_348);
nor U209 (N_209,In_858,In_933);
nor U210 (N_210,N_139,In_540);
nand U211 (N_211,N_196,In_147);
and U212 (N_212,In_930,In_199);
nand U213 (N_213,In_738,N_192);
or U214 (N_214,In_614,N_162);
nand U215 (N_215,In_923,In_883);
nor U216 (N_216,In_409,In_739);
or U217 (N_217,In_377,In_443);
nor U218 (N_218,In_224,In_487);
or U219 (N_219,N_38,In_691);
nand U220 (N_220,N_125,In_76);
nor U221 (N_221,In_867,In_725);
or U222 (N_222,N_71,N_48);
nand U223 (N_223,In_139,In_670);
nor U224 (N_224,In_651,In_775);
or U225 (N_225,In_271,In_958);
and U226 (N_226,N_183,In_784);
nand U227 (N_227,In_25,N_143);
and U228 (N_228,N_36,In_925);
and U229 (N_229,In_798,N_42);
nor U230 (N_230,In_871,In_191);
xnor U231 (N_231,N_103,In_605);
nor U232 (N_232,In_982,In_119);
or U233 (N_233,N_189,In_594);
xnor U234 (N_234,In_282,In_578);
nand U235 (N_235,N_101,In_745);
nor U236 (N_236,N_132,In_351);
nand U237 (N_237,In_483,In_766);
xor U238 (N_238,In_120,N_43);
nand U239 (N_239,N_146,In_190);
nand U240 (N_240,N_28,In_729);
xnor U241 (N_241,In_165,In_270);
xnor U242 (N_242,In_444,In_960);
nand U243 (N_243,N_83,N_124);
or U244 (N_244,In_583,In_197);
xnor U245 (N_245,In_129,N_138);
and U246 (N_246,N_93,In_362);
and U247 (N_247,In_822,In_904);
and U248 (N_248,N_69,N_170);
and U249 (N_249,N_47,In_973);
xor U250 (N_250,In_126,In_248);
or U251 (N_251,N_153,In_506);
and U252 (N_252,In_182,In_815);
nor U253 (N_253,In_15,In_684);
xor U254 (N_254,In_92,N_13);
or U255 (N_255,In_143,N_96);
and U256 (N_256,In_603,In_227);
or U257 (N_257,In_635,In_141);
nand U258 (N_258,In_615,In_955);
nor U259 (N_259,In_363,In_934);
or U260 (N_260,In_422,In_464);
nand U261 (N_261,In_366,In_168);
nand U262 (N_262,In_344,In_255);
or U263 (N_263,In_194,N_12);
nand U264 (N_264,In_727,In_792);
nand U265 (N_265,In_547,In_896);
xor U266 (N_266,In_748,In_643);
xor U267 (N_267,In_413,In_214);
nand U268 (N_268,N_4,In_914);
nor U269 (N_269,In_4,N_44);
nand U270 (N_270,In_112,In_172);
or U271 (N_271,In_211,In_807);
nor U272 (N_272,N_11,In_355);
and U273 (N_273,In_584,In_205);
nand U274 (N_274,In_421,In_769);
xor U275 (N_275,In_331,In_654);
nand U276 (N_276,In_19,In_556);
xnor U277 (N_277,In_818,In_949);
nand U278 (N_278,In_108,N_168);
and U279 (N_279,In_277,In_289);
or U280 (N_280,In_595,In_921);
xnor U281 (N_281,In_561,In_13);
or U282 (N_282,N_86,In_597);
and U283 (N_283,In_391,In_479);
xnor U284 (N_284,N_75,In_987);
and U285 (N_285,In_433,In_568);
nand U286 (N_286,In_668,In_360);
or U287 (N_287,In_842,In_375);
nand U288 (N_288,In_61,In_582);
nand U289 (N_289,In_269,In_440);
xnor U290 (N_290,N_193,In_814);
and U291 (N_291,N_131,In_657);
and U292 (N_292,In_436,N_166);
and U293 (N_293,N_19,In_327);
nor U294 (N_294,N_128,In_932);
nand U295 (N_295,In_262,N_187);
nand U296 (N_296,N_195,N_155);
or U297 (N_297,N_50,In_844);
and U298 (N_298,In_531,In_91);
xor U299 (N_299,In_697,In_752);
and U300 (N_300,N_41,In_412);
and U301 (N_301,In_699,In_704);
nor U302 (N_302,In_917,In_717);
xnor U303 (N_303,In_475,In_272);
nor U304 (N_304,In_589,In_38);
and U305 (N_305,N_30,In_808);
xor U306 (N_306,N_102,In_340);
nor U307 (N_307,N_58,In_669);
nand U308 (N_308,In_122,In_880);
and U309 (N_309,In_503,In_534);
nand U310 (N_310,In_523,N_45);
nand U311 (N_311,In_7,N_99);
or U312 (N_312,In_459,In_185);
or U313 (N_313,In_389,N_84);
xnor U314 (N_314,In_315,In_740);
nor U315 (N_315,N_154,In_994);
xnor U316 (N_316,In_514,In_667);
nand U317 (N_317,In_983,In_56);
nand U318 (N_318,In_127,In_332);
or U319 (N_319,In_937,In_972);
nor U320 (N_320,In_286,In_854);
nor U321 (N_321,N_29,In_601);
and U322 (N_322,N_180,In_417);
or U323 (N_323,In_833,In_109);
or U324 (N_324,N_35,N_0);
nor U325 (N_325,In_384,In_820);
xnor U326 (N_326,In_800,N_23);
nand U327 (N_327,In_881,In_901);
and U328 (N_328,N_57,N_191);
xnor U329 (N_329,In_411,N_70);
or U330 (N_330,N_16,In_637);
xor U331 (N_331,In_875,In_586);
xor U332 (N_332,In_12,In_103);
and U333 (N_333,In_225,N_39);
nand U334 (N_334,N_89,In_505);
nand U335 (N_335,In_48,In_77);
xor U336 (N_336,In_865,N_127);
and U337 (N_337,In_712,In_777);
nor U338 (N_338,In_406,In_734);
nor U339 (N_339,In_229,N_18);
or U340 (N_340,In_675,In_870);
nor U341 (N_341,In_970,In_794);
or U342 (N_342,In_560,In_876);
nand U343 (N_343,N_74,In_843);
nand U344 (N_344,In_710,In_447);
and U345 (N_345,In_995,In_142);
and U346 (N_346,In_27,In_477);
and U347 (N_347,In_787,In_294);
or U348 (N_348,In_268,In_517);
nand U349 (N_349,In_884,In_105);
nand U350 (N_350,In_357,In_465);
xor U351 (N_351,In_428,In_35);
and U352 (N_352,In_28,N_113);
nand U353 (N_353,In_795,In_848);
nand U354 (N_354,In_353,In_11);
or U355 (N_355,In_634,In_851);
nor U356 (N_356,In_418,In_170);
xor U357 (N_357,In_799,In_990);
or U358 (N_358,In_655,In_924);
and U359 (N_359,In_221,In_338);
xor U360 (N_360,N_110,N_120);
nand U361 (N_361,In_855,In_132);
xnor U362 (N_362,In_962,In_74);
or U363 (N_363,In_107,In_811);
nand U364 (N_364,In_796,In_179);
or U365 (N_365,N_56,In_8);
and U366 (N_366,In_144,In_889);
nor U367 (N_367,In_533,N_63);
nand U368 (N_368,N_53,N_179);
nand U369 (N_369,In_863,In_544);
and U370 (N_370,N_158,In_153);
or U371 (N_371,In_894,In_280);
nor U372 (N_372,In_877,N_165);
and U373 (N_373,In_274,In_267);
xnor U374 (N_374,In_281,In_75);
nor U375 (N_375,In_673,N_159);
and U376 (N_376,N_181,In_663);
nor U377 (N_377,N_134,In_218);
and U378 (N_378,N_91,In_192);
and U379 (N_379,N_136,In_644);
or U380 (N_380,In_356,In_152);
xor U381 (N_381,In_257,In_288);
and U382 (N_382,N_148,In_847);
xnor U383 (N_383,N_145,In_957);
nor U384 (N_384,In_55,N_33);
xor U385 (N_385,N_6,In_749);
and U386 (N_386,In_186,In_226);
nor U387 (N_387,In_944,In_480);
nor U388 (N_388,In_658,In_853);
and U389 (N_389,N_52,N_64);
and U390 (N_390,N_172,In_323);
or U391 (N_391,N_34,In_980);
nor U392 (N_392,In_39,In_694);
nor U393 (N_393,In_611,N_7);
and U394 (N_394,N_119,In_981);
and U395 (N_395,N_72,In_715);
nand U396 (N_396,In_81,In_878);
or U397 (N_397,In_115,In_978);
nor U398 (N_398,In_659,In_216);
nand U399 (N_399,In_553,In_240);
and U400 (N_400,N_368,N_353);
nor U401 (N_401,N_303,N_285);
and U402 (N_402,N_237,In_996);
and U403 (N_403,N_261,N_121);
and U404 (N_404,In_780,In_542);
nand U405 (N_405,N_130,N_321);
xnor U406 (N_406,In_522,N_325);
and U407 (N_407,In_383,In_432);
and U408 (N_408,In_212,In_5);
xnor U409 (N_409,N_256,N_314);
xor U410 (N_410,In_789,In_73);
and U411 (N_411,In_860,N_177);
nand U412 (N_412,N_278,In_309);
and U413 (N_413,N_308,N_333);
and U414 (N_414,In_219,N_253);
xnor U415 (N_415,N_240,N_306);
xor U416 (N_416,In_200,In_676);
and U417 (N_417,N_334,N_87);
nor U418 (N_418,N_32,N_222);
or U419 (N_419,In_588,In_82);
or U420 (N_420,In_50,N_197);
nor U421 (N_421,N_167,N_397);
nand U422 (N_422,In_463,In_207);
nor U423 (N_423,In_810,In_639);
xnor U424 (N_424,In_648,N_194);
and U425 (N_425,In_285,N_27);
and U426 (N_426,N_178,N_244);
and U427 (N_427,In_767,In_742);
nor U428 (N_428,In_864,In_541);
xor U429 (N_429,In_532,N_26);
and U430 (N_430,N_8,In_626);
or U431 (N_431,N_269,In_674);
and U432 (N_432,In_469,In_570);
xor U433 (N_433,In_1,N_272);
and U434 (N_434,In_773,In_231);
xnor U435 (N_435,N_383,In_114);
nand U436 (N_436,In_638,N_266);
xnor U437 (N_437,N_287,In_254);
or U438 (N_438,In_713,N_203);
or U439 (N_439,N_210,In_496);
xnor U440 (N_440,In_629,In_683);
and U441 (N_441,In_793,In_518);
nor U442 (N_442,N_310,In_755);
and U443 (N_443,N_1,N_219);
xnor U444 (N_444,N_280,N_396);
or U445 (N_445,N_296,N_14);
nand U446 (N_446,N_363,In_249);
nand U447 (N_447,N_298,N_216);
and U448 (N_448,N_384,In_661);
or U449 (N_449,In_215,N_270);
and U450 (N_450,N_336,N_141);
or U451 (N_451,In_647,In_297);
and U452 (N_452,In_999,In_405);
nand U453 (N_453,In_293,In_46);
nor U454 (N_454,N_346,In_342);
and U455 (N_455,In_897,In_587);
nor U456 (N_456,N_264,In_602);
xnor U457 (N_457,N_283,In_936);
nand U458 (N_458,In_54,In_310);
xor U459 (N_459,In_265,N_326);
xnor U460 (N_460,N_212,In_302);
or U461 (N_461,In_110,N_376);
nor U462 (N_462,In_402,N_263);
and U463 (N_463,N_289,In_359);
and U464 (N_464,In_408,In_585);
and U465 (N_465,N_67,In_419);
nand U466 (N_466,N_232,In_52);
xor U467 (N_467,In_913,In_16);
and U468 (N_468,In_912,In_66);
nor U469 (N_469,N_215,In_258);
and U470 (N_470,In_834,In_720);
and U471 (N_471,N_340,In_525);
or U472 (N_472,N_151,N_235);
nand U473 (N_473,In_78,N_271);
xnor U474 (N_474,In_329,In_671);
and U475 (N_475,N_5,N_273);
or U476 (N_476,N_312,In_490);
and U477 (N_477,In_782,N_169);
xnor U478 (N_478,In_827,N_351);
nand U479 (N_479,In_857,N_228);
and U480 (N_480,N_341,In_234);
nand U481 (N_481,In_554,N_284);
nor U482 (N_482,N_335,N_224);
nand U483 (N_483,N_372,N_239);
nand U484 (N_484,In_275,In_44);
or U485 (N_485,N_62,N_286);
and U486 (N_486,In_159,In_770);
or U487 (N_487,N_207,N_175);
nand U488 (N_488,N_374,In_273);
and U489 (N_489,In_722,N_316);
xnor U490 (N_490,N_343,N_186);
nand U491 (N_491,In_624,In_206);
and U492 (N_492,N_347,In_966);
or U493 (N_493,In_138,In_527);
nor U494 (N_494,In_251,In_250);
nor U495 (N_495,In_86,In_368);
nor U496 (N_496,In_736,In_569);
xnor U497 (N_497,In_118,In_846);
nand U498 (N_498,In_158,N_388);
or U499 (N_499,In_757,N_229);
or U500 (N_500,N_332,In_768);
nand U501 (N_501,In_410,N_78);
or U502 (N_502,N_60,In_772);
nor U503 (N_503,N_135,In_94);
nor U504 (N_504,In_424,N_288);
or U505 (N_505,In_926,In_785);
nand U506 (N_506,In_916,In_316);
nand U507 (N_507,In_65,In_512);
xor U508 (N_508,N_217,In_719);
or U509 (N_509,N_390,N_281);
xnor U510 (N_510,N_257,In_431);
nor U511 (N_511,In_462,In_36);
or U512 (N_512,In_565,N_22);
or U513 (N_513,In_753,In_395);
xor U514 (N_514,N_367,In_372);
nor U515 (N_515,N_152,N_137);
or U516 (N_516,In_809,N_160);
or U517 (N_517,N_129,In_32);
or U518 (N_518,N_277,N_25);
xnor U519 (N_519,N_249,N_399);
nand U520 (N_520,N_156,In_407);
or U521 (N_521,N_320,N_123);
nor U522 (N_522,In_632,N_323);
nand U523 (N_523,N_369,In_776);
or U524 (N_524,N_313,N_107);
and U525 (N_525,N_37,N_61);
nor U526 (N_526,N_90,In_99);
xor U527 (N_527,N_55,N_190);
and U528 (N_528,In_929,N_49);
or U529 (N_529,In_352,In_321);
or U530 (N_530,N_342,In_779);
xnor U531 (N_531,N_234,N_81);
and U532 (N_532,In_945,N_114);
nand U533 (N_533,N_381,N_20);
nor U534 (N_534,N_339,In_177);
and U535 (N_535,N_377,N_246);
or U536 (N_536,In_334,N_95);
or U537 (N_537,In_241,N_238);
xor U538 (N_538,In_572,In_946);
xnor U539 (N_539,N_149,In_672);
and U540 (N_540,N_21,N_360);
or U541 (N_541,N_295,In_450);
nor U542 (N_542,N_211,N_392);
xor U543 (N_543,N_327,In_803);
and U544 (N_544,In_935,In_222);
xor U545 (N_545,In_682,N_259);
nand U546 (N_546,N_115,In_515);
and U547 (N_547,N_199,N_225);
nor U548 (N_548,N_221,In_166);
nor U549 (N_549,N_389,In_948);
xnor U550 (N_550,In_774,In_435);
or U551 (N_551,In_455,In_941);
or U552 (N_552,N_100,N_337);
and U553 (N_553,N_366,N_248);
nor U554 (N_554,In_427,In_339);
xnor U555 (N_555,In_599,In_690);
and U556 (N_556,In_645,N_359);
and U557 (N_557,N_218,In_905);
xnor U558 (N_558,In_283,In_617);
and U559 (N_559,N_233,N_251);
and U560 (N_560,N_385,N_304);
or U561 (N_561,N_24,In_390);
xnor U562 (N_562,In_429,In_371);
nand U563 (N_563,In_906,N_393);
xnor U564 (N_564,N_362,N_147);
or U565 (N_565,N_324,N_164);
nor U566 (N_566,In_679,N_198);
xor U567 (N_567,In_900,N_208);
nand U568 (N_568,In_70,N_97);
nor U569 (N_569,In_828,N_395);
or U570 (N_570,N_202,In_781);
or U571 (N_571,In_965,In_174);
or U572 (N_572,N_209,In_640);
and U573 (N_573,N_394,In_484);
and U574 (N_574,N_220,In_388);
nor U575 (N_575,N_140,N_184);
or U576 (N_576,N_109,In_718);
nand U577 (N_577,N_322,N_204);
and U578 (N_578,In_908,In_507);
xnor U579 (N_579,N_213,N_260);
nor U580 (N_580,In_394,In_102);
nor U581 (N_581,In_549,In_887);
or U582 (N_582,N_242,N_82);
xor U583 (N_583,N_133,In_555);
and U584 (N_584,N_65,N_292);
nor U585 (N_585,In_137,N_302);
nand U586 (N_586,In_104,N_380);
or U587 (N_587,In_598,N_254);
nor U588 (N_588,In_298,N_144);
or U589 (N_589,N_373,N_10);
nand U590 (N_590,N_317,N_46);
and U591 (N_591,In_284,In_730);
nand U592 (N_592,In_563,In_100);
nor U593 (N_593,N_252,N_243);
xor U594 (N_594,In_665,N_227);
nor U595 (N_595,N_236,N_349);
nor U596 (N_596,N_77,N_267);
and U597 (N_597,N_223,In_495);
nor U598 (N_598,In_849,N_105);
nand U599 (N_599,N_173,In_167);
or U600 (N_600,N_427,In_63);
nor U601 (N_601,In_71,N_565);
and U602 (N_602,N_508,N_299);
or U603 (N_603,N_430,N_495);
and U604 (N_604,N_315,N_560);
xor U605 (N_605,N_398,N_421);
and U606 (N_606,N_450,N_534);
xnor U607 (N_607,N_557,N_441);
nand U608 (N_608,N_386,N_485);
and U609 (N_609,N_516,N_535);
nand U610 (N_610,N_418,In_891);
xor U611 (N_611,N_126,N_596);
xor U612 (N_612,In_984,N_539);
or U613 (N_613,N_463,N_501);
and U614 (N_614,N_301,N_300);
or U615 (N_615,N_344,N_357);
nor U616 (N_616,N_584,N_478);
and U617 (N_617,N_540,N_226);
nand U618 (N_618,In_552,N_345);
or U619 (N_619,N_305,In_133);
and U620 (N_620,In_786,In_716);
or U621 (N_621,N_403,In_692);
nor U622 (N_622,N_473,In_687);
or U623 (N_623,N_406,N_590);
nand U624 (N_624,N_459,N_443);
nor U625 (N_625,N_471,In_919);
nor U626 (N_626,N_258,N_537);
and U627 (N_627,In_33,N_435);
nand U628 (N_628,N_583,In_630);
nand U629 (N_629,N_581,N_521);
nor U630 (N_630,N_489,N_182);
xor U631 (N_631,N_328,N_432);
xor U632 (N_632,N_594,N_429);
or U633 (N_633,In_180,N_523);
or U634 (N_634,N_290,N_526);
nor U635 (N_635,N_51,N_3);
nand U636 (N_636,In_245,N_502);
xor U637 (N_637,N_447,N_311);
nand U638 (N_638,In_622,N_456);
and U639 (N_639,N_460,N_245);
and U640 (N_640,N_448,N_407);
and U641 (N_641,N_493,N_554);
nor U642 (N_642,N_514,N_519);
nand U643 (N_643,N_547,N_206);
or U644 (N_644,N_438,N_188);
nand U645 (N_645,N_453,N_474);
nor U646 (N_646,N_157,N_506);
xnor U647 (N_647,N_484,N_551);
nor U648 (N_648,N_262,In_619);
xnor U649 (N_649,N_597,In_87);
or U650 (N_650,N_472,N_417);
nand U651 (N_651,N_462,N_503);
nor U652 (N_652,In_0,N_582);
or U653 (N_653,N_282,N_401);
and U654 (N_654,N_513,N_571);
nand U655 (N_655,N_436,In_840);
xor U656 (N_656,N_545,N_358);
or U657 (N_657,N_444,In_189);
xor U658 (N_658,In_416,In_910);
nand U659 (N_659,N_580,N_598);
or U660 (N_660,In_457,N_445);
or U661 (N_661,N_550,N_576);
or U662 (N_662,N_201,N_546);
xor U663 (N_663,N_108,N_556);
xor U664 (N_664,N_455,In_6);
nor U665 (N_665,N_528,N_112);
xnor U666 (N_666,N_538,N_370);
xor U667 (N_667,In_956,N_520);
and U668 (N_668,N_352,N_354);
nand U669 (N_669,In_69,N_488);
and U670 (N_670,In_650,N_449);
nand U671 (N_671,N_423,N_364);
xor U672 (N_672,N_80,N_76);
or U673 (N_673,In_96,N_543);
xnor U674 (N_674,In_173,N_85);
nor U675 (N_675,N_588,N_265);
nand U676 (N_676,N_525,N_31);
or U677 (N_677,N_492,N_433);
and U678 (N_678,In_511,N_241);
xnor U679 (N_679,N_94,In_790);
nand U680 (N_680,N_338,In_60);
xnor U681 (N_681,N_412,N_200);
and U682 (N_682,In_979,N_118);
nand U683 (N_683,N_575,N_425);
nor U684 (N_684,N_276,N_309);
and U685 (N_685,In_961,N_465);
nand U686 (N_686,In_426,N_593);
nand U687 (N_687,N_428,N_411);
or U688 (N_688,N_422,N_424);
nor U689 (N_689,In_213,N_599);
nand U690 (N_690,N_98,N_275);
or U691 (N_691,N_161,N_589);
and U692 (N_692,N_482,N_585);
xnor U693 (N_693,N_413,In_468);
nand U694 (N_694,N_382,N_185);
and U695 (N_695,N_176,N_318);
xor U696 (N_696,N_59,In_208);
or U697 (N_697,N_434,N_511);
xnor U698 (N_698,N_350,In_992);
and U699 (N_699,N_587,N_255);
nand U700 (N_700,In_449,In_62);
xnor U701 (N_701,N_568,N_330);
or U702 (N_702,N_355,N_419);
and U703 (N_703,N_497,N_171);
nor U704 (N_704,In_154,In_998);
nand U705 (N_705,N_409,In_501);
and U706 (N_706,N_457,N_552);
nand U707 (N_707,N_481,N_378);
and U708 (N_708,In_564,N_490);
xor U709 (N_709,In_604,N_527);
xor U710 (N_710,In_764,N_561);
nor U711 (N_711,N_559,In_580);
nor U712 (N_712,N_592,In_596);
and U713 (N_713,N_437,N_106);
xor U714 (N_714,N_451,In_83);
nor U715 (N_715,N_553,N_66);
nor U716 (N_716,N_510,N_533);
and U717 (N_717,N_466,In_550);
nand U718 (N_718,N_452,In_184);
nor U719 (N_719,N_250,N_348);
and U720 (N_720,N_365,N_567);
or U721 (N_721,N_591,N_454);
nor U722 (N_722,N_500,In_952);
and U723 (N_723,N_496,N_555);
nand U724 (N_724,In_401,In_765);
nor U725 (N_725,N_498,N_294);
or U726 (N_726,In_892,N_446);
nand U727 (N_727,In_504,In_859);
xor U728 (N_728,In_708,N_532);
nand U729 (N_729,In_508,N_491);
and U730 (N_730,In_47,N_142);
or U731 (N_731,N_307,N_505);
xor U732 (N_732,In_220,In_825);
or U733 (N_733,N_518,N_461);
or U734 (N_734,N_548,N_379);
and U735 (N_735,N_586,In_845);
xor U736 (N_736,In_751,N_544);
or U737 (N_737,N_88,N_504);
or U738 (N_738,N_541,N_536);
and U739 (N_739,N_573,N_297);
nor U740 (N_740,N_464,N_475);
nor U741 (N_741,N_416,N_356);
nand U742 (N_742,In_928,N_507);
nand U743 (N_743,N_530,In_641);
nor U744 (N_744,N_574,N_9);
and U745 (N_745,N_400,N_329);
and U746 (N_746,N_439,N_549);
nor U747 (N_747,In_536,N_117);
and U748 (N_748,N_319,N_150);
xnor U749 (N_749,In_330,N_499);
and U750 (N_750,In_911,N_15);
and U751 (N_751,N_79,In_64);
xor U752 (N_752,In_292,N_468);
and U753 (N_753,N_274,N_111);
and U754 (N_754,In_242,In_698);
nor U755 (N_755,N_431,N_291);
xnor U756 (N_756,N_480,N_391);
and U757 (N_757,N_405,N_577);
or U758 (N_758,N_469,N_408);
and U759 (N_759,N_73,N_414);
nor U760 (N_760,N_558,N_420);
xnor U761 (N_761,N_415,N_404);
and U762 (N_762,N_375,N_205);
xor U763 (N_763,In_111,N_410);
nor U764 (N_764,N_517,N_570);
and U765 (N_765,N_531,In_445);
xnor U766 (N_766,In_724,N_40);
nand U767 (N_767,N_361,N_487);
or U768 (N_768,N_569,N_579);
xnor U769 (N_769,In_59,N_486);
xor U770 (N_770,N_371,In_238);
or U771 (N_771,In_964,N_467);
or U772 (N_772,N_104,N_279);
xnor U773 (N_773,N_293,N_476);
and U774 (N_774,N_268,N_529);
nor U775 (N_775,In_510,N_68);
or U776 (N_776,N_387,N_509);
or U777 (N_777,N_214,N_572);
nor U778 (N_778,N_470,N_458);
and U779 (N_779,In_482,N_522);
and U780 (N_780,N_566,In_169);
xor U781 (N_781,N_426,N_231);
nor U782 (N_782,In_971,N_479);
xor U783 (N_783,N_17,N_116);
or U784 (N_784,N_402,In_466);
and U785 (N_785,N_512,N_562);
and U786 (N_786,In_246,N_563);
nand U787 (N_787,N_442,In_67);
and U788 (N_788,N_230,In_931);
and U789 (N_789,In_886,In_895);
nor U790 (N_790,N_440,In_976);
and U791 (N_791,In_467,N_247);
nor U792 (N_792,In_21,N_331);
xor U793 (N_793,In_631,N_524);
nand U794 (N_794,N_578,N_477);
nor U795 (N_795,In_85,N_122);
or U796 (N_796,N_564,N_542);
or U797 (N_797,N_595,N_494);
nand U798 (N_798,In_750,In_291);
nand U799 (N_799,N_483,N_515);
nand U800 (N_800,N_796,N_696);
nand U801 (N_801,N_642,N_618);
xnor U802 (N_802,N_793,N_620);
or U803 (N_803,N_727,N_736);
xor U804 (N_804,N_776,N_629);
nand U805 (N_805,N_626,N_713);
nor U806 (N_806,N_765,N_783);
nor U807 (N_807,N_746,N_656);
xor U808 (N_808,N_678,N_681);
or U809 (N_809,N_634,N_700);
nand U810 (N_810,N_738,N_606);
or U811 (N_811,N_777,N_773);
nor U812 (N_812,N_770,N_680);
nor U813 (N_813,N_639,N_646);
and U814 (N_814,N_645,N_655);
xor U815 (N_815,N_616,N_692);
or U816 (N_816,N_797,N_754);
nand U817 (N_817,N_665,N_759);
or U818 (N_818,N_728,N_615);
or U819 (N_819,N_747,N_689);
xor U820 (N_820,N_701,N_602);
xnor U821 (N_821,N_752,N_660);
xor U822 (N_822,N_695,N_785);
nor U823 (N_823,N_674,N_624);
or U824 (N_824,N_791,N_702);
or U825 (N_825,N_654,N_679);
nor U826 (N_826,N_730,N_651);
or U827 (N_827,N_698,N_610);
nor U828 (N_828,N_650,N_794);
or U829 (N_829,N_627,N_719);
nand U830 (N_830,N_649,N_737);
nand U831 (N_831,N_710,N_672);
nand U832 (N_832,N_760,N_677);
nand U833 (N_833,N_758,N_611);
xnor U834 (N_834,N_789,N_771);
nor U835 (N_835,N_687,N_751);
xor U836 (N_836,N_653,N_613);
nor U837 (N_837,N_722,N_670);
xnor U838 (N_838,N_742,N_724);
or U839 (N_839,N_731,N_675);
and U840 (N_840,N_658,N_682);
and U841 (N_841,N_647,N_782);
nor U842 (N_842,N_690,N_799);
nand U843 (N_843,N_635,N_694);
xnor U844 (N_844,N_683,N_663);
or U845 (N_845,N_693,N_664);
or U846 (N_846,N_715,N_600);
nor U847 (N_847,N_684,N_720);
or U848 (N_848,N_644,N_784);
and U849 (N_849,N_621,N_774);
nor U850 (N_850,N_711,N_735);
nor U851 (N_851,N_723,N_623);
nor U852 (N_852,N_762,N_767);
nand U853 (N_853,N_659,N_601);
nor U854 (N_854,N_709,N_703);
xor U855 (N_855,N_733,N_732);
xnor U856 (N_856,N_778,N_657);
xnor U857 (N_857,N_764,N_637);
or U858 (N_858,N_640,N_798);
xnor U859 (N_859,N_603,N_755);
nor U860 (N_860,N_761,N_638);
and U861 (N_861,N_666,N_707);
xor U862 (N_862,N_795,N_775);
xnor U863 (N_863,N_788,N_792);
nor U864 (N_864,N_704,N_617);
and U865 (N_865,N_779,N_766);
nor U866 (N_866,N_780,N_673);
nor U867 (N_867,N_741,N_706);
or U868 (N_868,N_628,N_745);
and U869 (N_869,N_632,N_609);
and U870 (N_870,N_787,N_671);
and U871 (N_871,N_641,N_622);
or U872 (N_872,N_748,N_753);
nand U873 (N_873,N_749,N_721);
nor U874 (N_874,N_740,N_712);
xnor U875 (N_875,N_608,N_750);
or U876 (N_876,N_790,N_676);
nand U877 (N_877,N_686,N_708);
or U878 (N_878,N_772,N_763);
xnor U879 (N_879,N_688,N_605);
xor U880 (N_880,N_662,N_786);
xor U881 (N_881,N_614,N_743);
nand U882 (N_882,N_697,N_734);
nor U883 (N_883,N_648,N_685);
xnor U884 (N_884,N_631,N_725);
and U885 (N_885,N_669,N_636);
nor U886 (N_886,N_652,N_612);
or U887 (N_887,N_726,N_729);
or U888 (N_888,N_604,N_630);
xnor U889 (N_889,N_667,N_739);
or U890 (N_890,N_607,N_699);
xor U891 (N_891,N_691,N_744);
nand U892 (N_892,N_781,N_716);
or U893 (N_893,N_714,N_643);
nand U894 (N_894,N_668,N_769);
and U895 (N_895,N_705,N_718);
xnor U896 (N_896,N_661,N_625);
nand U897 (N_897,N_768,N_757);
and U898 (N_898,N_717,N_619);
nand U899 (N_899,N_756,N_633);
and U900 (N_900,N_708,N_754);
or U901 (N_901,N_623,N_711);
or U902 (N_902,N_793,N_734);
or U903 (N_903,N_742,N_790);
nor U904 (N_904,N_765,N_798);
and U905 (N_905,N_752,N_665);
and U906 (N_906,N_631,N_720);
nand U907 (N_907,N_624,N_761);
or U908 (N_908,N_752,N_647);
xor U909 (N_909,N_633,N_687);
xnor U910 (N_910,N_630,N_610);
and U911 (N_911,N_796,N_693);
nand U912 (N_912,N_712,N_617);
and U913 (N_913,N_664,N_673);
nor U914 (N_914,N_617,N_764);
nand U915 (N_915,N_631,N_751);
nand U916 (N_916,N_700,N_641);
xnor U917 (N_917,N_654,N_622);
and U918 (N_918,N_672,N_636);
and U919 (N_919,N_799,N_730);
nand U920 (N_920,N_777,N_658);
nor U921 (N_921,N_717,N_728);
and U922 (N_922,N_636,N_660);
nor U923 (N_923,N_666,N_713);
and U924 (N_924,N_646,N_659);
and U925 (N_925,N_780,N_789);
nand U926 (N_926,N_684,N_724);
xnor U927 (N_927,N_746,N_707);
xnor U928 (N_928,N_621,N_739);
xnor U929 (N_929,N_737,N_714);
xnor U930 (N_930,N_618,N_615);
nor U931 (N_931,N_746,N_723);
nand U932 (N_932,N_759,N_669);
and U933 (N_933,N_777,N_619);
xor U934 (N_934,N_603,N_720);
nor U935 (N_935,N_729,N_609);
and U936 (N_936,N_684,N_782);
nand U937 (N_937,N_664,N_731);
xnor U938 (N_938,N_728,N_665);
nor U939 (N_939,N_689,N_678);
nor U940 (N_940,N_676,N_795);
nor U941 (N_941,N_651,N_758);
and U942 (N_942,N_772,N_620);
or U943 (N_943,N_683,N_679);
or U944 (N_944,N_746,N_660);
or U945 (N_945,N_737,N_666);
nor U946 (N_946,N_738,N_672);
xnor U947 (N_947,N_714,N_652);
xor U948 (N_948,N_774,N_695);
and U949 (N_949,N_709,N_619);
nor U950 (N_950,N_682,N_713);
xor U951 (N_951,N_655,N_769);
nor U952 (N_952,N_734,N_782);
or U953 (N_953,N_763,N_707);
and U954 (N_954,N_645,N_755);
nand U955 (N_955,N_775,N_747);
xor U956 (N_956,N_681,N_689);
xnor U957 (N_957,N_726,N_747);
nand U958 (N_958,N_761,N_652);
nor U959 (N_959,N_627,N_708);
and U960 (N_960,N_754,N_735);
xnor U961 (N_961,N_784,N_785);
nor U962 (N_962,N_672,N_775);
nor U963 (N_963,N_782,N_609);
nor U964 (N_964,N_634,N_655);
and U965 (N_965,N_739,N_736);
and U966 (N_966,N_613,N_681);
nor U967 (N_967,N_756,N_688);
or U968 (N_968,N_687,N_644);
or U969 (N_969,N_640,N_737);
xor U970 (N_970,N_612,N_798);
or U971 (N_971,N_683,N_675);
nand U972 (N_972,N_669,N_719);
nand U973 (N_973,N_703,N_751);
nand U974 (N_974,N_681,N_727);
nor U975 (N_975,N_630,N_759);
nor U976 (N_976,N_681,N_710);
or U977 (N_977,N_680,N_709);
and U978 (N_978,N_679,N_697);
and U979 (N_979,N_795,N_616);
xnor U980 (N_980,N_615,N_634);
xnor U981 (N_981,N_792,N_631);
nor U982 (N_982,N_752,N_683);
nand U983 (N_983,N_600,N_722);
xor U984 (N_984,N_774,N_652);
or U985 (N_985,N_764,N_739);
xnor U986 (N_986,N_666,N_797);
xnor U987 (N_987,N_657,N_764);
xor U988 (N_988,N_674,N_615);
nand U989 (N_989,N_754,N_669);
or U990 (N_990,N_614,N_666);
nand U991 (N_991,N_684,N_737);
nor U992 (N_992,N_753,N_683);
or U993 (N_993,N_711,N_792);
xor U994 (N_994,N_674,N_699);
nand U995 (N_995,N_666,N_743);
xnor U996 (N_996,N_662,N_711);
and U997 (N_997,N_727,N_737);
nor U998 (N_998,N_791,N_680);
or U999 (N_999,N_653,N_753);
and U1000 (N_1000,N_920,N_970);
nor U1001 (N_1001,N_855,N_984);
xor U1002 (N_1002,N_801,N_832);
xor U1003 (N_1003,N_858,N_968);
xor U1004 (N_1004,N_999,N_802);
nand U1005 (N_1005,N_965,N_837);
nor U1006 (N_1006,N_844,N_897);
xnor U1007 (N_1007,N_865,N_946);
and U1008 (N_1008,N_845,N_963);
or U1009 (N_1009,N_941,N_905);
nand U1010 (N_1010,N_969,N_835);
nor U1011 (N_1011,N_871,N_981);
xor U1012 (N_1012,N_888,N_924);
xor U1013 (N_1013,N_904,N_867);
or U1014 (N_1014,N_995,N_883);
or U1015 (N_1015,N_959,N_836);
and U1016 (N_1016,N_948,N_913);
or U1017 (N_1017,N_919,N_964);
nand U1018 (N_1018,N_917,N_911);
nor U1019 (N_1019,N_975,N_820);
xor U1020 (N_1020,N_928,N_908);
nor U1021 (N_1021,N_866,N_982);
nand U1022 (N_1022,N_822,N_932);
or U1023 (N_1023,N_921,N_955);
nor U1024 (N_1024,N_848,N_891);
and U1025 (N_1025,N_890,N_900);
xnor U1026 (N_1026,N_872,N_885);
and U1027 (N_1027,N_952,N_925);
or U1028 (N_1028,N_990,N_958);
nor U1029 (N_1029,N_869,N_956);
and U1030 (N_1030,N_831,N_876);
or U1031 (N_1031,N_825,N_863);
and U1032 (N_1032,N_812,N_962);
nor U1033 (N_1033,N_988,N_824);
and U1034 (N_1034,N_915,N_852);
and U1035 (N_1035,N_854,N_814);
or U1036 (N_1036,N_980,N_934);
and U1037 (N_1037,N_927,N_808);
or U1038 (N_1038,N_971,N_838);
nor U1039 (N_1039,N_972,N_849);
or U1040 (N_1040,N_819,N_877);
and U1041 (N_1041,N_873,N_994);
xor U1042 (N_1042,N_910,N_935);
or U1043 (N_1043,N_823,N_987);
xor U1044 (N_1044,N_940,N_813);
nor U1045 (N_1045,N_985,N_875);
or U1046 (N_1046,N_878,N_998);
nor U1047 (N_1047,N_951,N_944);
nor U1048 (N_1048,N_827,N_979);
xor U1049 (N_1049,N_986,N_974);
nand U1050 (N_1050,N_939,N_926);
or U1051 (N_1051,N_887,N_899);
xnor U1052 (N_1052,N_997,N_991);
nor U1053 (N_1053,N_879,N_803);
or U1054 (N_1054,N_950,N_978);
xor U1055 (N_1055,N_923,N_886);
and U1056 (N_1056,N_936,N_850);
or U1057 (N_1057,N_843,N_842);
and U1058 (N_1058,N_804,N_902);
nor U1059 (N_1059,N_945,N_929);
and U1060 (N_1060,N_816,N_943);
or U1061 (N_1061,N_806,N_947);
and U1062 (N_1062,N_909,N_821);
nor U1063 (N_1063,N_807,N_861);
nand U1064 (N_1064,N_967,N_853);
xnor U1065 (N_1065,N_993,N_893);
nand U1066 (N_1066,N_884,N_903);
xnor U1067 (N_1067,N_957,N_846);
or U1068 (N_1068,N_907,N_914);
nor U1069 (N_1069,N_906,N_847);
nand U1070 (N_1070,N_800,N_942);
and U1071 (N_1071,N_868,N_809);
nand U1072 (N_1072,N_839,N_930);
nand U1073 (N_1073,N_996,N_901);
and U1074 (N_1074,N_834,N_817);
nand U1075 (N_1075,N_895,N_864);
nor U1076 (N_1076,N_961,N_857);
nand U1077 (N_1077,N_840,N_892);
or U1078 (N_1078,N_815,N_973);
xnor U1079 (N_1079,N_851,N_938);
nand U1080 (N_1080,N_881,N_860);
or U1081 (N_1081,N_870,N_859);
nand U1082 (N_1082,N_931,N_874);
nand U1083 (N_1083,N_922,N_810);
and U1084 (N_1084,N_805,N_889);
nand U1085 (N_1085,N_966,N_830);
nor U1086 (N_1086,N_916,N_953);
xnor U1087 (N_1087,N_826,N_977);
nand U1088 (N_1088,N_949,N_862);
xnor U1089 (N_1089,N_918,N_882);
nor U1090 (N_1090,N_818,N_937);
or U1091 (N_1091,N_829,N_912);
nor U1092 (N_1092,N_828,N_833);
nand U1093 (N_1093,N_960,N_983);
and U1094 (N_1094,N_992,N_933);
or U1095 (N_1095,N_880,N_976);
nor U1096 (N_1096,N_989,N_898);
and U1097 (N_1097,N_841,N_811);
xnor U1098 (N_1098,N_896,N_894);
and U1099 (N_1099,N_954,N_856);
or U1100 (N_1100,N_808,N_943);
nand U1101 (N_1101,N_998,N_891);
nand U1102 (N_1102,N_910,N_992);
and U1103 (N_1103,N_913,N_910);
nand U1104 (N_1104,N_930,N_948);
xnor U1105 (N_1105,N_990,N_997);
xnor U1106 (N_1106,N_961,N_948);
nand U1107 (N_1107,N_893,N_964);
or U1108 (N_1108,N_864,N_851);
nand U1109 (N_1109,N_965,N_904);
xor U1110 (N_1110,N_995,N_996);
and U1111 (N_1111,N_938,N_951);
nand U1112 (N_1112,N_865,N_935);
or U1113 (N_1113,N_980,N_847);
and U1114 (N_1114,N_922,N_809);
or U1115 (N_1115,N_879,N_807);
nand U1116 (N_1116,N_950,N_849);
nand U1117 (N_1117,N_883,N_920);
and U1118 (N_1118,N_935,N_955);
xor U1119 (N_1119,N_933,N_990);
and U1120 (N_1120,N_902,N_888);
xor U1121 (N_1121,N_960,N_882);
nand U1122 (N_1122,N_891,N_832);
xnor U1123 (N_1123,N_801,N_841);
xor U1124 (N_1124,N_888,N_932);
and U1125 (N_1125,N_986,N_913);
xor U1126 (N_1126,N_820,N_962);
and U1127 (N_1127,N_941,N_979);
nand U1128 (N_1128,N_924,N_825);
xor U1129 (N_1129,N_890,N_866);
xor U1130 (N_1130,N_971,N_857);
xor U1131 (N_1131,N_805,N_853);
nor U1132 (N_1132,N_852,N_838);
nor U1133 (N_1133,N_806,N_800);
and U1134 (N_1134,N_845,N_811);
xnor U1135 (N_1135,N_864,N_848);
nand U1136 (N_1136,N_813,N_992);
and U1137 (N_1137,N_949,N_986);
nor U1138 (N_1138,N_953,N_931);
and U1139 (N_1139,N_909,N_973);
nor U1140 (N_1140,N_881,N_890);
nor U1141 (N_1141,N_862,N_910);
nand U1142 (N_1142,N_917,N_894);
xor U1143 (N_1143,N_925,N_969);
xnor U1144 (N_1144,N_950,N_904);
xor U1145 (N_1145,N_992,N_999);
xor U1146 (N_1146,N_822,N_800);
nand U1147 (N_1147,N_922,N_840);
nor U1148 (N_1148,N_962,N_903);
xnor U1149 (N_1149,N_802,N_941);
nor U1150 (N_1150,N_888,N_844);
and U1151 (N_1151,N_945,N_859);
nand U1152 (N_1152,N_896,N_816);
xor U1153 (N_1153,N_825,N_985);
or U1154 (N_1154,N_927,N_870);
nand U1155 (N_1155,N_833,N_988);
nor U1156 (N_1156,N_867,N_839);
xnor U1157 (N_1157,N_971,N_827);
nor U1158 (N_1158,N_952,N_862);
or U1159 (N_1159,N_820,N_879);
and U1160 (N_1160,N_952,N_877);
xor U1161 (N_1161,N_881,N_812);
or U1162 (N_1162,N_989,N_856);
and U1163 (N_1163,N_969,N_967);
nand U1164 (N_1164,N_873,N_878);
xnor U1165 (N_1165,N_973,N_935);
or U1166 (N_1166,N_882,N_964);
or U1167 (N_1167,N_871,N_812);
nand U1168 (N_1168,N_803,N_949);
nor U1169 (N_1169,N_937,N_875);
nand U1170 (N_1170,N_964,N_968);
or U1171 (N_1171,N_866,N_976);
and U1172 (N_1172,N_906,N_953);
and U1173 (N_1173,N_954,N_922);
or U1174 (N_1174,N_999,N_941);
nor U1175 (N_1175,N_846,N_834);
or U1176 (N_1176,N_940,N_883);
and U1177 (N_1177,N_947,N_831);
xor U1178 (N_1178,N_990,N_971);
nor U1179 (N_1179,N_961,N_992);
nand U1180 (N_1180,N_912,N_827);
or U1181 (N_1181,N_845,N_892);
nor U1182 (N_1182,N_853,N_864);
or U1183 (N_1183,N_968,N_819);
nand U1184 (N_1184,N_835,N_854);
and U1185 (N_1185,N_871,N_876);
nand U1186 (N_1186,N_891,N_925);
xor U1187 (N_1187,N_853,N_931);
xnor U1188 (N_1188,N_989,N_817);
or U1189 (N_1189,N_926,N_925);
nor U1190 (N_1190,N_883,N_951);
nor U1191 (N_1191,N_806,N_959);
nor U1192 (N_1192,N_940,N_822);
nand U1193 (N_1193,N_953,N_993);
or U1194 (N_1194,N_888,N_941);
or U1195 (N_1195,N_862,N_876);
or U1196 (N_1196,N_906,N_891);
nand U1197 (N_1197,N_813,N_920);
and U1198 (N_1198,N_918,N_824);
nand U1199 (N_1199,N_815,N_996);
nand U1200 (N_1200,N_1092,N_1068);
nor U1201 (N_1201,N_1036,N_1009);
xnor U1202 (N_1202,N_1028,N_1001);
and U1203 (N_1203,N_1152,N_1109);
nor U1204 (N_1204,N_1065,N_1054);
xnor U1205 (N_1205,N_1189,N_1084);
nor U1206 (N_1206,N_1062,N_1097);
nand U1207 (N_1207,N_1067,N_1014);
and U1208 (N_1208,N_1002,N_1116);
xnor U1209 (N_1209,N_1031,N_1126);
nand U1210 (N_1210,N_1087,N_1190);
nor U1211 (N_1211,N_1158,N_1023);
nand U1212 (N_1212,N_1156,N_1198);
nand U1213 (N_1213,N_1008,N_1111);
nand U1214 (N_1214,N_1091,N_1179);
nor U1215 (N_1215,N_1021,N_1010);
nor U1216 (N_1216,N_1141,N_1027);
or U1217 (N_1217,N_1080,N_1165);
xnor U1218 (N_1218,N_1180,N_1032);
and U1219 (N_1219,N_1185,N_1045);
or U1220 (N_1220,N_1105,N_1187);
and U1221 (N_1221,N_1000,N_1121);
nor U1222 (N_1222,N_1071,N_1130);
and U1223 (N_1223,N_1137,N_1094);
and U1224 (N_1224,N_1132,N_1012);
xor U1225 (N_1225,N_1154,N_1188);
and U1226 (N_1226,N_1175,N_1022);
nor U1227 (N_1227,N_1128,N_1142);
xnor U1228 (N_1228,N_1192,N_1069);
nor U1229 (N_1229,N_1170,N_1043);
and U1230 (N_1230,N_1020,N_1129);
xor U1231 (N_1231,N_1114,N_1144);
or U1232 (N_1232,N_1193,N_1178);
and U1233 (N_1233,N_1146,N_1090);
or U1234 (N_1234,N_1153,N_1186);
nand U1235 (N_1235,N_1167,N_1024);
xnor U1236 (N_1236,N_1052,N_1136);
and U1237 (N_1237,N_1115,N_1074);
and U1238 (N_1238,N_1082,N_1118);
xnor U1239 (N_1239,N_1174,N_1095);
nand U1240 (N_1240,N_1149,N_1195);
and U1241 (N_1241,N_1127,N_1063);
nand U1242 (N_1242,N_1075,N_1124);
xnor U1243 (N_1243,N_1183,N_1182);
nor U1244 (N_1244,N_1176,N_1072);
xnor U1245 (N_1245,N_1162,N_1138);
nand U1246 (N_1246,N_1026,N_1085);
nor U1247 (N_1247,N_1135,N_1064);
xor U1248 (N_1248,N_1005,N_1061);
nor U1249 (N_1249,N_1139,N_1046);
and U1250 (N_1250,N_1169,N_1004);
nor U1251 (N_1251,N_1047,N_1060);
and U1252 (N_1252,N_1044,N_1112);
xnor U1253 (N_1253,N_1081,N_1196);
nand U1254 (N_1254,N_1058,N_1059);
or U1255 (N_1255,N_1113,N_1101);
and U1256 (N_1256,N_1089,N_1157);
nor U1257 (N_1257,N_1155,N_1018);
and U1258 (N_1258,N_1108,N_1177);
and U1259 (N_1259,N_1103,N_1029);
nor U1260 (N_1260,N_1166,N_1140);
nor U1261 (N_1261,N_1025,N_1122);
and U1262 (N_1262,N_1197,N_1070);
nand U1263 (N_1263,N_1053,N_1051);
and U1264 (N_1264,N_1151,N_1133);
nor U1265 (N_1265,N_1199,N_1040);
nand U1266 (N_1266,N_1038,N_1119);
xor U1267 (N_1267,N_1033,N_1019);
nor U1268 (N_1268,N_1098,N_1168);
xnor U1269 (N_1269,N_1184,N_1055);
and U1270 (N_1270,N_1078,N_1161);
nor U1271 (N_1271,N_1035,N_1134);
nand U1272 (N_1272,N_1076,N_1145);
and U1273 (N_1273,N_1037,N_1099);
nand U1274 (N_1274,N_1030,N_1171);
nor U1275 (N_1275,N_1007,N_1096);
and U1276 (N_1276,N_1120,N_1006);
nor U1277 (N_1277,N_1057,N_1049);
or U1278 (N_1278,N_1106,N_1104);
and U1279 (N_1279,N_1147,N_1150);
nand U1280 (N_1280,N_1034,N_1086);
or U1281 (N_1281,N_1110,N_1048);
and U1282 (N_1282,N_1011,N_1163);
xnor U1283 (N_1283,N_1159,N_1191);
and U1284 (N_1284,N_1056,N_1143);
and U1285 (N_1285,N_1173,N_1100);
xor U1286 (N_1286,N_1102,N_1160);
or U1287 (N_1287,N_1042,N_1107);
or U1288 (N_1288,N_1117,N_1079);
nand U1289 (N_1289,N_1181,N_1066);
and U1290 (N_1290,N_1013,N_1088);
and U1291 (N_1291,N_1077,N_1041);
and U1292 (N_1292,N_1194,N_1050);
and U1293 (N_1293,N_1073,N_1015);
or U1294 (N_1294,N_1172,N_1164);
xor U1295 (N_1295,N_1017,N_1148);
nor U1296 (N_1296,N_1131,N_1093);
nor U1297 (N_1297,N_1125,N_1039);
nor U1298 (N_1298,N_1016,N_1123);
nand U1299 (N_1299,N_1003,N_1083);
nor U1300 (N_1300,N_1187,N_1035);
and U1301 (N_1301,N_1082,N_1043);
xor U1302 (N_1302,N_1143,N_1066);
and U1303 (N_1303,N_1052,N_1022);
and U1304 (N_1304,N_1114,N_1087);
nor U1305 (N_1305,N_1031,N_1079);
or U1306 (N_1306,N_1077,N_1110);
nand U1307 (N_1307,N_1017,N_1184);
or U1308 (N_1308,N_1078,N_1076);
or U1309 (N_1309,N_1102,N_1043);
and U1310 (N_1310,N_1082,N_1162);
or U1311 (N_1311,N_1038,N_1157);
nor U1312 (N_1312,N_1145,N_1064);
nand U1313 (N_1313,N_1100,N_1143);
and U1314 (N_1314,N_1193,N_1157);
and U1315 (N_1315,N_1064,N_1125);
nand U1316 (N_1316,N_1162,N_1129);
and U1317 (N_1317,N_1090,N_1167);
nand U1318 (N_1318,N_1194,N_1064);
nor U1319 (N_1319,N_1184,N_1114);
or U1320 (N_1320,N_1079,N_1148);
nor U1321 (N_1321,N_1187,N_1018);
nand U1322 (N_1322,N_1054,N_1012);
or U1323 (N_1323,N_1167,N_1037);
nand U1324 (N_1324,N_1011,N_1167);
or U1325 (N_1325,N_1036,N_1038);
and U1326 (N_1326,N_1131,N_1118);
nor U1327 (N_1327,N_1066,N_1030);
nand U1328 (N_1328,N_1023,N_1071);
and U1329 (N_1329,N_1074,N_1139);
nor U1330 (N_1330,N_1161,N_1151);
or U1331 (N_1331,N_1016,N_1060);
and U1332 (N_1332,N_1096,N_1038);
or U1333 (N_1333,N_1094,N_1190);
and U1334 (N_1334,N_1151,N_1182);
xnor U1335 (N_1335,N_1089,N_1036);
xor U1336 (N_1336,N_1118,N_1013);
xnor U1337 (N_1337,N_1092,N_1102);
xor U1338 (N_1338,N_1086,N_1043);
nand U1339 (N_1339,N_1177,N_1039);
nand U1340 (N_1340,N_1176,N_1175);
xnor U1341 (N_1341,N_1060,N_1069);
nand U1342 (N_1342,N_1127,N_1166);
and U1343 (N_1343,N_1173,N_1142);
or U1344 (N_1344,N_1050,N_1103);
xor U1345 (N_1345,N_1148,N_1143);
and U1346 (N_1346,N_1100,N_1164);
or U1347 (N_1347,N_1126,N_1077);
or U1348 (N_1348,N_1041,N_1171);
or U1349 (N_1349,N_1148,N_1150);
nor U1350 (N_1350,N_1015,N_1138);
nand U1351 (N_1351,N_1124,N_1039);
or U1352 (N_1352,N_1145,N_1053);
and U1353 (N_1353,N_1062,N_1050);
xor U1354 (N_1354,N_1189,N_1190);
nor U1355 (N_1355,N_1127,N_1146);
or U1356 (N_1356,N_1048,N_1159);
and U1357 (N_1357,N_1147,N_1182);
and U1358 (N_1358,N_1158,N_1033);
xor U1359 (N_1359,N_1165,N_1040);
and U1360 (N_1360,N_1191,N_1154);
and U1361 (N_1361,N_1045,N_1119);
nor U1362 (N_1362,N_1104,N_1167);
nor U1363 (N_1363,N_1191,N_1199);
or U1364 (N_1364,N_1041,N_1187);
xnor U1365 (N_1365,N_1181,N_1003);
nor U1366 (N_1366,N_1027,N_1189);
or U1367 (N_1367,N_1151,N_1026);
nand U1368 (N_1368,N_1010,N_1092);
or U1369 (N_1369,N_1026,N_1119);
and U1370 (N_1370,N_1031,N_1010);
xor U1371 (N_1371,N_1147,N_1157);
xor U1372 (N_1372,N_1046,N_1140);
or U1373 (N_1373,N_1012,N_1089);
xor U1374 (N_1374,N_1034,N_1089);
or U1375 (N_1375,N_1044,N_1055);
xor U1376 (N_1376,N_1080,N_1101);
nand U1377 (N_1377,N_1122,N_1125);
nor U1378 (N_1378,N_1122,N_1102);
and U1379 (N_1379,N_1021,N_1138);
nand U1380 (N_1380,N_1155,N_1151);
and U1381 (N_1381,N_1007,N_1017);
nand U1382 (N_1382,N_1159,N_1139);
or U1383 (N_1383,N_1151,N_1199);
or U1384 (N_1384,N_1168,N_1018);
or U1385 (N_1385,N_1181,N_1138);
xnor U1386 (N_1386,N_1034,N_1194);
and U1387 (N_1387,N_1004,N_1154);
nor U1388 (N_1388,N_1102,N_1180);
nor U1389 (N_1389,N_1173,N_1068);
or U1390 (N_1390,N_1112,N_1182);
and U1391 (N_1391,N_1120,N_1025);
and U1392 (N_1392,N_1135,N_1001);
xnor U1393 (N_1393,N_1092,N_1126);
or U1394 (N_1394,N_1087,N_1188);
or U1395 (N_1395,N_1198,N_1024);
nand U1396 (N_1396,N_1140,N_1053);
nor U1397 (N_1397,N_1174,N_1121);
xnor U1398 (N_1398,N_1086,N_1031);
and U1399 (N_1399,N_1010,N_1192);
nand U1400 (N_1400,N_1325,N_1230);
and U1401 (N_1401,N_1290,N_1350);
nand U1402 (N_1402,N_1251,N_1388);
nor U1403 (N_1403,N_1320,N_1259);
and U1404 (N_1404,N_1305,N_1393);
nand U1405 (N_1405,N_1318,N_1294);
and U1406 (N_1406,N_1313,N_1367);
or U1407 (N_1407,N_1341,N_1256);
nand U1408 (N_1408,N_1205,N_1346);
nand U1409 (N_1409,N_1277,N_1287);
nor U1410 (N_1410,N_1208,N_1394);
or U1411 (N_1411,N_1239,N_1337);
or U1412 (N_1412,N_1399,N_1348);
and U1413 (N_1413,N_1371,N_1324);
and U1414 (N_1414,N_1391,N_1232);
nand U1415 (N_1415,N_1303,N_1296);
nor U1416 (N_1416,N_1357,N_1266);
and U1417 (N_1417,N_1240,N_1356);
nand U1418 (N_1418,N_1212,N_1340);
nor U1419 (N_1419,N_1336,N_1210);
or U1420 (N_1420,N_1322,N_1223);
nand U1421 (N_1421,N_1274,N_1258);
and U1422 (N_1422,N_1219,N_1269);
and U1423 (N_1423,N_1321,N_1301);
or U1424 (N_1424,N_1334,N_1363);
xor U1425 (N_1425,N_1300,N_1309);
xnor U1426 (N_1426,N_1200,N_1222);
xor U1427 (N_1427,N_1271,N_1331);
nand U1428 (N_1428,N_1280,N_1272);
nand U1429 (N_1429,N_1355,N_1338);
xnor U1430 (N_1430,N_1374,N_1328);
nand U1431 (N_1431,N_1304,N_1268);
or U1432 (N_1432,N_1329,N_1255);
and U1433 (N_1433,N_1207,N_1261);
and U1434 (N_1434,N_1395,N_1265);
xnor U1435 (N_1435,N_1242,N_1323);
xnor U1436 (N_1436,N_1270,N_1264);
nand U1437 (N_1437,N_1358,N_1282);
or U1438 (N_1438,N_1228,N_1335);
xnor U1439 (N_1439,N_1216,N_1227);
xnor U1440 (N_1440,N_1342,N_1368);
xor U1441 (N_1441,N_1248,N_1306);
xor U1442 (N_1442,N_1299,N_1387);
nand U1443 (N_1443,N_1352,N_1224);
xnor U1444 (N_1444,N_1285,N_1312);
and U1445 (N_1445,N_1246,N_1382);
or U1446 (N_1446,N_1234,N_1267);
and U1447 (N_1447,N_1247,N_1273);
xor U1448 (N_1448,N_1260,N_1288);
xor U1449 (N_1449,N_1345,N_1370);
or U1450 (N_1450,N_1377,N_1381);
nand U1451 (N_1451,N_1279,N_1241);
xor U1452 (N_1452,N_1353,N_1218);
nor U1453 (N_1453,N_1364,N_1202);
and U1454 (N_1454,N_1281,N_1362);
and U1455 (N_1455,N_1384,N_1385);
nor U1456 (N_1456,N_1347,N_1220);
or U1457 (N_1457,N_1201,N_1284);
nand U1458 (N_1458,N_1263,N_1369);
and U1459 (N_1459,N_1398,N_1302);
nand U1460 (N_1460,N_1235,N_1226);
and U1461 (N_1461,N_1225,N_1209);
or U1462 (N_1462,N_1389,N_1317);
nor U1463 (N_1463,N_1311,N_1339);
nor U1464 (N_1464,N_1307,N_1376);
or U1465 (N_1465,N_1236,N_1206);
or U1466 (N_1466,N_1278,N_1229);
or U1467 (N_1467,N_1237,N_1344);
nand U1468 (N_1468,N_1310,N_1383);
xor U1469 (N_1469,N_1379,N_1254);
or U1470 (N_1470,N_1349,N_1250);
nand U1471 (N_1471,N_1286,N_1308);
xor U1472 (N_1472,N_1330,N_1380);
or U1473 (N_1473,N_1365,N_1392);
nand U1474 (N_1474,N_1327,N_1244);
and U1475 (N_1475,N_1291,N_1275);
nand U1476 (N_1476,N_1332,N_1249);
and U1477 (N_1477,N_1295,N_1204);
and U1478 (N_1478,N_1298,N_1211);
and U1479 (N_1479,N_1289,N_1354);
or U1480 (N_1480,N_1361,N_1319);
xnor U1481 (N_1481,N_1283,N_1253);
nand U1482 (N_1482,N_1297,N_1360);
or U1483 (N_1483,N_1351,N_1215);
xor U1484 (N_1484,N_1213,N_1397);
nor U1485 (N_1485,N_1390,N_1372);
or U1486 (N_1486,N_1252,N_1333);
nor U1487 (N_1487,N_1262,N_1276);
or U1488 (N_1488,N_1378,N_1221);
nor U1489 (N_1489,N_1243,N_1326);
nand U1490 (N_1490,N_1316,N_1373);
or U1491 (N_1491,N_1375,N_1343);
xor U1492 (N_1492,N_1359,N_1233);
or U1493 (N_1493,N_1231,N_1214);
nand U1494 (N_1494,N_1245,N_1217);
and U1495 (N_1495,N_1386,N_1396);
xor U1496 (N_1496,N_1314,N_1292);
nor U1497 (N_1497,N_1203,N_1315);
nand U1498 (N_1498,N_1238,N_1293);
and U1499 (N_1499,N_1366,N_1257);
nor U1500 (N_1500,N_1248,N_1351);
and U1501 (N_1501,N_1310,N_1367);
nor U1502 (N_1502,N_1209,N_1328);
and U1503 (N_1503,N_1234,N_1211);
nor U1504 (N_1504,N_1392,N_1344);
xnor U1505 (N_1505,N_1320,N_1308);
xnor U1506 (N_1506,N_1339,N_1351);
xor U1507 (N_1507,N_1310,N_1258);
nor U1508 (N_1508,N_1216,N_1303);
or U1509 (N_1509,N_1216,N_1284);
nor U1510 (N_1510,N_1254,N_1326);
and U1511 (N_1511,N_1256,N_1233);
or U1512 (N_1512,N_1259,N_1366);
and U1513 (N_1513,N_1388,N_1398);
or U1514 (N_1514,N_1234,N_1246);
xnor U1515 (N_1515,N_1272,N_1238);
xnor U1516 (N_1516,N_1293,N_1246);
and U1517 (N_1517,N_1372,N_1358);
or U1518 (N_1518,N_1345,N_1349);
and U1519 (N_1519,N_1280,N_1373);
or U1520 (N_1520,N_1370,N_1273);
nor U1521 (N_1521,N_1227,N_1287);
and U1522 (N_1522,N_1358,N_1348);
nor U1523 (N_1523,N_1375,N_1320);
and U1524 (N_1524,N_1319,N_1344);
nand U1525 (N_1525,N_1259,N_1327);
nand U1526 (N_1526,N_1330,N_1222);
xor U1527 (N_1527,N_1326,N_1322);
xnor U1528 (N_1528,N_1204,N_1291);
and U1529 (N_1529,N_1397,N_1214);
nor U1530 (N_1530,N_1210,N_1236);
and U1531 (N_1531,N_1225,N_1342);
nor U1532 (N_1532,N_1304,N_1388);
nand U1533 (N_1533,N_1347,N_1278);
nand U1534 (N_1534,N_1230,N_1270);
xnor U1535 (N_1535,N_1256,N_1258);
and U1536 (N_1536,N_1279,N_1320);
or U1537 (N_1537,N_1214,N_1322);
and U1538 (N_1538,N_1235,N_1282);
nor U1539 (N_1539,N_1215,N_1231);
xnor U1540 (N_1540,N_1392,N_1233);
nor U1541 (N_1541,N_1294,N_1286);
or U1542 (N_1542,N_1274,N_1327);
or U1543 (N_1543,N_1325,N_1378);
nor U1544 (N_1544,N_1345,N_1273);
or U1545 (N_1545,N_1390,N_1304);
nand U1546 (N_1546,N_1222,N_1225);
and U1547 (N_1547,N_1339,N_1380);
or U1548 (N_1548,N_1363,N_1279);
and U1549 (N_1549,N_1252,N_1211);
xnor U1550 (N_1550,N_1252,N_1229);
and U1551 (N_1551,N_1348,N_1274);
or U1552 (N_1552,N_1372,N_1202);
or U1553 (N_1553,N_1369,N_1384);
nor U1554 (N_1554,N_1200,N_1280);
xnor U1555 (N_1555,N_1254,N_1352);
and U1556 (N_1556,N_1229,N_1365);
nand U1557 (N_1557,N_1250,N_1350);
nand U1558 (N_1558,N_1392,N_1340);
xnor U1559 (N_1559,N_1237,N_1211);
and U1560 (N_1560,N_1223,N_1276);
and U1561 (N_1561,N_1286,N_1320);
xor U1562 (N_1562,N_1334,N_1323);
or U1563 (N_1563,N_1219,N_1241);
or U1564 (N_1564,N_1325,N_1275);
and U1565 (N_1565,N_1371,N_1312);
nand U1566 (N_1566,N_1224,N_1312);
and U1567 (N_1567,N_1249,N_1349);
and U1568 (N_1568,N_1233,N_1375);
xor U1569 (N_1569,N_1274,N_1251);
nand U1570 (N_1570,N_1337,N_1344);
xor U1571 (N_1571,N_1394,N_1260);
or U1572 (N_1572,N_1319,N_1398);
nor U1573 (N_1573,N_1218,N_1391);
or U1574 (N_1574,N_1321,N_1375);
and U1575 (N_1575,N_1266,N_1325);
xor U1576 (N_1576,N_1315,N_1389);
nor U1577 (N_1577,N_1277,N_1205);
or U1578 (N_1578,N_1327,N_1346);
and U1579 (N_1579,N_1286,N_1224);
and U1580 (N_1580,N_1242,N_1287);
and U1581 (N_1581,N_1219,N_1283);
and U1582 (N_1582,N_1252,N_1395);
and U1583 (N_1583,N_1338,N_1225);
xor U1584 (N_1584,N_1211,N_1399);
and U1585 (N_1585,N_1354,N_1213);
nand U1586 (N_1586,N_1320,N_1301);
xnor U1587 (N_1587,N_1278,N_1310);
xnor U1588 (N_1588,N_1335,N_1362);
xnor U1589 (N_1589,N_1397,N_1370);
and U1590 (N_1590,N_1331,N_1296);
nor U1591 (N_1591,N_1265,N_1373);
nor U1592 (N_1592,N_1302,N_1385);
xor U1593 (N_1593,N_1262,N_1246);
xor U1594 (N_1594,N_1216,N_1324);
nand U1595 (N_1595,N_1203,N_1340);
xnor U1596 (N_1596,N_1231,N_1307);
nand U1597 (N_1597,N_1328,N_1368);
and U1598 (N_1598,N_1315,N_1243);
nand U1599 (N_1599,N_1291,N_1280);
nor U1600 (N_1600,N_1482,N_1408);
nand U1601 (N_1601,N_1527,N_1459);
nand U1602 (N_1602,N_1471,N_1457);
and U1603 (N_1603,N_1575,N_1590);
xnor U1604 (N_1604,N_1544,N_1450);
or U1605 (N_1605,N_1487,N_1550);
and U1606 (N_1606,N_1489,N_1571);
xor U1607 (N_1607,N_1474,N_1455);
or U1608 (N_1608,N_1593,N_1461);
and U1609 (N_1609,N_1444,N_1421);
nand U1610 (N_1610,N_1418,N_1448);
and U1611 (N_1611,N_1599,N_1522);
xor U1612 (N_1612,N_1507,N_1557);
and U1613 (N_1613,N_1484,N_1402);
or U1614 (N_1614,N_1485,N_1486);
nand U1615 (N_1615,N_1505,N_1534);
and U1616 (N_1616,N_1436,N_1528);
nand U1617 (N_1617,N_1560,N_1465);
xor U1618 (N_1618,N_1462,N_1532);
and U1619 (N_1619,N_1401,N_1563);
or U1620 (N_1620,N_1502,N_1515);
nand U1621 (N_1621,N_1434,N_1420);
nor U1622 (N_1622,N_1517,N_1556);
and U1623 (N_1623,N_1539,N_1536);
or U1624 (N_1624,N_1520,N_1558);
xor U1625 (N_1625,N_1537,N_1463);
nor U1626 (N_1626,N_1559,N_1498);
or U1627 (N_1627,N_1501,N_1430);
nand U1628 (N_1628,N_1577,N_1549);
nand U1629 (N_1629,N_1578,N_1404);
xnor U1630 (N_1630,N_1415,N_1525);
or U1631 (N_1631,N_1460,N_1592);
nand U1632 (N_1632,N_1542,N_1546);
nor U1633 (N_1633,N_1409,N_1519);
or U1634 (N_1634,N_1424,N_1586);
nand U1635 (N_1635,N_1561,N_1456);
nand U1636 (N_1636,N_1545,N_1552);
or U1637 (N_1637,N_1447,N_1597);
nand U1638 (N_1638,N_1412,N_1548);
nor U1639 (N_1639,N_1429,N_1425);
nor U1640 (N_1640,N_1446,N_1508);
nand U1641 (N_1641,N_1510,N_1411);
nand U1642 (N_1642,N_1538,N_1530);
xor U1643 (N_1643,N_1580,N_1506);
and U1644 (N_1644,N_1574,N_1466);
and U1645 (N_1645,N_1454,N_1467);
nor U1646 (N_1646,N_1531,N_1477);
and U1647 (N_1647,N_1405,N_1400);
or U1648 (N_1648,N_1523,N_1449);
xor U1649 (N_1649,N_1595,N_1504);
or U1650 (N_1650,N_1582,N_1569);
nand U1651 (N_1651,N_1540,N_1441);
xnor U1652 (N_1652,N_1493,N_1416);
or U1653 (N_1653,N_1438,N_1562);
and U1654 (N_1654,N_1514,N_1570);
nor U1655 (N_1655,N_1588,N_1494);
nand U1656 (N_1656,N_1589,N_1598);
nand U1657 (N_1657,N_1572,N_1594);
nor U1658 (N_1658,N_1553,N_1407);
or U1659 (N_1659,N_1426,N_1555);
and U1660 (N_1660,N_1473,N_1497);
or U1661 (N_1661,N_1496,N_1458);
or U1662 (N_1662,N_1432,N_1541);
xnor U1663 (N_1663,N_1480,N_1413);
xnor U1664 (N_1664,N_1451,N_1521);
nand U1665 (N_1665,N_1453,N_1568);
or U1666 (N_1666,N_1435,N_1472);
and U1667 (N_1667,N_1512,N_1499);
nand U1668 (N_1668,N_1481,N_1437);
xnor U1669 (N_1669,N_1591,N_1410);
or U1670 (N_1670,N_1535,N_1583);
and U1671 (N_1671,N_1442,N_1547);
and U1672 (N_1672,N_1516,N_1470);
and U1673 (N_1673,N_1526,N_1524);
nor U1674 (N_1674,N_1427,N_1576);
nor U1675 (N_1675,N_1428,N_1488);
xor U1676 (N_1676,N_1511,N_1551);
nor U1677 (N_1677,N_1495,N_1509);
xor U1678 (N_1678,N_1584,N_1478);
or U1679 (N_1679,N_1500,N_1483);
xnor U1680 (N_1680,N_1513,N_1439);
and U1681 (N_1681,N_1518,N_1567);
xor U1682 (N_1682,N_1468,N_1596);
nand U1683 (N_1683,N_1452,N_1581);
nor U1684 (N_1684,N_1479,N_1579);
xor U1685 (N_1685,N_1554,N_1464);
xnor U1686 (N_1686,N_1423,N_1573);
xnor U1687 (N_1687,N_1503,N_1443);
nor U1688 (N_1688,N_1476,N_1585);
nand U1689 (N_1689,N_1469,N_1433);
and U1690 (N_1690,N_1440,N_1587);
or U1691 (N_1691,N_1417,N_1419);
and U1692 (N_1692,N_1445,N_1564);
nand U1693 (N_1693,N_1414,N_1543);
nor U1694 (N_1694,N_1422,N_1565);
nand U1695 (N_1695,N_1529,N_1403);
nand U1696 (N_1696,N_1533,N_1491);
or U1697 (N_1697,N_1490,N_1475);
nor U1698 (N_1698,N_1566,N_1431);
xor U1699 (N_1699,N_1492,N_1406);
and U1700 (N_1700,N_1477,N_1457);
nand U1701 (N_1701,N_1566,N_1444);
xnor U1702 (N_1702,N_1406,N_1497);
nor U1703 (N_1703,N_1539,N_1517);
nor U1704 (N_1704,N_1536,N_1529);
and U1705 (N_1705,N_1502,N_1513);
and U1706 (N_1706,N_1533,N_1585);
or U1707 (N_1707,N_1590,N_1531);
nand U1708 (N_1708,N_1566,N_1557);
xnor U1709 (N_1709,N_1500,N_1514);
nand U1710 (N_1710,N_1511,N_1426);
nor U1711 (N_1711,N_1542,N_1590);
and U1712 (N_1712,N_1593,N_1469);
or U1713 (N_1713,N_1583,N_1576);
xnor U1714 (N_1714,N_1540,N_1498);
nor U1715 (N_1715,N_1499,N_1487);
xnor U1716 (N_1716,N_1489,N_1511);
nand U1717 (N_1717,N_1548,N_1481);
nor U1718 (N_1718,N_1549,N_1515);
and U1719 (N_1719,N_1419,N_1565);
or U1720 (N_1720,N_1462,N_1416);
or U1721 (N_1721,N_1544,N_1460);
nand U1722 (N_1722,N_1530,N_1493);
nand U1723 (N_1723,N_1581,N_1563);
nand U1724 (N_1724,N_1463,N_1470);
or U1725 (N_1725,N_1576,N_1570);
and U1726 (N_1726,N_1594,N_1541);
or U1727 (N_1727,N_1499,N_1448);
nor U1728 (N_1728,N_1478,N_1445);
and U1729 (N_1729,N_1446,N_1435);
xor U1730 (N_1730,N_1573,N_1480);
or U1731 (N_1731,N_1444,N_1467);
nand U1732 (N_1732,N_1503,N_1491);
nor U1733 (N_1733,N_1538,N_1565);
or U1734 (N_1734,N_1545,N_1447);
nor U1735 (N_1735,N_1589,N_1409);
nand U1736 (N_1736,N_1407,N_1574);
nand U1737 (N_1737,N_1457,N_1541);
or U1738 (N_1738,N_1469,N_1465);
and U1739 (N_1739,N_1595,N_1405);
and U1740 (N_1740,N_1492,N_1401);
and U1741 (N_1741,N_1592,N_1566);
nand U1742 (N_1742,N_1523,N_1411);
xor U1743 (N_1743,N_1537,N_1505);
xor U1744 (N_1744,N_1531,N_1528);
nand U1745 (N_1745,N_1409,N_1523);
and U1746 (N_1746,N_1412,N_1539);
and U1747 (N_1747,N_1580,N_1441);
or U1748 (N_1748,N_1404,N_1514);
xnor U1749 (N_1749,N_1462,N_1526);
or U1750 (N_1750,N_1510,N_1582);
and U1751 (N_1751,N_1542,N_1428);
or U1752 (N_1752,N_1499,N_1492);
xor U1753 (N_1753,N_1415,N_1414);
nand U1754 (N_1754,N_1468,N_1569);
and U1755 (N_1755,N_1416,N_1538);
and U1756 (N_1756,N_1438,N_1525);
and U1757 (N_1757,N_1539,N_1402);
or U1758 (N_1758,N_1539,N_1483);
or U1759 (N_1759,N_1554,N_1521);
or U1760 (N_1760,N_1509,N_1543);
and U1761 (N_1761,N_1475,N_1409);
xor U1762 (N_1762,N_1408,N_1558);
and U1763 (N_1763,N_1473,N_1498);
nor U1764 (N_1764,N_1458,N_1549);
nand U1765 (N_1765,N_1417,N_1407);
and U1766 (N_1766,N_1521,N_1583);
or U1767 (N_1767,N_1491,N_1453);
xnor U1768 (N_1768,N_1496,N_1512);
nand U1769 (N_1769,N_1548,N_1552);
xnor U1770 (N_1770,N_1497,N_1477);
and U1771 (N_1771,N_1494,N_1573);
and U1772 (N_1772,N_1511,N_1598);
nand U1773 (N_1773,N_1596,N_1474);
and U1774 (N_1774,N_1589,N_1470);
nand U1775 (N_1775,N_1470,N_1580);
and U1776 (N_1776,N_1492,N_1479);
and U1777 (N_1777,N_1500,N_1420);
or U1778 (N_1778,N_1417,N_1500);
nand U1779 (N_1779,N_1447,N_1423);
nor U1780 (N_1780,N_1596,N_1439);
xnor U1781 (N_1781,N_1456,N_1572);
or U1782 (N_1782,N_1466,N_1580);
nor U1783 (N_1783,N_1493,N_1548);
and U1784 (N_1784,N_1568,N_1598);
or U1785 (N_1785,N_1597,N_1410);
nor U1786 (N_1786,N_1499,N_1510);
nor U1787 (N_1787,N_1529,N_1506);
xnor U1788 (N_1788,N_1453,N_1403);
xor U1789 (N_1789,N_1434,N_1433);
xnor U1790 (N_1790,N_1401,N_1571);
xnor U1791 (N_1791,N_1584,N_1492);
and U1792 (N_1792,N_1483,N_1453);
xnor U1793 (N_1793,N_1417,N_1511);
nor U1794 (N_1794,N_1411,N_1525);
nand U1795 (N_1795,N_1462,N_1426);
or U1796 (N_1796,N_1456,N_1448);
and U1797 (N_1797,N_1515,N_1573);
and U1798 (N_1798,N_1424,N_1482);
or U1799 (N_1799,N_1461,N_1440);
or U1800 (N_1800,N_1600,N_1745);
and U1801 (N_1801,N_1603,N_1721);
nand U1802 (N_1802,N_1699,N_1679);
nor U1803 (N_1803,N_1642,N_1734);
or U1804 (N_1804,N_1615,N_1628);
xnor U1805 (N_1805,N_1633,N_1713);
and U1806 (N_1806,N_1617,N_1666);
and U1807 (N_1807,N_1724,N_1761);
xor U1808 (N_1808,N_1795,N_1712);
xnor U1809 (N_1809,N_1657,N_1709);
and U1810 (N_1810,N_1634,N_1707);
xor U1811 (N_1811,N_1790,N_1669);
xor U1812 (N_1812,N_1613,N_1741);
nand U1813 (N_1813,N_1706,N_1694);
xnor U1814 (N_1814,N_1665,N_1675);
or U1815 (N_1815,N_1775,N_1607);
nor U1816 (N_1816,N_1701,N_1744);
or U1817 (N_1817,N_1729,N_1755);
nand U1818 (N_1818,N_1683,N_1627);
nor U1819 (N_1819,N_1614,N_1636);
and U1820 (N_1820,N_1635,N_1770);
nand U1821 (N_1821,N_1749,N_1681);
xnor U1822 (N_1822,N_1791,N_1677);
nor U1823 (N_1823,N_1786,N_1726);
or U1824 (N_1824,N_1710,N_1758);
xor U1825 (N_1825,N_1774,N_1624);
or U1826 (N_1826,N_1678,N_1640);
and U1827 (N_1827,N_1605,N_1731);
xor U1828 (N_1828,N_1757,N_1672);
nand U1829 (N_1829,N_1716,N_1697);
and U1830 (N_1830,N_1663,N_1644);
xor U1831 (N_1831,N_1739,N_1736);
nand U1832 (N_1832,N_1629,N_1743);
and U1833 (N_1833,N_1771,N_1751);
nor U1834 (N_1834,N_1652,N_1647);
nand U1835 (N_1835,N_1784,N_1610);
nand U1836 (N_1836,N_1655,N_1674);
and U1837 (N_1837,N_1623,N_1715);
nand U1838 (N_1838,N_1703,N_1718);
nand U1839 (N_1839,N_1714,N_1648);
xor U1840 (N_1840,N_1651,N_1686);
and U1841 (N_1841,N_1684,N_1766);
nand U1842 (N_1842,N_1602,N_1732);
nand U1843 (N_1843,N_1711,N_1671);
and U1844 (N_1844,N_1772,N_1781);
xnor U1845 (N_1845,N_1619,N_1753);
or U1846 (N_1846,N_1612,N_1782);
xor U1847 (N_1847,N_1685,N_1785);
nor U1848 (N_1848,N_1689,N_1763);
and U1849 (N_1849,N_1787,N_1611);
nor U1850 (N_1850,N_1777,N_1680);
nor U1851 (N_1851,N_1720,N_1691);
nor U1852 (N_1852,N_1606,N_1779);
nor U1853 (N_1853,N_1727,N_1760);
xnor U1854 (N_1854,N_1705,N_1673);
xnor U1855 (N_1855,N_1696,N_1667);
nand U1856 (N_1856,N_1661,N_1631);
and U1857 (N_1857,N_1654,N_1735);
nor U1858 (N_1858,N_1670,N_1659);
xnor U1859 (N_1859,N_1719,N_1643);
or U1860 (N_1860,N_1740,N_1658);
and U1861 (N_1861,N_1778,N_1622);
nor U1862 (N_1862,N_1796,N_1682);
nand U1863 (N_1863,N_1645,N_1730);
nand U1864 (N_1864,N_1797,N_1793);
or U1865 (N_1865,N_1768,N_1641);
nor U1866 (N_1866,N_1653,N_1733);
nor U1867 (N_1867,N_1687,N_1792);
nand U1868 (N_1868,N_1637,N_1752);
and U1869 (N_1869,N_1626,N_1649);
nand U1870 (N_1870,N_1692,N_1688);
xor U1871 (N_1871,N_1767,N_1601);
xor U1872 (N_1872,N_1620,N_1656);
xnor U1873 (N_1873,N_1765,N_1738);
xor U1874 (N_1874,N_1695,N_1723);
nor U1875 (N_1875,N_1754,N_1748);
xnor U1876 (N_1876,N_1632,N_1630);
or U1877 (N_1877,N_1646,N_1788);
xnor U1878 (N_1878,N_1783,N_1717);
nor U1879 (N_1879,N_1728,N_1604);
nor U1880 (N_1880,N_1780,N_1700);
or U1881 (N_1881,N_1750,N_1693);
or U1882 (N_1882,N_1794,N_1722);
and U1883 (N_1883,N_1725,N_1776);
nand U1884 (N_1884,N_1756,N_1708);
nand U1885 (N_1885,N_1704,N_1676);
xor U1886 (N_1886,N_1702,N_1746);
nand U1887 (N_1887,N_1737,N_1608);
nor U1888 (N_1888,N_1639,N_1668);
nand U1889 (N_1889,N_1762,N_1638);
or U1890 (N_1890,N_1662,N_1742);
xor U1891 (N_1891,N_1625,N_1747);
or U1892 (N_1892,N_1609,N_1618);
and U1893 (N_1893,N_1616,N_1769);
or U1894 (N_1894,N_1660,N_1650);
xnor U1895 (N_1895,N_1621,N_1799);
nand U1896 (N_1896,N_1664,N_1764);
and U1897 (N_1897,N_1690,N_1798);
nand U1898 (N_1898,N_1698,N_1759);
nor U1899 (N_1899,N_1773,N_1789);
nor U1900 (N_1900,N_1706,N_1656);
and U1901 (N_1901,N_1652,N_1663);
nand U1902 (N_1902,N_1743,N_1657);
or U1903 (N_1903,N_1707,N_1708);
xnor U1904 (N_1904,N_1761,N_1686);
nand U1905 (N_1905,N_1711,N_1757);
nor U1906 (N_1906,N_1670,N_1600);
xor U1907 (N_1907,N_1618,N_1708);
or U1908 (N_1908,N_1630,N_1696);
and U1909 (N_1909,N_1723,N_1604);
or U1910 (N_1910,N_1642,N_1765);
nand U1911 (N_1911,N_1719,N_1672);
or U1912 (N_1912,N_1790,N_1712);
or U1913 (N_1913,N_1787,N_1656);
or U1914 (N_1914,N_1739,N_1676);
nor U1915 (N_1915,N_1642,N_1770);
nand U1916 (N_1916,N_1650,N_1667);
or U1917 (N_1917,N_1669,N_1698);
nor U1918 (N_1918,N_1720,N_1688);
nand U1919 (N_1919,N_1753,N_1644);
nor U1920 (N_1920,N_1656,N_1674);
and U1921 (N_1921,N_1630,N_1670);
nand U1922 (N_1922,N_1727,N_1613);
or U1923 (N_1923,N_1639,N_1600);
or U1924 (N_1924,N_1765,N_1627);
and U1925 (N_1925,N_1762,N_1702);
and U1926 (N_1926,N_1751,N_1691);
and U1927 (N_1927,N_1665,N_1699);
xnor U1928 (N_1928,N_1720,N_1664);
nor U1929 (N_1929,N_1788,N_1796);
nor U1930 (N_1930,N_1686,N_1642);
nand U1931 (N_1931,N_1634,N_1686);
xnor U1932 (N_1932,N_1706,N_1763);
xnor U1933 (N_1933,N_1773,N_1696);
and U1934 (N_1934,N_1723,N_1642);
or U1935 (N_1935,N_1703,N_1635);
and U1936 (N_1936,N_1775,N_1695);
nand U1937 (N_1937,N_1654,N_1797);
xor U1938 (N_1938,N_1606,N_1611);
and U1939 (N_1939,N_1693,N_1699);
or U1940 (N_1940,N_1681,N_1604);
and U1941 (N_1941,N_1651,N_1792);
and U1942 (N_1942,N_1690,N_1682);
nor U1943 (N_1943,N_1698,N_1605);
nand U1944 (N_1944,N_1789,N_1710);
xnor U1945 (N_1945,N_1671,N_1736);
and U1946 (N_1946,N_1777,N_1699);
nand U1947 (N_1947,N_1726,N_1698);
xor U1948 (N_1948,N_1690,N_1674);
or U1949 (N_1949,N_1728,N_1741);
or U1950 (N_1950,N_1788,N_1619);
and U1951 (N_1951,N_1653,N_1774);
and U1952 (N_1952,N_1788,N_1789);
and U1953 (N_1953,N_1742,N_1761);
nand U1954 (N_1954,N_1610,N_1732);
nor U1955 (N_1955,N_1650,N_1620);
nand U1956 (N_1956,N_1770,N_1656);
or U1957 (N_1957,N_1783,N_1646);
or U1958 (N_1958,N_1685,N_1719);
nand U1959 (N_1959,N_1692,N_1732);
or U1960 (N_1960,N_1642,N_1662);
and U1961 (N_1961,N_1741,N_1756);
nand U1962 (N_1962,N_1727,N_1685);
xnor U1963 (N_1963,N_1727,N_1654);
xnor U1964 (N_1964,N_1663,N_1773);
and U1965 (N_1965,N_1710,N_1716);
xnor U1966 (N_1966,N_1734,N_1776);
xor U1967 (N_1967,N_1786,N_1784);
nand U1968 (N_1968,N_1738,N_1697);
nand U1969 (N_1969,N_1794,N_1611);
or U1970 (N_1970,N_1652,N_1635);
xor U1971 (N_1971,N_1629,N_1622);
xnor U1972 (N_1972,N_1602,N_1786);
nor U1973 (N_1973,N_1790,N_1747);
xor U1974 (N_1974,N_1710,N_1697);
and U1975 (N_1975,N_1608,N_1699);
nand U1976 (N_1976,N_1656,N_1778);
xor U1977 (N_1977,N_1764,N_1711);
or U1978 (N_1978,N_1682,N_1732);
or U1979 (N_1979,N_1612,N_1668);
or U1980 (N_1980,N_1729,N_1624);
or U1981 (N_1981,N_1790,N_1670);
nand U1982 (N_1982,N_1655,N_1780);
or U1983 (N_1983,N_1751,N_1670);
xor U1984 (N_1984,N_1781,N_1659);
nor U1985 (N_1985,N_1614,N_1658);
or U1986 (N_1986,N_1706,N_1734);
xnor U1987 (N_1987,N_1745,N_1612);
and U1988 (N_1988,N_1788,N_1756);
and U1989 (N_1989,N_1725,N_1787);
or U1990 (N_1990,N_1667,N_1775);
nand U1991 (N_1991,N_1702,N_1743);
nor U1992 (N_1992,N_1677,N_1794);
or U1993 (N_1993,N_1731,N_1797);
or U1994 (N_1994,N_1664,N_1673);
or U1995 (N_1995,N_1657,N_1726);
or U1996 (N_1996,N_1639,N_1727);
nor U1997 (N_1997,N_1794,N_1676);
nor U1998 (N_1998,N_1654,N_1676);
and U1999 (N_1999,N_1646,N_1765);
nor U2000 (N_2000,N_1977,N_1868);
nor U2001 (N_2001,N_1955,N_1820);
or U2002 (N_2002,N_1870,N_1986);
and U2003 (N_2003,N_1865,N_1834);
xnor U2004 (N_2004,N_1911,N_1860);
or U2005 (N_2005,N_1824,N_1928);
and U2006 (N_2006,N_1972,N_1937);
nand U2007 (N_2007,N_1866,N_1848);
or U2008 (N_2008,N_1832,N_1996);
nor U2009 (N_2009,N_1948,N_1959);
nor U2010 (N_2010,N_1927,N_1828);
xor U2011 (N_2011,N_1920,N_1817);
nand U2012 (N_2012,N_1953,N_1852);
nand U2013 (N_2013,N_1898,N_1935);
xnor U2014 (N_2014,N_1992,N_1932);
nor U2015 (N_2015,N_1821,N_1809);
or U2016 (N_2016,N_1900,N_1819);
or U2017 (N_2017,N_1889,N_1947);
nand U2018 (N_2018,N_1874,N_1843);
and U2019 (N_2019,N_1966,N_1867);
nor U2020 (N_2020,N_1837,N_1940);
nor U2021 (N_2021,N_1985,N_1905);
or U2022 (N_2022,N_1897,N_1842);
nor U2023 (N_2023,N_1855,N_1857);
and U2024 (N_2024,N_1805,N_1949);
nor U2025 (N_2025,N_1831,N_1983);
nand U2026 (N_2026,N_1803,N_1894);
nor U2027 (N_2027,N_1896,N_1929);
and U2028 (N_2028,N_1850,N_1906);
and U2029 (N_2029,N_1862,N_1825);
xor U2030 (N_2030,N_1919,N_1933);
and U2031 (N_2031,N_1816,N_1875);
nor U2032 (N_2032,N_1807,N_1808);
xnor U2033 (N_2033,N_1962,N_1987);
xnor U2034 (N_2034,N_1886,N_1901);
and U2035 (N_2035,N_1846,N_1892);
or U2036 (N_2036,N_1888,N_1995);
xor U2037 (N_2037,N_1936,N_1956);
or U2038 (N_2038,N_1941,N_1934);
and U2039 (N_2039,N_1810,N_1858);
and U2040 (N_2040,N_1943,N_1993);
xor U2041 (N_2041,N_1957,N_1944);
xnor U2042 (N_2042,N_1801,N_1904);
xnor U2043 (N_2043,N_1954,N_1938);
nor U2044 (N_2044,N_1836,N_1835);
or U2045 (N_2045,N_1833,N_1881);
and U2046 (N_2046,N_1980,N_1890);
nand U2047 (N_2047,N_1974,N_1965);
or U2048 (N_2048,N_1829,N_1970);
xnor U2049 (N_2049,N_1907,N_1856);
or U2050 (N_2050,N_1984,N_1840);
nand U2051 (N_2051,N_1861,N_1961);
xnor U2052 (N_2052,N_1818,N_1945);
or U2053 (N_2053,N_1998,N_1990);
xnor U2054 (N_2054,N_1916,N_1849);
and U2055 (N_2055,N_1981,N_1847);
nand U2056 (N_2056,N_1978,N_1882);
xor U2057 (N_2057,N_1899,N_1815);
and U2058 (N_2058,N_1921,N_1909);
nand U2059 (N_2059,N_1991,N_1873);
and U2060 (N_2060,N_1902,N_1924);
nand U2061 (N_2061,N_1878,N_1960);
or U2062 (N_2062,N_1925,N_1922);
and U2063 (N_2063,N_1917,N_1811);
nor U2064 (N_2064,N_1964,N_1913);
and U2065 (N_2065,N_1872,N_1876);
nor U2066 (N_2066,N_1958,N_1999);
and U2067 (N_2067,N_1891,N_1931);
xnor U2068 (N_2068,N_1883,N_1885);
nor U2069 (N_2069,N_1839,N_1830);
or U2070 (N_2070,N_1826,N_1994);
xor U2071 (N_2071,N_1942,N_1869);
nand U2072 (N_2072,N_1841,N_1845);
and U2073 (N_2073,N_1879,N_1908);
xor U2074 (N_2074,N_1884,N_1814);
nor U2075 (N_2075,N_1915,N_1968);
nor U2076 (N_2076,N_1880,N_1950);
xor U2077 (N_2077,N_1822,N_1853);
and U2078 (N_2078,N_1895,N_1975);
nor U2079 (N_2079,N_1806,N_1813);
and U2080 (N_2080,N_1887,N_1989);
and U2081 (N_2081,N_1971,N_1914);
xor U2082 (N_2082,N_1812,N_1923);
or U2083 (N_2083,N_1804,N_1973);
and U2084 (N_2084,N_1800,N_1802);
and U2085 (N_2085,N_1838,N_1859);
or U2086 (N_2086,N_1926,N_1951);
xnor U2087 (N_2087,N_1863,N_1930);
nor U2088 (N_2088,N_1979,N_1893);
and U2089 (N_2089,N_1997,N_1823);
nand U2090 (N_2090,N_1939,N_1967);
and U2091 (N_2091,N_1969,N_1877);
xnor U2092 (N_2092,N_1871,N_1963);
xnor U2093 (N_2093,N_1918,N_1946);
nand U2094 (N_2094,N_1827,N_1982);
nor U2095 (N_2095,N_1844,N_1988);
nor U2096 (N_2096,N_1864,N_1910);
nand U2097 (N_2097,N_1976,N_1851);
xnor U2098 (N_2098,N_1903,N_1952);
nand U2099 (N_2099,N_1912,N_1854);
xor U2100 (N_2100,N_1926,N_1999);
and U2101 (N_2101,N_1948,N_1898);
nand U2102 (N_2102,N_1873,N_1912);
and U2103 (N_2103,N_1830,N_1954);
or U2104 (N_2104,N_1932,N_1848);
and U2105 (N_2105,N_1916,N_1967);
nor U2106 (N_2106,N_1995,N_1939);
xor U2107 (N_2107,N_1839,N_1928);
nand U2108 (N_2108,N_1922,N_1957);
and U2109 (N_2109,N_1922,N_1868);
xor U2110 (N_2110,N_1951,N_1806);
nor U2111 (N_2111,N_1986,N_1811);
nor U2112 (N_2112,N_1952,N_1955);
nand U2113 (N_2113,N_1801,N_1949);
and U2114 (N_2114,N_1920,N_1826);
nor U2115 (N_2115,N_1950,N_1850);
xnor U2116 (N_2116,N_1845,N_1956);
and U2117 (N_2117,N_1832,N_1813);
nor U2118 (N_2118,N_1879,N_1942);
xnor U2119 (N_2119,N_1931,N_1989);
or U2120 (N_2120,N_1999,N_1970);
nor U2121 (N_2121,N_1973,N_1832);
and U2122 (N_2122,N_1891,N_1904);
or U2123 (N_2123,N_1917,N_1994);
xnor U2124 (N_2124,N_1978,N_1935);
xor U2125 (N_2125,N_1945,N_1832);
or U2126 (N_2126,N_1927,N_1929);
xnor U2127 (N_2127,N_1855,N_1937);
xnor U2128 (N_2128,N_1983,N_1920);
and U2129 (N_2129,N_1808,N_1916);
or U2130 (N_2130,N_1884,N_1926);
nand U2131 (N_2131,N_1812,N_1870);
xor U2132 (N_2132,N_1905,N_1804);
xor U2133 (N_2133,N_1890,N_1880);
nor U2134 (N_2134,N_1900,N_1860);
nor U2135 (N_2135,N_1873,N_1993);
xnor U2136 (N_2136,N_1868,N_1899);
nand U2137 (N_2137,N_1875,N_1883);
or U2138 (N_2138,N_1907,N_1948);
xnor U2139 (N_2139,N_1810,N_1868);
and U2140 (N_2140,N_1888,N_1988);
nor U2141 (N_2141,N_1817,N_1970);
nand U2142 (N_2142,N_1920,N_1912);
nand U2143 (N_2143,N_1957,N_1836);
nor U2144 (N_2144,N_1836,N_1949);
nor U2145 (N_2145,N_1825,N_1934);
nor U2146 (N_2146,N_1999,N_1971);
and U2147 (N_2147,N_1834,N_1803);
and U2148 (N_2148,N_1971,N_1985);
xor U2149 (N_2149,N_1822,N_1940);
nor U2150 (N_2150,N_1849,N_1851);
nor U2151 (N_2151,N_1992,N_1888);
xor U2152 (N_2152,N_1851,N_1886);
nor U2153 (N_2153,N_1954,N_1871);
nand U2154 (N_2154,N_1959,N_1966);
nor U2155 (N_2155,N_1962,N_1938);
nand U2156 (N_2156,N_1942,N_1900);
and U2157 (N_2157,N_1939,N_1907);
nor U2158 (N_2158,N_1866,N_1873);
nand U2159 (N_2159,N_1871,N_1886);
nor U2160 (N_2160,N_1889,N_1911);
nor U2161 (N_2161,N_1892,N_1923);
and U2162 (N_2162,N_1857,N_1905);
or U2163 (N_2163,N_1993,N_1820);
nand U2164 (N_2164,N_1914,N_1844);
xnor U2165 (N_2165,N_1813,N_1914);
xnor U2166 (N_2166,N_1880,N_1852);
or U2167 (N_2167,N_1864,N_1894);
nand U2168 (N_2168,N_1906,N_1820);
xor U2169 (N_2169,N_1985,N_1955);
nor U2170 (N_2170,N_1844,N_1964);
nand U2171 (N_2171,N_1856,N_1909);
and U2172 (N_2172,N_1890,N_1843);
xnor U2173 (N_2173,N_1866,N_1918);
xnor U2174 (N_2174,N_1916,N_1930);
or U2175 (N_2175,N_1923,N_1911);
nand U2176 (N_2176,N_1830,N_1874);
or U2177 (N_2177,N_1992,N_1864);
or U2178 (N_2178,N_1957,N_1994);
or U2179 (N_2179,N_1968,N_1898);
nand U2180 (N_2180,N_1950,N_1894);
and U2181 (N_2181,N_1880,N_1911);
nor U2182 (N_2182,N_1922,N_1851);
and U2183 (N_2183,N_1901,N_1884);
nand U2184 (N_2184,N_1995,N_1942);
and U2185 (N_2185,N_1952,N_1904);
xor U2186 (N_2186,N_1931,N_1827);
and U2187 (N_2187,N_1891,N_1824);
nand U2188 (N_2188,N_1954,N_1924);
nand U2189 (N_2189,N_1845,N_1867);
or U2190 (N_2190,N_1999,N_1916);
nand U2191 (N_2191,N_1887,N_1943);
or U2192 (N_2192,N_1818,N_1912);
or U2193 (N_2193,N_1875,N_1839);
nand U2194 (N_2194,N_1936,N_1809);
or U2195 (N_2195,N_1892,N_1930);
and U2196 (N_2196,N_1845,N_1801);
or U2197 (N_2197,N_1891,N_1897);
and U2198 (N_2198,N_1990,N_1932);
or U2199 (N_2199,N_1891,N_1985);
and U2200 (N_2200,N_2040,N_2139);
nand U2201 (N_2201,N_2008,N_2001);
nor U2202 (N_2202,N_2029,N_2034);
and U2203 (N_2203,N_2180,N_2030);
nand U2204 (N_2204,N_2094,N_2053);
nor U2205 (N_2205,N_2010,N_2113);
and U2206 (N_2206,N_2133,N_2088);
nand U2207 (N_2207,N_2079,N_2099);
or U2208 (N_2208,N_2157,N_2130);
and U2209 (N_2209,N_2061,N_2036);
nor U2210 (N_2210,N_2059,N_2006);
nand U2211 (N_2211,N_2039,N_2116);
or U2212 (N_2212,N_2048,N_2177);
and U2213 (N_2213,N_2056,N_2024);
nand U2214 (N_2214,N_2120,N_2102);
nand U2215 (N_2215,N_2142,N_2109);
or U2216 (N_2216,N_2032,N_2162);
or U2217 (N_2217,N_2075,N_2161);
and U2218 (N_2218,N_2035,N_2178);
nand U2219 (N_2219,N_2123,N_2082);
nor U2220 (N_2220,N_2141,N_2144);
nand U2221 (N_2221,N_2004,N_2044);
or U2222 (N_2222,N_2000,N_2012);
nand U2223 (N_2223,N_2126,N_2045);
nor U2224 (N_2224,N_2092,N_2132);
nand U2225 (N_2225,N_2190,N_2009);
or U2226 (N_2226,N_2191,N_2192);
nor U2227 (N_2227,N_2063,N_2086);
nor U2228 (N_2228,N_2124,N_2081);
or U2229 (N_2229,N_2198,N_2050);
and U2230 (N_2230,N_2149,N_2005);
xnor U2231 (N_2231,N_2041,N_2026);
nor U2232 (N_2232,N_2080,N_2084);
or U2233 (N_2233,N_2154,N_2076);
nand U2234 (N_2234,N_2135,N_2066);
nand U2235 (N_2235,N_2042,N_2196);
and U2236 (N_2236,N_2060,N_2051);
nor U2237 (N_2237,N_2095,N_2007);
nand U2238 (N_2238,N_2020,N_2171);
nand U2239 (N_2239,N_2110,N_2011);
nor U2240 (N_2240,N_2098,N_2121);
or U2241 (N_2241,N_2071,N_2025);
or U2242 (N_2242,N_2166,N_2115);
nor U2243 (N_2243,N_2176,N_2072);
nand U2244 (N_2244,N_2114,N_2002);
nor U2245 (N_2245,N_2182,N_2138);
and U2246 (N_2246,N_2065,N_2043);
or U2247 (N_2247,N_2125,N_2188);
nor U2248 (N_2248,N_2021,N_2189);
or U2249 (N_2249,N_2159,N_2147);
nand U2250 (N_2250,N_2090,N_2073);
nand U2251 (N_2251,N_2187,N_2105);
nand U2252 (N_2252,N_2155,N_2019);
and U2253 (N_2253,N_2055,N_2070);
nor U2254 (N_2254,N_2134,N_2028);
nor U2255 (N_2255,N_2104,N_2103);
xor U2256 (N_2256,N_2127,N_2118);
nand U2257 (N_2257,N_2184,N_2186);
nand U2258 (N_2258,N_2137,N_2089);
xor U2259 (N_2259,N_2146,N_2100);
nand U2260 (N_2260,N_2129,N_2172);
xor U2261 (N_2261,N_2093,N_2068);
and U2262 (N_2262,N_2195,N_2163);
or U2263 (N_2263,N_2122,N_2153);
nor U2264 (N_2264,N_2181,N_2033);
xor U2265 (N_2265,N_2049,N_2128);
or U2266 (N_2266,N_2015,N_2062);
xor U2267 (N_2267,N_2143,N_2197);
and U2268 (N_2268,N_2087,N_2031);
xor U2269 (N_2269,N_2047,N_2194);
xor U2270 (N_2270,N_2052,N_2136);
nand U2271 (N_2271,N_2111,N_2077);
nor U2272 (N_2272,N_2046,N_2064);
or U2273 (N_2273,N_2151,N_2106);
or U2274 (N_2274,N_2027,N_2023);
nand U2275 (N_2275,N_2183,N_2174);
nor U2276 (N_2276,N_2091,N_2078);
and U2277 (N_2277,N_2170,N_2168);
nor U2278 (N_2278,N_2107,N_2156);
nor U2279 (N_2279,N_2119,N_2117);
or U2280 (N_2280,N_2185,N_2179);
xnor U2281 (N_2281,N_2096,N_2108);
and U2282 (N_2282,N_2038,N_2022);
xor U2283 (N_2283,N_2158,N_2131);
or U2284 (N_2284,N_2152,N_2083);
nor U2285 (N_2285,N_2069,N_2193);
nand U2286 (N_2286,N_2054,N_2085);
or U2287 (N_2287,N_2017,N_2097);
and U2288 (N_2288,N_2037,N_2175);
nand U2289 (N_2289,N_2164,N_2199);
and U2290 (N_2290,N_2173,N_2067);
nor U2291 (N_2291,N_2112,N_2160);
or U2292 (N_2292,N_2148,N_2018);
nor U2293 (N_2293,N_2013,N_2003);
nand U2294 (N_2294,N_2058,N_2140);
nand U2295 (N_2295,N_2165,N_2014);
or U2296 (N_2296,N_2150,N_2074);
or U2297 (N_2297,N_2101,N_2145);
nand U2298 (N_2298,N_2016,N_2057);
or U2299 (N_2299,N_2169,N_2167);
xor U2300 (N_2300,N_2056,N_2151);
xor U2301 (N_2301,N_2091,N_2105);
xnor U2302 (N_2302,N_2032,N_2193);
xnor U2303 (N_2303,N_2138,N_2040);
nor U2304 (N_2304,N_2061,N_2173);
xor U2305 (N_2305,N_2148,N_2133);
and U2306 (N_2306,N_2199,N_2051);
xor U2307 (N_2307,N_2137,N_2124);
nand U2308 (N_2308,N_2123,N_2034);
nor U2309 (N_2309,N_2087,N_2128);
nand U2310 (N_2310,N_2167,N_2178);
and U2311 (N_2311,N_2129,N_2198);
or U2312 (N_2312,N_2102,N_2197);
nand U2313 (N_2313,N_2047,N_2003);
nor U2314 (N_2314,N_2086,N_2126);
nand U2315 (N_2315,N_2045,N_2075);
xnor U2316 (N_2316,N_2012,N_2133);
or U2317 (N_2317,N_2068,N_2193);
nor U2318 (N_2318,N_2041,N_2060);
or U2319 (N_2319,N_2160,N_2123);
or U2320 (N_2320,N_2174,N_2151);
and U2321 (N_2321,N_2044,N_2107);
or U2322 (N_2322,N_2194,N_2017);
nand U2323 (N_2323,N_2030,N_2142);
or U2324 (N_2324,N_2193,N_2146);
or U2325 (N_2325,N_2189,N_2017);
and U2326 (N_2326,N_2177,N_2016);
or U2327 (N_2327,N_2137,N_2101);
and U2328 (N_2328,N_2123,N_2052);
and U2329 (N_2329,N_2196,N_2157);
or U2330 (N_2330,N_2056,N_2166);
nor U2331 (N_2331,N_2075,N_2083);
nand U2332 (N_2332,N_2128,N_2040);
or U2333 (N_2333,N_2016,N_2075);
and U2334 (N_2334,N_2026,N_2084);
or U2335 (N_2335,N_2147,N_2003);
nor U2336 (N_2336,N_2189,N_2130);
nor U2337 (N_2337,N_2045,N_2068);
and U2338 (N_2338,N_2122,N_2062);
nand U2339 (N_2339,N_2110,N_2033);
nand U2340 (N_2340,N_2036,N_2161);
and U2341 (N_2341,N_2073,N_2199);
or U2342 (N_2342,N_2036,N_2151);
nand U2343 (N_2343,N_2120,N_2079);
nand U2344 (N_2344,N_2103,N_2033);
nor U2345 (N_2345,N_2025,N_2174);
nand U2346 (N_2346,N_2083,N_2060);
nand U2347 (N_2347,N_2019,N_2106);
nand U2348 (N_2348,N_2087,N_2092);
xnor U2349 (N_2349,N_2053,N_2025);
or U2350 (N_2350,N_2089,N_2053);
nor U2351 (N_2351,N_2096,N_2127);
xor U2352 (N_2352,N_2029,N_2010);
nand U2353 (N_2353,N_2185,N_2109);
or U2354 (N_2354,N_2041,N_2021);
or U2355 (N_2355,N_2124,N_2088);
nor U2356 (N_2356,N_2132,N_2033);
nand U2357 (N_2357,N_2141,N_2106);
and U2358 (N_2358,N_2151,N_2014);
nand U2359 (N_2359,N_2039,N_2094);
nand U2360 (N_2360,N_2110,N_2004);
and U2361 (N_2361,N_2027,N_2121);
xnor U2362 (N_2362,N_2051,N_2095);
xor U2363 (N_2363,N_2184,N_2008);
nor U2364 (N_2364,N_2044,N_2093);
xor U2365 (N_2365,N_2032,N_2192);
nand U2366 (N_2366,N_2008,N_2183);
xor U2367 (N_2367,N_2061,N_2019);
xnor U2368 (N_2368,N_2054,N_2157);
nor U2369 (N_2369,N_2194,N_2093);
nand U2370 (N_2370,N_2095,N_2018);
or U2371 (N_2371,N_2069,N_2099);
xnor U2372 (N_2372,N_2129,N_2059);
and U2373 (N_2373,N_2152,N_2036);
and U2374 (N_2374,N_2109,N_2074);
nor U2375 (N_2375,N_2195,N_2143);
nor U2376 (N_2376,N_2104,N_2092);
nor U2377 (N_2377,N_2131,N_2083);
nor U2378 (N_2378,N_2054,N_2136);
xnor U2379 (N_2379,N_2051,N_2193);
nand U2380 (N_2380,N_2170,N_2130);
or U2381 (N_2381,N_2099,N_2041);
xnor U2382 (N_2382,N_2041,N_2027);
nand U2383 (N_2383,N_2035,N_2109);
nor U2384 (N_2384,N_2147,N_2174);
or U2385 (N_2385,N_2194,N_2045);
and U2386 (N_2386,N_2123,N_2177);
nand U2387 (N_2387,N_2123,N_2195);
xnor U2388 (N_2388,N_2095,N_2127);
nand U2389 (N_2389,N_2192,N_2067);
xnor U2390 (N_2390,N_2027,N_2154);
xor U2391 (N_2391,N_2014,N_2135);
nor U2392 (N_2392,N_2016,N_2020);
and U2393 (N_2393,N_2086,N_2027);
or U2394 (N_2394,N_2014,N_2118);
nor U2395 (N_2395,N_2182,N_2178);
xor U2396 (N_2396,N_2187,N_2039);
nor U2397 (N_2397,N_2176,N_2077);
nand U2398 (N_2398,N_2138,N_2197);
nor U2399 (N_2399,N_2199,N_2010);
and U2400 (N_2400,N_2355,N_2268);
xnor U2401 (N_2401,N_2346,N_2212);
nor U2402 (N_2402,N_2226,N_2386);
xnor U2403 (N_2403,N_2250,N_2331);
or U2404 (N_2404,N_2223,N_2233);
nor U2405 (N_2405,N_2351,N_2279);
and U2406 (N_2406,N_2258,N_2265);
xnor U2407 (N_2407,N_2382,N_2254);
and U2408 (N_2408,N_2242,N_2243);
or U2409 (N_2409,N_2240,N_2311);
nor U2410 (N_2410,N_2363,N_2318);
xnor U2411 (N_2411,N_2367,N_2389);
nand U2412 (N_2412,N_2257,N_2287);
xor U2413 (N_2413,N_2307,N_2304);
nor U2414 (N_2414,N_2319,N_2251);
or U2415 (N_2415,N_2353,N_2201);
or U2416 (N_2416,N_2217,N_2350);
and U2417 (N_2417,N_2221,N_2327);
nand U2418 (N_2418,N_2234,N_2248);
xor U2419 (N_2419,N_2393,N_2230);
nor U2420 (N_2420,N_2317,N_2381);
and U2421 (N_2421,N_2328,N_2280);
nor U2422 (N_2422,N_2344,N_2361);
xor U2423 (N_2423,N_2369,N_2371);
nor U2424 (N_2424,N_2272,N_2309);
nand U2425 (N_2425,N_2235,N_2333);
and U2426 (N_2426,N_2261,N_2338);
and U2427 (N_2427,N_2262,N_2335);
and U2428 (N_2428,N_2300,N_2368);
nor U2429 (N_2429,N_2246,N_2339);
nand U2430 (N_2430,N_2360,N_2219);
or U2431 (N_2431,N_2334,N_2378);
xnor U2432 (N_2432,N_2271,N_2241);
nor U2433 (N_2433,N_2380,N_2253);
and U2434 (N_2434,N_2207,N_2315);
or U2435 (N_2435,N_2312,N_2299);
and U2436 (N_2436,N_2236,N_2372);
nand U2437 (N_2437,N_2362,N_2256);
and U2438 (N_2438,N_2216,N_2204);
or U2439 (N_2439,N_2237,N_2354);
nor U2440 (N_2440,N_2316,N_2388);
nand U2441 (N_2441,N_2352,N_2208);
xor U2442 (N_2442,N_2245,N_2231);
nand U2443 (N_2443,N_2284,N_2247);
nor U2444 (N_2444,N_2275,N_2213);
xnor U2445 (N_2445,N_2281,N_2264);
or U2446 (N_2446,N_2347,N_2323);
nand U2447 (N_2447,N_2278,N_2290);
or U2448 (N_2448,N_2283,N_2301);
nor U2449 (N_2449,N_2293,N_2282);
or U2450 (N_2450,N_2342,N_2377);
nor U2451 (N_2451,N_2374,N_2297);
nor U2452 (N_2452,N_2383,N_2375);
and U2453 (N_2453,N_2358,N_2392);
and U2454 (N_2454,N_2337,N_2340);
nor U2455 (N_2455,N_2203,N_2209);
and U2456 (N_2456,N_2266,N_2210);
or U2457 (N_2457,N_2259,N_2286);
xor U2458 (N_2458,N_2291,N_2332);
nand U2459 (N_2459,N_2321,N_2390);
or U2460 (N_2460,N_2343,N_2289);
and U2461 (N_2461,N_2399,N_2379);
nor U2462 (N_2462,N_2229,N_2228);
or U2463 (N_2463,N_2345,N_2324);
nand U2464 (N_2464,N_2288,N_2364);
nor U2465 (N_2465,N_2249,N_2314);
nand U2466 (N_2466,N_2396,N_2263);
and U2467 (N_2467,N_2292,N_2349);
xnor U2468 (N_2468,N_2366,N_2326);
and U2469 (N_2469,N_2296,N_2211);
nor U2470 (N_2470,N_2306,N_2270);
or U2471 (N_2471,N_2202,N_2397);
nor U2472 (N_2472,N_2370,N_2398);
xnor U2473 (N_2473,N_2308,N_2232);
nand U2474 (N_2474,N_2239,N_2322);
xnor U2475 (N_2475,N_2244,N_2225);
xnor U2476 (N_2476,N_2224,N_2273);
xor U2477 (N_2477,N_2252,N_2330);
nand U2478 (N_2478,N_2218,N_2285);
nor U2479 (N_2479,N_2303,N_2373);
and U2480 (N_2480,N_2359,N_2302);
xor U2481 (N_2481,N_2274,N_2222);
nand U2482 (N_2482,N_2387,N_2269);
xnor U2483 (N_2483,N_2205,N_2329);
nor U2484 (N_2484,N_2255,N_2220);
xor U2485 (N_2485,N_2276,N_2395);
nor U2486 (N_2486,N_2238,N_2385);
nor U2487 (N_2487,N_2227,N_2206);
and U2488 (N_2488,N_2313,N_2336);
and U2489 (N_2489,N_2294,N_2348);
nand U2490 (N_2490,N_2391,N_2357);
or U2491 (N_2491,N_2200,N_2376);
nor U2492 (N_2492,N_2356,N_2260);
nand U2493 (N_2493,N_2298,N_2365);
nand U2494 (N_2494,N_2267,N_2325);
and U2495 (N_2495,N_2215,N_2310);
or U2496 (N_2496,N_2320,N_2394);
nor U2497 (N_2497,N_2214,N_2384);
xnor U2498 (N_2498,N_2341,N_2277);
and U2499 (N_2499,N_2305,N_2295);
or U2500 (N_2500,N_2255,N_2331);
xnor U2501 (N_2501,N_2386,N_2244);
xor U2502 (N_2502,N_2366,N_2271);
nor U2503 (N_2503,N_2292,N_2340);
and U2504 (N_2504,N_2279,N_2221);
or U2505 (N_2505,N_2227,N_2376);
or U2506 (N_2506,N_2217,N_2398);
nand U2507 (N_2507,N_2223,N_2215);
nand U2508 (N_2508,N_2329,N_2388);
or U2509 (N_2509,N_2385,N_2267);
xor U2510 (N_2510,N_2242,N_2206);
or U2511 (N_2511,N_2275,N_2367);
nand U2512 (N_2512,N_2239,N_2267);
xor U2513 (N_2513,N_2258,N_2391);
and U2514 (N_2514,N_2293,N_2387);
nor U2515 (N_2515,N_2327,N_2230);
nor U2516 (N_2516,N_2334,N_2365);
and U2517 (N_2517,N_2259,N_2387);
nor U2518 (N_2518,N_2266,N_2287);
xor U2519 (N_2519,N_2320,N_2304);
or U2520 (N_2520,N_2356,N_2214);
nor U2521 (N_2521,N_2237,N_2303);
nand U2522 (N_2522,N_2218,N_2214);
and U2523 (N_2523,N_2214,N_2370);
nand U2524 (N_2524,N_2329,N_2290);
and U2525 (N_2525,N_2366,N_2200);
nor U2526 (N_2526,N_2321,N_2359);
nand U2527 (N_2527,N_2303,N_2200);
xor U2528 (N_2528,N_2394,N_2283);
or U2529 (N_2529,N_2335,N_2385);
nand U2530 (N_2530,N_2304,N_2373);
nor U2531 (N_2531,N_2244,N_2363);
nand U2532 (N_2532,N_2290,N_2225);
nand U2533 (N_2533,N_2236,N_2285);
nand U2534 (N_2534,N_2292,N_2306);
nand U2535 (N_2535,N_2271,N_2214);
xor U2536 (N_2536,N_2317,N_2335);
xnor U2537 (N_2537,N_2204,N_2254);
and U2538 (N_2538,N_2291,N_2339);
nand U2539 (N_2539,N_2375,N_2395);
nor U2540 (N_2540,N_2298,N_2377);
nor U2541 (N_2541,N_2222,N_2361);
nor U2542 (N_2542,N_2217,N_2238);
and U2543 (N_2543,N_2373,N_2201);
nor U2544 (N_2544,N_2302,N_2237);
nor U2545 (N_2545,N_2266,N_2215);
xnor U2546 (N_2546,N_2301,N_2297);
nor U2547 (N_2547,N_2266,N_2399);
xnor U2548 (N_2548,N_2370,N_2333);
xnor U2549 (N_2549,N_2289,N_2258);
and U2550 (N_2550,N_2364,N_2334);
and U2551 (N_2551,N_2234,N_2277);
nand U2552 (N_2552,N_2317,N_2206);
and U2553 (N_2553,N_2377,N_2286);
xnor U2554 (N_2554,N_2267,N_2246);
nand U2555 (N_2555,N_2225,N_2275);
nand U2556 (N_2556,N_2289,N_2336);
and U2557 (N_2557,N_2385,N_2206);
nand U2558 (N_2558,N_2351,N_2349);
xnor U2559 (N_2559,N_2205,N_2313);
nand U2560 (N_2560,N_2359,N_2319);
xor U2561 (N_2561,N_2376,N_2237);
xor U2562 (N_2562,N_2313,N_2398);
nand U2563 (N_2563,N_2307,N_2254);
nand U2564 (N_2564,N_2247,N_2293);
or U2565 (N_2565,N_2250,N_2261);
or U2566 (N_2566,N_2306,N_2262);
or U2567 (N_2567,N_2346,N_2334);
nor U2568 (N_2568,N_2286,N_2378);
and U2569 (N_2569,N_2208,N_2389);
xnor U2570 (N_2570,N_2271,N_2303);
nand U2571 (N_2571,N_2368,N_2338);
and U2572 (N_2572,N_2244,N_2289);
and U2573 (N_2573,N_2376,N_2347);
xnor U2574 (N_2574,N_2216,N_2297);
nand U2575 (N_2575,N_2313,N_2233);
or U2576 (N_2576,N_2314,N_2251);
nor U2577 (N_2577,N_2359,N_2383);
xnor U2578 (N_2578,N_2231,N_2317);
nor U2579 (N_2579,N_2327,N_2354);
nor U2580 (N_2580,N_2389,N_2334);
and U2581 (N_2581,N_2341,N_2229);
nand U2582 (N_2582,N_2270,N_2350);
or U2583 (N_2583,N_2275,N_2383);
nand U2584 (N_2584,N_2282,N_2262);
or U2585 (N_2585,N_2252,N_2344);
and U2586 (N_2586,N_2290,N_2281);
or U2587 (N_2587,N_2259,N_2349);
and U2588 (N_2588,N_2335,N_2266);
xnor U2589 (N_2589,N_2207,N_2356);
xor U2590 (N_2590,N_2378,N_2344);
nand U2591 (N_2591,N_2357,N_2332);
or U2592 (N_2592,N_2230,N_2342);
nor U2593 (N_2593,N_2273,N_2334);
nor U2594 (N_2594,N_2337,N_2203);
xor U2595 (N_2595,N_2347,N_2334);
nor U2596 (N_2596,N_2219,N_2281);
xor U2597 (N_2597,N_2215,N_2331);
nor U2598 (N_2598,N_2304,N_2358);
or U2599 (N_2599,N_2281,N_2397);
and U2600 (N_2600,N_2476,N_2586);
or U2601 (N_2601,N_2520,N_2511);
nor U2602 (N_2602,N_2430,N_2594);
nand U2603 (N_2603,N_2436,N_2522);
nor U2604 (N_2604,N_2593,N_2585);
and U2605 (N_2605,N_2445,N_2518);
nand U2606 (N_2606,N_2563,N_2583);
and U2607 (N_2607,N_2587,N_2566);
nor U2608 (N_2608,N_2559,N_2442);
or U2609 (N_2609,N_2453,N_2550);
xnor U2610 (N_2610,N_2501,N_2406);
nand U2611 (N_2611,N_2508,N_2515);
nor U2612 (N_2612,N_2492,N_2537);
xnor U2613 (N_2613,N_2580,N_2578);
nand U2614 (N_2614,N_2534,N_2485);
nand U2615 (N_2615,N_2403,N_2452);
nand U2616 (N_2616,N_2405,N_2547);
xor U2617 (N_2617,N_2444,N_2551);
xor U2618 (N_2618,N_2472,N_2431);
xnor U2619 (N_2619,N_2419,N_2568);
xor U2620 (N_2620,N_2422,N_2465);
xor U2621 (N_2621,N_2443,N_2415);
nor U2622 (N_2622,N_2541,N_2425);
xor U2623 (N_2623,N_2408,N_2544);
nor U2624 (N_2624,N_2531,N_2486);
xor U2625 (N_2625,N_2592,N_2502);
xor U2626 (N_2626,N_2536,N_2451);
and U2627 (N_2627,N_2413,N_2423);
or U2628 (N_2628,N_2483,N_2416);
and U2629 (N_2629,N_2554,N_2523);
or U2630 (N_2630,N_2527,N_2482);
nand U2631 (N_2631,N_2595,N_2571);
nor U2632 (N_2632,N_2473,N_2506);
xnor U2633 (N_2633,N_2572,N_2456);
nor U2634 (N_2634,N_2454,N_2498);
or U2635 (N_2635,N_2589,N_2426);
xor U2636 (N_2636,N_2496,N_2464);
nand U2637 (N_2637,N_2468,N_2562);
nor U2638 (N_2638,N_2567,N_2548);
nand U2639 (N_2639,N_2446,N_2532);
xnor U2640 (N_2640,N_2424,N_2543);
nand U2641 (N_2641,N_2598,N_2525);
and U2642 (N_2642,N_2457,N_2478);
nor U2643 (N_2643,N_2521,N_2561);
and U2644 (N_2644,N_2558,N_2433);
and U2645 (N_2645,N_2462,N_2488);
nor U2646 (N_2646,N_2553,N_2517);
nor U2647 (N_2647,N_2491,N_2458);
nand U2648 (N_2648,N_2574,N_2440);
nand U2649 (N_2649,N_2509,N_2467);
xnor U2650 (N_2650,N_2557,N_2493);
or U2651 (N_2651,N_2516,N_2570);
nand U2652 (N_2652,N_2421,N_2577);
nand U2653 (N_2653,N_2432,N_2549);
and U2654 (N_2654,N_2539,N_2448);
or U2655 (N_2655,N_2576,N_2497);
nor U2656 (N_2656,N_2528,N_2489);
nand U2657 (N_2657,N_2530,N_2449);
and U2658 (N_2658,N_2490,N_2484);
or U2659 (N_2659,N_2579,N_2510);
nand U2660 (N_2660,N_2552,N_2569);
or U2661 (N_2661,N_2526,N_2519);
nor U2662 (N_2662,N_2418,N_2417);
and U2663 (N_2663,N_2581,N_2535);
or U2664 (N_2664,N_2400,N_2538);
nand U2665 (N_2665,N_2466,N_2463);
xor U2666 (N_2666,N_2540,N_2505);
nor U2667 (N_2667,N_2584,N_2599);
xnor U2668 (N_2668,N_2533,N_2582);
or U2669 (N_2669,N_2470,N_2503);
xor U2670 (N_2670,N_2471,N_2428);
xnor U2671 (N_2671,N_2500,N_2545);
and U2672 (N_2672,N_2409,N_2542);
or U2673 (N_2673,N_2439,N_2477);
nand U2674 (N_2674,N_2434,N_2479);
nand U2675 (N_2675,N_2474,N_2450);
xor U2676 (N_2676,N_2481,N_2514);
or U2677 (N_2677,N_2487,N_2407);
and U2678 (N_2678,N_2414,N_2564);
nor U2679 (N_2679,N_2460,N_2459);
or U2680 (N_2680,N_2495,N_2401);
nand U2681 (N_2681,N_2504,N_2427);
nand U2682 (N_2682,N_2475,N_2529);
nor U2683 (N_2683,N_2441,N_2597);
or U2684 (N_2684,N_2560,N_2447);
and U2685 (N_2685,N_2513,N_2524);
and U2686 (N_2686,N_2404,N_2591);
nor U2687 (N_2687,N_2494,N_2438);
nor U2688 (N_2688,N_2588,N_2410);
nor U2689 (N_2689,N_2402,N_2411);
nand U2690 (N_2690,N_2546,N_2420);
nor U2691 (N_2691,N_2556,N_2435);
or U2692 (N_2692,N_2555,N_2461);
xor U2693 (N_2693,N_2575,N_2590);
nor U2694 (N_2694,N_2499,N_2573);
xor U2695 (N_2695,N_2455,N_2437);
xor U2696 (N_2696,N_2429,N_2565);
xor U2697 (N_2697,N_2507,N_2469);
nand U2698 (N_2698,N_2512,N_2480);
and U2699 (N_2699,N_2596,N_2412);
nand U2700 (N_2700,N_2559,N_2542);
nand U2701 (N_2701,N_2415,N_2594);
and U2702 (N_2702,N_2442,N_2584);
or U2703 (N_2703,N_2462,N_2446);
nand U2704 (N_2704,N_2447,N_2578);
and U2705 (N_2705,N_2438,N_2543);
or U2706 (N_2706,N_2566,N_2474);
or U2707 (N_2707,N_2472,N_2539);
and U2708 (N_2708,N_2552,N_2535);
nor U2709 (N_2709,N_2431,N_2594);
or U2710 (N_2710,N_2495,N_2574);
nand U2711 (N_2711,N_2415,N_2589);
and U2712 (N_2712,N_2409,N_2521);
and U2713 (N_2713,N_2419,N_2597);
or U2714 (N_2714,N_2423,N_2481);
nand U2715 (N_2715,N_2507,N_2450);
nand U2716 (N_2716,N_2400,N_2550);
nor U2717 (N_2717,N_2404,N_2429);
or U2718 (N_2718,N_2549,N_2554);
nand U2719 (N_2719,N_2461,N_2463);
nand U2720 (N_2720,N_2570,N_2580);
and U2721 (N_2721,N_2402,N_2439);
or U2722 (N_2722,N_2528,N_2559);
or U2723 (N_2723,N_2478,N_2512);
nor U2724 (N_2724,N_2490,N_2553);
and U2725 (N_2725,N_2418,N_2477);
xor U2726 (N_2726,N_2575,N_2466);
and U2727 (N_2727,N_2528,N_2576);
and U2728 (N_2728,N_2532,N_2556);
nor U2729 (N_2729,N_2410,N_2539);
xnor U2730 (N_2730,N_2454,N_2441);
nor U2731 (N_2731,N_2461,N_2447);
nand U2732 (N_2732,N_2588,N_2521);
nor U2733 (N_2733,N_2580,N_2535);
and U2734 (N_2734,N_2485,N_2549);
xnor U2735 (N_2735,N_2563,N_2471);
or U2736 (N_2736,N_2407,N_2406);
or U2737 (N_2737,N_2542,N_2469);
nor U2738 (N_2738,N_2509,N_2479);
or U2739 (N_2739,N_2439,N_2475);
and U2740 (N_2740,N_2530,N_2521);
nor U2741 (N_2741,N_2529,N_2509);
nor U2742 (N_2742,N_2551,N_2487);
nor U2743 (N_2743,N_2505,N_2515);
xor U2744 (N_2744,N_2585,N_2594);
xnor U2745 (N_2745,N_2597,N_2573);
or U2746 (N_2746,N_2564,N_2543);
nand U2747 (N_2747,N_2584,N_2498);
nand U2748 (N_2748,N_2402,N_2479);
and U2749 (N_2749,N_2567,N_2551);
xor U2750 (N_2750,N_2471,N_2521);
nor U2751 (N_2751,N_2485,N_2420);
nand U2752 (N_2752,N_2413,N_2524);
nand U2753 (N_2753,N_2481,N_2529);
nand U2754 (N_2754,N_2592,N_2518);
nand U2755 (N_2755,N_2522,N_2417);
and U2756 (N_2756,N_2493,N_2558);
nand U2757 (N_2757,N_2582,N_2501);
nand U2758 (N_2758,N_2523,N_2431);
or U2759 (N_2759,N_2478,N_2532);
or U2760 (N_2760,N_2596,N_2458);
nor U2761 (N_2761,N_2552,N_2555);
and U2762 (N_2762,N_2402,N_2434);
and U2763 (N_2763,N_2501,N_2503);
nor U2764 (N_2764,N_2578,N_2511);
or U2765 (N_2765,N_2461,N_2526);
xnor U2766 (N_2766,N_2512,N_2418);
or U2767 (N_2767,N_2532,N_2597);
or U2768 (N_2768,N_2421,N_2563);
nor U2769 (N_2769,N_2434,N_2509);
nand U2770 (N_2770,N_2405,N_2458);
or U2771 (N_2771,N_2460,N_2550);
or U2772 (N_2772,N_2469,N_2572);
nand U2773 (N_2773,N_2577,N_2477);
nand U2774 (N_2774,N_2490,N_2434);
or U2775 (N_2775,N_2528,N_2598);
and U2776 (N_2776,N_2596,N_2459);
nand U2777 (N_2777,N_2563,N_2492);
and U2778 (N_2778,N_2412,N_2473);
nor U2779 (N_2779,N_2523,N_2560);
xnor U2780 (N_2780,N_2599,N_2401);
or U2781 (N_2781,N_2583,N_2518);
nor U2782 (N_2782,N_2443,N_2455);
xnor U2783 (N_2783,N_2593,N_2540);
nand U2784 (N_2784,N_2507,N_2513);
and U2785 (N_2785,N_2579,N_2436);
or U2786 (N_2786,N_2416,N_2581);
nand U2787 (N_2787,N_2549,N_2401);
nand U2788 (N_2788,N_2475,N_2544);
xor U2789 (N_2789,N_2471,N_2472);
nand U2790 (N_2790,N_2403,N_2440);
nand U2791 (N_2791,N_2472,N_2566);
and U2792 (N_2792,N_2480,N_2513);
and U2793 (N_2793,N_2553,N_2599);
and U2794 (N_2794,N_2485,N_2599);
nand U2795 (N_2795,N_2567,N_2534);
nor U2796 (N_2796,N_2432,N_2490);
nand U2797 (N_2797,N_2484,N_2437);
and U2798 (N_2798,N_2419,N_2474);
and U2799 (N_2799,N_2441,N_2549);
xor U2800 (N_2800,N_2619,N_2630);
and U2801 (N_2801,N_2755,N_2778);
nor U2802 (N_2802,N_2662,N_2753);
xor U2803 (N_2803,N_2668,N_2752);
or U2804 (N_2804,N_2603,N_2735);
and U2805 (N_2805,N_2697,N_2635);
and U2806 (N_2806,N_2645,N_2764);
nor U2807 (N_2807,N_2793,N_2669);
nand U2808 (N_2808,N_2714,N_2677);
nand U2809 (N_2809,N_2719,N_2736);
xnor U2810 (N_2810,N_2622,N_2798);
nor U2811 (N_2811,N_2713,N_2676);
nand U2812 (N_2812,N_2711,N_2791);
nor U2813 (N_2813,N_2650,N_2608);
xor U2814 (N_2814,N_2682,N_2756);
and U2815 (N_2815,N_2782,N_2656);
or U2816 (N_2816,N_2671,N_2691);
nor U2817 (N_2817,N_2685,N_2768);
xnor U2818 (N_2818,N_2642,N_2796);
nand U2819 (N_2819,N_2649,N_2655);
and U2820 (N_2820,N_2727,N_2770);
or U2821 (N_2821,N_2695,N_2661);
and U2822 (N_2822,N_2698,N_2627);
nand U2823 (N_2823,N_2767,N_2721);
nor U2824 (N_2824,N_2632,N_2785);
nor U2825 (N_2825,N_2734,N_2688);
and U2826 (N_2826,N_2724,N_2732);
xnor U2827 (N_2827,N_2747,N_2610);
xnor U2828 (N_2828,N_2605,N_2634);
nor U2829 (N_2829,N_2717,N_2667);
nor U2830 (N_2830,N_2620,N_2751);
nand U2831 (N_2831,N_2799,N_2703);
xnor U2832 (N_2832,N_2750,N_2616);
xnor U2833 (N_2833,N_2673,N_2766);
and U2834 (N_2834,N_2646,N_2797);
or U2835 (N_2835,N_2657,N_2777);
nand U2836 (N_2836,N_2612,N_2761);
and U2837 (N_2837,N_2749,N_2683);
or U2838 (N_2838,N_2771,N_2789);
xor U2839 (N_2839,N_2659,N_2660);
nand U2840 (N_2840,N_2737,N_2729);
nand U2841 (N_2841,N_2600,N_2638);
nand U2842 (N_2842,N_2607,N_2776);
nor U2843 (N_2843,N_2774,N_2718);
nand U2844 (N_2844,N_2788,N_2687);
and U2845 (N_2845,N_2786,N_2644);
or U2846 (N_2846,N_2733,N_2626);
and U2847 (N_2847,N_2614,N_2670);
nor U2848 (N_2848,N_2694,N_2762);
xnor U2849 (N_2849,N_2633,N_2666);
nor U2850 (N_2850,N_2617,N_2744);
xor U2851 (N_2851,N_2728,N_2672);
nor U2852 (N_2852,N_2730,N_2615);
nand U2853 (N_2853,N_2654,N_2702);
nor U2854 (N_2854,N_2725,N_2704);
xor U2855 (N_2855,N_2641,N_2613);
nand U2856 (N_2856,N_2705,N_2739);
nor U2857 (N_2857,N_2790,N_2763);
xnor U2858 (N_2858,N_2765,N_2696);
nand U2859 (N_2859,N_2611,N_2759);
nor U2860 (N_2860,N_2623,N_2674);
nand U2861 (N_2861,N_2621,N_2760);
or U2862 (N_2862,N_2625,N_2783);
xnor U2863 (N_2863,N_2680,N_2618);
nand U2864 (N_2864,N_2637,N_2708);
and U2865 (N_2865,N_2781,N_2664);
nor U2866 (N_2866,N_2710,N_2665);
and U2867 (N_2867,N_2743,N_2742);
nor U2868 (N_2868,N_2681,N_2731);
xor U2869 (N_2869,N_2720,N_2748);
and U2870 (N_2870,N_2746,N_2643);
and U2871 (N_2871,N_2772,N_2602);
or U2872 (N_2872,N_2658,N_2604);
xnor U2873 (N_2873,N_2723,N_2699);
xnor U2874 (N_2874,N_2693,N_2651);
nand U2875 (N_2875,N_2745,N_2787);
xor U2876 (N_2876,N_2754,N_2628);
nand U2877 (N_2877,N_2663,N_2684);
xnor U2878 (N_2878,N_2629,N_2701);
or U2879 (N_2879,N_2740,N_2709);
nand U2880 (N_2880,N_2601,N_2792);
and U2881 (N_2881,N_2773,N_2606);
nand U2882 (N_2882,N_2624,N_2689);
xnor U2883 (N_2883,N_2631,N_2675);
nand U2884 (N_2884,N_2715,N_2726);
nor U2885 (N_2885,N_2692,N_2648);
nand U2886 (N_2886,N_2757,N_2678);
and U2887 (N_2887,N_2775,N_2769);
xor U2888 (N_2888,N_2706,N_2647);
nand U2889 (N_2889,N_2758,N_2652);
and U2890 (N_2890,N_2700,N_2741);
nor U2891 (N_2891,N_2636,N_2738);
and U2892 (N_2892,N_2653,N_2679);
or U2893 (N_2893,N_2780,N_2609);
or U2894 (N_2894,N_2716,N_2784);
nor U2895 (N_2895,N_2639,N_2794);
nand U2896 (N_2896,N_2686,N_2707);
nor U2897 (N_2897,N_2795,N_2640);
and U2898 (N_2898,N_2690,N_2722);
xnor U2899 (N_2899,N_2779,N_2712);
and U2900 (N_2900,N_2726,N_2738);
and U2901 (N_2901,N_2767,N_2683);
xor U2902 (N_2902,N_2796,N_2614);
or U2903 (N_2903,N_2605,N_2698);
or U2904 (N_2904,N_2675,N_2735);
and U2905 (N_2905,N_2751,N_2750);
nand U2906 (N_2906,N_2654,N_2638);
and U2907 (N_2907,N_2631,N_2677);
or U2908 (N_2908,N_2670,N_2624);
and U2909 (N_2909,N_2684,N_2622);
nand U2910 (N_2910,N_2745,N_2619);
nor U2911 (N_2911,N_2757,N_2786);
xor U2912 (N_2912,N_2737,N_2680);
xnor U2913 (N_2913,N_2774,N_2715);
nor U2914 (N_2914,N_2717,N_2670);
and U2915 (N_2915,N_2771,N_2676);
nand U2916 (N_2916,N_2660,N_2797);
nor U2917 (N_2917,N_2704,N_2710);
nor U2918 (N_2918,N_2725,N_2716);
xor U2919 (N_2919,N_2636,N_2630);
xnor U2920 (N_2920,N_2773,N_2626);
or U2921 (N_2921,N_2643,N_2787);
nor U2922 (N_2922,N_2624,N_2765);
nor U2923 (N_2923,N_2732,N_2614);
nor U2924 (N_2924,N_2774,N_2641);
or U2925 (N_2925,N_2692,N_2736);
xor U2926 (N_2926,N_2795,N_2774);
or U2927 (N_2927,N_2688,N_2669);
nand U2928 (N_2928,N_2667,N_2709);
nor U2929 (N_2929,N_2741,N_2718);
nor U2930 (N_2930,N_2730,N_2638);
nand U2931 (N_2931,N_2732,N_2678);
or U2932 (N_2932,N_2753,N_2711);
xnor U2933 (N_2933,N_2622,N_2776);
nand U2934 (N_2934,N_2779,N_2658);
nand U2935 (N_2935,N_2698,N_2775);
and U2936 (N_2936,N_2676,N_2623);
xor U2937 (N_2937,N_2752,N_2717);
nand U2938 (N_2938,N_2627,N_2624);
and U2939 (N_2939,N_2617,N_2741);
nor U2940 (N_2940,N_2744,N_2709);
or U2941 (N_2941,N_2630,N_2673);
and U2942 (N_2942,N_2786,N_2694);
xor U2943 (N_2943,N_2714,N_2687);
nor U2944 (N_2944,N_2748,N_2677);
nor U2945 (N_2945,N_2689,N_2656);
nor U2946 (N_2946,N_2751,N_2747);
or U2947 (N_2947,N_2758,N_2704);
xor U2948 (N_2948,N_2772,N_2752);
or U2949 (N_2949,N_2694,N_2692);
and U2950 (N_2950,N_2649,N_2691);
nand U2951 (N_2951,N_2630,N_2754);
nand U2952 (N_2952,N_2717,N_2652);
and U2953 (N_2953,N_2774,N_2600);
and U2954 (N_2954,N_2772,N_2601);
or U2955 (N_2955,N_2617,N_2757);
or U2956 (N_2956,N_2620,N_2729);
and U2957 (N_2957,N_2696,N_2614);
or U2958 (N_2958,N_2663,N_2689);
nand U2959 (N_2959,N_2768,N_2790);
and U2960 (N_2960,N_2765,N_2671);
xor U2961 (N_2961,N_2784,N_2760);
and U2962 (N_2962,N_2725,N_2769);
nand U2963 (N_2963,N_2724,N_2643);
nor U2964 (N_2964,N_2747,N_2755);
nor U2965 (N_2965,N_2673,N_2763);
xnor U2966 (N_2966,N_2674,N_2621);
nand U2967 (N_2967,N_2622,N_2662);
xnor U2968 (N_2968,N_2694,N_2615);
xnor U2969 (N_2969,N_2626,N_2714);
nand U2970 (N_2970,N_2770,N_2655);
xor U2971 (N_2971,N_2698,N_2623);
nor U2972 (N_2972,N_2606,N_2781);
and U2973 (N_2973,N_2661,N_2737);
or U2974 (N_2974,N_2754,N_2682);
nor U2975 (N_2975,N_2675,N_2780);
and U2976 (N_2976,N_2778,N_2763);
or U2977 (N_2977,N_2683,N_2665);
xor U2978 (N_2978,N_2638,N_2781);
nor U2979 (N_2979,N_2724,N_2604);
nor U2980 (N_2980,N_2722,N_2742);
and U2981 (N_2981,N_2639,N_2700);
or U2982 (N_2982,N_2653,N_2739);
nor U2983 (N_2983,N_2705,N_2678);
or U2984 (N_2984,N_2707,N_2606);
nor U2985 (N_2985,N_2668,N_2751);
or U2986 (N_2986,N_2728,N_2762);
nand U2987 (N_2987,N_2770,N_2765);
nand U2988 (N_2988,N_2694,N_2674);
or U2989 (N_2989,N_2772,N_2637);
nand U2990 (N_2990,N_2690,N_2790);
or U2991 (N_2991,N_2625,N_2713);
nor U2992 (N_2992,N_2793,N_2773);
xor U2993 (N_2993,N_2799,N_2758);
nand U2994 (N_2994,N_2708,N_2711);
nor U2995 (N_2995,N_2605,N_2770);
and U2996 (N_2996,N_2658,N_2617);
nand U2997 (N_2997,N_2792,N_2636);
and U2998 (N_2998,N_2600,N_2736);
nand U2999 (N_2999,N_2708,N_2733);
nand U3000 (N_3000,N_2873,N_2804);
xnor U3001 (N_3001,N_2986,N_2836);
and U3002 (N_3002,N_2910,N_2980);
nand U3003 (N_3003,N_2975,N_2865);
nand U3004 (N_3004,N_2911,N_2897);
xor U3005 (N_3005,N_2818,N_2892);
and U3006 (N_3006,N_2838,N_2811);
or U3007 (N_3007,N_2983,N_2960);
or U3008 (N_3008,N_2958,N_2913);
nor U3009 (N_3009,N_2821,N_2823);
xor U3010 (N_3010,N_2809,N_2852);
nor U3011 (N_3011,N_2850,N_2909);
and U3012 (N_3012,N_2807,N_2893);
and U3013 (N_3013,N_2924,N_2976);
nand U3014 (N_3014,N_2982,N_2937);
or U3015 (N_3015,N_2946,N_2843);
nor U3016 (N_3016,N_2801,N_2888);
and U3017 (N_3017,N_2954,N_2845);
xnor U3018 (N_3018,N_2837,N_2844);
or U3019 (N_3019,N_2854,N_2941);
xnor U3020 (N_3020,N_2921,N_2882);
or U3021 (N_3021,N_2842,N_2816);
and U3022 (N_3022,N_2827,N_2808);
xnor U3023 (N_3023,N_2890,N_2952);
nand U3024 (N_3024,N_2832,N_2858);
nor U3025 (N_3025,N_2918,N_2814);
and U3026 (N_3026,N_2908,N_2919);
xnor U3027 (N_3027,N_2864,N_2889);
xnor U3028 (N_3028,N_2833,N_2805);
nor U3029 (N_3029,N_2934,N_2912);
nor U3030 (N_3030,N_2926,N_2933);
or U3031 (N_3031,N_2899,N_2974);
and U3032 (N_3032,N_2880,N_2964);
and U3033 (N_3033,N_2853,N_2851);
nor U3034 (N_3034,N_2922,N_2942);
nand U3035 (N_3035,N_2917,N_2957);
xor U3036 (N_3036,N_2884,N_2861);
nand U3037 (N_3037,N_2819,N_2802);
nand U3038 (N_3038,N_2841,N_2956);
or U3039 (N_3039,N_2969,N_2927);
or U3040 (N_3040,N_2966,N_2961);
or U3041 (N_3041,N_2992,N_2936);
xnor U3042 (N_3042,N_2869,N_2900);
nor U3043 (N_3043,N_2993,N_2995);
or U3044 (N_3044,N_2978,N_2943);
xnor U3045 (N_3045,N_2968,N_2876);
nor U3046 (N_3046,N_2829,N_2863);
xnor U3047 (N_3047,N_2839,N_2887);
nand U3048 (N_3048,N_2859,N_2870);
xnor U3049 (N_3049,N_2984,N_2951);
nand U3050 (N_3050,N_2903,N_2867);
nand U3051 (N_3051,N_2962,N_2938);
nand U3052 (N_3052,N_2813,N_2998);
and U3053 (N_3053,N_2860,N_2855);
xnor U3054 (N_3054,N_2895,N_2944);
xnor U3055 (N_3055,N_2848,N_2967);
xor U3056 (N_3056,N_2875,N_2945);
xor U3057 (N_3057,N_2886,N_2830);
or U3058 (N_3058,N_2906,N_2902);
xnor U3059 (N_3059,N_2925,N_2959);
nor U3060 (N_3060,N_2896,N_2815);
xor U3061 (N_3061,N_2988,N_2856);
xor U3062 (N_3062,N_2947,N_2999);
xnor U3063 (N_3063,N_2997,N_2935);
xnor U3064 (N_3064,N_2831,N_2868);
nand U3065 (N_3065,N_2916,N_2904);
or U3066 (N_3066,N_2872,N_2847);
xnor U3067 (N_3067,N_2972,N_2835);
nand U3068 (N_3068,N_2970,N_2826);
nor U3069 (N_3069,N_2883,N_2987);
or U3070 (N_3070,N_2866,N_2915);
nand U3071 (N_3071,N_2923,N_2828);
or U3072 (N_3072,N_2878,N_2973);
nor U3073 (N_3073,N_2898,N_2990);
and U3074 (N_3074,N_2820,N_2803);
or U3075 (N_3075,N_2939,N_2931);
xnor U3076 (N_3076,N_2981,N_2929);
nor U3077 (N_3077,N_2862,N_2971);
xnor U3078 (N_3078,N_2953,N_2930);
and U3079 (N_3079,N_2877,N_2879);
and U3080 (N_3080,N_2949,N_2928);
nand U3081 (N_3081,N_2846,N_2810);
nand U3082 (N_3082,N_2822,N_2963);
and U3083 (N_3083,N_2979,N_2991);
and U3084 (N_3084,N_2955,N_2874);
xnor U3085 (N_3085,N_2800,N_2905);
nand U3086 (N_3086,N_2825,N_2824);
and U3087 (N_3087,N_2940,N_2891);
nor U3088 (N_3088,N_2881,N_2834);
nor U3089 (N_3089,N_2901,N_2812);
or U3090 (N_3090,N_2977,N_2914);
or U3091 (N_3091,N_2871,N_2849);
nor U3092 (N_3092,N_2996,N_2932);
or U3093 (N_3093,N_2948,N_2806);
or U3094 (N_3094,N_2985,N_2994);
and U3095 (N_3095,N_2989,N_2885);
nand U3096 (N_3096,N_2817,N_2950);
or U3097 (N_3097,N_2965,N_2907);
nor U3098 (N_3098,N_2920,N_2840);
nor U3099 (N_3099,N_2857,N_2894);
or U3100 (N_3100,N_2890,N_2922);
or U3101 (N_3101,N_2904,N_2918);
xor U3102 (N_3102,N_2816,N_2844);
or U3103 (N_3103,N_2921,N_2990);
or U3104 (N_3104,N_2826,N_2927);
nand U3105 (N_3105,N_2922,N_2884);
nor U3106 (N_3106,N_2996,N_2839);
xor U3107 (N_3107,N_2841,N_2817);
nand U3108 (N_3108,N_2854,N_2981);
and U3109 (N_3109,N_2930,N_2878);
nor U3110 (N_3110,N_2964,N_2874);
or U3111 (N_3111,N_2853,N_2945);
nand U3112 (N_3112,N_2828,N_2867);
nand U3113 (N_3113,N_2857,N_2879);
and U3114 (N_3114,N_2985,N_2835);
xnor U3115 (N_3115,N_2841,N_2976);
nor U3116 (N_3116,N_2984,N_2846);
and U3117 (N_3117,N_2819,N_2964);
xnor U3118 (N_3118,N_2948,N_2906);
nor U3119 (N_3119,N_2899,N_2800);
xnor U3120 (N_3120,N_2998,N_2957);
or U3121 (N_3121,N_2983,N_2897);
xor U3122 (N_3122,N_2949,N_2883);
nor U3123 (N_3123,N_2965,N_2802);
and U3124 (N_3124,N_2988,N_2920);
nor U3125 (N_3125,N_2981,N_2905);
and U3126 (N_3126,N_2876,N_2804);
and U3127 (N_3127,N_2927,N_2878);
and U3128 (N_3128,N_2826,N_2896);
or U3129 (N_3129,N_2906,N_2970);
nor U3130 (N_3130,N_2866,N_2972);
and U3131 (N_3131,N_2972,N_2838);
or U3132 (N_3132,N_2952,N_2812);
nor U3133 (N_3133,N_2881,N_2886);
xnor U3134 (N_3134,N_2854,N_2964);
nand U3135 (N_3135,N_2898,N_2820);
nor U3136 (N_3136,N_2890,N_2959);
nand U3137 (N_3137,N_2992,N_2838);
or U3138 (N_3138,N_2824,N_2816);
nor U3139 (N_3139,N_2828,N_2898);
and U3140 (N_3140,N_2875,N_2909);
or U3141 (N_3141,N_2887,N_2842);
nor U3142 (N_3142,N_2933,N_2936);
and U3143 (N_3143,N_2893,N_2916);
nor U3144 (N_3144,N_2968,N_2987);
and U3145 (N_3145,N_2920,N_2962);
and U3146 (N_3146,N_2807,N_2802);
or U3147 (N_3147,N_2927,N_2916);
nor U3148 (N_3148,N_2902,N_2842);
and U3149 (N_3149,N_2944,N_2947);
nand U3150 (N_3150,N_2843,N_2830);
xnor U3151 (N_3151,N_2852,N_2885);
nand U3152 (N_3152,N_2808,N_2823);
and U3153 (N_3153,N_2875,N_2929);
and U3154 (N_3154,N_2824,N_2807);
nand U3155 (N_3155,N_2980,N_2815);
xor U3156 (N_3156,N_2910,N_2955);
xnor U3157 (N_3157,N_2971,N_2839);
nand U3158 (N_3158,N_2865,N_2886);
nor U3159 (N_3159,N_2823,N_2954);
or U3160 (N_3160,N_2958,N_2936);
or U3161 (N_3161,N_2984,N_2818);
nand U3162 (N_3162,N_2933,N_2957);
and U3163 (N_3163,N_2962,N_2926);
and U3164 (N_3164,N_2906,N_2810);
xnor U3165 (N_3165,N_2962,N_2833);
and U3166 (N_3166,N_2898,N_2977);
nor U3167 (N_3167,N_2883,N_2881);
nand U3168 (N_3168,N_2814,N_2878);
and U3169 (N_3169,N_2882,N_2841);
nor U3170 (N_3170,N_2875,N_2820);
and U3171 (N_3171,N_2874,N_2932);
and U3172 (N_3172,N_2846,N_2843);
nor U3173 (N_3173,N_2813,N_2960);
nand U3174 (N_3174,N_2825,N_2979);
or U3175 (N_3175,N_2976,N_2882);
or U3176 (N_3176,N_2934,N_2821);
or U3177 (N_3177,N_2868,N_2832);
or U3178 (N_3178,N_2897,N_2920);
nand U3179 (N_3179,N_2892,N_2850);
nor U3180 (N_3180,N_2934,N_2918);
nand U3181 (N_3181,N_2841,N_2975);
xor U3182 (N_3182,N_2965,N_2813);
nor U3183 (N_3183,N_2908,N_2986);
or U3184 (N_3184,N_2842,N_2863);
xnor U3185 (N_3185,N_2838,N_2951);
or U3186 (N_3186,N_2928,N_2868);
nand U3187 (N_3187,N_2876,N_2917);
nand U3188 (N_3188,N_2950,N_2863);
or U3189 (N_3189,N_2844,N_2918);
xor U3190 (N_3190,N_2830,N_2964);
nor U3191 (N_3191,N_2929,N_2853);
xor U3192 (N_3192,N_2855,N_2893);
nor U3193 (N_3193,N_2808,N_2804);
and U3194 (N_3194,N_2911,N_2848);
and U3195 (N_3195,N_2995,N_2967);
or U3196 (N_3196,N_2897,N_2828);
or U3197 (N_3197,N_2946,N_2955);
xnor U3198 (N_3198,N_2884,N_2900);
or U3199 (N_3199,N_2836,N_2901);
and U3200 (N_3200,N_3091,N_3000);
xor U3201 (N_3201,N_3033,N_3196);
and U3202 (N_3202,N_3011,N_3081);
and U3203 (N_3203,N_3045,N_3180);
nor U3204 (N_3204,N_3141,N_3082);
nand U3205 (N_3205,N_3042,N_3143);
xnor U3206 (N_3206,N_3068,N_3005);
nand U3207 (N_3207,N_3046,N_3020);
xor U3208 (N_3208,N_3099,N_3022);
nor U3209 (N_3209,N_3156,N_3173);
nor U3210 (N_3210,N_3182,N_3012);
nor U3211 (N_3211,N_3043,N_3199);
nand U3212 (N_3212,N_3014,N_3070);
or U3213 (N_3213,N_3017,N_3088);
nand U3214 (N_3214,N_3194,N_3096);
or U3215 (N_3215,N_3154,N_3047);
nand U3216 (N_3216,N_3061,N_3151);
and U3217 (N_3217,N_3031,N_3144);
and U3218 (N_3218,N_3197,N_3076);
nand U3219 (N_3219,N_3158,N_3095);
or U3220 (N_3220,N_3078,N_3146);
nand U3221 (N_3221,N_3170,N_3059);
xnor U3222 (N_3222,N_3009,N_3181);
and U3223 (N_3223,N_3121,N_3172);
xor U3224 (N_3224,N_3177,N_3161);
nor U3225 (N_3225,N_3030,N_3118);
or U3226 (N_3226,N_3124,N_3187);
and U3227 (N_3227,N_3114,N_3002);
nand U3228 (N_3228,N_3074,N_3108);
nand U3229 (N_3229,N_3038,N_3019);
and U3230 (N_3230,N_3063,N_3185);
nor U3231 (N_3231,N_3184,N_3062);
xor U3232 (N_3232,N_3175,N_3035);
nor U3233 (N_3233,N_3157,N_3129);
or U3234 (N_3234,N_3058,N_3135);
or U3235 (N_3235,N_3117,N_3119);
xnor U3236 (N_3236,N_3086,N_3127);
and U3237 (N_3237,N_3052,N_3125);
nand U3238 (N_3238,N_3178,N_3089);
or U3239 (N_3239,N_3136,N_3130);
nand U3240 (N_3240,N_3189,N_3164);
or U3241 (N_3241,N_3067,N_3128);
or U3242 (N_3242,N_3113,N_3137);
xnor U3243 (N_3243,N_3021,N_3015);
nand U3244 (N_3244,N_3040,N_3028);
nand U3245 (N_3245,N_3050,N_3131);
nand U3246 (N_3246,N_3049,N_3003);
xnor U3247 (N_3247,N_3153,N_3191);
nand U3248 (N_3248,N_3006,N_3132);
xor U3249 (N_3249,N_3065,N_3142);
or U3250 (N_3250,N_3071,N_3083);
nand U3251 (N_3251,N_3025,N_3183);
xnor U3252 (N_3252,N_3159,N_3123);
nor U3253 (N_3253,N_3167,N_3162);
nor U3254 (N_3254,N_3013,N_3079);
and U3255 (N_3255,N_3018,N_3171);
and U3256 (N_3256,N_3004,N_3106);
nand U3257 (N_3257,N_3111,N_3069);
and U3258 (N_3258,N_3105,N_3112);
or U3259 (N_3259,N_3055,N_3066);
or U3260 (N_3260,N_3016,N_3190);
and U3261 (N_3261,N_3192,N_3080);
and U3262 (N_3262,N_3057,N_3051);
nand U3263 (N_3263,N_3090,N_3149);
nand U3264 (N_3264,N_3155,N_3140);
nand U3265 (N_3265,N_3165,N_3126);
nand U3266 (N_3266,N_3103,N_3075);
nand U3267 (N_3267,N_3085,N_3195);
xor U3268 (N_3268,N_3168,N_3104);
and U3269 (N_3269,N_3060,N_3027);
nor U3270 (N_3270,N_3054,N_3102);
nor U3271 (N_3271,N_3109,N_3041);
and U3272 (N_3272,N_3024,N_3138);
xnor U3273 (N_3273,N_3039,N_3152);
xnor U3274 (N_3274,N_3147,N_3120);
xor U3275 (N_3275,N_3148,N_3163);
nor U3276 (N_3276,N_3139,N_3160);
xnor U3277 (N_3277,N_3026,N_3001);
nor U3278 (N_3278,N_3007,N_3092);
or U3279 (N_3279,N_3097,N_3198);
and U3280 (N_3280,N_3029,N_3032);
nand U3281 (N_3281,N_3150,N_3036);
nor U3282 (N_3282,N_3169,N_3166);
nand U3283 (N_3283,N_3115,N_3122);
nand U3284 (N_3284,N_3010,N_3186);
nor U3285 (N_3285,N_3101,N_3188);
nor U3286 (N_3286,N_3034,N_3193);
nand U3287 (N_3287,N_3087,N_3100);
xor U3288 (N_3288,N_3176,N_3179);
nor U3289 (N_3289,N_3044,N_3064);
and U3290 (N_3290,N_3174,N_3133);
xor U3291 (N_3291,N_3084,N_3053);
or U3292 (N_3292,N_3107,N_3077);
or U3293 (N_3293,N_3094,N_3056);
nor U3294 (N_3294,N_3116,N_3134);
nor U3295 (N_3295,N_3023,N_3037);
xnor U3296 (N_3296,N_3008,N_3110);
and U3297 (N_3297,N_3145,N_3048);
and U3298 (N_3298,N_3098,N_3073);
and U3299 (N_3299,N_3072,N_3093);
and U3300 (N_3300,N_3084,N_3043);
xor U3301 (N_3301,N_3047,N_3152);
and U3302 (N_3302,N_3174,N_3002);
nor U3303 (N_3303,N_3041,N_3090);
xnor U3304 (N_3304,N_3102,N_3055);
nand U3305 (N_3305,N_3132,N_3081);
or U3306 (N_3306,N_3064,N_3086);
nand U3307 (N_3307,N_3160,N_3014);
and U3308 (N_3308,N_3162,N_3043);
nand U3309 (N_3309,N_3113,N_3019);
or U3310 (N_3310,N_3144,N_3178);
or U3311 (N_3311,N_3038,N_3178);
xor U3312 (N_3312,N_3107,N_3190);
nand U3313 (N_3313,N_3116,N_3091);
nand U3314 (N_3314,N_3088,N_3195);
or U3315 (N_3315,N_3030,N_3136);
nor U3316 (N_3316,N_3046,N_3157);
nor U3317 (N_3317,N_3054,N_3179);
nand U3318 (N_3318,N_3182,N_3162);
and U3319 (N_3319,N_3074,N_3010);
xor U3320 (N_3320,N_3185,N_3057);
nand U3321 (N_3321,N_3013,N_3031);
nor U3322 (N_3322,N_3076,N_3048);
and U3323 (N_3323,N_3086,N_3152);
nor U3324 (N_3324,N_3071,N_3136);
or U3325 (N_3325,N_3032,N_3137);
nand U3326 (N_3326,N_3094,N_3147);
nand U3327 (N_3327,N_3060,N_3106);
xor U3328 (N_3328,N_3037,N_3035);
nand U3329 (N_3329,N_3104,N_3120);
nor U3330 (N_3330,N_3068,N_3021);
nand U3331 (N_3331,N_3157,N_3095);
nor U3332 (N_3332,N_3198,N_3148);
xor U3333 (N_3333,N_3103,N_3162);
or U3334 (N_3334,N_3117,N_3095);
nor U3335 (N_3335,N_3186,N_3132);
nand U3336 (N_3336,N_3136,N_3154);
xnor U3337 (N_3337,N_3195,N_3003);
nor U3338 (N_3338,N_3036,N_3103);
or U3339 (N_3339,N_3053,N_3014);
and U3340 (N_3340,N_3107,N_3146);
xor U3341 (N_3341,N_3047,N_3012);
nor U3342 (N_3342,N_3072,N_3082);
xnor U3343 (N_3343,N_3117,N_3033);
or U3344 (N_3344,N_3065,N_3043);
xnor U3345 (N_3345,N_3137,N_3097);
nand U3346 (N_3346,N_3017,N_3199);
nand U3347 (N_3347,N_3019,N_3049);
and U3348 (N_3348,N_3087,N_3139);
and U3349 (N_3349,N_3089,N_3015);
nor U3350 (N_3350,N_3084,N_3127);
nor U3351 (N_3351,N_3165,N_3023);
or U3352 (N_3352,N_3164,N_3001);
nor U3353 (N_3353,N_3068,N_3123);
nor U3354 (N_3354,N_3173,N_3057);
and U3355 (N_3355,N_3092,N_3138);
xor U3356 (N_3356,N_3091,N_3149);
nand U3357 (N_3357,N_3101,N_3113);
nand U3358 (N_3358,N_3128,N_3146);
nor U3359 (N_3359,N_3022,N_3081);
nand U3360 (N_3360,N_3068,N_3117);
nor U3361 (N_3361,N_3076,N_3036);
nor U3362 (N_3362,N_3092,N_3162);
or U3363 (N_3363,N_3119,N_3041);
and U3364 (N_3364,N_3037,N_3162);
nand U3365 (N_3365,N_3160,N_3064);
nand U3366 (N_3366,N_3063,N_3082);
or U3367 (N_3367,N_3085,N_3187);
nor U3368 (N_3368,N_3141,N_3073);
nor U3369 (N_3369,N_3096,N_3121);
nor U3370 (N_3370,N_3117,N_3078);
and U3371 (N_3371,N_3186,N_3045);
nand U3372 (N_3372,N_3060,N_3019);
xnor U3373 (N_3373,N_3082,N_3085);
or U3374 (N_3374,N_3052,N_3151);
nand U3375 (N_3375,N_3008,N_3017);
and U3376 (N_3376,N_3143,N_3178);
or U3377 (N_3377,N_3120,N_3054);
xor U3378 (N_3378,N_3160,N_3130);
or U3379 (N_3379,N_3075,N_3115);
or U3380 (N_3380,N_3097,N_3002);
nand U3381 (N_3381,N_3141,N_3109);
nand U3382 (N_3382,N_3059,N_3147);
and U3383 (N_3383,N_3165,N_3097);
and U3384 (N_3384,N_3192,N_3186);
nor U3385 (N_3385,N_3151,N_3141);
or U3386 (N_3386,N_3198,N_3092);
nor U3387 (N_3387,N_3154,N_3093);
xor U3388 (N_3388,N_3070,N_3131);
nand U3389 (N_3389,N_3131,N_3018);
nor U3390 (N_3390,N_3018,N_3103);
and U3391 (N_3391,N_3079,N_3035);
or U3392 (N_3392,N_3137,N_3030);
or U3393 (N_3393,N_3111,N_3015);
and U3394 (N_3394,N_3052,N_3157);
or U3395 (N_3395,N_3058,N_3169);
or U3396 (N_3396,N_3093,N_3132);
and U3397 (N_3397,N_3125,N_3153);
xor U3398 (N_3398,N_3036,N_3030);
nor U3399 (N_3399,N_3004,N_3035);
or U3400 (N_3400,N_3236,N_3209);
or U3401 (N_3401,N_3327,N_3311);
or U3402 (N_3402,N_3266,N_3337);
and U3403 (N_3403,N_3218,N_3282);
xor U3404 (N_3404,N_3344,N_3211);
nand U3405 (N_3405,N_3392,N_3376);
or U3406 (N_3406,N_3329,N_3326);
nand U3407 (N_3407,N_3271,N_3317);
and U3408 (N_3408,N_3339,N_3290);
and U3409 (N_3409,N_3221,N_3220);
nand U3410 (N_3410,N_3275,N_3368);
nand U3411 (N_3411,N_3255,N_3273);
xor U3412 (N_3412,N_3362,N_3371);
nor U3413 (N_3413,N_3281,N_3265);
xnor U3414 (N_3414,N_3309,N_3351);
xor U3415 (N_3415,N_3358,N_3380);
or U3416 (N_3416,N_3297,N_3389);
xnor U3417 (N_3417,N_3398,N_3205);
nand U3418 (N_3418,N_3335,N_3237);
xnor U3419 (N_3419,N_3269,N_3246);
or U3420 (N_3420,N_3330,N_3222);
xnor U3421 (N_3421,N_3391,N_3251);
xnor U3422 (N_3422,N_3373,N_3261);
xnor U3423 (N_3423,N_3388,N_3259);
nor U3424 (N_3424,N_3383,N_3206);
and U3425 (N_3425,N_3369,N_3258);
nor U3426 (N_3426,N_3232,N_3319);
and U3427 (N_3427,N_3316,N_3374);
xnor U3428 (N_3428,N_3382,N_3338);
xnor U3429 (N_3429,N_3253,N_3336);
nor U3430 (N_3430,N_3315,N_3288);
nor U3431 (N_3431,N_3280,N_3352);
nor U3432 (N_3432,N_3227,N_3390);
nand U3433 (N_3433,N_3360,N_3249);
or U3434 (N_3434,N_3277,N_3276);
nand U3435 (N_3435,N_3322,N_3379);
nand U3436 (N_3436,N_3370,N_3225);
xnor U3437 (N_3437,N_3292,N_3294);
xor U3438 (N_3438,N_3303,N_3248);
nand U3439 (N_3439,N_3289,N_3257);
xor U3440 (N_3440,N_3384,N_3264);
nand U3441 (N_3441,N_3325,N_3262);
nand U3442 (N_3442,N_3377,N_3238);
nand U3443 (N_3443,N_3279,N_3298);
nand U3444 (N_3444,N_3350,N_3313);
and U3445 (N_3445,N_3356,N_3354);
and U3446 (N_3446,N_3310,N_3302);
xnor U3447 (N_3447,N_3234,N_3372);
xnor U3448 (N_3448,N_3345,N_3348);
and U3449 (N_3449,N_3226,N_3363);
nand U3450 (N_3450,N_3361,N_3239);
xnor U3451 (N_3451,N_3375,N_3387);
nand U3452 (N_3452,N_3244,N_3340);
xor U3453 (N_3453,N_3252,N_3320);
xor U3454 (N_3454,N_3346,N_3342);
and U3455 (N_3455,N_3365,N_3216);
xor U3456 (N_3456,N_3268,N_3285);
nor U3457 (N_3457,N_3399,N_3355);
and U3458 (N_3458,N_3233,N_3343);
and U3459 (N_3459,N_3217,N_3299);
and U3460 (N_3460,N_3208,N_3386);
xor U3461 (N_3461,N_3334,N_3295);
nand U3462 (N_3462,N_3366,N_3204);
nor U3463 (N_3463,N_3229,N_3215);
nor U3464 (N_3464,N_3349,N_3283);
nand U3465 (N_3465,N_3260,N_3306);
nand U3466 (N_3466,N_3307,N_3367);
xnor U3467 (N_3467,N_3256,N_3224);
or U3468 (N_3468,N_3378,N_3245);
or U3469 (N_3469,N_3323,N_3263);
xnor U3470 (N_3470,N_3212,N_3254);
nor U3471 (N_3471,N_3270,N_3331);
or U3472 (N_3472,N_3223,N_3318);
or U3473 (N_3473,N_3296,N_3359);
nor U3474 (N_3474,N_3240,N_3304);
or U3475 (N_3475,N_3243,N_3287);
or U3476 (N_3476,N_3235,N_3291);
nor U3477 (N_3477,N_3202,N_3267);
xnor U3478 (N_3478,N_3333,N_3321);
and U3479 (N_3479,N_3328,N_3305);
nand U3480 (N_3480,N_3274,N_3397);
and U3481 (N_3481,N_3332,N_3213);
or U3482 (N_3482,N_3393,N_3381);
xnor U3483 (N_3483,N_3250,N_3353);
nand U3484 (N_3484,N_3278,N_3230);
or U3485 (N_3485,N_3200,N_3364);
xnor U3486 (N_3486,N_3247,N_3207);
or U3487 (N_3487,N_3272,N_3214);
xnor U3488 (N_3488,N_3341,N_3301);
nand U3489 (N_3489,N_3228,N_3300);
nor U3490 (N_3490,N_3357,N_3314);
nor U3491 (N_3491,N_3203,N_3231);
and U3492 (N_3492,N_3242,N_3241);
nor U3493 (N_3493,N_3308,N_3210);
or U3494 (N_3494,N_3201,N_3385);
or U3495 (N_3495,N_3324,N_3284);
xor U3496 (N_3496,N_3219,N_3286);
or U3497 (N_3497,N_3394,N_3396);
and U3498 (N_3498,N_3395,N_3347);
xnor U3499 (N_3499,N_3312,N_3293);
and U3500 (N_3500,N_3310,N_3226);
and U3501 (N_3501,N_3381,N_3355);
and U3502 (N_3502,N_3323,N_3348);
xor U3503 (N_3503,N_3356,N_3223);
or U3504 (N_3504,N_3302,N_3330);
or U3505 (N_3505,N_3337,N_3305);
and U3506 (N_3506,N_3342,N_3303);
nor U3507 (N_3507,N_3226,N_3372);
nand U3508 (N_3508,N_3265,N_3326);
nor U3509 (N_3509,N_3302,N_3306);
nand U3510 (N_3510,N_3385,N_3282);
nand U3511 (N_3511,N_3371,N_3230);
nor U3512 (N_3512,N_3364,N_3355);
or U3513 (N_3513,N_3241,N_3380);
nor U3514 (N_3514,N_3292,N_3230);
xnor U3515 (N_3515,N_3349,N_3384);
and U3516 (N_3516,N_3304,N_3356);
nor U3517 (N_3517,N_3321,N_3350);
nor U3518 (N_3518,N_3238,N_3296);
and U3519 (N_3519,N_3375,N_3294);
nand U3520 (N_3520,N_3243,N_3213);
xor U3521 (N_3521,N_3241,N_3308);
or U3522 (N_3522,N_3204,N_3334);
xnor U3523 (N_3523,N_3362,N_3338);
nor U3524 (N_3524,N_3272,N_3307);
xnor U3525 (N_3525,N_3325,N_3240);
and U3526 (N_3526,N_3212,N_3338);
nor U3527 (N_3527,N_3221,N_3308);
xor U3528 (N_3528,N_3336,N_3341);
nor U3529 (N_3529,N_3276,N_3367);
nor U3530 (N_3530,N_3397,N_3284);
nor U3531 (N_3531,N_3273,N_3337);
or U3532 (N_3532,N_3226,N_3340);
nand U3533 (N_3533,N_3280,N_3383);
and U3534 (N_3534,N_3341,N_3317);
nand U3535 (N_3535,N_3220,N_3203);
and U3536 (N_3536,N_3265,N_3214);
and U3537 (N_3537,N_3268,N_3397);
xor U3538 (N_3538,N_3298,N_3264);
xor U3539 (N_3539,N_3209,N_3382);
xnor U3540 (N_3540,N_3374,N_3340);
xnor U3541 (N_3541,N_3218,N_3265);
xor U3542 (N_3542,N_3224,N_3252);
nor U3543 (N_3543,N_3224,N_3319);
nand U3544 (N_3544,N_3278,N_3267);
nor U3545 (N_3545,N_3278,N_3242);
and U3546 (N_3546,N_3238,N_3282);
nand U3547 (N_3547,N_3259,N_3251);
or U3548 (N_3548,N_3398,N_3387);
or U3549 (N_3549,N_3216,N_3387);
and U3550 (N_3550,N_3368,N_3376);
and U3551 (N_3551,N_3306,N_3364);
or U3552 (N_3552,N_3334,N_3297);
and U3553 (N_3553,N_3303,N_3281);
and U3554 (N_3554,N_3317,N_3331);
and U3555 (N_3555,N_3259,N_3394);
nor U3556 (N_3556,N_3200,N_3368);
xnor U3557 (N_3557,N_3289,N_3380);
or U3558 (N_3558,N_3380,N_3268);
nor U3559 (N_3559,N_3271,N_3277);
or U3560 (N_3560,N_3218,N_3341);
and U3561 (N_3561,N_3382,N_3322);
xor U3562 (N_3562,N_3292,N_3269);
or U3563 (N_3563,N_3240,N_3268);
nand U3564 (N_3564,N_3240,N_3210);
and U3565 (N_3565,N_3300,N_3319);
and U3566 (N_3566,N_3323,N_3327);
or U3567 (N_3567,N_3234,N_3364);
nor U3568 (N_3568,N_3294,N_3327);
nand U3569 (N_3569,N_3228,N_3260);
or U3570 (N_3570,N_3309,N_3380);
nand U3571 (N_3571,N_3347,N_3381);
nand U3572 (N_3572,N_3256,N_3234);
and U3573 (N_3573,N_3343,N_3251);
or U3574 (N_3574,N_3380,N_3329);
and U3575 (N_3575,N_3329,N_3370);
nor U3576 (N_3576,N_3308,N_3370);
xor U3577 (N_3577,N_3260,N_3315);
or U3578 (N_3578,N_3223,N_3215);
and U3579 (N_3579,N_3323,N_3317);
xor U3580 (N_3580,N_3244,N_3389);
nor U3581 (N_3581,N_3309,N_3262);
and U3582 (N_3582,N_3240,N_3345);
xor U3583 (N_3583,N_3341,N_3262);
xnor U3584 (N_3584,N_3309,N_3269);
and U3585 (N_3585,N_3382,N_3339);
nand U3586 (N_3586,N_3207,N_3210);
and U3587 (N_3587,N_3361,N_3314);
and U3588 (N_3588,N_3247,N_3343);
or U3589 (N_3589,N_3275,N_3379);
nor U3590 (N_3590,N_3271,N_3387);
or U3591 (N_3591,N_3337,N_3317);
and U3592 (N_3592,N_3261,N_3262);
and U3593 (N_3593,N_3304,N_3336);
and U3594 (N_3594,N_3312,N_3274);
or U3595 (N_3595,N_3321,N_3316);
or U3596 (N_3596,N_3224,N_3383);
or U3597 (N_3597,N_3203,N_3317);
or U3598 (N_3598,N_3249,N_3264);
xor U3599 (N_3599,N_3242,N_3382);
xnor U3600 (N_3600,N_3526,N_3534);
nor U3601 (N_3601,N_3429,N_3483);
and U3602 (N_3602,N_3578,N_3589);
xor U3603 (N_3603,N_3508,N_3458);
xnor U3604 (N_3604,N_3535,N_3528);
and U3605 (N_3605,N_3465,N_3512);
nand U3606 (N_3606,N_3435,N_3489);
and U3607 (N_3607,N_3511,N_3568);
nor U3608 (N_3608,N_3538,N_3434);
or U3609 (N_3609,N_3407,N_3466);
or U3610 (N_3610,N_3586,N_3510);
xor U3611 (N_3611,N_3427,N_3420);
and U3612 (N_3612,N_3468,N_3591);
nor U3613 (N_3613,N_3577,N_3492);
nor U3614 (N_3614,N_3562,N_3452);
and U3615 (N_3615,N_3515,N_3462);
or U3616 (N_3616,N_3597,N_3503);
and U3617 (N_3617,N_3487,N_3472);
nand U3618 (N_3618,N_3495,N_3422);
nand U3619 (N_3619,N_3554,N_3410);
xnor U3620 (N_3620,N_3556,N_3533);
nand U3621 (N_3621,N_3445,N_3469);
or U3622 (N_3622,N_3550,N_3502);
xor U3623 (N_3623,N_3457,N_3572);
xnor U3624 (N_3624,N_3497,N_3529);
nor U3625 (N_3625,N_3588,N_3546);
xor U3626 (N_3626,N_3401,N_3485);
xor U3627 (N_3627,N_3573,N_3426);
nor U3628 (N_3628,N_3455,N_3412);
or U3629 (N_3629,N_3408,N_3431);
xor U3630 (N_3630,N_3405,N_3579);
nand U3631 (N_3631,N_3415,N_3481);
nor U3632 (N_3632,N_3490,N_3482);
and U3633 (N_3633,N_3500,N_3553);
and U3634 (N_3634,N_3473,N_3599);
nand U3635 (N_3635,N_3517,N_3499);
or U3636 (N_3636,N_3551,N_3594);
nand U3637 (N_3637,N_3513,N_3461);
nor U3638 (N_3638,N_3560,N_3456);
and U3639 (N_3639,N_3527,N_3436);
nor U3640 (N_3640,N_3575,N_3574);
nand U3641 (N_3641,N_3537,N_3491);
or U3642 (N_3642,N_3438,N_3516);
or U3643 (N_3643,N_3581,N_3571);
nand U3644 (N_3644,N_3549,N_3479);
xnor U3645 (N_3645,N_3403,N_3564);
and U3646 (N_3646,N_3530,N_3449);
nand U3647 (N_3647,N_3584,N_3505);
or U3648 (N_3648,N_3598,N_3402);
xor U3649 (N_3649,N_3476,N_3518);
or U3650 (N_3650,N_3506,N_3411);
nand U3651 (N_3651,N_3557,N_3444);
nor U3652 (N_3652,N_3555,N_3488);
nor U3653 (N_3653,N_3443,N_3437);
nor U3654 (N_3654,N_3563,N_3541);
or U3655 (N_3655,N_3442,N_3467);
xor U3656 (N_3656,N_3484,N_3587);
or U3657 (N_3657,N_3561,N_3433);
and U3658 (N_3658,N_3544,N_3486);
nor U3659 (N_3659,N_3520,N_3448);
nand U3660 (N_3660,N_3414,N_3539);
or U3661 (N_3661,N_3507,N_3471);
nor U3662 (N_3662,N_3514,N_3524);
and U3663 (N_3663,N_3593,N_3566);
or U3664 (N_3664,N_3480,N_3425);
or U3665 (N_3665,N_3441,N_3417);
or U3666 (N_3666,N_3558,N_3447);
nor U3667 (N_3667,N_3428,N_3446);
nand U3668 (N_3668,N_3523,N_3547);
and U3669 (N_3669,N_3543,N_3404);
xnor U3670 (N_3670,N_3583,N_3525);
nand U3671 (N_3671,N_3570,N_3423);
xor U3672 (N_3672,N_3406,N_3400);
and U3673 (N_3673,N_3464,N_3440);
nand U3674 (N_3674,N_3450,N_3585);
or U3675 (N_3675,N_3536,N_3545);
and U3676 (N_3676,N_3498,N_3418);
or U3677 (N_3677,N_3475,N_3565);
nand U3678 (N_3678,N_3567,N_3552);
nor U3679 (N_3679,N_3532,N_3504);
nand U3680 (N_3680,N_3595,N_3592);
nand U3681 (N_3681,N_3590,N_3470);
or U3682 (N_3682,N_3451,N_3531);
and U3683 (N_3683,N_3453,N_3459);
nor U3684 (N_3684,N_3460,N_3519);
nor U3685 (N_3685,N_3494,N_3569);
and U3686 (N_3686,N_3439,N_3559);
or U3687 (N_3687,N_3474,N_3496);
nor U3688 (N_3688,N_3542,N_3493);
or U3689 (N_3689,N_3582,N_3596);
and U3690 (N_3690,N_3409,N_3501);
xnor U3691 (N_3691,N_3580,N_3430);
or U3692 (N_3692,N_3509,N_3463);
nor U3693 (N_3693,N_3432,N_3421);
xor U3694 (N_3694,N_3478,N_3416);
nor U3695 (N_3695,N_3419,N_3477);
or U3696 (N_3696,N_3548,N_3454);
nand U3697 (N_3697,N_3413,N_3540);
nor U3698 (N_3698,N_3521,N_3424);
nand U3699 (N_3699,N_3522,N_3576);
or U3700 (N_3700,N_3520,N_3464);
and U3701 (N_3701,N_3593,N_3554);
or U3702 (N_3702,N_3489,N_3424);
and U3703 (N_3703,N_3583,N_3537);
or U3704 (N_3704,N_3460,N_3456);
or U3705 (N_3705,N_3506,N_3474);
nand U3706 (N_3706,N_3415,N_3486);
nor U3707 (N_3707,N_3598,N_3568);
xor U3708 (N_3708,N_3524,N_3504);
and U3709 (N_3709,N_3468,N_3501);
or U3710 (N_3710,N_3465,N_3529);
nor U3711 (N_3711,N_3444,N_3544);
and U3712 (N_3712,N_3497,N_3560);
or U3713 (N_3713,N_3432,N_3560);
xnor U3714 (N_3714,N_3509,N_3473);
nor U3715 (N_3715,N_3465,N_3574);
nor U3716 (N_3716,N_3446,N_3457);
and U3717 (N_3717,N_3549,N_3474);
xor U3718 (N_3718,N_3560,N_3450);
and U3719 (N_3719,N_3432,N_3514);
nand U3720 (N_3720,N_3441,N_3460);
xor U3721 (N_3721,N_3489,N_3447);
nor U3722 (N_3722,N_3545,N_3546);
nand U3723 (N_3723,N_3506,N_3465);
and U3724 (N_3724,N_3527,N_3438);
nor U3725 (N_3725,N_3535,N_3445);
or U3726 (N_3726,N_3489,N_3590);
nor U3727 (N_3727,N_3407,N_3463);
nor U3728 (N_3728,N_3450,N_3477);
and U3729 (N_3729,N_3470,N_3519);
and U3730 (N_3730,N_3414,N_3555);
nand U3731 (N_3731,N_3465,N_3492);
nand U3732 (N_3732,N_3458,N_3592);
and U3733 (N_3733,N_3576,N_3571);
nand U3734 (N_3734,N_3411,N_3448);
nor U3735 (N_3735,N_3439,N_3490);
or U3736 (N_3736,N_3488,N_3539);
xnor U3737 (N_3737,N_3539,N_3530);
xnor U3738 (N_3738,N_3476,N_3455);
nor U3739 (N_3739,N_3598,N_3470);
xor U3740 (N_3740,N_3413,N_3414);
nand U3741 (N_3741,N_3483,N_3596);
xor U3742 (N_3742,N_3595,N_3447);
nor U3743 (N_3743,N_3498,N_3485);
and U3744 (N_3744,N_3411,N_3525);
and U3745 (N_3745,N_3501,N_3450);
or U3746 (N_3746,N_3561,N_3502);
and U3747 (N_3747,N_3571,N_3408);
or U3748 (N_3748,N_3472,N_3450);
or U3749 (N_3749,N_3496,N_3463);
or U3750 (N_3750,N_3546,N_3450);
nand U3751 (N_3751,N_3538,N_3548);
and U3752 (N_3752,N_3501,N_3504);
nand U3753 (N_3753,N_3435,N_3503);
or U3754 (N_3754,N_3484,N_3501);
or U3755 (N_3755,N_3439,N_3516);
nand U3756 (N_3756,N_3505,N_3487);
nand U3757 (N_3757,N_3447,N_3594);
or U3758 (N_3758,N_3596,N_3438);
and U3759 (N_3759,N_3540,N_3404);
nor U3760 (N_3760,N_3569,N_3506);
nand U3761 (N_3761,N_3595,N_3502);
or U3762 (N_3762,N_3507,N_3599);
nand U3763 (N_3763,N_3469,N_3487);
nor U3764 (N_3764,N_3508,N_3534);
xor U3765 (N_3765,N_3487,N_3530);
or U3766 (N_3766,N_3477,N_3414);
and U3767 (N_3767,N_3509,N_3435);
nand U3768 (N_3768,N_3461,N_3501);
and U3769 (N_3769,N_3423,N_3499);
or U3770 (N_3770,N_3504,N_3459);
nand U3771 (N_3771,N_3447,N_3544);
and U3772 (N_3772,N_3404,N_3499);
or U3773 (N_3773,N_3451,N_3507);
nand U3774 (N_3774,N_3432,N_3516);
nor U3775 (N_3775,N_3554,N_3451);
nand U3776 (N_3776,N_3520,N_3408);
xnor U3777 (N_3777,N_3513,N_3475);
nand U3778 (N_3778,N_3418,N_3429);
or U3779 (N_3779,N_3573,N_3541);
nand U3780 (N_3780,N_3544,N_3527);
and U3781 (N_3781,N_3464,N_3408);
nor U3782 (N_3782,N_3400,N_3595);
xnor U3783 (N_3783,N_3511,N_3545);
or U3784 (N_3784,N_3406,N_3558);
or U3785 (N_3785,N_3449,N_3501);
and U3786 (N_3786,N_3424,N_3488);
nand U3787 (N_3787,N_3591,N_3595);
xor U3788 (N_3788,N_3436,N_3430);
nand U3789 (N_3789,N_3599,N_3424);
xnor U3790 (N_3790,N_3541,N_3453);
xor U3791 (N_3791,N_3576,N_3451);
and U3792 (N_3792,N_3463,N_3440);
nor U3793 (N_3793,N_3565,N_3491);
nor U3794 (N_3794,N_3537,N_3421);
nand U3795 (N_3795,N_3426,N_3455);
nand U3796 (N_3796,N_3500,N_3505);
and U3797 (N_3797,N_3404,N_3596);
nor U3798 (N_3798,N_3448,N_3542);
nand U3799 (N_3799,N_3531,N_3410);
nor U3800 (N_3800,N_3654,N_3697);
xnor U3801 (N_3801,N_3724,N_3776);
nand U3802 (N_3802,N_3646,N_3717);
nor U3803 (N_3803,N_3659,N_3752);
nor U3804 (N_3804,N_3634,N_3772);
or U3805 (N_3805,N_3608,N_3718);
nor U3806 (N_3806,N_3710,N_3685);
nor U3807 (N_3807,N_3709,N_3641);
nor U3808 (N_3808,N_3622,N_3680);
nor U3809 (N_3809,N_3773,N_3765);
xnor U3810 (N_3810,N_3693,N_3715);
nor U3811 (N_3811,N_3667,N_3785);
or U3812 (N_3812,N_3643,N_3676);
and U3813 (N_3813,N_3739,N_3742);
nor U3814 (N_3814,N_3781,N_3611);
nor U3815 (N_3815,N_3777,N_3764);
xnor U3816 (N_3816,N_3758,N_3789);
and U3817 (N_3817,N_3616,N_3651);
or U3818 (N_3818,N_3795,N_3649);
or U3819 (N_3819,N_3759,N_3627);
nor U3820 (N_3820,N_3652,N_3656);
and U3821 (N_3821,N_3658,N_3686);
nand U3822 (N_3822,N_3607,N_3762);
nor U3823 (N_3823,N_3691,N_3712);
nor U3824 (N_3824,N_3760,N_3769);
and U3825 (N_3825,N_3730,N_3791);
nor U3826 (N_3826,N_3696,N_3601);
nor U3827 (N_3827,N_3726,N_3683);
nand U3828 (N_3828,N_3783,N_3745);
nand U3829 (N_3829,N_3630,N_3719);
nand U3830 (N_3830,N_3723,N_3653);
xor U3831 (N_3831,N_3665,N_3631);
and U3832 (N_3832,N_3728,N_3740);
and U3833 (N_3833,N_3793,N_3792);
nor U3834 (N_3834,N_3736,N_3695);
and U3835 (N_3835,N_3700,N_3675);
nor U3836 (N_3836,N_3731,N_3734);
nor U3837 (N_3837,N_3711,N_3716);
or U3838 (N_3838,N_3604,N_3722);
or U3839 (N_3839,N_3771,N_3755);
xnor U3840 (N_3840,N_3778,N_3632);
and U3841 (N_3841,N_3637,N_3682);
nand U3842 (N_3842,N_3624,N_3703);
and U3843 (N_3843,N_3798,N_3708);
nand U3844 (N_3844,N_3636,N_3662);
nor U3845 (N_3845,N_3784,N_3678);
xnor U3846 (N_3846,N_3725,N_3689);
nor U3847 (N_3847,N_3629,N_3625);
xnor U3848 (N_3848,N_3747,N_3767);
nand U3849 (N_3849,N_3699,N_3770);
and U3850 (N_3850,N_3757,N_3744);
nand U3851 (N_3851,N_3602,N_3600);
or U3852 (N_3852,N_3790,N_3645);
and U3853 (N_3853,N_3797,N_3753);
nand U3854 (N_3854,N_3763,N_3706);
xor U3855 (N_3855,N_3690,N_3729);
xnor U3856 (N_3856,N_3794,N_3603);
nor U3857 (N_3857,N_3743,N_3639);
nor U3858 (N_3858,N_3628,N_3749);
nand U3859 (N_3859,N_3782,N_3768);
nor U3860 (N_3860,N_3766,N_3774);
nor U3861 (N_3861,N_3638,N_3732);
nand U3862 (N_3862,N_3650,N_3666);
or U3863 (N_3863,N_3787,N_3664);
or U3864 (N_3864,N_3704,N_3672);
nand U3865 (N_3865,N_3721,N_3621);
xnor U3866 (N_3866,N_3761,N_3779);
or U3867 (N_3867,N_3614,N_3741);
nand U3868 (N_3868,N_3605,N_3788);
nand U3869 (N_3869,N_3799,N_3633);
nand U3870 (N_3870,N_3620,N_3688);
nor U3871 (N_3871,N_3705,N_3619);
xnor U3872 (N_3872,N_3610,N_3780);
and U3873 (N_3873,N_3617,N_3727);
nor U3874 (N_3874,N_3671,N_3796);
nor U3875 (N_3875,N_3684,N_3702);
nand U3876 (N_3876,N_3692,N_3668);
nor U3877 (N_3877,N_3775,N_3648);
and U3878 (N_3878,N_3661,N_3615);
xor U3879 (N_3879,N_3609,N_3612);
or U3880 (N_3880,N_3751,N_3663);
and U3881 (N_3881,N_3679,N_3714);
nand U3882 (N_3882,N_3642,N_3618);
and U3883 (N_3883,N_3786,N_3681);
xor U3884 (N_3884,N_3657,N_3655);
nor U3885 (N_3885,N_3737,N_3707);
nand U3886 (N_3886,N_3750,N_3674);
or U3887 (N_3887,N_3746,N_3647);
nor U3888 (N_3888,N_3694,N_3623);
or U3889 (N_3889,N_3626,N_3606);
and U3890 (N_3890,N_3613,N_3733);
or U3891 (N_3891,N_3720,N_3660);
nor U3892 (N_3892,N_3687,N_3669);
or U3893 (N_3893,N_3677,N_3748);
or U3894 (N_3894,N_3644,N_3701);
or U3895 (N_3895,N_3754,N_3735);
nor U3896 (N_3896,N_3756,N_3640);
xor U3897 (N_3897,N_3673,N_3713);
and U3898 (N_3898,N_3635,N_3738);
or U3899 (N_3899,N_3670,N_3698);
nor U3900 (N_3900,N_3674,N_3620);
or U3901 (N_3901,N_3758,N_3694);
nand U3902 (N_3902,N_3686,N_3797);
xor U3903 (N_3903,N_3758,N_3601);
xnor U3904 (N_3904,N_3663,N_3632);
xnor U3905 (N_3905,N_3664,N_3629);
nand U3906 (N_3906,N_3719,N_3789);
xor U3907 (N_3907,N_3785,N_3665);
or U3908 (N_3908,N_3647,N_3739);
or U3909 (N_3909,N_3718,N_3755);
or U3910 (N_3910,N_3657,N_3703);
nand U3911 (N_3911,N_3773,N_3740);
or U3912 (N_3912,N_3665,N_3745);
nor U3913 (N_3913,N_3690,N_3760);
nand U3914 (N_3914,N_3720,N_3623);
nand U3915 (N_3915,N_3727,N_3676);
nor U3916 (N_3916,N_3637,N_3771);
and U3917 (N_3917,N_3775,N_3633);
xor U3918 (N_3918,N_3710,N_3639);
or U3919 (N_3919,N_3719,N_3724);
nand U3920 (N_3920,N_3624,N_3778);
xnor U3921 (N_3921,N_3758,N_3620);
xor U3922 (N_3922,N_3797,N_3664);
xnor U3923 (N_3923,N_3719,N_3686);
or U3924 (N_3924,N_3659,N_3698);
nor U3925 (N_3925,N_3727,N_3609);
nor U3926 (N_3926,N_3623,N_3672);
xor U3927 (N_3927,N_3612,N_3750);
xnor U3928 (N_3928,N_3615,N_3744);
nand U3929 (N_3929,N_3750,N_3638);
nand U3930 (N_3930,N_3685,N_3761);
nand U3931 (N_3931,N_3659,N_3681);
nand U3932 (N_3932,N_3671,N_3602);
nor U3933 (N_3933,N_3708,N_3748);
and U3934 (N_3934,N_3761,N_3755);
nor U3935 (N_3935,N_3741,N_3798);
xnor U3936 (N_3936,N_3751,N_3633);
and U3937 (N_3937,N_3774,N_3784);
xnor U3938 (N_3938,N_3781,N_3642);
nor U3939 (N_3939,N_3716,N_3649);
xnor U3940 (N_3940,N_3612,N_3725);
xor U3941 (N_3941,N_3732,N_3761);
nand U3942 (N_3942,N_3764,N_3771);
and U3943 (N_3943,N_3750,N_3722);
xor U3944 (N_3944,N_3746,N_3623);
and U3945 (N_3945,N_3730,N_3690);
xor U3946 (N_3946,N_3708,N_3797);
and U3947 (N_3947,N_3665,N_3661);
or U3948 (N_3948,N_3628,N_3662);
nand U3949 (N_3949,N_3682,N_3745);
nand U3950 (N_3950,N_3780,N_3793);
and U3951 (N_3951,N_3772,N_3648);
nand U3952 (N_3952,N_3613,N_3674);
nor U3953 (N_3953,N_3797,N_3671);
nand U3954 (N_3954,N_3648,N_3758);
nand U3955 (N_3955,N_3733,N_3626);
and U3956 (N_3956,N_3687,N_3780);
nor U3957 (N_3957,N_3760,N_3684);
xnor U3958 (N_3958,N_3732,N_3767);
or U3959 (N_3959,N_3640,N_3790);
xnor U3960 (N_3960,N_3698,N_3682);
nand U3961 (N_3961,N_3676,N_3699);
nor U3962 (N_3962,N_3752,N_3777);
nor U3963 (N_3963,N_3742,N_3718);
and U3964 (N_3964,N_3688,N_3736);
or U3965 (N_3965,N_3600,N_3776);
nand U3966 (N_3966,N_3716,N_3690);
xnor U3967 (N_3967,N_3774,N_3699);
nor U3968 (N_3968,N_3672,N_3740);
xnor U3969 (N_3969,N_3612,N_3604);
xnor U3970 (N_3970,N_3729,N_3737);
nand U3971 (N_3971,N_3760,N_3730);
and U3972 (N_3972,N_3606,N_3725);
nor U3973 (N_3973,N_3692,N_3610);
and U3974 (N_3974,N_3615,N_3642);
or U3975 (N_3975,N_3769,N_3652);
xnor U3976 (N_3976,N_3746,N_3763);
or U3977 (N_3977,N_3760,N_3669);
or U3978 (N_3978,N_3623,N_3631);
and U3979 (N_3979,N_3765,N_3771);
or U3980 (N_3980,N_3787,N_3728);
and U3981 (N_3981,N_3634,N_3762);
or U3982 (N_3982,N_3705,N_3645);
and U3983 (N_3983,N_3618,N_3733);
nand U3984 (N_3984,N_3765,N_3644);
or U3985 (N_3985,N_3753,N_3708);
and U3986 (N_3986,N_3796,N_3659);
xor U3987 (N_3987,N_3655,N_3679);
xnor U3988 (N_3988,N_3770,N_3661);
or U3989 (N_3989,N_3715,N_3753);
and U3990 (N_3990,N_3711,N_3725);
or U3991 (N_3991,N_3774,N_3739);
nand U3992 (N_3992,N_3763,N_3748);
nor U3993 (N_3993,N_3629,N_3681);
xnor U3994 (N_3994,N_3695,N_3656);
xnor U3995 (N_3995,N_3729,N_3749);
nor U3996 (N_3996,N_3607,N_3677);
and U3997 (N_3997,N_3730,N_3784);
nand U3998 (N_3998,N_3748,N_3633);
nor U3999 (N_3999,N_3702,N_3687);
xor U4000 (N_4000,N_3822,N_3944);
nand U4001 (N_4001,N_3957,N_3945);
nor U4002 (N_4002,N_3948,N_3804);
nand U4003 (N_4003,N_3995,N_3835);
and U4004 (N_4004,N_3908,N_3926);
and U4005 (N_4005,N_3832,N_3994);
nand U4006 (N_4006,N_3865,N_3953);
nand U4007 (N_4007,N_3837,N_3936);
or U4008 (N_4008,N_3928,N_3918);
xnor U4009 (N_4009,N_3911,N_3902);
and U4010 (N_4010,N_3987,N_3849);
xnor U4011 (N_4011,N_3990,N_3819);
and U4012 (N_4012,N_3874,N_3909);
and U4013 (N_4013,N_3973,N_3862);
and U4014 (N_4014,N_3806,N_3976);
or U4015 (N_4015,N_3814,N_3888);
nand U4016 (N_4016,N_3823,N_3979);
or U4017 (N_4017,N_3892,N_3811);
nand U4018 (N_4018,N_3815,N_3839);
nor U4019 (N_4019,N_3840,N_3986);
nand U4020 (N_4020,N_3877,N_3807);
and U4021 (N_4021,N_3803,N_3962);
nand U4022 (N_4022,N_3989,N_3846);
xor U4023 (N_4023,N_3817,N_3861);
nand U4024 (N_4024,N_3988,N_3825);
and U4025 (N_4025,N_3982,N_3913);
xor U4026 (N_4026,N_3929,N_3966);
and U4027 (N_4027,N_3935,N_3800);
nand U4028 (N_4028,N_3828,N_3879);
nand U4029 (N_4029,N_3830,N_3974);
xnor U4030 (N_4030,N_3852,N_3933);
xnor U4031 (N_4031,N_3853,N_3821);
and U4032 (N_4032,N_3880,N_3808);
and U4033 (N_4033,N_3922,N_3802);
xnor U4034 (N_4034,N_3967,N_3897);
xnor U4035 (N_4035,N_3857,N_3985);
xor U4036 (N_4036,N_3927,N_3810);
nand U4037 (N_4037,N_3934,N_3931);
or U4038 (N_4038,N_3873,N_3854);
xor U4039 (N_4039,N_3983,N_3812);
xor U4040 (N_4040,N_3827,N_3993);
nand U4041 (N_4041,N_3870,N_3831);
nand U4042 (N_4042,N_3882,N_3940);
and U4043 (N_4043,N_3904,N_3847);
nand U4044 (N_4044,N_3842,N_3875);
and U4045 (N_4045,N_3968,N_3903);
nor U4046 (N_4046,N_3884,N_3951);
and U4047 (N_4047,N_3829,N_3930);
and U4048 (N_4048,N_3889,N_3932);
nand U4049 (N_4049,N_3864,N_3965);
xor U4050 (N_4050,N_3900,N_3921);
nand U4051 (N_4051,N_3894,N_3942);
xnor U4052 (N_4052,N_3938,N_3912);
xor U4053 (N_4053,N_3937,N_3964);
or U4054 (N_4054,N_3855,N_3991);
nand U4055 (N_4055,N_3848,N_3868);
xnor U4056 (N_4056,N_3898,N_3863);
or U4057 (N_4057,N_3885,N_3896);
nand U4058 (N_4058,N_3833,N_3891);
xnor U4059 (N_4059,N_3923,N_3843);
xnor U4060 (N_4060,N_3867,N_3826);
or U4061 (N_4061,N_3824,N_3836);
nor U4062 (N_4062,N_3943,N_3818);
nand U4063 (N_4063,N_3876,N_3981);
xnor U4064 (N_4064,N_3845,N_3941);
or U4065 (N_4065,N_3963,N_3975);
or U4066 (N_4066,N_3984,N_3820);
and U4067 (N_4067,N_3856,N_3950);
and U4068 (N_4068,N_3869,N_3901);
nand U4069 (N_4069,N_3961,N_3916);
and U4070 (N_4070,N_3890,N_3992);
or U4071 (N_4071,N_3878,N_3924);
nor U4072 (N_4072,N_3809,N_3851);
or U4073 (N_4073,N_3956,N_3996);
or U4074 (N_4074,N_3860,N_3958);
and U4075 (N_4075,N_3841,N_3910);
or U4076 (N_4076,N_3998,N_3978);
and U4077 (N_4077,N_3834,N_3850);
xnor U4078 (N_4078,N_3871,N_3919);
or U4079 (N_4079,N_3881,N_3907);
or U4080 (N_4080,N_3905,N_3844);
nor U4081 (N_4081,N_3969,N_3893);
nor U4082 (N_4082,N_3972,N_3859);
and U4083 (N_4083,N_3977,N_3886);
xnor U4084 (N_4084,N_3955,N_3801);
xnor U4085 (N_4085,N_3866,N_3997);
nor U4086 (N_4086,N_3949,N_3816);
nor U4087 (N_4087,N_3946,N_3883);
xnor U4088 (N_4088,N_3939,N_3971);
nor U4089 (N_4089,N_3952,N_3813);
xor U4090 (N_4090,N_3920,N_3805);
and U4091 (N_4091,N_3959,N_3954);
nand U4092 (N_4092,N_3970,N_3872);
and U4093 (N_4093,N_3947,N_3899);
nand U4094 (N_4094,N_3914,N_3917);
nor U4095 (N_4095,N_3858,N_3838);
nand U4096 (N_4096,N_3915,N_3895);
nor U4097 (N_4097,N_3906,N_3980);
xor U4098 (N_4098,N_3887,N_3960);
nor U4099 (N_4099,N_3999,N_3925);
nor U4100 (N_4100,N_3892,N_3989);
nand U4101 (N_4101,N_3958,N_3905);
and U4102 (N_4102,N_3950,N_3833);
nand U4103 (N_4103,N_3909,N_3999);
and U4104 (N_4104,N_3894,N_3961);
nor U4105 (N_4105,N_3841,N_3960);
nand U4106 (N_4106,N_3926,N_3971);
nand U4107 (N_4107,N_3973,N_3934);
nor U4108 (N_4108,N_3813,N_3890);
or U4109 (N_4109,N_3930,N_3830);
and U4110 (N_4110,N_3919,N_3895);
and U4111 (N_4111,N_3830,N_3965);
nand U4112 (N_4112,N_3972,N_3883);
nand U4113 (N_4113,N_3842,N_3917);
and U4114 (N_4114,N_3956,N_3942);
nor U4115 (N_4115,N_3970,N_3888);
xnor U4116 (N_4116,N_3994,N_3969);
and U4117 (N_4117,N_3892,N_3973);
xnor U4118 (N_4118,N_3838,N_3807);
xnor U4119 (N_4119,N_3932,N_3881);
nand U4120 (N_4120,N_3918,N_3851);
nor U4121 (N_4121,N_3946,N_3931);
or U4122 (N_4122,N_3811,N_3969);
nor U4123 (N_4123,N_3969,N_3868);
nor U4124 (N_4124,N_3804,N_3986);
and U4125 (N_4125,N_3925,N_3851);
xnor U4126 (N_4126,N_3978,N_3964);
nor U4127 (N_4127,N_3802,N_3891);
and U4128 (N_4128,N_3889,N_3966);
or U4129 (N_4129,N_3838,N_3917);
nor U4130 (N_4130,N_3820,N_3946);
nand U4131 (N_4131,N_3930,N_3957);
or U4132 (N_4132,N_3936,N_3880);
nor U4133 (N_4133,N_3823,N_3832);
or U4134 (N_4134,N_3968,N_3916);
nand U4135 (N_4135,N_3805,N_3917);
xnor U4136 (N_4136,N_3858,N_3965);
nand U4137 (N_4137,N_3930,N_3865);
nor U4138 (N_4138,N_3809,N_3802);
or U4139 (N_4139,N_3848,N_3971);
nor U4140 (N_4140,N_3988,N_3942);
and U4141 (N_4141,N_3862,N_3897);
nand U4142 (N_4142,N_3911,N_3951);
xnor U4143 (N_4143,N_3920,N_3875);
or U4144 (N_4144,N_3822,N_3834);
and U4145 (N_4145,N_3935,N_3927);
and U4146 (N_4146,N_3926,N_3888);
and U4147 (N_4147,N_3895,N_3965);
xor U4148 (N_4148,N_3908,N_3983);
xnor U4149 (N_4149,N_3821,N_3921);
nor U4150 (N_4150,N_3835,N_3958);
nand U4151 (N_4151,N_3932,N_3946);
nand U4152 (N_4152,N_3904,N_3856);
nand U4153 (N_4153,N_3979,N_3938);
xor U4154 (N_4154,N_3867,N_3974);
and U4155 (N_4155,N_3906,N_3941);
or U4156 (N_4156,N_3977,N_3803);
nand U4157 (N_4157,N_3873,N_3875);
xor U4158 (N_4158,N_3977,N_3979);
nor U4159 (N_4159,N_3880,N_3959);
xnor U4160 (N_4160,N_3843,N_3950);
or U4161 (N_4161,N_3975,N_3944);
xor U4162 (N_4162,N_3903,N_3800);
nor U4163 (N_4163,N_3865,N_3972);
nor U4164 (N_4164,N_3902,N_3842);
nand U4165 (N_4165,N_3822,N_3894);
or U4166 (N_4166,N_3910,N_3823);
or U4167 (N_4167,N_3850,N_3863);
and U4168 (N_4168,N_3933,N_3958);
nor U4169 (N_4169,N_3992,N_3978);
and U4170 (N_4170,N_3836,N_3941);
nand U4171 (N_4171,N_3979,N_3906);
nand U4172 (N_4172,N_3858,N_3994);
nand U4173 (N_4173,N_3984,N_3813);
xnor U4174 (N_4174,N_3859,N_3998);
and U4175 (N_4175,N_3996,N_3923);
xnor U4176 (N_4176,N_3887,N_3864);
or U4177 (N_4177,N_3860,N_3912);
xor U4178 (N_4178,N_3803,N_3889);
and U4179 (N_4179,N_3821,N_3802);
xor U4180 (N_4180,N_3881,N_3924);
nor U4181 (N_4181,N_3888,N_3852);
nand U4182 (N_4182,N_3995,N_3983);
nor U4183 (N_4183,N_3877,N_3856);
nor U4184 (N_4184,N_3979,N_3856);
or U4185 (N_4185,N_3968,N_3890);
xor U4186 (N_4186,N_3801,N_3832);
nand U4187 (N_4187,N_3918,N_3822);
nor U4188 (N_4188,N_3942,N_3994);
nand U4189 (N_4189,N_3949,N_3829);
or U4190 (N_4190,N_3903,N_3943);
nor U4191 (N_4191,N_3881,N_3801);
nand U4192 (N_4192,N_3807,N_3909);
or U4193 (N_4193,N_3982,N_3958);
or U4194 (N_4194,N_3884,N_3978);
nor U4195 (N_4195,N_3844,N_3901);
or U4196 (N_4196,N_3989,N_3897);
or U4197 (N_4197,N_3908,N_3879);
nand U4198 (N_4198,N_3873,N_3850);
nor U4199 (N_4199,N_3811,N_3857);
nand U4200 (N_4200,N_4024,N_4021);
nand U4201 (N_4201,N_4088,N_4064);
xor U4202 (N_4202,N_4149,N_4072);
or U4203 (N_4203,N_4125,N_4087);
nand U4204 (N_4204,N_4100,N_4075);
nor U4205 (N_4205,N_4077,N_4198);
and U4206 (N_4206,N_4124,N_4120);
nor U4207 (N_4207,N_4096,N_4029);
or U4208 (N_4208,N_4161,N_4113);
nand U4209 (N_4209,N_4111,N_4193);
xnor U4210 (N_4210,N_4162,N_4171);
nor U4211 (N_4211,N_4074,N_4079);
or U4212 (N_4212,N_4164,N_4176);
xor U4213 (N_4213,N_4151,N_4082);
xnor U4214 (N_4214,N_4032,N_4117);
or U4215 (N_4215,N_4057,N_4078);
nand U4216 (N_4216,N_4156,N_4060);
and U4217 (N_4217,N_4005,N_4007);
xor U4218 (N_4218,N_4013,N_4009);
xor U4219 (N_4219,N_4015,N_4014);
xor U4220 (N_4220,N_4002,N_4101);
nor U4221 (N_4221,N_4065,N_4146);
xor U4222 (N_4222,N_4140,N_4155);
or U4223 (N_4223,N_4027,N_4073);
nor U4224 (N_4224,N_4090,N_4030);
nor U4225 (N_4225,N_4043,N_4139);
xnor U4226 (N_4226,N_4016,N_4138);
or U4227 (N_4227,N_4046,N_4040);
xor U4228 (N_4228,N_4180,N_4160);
nor U4229 (N_4229,N_4006,N_4108);
xor U4230 (N_4230,N_4058,N_4035);
or U4231 (N_4231,N_4091,N_4053);
nand U4232 (N_4232,N_4026,N_4086);
nor U4233 (N_4233,N_4179,N_4131);
and U4234 (N_4234,N_4150,N_4039);
nor U4235 (N_4235,N_4056,N_4187);
xnor U4236 (N_4236,N_4092,N_4037);
xnor U4237 (N_4237,N_4188,N_4051);
nand U4238 (N_4238,N_4052,N_4054);
nand U4239 (N_4239,N_4134,N_4083);
nand U4240 (N_4240,N_4059,N_4038);
nand U4241 (N_4241,N_4033,N_4145);
xnor U4242 (N_4242,N_4197,N_4095);
nand U4243 (N_4243,N_4011,N_4069);
and U4244 (N_4244,N_4103,N_4104);
or U4245 (N_4245,N_4050,N_4094);
or U4246 (N_4246,N_4122,N_4135);
and U4247 (N_4247,N_4019,N_4110);
nand U4248 (N_4248,N_4148,N_4047);
xnor U4249 (N_4249,N_4128,N_4178);
or U4250 (N_4250,N_4012,N_4070);
nor U4251 (N_4251,N_4097,N_4173);
or U4252 (N_4252,N_4084,N_4185);
and U4253 (N_4253,N_4194,N_4022);
xor U4254 (N_4254,N_4042,N_4099);
or U4255 (N_4255,N_4031,N_4063);
or U4256 (N_4256,N_4023,N_4004);
xnor U4257 (N_4257,N_4020,N_4199);
or U4258 (N_4258,N_4067,N_4196);
or U4259 (N_4259,N_4028,N_4141);
nor U4260 (N_4260,N_4000,N_4085);
nand U4261 (N_4261,N_4010,N_4169);
nand U4262 (N_4262,N_4017,N_4089);
and U4263 (N_4263,N_4163,N_4093);
nand U4264 (N_4264,N_4183,N_4003);
xnor U4265 (N_4265,N_4142,N_4102);
and U4266 (N_4266,N_4066,N_4172);
and U4267 (N_4267,N_4129,N_4154);
and U4268 (N_4268,N_4132,N_4076);
and U4269 (N_4269,N_4175,N_4192);
and U4270 (N_4270,N_4152,N_4123);
or U4271 (N_4271,N_4158,N_4190);
or U4272 (N_4272,N_4177,N_4044);
xnor U4273 (N_4273,N_4191,N_4045);
xor U4274 (N_4274,N_4130,N_4112);
xnor U4275 (N_4275,N_4080,N_4001);
and U4276 (N_4276,N_4144,N_4181);
and U4277 (N_4277,N_4127,N_4157);
or U4278 (N_4278,N_4186,N_4114);
nand U4279 (N_4279,N_4195,N_4167);
nand U4280 (N_4280,N_4126,N_4121);
and U4281 (N_4281,N_4133,N_4116);
and U4282 (N_4282,N_4143,N_4041);
xor U4283 (N_4283,N_4018,N_4159);
nand U4284 (N_4284,N_4107,N_4008);
nor U4285 (N_4285,N_4025,N_4061);
xnor U4286 (N_4286,N_4115,N_4118);
and U4287 (N_4287,N_4189,N_4106);
xnor U4288 (N_4288,N_4136,N_4048);
and U4289 (N_4289,N_4049,N_4109);
and U4290 (N_4290,N_4174,N_4147);
and U4291 (N_4291,N_4184,N_4105);
or U4292 (N_4292,N_4098,N_4170);
xor U4293 (N_4293,N_4068,N_4119);
xnor U4294 (N_4294,N_4034,N_4153);
or U4295 (N_4295,N_4165,N_4071);
xnor U4296 (N_4296,N_4081,N_4166);
xnor U4297 (N_4297,N_4137,N_4062);
xnor U4298 (N_4298,N_4168,N_4182);
and U4299 (N_4299,N_4055,N_4036);
xnor U4300 (N_4300,N_4034,N_4022);
xor U4301 (N_4301,N_4020,N_4182);
xor U4302 (N_4302,N_4163,N_4197);
nor U4303 (N_4303,N_4019,N_4035);
or U4304 (N_4304,N_4120,N_4138);
or U4305 (N_4305,N_4018,N_4130);
xnor U4306 (N_4306,N_4153,N_4161);
nand U4307 (N_4307,N_4096,N_4032);
nand U4308 (N_4308,N_4023,N_4088);
xor U4309 (N_4309,N_4033,N_4158);
nand U4310 (N_4310,N_4193,N_4014);
nand U4311 (N_4311,N_4180,N_4052);
xnor U4312 (N_4312,N_4000,N_4055);
and U4313 (N_4313,N_4149,N_4120);
nand U4314 (N_4314,N_4194,N_4186);
xor U4315 (N_4315,N_4147,N_4107);
nor U4316 (N_4316,N_4069,N_4159);
or U4317 (N_4317,N_4088,N_4053);
nand U4318 (N_4318,N_4188,N_4190);
xnor U4319 (N_4319,N_4163,N_4047);
or U4320 (N_4320,N_4152,N_4064);
or U4321 (N_4321,N_4190,N_4168);
nor U4322 (N_4322,N_4047,N_4195);
nand U4323 (N_4323,N_4085,N_4178);
xnor U4324 (N_4324,N_4050,N_4000);
or U4325 (N_4325,N_4087,N_4080);
xor U4326 (N_4326,N_4104,N_4186);
nand U4327 (N_4327,N_4088,N_4193);
xnor U4328 (N_4328,N_4145,N_4103);
and U4329 (N_4329,N_4095,N_4161);
and U4330 (N_4330,N_4167,N_4033);
nand U4331 (N_4331,N_4147,N_4025);
xnor U4332 (N_4332,N_4026,N_4142);
and U4333 (N_4333,N_4181,N_4015);
or U4334 (N_4334,N_4076,N_4094);
and U4335 (N_4335,N_4028,N_4132);
nand U4336 (N_4336,N_4009,N_4052);
nor U4337 (N_4337,N_4181,N_4076);
nor U4338 (N_4338,N_4010,N_4060);
nand U4339 (N_4339,N_4194,N_4145);
xnor U4340 (N_4340,N_4047,N_4056);
nand U4341 (N_4341,N_4076,N_4153);
or U4342 (N_4342,N_4103,N_4023);
nand U4343 (N_4343,N_4097,N_4036);
nor U4344 (N_4344,N_4036,N_4019);
or U4345 (N_4345,N_4026,N_4113);
xnor U4346 (N_4346,N_4044,N_4156);
nand U4347 (N_4347,N_4197,N_4086);
or U4348 (N_4348,N_4078,N_4018);
nor U4349 (N_4349,N_4062,N_4078);
or U4350 (N_4350,N_4139,N_4108);
or U4351 (N_4351,N_4071,N_4126);
nand U4352 (N_4352,N_4186,N_4190);
and U4353 (N_4353,N_4057,N_4016);
nor U4354 (N_4354,N_4038,N_4131);
xnor U4355 (N_4355,N_4041,N_4070);
or U4356 (N_4356,N_4136,N_4122);
and U4357 (N_4357,N_4068,N_4048);
nand U4358 (N_4358,N_4150,N_4165);
nor U4359 (N_4359,N_4030,N_4023);
nor U4360 (N_4360,N_4193,N_4013);
nand U4361 (N_4361,N_4087,N_4166);
nor U4362 (N_4362,N_4167,N_4134);
nor U4363 (N_4363,N_4006,N_4101);
nand U4364 (N_4364,N_4027,N_4041);
nand U4365 (N_4365,N_4059,N_4091);
xnor U4366 (N_4366,N_4075,N_4024);
xor U4367 (N_4367,N_4091,N_4153);
or U4368 (N_4368,N_4054,N_4117);
nand U4369 (N_4369,N_4161,N_4192);
or U4370 (N_4370,N_4092,N_4129);
xnor U4371 (N_4371,N_4177,N_4099);
or U4372 (N_4372,N_4028,N_4183);
or U4373 (N_4373,N_4078,N_4003);
nand U4374 (N_4374,N_4050,N_4154);
or U4375 (N_4375,N_4168,N_4069);
nand U4376 (N_4376,N_4140,N_4161);
or U4377 (N_4377,N_4190,N_4159);
or U4378 (N_4378,N_4157,N_4105);
and U4379 (N_4379,N_4147,N_4151);
or U4380 (N_4380,N_4125,N_4107);
nor U4381 (N_4381,N_4147,N_4087);
nor U4382 (N_4382,N_4031,N_4185);
and U4383 (N_4383,N_4105,N_4177);
nand U4384 (N_4384,N_4095,N_4117);
and U4385 (N_4385,N_4171,N_4060);
xnor U4386 (N_4386,N_4102,N_4127);
xnor U4387 (N_4387,N_4088,N_4087);
and U4388 (N_4388,N_4010,N_4189);
xnor U4389 (N_4389,N_4163,N_4154);
and U4390 (N_4390,N_4161,N_4150);
and U4391 (N_4391,N_4025,N_4053);
and U4392 (N_4392,N_4028,N_4083);
nor U4393 (N_4393,N_4051,N_4138);
and U4394 (N_4394,N_4128,N_4147);
nor U4395 (N_4395,N_4036,N_4007);
nor U4396 (N_4396,N_4117,N_4128);
nand U4397 (N_4397,N_4183,N_4113);
xor U4398 (N_4398,N_4192,N_4120);
nand U4399 (N_4399,N_4002,N_4181);
and U4400 (N_4400,N_4288,N_4251);
and U4401 (N_4401,N_4321,N_4216);
nor U4402 (N_4402,N_4232,N_4294);
nor U4403 (N_4403,N_4206,N_4241);
xor U4404 (N_4404,N_4276,N_4371);
nor U4405 (N_4405,N_4240,N_4345);
nor U4406 (N_4406,N_4282,N_4360);
or U4407 (N_4407,N_4292,N_4304);
or U4408 (N_4408,N_4222,N_4226);
or U4409 (N_4409,N_4225,N_4395);
nand U4410 (N_4410,N_4265,N_4387);
nor U4411 (N_4411,N_4388,N_4355);
nand U4412 (N_4412,N_4249,N_4394);
or U4413 (N_4413,N_4390,N_4363);
or U4414 (N_4414,N_4343,N_4309);
or U4415 (N_4415,N_4380,N_4237);
xnor U4416 (N_4416,N_4376,N_4213);
nand U4417 (N_4417,N_4257,N_4381);
or U4418 (N_4418,N_4305,N_4219);
nor U4419 (N_4419,N_4353,N_4378);
or U4420 (N_4420,N_4379,N_4324);
nand U4421 (N_4421,N_4272,N_4382);
xor U4422 (N_4422,N_4215,N_4341);
nor U4423 (N_4423,N_4260,N_4220);
and U4424 (N_4424,N_4366,N_4290);
nand U4425 (N_4425,N_4253,N_4359);
xnor U4426 (N_4426,N_4296,N_4263);
or U4427 (N_4427,N_4383,N_4227);
or U4428 (N_4428,N_4342,N_4233);
xor U4429 (N_4429,N_4391,N_4370);
or U4430 (N_4430,N_4362,N_4392);
and U4431 (N_4431,N_4397,N_4223);
nor U4432 (N_4432,N_4331,N_4314);
or U4433 (N_4433,N_4350,N_4361);
and U4434 (N_4434,N_4268,N_4386);
xnor U4435 (N_4435,N_4235,N_4357);
nor U4436 (N_4436,N_4340,N_4334);
nand U4437 (N_4437,N_4330,N_4356);
nor U4438 (N_4438,N_4275,N_4325);
nand U4439 (N_4439,N_4308,N_4218);
or U4440 (N_4440,N_4283,N_4238);
or U4441 (N_4441,N_4393,N_4254);
xor U4442 (N_4442,N_4295,N_4312);
or U4443 (N_4443,N_4313,N_4320);
or U4444 (N_4444,N_4259,N_4236);
and U4445 (N_4445,N_4375,N_4245);
xnor U4446 (N_4446,N_4248,N_4372);
and U4447 (N_4447,N_4205,N_4246);
nor U4448 (N_4448,N_4270,N_4298);
xor U4449 (N_4449,N_4211,N_4317);
nor U4450 (N_4450,N_4396,N_4347);
nor U4451 (N_4451,N_4207,N_4374);
xor U4452 (N_4452,N_4252,N_4250);
or U4453 (N_4453,N_4293,N_4287);
or U4454 (N_4454,N_4255,N_4316);
or U4455 (N_4455,N_4285,N_4289);
xor U4456 (N_4456,N_4299,N_4351);
and U4457 (N_4457,N_4369,N_4318);
nand U4458 (N_4458,N_4297,N_4367);
nand U4459 (N_4459,N_4291,N_4322);
nand U4460 (N_4460,N_4337,N_4203);
nor U4461 (N_4461,N_4224,N_4242);
and U4462 (N_4462,N_4271,N_4286);
or U4463 (N_4463,N_4239,N_4373);
nor U4464 (N_4464,N_4258,N_4365);
or U4465 (N_4465,N_4349,N_4210);
and U4466 (N_4466,N_4384,N_4319);
and U4467 (N_4467,N_4266,N_4310);
nor U4468 (N_4468,N_4354,N_4221);
nand U4469 (N_4469,N_4230,N_4280);
and U4470 (N_4470,N_4368,N_4329);
nor U4471 (N_4471,N_4311,N_4267);
xor U4472 (N_4472,N_4214,N_4323);
or U4473 (N_4473,N_4303,N_4256);
xnor U4474 (N_4474,N_4389,N_4302);
or U4475 (N_4475,N_4228,N_4358);
and U4476 (N_4476,N_4243,N_4307);
nor U4477 (N_4477,N_4247,N_4281);
and U4478 (N_4478,N_4332,N_4244);
or U4479 (N_4479,N_4277,N_4273);
or U4480 (N_4480,N_4279,N_4333);
and U4481 (N_4481,N_4399,N_4264);
nor U4482 (N_4482,N_4202,N_4326);
xnor U4483 (N_4483,N_4339,N_4377);
or U4484 (N_4484,N_4278,N_4327);
nand U4485 (N_4485,N_4364,N_4209);
xnor U4486 (N_4486,N_4346,N_4398);
nand U4487 (N_4487,N_4208,N_4229);
or U4488 (N_4488,N_4200,N_4212);
nor U4489 (N_4489,N_4385,N_4262);
nor U4490 (N_4490,N_4217,N_4335);
and U4491 (N_4491,N_4201,N_4301);
xnor U4492 (N_4492,N_4234,N_4348);
or U4493 (N_4493,N_4352,N_4336);
nor U4494 (N_4494,N_4261,N_4269);
and U4495 (N_4495,N_4306,N_4344);
nand U4496 (N_4496,N_4328,N_4300);
or U4497 (N_4497,N_4338,N_4284);
xnor U4498 (N_4498,N_4204,N_4274);
nor U4499 (N_4499,N_4315,N_4231);
xor U4500 (N_4500,N_4278,N_4213);
or U4501 (N_4501,N_4293,N_4244);
or U4502 (N_4502,N_4328,N_4314);
nor U4503 (N_4503,N_4213,N_4335);
and U4504 (N_4504,N_4362,N_4354);
nor U4505 (N_4505,N_4391,N_4205);
or U4506 (N_4506,N_4213,N_4248);
nand U4507 (N_4507,N_4299,N_4358);
nor U4508 (N_4508,N_4336,N_4285);
xor U4509 (N_4509,N_4349,N_4268);
and U4510 (N_4510,N_4327,N_4261);
nor U4511 (N_4511,N_4246,N_4305);
and U4512 (N_4512,N_4340,N_4318);
nand U4513 (N_4513,N_4365,N_4215);
and U4514 (N_4514,N_4312,N_4398);
or U4515 (N_4515,N_4247,N_4344);
and U4516 (N_4516,N_4356,N_4288);
nand U4517 (N_4517,N_4373,N_4292);
nor U4518 (N_4518,N_4236,N_4230);
or U4519 (N_4519,N_4318,N_4259);
or U4520 (N_4520,N_4322,N_4247);
or U4521 (N_4521,N_4289,N_4346);
or U4522 (N_4522,N_4249,N_4350);
and U4523 (N_4523,N_4336,N_4387);
or U4524 (N_4524,N_4210,N_4235);
and U4525 (N_4525,N_4316,N_4281);
xnor U4526 (N_4526,N_4344,N_4239);
nand U4527 (N_4527,N_4262,N_4272);
xor U4528 (N_4528,N_4340,N_4337);
nor U4529 (N_4529,N_4382,N_4381);
nand U4530 (N_4530,N_4252,N_4348);
nand U4531 (N_4531,N_4289,N_4284);
xnor U4532 (N_4532,N_4396,N_4269);
nand U4533 (N_4533,N_4217,N_4249);
nand U4534 (N_4534,N_4260,N_4377);
and U4535 (N_4535,N_4274,N_4283);
and U4536 (N_4536,N_4291,N_4245);
and U4537 (N_4537,N_4395,N_4373);
nor U4538 (N_4538,N_4328,N_4288);
nor U4539 (N_4539,N_4300,N_4290);
and U4540 (N_4540,N_4275,N_4208);
and U4541 (N_4541,N_4256,N_4227);
nand U4542 (N_4542,N_4266,N_4384);
and U4543 (N_4543,N_4397,N_4336);
nand U4544 (N_4544,N_4212,N_4259);
nand U4545 (N_4545,N_4202,N_4337);
and U4546 (N_4546,N_4317,N_4364);
or U4547 (N_4547,N_4234,N_4379);
nand U4548 (N_4548,N_4297,N_4225);
xnor U4549 (N_4549,N_4275,N_4323);
nor U4550 (N_4550,N_4226,N_4372);
nor U4551 (N_4551,N_4309,N_4370);
nand U4552 (N_4552,N_4334,N_4324);
xnor U4553 (N_4553,N_4301,N_4300);
or U4554 (N_4554,N_4213,N_4221);
or U4555 (N_4555,N_4242,N_4291);
xnor U4556 (N_4556,N_4319,N_4242);
and U4557 (N_4557,N_4336,N_4343);
nor U4558 (N_4558,N_4231,N_4256);
xnor U4559 (N_4559,N_4266,N_4232);
or U4560 (N_4560,N_4228,N_4348);
or U4561 (N_4561,N_4321,N_4306);
xor U4562 (N_4562,N_4248,N_4204);
nand U4563 (N_4563,N_4378,N_4372);
nor U4564 (N_4564,N_4225,N_4348);
and U4565 (N_4565,N_4396,N_4338);
nor U4566 (N_4566,N_4335,N_4324);
nor U4567 (N_4567,N_4299,N_4319);
and U4568 (N_4568,N_4315,N_4266);
nor U4569 (N_4569,N_4259,N_4330);
and U4570 (N_4570,N_4243,N_4246);
xnor U4571 (N_4571,N_4359,N_4277);
nor U4572 (N_4572,N_4231,N_4335);
or U4573 (N_4573,N_4226,N_4286);
nand U4574 (N_4574,N_4319,N_4392);
xor U4575 (N_4575,N_4351,N_4257);
and U4576 (N_4576,N_4338,N_4272);
xor U4577 (N_4577,N_4222,N_4333);
and U4578 (N_4578,N_4347,N_4226);
and U4579 (N_4579,N_4307,N_4372);
and U4580 (N_4580,N_4240,N_4286);
and U4581 (N_4581,N_4324,N_4261);
nand U4582 (N_4582,N_4334,N_4365);
or U4583 (N_4583,N_4273,N_4365);
xor U4584 (N_4584,N_4367,N_4379);
and U4585 (N_4585,N_4376,N_4237);
xor U4586 (N_4586,N_4374,N_4200);
xor U4587 (N_4587,N_4310,N_4343);
or U4588 (N_4588,N_4335,N_4379);
or U4589 (N_4589,N_4243,N_4233);
nand U4590 (N_4590,N_4224,N_4280);
or U4591 (N_4591,N_4278,N_4269);
nand U4592 (N_4592,N_4329,N_4208);
nor U4593 (N_4593,N_4330,N_4241);
xor U4594 (N_4594,N_4311,N_4269);
nor U4595 (N_4595,N_4317,N_4206);
and U4596 (N_4596,N_4396,N_4316);
and U4597 (N_4597,N_4262,N_4319);
xor U4598 (N_4598,N_4358,N_4322);
or U4599 (N_4599,N_4212,N_4252);
xor U4600 (N_4600,N_4580,N_4578);
nor U4601 (N_4601,N_4450,N_4498);
or U4602 (N_4602,N_4454,N_4595);
or U4603 (N_4603,N_4509,N_4572);
or U4604 (N_4604,N_4539,N_4582);
nor U4605 (N_4605,N_4500,N_4585);
xnor U4606 (N_4606,N_4508,N_4577);
nand U4607 (N_4607,N_4431,N_4594);
nor U4608 (N_4608,N_4523,N_4567);
nand U4609 (N_4609,N_4401,N_4404);
xnor U4610 (N_4610,N_4546,N_4552);
and U4611 (N_4611,N_4569,N_4525);
nor U4612 (N_4612,N_4441,N_4427);
nand U4613 (N_4613,N_4415,N_4571);
and U4614 (N_4614,N_4583,N_4501);
or U4615 (N_4615,N_4403,N_4471);
nor U4616 (N_4616,N_4599,N_4545);
xor U4617 (N_4617,N_4570,N_4531);
and U4618 (N_4618,N_4555,N_4432);
and U4619 (N_4619,N_4414,N_4452);
and U4620 (N_4620,N_4557,N_4460);
xnor U4621 (N_4621,N_4444,N_4536);
or U4622 (N_4622,N_4544,N_4458);
nor U4623 (N_4623,N_4436,N_4459);
or U4624 (N_4624,N_4475,N_4521);
nor U4625 (N_4625,N_4519,N_4413);
and U4626 (N_4626,N_4439,N_4514);
nor U4627 (N_4627,N_4551,N_4487);
nor U4628 (N_4628,N_4425,N_4474);
nor U4629 (N_4629,N_4596,N_4517);
nand U4630 (N_4630,N_4532,N_4593);
or U4631 (N_4631,N_4479,N_4575);
nor U4632 (N_4632,N_4476,N_4558);
or U4633 (N_4633,N_4402,N_4467);
or U4634 (N_4634,N_4563,N_4576);
nor U4635 (N_4635,N_4535,N_4507);
nor U4636 (N_4636,N_4482,N_4559);
or U4637 (N_4637,N_4588,N_4520);
or U4638 (N_4638,N_4416,N_4579);
and U4639 (N_4639,N_4455,N_4481);
and U4640 (N_4640,N_4472,N_4564);
nor U4641 (N_4641,N_4527,N_4574);
xor U4642 (N_4642,N_4448,N_4524);
xor U4643 (N_4643,N_4549,N_4589);
nand U4644 (N_4644,N_4473,N_4463);
nor U4645 (N_4645,N_4518,N_4566);
nand U4646 (N_4646,N_4543,N_4541);
nor U4647 (N_4647,N_4438,N_4503);
xnor U4648 (N_4648,N_4483,N_4417);
nand U4649 (N_4649,N_4429,N_4548);
and U4650 (N_4650,N_4553,N_4499);
nand U4651 (N_4651,N_4485,N_4464);
nand U4652 (N_4652,N_4528,N_4491);
nor U4653 (N_4653,N_4550,N_4470);
xnor U4654 (N_4654,N_4408,N_4540);
nor U4655 (N_4655,N_4469,N_4405);
nand U4656 (N_4656,N_4443,N_4573);
and U4657 (N_4657,N_4530,N_4445);
and U4658 (N_4658,N_4592,N_4440);
nor U4659 (N_4659,N_4480,N_4490);
nor U4660 (N_4660,N_4465,N_4492);
or U4661 (N_4661,N_4495,N_4468);
or U4662 (N_4662,N_4554,N_4505);
or U4663 (N_4663,N_4598,N_4462);
nor U4664 (N_4664,N_4494,N_4420);
nand U4665 (N_4665,N_4510,N_4533);
or U4666 (N_4666,N_4424,N_4561);
nor U4667 (N_4667,N_4502,N_4496);
or U4668 (N_4668,N_4457,N_4449);
and U4669 (N_4669,N_4437,N_4506);
nor U4670 (N_4670,N_4581,N_4542);
and U4671 (N_4671,N_4400,N_4522);
and U4672 (N_4672,N_4422,N_4421);
nor U4673 (N_4673,N_4537,N_4466);
xor U4674 (N_4674,N_4419,N_4504);
or U4675 (N_4675,N_4586,N_4411);
xor U4676 (N_4676,N_4410,N_4512);
nand U4677 (N_4677,N_4513,N_4516);
nor U4678 (N_4678,N_4461,N_4515);
or U4679 (N_4679,N_4456,N_4547);
xnor U4680 (N_4680,N_4562,N_4434);
nand U4681 (N_4681,N_4591,N_4560);
and U4682 (N_4682,N_4584,N_4477);
and U4683 (N_4683,N_4478,N_4407);
or U4684 (N_4684,N_4428,N_4409);
nand U4685 (N_4685,N_4426,N_4534);
nand U4686 (N_4686,N_4430,N_4511);
and U4687 (N_4687,N_4568,N_4423);
xor U4688 (N_4688,N_4442,N_4526);
nor U4689 (N_4689,N_4486,N_4451);
nand U4690 (N_4690,N_4488,N_4587);
nor U4691 (N_4691,N_4433,N_4412);
xnor U4692 (N_4692,N_4446,N_4418);
xnor U4693 (N_4693,N_4435,N_4453);
nand U4694 (N_4694,N_4538,N_4565);
or U4695 (N_4695,N_4556,N_4493);
xnor U4696 (N_4696,N_4484,N_4447);
nor U4697 (N_4697,N_4406,N_4590);
and U4698 (N_4698,N_4497,N_4529);
nand U4699 (N_4699,N_4489,N_4597);
xor U4700 (N_4700,N_4549,N_4507);
nor U4701 (N_4701,N_4431,N_4574);
and U4702 (N_4702,N_4468,N_4580);
nor U4703 (N_4703,N_4437,N_4556);
nor U4704 (N_4704,N_4452,N_4537);
and U4705 (N_4705,N_4454,N_4446);
xnor U4706 (N_4706,N_4404,N_4580);
and U4707 (N_4707,N_4522,N_4555);
or U4708 (N_4708,N_4424,N_4497);
nor U4709 (N_4709,N_4448,N_4523);
nand U4710 (N_4710,N_4413,N_4406);
or U4711 (N_4711,N_4537,N_4494);
xor U4712 (N_4712,N_4411,N_4590);
nand U4713 (N_4713,N_4504,N_4421);
nand U4714 (N_4714,N_4537,N_4423);
nor U4715 (N_4715,N_4484,N_4511);
xor U4716 (N_4716,N_4554,N_4424);
and U4717 (N_4717,N_4439,N_4447);
and U4718 (N_4718,N_4560,N_4476);
xnor U4719 (N_4719,N_4524,N_4590);
nand U4720 (N_4720,N_4554,N_4460);
and U4721 (N_4721,N_4426,N_4561);
or U4722 (N_4722,N_4402,N_4407);
and U4723 (N_4723,N_4555,N_4419);
and U4724 (N_4724,N_4512,N_4543);
nor U4725 (N_4725,N_4592,N_4547);
nand U4726 (N_4726,N_4547,N_4420);
nor U4727 (N_4727,N_4483,N_4555);
and U4728 (N_4728,N_4517,N_4541);
xor U4729 (N_4729,N_4563,N_4402);
or U4730 (N_4730,N_4591,N_4461);
or U4731 (N_4731,N_4456,N_4421);
and U4732 (N_4732,N_4574,N_4487);
or U4733 (N_4733,N_4511,N_4464);
xor U4734 (N_4734,N_4487,N_4521);
or U4735 (N_4735,N_4543,N_4425);
or U4736 (N_4736,N_4537,N_4536);
xnor U4737 (N_4737,N_4553,N_4470);
xor U4738 (N_4738,N_4452,N_4518);
and U4739 (N_4739,N_4588,N_4504);
nor U4740 (N_4740,N_4406,N_4581);
or U4741 (N_4741,N_4426,N_4493);
xor U4742 (N_4742,N_4539,N_4467);
and U4743 (N_4743,N_4495,N_4426);
and U4744 (N_4744,N_4449,N_4414);
or U4745 (N_4745,N_4560,N_4571);
and U4746 (N_4746,N_4514,N_4461);
nor U4747 (N_4747,N_4416,N_4489);
nor U4748 (N_4748,N_4585,N_4484);
and U4749 (N_4749,N_4584,N_4543);
xor U4750 (N_4750,N_4478,N_4529);
and U4751 (N_4751,N_4471,N_4470);
nor U4752 (N_4752,N_4595,N_4459);
and U4753 (N_4753,N_4482,N_4551);
nor U4754 (N_4754,N_4501,N_4450);
and U4755 (N_4755,N_4400,N_4596);
and U4756 (N_4756,N_4437,N_4401);
nand U4757 (N_4757,N_4488,N_4440);
and U4758 (N_4758,N_4471,N_4410);
xnor U4759 (N_4759,N_4500,N_4535);
nand U4760 (N_4760,N_4497,N_4554);
or U4761 (N_4761,N_4466,N_4458);
nor U4762 (N_4762,N_4509,N_4521);
nor U4763 (N_4763,N_4508,N_4488);
nor U4764 (N_4764,N_4416,N_4566);
nand U4765 (N_4765,N_4549,N_4560);
xnor U4766 (N_4766,N_4554,N_4431);
xor U4767 (N_4767,N_4455,N_4464);
and U4768 (N_4768,N_4580,N_4467);
nand U4769 (N_4769,N_4435,N_4417);
and U4770 (N_4770,N_4583,N_4409);
nand U4771 (N_4771,N_4461,N_4403);
nand U4772 (N_4772,N_4495,N_4404);
and U4773 (N_4773,N_4509,N_4567);
nor U4774 (N_4774,N_4417,N_4541);
or U4775 (N_4775,N_4441,N_4417);
nand U4776 (N_4776,N_4556,N_4463);
xor U4777 (N_4777,N_4554,N_4514);
and U4778 (N_4778,N_4530,N_4430);
or U4779 (N_4779,N_4560,N_4410);
nor U4780 (N_4780,N_4448,N_4541);
nor U4781 (N_4781,N_4461,N_4586);
nand U4782 (N_4782,N_4444,N_4510);
or U4783 (N_4783,N_4495,N_4503);
nand U4784 (N_4784,N_4510,N_4528);
or U4785 (N_4785,N_4472,N_4420);
nor U4786 (N_4786,N_4554,N_4563);
nand U4787 (N_4787,N_4519,N_4515);
xnor U4788 (N_4788,N_4483,N_4442);
xor U4789 (N_4789,N_4503,N_4436);
and U4790 (N_4790,N_4481,N_4509);
xnor U4791 (N_4791,N_4577,N_4471);
or U4792 (N_4792,N_4490,N_4477);
and U4793 (N_4793,N_4415,N_4577);
xnor U4794 (N_4794,N_4537,N_4442);
and U4795 (N_4795,N_4598,N_4529);
nor U4796 (N_4796,N_4524,N_4556);
xnor U4797 (N_4797,N_4450,N_4594);
xor U4798 (N_4798,N_4413,N_4581);
or U4799 (N_4799,N_4473,N_4436);
xor U4800 (N_4800,N_4734,N_4687);
nand U4801 (N_4801,N_4602,N_4711);
and U4802 (N_4802,N_4788,N_4759);
and U4803 (N_4803,N_4621,N_4681);
and U4804 (N_4804,N_4715,N_4749);
and U4805 (N_4805,N_4771,N_4737);
xor U4806 (N_4806,N_4779,N_4689);
nand U4807 (N_4807,N_4696,N_4694);
nor U4808 (N_4808,N_4667,N_4656);
or U4809 (N_4809,N_4795,N_4730);
nand U4810 (N_4810,N_4692,N_4635);
nor U4811 (N_4811,N_4792,N_4761);
xnor U4812 (N_4812,N_4740,N_4723);
nand U4813 (N_4813,N_4733,N_4695);
or U4814 (N_4814,N_4618,N_4698);
nor U4815 (N_4815,N_4744,N_4796);
or U4816 (N_4816,N_4630,N_4799);
nor U4817 (N_4817,N_4606,N_4641);
nor U4818 (N_4818,N_4646,N_4678);
and U4819 (N_4819,N_4751,N_4676);
nand U4820 (N_4820,N_4775,N_4750);
and U4821 (N_4821,N_4739,N_4600);
nor U4822 (N_4822,N_4701,N_4728);
nand U4823 (N_4823,N_4679,N_4675);
or U4824 (N_4824,N_4755,N_4607);
or U4825 (N_4825,N_4706,N_4768);
nand U4826 (N_4826,N_4625,N_4639);
or U4827 (N_4827,N_4713,N_4791);
xnor U4828 (N_4828,N_4662,N_4651);
or U4829 (N_4829,N_4727,N_4649);
xnor U4830 (N_4830,N_4721,N_4684);
nor U4831 (N_4831,N_4783,N_4738);
xor U4832 (N_4832,N_4622,N_4620);
nor U4833 (N_4833,N_4798,N_4729);
and U4834 (N_4834,N_4619,N_4776);
or U4835 (N_4835,N_4781,N_4793);
and U4836 (N_4836,N_4627,N_4677);
xnor U4837 (N_4837,N_4797,N_4787);
nor U4838 (N_4838,N_4611,N_4688);
xor U4839 (N_4839,N_4774,N_4609);
and U4840 (N_4840,N_4770,N_4608);
and U4841 (N_4841,N_4741,N_4682);
and U4842 (N_4842,N_4605,N_4708);
or U4843 (N_4843,N_4742,N_4754);
and U4844 (N_4844,N_4665,N_4642);
xor U4845 (N_4845,N_4648,N_4702);
nand U4846 (N_4846,N_4636,N_4716);
or U4847 (N_4847,N_4780,N_4757);
or U4848 (N_4848,N_4637,N_4617);
nor U4849 (N_4849,N_4722,N_4731);
or U4850 (N_4850,N_4735,N_4743);
and U4851 (N_4851,N_4640,N_4720);
xor U4852 (N_4852,N_4707,N_4683);
xnor U4853 (N_4853,N_4659,N_4736);
or U4854 (N_4854,N_4756,N_4714);
xnor U4855 (N_4855,N_4745,N_4645);
or U4856 (N_4856,N_4763,N_4658);
or U4857 (N_4857,N_4686,N_4638);
or U4858 (N_4858,N_4670,N_4657);
xor U4859 (N_4859,N_4712,N_4612);
nand U4860 (N_4860,N_4685,N_4760);
or U4861 (N_4861,N_4786,N_4710);
and U4862 (N_4862,N_4614,N_4747);
or U4863 (N_4863,N_4664,N_4601);
and U4864 (N_4864,N_4691,N_4703);
and U4865 (N_4865,N_4752,N_4690);
nand U4866 (N_4866,N_4704,N_4773);
or U4867 (N_4867,N_4753,N_4652);
xnor U4868 (N_4868,N_4661,N_4623);
nand U4869 (N_4869,N_4697,N_4766);
nand U4870 (N_4870,N_4785,N_4671);
nor U4871 (N_4871,N_4790,N_4650);
xnor U4872 (N_4872,N_4655,N_4724);
and U4873 (N_4873,N_4604,N_4789);
nor U4874 (N_4874,N_4719,N_4748);
and U4875 (N_4875,N_4772,N_4647);
nor U4876 (N_4876,N_4634,N_4767);
or U4877 (N_4877,N_4699,N_4643);
and U4878 (N_4878,N_4633,N_4709);
or U4879 (N_4879,N_4764,N_4717);
xnor U4880 (N_4880,N_4732,N_4718);
or U4881 (N_4881,N_4680,N_4654);
nand U4882 (N_4882,N_4610,N_4624);
nand U4883 (N_4883,N_4626,N_4725);
or U4884 (N_4884,N_4663,N_4631);
xor U4885 (N_4885,N_4758,N_4616);
nand U4886 (N_4886,N_4660,N_4784);
and U4887 (N_4887,N_4782,N_4632);
nand U4888 (N_4888,N_4726,N_4700);
nand U4889 (N_4889,N_4705,N_4673);
xnor U4890 (N_4890,N_4628,N_4746);
or U4891 (N_4891,N_4672,N_4668);
or U4892 (N_4892,N_4778,N_4666);
or U4893 (N_4893,N_4613,N_4769);
nor U4894 (N_4894,N_4629,N_4674);
and U4895 (N_4895,N_4765,N_4693);
nand U4896 (N_4896,N_4653,N_4615);
or U4897 (N_4897,N_4644,N_4669);
nand U4898 (N_4898,N_4762,N_4777);
nand U4899 (N_4899,N_4603,N_4794);
and U4900 (N_4900,N_4641,N_4692);
xor U4901 (N_4901,N_4621,N_4760);
xnor U4902 (N_4902,N_4735,N_4699);
or U4903 (N_4903,N_4775,N_4675);
or U4904 (N_4904,N_4642,N_4779);
xnor U4905 (N_4905,N_4652,N_4682);
and U4906 (N_4906,N_4758,N_4700);
or U4907 (N_4907,N_4782,N_4684);
nand U4908 (N_4908,N_4636,N_4619);
or U4909 (N_4909,N_4728,N_4730);
nor U4910 (N_4910,N_4663,N_4655);
nand U4911 (N_4911,N_4604,N_4761);
or U4912 (N_4912,N_4713,N_4673);
xor U4913 (N_4913,N_4642,N_4620);
or U4914 (N_4914,N_4723,N_4636);
nand U4915 (N_4915,N_4785,N_4747);
nand U4916 (N_4916,N_4680,N_4646);
or U4917 (N_4917,N_4680,N_4709);
nand U4918 (N_4918,N_4787,N_4657);
or U4919 (N_4919,N_4789,N_4603);
and U4920 (N_4920,N_4798,N_4649);
nand U4921 (N_4921,N_4605,N_4734);
xnor U4922 (N_4922,N_4739,N_4636);
or U4923 (N_4923,N_4608,N_4702);
and U4924 (N_4924,N_4627,N_4766);
or U4925 (N_4925,N_4625,N_4768);
nor U4926 (N_4926,N_4659,N_4667);
xor U4927 (N_4927,N_4799,N_4680);
nor U4928 (N_4928,N_4678,N_4773);
or U4929 (N_4929,N_4616,N_4608);
and U4930 (N_4930,N_4791,N_4620);
or U4931 (N_4931,N_4603,N_4671);
xor U4932 (N_4932,N_4687,N_4793);
nor U4933 (N_4933,N_4796,N_4733);
nand U4934 (N_4934,N_4692,N_4688);
nor U4935 (N_4935,N_4788,N_4776);
nand U4936 (N_4936,N_4680,N_4762);
or U4937 (N_4937,N_4789,N_4658);
nor U4938 (N_4938,N_4756,N_4668);
or U4939 (N_4939,N_4619,N_4631);
nand U4940 (N_4940,N_4653,N_4728);
nand U4941 (N_4941,N_4724,N_4658);
nand U4942 (N_4942,N_4711,N_4665);
and U4943 (N_4943,N_4673,N_4610);
xnor U4944 (N_4944,N_4702,N_4635);
or U4945 (N_4945,N_4789,N_4715);
or U4946 (N_4946,N_4612,N_4605);
and U4947 (N_4947,N_4681,N_4781);
and U4948 (N_4948,N_4745,N_4779);
and U4949 (N_4949,N_4672,N_4690);
nor U4950 (N_4950,N_4769,N_4788);
and U4951 (N_4951,N_4692,N_4639);
or U4952 (N_4952,N_4694,N_4732);
nand U4953 (N_4953,N_4775,N_4680);
or U4954 (N_4954,N_4608,N_4710);
and U4955 (N_4955,N_4610,N_4725);
or U4956 (N_4956,N_4676,N_4669);
xnor U4957 (N_4957,N_4714,N_4663);
xor U4958 (N_4958,N_4678,N_4709);
and U4959 (N_4959,N_4600,N_4724);
nor U4960 (N_4960,N_4694,N_4741);
nand U4961 (N_4961,N_4612,N_4692);
nand U4962 (N_4962,N_4635,N_4753);
nand U4963 (N_4963,N_4720,N_4648);
nor U4964 (N_4964,N_4728,N_4702);
or U4965 (N_4965,N_4749,N_4614);
xnor U4966 (N_4966,N_4680,N_4759);
and U4967 (N_4967,N_4706,N_4730);
nor U4968 (N_4968,N_4625,N_4700);
xnor U4969 (N_4969,N_4782,N_4761);
nand U4970 (N_4970,N_4706,N_4753);
nor U4971 (N_4971,N_4635,N_4639);
xor U4972 (N_4972,N_4767,N_4768);
nor U4973 (N_4973,N_4705,N_4631);
nand U4974 (N_4974,N_4793,N_4795);
or U4975 (N_4975,N_4737,N_4664);
nor U4976 (N_4976,N_4601,N_4630);
nor U4977 (N_4977,N_4608,N_4651);
xnor U4978 (N_4978,N_4748,N_4662);
and U4979 (N_4979,N_4736,N_4676);
xnor U4980 (N_4980,N_4685,N_4730);
or U4981 (N_4981,N_4716,N_4760);
and U4982 (N_4982,N_4714,N_4655);
and U4983 (N_4983,N_4718,N_4723);
nor U4984 (N_4984,N_4700,N_4799);
nand U4985 (N_4985,N_4712,N_4791);
xnor U4986 (N_4986,N_4626,N_4640);
or U4987 (N_4987,N_4742,N_4705);
xnor U4988 (N_4988,N_4616,N_4710);
or U4989 (N_4989,N_4751,N_4694);
nor U4990 (N_4990,N_4621,N_4748);
nand U4991 (N_4991,N_4711,N_4679);
nand U4992 (N_4992,N_4764,N_4713);
nand U4993 (N_4993,N_4601,N_4613);
xnor U4994 (N_4994,N_4741,N_4634);
and U4995 (N_4995,N_4714,N_4694);
nor U4996 (N_4996,N_4753,N_4768);
nand U4997 (N_4997,N_4732,N_4778);
or U4998 (N_4998,N_4760,N_4754);
or U4999 (N_4999,N_4666,N_4652);
nor U5000 (N_5000,N_4898,N_4843);
and U5001 (N_5001,N_4902,N_4861);
nand U5002 (N_5002,N_4872,N_4897);
nor U5003 (N_5003,N_4839,N_4914);
or U5004 (N_5004,N_4808,N_4908);
nand U5005 (N_5005,N_4998,N_4852);
xnor U5006 (N_5006,N_4821,N_4804);
xor U5007 (N_5007,N_4960,N_4833);
nand U5008 (N_5008,N_4819,N_4915);
xnor U5009 (N_5009,N_4928,N_4987);
and U5010 (N_5010,N_4857,N_4801);
nor U5011 (N_5011,N_4952,N_4965);
and U5012 (N_5012,N_4919,N_4936);
nor U5013 (N_5013,N_4943,N_4997);
and U5014 (N_5014,N_4812,N_4890);
or U5015 (N_5015,N_4920,N_4803);
nor U5016 (N_5016,N_4903,N_4967);
nand U5017 (N_5017,N_4962,N_4996);
nor U5018 (N_5018,N_4956,N_4961);
nand U5019 (N_5019,N_4873,N_4811);
xor U5020 (N_5020,N_4900,N_4989);
or U5021 (N_5021,N_4846,N_4863);
nor U5022 (N_5022,N_4932,N_4993);
xnor U5023 (N_5023,N_4854,N_4935);
and U5024 (N_5024,N_4830,N_4842);
nor U5025 (N_5025,N_4927,N_4972);
nor U5026 (N_5026,N_4921,N_4938);
and U5027 (N_5027,N_4939,N_4858);
and U5028 (N_5028,N_4866,N_4925);
or U5029 (N_5029,N_4879,N_4822);
and U5030 (N_5030,N_4845,N_4999);
nor U5031 (N_5031,N_4849,N_4886);
and U5032 (N_5032,N_4817,N_4901);
nand U5033 (N_5033,N_4869,N_4836);
nor U5034 (N_5034,N_4951,N_4966);
nor U5035 (N_5035,N_4992,N_4995);
and U5036 (N_5036,N_4815,N_4970);
and U5037 (N_5037,N_4916,N_4875);
nand U5038 (N_5038,N_4884,N_4802);
nor U5039 (N_5039,N_4885,N_4805);
nor U5040 (N_5040,N_4982,N_4899);
xnor U5041 (N_5041,N_4838,N_4953);
nand U5042 (N_5042,N_4933,N_4964);
nand U5043 (N_5043,N_4931,N_4963);
xnor U5044 (N_5044,N_4874,N_4904);
and U5045 (N_5045,N_4831,N_4926);
nor U5046 (N_5046,N_4945,N_4880);
xnor U5047 (N_5047,N_4823,N_4895);
and U5048 (N_5048,N_4971,N_4834);
xnor U5049 (N_5049,N_4813,N_4832);
xnor U5050 (N_5050,N_4950,N_4825);
and U5051 (N_5051,N_4855,N_4878);
nor U5052 (N_5052,N_4840,N_4969);
nor U5053 (N_5053,N_4824,N_4814);
xnor U5054 (N_5054,N_4923,N_4912);
xor U5055 (N_5055,N_4949,N_4918);
and U5056 (N_5056,N_4942,N_4922);
nand U5057 (N_5057,N_4841,N_4862);
or U5058 (N_5058,N_4975,N_4978);
nor U5059 (N_5059,N_4892,N_4958);
and U5060 (N_5060,N_4870,N_4907);
nor U5061 (N_5061,N_4959,N_4913);
xor U5062 (N_5062,N_4887,N_4976);
nor U5063 (N_5063,N_4979,N_4981);
nor U5064 (N_5064,N_4851,N_4957);
nor U5065 (N_5065,N_4827,N_4974);
nand U5066 (N_5066,N_4864,N_4818);
nor U5067 (N_5067,N_4948,N_4835);
and U5068 (N_5068,N_4844,N_4820);
nor U5069 (N_5069,N_4944,N_4882);
nand U5070 (N_5070,N_4889,N_4896);
or U5071 (N_5071,N_4980,N_4893);
and U5072 (N_5072,N_4946,N_4991);
or U5073 (N_5073,N_4837,N_4807);
xnor U5074 (N_5074,N_4865,N_4850);
or U5075 (N_5075,N_4881,N_4930);
nand U5076 (N_5076,N_4891,N_4806);
and U5077 (N_5077,N_4910,N_4909);
nor U5078 (N_5078,N_4941,N_4990);
nand U5079 (N_5079,N_4973,N_4934);
xnor U5080 (N_5080,N_4883,N_4917);
nand U5081 (N_5081,N_4947,N_4859);
or U5082 (N_5082,N_4955,N_4860);
or U5083 (N_5083,N_4826,N_4924);
or U5084 (N_5084,N_4829,N_4871);
nor U5085 (N_5085,N_4876,N_4929);
or U5086 (N_5086,N_4994,N_4856);
or U5087 (N_5087,N_4810,N_4868);
or U5088 (N_5088,N_4853,N_4867);
nand U5089 (N_5089,N_4937,N_4968);
nand U5090 (N_5090,N_4894,N_4816);
nand U5091 (N_5091,N_4984,N_4986);
and U5092 (N_5092,N_4977,N_4888);
nand U5093 (N_5093,N_4988,N_4847);
or U5094 (N_5094,N_4985,N_4877);
nor U5095 (N_5095,N_4906,N_4809);
nand U5096 (N_5096,N_4911,N_4954);
xnor U5097 (N_5097,N_4848,N_4983);
nor U5098 (N_5098,N_4940,N_4905);
nand U5099 (N_5099,N_4828,N_4800);
nand U5100 (N_5100,N_4862,N_4847);
nor U5101 (N_5101,N_4800,N_4879);
nor U5102 (N_5102,N_4858,N_4805);
nor U5103 (N_5103,N_4895,N_4955);
nor U5104 (N_5104,N_4999,N_4938);
or U5105 (N_5105,N_4934,N_4994);
nand U5106 (N_5106,N_4891,N_4834);
and U5107 (N_5107,N_4980,N_4885);
or U5108 (N_5108,N_4857,N_4905);
nor U5109 (N_5109,N_4962,N_4805);
xor U5110 (N_5110,N_4871,N_4956);
nand U5111 (N_5111,N_4843,N_4889);
nand U5112 (N_5112,N_4920,N_4937);
or U5113 (N_5113,N_4800,N_4802);
nor U5114 (N_5114,N_4836,N_4880);
or U5115 (N_5115,N_4821,N_4911);
nor U5116 (N_5116,N_4807,N_4987);
or U5117 (N_5117,N_4972,N_4928);
or U5118 (N_5118,N_4905,N_4864);
nand U5119 (N_5119,N_4816,N_4896);
nor U5120 (N_5120,N_4875,N_4818);
nand U5121 (N_5121,N_4804,N_4947);
and U5122 (N_5122,N_4828,N_4927);
and U5123 (N_5123,N_4829,N_4885);
or U5124 (N_5124,N_4813,N_4965);
nand U5125 (N_5125,N_4914,N_4976);
nor U5126 (N_5126,N_4926,N_4817);
or U5127 (N_5127,N_4856,N_4993);
and U5128 (N_5128,N_4882,N_4856);
nand U5129 (N_5129,N_4880,N_4944);
and U5130 (N_5130,N_4894,N_4900);
xnor U5131 (N_5131,N_4940,N_4871);
and U5132 (N_5132,N_4801,N_4930);
nand U5133 (N_5133,N_4840,N_4832);
nand U5134 (N_5134,N_4811,N_4877);
nand U5135 (N_5135,N_4883,N_4893);
nand U5136 (N_5136,N_4846,N_4952);
xnor U5137 (N_5137,N_4914,N_4896);
and U5138 (N_5138,N_4842,N_4884);
and U5139 (N_5139,N_4809,N_4862);
nor U5140 (N_5140,N_4895,N_4991);
and U5141 (N_5141,N_4888,N_4929);
nor U5142 (N_5142,N_4867,N_4932);
xor U5143 (N_5143,N_4945,N_4972);
xor U5144 (N_5144,N_4930,N_4871);
nor U5145 (N_5145,N_4808,N_4994);
and U5146 (N_5146,N_4814,N_4849);
and U5147 (N_5147,N_4997,N_4877);
xor U5148 (N_5148,N_4868,N_4841);
xor U5149 (N_5149,N_4875,N_4952);
nand U5150 (N_5150,N_4890,N_4836);
nor U5151 (N_5151,N_4879,N_4805);
nor U5152 (N_5152,N_4972,N_4935);
or U5153 (N_5153,N_4815,N_4913);
and U5154 (N_5154,N_4945,N_4814);
nor U5155 (N_5155,N_4850,N_4820);
or U5156 (N_5156,N_4965,N_4931);
or U5157 (N_5157,N_4957,N_4876);
nor U5158 (N_5158,N_4967,N_4966);
and U5159 (N_5159,N_4941,N_4879);
and U5160 (N_5160,N_4928,N_4800);
xor U5161 (N_5161,N_4889,N_4924);
or U5162 (N_5162,N_4990,N_4895);
nor U5163 (N_5163,N_4947,N_4871);
xor U5164 (N_5164,N_4934,N_4988);
and U5165 (N_5165,N_4819,N_4872);
and U5166 (N_5166,N_4992,N_4851);
and U5167 (N_5167,N_4912,N_4873);
nand U5168 (N_5168,N_4873,N_4901);
nor U5169 (N_5169,N_4966,N_4888);
or U5170 (N_5170,N_4949,N_4960);
or U5171 (N_5171,N_4862,N_4917);
xor U5172 (N_5172,N_4986,N_4995);
nor U5173 (N_5173,N_4999,N_4836);
xnor U5174 (N_5174,N_4823,N_4915);
xnor U5175 (N_5175,N_4983,N_4875);
or U5176 (N_5176,N_4922,N_4837);
nor U5177 (N_5177,N_4809,N_4859);
xnor U5178 (N_5178,N_4944,N_4940);
and U5179 (N_5179,N_4900,N_4924);
nor U5180 (N_5180,N_4880,N_4961);
and U5181 (N_5181,N_4940,N_4853);
and U5182 (N_5182,N_4877,N_4948);
nor U5183 (N_5183,N_4882,N_4982);
nand U5184 (N_5184,N_4801,N_4965);
xor U5185 (N_5185,N_4948,N_4853);
and U5186 (N_5186,N_4861,N_4933);
or U5187 (N_5187,N_4896,N_4907);
nor U5188 (N_5188,N_4982,N_4837);
nand U5189 (N_5189,N_4843,N_4833);
xor U5190 (N_5190,N_4914,N_4865);
nand U5191 (N_5191,N_4869,N_4831);
and U5192 (N_5192,N_4871,N_4963);
xor U5193 (N_5193,N_4848,N_4998);
xnor U5194 (N_5194,N_4803,N_4937);
or U5195 (N_5195,N_4939,N_4919);
or U5196 (N_5196,N_4928,N_4899);
nand U5197 (N_5197,N_4973,N_4971);
or U5198 (N_5198,N_4944,N_4904);
nand U5199 (N_5199,N_4818,N_4959);
or U5200 (N_5200,N_5072,N_5087);
and U5201 (N_5201,N_5076,N_5035);
xnor U5202 (N_5202,N_5181,N_5158);
xnor U5203 (N_5203,N_5125,N_5152);
nor U5204 (N_5204,N_5126,N_5095);
or U5205 (N_5205,N_5029,N_5056);
xnor U5206 (N_5206,N_5092,N_5044);
nand U5207 (N_5207,N_5010,N_5071);
xnor U5208 (N_5208,N_5077,N_5188);
and U5209 (N_5209,N_5175,N_5178);
and U5210 (N_5210,N_5047,N_5098);
nor U5211 (N_5211,N_5068,N_5094);
or U5212 (N_5212,N_5174,N_5101);
or U5213 (N_5213,N_5083,N_5136);
nand U5214 (N_5214,N_5189,N_5153);
xnor U5215 (N_5215,N_5194,N_5073);
nor U5216 (N_5216,N_5166,N_5046);
nor U5217 (N_5217,N_5084,N_5100);
nor U5218 (N_5218,N_5163,N_5172);
or U5219 (N_5219,N_5004,N_5130);
or U5220 (N_5220,N_5051,N_5021);
or U5221 (N_5221,N_5042,N_5161);
or U5222 (N_5222,N_5167,N_5013);
nor U5223 (N_5223,N_5064,N_5143);
and U5224 (N_5224,N_5054,N_5030);
nor U5225 (N_5225,N_5082,N_5150);
and U5226 (N_5226,N_5144,N_5198);
xor U5227 (N_5227,N_5184,N_5176);
nor U5228 (N_5228,N_5199,N_5055);
or U5229 (N_5229,N_5159,N_5052);
and U5230 (N_5230,N_5164,N_5061);
xnor U5231 (N_5231,N_5034,N_5156);
and U5232 (N_5232,N_5040,N_5187);
nand U5233 (N_5233,N_5093,N_5090);
nand U5234 (N_5234,N_5186,N_5131);
nand U5235 (N_5235,N_5036,N_5104);
xor U5236 (N_5236,N_5058,N_5160);
nand U5237 (N_5237,N_5171,N_5025);
nor U5238 (N_5238,N_5028,N_5041);
and U5239 (N_5239,N_5020,N_5197);
nand U5240 (N_5240,N_5140,N_5133);
and U5241 (N_5241,N_5124,N_5015);
or U5242 (N_5242,N_5147,N_5012);
nand U5243 (N_5243,N_5059,N_5107);
and U5244 (N_5244,N_5113,N_5078);
xnor U5245 (N_5245,N_5018,N_5129);
or U5246 (N_5246,N_5112,N_5118);
or U5247 (N_5247,N_5135,N_5066);
and U5248 (N_5248,N_5127,N_5099);
nand U5249 (N_5249,N_5193,N_5177);
nor U5250 (N_5250,N_5019,N_5116);
nor U5251 (N_5251,N_5070,N_5048);
and U5252 (N_5252,N_5173,N_5179);
xnor U5253 (N_5253,N_5085,N_5110);
xnor U5254 (N_5254,N_5023,N_5154);
or U5255 (N_5255,N_5043,N_5155);
nor U5256 (N_5256,N_5031,N_5109);
nor U5257 (N_5257,N_5192,N_5022);
nand U5258 (N_5258,N_5045,N_5011);
or U5259 (N_5259,N_5060,N_5102);
nand U5260 (N_5260,N_5111,N_5032);
or U5261 (N_5261,N_5014,N_5089);
nand U5262 (N_5262,N_5057,N_5017);
nand U5263 (N_5263,N_5065,N_5027);
xor U5264 (N_5264,N_5063,N_5117);
nor U5265 (N_5265,N_5086,N_5185);
xnor U5266 (N_5266,N_5141,N_5134);
xnor U5267 (N_5267,N_5038,N_5149);
nand U5268 (N_5268,N_5000,N_5145);
nor U5269 (N_5269,N_5132,N_5138);
nor U5270 (N_5270,N_5003,N_5050);
or U5271 (N_5271,N_5039,N_5142);
or U5272 (N_5272,N_5069,N_5123);
and U5273 (N_5273,N_5151,N_5079);
or U5274 (N_5274,N_5097,N_5075);
nand U5275 (N_5275,N_5006,N_5157);
nand U5276 (N_5276,N_5139,N_5062);
nand U5277 (N_5277,N_5080,N_5137);
nor U5278 (N_5278,N_5168,N_5180);
nor U5279 (N_5279,N_5119,N_5182);
or U5280 (N_5280,N_5091,N_5049);
nand U5281 (N_5281,N_5033,N_5148);
nand U5282 (N_5282,N_5191,N_5026);
nor U5283 (N_5283,N_5183,N_5165);
or U5284 (N_5284,N_5024,N_5016);
xor U5285 (N_5285,N_5001,N_5074);
xor U5286 (N_5286,N_5105,N_5190);
or U5287 (N_5287,N_5121,N_5128);
nor U5288 (N_5288,N_5005,N_5162);
and U5289 (N_5289,N_5103,N_5053);
or U5290 (N_5290,N_5002,N_5037);
xor U5291 (N_5291,N_5114,N_5108);
nor U5292 (N_5292,N_5170,N_5067);
or U5293 (N_5293,N_5096,N_5196);
xor U5294 (N_5294,N_5007,N_5009);
nor U5295 (N_5295,N_5195,N_5122);
and U5296 (N_5296,N_5088,N_5008);
xnor U5297 (N_5297,N_5081,N_5120);
xor U5298 (N_5298,N_5169,N_5106);
nor U5299 (N_5299,N_5146,N_5115);
or U5300 (N_5300,N_5140,N_5052);
xor U5301 (N_5301,N_5098,N_5001);
nand U5302 (N_5302,N_5003,N_5109);
and U5303 (N_5303,N_5036,N_5012);
nand U5304 (N_5304,N_5192,N_5140);
nand U5305 (N_5305,N_5029,N_5106);
nor U5306 (N_5306,N_5020,N_5102);
nand U5307 (N_5307,N_5089,N_5168);
or U5308 (N_5308,N_5073,N_5147);
nor U5309 (N_5309,N_5141,N_5158);
and U5310 (N_5310,N_5023,N_5056);
or U5311 (N_5311,N_5098,N_5159);
nand U5312 (N_5312,N_5060,N_5163);
xnor U5313 (N_5313,N_5146,N_5155);
and U5314 (N_5314,N_5092,N_5048);
nor U5315 (N_5315,N_5038,N_5159);
xnor U5316 (N_5316,N_5065,N_5080);
xnor U5317 (N_5317,N_5078,N_5068);
or U5318 (N_5318,N_5053,N_5157);
and U5319 (N_5319,N_5144,N_5091);
or U5320 (N_5320,N_5097,N_5009);
or U5321 (N_5321,N_5179,N_5140);
and U5322 (N_5322,N_5083,N_5125);
or U5323 (N_5323,N_5114,N_5045);
or U5324 (N_5324,N_5174,N_5079);
xnor U5325 (N_5325,N_5131,N_5184);
xnor U5326 (N_5326,N_5164,N_5024);
xnor U5327 (N_5327,N_5178,N_5069);
nor U5328 (N_5328,N_5085,N_5011);
or U5329 (N_5329,N_5108,N_5032);
xor U5330 (N_5330,N_5060,N_5027);
or U5331 (N_5331,N_5127,N_5124);
nand U5332 (N_5332,N_5004,N_5021);
xnor U5333 (N_5333,N_5013,N_5004);
or U5334 (N_5334,N_5185,N_5043);
nand U5335 (N_5335,N_5062,N_5069);
nand U5336 (N_5336,N_5191,N_5094);
nor U5337 (N_5337,N_5179,N_5141);
or U5338 (N_5338,N_5083,N_5067);
xor U5339 (N_5339,N_5134,N_5119);
or U5340 (N_5340,N_5134,N_5100);
nand U5341 (N_5341,N_5150,N_5054);
and U5342 (N_5342,N_5129,N_5069);
or U5343 (N_5343,N_5182,N_5029);
and U5344 (N_5344,N_5168,N_5031);
xnor U5345 (N_5345,N_5174,N_5140);
nor U5346 (N_5346,N_5124,N_5061);
nand U5347 (N_5347,N_5117,N_5179);
and U5348 (N_5348,N_5195,N_5147);
nand U5349 (N_5349,N_5133,N_5012);
xnor U5350 (N_5350,N_5016,N_5059);
or U5351 (N_5351,N_5199,N_5005);
or U5352 (N_5352,N_5040,N_5033);
xnor U5353 (N_5353,N_5177,N_5098);
nand U5354 (N_5354,N_5035,N_5119);
xor U5355 (N_5355,N_5093,N_5185);
and U5356 (N_5356,N_5082,N_5034);
xor U5357 (N_5357,N_5026,N_5001);
or U5358 (N_5358,N_5088,N_5054);
nand U5359 (N_5359,N_5149,N_5138);
nor U5360 (N_5360,N_5012,N_5193);
and U5361 (N_5361,N_5007,N_5044);
or U5362 (N_5362,N_5181,N_5189);
and U5363 (N_5363,N_5090,N_5184);
xnor U5364 (N_5364,N_5125,N_5105);
nand U5365 (N_5365,N_5142,N_5164);
nor U5366 (N_5366,N_5012,N_5186);
nor U5367 (N_5367,N_5189,N_5067);
nand U5368 (N_5368,N_5184,N_5189);
nor U5369 (N_5369,N_5048,N_5077);
nand U5370 (N_5370,N_5030,N_5094);
nand U5371 (N_5371,N_5115,N_5055);
or U5372 (N_5372,N_5010,N_5058);
and U5373 (N_5373,N_5195,N_5126);
nand U5374 (N_5374,N_5075,N_5167);
or U5375 (N_5375,N_5047,N_5086);
xor U5376 (N_5376,N_5117,N_5136);
nand U5377 (N_5377,N_5044,N_5079);
and U5378 (N_5378,N_5076,N_5185);
or U5379 (N_5379,N_5112,N_5028);
or U5380 (N_5380,N_5106,N_5055);
xnor U5381 (N_5381,N_5191,N_5131);
nand U5382 (N_5382,N_5012,N_5041);
or U5383 (N_5383,N_5053,N_5077);
nand U5384 (N_5384,N_5093,N_5033);
or U5385 (N_5385,N_5175,N_5086);
nand U5386 (N_5386,N_5064,N_5128);
nor U5387 (N_5387,N_5021,N_5108);
xor U5388 (N_5388,N_5185,N_5194);
or U5389 (N_5389,N_5163,N_5045);
nand U5390 (N_5390,N_5117,N_5195);
and U5391 (N_5391,N_5073,N_5040);
nand U5392 (N_5392,N_5185,N_5081);
and U5393 (N_5393,N_5129,N_5077);
or U5394 (N_5394,N_5091,N_5198);
nand U5395 (N_5395,N_5159,N_5197);
or U5396 (N_5396,N_5111,N_5134);
nand U5397 (N_5397,N_5099,N_5005);
and U5398 (N_5398,N_5051,N_5037);
xor U5399 (N_5399,N_5125,N_5078);
xor U5400 (N_5400,N_5266,N_5340);
xnor U5401 (N_5401,N_5344,N_5277);
and U5402 (N_5402,N_5238,N_5264);
or U5403 (N_5403,N_5318,N_5382);
xnor U5404 (N_5404,N_5254,N_5251);
and U5405 (N_5405,N_5365,N_5246);
and U5406 (N_5406,N_5351,N_5240);
nand U5407 (N_5407,N_5386,N_5262);
and U5408 (N_5408,N_5270,N_5215);
or U5409 (N_5409,N_5360,N_5212);
xnor U5410 (N_5410,N_5304,N_5338);
and U5411 (N_5411,N_5392,N_5265);
nand U5412 (N_5412,N_5204,N_5288);
nand U5413 (N_5413,N_5383,N_5397);
and U5414 (N_5414,N_5244,N_5203);
nor U5415 (N_5415,N_5243,N_5379);
and U5416 (N_5416,N_5259,N_5253);
nor U5417 (N_5417,N_5346,N_5358);
xnor U5418 (N_5418,N_5384,N_5209);
nand U5419 (N_5419,N_5333,N_5218);
nor U5420 (N_5420,N_5260,N_5242);
or U5421 (N_5421,N_5208,N_5343);
nor U5422 (N_5422,N_5322,N_5285);
nand U5423 (N_5423,N_5241,N_5380);
xor U5424 (N_5424,N_5257,N_5228);
nand U5425 (N_5425,N_5361,N_5237);
xor U5426 (N_5426,N_5387,N_5306);
xnor U5427 (N_5427,N_5357,N_5230);
nor U5428 (N_5428,N_5308,N_5388);
nand U5429 (N_5429,N_5309,N_5367);
or U5430 (N_5430,N_5349,N_5315);
xor U5431 (N_5431,N_5305,N_5341);
nand U5432 (N_5432,N_5289,N_5396);
nor U5433 (N_5433,N_5297,N_5345);
or U5434 (N_5434,N_5398,N_5200);
xnor U5435 (N_5435,N_5227,N_5281);
nor U5436 (N_5436,N_5219,N_5353);
nand U5437 (N_5437,N_5222,N_5295);
and U5438 (N_5438,N_5325,N_5332);
nor U5439 (N_5439,N_5236,N_5326);
xor U5440 (N_5440,N_5362,N_5279);
or U5441 (N_5441,N_5286,N_5255);
or U5442 (N_5442,N_5258,N_5275);
xnor U5443 (N_5443,N_5327,N_5231);
xnor U5444 (N_5444,N_5303,N_5378);
or U5445 (N_5445,N_5268,N_5370);
xor U5446 (N_5446,N_5296,N_5313);
or U5447 (N_5447,N_5377,N_5371);
and U5448 (N_5448,N_5336,N_5263);
xor U5449 (N_5449,N_5217,N_5252);
nor U5450 (N_5450,N_5324,N_5206);
xor U5451 (N_5451,N_5249,N_5293);
nand U5452 (N_5452,N_5368,N_5226);
nor U5453 (N_5453,N_5339,N_5271);
nor U5454 (N_5454,N_5359,N_5210);
and U5455 (N_5455,N_5393,N_5376);
nor U5456 (N_5456,N_5273,N_5356);
nor U5457 (N_5457,N_5261,N_5233);
xnor U5458 (N_5458,N_5350,N_5394);
and U5459 (N_5459,N_5330,N_5224);
xnor U5460 (N_5460,N_5355,N_5287);
xnor U5461 (N_5461,N_5267,N_5385);
nor U5462 (N_5462,N_5248,N_5232);
xor U5463 (N_5463,N_5395,N_5211);
xor U5464 (N_5464,N_5216,N_5334);
nor U5465 (N_5465,N_5373,N_5316);
nor U5466 (N_5466,N_5283,N_5284);
and U5467 (N_5467,N_5225,N_5202);
nor U5468 (N_5468,N_5301,N_5207);
nand U5469 (N_5469,N_5298,N_5302);
nor U5470 (N_5470,N_5369,N_5323);
or U5471 (N_5471,N_5229,N_5381);
xor U5472 (N_5472,N_5299,N_5352);
nand U5473 (N_5473,N_5310,N_5342);
nand U5474 (N_5474,N_5364,N_5213);
nand U5475 (N_5475,N_5366,N_5294);
or U5476 (N_5476,N_5329,N_5220);
nor U5477 (N_5477,N_5278,N_5239);
nor U5478 (N_5478,N_5221,N_5201);
or U5479 (N_5479,N_5347,N_5256);
xnor U5480 (N_5480,N_5245,N_5269);
nand U5481 (N_5481,N_5274,N_5312);
nand U5482 (N_5482,N_5290,N_5348);
nand U5483 (N_5483,N_5375,N_5363);
and U5484 (N_5484,N_5319,N_5300);
nor U5485 (N_5485,N_5399,N_5321);
xor U5486 (N_5486,N_5314,N_5205);
and U5487 (N_5487,N_5328,N_5292);
or U5488 (N_5488,N_5282,N_5331);
nand U5489 (N_5489,N_5235,N_5250);
or U5490 (N_5490,N_5354,N_5374);
and U5491 (N_5491,N_5389,N_5276);
nand U5492 (N_5492,N_5372,N_5320);
xnor U5493 (N_5493,N_5307,N_5214);
and U5494 (N_5494,N_5390,N_5291);
nand U5495 (N_5495,N_5391,N_5280);
nor U5496 (N_5496,N_5234,N_5317);
or U5497 (N_5497,N_5337,N_5335);
and U5498 (N_5498,N_5223,N_5247);
nor U5499 (N_5499,N_5311,N_5272);
xnor U5500 (N_5500,N_5361,N_5275);
nor U5501 (N_5501,N_5323,N_5383);
nor U5502 (N_5502,N_5337,N_5214);
xor U5503 (N_5503,N_5287,N_5399);
nand U5504 (N_5504,N_5336,N_5329);
xnor U5505 (N_5505,N_5236,N_5233);
and U5506 (N_5506,N_5230,N_5354);
and U5507 (N_5507,N_5366,N_5254);
nor U5508 (N_5508,N_5213,N_5261);
nor U5509 (N_5509,N_5398,N_5288);
xor U5510 (N_5510,N_5357,N_5202);
and U5511 (N_5511,N_5310,N_5279);
nand U5512 (N_5512,N_5338,N_5266);
xor U5513 (N_5513,N_5302,N_5237);
or U5514 (N_5514,N_5399,N_5380);
nand U5515 (N_5515,N_5373,N_5242);
nor U5516 (N_5516,N_5236,N_5293);
xor U5517 (N_5517,N_5308,N_5322);
nor U5518 (N_5518,N_5353,N_5259);
nand U5519 (N_5519,N_5382,N_5256);
and U5520 (N_5520,N_5316,N_5340);
xor U5521 (N_5521,N_5346,N_5233);
nand U5522 (N_5522,N_5361,N_5279);
or U5523 (N_5523,N_5246,N_5201);
nand U5524 (N_5524,N_5344,N_5260);
or U5525 (N_5525,N_5200,N_5332);
xor U5526 (N_5526,N_5399,N_5215);
nand U5527 (N_5527,N_5341,N_5396);
or U5528 (N_5528,N_5309,N_5218);
nand U5529 (N_5529,N_5328,N_5275);
or U5530 (N_5530,N_5281,N_5240);
and U5531 (N_5531,N_5384,N_5328);
nand U5532 (N_5532,N_5262,N_5339);
or U5533 (N_5533,N_5273,N_5247);
nor U5534 (N_5534,N_5221,N_5206);
xor U5535 (N_5535,N_5266,N_5364);
nor U5536 (N_5536,N_5284,N_5323);
nand U5537 (N_5537,N_5374,N_5385);
xor U5538 (N_5538,N_5264,N_5206);
and U5539 (N_5539,N_5387,N_5216);
and U5540 (N_5540,N_5245,N_5303);
and U5541 (N_5541,N_5360,N_5324);
and U5542 (N_5542,N_5248,N_5256);
xor U5543 (N_5543,N_5339,N_5276);
nor U5544 (N_5544,N_5244,N_5214);
nand U5545 (N_5545,N_5332,N_5217);
and U5546 (N_5546,N_5289,N_5379);
nand U5547 (N_5547,N_5232,N_5293);
xnor U5548 (N_5548,N_5212,N_5278);
nand U5549 (N_5549,N_5275,N_5207);
xor U5550 (N_5550,N_5201,N_5211);
or U5551 (N_5551,N_5380,N_5211);
nor U5552 (N_5552,N_5362,N_5380);
nor U5553 (N_5553,N_5223,N_5208);
xor U5554 (N_5554,N_5355,N_5248);
xnor U5555 (N_5555,N_5230,N_5367);
and U5556 (N_5556,N_5256,N_5200);
and U5557 (N_5557,N_5270,N_5373);
xor U5558 (N_5558,N_5233,N_5343);
xor U5559 (N_5559,N_5376,N_5375);
nand U5560 (N_5560,N_5371,N_5389);
nor U5561 (N_5561,N_5287,N_5278);
or U5562 (N_5562,N_5296,N_5376);
or U5563 (N_5563,N_5316,N_5384);
nor U5564 (N_5564,N_5235,N_5280);
nand U5565 (N_5565,N_5209,N_5369);
xor U5566 (N_5566,N_5217,N_5208);
xnor U5567 (N_5567,N_5353,N_5249);
xnor U5568 (N_5568,N_5268,N_5228);
nor U5569 (N_5569,N_5290,N_5272);
xor U5570 (N_5570,N_5235,N_5299);
nor U5571 (N_5571,N_5259,N_5332);
nand U5572 (N_5572,N_5309,N_5258);
nor U5573 (N_5573,N_5231,N_5260);
nor U5574 (N_5574,N_5368,N_5264);
and U5575 (N_5575,N_5249,N_5224);
or U5576 (N_5576,N_5352,N_5223);
nand U5577 (N_5577,N_5293,N_5317);
nand U5578 (N_5578,N_5213,N_5349);
xnor U5579 (N_5579,N_5375,N_5275);
and U5580 (N_5580,N_5231,N_5265);
or U5581 (N_5581,N_5292,N_5327);
nor U5582 (N_5582,N_5287,N_5281);
nor U5583 (N_5583,N_5216,N_5374);
and U5584 (N_5584,N_5204,N_5265);
nand U5585 (N_5585,N_5242,N_5270);
xnor U5586 (N_5586,N_5329,N_5287);
xnor U5587 (N_5587,N_5393,N_5245);
xnor U5588 (N_5588,N_5205,N_5352);
and U5589 (N_5589,N_5223,N_5305);
nand U5590 (N_5590,N_5393,N_5261);
nor U5591 (N_5591,N_5203,N_5218);
nor U5592 (N_5592,N_5330,N_5286);
and U5593 (N_5593,N_5224,N_5386);
xor U5594 (N_5594,N_5373,N_5362);
nand U5595 (N_5595,N_5233,N_5272);
and U5596 (N_5596,N_5388,N_5324);
nor U5597 (N_5597,N_5246,N_5304);
and U5598 (N_5598,N_5220,N_5399);
xnor U5599 (N_5599,N_5328,N_5364);
or U5600 (N_5600,N_5542,N_5587);
and U5601 (N_5601,N_5570,N_5411);
or U5602 (N_5602,N_5592,N_5585);
xor U5603 (N_5603,N_5433,N_5599);
nand U5604 (N_5604,N_5458,N_5418);
xnor U5605 (N_5605,N_5593,N_5461);
nor U5606 (N_5606,N_5424,N_5510);
nand U5607 (N_5607,N_5466,N_5590);
nor U5608 (N_5608,N_5423,N_5499);
nand U5609 (N_5609,N_5505,N_5576);
and U5610 (N_5610,N_5457,N_5583);
or U5611 (N_5611,N_5470,N_5415);
nand U5612 (N_5612,N_5496,N_5462);
xnor U5613 (N_5613,N_5494,N_5555);
xnor U5614 (N_5614,N_5440,N_5572);
or U5615 (N_5615,N_5547,N_5492);
nor U5616 (N_5616,N_5454,N_5552);
xnor U5617 (N_5617,N_5586,N_5422);
nor U5618 (N_5618,N_5459,N_5589);
or U5619 (N_5619,N_5482,N_5568);
nor U5620 (N_5620,N_5513,N_5571);
xnor U5621 (N_5621,N_5420,N_5404);
nand U5622 (N_5622,N_5524,N_5400);
and U5623 (N_5623,N_5408,N_5535);
or U5624 (N_5624,N_5497,N_5532);
nand U5625 (N_5625,N_5591,N_5453);
and U5626 (N_5626,N_5543,N_5429);
nand U5627 (N_5627,N_5435,N_5443);
or U5628 (N_5628,N_5598,N_5569);
and U5629 (N_5629,N_5538,N_5525);
nor U5630 (N_5630,N_5448,N_5486);
nand U5631 (N_5631,N_5413,N_5563);
and U5632 (N_5632,N_5437,N_5527);
xor U5633 (N_5633,N_5485,N_5476);
or U5634 (N_5634,N_5551,N_5446);
and U5635 (N_5635,N_5562,N_5530);
xor U5636 (N_5636,N_5444,N_5516);
and U5637 (N_5637,N_5417,N_5447);
nand U5638 (N_5638,N_5480,N_5521);
nor U5639 (N_5639,N_5549,N_5465);
xor U5640 (N_5640,N_5469,N_5577);
or U5641 (N_5641,N_5534,N_5581);
xnor U5642 (N_5642,N_5506,N_5456);
nand U5643 (N_5643,N_5401,N_5550);
nor U5644 (N_5644,N_5537,N_5464);
nand U5645 (N_5645,N_5436,N_5483);
nor U5646 (N_5646,N_5545,N_5514);
nor U5647 (N_5647,N_5427,N_5451);
and U5648 (N_5648,N_5430,N_5402);
nand U5649 (N_5649,N_5553,N_5502);
and U5650 (N_5650,N_5426,N_5428);
and U5651 (N_5651,N_5495,N_5479);
or U5652 (N_5652,N_5475,N_5491);
and U5653 (N_5653,N_5529,N_5425);
xnor U5654 (N_5654,N_5564,N_5452);
or U5655 (N_5655,N_5540,N_5438);
nor U5656 (N_5656,N_5582,N_5539);
xnor U5657 (N_5657,N_5442,N_5504);
and U5658 (N_5658,N_5518,N_5445);
and U5659 (N_5659,N_5507,N_5519);
or U5660 (N_5660,N_5431,N_5487);
nor U5661 (N_5661,N_5471,N_5403);
xnor U5662 (N_5662,N_5575,N_5477);
xor U5663 (N_5663,N_5500,N_5544);
nand U5664 (N_5664,N_5449,N_5512);
nand U5665 (N_5665,N_5574,N_5548);
xnor U5666 (N_5666,N_5405,N_5509);
xor U5667 (N_5667,N_5455,N_5488);
or U5668 (N_5668,N_5501,N_5450);
or U5669 (N_5669,N_5467,N_5580);
xor U5670 (N_5670,N_5434,N_5517);
and U5671 (N_5671,N_5409,N_5493);
nor U5672 (N_5672,N_5566,N_5594);
and U5673 (N_5673,N_5416,N_5490);
xnor U5674 (N_5674,N_5561,N_5565);
nand U5675 (N_5675,N_5556,N_5460);
and U5676 (N_5676,N_5573,N_5498);
or U5677 (N_5677,N_5414,N_5546);
and U5678 (N_5678,N_5441,N_5503);
or U5679 (N_5679,N_5515,N_5523);
nand U5680 (N_5680,N_5520,N_5421);
nand U5681 (N_5681,N_5541,N_5588);
or U5682 (N_5682,N_5463,N_5474);
nor U5683 (N_5683,N_5522,N_5419);
xnor U5684 (N_5684,N_5597,N_5558);
xor U5685 (N_5685,N_5406,N_5478);
or U5686 (N_5686,N_5410,N_5439);
nor U5687 (N_5687,N_5508,N_5489);
or U5688 (N_5688,N_5468,N_5536);
and U5689 (N_5689,N_5567,N_5579);
xnor U5690 (N_5690,N_5528,N_5596);
or U5691 (N_5691,N_5511,N_5559);
nand U5692 (N_5692,N_5526,N_5595);
xnor U5693 (N_5693,N_5432,N_5531);
or U5694 (N_5694,N_5407,N_5484);
or U5695 (N_5695,N_5481,N_5560);
or U5696 (N_5696,N_5578,N_5473);
and U5697 (N_5697,N_5533,N_5554);
xor U5698 (N_5698,N_5584,N_5412);
nand U5699 (N_5699,N_5472,N_5557);
nor U5700 (N_5700,N_5560,N_5492);
or U5701 (N_5701,N_5422,N_5552);
xor U5702 (N_5702,N_5574,N_5472);
nand U5703 (N_5703,N_5484,N_5429);
nand U5704 (N_5704,N_5423,N_5453);
xnor U5705 (N_5705,N_5483,N_5443);
nor U5706 (N_5706,N_5568,N_5584);
nor U5707 (N_5707,N_5431,N_5566);
xnor U5708 (N_5708,N_5588,N_5534);
xnor U5709 (N_5709,N_5530,N_5434);
nand U5710 (N_5710,N_5473,N_5504);
nor U5711 (N_5711,N_5452,N_5532);
and U5712 (N_5712,N_5441,N_5554);
nand U5713 (N_5713,N_5542,N_5515);
and U5714 (N_5714,N_5493,N_5584);
or U5715 (N_5715,N_5452,N_5590);
or U5716 (N_5716,N_5538,N_5474);
nor U5717 (N_5717,N_5461,N_5408);
or U5718 (N_5718,N_5521,N_5598);
nor U5719 (N_5719,N_5571,N_5495);
and U5720 (N_5720,N_5576,N_5515);
and U5721 (N_5721,N_5593,N_5590);
and U5722 (N_5722,N_5455,N_5559);
nand U5723 (N_5723,N_5479,N_5461);
nand U5724 (N_5724,N_5422,N_5580);
and U5725 (N_5725,N_5458,N_5570);
nor U5726 (N_5726,N_5450,N_5429);
and U5727 (N_5727,N_5509,N_5450);
nand U5728 (N_5728,N_5434,N_5482);
xnor U5729 (N_5729,N_5506,N_5541);
or U5730 (N_5730,N_5506,N_5507);
and U5731 (N_5731,N_5403,N_5542);
and U5732 (N_5732,N_5441,N_5488);
nand U5733 (N_5733,N_5495,N_5551);
or U5734 (N_5734,N_5425,N_5489);
nand U5735 (N_5735,N_5481,N_5446);
and U5736 (N_5736,N_5522,N_5430);
nor U5737 (N_5737,N_5484,N_5543);
and U5738 (N_5738,N_5569,N_5431);
nand U5739 (N_5739,N_5531,N_5573);
or U5740 (N_5740,N_5420,N_5434);
or U5741 (N_5741,N_5401,N_5434);
and U5742 (N_5742,N_5520,N_5549);
xnor U5743 (N_5743,N_5558,N_5462);
nand U5744 (N_5744,N_5450,N_5589);
and U5745 (N_5745,N_5488,N_5511);
xnor U5746 (N_5746,N_5524,N_5456);
nand U5747 (N_5747,N_5472,N_5532);
or U5748 (N_5748,N_5483,N_5404);
and U5749 (N_5749,N_5594,N_5584);
and U5750 (N_5750,N_5423,N_5434);
and U5751 (N_5751,N_5561,N_5443);
and U5752 (N_5752,N_5504,N_5491);
xnor U5753 (N_5753,N_5530,N_5511);
xnor U5754 (N_5754,N_5417,N_5550);
or U5755 (N_5755,N_5414,N_5458);
xor U5756 (N_5756,N_5436,N_5597);
xnor U5757 (N_5757,N_5534,N_5591);
nand U5758 (N_5758,N_5584,N_5471);
xor U5759 (N_5759,N_5597,N_5487);
or U5760 (N_5760,N_5480,N_5418);
xnor U5761 (N_5761,N_5465,N_5441);
nor U5762 (N_5762,N_5431,N_5599);
xor U5763 (N_5763,N_5472,N_5567);
nor U5764 (N_5764,N_5591,N_5588);
nand U5765 (N_5765,N_5573,N_5439);
or U5766 (N_5766,N_5429,N_5550);
xnor U5767 (N_5767,N_5540,N_5445);
xnor U5768 (N_5768,N_5564,N_5412);
or U5769 (N_5769,N_5456,N_5491);
nand U5770 (N_5770,N_5575,N_5536);
xnor U5771 (N_5771,N_5512,N_5403);
and U5772 (N_5772,N_5422,N_5519);
and U5773 (N_5773,N_5537,N_5482);
nor U5774 (N_5774,N_5487,N_5589);
nand U5775 (N_5775,N_5485,N_5462);
and U5776 (N_5776,N_5599,N_5539);
nor U5777 (N_5777,N_5419,N_5578);
xor U5778 (N_5778,N_5526,N_5499);
xnor U5779 (N_5779,N_5538,N_5492);
or U5780 (N_5780,N_5572,N_5506);
xor U5781 (N_5781,N_5585,N_5440);
nor U5782 (N_5782,N_5479,N_5521);
nor U5783 (N_5783,N_5443,N_5517);
nor U5784 (N_5784,N_5535,N_5570);
nor U5785 (N_5785,N_5574,N_5537);
and U5786 (N_5786,N_5593,N_5429);
and U5787 (N_5787,N_5461,N_5456);
nand U5788 (N_5788,N_5457,N_5472);
xnor U5789 (N_5789,N_5463,N_5519);
xnor U5790 (N_5790,N_5514,N_5456);
nor U5791 (N_5791,N_5459,N_5405);
and U5792 (N_5792,N_5445,N_5568);
and U5793 (N_5793,N_5504,N_5597);
nor U5794 (N_5794,N_5484,N_5533);
nor U5795 (N_5795,N_5442,N_5495);
xnor U5796 (N_5796,N_5423,N_5540);
nor U5797 (N_5797,N_5594,N_5576);
nand U5798 (N_5798,N_5574,N_5463);
xnor U5799 (N_5799,N_5503,N_5535);
or U5800 (N_5800,N_5706,N_5713);
xnor U5801 (N_5801,N_5744,N_5679);
nor U5802 (N_5802,N_5761,N_5703);
nor U5803 (N_5803,N_5776,N_5632);
or U5804 (N_5804,N_5664,N_5652);
nor U5805 (N_5805,N_5638,N_5611);
nand U5806 (N_5806,N_5773,N_5667);
and U5807 (N_5807,N_5672,N_5648);
xnor U5808 (N_5808,N_5689,N_5657);
nor U5809 (N_5809,N_5688,N_5740);
nand U5810 (N_5810,N_5647,N_5791);
xor U5811 (N_5811,N_5694,N_5747);
xnor U5812 (N_5812,N_5784,N_5691);
nor U5813 (N_5813,N_5675,N_5643);
nand U5814 (N_5814,N_5602,N_5697);
and U5815 (N_5815,N_5721,N_5790);
nand U5816 (N_5816,N_5777,N_5645);
nor U5817 (N_5817,N_5624,N_5685);
or U5818 (N_5818,N_5686,N_5771);
nand U5819 (N_5819,N_5782,N_5764);
nand U5820 (N_5820,N_5725,N_5753);
and U5821 (N_5821,N_5738,N_5717);
or U5822 (N_5822,N_5662,N_5795);
or U5823 (N_5823,N_5718,N_5609);
nand U5824 (N_5824,N_5620,N_5627);
nor U5825 (N_5825,N_5799,N_5653);
and U5826 (N_5826,N_5702,N_5716);
and U5827 (N_5827,N_5607,N_5678);
xor U5828 (N_5828,N_5644,N_5655);
nor U5829 (N_5829,N_5749,N_5637);
or U5830 (N_5830,N_5666,N_5646);
and U5831 (N_5831,N_5714,N_5635);
xor U5832 (N_5832,N_5668,N_5735);
or U5833 (N_5833,N_5612,N_5732);
and U5834 (N_5834,N_5755,N_5733);
nand U5835 (N_5835,N_5621,N_5654);
or U5836 (N_5836,N_5700,N_5701);
nand U5837 (N_5837,N_5629,N_5683);
nand U5838 (N_5838,N_5628,N_5673);
and U5839 (N_5839,N_5677,N_5766);
nand U5840 (N_5840,N_5695,N_5727);
nor U5841 (N_5841,N_5658,N_5669);
nand U5842 (N_5842,N_5734,N_5785);
nor U5843 (N_5843,N_5670,N_5601);
or U5844 (N_5844,N_5661,N_5796);
xor U5845 (N_5845,N_5606,N_5754);
or U5846 (N_5846,N_5699,N_5786);
or U5847 (N_5847,N_5715,N_5711);
nand U5848 (N_5848,N_5680,N_5650);
nand U5849 (N_5849,N_5600,N_5640);
or U5850 (N_5850,N_5710,N_5639);
or U5851 (N_5851,N_5617,N_5719);
xor U5852 (N_5852,N_5704,N_5765);
or U5853 (N_5853,N_5760,N_5724);
and U5854 (N_5854,N_5613,N_5615);
nand U5855 (N_5855,N_5729,N_5758);
nor U5856 (N_5856,N_5745,N_5698);
and U5857 (N_5857,N_5723,N_5748);
or U5858 (N_5858,N_5618,N_5780);
nor U5859 (N_5859,N_5625,N_5610);
and U5860 (N_5860,N_5737,N_5696);
or U5861 (N_5861,N_5622,N_5779);
nand U5862 (N_5862,N_5731,N_5775);
nand U5863 (N_5863,N_5788,N_5756);
xnor U5864 (N_5864,N_5787,N_5619);
xor U5865 (N_5865,N_5705,N_5726);
or U5866 (N_5866,N_5623,N_5739);
or U5867 (N_5867,N_5752,N_5708);
xnor U5868 (N_5868,N_5692,N_5722);
xor U5869 (N_5869,N_5743,N_5649);
nor U5870 (N_5870,N_5730,N_5789);
nand U5871 (N_5871,N_5665,N_5736);
nor U5872 (N_5872,N_5608,N_5651);
nor U5873 (N_5873,N_5690,N_5772);
and U5874 (N_5874,N_5742,N_5720);
nor U5875 (N_5875,N_5741,N_5728);
nor U5876 (N_5876,N_5757,N_5793);
xor U5877 (N_5877,N_5783,N_5631);
nor U5878 (N_5878,N_5656,N_5634);
or U5879 (N_5879,N_5794,N_5687);
or U5880 (N_5880,N_5759,N_5674);
nand U5881 (N_5881,N_5636,N_5709);
nand U5882 (N_5882,N_5605,N_5642);
nor U5883 (N_5883,N_5676,N_5778);
nor U5884 (N_5884,N_5750,N_5770);
and U5885 (N_5885,N_5659,N_5751);
nor U5886 (N_5886,N_5707,N_5663);
and U5887 (N_5887,N_5660,N_5626);
or U5888 (N_5888,N_5671,N_5693);
nor U5889 (N_5889,N_5767,N_5603);
and U5890 (N_5890,N_5762,N_5616);
nor U5891 (N_5891,N_5682,N_5768);
xor U5892 (N_5892,N_5774,N_5763);
nand U5893 (N_5893,N_5781,N_5712);
or U5894 (N_5894,N_5769,N_5684);
and U5895 (N_5895,N_5681,N_5746);
and U5896 (N_5896,N_5792,N_5798);
and U5897 (N_5897,N_5630,N_5641);
nand U5898 (N_5898,N_5633,N_5614);
and U5899 (N_5899,N_5604,N_5797);
xor U5900 (N_5900,N_5758,N_5740);
nor U5901 (N_5901,N_5696,N_5710);
and U5902 (N_5902,N_5610,N_5696);
nor U5903 (N_5903,N_5674,N_5726);
and U5904 (N_5904,N_5765,N_5783);
and U5905 (N_5905,N_5766,N_5628);
nor U5906 (N_5906,N_5610,N_5619);
xor U5907 (N_5907,N_5742,N_5645);
nand U5908 (N_5908,N_5799,N_5763);
xor U5909 (N_5909,N_5720,N_5692);
or U5910 (N_5910,N_5651,N_5786);
and U5911 (N_5911,N_5756,N_5799);
nand U5912 (N_5912,N_5658,N_5793);
nand U5913 (N_5913,N_5611,N_5736);
nand U5914 (N_5914,N_5744,N_5772);
xnor U5915 (N_5915,N_5658,N_5764);
or U5916 (N_5916,N_5795,N_5622);
and U5917 (N_5917,N_5631,N_5695);
nand U5918 (N_5918,N_5661,N_5625);
and U5919 (N_5919,N_5702,N_5654);
and U5920 (N_5920,N_5704,N_5678);
nor U5921 (N_5921,N_5741,N_5795);
or U5922 (N_5922,N_5646,N_5708);
or U5923 (N_5923,N_5646,N_5706);
nor U5924 (N_5924,N_5661,N_5609);
and U5925 (N_5925,N_5698,N_5728);
and U5926 (N_5926,N_5709,N_5726);
xnor U5927 (N_5927,N_5618,N_5684);
or U5928 (N_5928,N_5766,N_5673);
nand U5929 (N_5929,N_5784,N_5664);
xor U5930 (N_5930,N_5641,N_5752);
xnor U5931 (N_5931,N_5780,N_5612);
nor U5932 (N_5932,N_5796,N_5731);
nor U5933 (N_5933,N_5689,N_5667);
nand U5934 (N_5934,N_5671,N_5610);
nor U5935 (N_5935,N_5670,N_5721);
xnor U5936 (N_5936,N_5601,N_5754);
nand U5937 (N_5937,N_5772,N_5767);
nand U5938 (N_5938,N_5706,N_5622);
and U5939 (N_5939,N_5776,N_5649);
nor U5940 (N_5940,N_5799,N_5636);
or U5941 (N_5941,N_5617,N_5670);
nand U5942 (N_5942,N_5638,N_5762);
nor U5943 (N_5943,N_5792,N_5661);
nand U5944 (N_5944,N_5715,N_5663);
nor U5945 (N_5945,N_5608,N_5658);
and U5946 (N_5946,N_5606,N_5727);
or U5947 (N_5947,N_5626,N_5739);
xor U5948 (N_5948,N_5652,N_5635);
and U5949 (N_5949,N_5623,N_5744);
or U5950 (N_5950,N_5685,N_5715);
nor U5951 (N_5951,N_5786,N_5640);
or U5952 (N_5952,N_5634,N_5755);
nor U5953 (N_5953,N_5686,N_5710);
and U5954 (N_5954,N_5640,N_5799);
xor U5955 (N_5955,N_5748,N_5648);
or U5956 (N_5956,N_5749,N_5702);
xnor U5957 (N_5957,N_5708,N_5642);
nand U5958 (N_5958,N_5772,N_5628);
or U5959 (N_5959,N_5721,N_5632);
or U5960 (N_5960,N_5780,N_5729);
or U5961 (N_5961,N_5733,N_5608);
and U5962 (N_5962,N_5716,N_5725);
xnor U5963 (N_5963,N_5604,N_5714);
xnor U5964 (N_5964,N_5689,N_5770);
xor U5965 (N_5965,N_5651,N_5739);
nand U5966 (N_5966,N_5774,N_5715);
and U5967 (N_5967,N_5745,N_5660);
nor U5968 (N_5968,N_5615,N_5605);
and U5969 (N_5969,N_5657,N_5736);
nor U5970 (N_5970,N_5696,N_5607);
nand U5971 (N_5971,N_5725,N_5693);
and U5972 (N_5972,N_5614,N_5609);
and U5973 (N_5973,N_5718,N_5613);
nor U5974 (N_5974,N_5606,N_5789);
nand U5975 (N_5975,N_5633,N_5737);
or U5976 (N_5976,N_5783,N_5640);
nand U5977 (N_5977,N_5720,N_5724);
and U5978 (N_5978,N_5657,N_5667);
xor U5979 (N_5979,N_5642,N_5600);
nor U5980 (N_5980,N_5689,N_5729);
nand U5981 (N_5981,N_5717,N_5609);
nor U5982 (N_5982,N_5669,N_5784);
xnor U5983 (N_5983,N_5783,N_5787);
xor U5984 (N_5984,N_5740,N_5767);
nor U5985 (N_5985,N_5634,N_5603);
xnor U5986 (N_5986,N_5679,N_5620);
nand U5987 (N_5987,N_5644,N_5670);
nor U5988 (N_5988,N_5650,N_5716);
xnor U5989 (N_5989,N_5791,N_5786);
xnor U5990 (N_5990,N_5647,N_5764);
and U5991 (N_5991,N_5650,N_5666);
nand U5992 (N_5992,N_5778,N_5660);
xor U5993 (N_5993,N_5778,N_5663);
nor U5994 (N_5994,N_5674,N_5615);
nand U5995 (N_5995,N_5639,N_5752);
or U5996 (N_5996,N_5624,N_5732);
or U5997 (N_5997,N_5691,N_5602);
nand U5998 (N_5998,N_5701,N_5613);
xor U5999 (N_5999,N_5785,N_5629);
nand U6000 (N_6000,N_5933,N_5847);
and U6001 (N_6001,N_5875,N_5824);
nor U6002 (N_6002,N_5894,N_5817);
nand U6003 (N_6003,N_5845,N_5970);
and U6004 (N_6004,N_5995,N_5890);
nand U6005 (N_6005,N_5803,N_5978);
or U6006 (N_6006,N_5841,N_5974);
and U6007 (N_6007,N_5812,N_5886);
or U6008 (N_6008,N_5919,N_5951);
nand U6009 (N_6009,N_5932,N_5916);
nor U6010 (N_6010,N_5975,N_5858);
and U6011 (N_6011,N_5800,N_5848);
nor U6012 (N_6012,N_5898,N_5866);
nand U6013 (N_6013,N_5954,N_5820);
and U6014 (N_6014,N_5815,N_5996);
nand U6015 (N_6015,N_5952,N_5833);
and U6016 (N_6016,N_5998,N_5994);
nor U6017 (N_6017,N_5910,N_5992);
xnor U6018 (N_6018,N_5895,N_5999);
xnor U6019 (N_6019,N_5826,N_5868);
nand U6020 (N_6020,N_5942,N_5948);
xnor U6021 (N_6021,N_5968,N_5984);
and U6022 (N_6022,N_5944,N_5806);
nor U6023 (N_6023,N_5973,N_5947);
nor U6024 (N_6024,N_5828,N_5901);
xnor U6025 (N_6025,N_5878,N_5856);
nor U6026 (N_6026,N_5989,N_5849);
nor U6027 (N_6027,N_5936,N_5854);
and U6028 (N_6028,N_5956,N_5962);
xor U6029 (N_6029,N_5872,N_5804);
or U6030 (N_6030,N_5988,N_5870);
xnor U6031 (N_6031,N_5809,N_5887);
and U6032 (N_6032,N_5885,N_5949);
nand U6033 (N_6033,N_5853,N_5939);
xor U6034 (N_6034,N_5850,N_5959);
or U6035 (N_6035,N_5857,N_5801);
nor U6036 (N_6036,N_5917,N_5938);
or U6037 (N_6037,N_5943,N_5888);
nand U6038 (N_6038,N_5863,N_5982);
nor U6039 (N_6039,N_5909,N_5834);
nor U6040 (N_6040,N_5813,N_5843);
xor U6041 (N_6041,N_5925,N_5964);
or U6042 (N_6042,N_5867,N_5810);
and U6043 (N_6043,N_5979,N_5805);
and U6044 (N_6044,N_5908,N_5922);
or U6045 (N_6045,N_5915,N_5980);
xor U6046 (N_6046,N_5827,N_5913);
xnor U6047 (N_6047,N_5929,N_5906);
and U6048 (N_6048,N_5821,N_5957);
xnor U6049 (N_6049,N_5941,N_5958);
xor U6050 (N_6050,N_5946,N_5864);
xnor U6051 (N_6051,N_5865,N_5883);
xnor U6052 (N_6052,N_5969,N_5912);
nor U6053 (N_6053,N_5884,N_5977);
nor U6054 (N_6054,N_5926,N_5940);
xor U6055 (N_6055,N_5823,N_5816);
nor U6056 (N_6056,N_5971,N_5839);
nor U6057 (N_6057,N_5923,N_5904);
nor U6058 (N_6058,N_5993,N_5931);
nand U6059 (N_6059,N_5880,N_5986);
xnor U6060 (N_6060,N_5882,N_5963);
xor U6061 (N_6061,N_5921,N_5950);
nand U6062 (N_6062,N_5881,N_5877);
and U6063 (N_6063,N_5937,N_5935);
nand U6064 (N_6064,N_5830,N_5892);
xnor U6065 (N_6065,N_5920,N_5891);
and U6066 (N_6066,N_5889,N_5972);
or U6067 (N_6067,N_5822,N_5897);
or U6068 (N_6068,N_5837,N_5852);
or U6069 (N_6069,N_5814,N_5918);
xor U6070 (N_6070,N_5967,N_5893);
or U6071 (N_6071,N_5905,N_5914);
and U6072 (N_6072,N_5871,N_5840);
nor U6073 (N_6073,N_5819,N_5842);
nand U6074 (N_6074,N_5945,N_5965);
xor U6075 (N_6075,N_5874,N_5927);
xnor U6076 (N_6076,N_5844,N_5900);
xnor U6077 (N_6077,N_5807,N_5808);
nand U6078 (N_6078,N_5879,N_5896);
nand U6079 (N_6079,N_5860,N_5832);
nor U6080 (N_6080,N_5831,N_5835);
xor U6081 (N_6081,N_5987,N_5990);
or U6082 (N_6082,N_5859,N_5869);
nor U6083 (N_6083,N_5818,N_5846);
or U6084 (N_6084,N_5873,N_5924);
xor U6085 (N_6085,N_5934,N_5911);
or U6086 (N_6086,N_5907,N_5961);
or U6087 (N_6087,N_5829,N_5966);
and U6088 (N_6088,N_5930,N_5811);
or U6089 (N_6089,N_5928,N_5802);
nor U6090 (N_6090,N_5855,N_5960);
xor U6091 (N_6091,N_5981,N_5876);
nand U6092 (N_6092,N_5899,N_5862);
nand U6093 (N_6093,N_5902,N_5851);
nor U6094 (N_6094,N_5991,N_5983);
xnor U6095 (N_6095,N_5861,N_5836);
nor U6096 (N_6096,N_5985,N_5953);
xnor U6097 (N_6097,N_5997,N_5955);
or U6098 (N_6098,N_5976,N_5838);
xor U6099 (N_6099,N_5825,N_5903);
or U6100 (N_6100,N_5820,N_5936);
or U6101 (N_6101,N_5842,N_5811);
or U6102 (N_6102,N_5968,N_5898);
or U6103 (N_6103,N_5998,N_5907);
nor U6104 (N_6104,N_5841,N_5860);
nand U6105 (N_6105,N_5837,N_5871);
nand U6106 (N_6106,N_5909,N_5940);
nor U6107 (N_6107,N_5868,N_5931);
xnor U6108 (N_6108,N_5841,N_5844);
and U6109 (N_6109,N_5901,N_5941);
xnor U6110 (N_6110,N_5843,N_5887);
xnor U6111 (N_6111,N_5864,N_5964);
or U6112 (N_6112,N_5870,N_5805);
or U6113 (N_6113,N_5979,N_5947);
nand U6114 (N_6114,N_5881,N_5906);
xnor U6115 (N_6115,N_5804,N_5803);
or U6116 (N_6116,N_5872,N_5809);
nand U6117 (N_6117,N_5832,N_5988);
nor U6118 (N_6118,N_5894,N_5971);
xnor U6119 (N_6119,N_5895,N_5890);
or U6120 (N_6120,N_5892,N_5863);
or U6121 (N_6121,N_5833,N_5891);
nor U6122 (N_6122,N_5827,N_5814);
nor U6123 (N_6123,N_5994,N_5824);
nor U6124 (N_6124,N_5836,N_5936);
nand U6125 (N_6125,N_5991,N_5934);
nand U6126 (N_6126,N_5819,N_5826);
and U6127 (N_6127,N_5870,N_5994);
and U6128 (N_6128,N_5837,N_5818);
or U6129 (N_6129,N_5805,N_5885);
nand U6130 (N_6130,N_5876,N_5869);
xnor U6131 (N_6131,N_5957,N_5824);
xnor U6132 (N_6132,N_5967,N_5830);
or U6133 (N_6133,N_5904,N_5837);
or U6134 (N_6134,N_5881,N_5987);
or U6135 (N_6135,N_5876,N_5810);
xor U6136 (N_6136,N_5907,N_5895);
and U6137 (N_6137,N_5916,N_5984);
and U6138 (N_6138,N_5948,N_5981);
xnor U6139 (N_6139,N_5942,N_5826);
and U6140 (N_6140,N_5922,N_5966);
or U6141 (N_6141,N_5899,N_5986);
nand U6142 (N_6142,N_5999,N_5927);
or U6143 (N_6143,N_5983,N_5807);
nand U6144 (N_6144,N_5884,N_5808);
nand U6145 (N_6145,N_5937,N_5992);
or U6146 (N_6146,N_5928,N_5867);
nand U6147 (N_6147,N_5926,N_5955);
and U6148 (N_6148,N_5904,N_5888);
or U6149 (N_6149,N_5844,N_5920);
nor U6150 (N_6150,N_5980,N_5992);
xor U6151 (N_6151,N_5925,N_5863);
nand U6152 (N_6152,N_5912,N_5804);
nand U6153 (N_6153,N_5904,N_5987);
and U6154 (N_6154,N_5885,N_5836);
and U6155 (N_6155,N_5876,N_5835);
and U6156 (N_6156,N_5999,N_5932);
and U6157 (N_6157,N_5914,N_5831);
or U6158 (N_6158,N_5979,N_5982);
nor U6159 (N_6159,N_5869,N_5817);
xor U6160 (N_6160,N_5917,N_5876);
or U6161 (N_6161,N_5902,N_5909);
or U6162 (N_6162,N_5873,N_5981);
or U6163 (N_6163,N_5876,N_5863);
nand U6164 (N_6164,N_5896,N_5994);
and U6165 (N_6165,N_5825,N_5946);
and U6166 (N_6166,N_5881,N_5826);
nand U6167 (N_6167,N_5903,N_5810);
and U6168 (N_6168,N_5849,N_5826);
nand U6169 (N_6169,N_5836,N_5997);
or U6170 (N_6170,N_5910,N_5897);
xnor U6171 (N_6171,N_5834,N_5918);
xor U6172 (N_6172,N_5892,N_5897);
nand U6173 (N_6173,N_5987,N_5927);
nand U6174 (N_6174,N_5891,N_5969);
or U6175 (N_6175,N_5929,N_5848);
or U6176 (N_6176,N_5866,N_5995);
or U6177 (N_6177,N_5858,N_5915);
nor U6178 (N_6178,N_5991,N_5851);
nand U6179 (N_6179,N_5941,N_5844);
nand U6180 (N_6180,N_5922,N_5814);
nand U6181 (N_6181,N_5899,N_5877);
xor U6182 (N_6182,N_5906,N_5811);
nand U6183 (N_6183,N_5939,N_5978);
or U6184 (N_6184,N_5814,N_5909);
and U6185 (N_6185,N_5807,N_5818);
and U6186 (N_6186,N_5927,N_5936);
and U6187 (N_6187,N_5834,N_5800);
nor U6188 (N_6188,N_5835,N_5966);
or U6189 (N_6189,N_5848,N_5892);
and U6190 (N_6190,N_5907,N_5947);
nand U6191 (N_6191,N_5883,N_5935);
xor U6192 (N_6192,N_5923,N_5994);
or U6193 (N_6193,N_5884,N_5878);
xor U6194 (N_6194,N_5800,N_5912);
nor U6195 (N_6195,N_5887,N_5987);
and U6196 (N_6196,N_5928,N_5919);
nor U6197 (N_6197,N_5975,N_5834);
xnor U6198 (N_6198,N_5917,N_5820);
and U6199 (N_6199,N_5989,N_5970);
and U6200 (N_6200,N_6085,N_6193);
nor U6201 (N_6201,N_6063,N_6092);
nor U6202 (N_6202,N_6024,N_6005);
and U6203 (N_6203,N_6181,N_6052);
nand U6204 (N_6204,N_6144,N_6164);
nand U6205 (N_6205,N_6019,N_6114);
or U6206 (N_6206,N_6040,N_6195);
nand U6207 (N_6207,N_6097,N_6069);
nand U6208 (N_6208,N_6119,N_6037);
and U6209 (N_6209,N_6031,N_6056);
nand U6210 (N_6210,N_6038,N_6065);
nor U6211 (N_6211,N_6192,N_6194);
or U6212 (N_6212,N_6143,N_6004);
xor U6213 (N_6213,N_6151,N_6084);
nor U6214 (N_6214,N_6032,N_6190);
xnor U6215 (N_6215,N_6107,N_6178);
nand U6216 (N_6216,N_6000,N_6157);
and U6217 (N_6217,N_6015,N_6007);
nand U6218 (N_6218,N_6075,N_6156);
nand U6219 (N_6219,N_6172,N_6011);
nor U6220 (N_6220,N_6021,N_6048);
nor U6221 (N_6221,N_6134,N_6154);
xor U6222 (N_6222,N_6146,N_6179);
xnor U6223 (N_6223,N_6016,N_6116);
or U6224 (N_6224,N_6028,N_6029);
nand U6225 (N_6225,N_6125,N_6036);
and U6226 (N_6226,N_6171,N_6077);
and U6227 (N_6227,N_6080,N_6177);
nand U6228 (N_6228,N_6051,N_6082);
xnor U6229 (N_6229,N_6197,N_6142);
nand U6230 (N_6230,N_6073,N_6128);
or U6231 (N_6231,N_6130,N_6072);
and U6232 (N_6232,N_6101,N_6033);
nand U6233 (N_6233,N_6137,N_6027);
or U6234 (N_6234,N_6138,N_6147);
and U6235 (N_6235,N_6159,N_6083);
nand U6236 (N_6236,N_6124,N_6168);
or U6237 (N_6237,N_6166,N_6078);
nand U6238 (N_6238,N_6175,N_6127);
xnor U6239 (N_6239,N_6022,N_6086);
xor U6240 (N_6240,N_6186,N_6041);
or U6241 (N_6241,N_6030,N_6003);
and U6242 (N_6242,N_6060,N_6012);
or U6243 (N_6243,N_6108,N_6162);
and U6244 (N_6244,N_6176,N_6161);
nor U6245 (N_6245,N_6199,N_6053);
xor U6246 (N_6246,N_6044,N_6126);
and U6247 (N_6247,N_6133,N_6009);
xor U6248 (N_6248,N_6183,N_6165);
and U6249 (N_6249,N_6020,N_6163);
or U6250 (N_6250,N_6095,N_6196);
and U6251 (N_6251,N_6185,N_6132);
xor U6252 (N_6252,N_6034,N_6198);
nor U6253 (N_6253,N_6170,N_6136);
and U6254 (N_6254,N_6099,N_6158);
xnor U6255 (N_6255,N_6062,N_6008);
nand U6256 (N_6256,N_6081,N_6071);
or U6257 (N_6257,N_6122,N_6123);
nor U6258 (N_6258,N_6068,N_6167);
nor U6259 (N_6259,N_6118,N_6064);
and U6260 (N_6260,N_6070,N_6105);
nor U6261 (N_6261,N_6025,N_6090);
nor U6262 (N_6262,N_6067,N_6045);
xor U6263 (N_6263,N_6010,N_6093);
and U6264 (N_6264,N_6102,N_6113);
xnor U6265 (N_6265,N_6191,N_6087);
nor U6266 (N_6266,N_6046,N_6121);
nor U6267 (N_6267,N_6035,N_6079);
nand U6268 (N_6268,N_6160,N_6094);
and U6269 (N_6269,N_6039,N_6141);
nor U6270 (N_6270,N_6111,N_6155);
nor U6271 (N_6271,N_6135,N_6100);
nand U6272 (N_6272,N_6184,N_6189);
and U6273 (N_6273,N_6149,N_6049);
nor U6274 (N_6274,N_6061,N_6109);
or U6275 (N_6275,N_6091,N_6188);
and U6276 (N_6276,N_6014,N_6187);
xor U6277 (N_6277,N_6006,N_6140);
xor U6278 (N_6278,N_6103,N_6018);
and U6279 (N_6279,N_6153,N_6088);
nand U6280 (N_6280,N_6120,N_6131);
nand U6281 (N_6281,N_6112,N_6174);
and U6282 (N_6282,N_6050,N_6047);
xnor U6283 (N_6283,N_6023,N_6173);
nand U6284 (N_6284,N_6058,N_6059);
xnor U6285 (N_6285,N_6002,N_6145);
or U6286 (N_6286,N_6013,N_6054);
nand U6287 (N_6287,N_6089,N_6055);
and U6288 (N_6288,N_6098,N_6150);
xnor U6289 (N_6289,N_6152,N_6057);
or U6290 (N_6290,N_6182,N_6042);
xnor U6291 (N_6291,N_6148,N_6169);
xnor U6292 (N_6292,N_6074,N_6139);
and U6293 (N_6293,N_6115,N_6066);
xor U6294 (N_6294,N_6017,N_6117);
xor U6295 (N_6295,N_6106,N_6026);
nor U6296 (N_6296,N_6043,N_6129);
nand U6297 (N_6297,N_6001,N_6076);
and U6298 (N_6298,N_6104,N_6180);
xor U6299 (N_6299,N_6096,N_6110);
or U6300 (N_6300,N_6020,N_6085);
xor U6301 (N_6301,N_6113,N_6173);
nor U6302 (N_6302,N_6093,N_6176);
and U6303 (N_6303,N_6081,N_6150);
xnor U6304 (N_6304,N_6038,N_6177);
or U6305 (N_6305,N_6008,N_6184);
nor U6306 (N_6306,N_6124,N_6183);
and U6307 (N_6307,N_6141,N_6190);
xor U6308 (N_6308,N_6051,N_6011);
nor U6309 (N_6309,N_6050,N_6029);
and U6310 (N_6310,N_6005,N_6009);
nand U6311 (N_6311,N_6027,N_6117);
xnor U6312 (N_6312,N_6187,N_6070);
nor U6313 (N_6313,N_6138,N_6199);
or U6314 (N_6314,N_6072,N_6122);
xnor U6315 (N_6315,N_6165,N_6124);
nor U6316 (N_6316,N_6080,N_6191);
or U6317 (N_6317,N_6134,N_6144);
and U6318 (N_6318,N_6018,N_6078);
nand U6319 (N_6319,N_6050,N_6165);
or U6320 (N_6320,N_6089,N_6155);
xnor U6321 (N_6321,N_6085,N_6162);
nand U6322 (N_6322,N_6164,N_6187);
or U6323 (N_6323,N_6044,N_6138);
nand U6324 (N_6324,N_6156,N_6178);
and U6325 (N_6325,N_6129,N_6061);
nand U6326 (N_6326,N_6143,N_6048);
nand U6327 (N_6327,N_6091,N_6185);
xor U6328 (N_6328,N_6055,N_6173);
and U6329 (N_6329,N_6131,N_6038);
nand U6330 (N_6330,N_6122,N_6073);
and U6331 (N_6331,N_6073,N_6070);
nand U6332 (N_6332,N_6177,N_6076);
xor U6333 (N_6333,N_6008,N_6148);
or U6334 (N_6334,N_6072,N_6159);
xor U6335 (N_6335,N_6175,N_6147);
nor U6336 (N_6336,N_6043,N_6095);
xor U6337 (N_6337,N_6075,N_6143);
or U6338 (N_6338,N_6032,N_6177);
nor U6339 (N_6339,N_6083,N_6157);
or U6340 (N_6340,N_6047,N_6133);
or U6341 (N_6341,N_6048,N_6102);
nand U6342 (N_6342,N_6186,N_6137);
and U6343 (N_6343,N_6068,N_6104);
and U6344 (N_6344,N_6076,N_6046);
or U6345 (N_6345,N_6173,N_6146);
xor U6346 (N_6346,N_6164,N_6028);
nand U6347 (N_6347,N_6121,N_6017);
and U6348 (N_6348,N_6041,N_6000);
nor U6349 (N_6349,N_6062,N_6012);
nand U6350 (N_6350,N_6139,N_6123);
xnor U6351 (N_6351,N_6004,N_6087);
nor U6352 (N_6352,N_6178,N_6167);
or U6353 (N_6353,N_6037,N_6117);
or U6354 (N_6354,N_6096,N_6007);
and U6355 (N_6355,N_6061,N_6106);
or U6356 (N_6356,N_6192,N_6024);
xor U6357 (N_6357,N_6176,N_6062);
or U6358 (N_6358,N_6038,N_6048);
or U6359 (N_6359,N_6070,N_6035);
nor U6360 (N_6360,N_6021,N_6148);
or U6361 (N_6361,N_6130,N_6057);
nor U6362 (N_6362,N_6076,N_6123);
nor U6363 (N_6363,N_6142,N_6198);
xor U6364 (N_6364,N_6146,N_6061);
and U6365 (N_6365,N_6151,N_6082);
nor U6366 (N_6366,N_6080,N_6086);
or U6367 (N_6367,N_6198,N_6134);
or U6368 (N_6368,N_6057,N_6006);
xor U6369 (N_6369,N_6056,N_6187);
nor U6370 (N_6370,N_6150,N_6067);
and U6371 (N_6371,N_6166,N_6051);
nand U6372 (N_6372,N_6128,N_6169);
or U6373 (N_6373,N_6180,N_6023);
nand U6374 (N_6374,N_6025,N_6099);
or U6375 (N_6375,N_6178,N_6051);
nor U6376 (N_6376,N_6105,N_6047);
or U6377 (N_6377,N_6169,N_6040);
nor U6378 (N_6378,N_6069,N_6065);
nor U6379 (N_6379,N_6075,N_6042);
or U6380 (N_6380,N_6097,N_6023);
nand U6381 (N_6381,N_6093,N_6129);
or U6382 (N_6382,N_6086,N_6100);
and U6383 (N_6383,N_6090,N_6190);
nand U6384 (N_6384,N_6000,N_6091);
nor U6385 (N_6385,N_6188,N_6183);
nor U6386 (N_6386,N_6183,N_6039);
xor U6387 (N_6387,N_6153,N_6196);
and U6388 (N_6388,N_6133,N_6054);
or U6389 (N_6389,N_6170,N_6065);
nor U6390 (N_6390,N_6160,N_6164);
or U6391 (N_6391,N_6169,N_6129);
nor U6392 (N_6392,N_6164,N_6031);
nor U6393 (N_6393,N_6104,N_6193);
xnor U6394 (N_6394,N_6081,N_6059);
or U6395 (N_6395,N_6030,N_6113);
nor U6396 (N_6396,N_6092,N_6109);
nor U6397 (N_6397,N_6057,N_6148);
nand U6398 (N_6398,N_6099,N_6118);
nor U6399 (N_6399,N_6000,N_6084);
xnor U6400 (N_6400,N_6352,N_6395);
and U6401 (N_6401,N_6323,N_6219);
and U6402 (N_6402,N_6391,N_6260);
and U6403 (N_6403,N_6293,N_6264);
nor U6404 (N_6404,N_6338,N_6257);
or U6405 (N_6405,N_6220,N_6292);
and U6406 (N_6406,N_6243,N_6289);
xnor U6407 (N_6407,N_6203,N_6349);
nand U6408 (N_6408,N_6319,N_6222);
or U6409 (N_6409,N_6344,N_6394);
or U6410 (N_6410,N_6230,N_6308);
or U6411 (N_6411,N_6254,N_6299);
nor U6412 (N_6412,N_6273,N_6302);
nor U6413 (N_6413,N_6268,N_6231);
nand U6414 (N_6414,N_6387,N_6378);
or U6415 (N_6415,N_6337,N_6350);
and U6416 (N_6416,N_6356,N_6331);
nand U6417 (N_6417,N_6225,N_6362);
xnor U6418 (N_6418,N_6345,N_6275);
xnor U6419 (N_6419,N_6246,N_6250);
or U6420 (N_6420,N_6259,N_6200);
nor U6421 (N_6421,N_6363,N_6272);
nand U6422 (N_6422,N_6239,N_6364);
nand U6423 (N_6423,N_6318,N_6388);
nor U6424 (N_6424,N_6255,N_6375);
xnor U6425 (N_6425,N_6303,N_6202);
nor U6426 (N_6426,N_6283,N_6351);
and U6427 (N_6427,N_6228,N_6277);
nand U6428 (N_6428,N_6321,N_6296);
nand U6429 (N_6429,N_6297,N_6227);
or U6430 (N_6430,N_6361,N_6305);
nand U6431 (N_6431,N_6282,N_6376);
xor U6432 (N_6432,N_6201,N_6269);
nor U6433 (N_6433,N_6348,N_6379);
or U6434 (N_6434,N_6358,N_6393);
or U6435 (N_6435,N_6256,N_6317);
nor U6436 (N_6436,N_6233,N_6382);
and U6437 (N_6437,N_6209,N_6380);
nor U6438 (N_6438,N_6327,N_6244);
nand U6439 (N_6439,N_6206,N_6329);
xnor U6440 (N_6440,N_6347,N_6328);
nor U6441 (N_6441,N_6399,N_6270);
nor U6442 (N_6442,N_6389,N_6336);
nor U6443 (N_6443,N_6267,N_6396);
or U6444 (N_6444,N_6218,N_6371);
and U6445 (N_6445,N_6367,N_6281);
nor U6446 (N_6446,N_6340,N_6377);
nor U6447 (N_6447,N_6221,N_6290);
xor U6448 (N_6448,N_6360,N_6313);
or U6449 (N_6449,N_6383,N_6291);
xnor U6450 (N_6450,N_6211,N_6324);
nand U6451 (N_6451,N_6251,N_6310);
nand U6452 (N_6452,N_6370,N_6284);
xor U6453 (N_6453,N_6335,N_6217);
nor U6454 (N_6454,N_6315,N_6253);
nor U6455 (N_6455,N_6384,N_6248);
or U6456 (N_6456,N_6369,N_6210);
xnor U6457 (N_6457,N_6359,N_6258);
and U6458 (N_6458,N_6374,N_6261);
nand U6459 (N_6459,N_6214,N_6286);
nand U6460 (N_6460,N_6245,N_6204);
and U6461 (N_6461,N_6354,N_6208);
xor U6462 (N_6462,N_6307,N_6224);
xnor U6463 (N_6463,N_6366,N_6242);
xnor U6464 (N_6464,N_6288,N_6332);
and U6465 (N_6465,N_6316,N_6368);
nand U6466 (N_6466,N_6397,N_6262);
and U6467 (N_6467,N_6341,N_6346);
and U6468 (N_6468,N_6274,N_6322);
or U6469 (N_6469,N_6365,N_6241);
or U6470 (N_6470,N_6386,N_6287);
xor U6471 (N_6471,N_6314,N_6249);
nor U6472 (N_6472,N_6325,N_6278);
nand U6473 (N_6473,N_6266,N_6326);
nand U6474 (N_6474,N_6353,N_6390);
xnor U6475 (N_6475,N_6392,N_6312);
and U6476 (N_6476,N_6263,N_6213);
or U6477 (N_6477,N_6311,N_6301);
nor U6478 (N_6478,N_6235,N_6223);
and U6479 (N_6479,N_6309,N_6306);
and U6480 (N_6480,N_6343,N_6398);
nor U6481 (N_6481,N_6238,N_6304);
or U6482 (N_6482,N_6205,N_6237);
xnor U6483 (N_6483,N_6279,N_6372);
xnor U6484 (N_6484,N_6320,N_6247);
and U6485 (N_6485,N_6236,N_6381);
and U6486 (N_6486,N_6234,N_6357);
xor U6487 (N_6487,N_6240,N_6226);
or U6488 (N_6488,N_6339,N_6252);
or U6489 (N_6489,N_6276,N_6334);
nor U6490 (N_6490,N_6330,N_6271);
xnor U6491 (N_6491,N_6333,N_6385);
nor U6492 (N_6492,N_6207,N_6355);
xor U6493 (N_6493,N_6298,N_6232);
or U6494 (N_6494,N_6373,N_6212);
and U6495 (N_6495,N_6294,N_6229);
xnor U6496 (N_6496,N_6265,N_6300);
and U6497 (N_6497,N_6342,N_6295);
xnor U6498 (N_6498,N_6216,N_6215);
xor U6499 (N_6499,N_6280,N_6285);
or U6500 (N_6500,N_6200,N_6232);
xnor U6501 (N_6501,N_6218,N_6215);
and U6502 (N_6502,N_6324,N_6372);
or U6503 (N_6503,N_6331,N_6344);
nand U6504 (N_6504,N_6263,N_6352);
and U6505 (N_6505,N_6297,N_6330);
nand U6506 (N_6506,N_6225,N_6354);
xnor U6507 (N_6507,N_6331,N_6322);
or U6508 (N_6508,N_6334,N_6389);
nand U6509 (N_6509,N_6361,N_6387);
nor U6510 (N_6510,N_6201,N_6262);
xor U6511 (N_6511,N_6288,N_6230);
and U6512 (N_6512,N_6322,N_6391);
and U6513 (N_6513,N_6252,N_6347);
and U6514 (N_6514,N_6252,N_6397);
xnor U6515 (N_6515,N_6258,N_6261);
xor U6516 (N_6516,N_6388,N_6219);
nand U6517 (N_6517,N_6385,N_6398);
nand U6518 (N_6518,N_6303,N_6271);
and U6519 (N_6519,N_6217,N_6395);
or U6520 (N_6520,N_6359,N_6283);
xor U6521 (N_6521,N_6352,N_6258);
nand U6522 (N_6522,N_6286,N_6315);
or U6523 (N_6523,N_6336,N_6342);
and U6524 (N_6524,N_6341,N_6354);
or U6525 (N_6525,N_6221,N_6303);
xnor U6526 (N_6526,N_6366,N_6257);
xor U6527 (N_6527,N_6273,N_6318);
xor U6528 (N_6528,N_6351,N_6339);
or U6529 (N_6529,N_6348,N_6233);
nor U6530 (N_6530,N_6384,N_6207);
nand U6531 (N_6531,N_6267,N_6390);
and U6532 (N_6532,N_6325,N_6217);
xor U6533 (N_6533,N_6268,N_6327);
nand U6534 (N_6534,N_6391,N_6314);
xor U6535 (N_6535,N_6288,N_6391);
xor U6536 (N_6536,N_6284,N_6209);
nand U6537 (N_6537,N_6234,N_6393);
nand U6538 (N_6538,N_6397,N_6218);
and U6539 (N_6539,N_6317,N_6311);
xor U6540 (N_6540,N_6272,N_6375);
and U6541 (N_6541,N_6298,N_6240);
nor U6542 (N_6542,N_6255,N_6345);
xor U6543 (N_6543,N_6399,N_6213);
nor U6544 (N_6544,N_6339,N_6300);
xor U6545 (N_6545,N_6260,N_6375);
or U6546 (N_6546,N_6243,N_6207);
and U6547 (N_6547,N_6379,N_6285);
nor U6548 (N_6548,N_6364,N_6234);
or U6549 (N_6549,N_6216,N_6238);
nor U6550 (N_6550,N_6283,N_6244);
nor U6551 (N_6551,N_6309,N_6204);
nand U6552 (N_6552,N_6329,N_6346);
xor U6553 (N_6553,N_6391,N_6285);
nand U6554 (N_6554,N_6376,N_6211);
xor U6555 (N_6555,N_6258,N_6319);
or U6556 (N_6556,N_6397,N_6316);
xnor U6557 (N_6557,N_6319,N_6396);
nand U6558 (N_6558,N_6317,N_6248);
nand U6559 (N_6559,N_6297,N_6245);
nand U6560 (N_6560,N_6370,N_6297);
xor U6561 (N_6561,N_6376,N_6384);
and U6562 (N_6562,N_6339,N_6364);
nor U6563 (N_6563,N_6354,N_6218);
and U6564 (N_6564,N_6227,N_6298);
and U6565 (N_6565,N_6306,N_6372);
and U6566 (N_6566,N_6390,N_6389);
nor U6567 (N_6567,N_6317,N_6378);
nand U6568 (N_6568,N_6203,N_6233);
nor U6569 (N_6569,N_6312,N_6323);
nand U6570 (N_6570,N_6217,N_6270);
nor U6571 (N_6571,N_6333,N_6238);
or U6572 (N_6572,N_6382,N_6323);
nor U6573 (N_6573,N_6200,N_6320);
nor U6574 (N_6574,N_6251,N_6373);
nor U6575 (N_6575,N_6382,N_6338);
and U6576 (N_6576,N_6334,N_6305);
nand U6577 (N_6577,N_6342,N_6270);
nand U6578 (N_6578,N_6337,N_6383);
xor U6579 (N_6579,N_6249,N_6214);
or U6580 (N_6580,N_6207,N_6302);
or U6581 (N_6581,N_6288,N_6261);
or U6582 (N_6582,N_6272,N_6378);
nand U6583 (N_6583,N_6225,N_6392);
and U6584 (N_6584,N_6209,N_6212);
and U6585 (N_6585,N_6220,N_6238);
xnor U6586 (N_6586,N_6238,N_6240);
nand U6587 (N_6587,N_6309,N_6232);
xor U6588 (N_6588,N_6342,N_6247);
xnor U6589 (N_6589,N_6384,N_6203);
nand U6590 (N_6590,N_6378,N_6348);
nor U6591 (N_6591,N_6332,N_6371);
xor U6592 (N_6592,N_6206,N_6397);
nand U6593 (N_6593,N_6239,N_6347);
or U6594 (N_6594,N_6303,N_6287);
nor U6595 (N_6595,N_6200,N_6344);
nor U6596 (N_6596,N_6367,N_6317);
and U6597 (N_6597,N_6372,N_6252);
nor U6598 (N_6598,N_6334,N_6300);
xor U6599 (N_6599,N_6288,N_6325);
nand U6600 (N_6600,N_6471,N_6589);
nor U6601 (N_6601,N_6561,N_6448);
and U6602 (N_6602,N_6553,N_6419);
nor U6603 (N_6603,N_6430,N_6400);
xor U6604 (N_6604,N_6435,N_6531);
or U6605 (N_6605,N_6425,N_6483);
or U6606 (N_6606,N_6597,N_6560);
nor U6607 (N_6607,N_6529,N_6422);
nor U6608 (N_6608,N_6403,N_6418);
nor U6609 (N_6609,N_6532,N_6514);
nand U6610 (N_6610,N_6451,N_6501);
nand U6611 (N_6611,N_6449,N_6512);
or U6612 (N_6612,N_6443,N_6562);
or U6613 (N_6613,N_6496,N_6506);
nor U6614 (N_6614,N_6580,N_6417);
or U6615 (N_6615,N_6568,N_6444);
nand U6616 (N_6616,N_6557,N_6416);
nor U6617 (N_6617,N_6564,N_6491);
xnor U6618 (N_6618,N_6478,N_6412);
nand U6619 (N_6619,N_6459,N_6549);
xor U6620 (N_6620,N_6413,N_6457);
nand U6621 (N_6621,N_6463,N_6526);
and U6622 (N_6622,N_6405,N_6467);
or U6623 (N_6623,N_6547,N_6466);
or U6624 (N_6624,N_6535,N_6598);
or U6625 (N_6625,N_6592,N_6528);
nand U6626 (N_6626,N_6508,N_6423);
or U6627 (N_6627,N_6479,N_6411);
nor U6628 (N_6628,N_6455,N_6517);
or U6629 (N_6629,N_6590,N_6576);
nor U6630 (N_6630,N_6585,N_6499);
xor U6631 (N_6631,N_6475,N_6461);
nor U6632 (N_6632,N_6476,N_6572);
nand U6633 (N_6633,N_6495,N_6550);
nand U6634 (N_6634,N_6481,N_6545);
nand U6635 (N_6635,N_6502,N_6484);
nor U6636 (N_6636,N_6498,N_6519);
nor U6637 (N_6637,N_6540,N_6410);
nor U6638 (N_6638,N_6599,N_6588);
xor U6639 (N_6639,N_6534,N_6437);
nor U6640 (N_6640,N_6445,N_6537);
nor U6641 (N_6641,N_6493,N_6402);
xnor U6642 (N_6642,N_6446,N_6460);
nand U6643 (N_6643,N_6421,N_6582);
nand U6644 (N_6644,N_6480,N_6439);
or U6645 (N_6645,N_6551,N_6504);
and U6646 (N_6646,N_6452,N_6567);
nand U6647 (N_6647,N_6472,N_6489);
or U6648 (N_6648,N_6447,N_6584);
or U6649 (N_6649,N_6456,N_6497);
nand U6650 (N_6650,N_6510,N_6541);
or U6651 (N_6651,N_6490,N_6486);
or U6652 (N_6652,N_6574,N_6468);
or U6653 (N_6653,N_6513,N_6442);
and U6654 (N_6654,N_6518,N_6465);
nand U6655 (N_6655,N_6453,N_6548);
and U6656 (N_6656,N_6533,N_6424);
and U6657 (N_6657,N_6523,N_6426);
nand U6658 (N_6658,N_6487,N_6524);
and U6659 (N_6659,N_6503,N_6593);
nand U6660 (N_6660,N_6462,N_6511);
and U6661 (N_6661,N_6409,N_6470);
nor U6662 (N_6662,N_6492,N_6522);
or U6663 (N_6663,N_6520,N_6500);
nand U6664 (N_6664,N_6433,N_6594);
xnor U6665 (N_6665,N_6414,N_6407);
and U6666 (N_6666,N_6515,N_6438);
and U6667 (N_6667,N_6440,N_6577);
and U6668 (N_6668,N_6555,N_6516);
and U6669 (N_6669,N_6596,N_6458);
xnor U6670 (N_6670,N_6527,N_6488);
or U6671 (N_6671,N_6595,N_6566);
nor U6672 (N_6672,N_6558,N_6554);
and U6673 (N_6673,N_6454,N_6473);
nor U6674 (N_6674,N_6581,N_6575);
or U6675 (N_6675,N_6404,N_6583);
nand U6676 (N_6676,N_6544,N_6570);
and U6677 (N_6677,N_6543,N_6573);
xor U6678 (N_6678,N_6530,N_6556);
or U6679 (N_6679,N_6521,N_6450);
and U6680 (N_6680,N_6427,N_6401);
and U6681 (N_6681,N_6579,N_6571);
nor U6682 (N_6682,N_6429,N_6507);
and U6683 (N_6683,N_6509,N_6477);
nand U6684 (N_6684,N_6464,N_6586);
or U6685 (N_6685,N_6408,N_6525);
or U6686 (N_6686,N_6565,N_6436);
nand U6687 (N_6687,N_6563,N_6420);
nor U6688 (N_6688,N_6559,N_6546);
and U6689 (N_6689,N_6552,N_6474);
nor U6690 (N_6690,N_6482,N_6441);
xnor U6691 (N_6691,N_6536,N_6578);
or U6692 (N_6692,N_6415,N_6428);
nor U6693 (N_6693,N_6431,N_6591);
nor U6694 (N_6694,N_6469,N_6434);
and U6695 (N_6695,N_6505,N_6587);
and U6696 (N_6696,N_6406,N_6542);
or U6697 (N_6697,N_6538,N_6569);
nor U6698 (N_6698,N_6539,N_6485);
nand U6699 (N_6699,N_6494,N_6432);
or U6700 (N_6700,N_6525,N_6573);
nand U6701 (N_6701,N_6511,N_6520);
or U6702 (N_6702,N_6443,N_6564);
or U6703 (N_6703,N_6587,N_6473);
nand U6704 (N_6704,N_6434,N_6534);
or U6705 (N_6705,N_6459,N_6565);
or U6706 (N_6706,N_6454,N_6578);
or U6707 (N_6707,N_6568,N_6573);
nand U6708 (N_6708,N_6472,N_6470);
nand U6709 (N_6709,N_6596,N_6498);
nor U6710 (N_6710,N_6591,N_6468);
nand U6711 (N_6711,N_6455,N_6555);
nand U6712 (N_6712,N_6407,N_6580);
nand U6713 (N_6713,N_6430,N_6515);
and U6714 (N_6714,N_6447,N_6535);
nor U6715 (N_6715,N_6516,N_6549);
or U6716 (N_6716,N_6466,N_6521);
or U6717 (N_6717,N_6502,N_6591);
xnor U6718 (N_6718,N_6413,N_6404);
nand U6719 (N_6719,N_6435,N_6429);
nor U6720 (N_6720,N_6543,N_6462);
xnor U6721 (N_6721,N_6531,N_6571);
nor U6722 (N_6722,N_6414,N_6453);
nand U6723 (N_6723,N_6568,N_6413);
nor U6724 (N_6724,N_6583,N_6452);
or U6725 (N_6725,N_6400,N_6507);
nand U6726 (N_6726,N_6499,N_6586);
or U6727 (N_6727,N_6507,N_6557);
and U6728 (N_6728,N_6522,N_6526);
xor U6729 (N_6729,N_6551,N_6506);
nor U6730 (N_6730,N_6522,N_6451);
nor U6731 (N_6731,N_6424,N_6579);
xnor U6732 (N_6732,N_6496,N_6547);
nand U6733 (N_6733,N_6552,N_6575);
nor U6734 (N_6734,N_6489,N_6547);
or U6735 (N_6735,N_6558,N_6490);
nor U6736 (N_6736,N_6535,N_6508);
xor U6737 (N_6737,N_6536,N_6491);
nand U6738 (N_6738,N_6410,N_6588);
nor U6739 (N_6739,N_6579,N_6594);
and U6740 (N_6740,N_6431,N_6409);
nand U6741 (N_6741,N_6447,N_6489);
nor U6742 (N_6742,N_6421,N_6563);
nand U6743 (N_6743,N_6470,N_6447);
and U6744 (N_6744,N_6449,N_6559);
and U6745 (N_6745,N_6497,N_6415);
and U6746 (N_6746,N_6466,N_6440);
or U6747 (N_6747,N_6512,N_6423);
nor U6748 (N_6748,N_6456,N_6501);
nand U6749 (N_6749,N_6556,N_6566);
xnor U6750 (N_6750,N_6516,N_6531);
and U6751 (N_6751,N_6446,N_6466);
or U6752 (N_6752,N_6436,N_6498);
nor U6753 (N_6753,N_6448,N_6530);
and U6754 (N_6754,N_6426,N_6464);
and U6755 (N_6755,N_6527,N_6561);
xor U6756 (N_6756,N_6414,N_6445);
nand U6757 (N_6757,N_6589,N_6417);
and U6758 (N_6758,N_6529,N_6414);
or U6759 (N_6759,N_6547,N_6415);
and U6760 (N_6760,N_6444,N_6458);
nor U6761 (N_6761,N_6512,N_6546);
xor U6762 (N_6762,N_6505,N_6456);
nand U6763 (N_6763,N_6455,N_6540);
nor U6764 (N_6764,N_6593,N_6411);
and U6765 (N_6765,N_6473,N_6430);
xnor U6766 (N_6766,N_6438,N_6401);
nor U6767 (N_6767,N_6486,N_6566);
nand U6768 (N_6768,N_6597,N_6423);
or U6769 (N_6769,N_6456,N_6495);
nor U6770 (N_6770,N_6445,N_6452);
nor U6771 (N_6771,N_6491,N_6534);
or U6772 (N_6772,N_6418,N_6599);
xor U6773 (N_6773,N_6448,N_6438);
and U6774 (N_6774,N_6541,N_6507);
or U6775 (N_6775,N_6537,N_6576);
xnor U6776 (N_6776,N_6519,N_6494);
or U6777 (N_6777,N_6559,N_6563);
nand U6778 (N_6778,N_6411,N_6477);
or U6779 (N_6779,N_6502,N_6458);
or U6780 (N_6780,N_6454,N_6492);
xnor U6781 (N_6781,N_6565,N_6541);
or U6782 (N_6782,N_6553,N_6547);
or U6783 (N_6783,N_6414,N_6589);
or U6784 (N_6784,N_6426,N_6432);
and U6785 (N_6785,N_6402,N_6421);
and U6786 (N_6786,N_6483,N_6509);
or U6787 (N_6787,N_6436,N_6578);
nor U6788 (N_6788,N_6580,N_6533);
or U6789 (N_6789,N_6440,N_6545);
nor U6790 (N_6790,N_6502,N_6559);
or U6791 (N_6791,N_6422,N_6575);
nor U6792 (N_6792,N_6452,N_6549);
xnor U6793 (N_6793,N_6545,N_6574);
nand U6794 (N_6794,N_6461,N_6480);
nor U6795 (N_6795,N_6528,N_6408);
nand U6796 (N_6796,N_6506,N_6499);
nand U6797 (N_6797,N_6523,N_6491);
xnor U6798 (N_6798,N_6444,N_6591);
or U6799 (N_6799,N_6400,N_6525);
and U6800 (N_6800,N_6769,N_6627);
or U6801 (N_6801,N_6709,N_6723);
and U6802 (N_6802,N_6736,N_6620);
nand U6803 (N_6803,N_6662,N_6694);
nor U6804 (N_6804,N_6677,N_6617);
nand U6805 (N_6805,N_6759,N_6765);
xnor U6806 (N_6806,N_6732,N_6643);
or U6807 (N_6807,N_6754,N_6685);
and U6808 (N_6808,N_6634,N_6738);
nand U6809 (N_6809,N_6644,N_6648);
and U6810 (N_6810,N_6719,N_6673);
xor U6811 (N_6811,N_6670,N_6761);
nand U6812 (N_6812,N_6680,N_6785);
nor U6813 (N_6813,N_6651,N_6602);
nor U6814 (N_6814,N_6607,N_6678);
nand U6815 (N_6815,N_6737,N_6797);
or U6816 (N_6816,N_6717,N_6609);
nor U6817 (N_6817,N_6778,N_6716);
or U6818 (N_6818,N_6749,N_6681);
xor U6819 (N_6819,N_6603,N_6640);
nand U6820 (N_6820,N_6652,N_6649);
or U6821 (N_6821,N_6713,N_6753);
or U6822 (N_6822,N_6608,N_6776);
and U6823 (N_6823,N_6714,N_6746);
xnor U6824 (N_6824,N_6625,N_6780);
nor U6825 (N_6825,N_6739,N_6725);
nor U6826 (N_6826,N_6614,N_6663);
nand U6827 (N_6827,N_6702,N_6711);
and U6828 (N_6828,N_6619,N_6696);
xnor U6829 (N_6829,N_6756,N_6744);
xor U6830 (N_6830,N_6600,N_6782);
or U6831 (N_6831,N_6612,N_6712);
or U6832 (N_6832,N_6624,N_6748);
and U6833 (N_6833,N_6667,N_6731);
nor U6834 (N_6834,N_6764,N_6691);
nor U6835 (N_6835,N_6653,N_6792);
xor U6836 (N_6836,N_6626,N_6770);
or U6837 (N_6837,N_6729,N_6639);
nand U6838 (N_6838,N_6798,N_6789);
nor U6839 (N_6839,N_6795,N_6724);
and U6840 (N_6840,N_6752,N_6772);
and U6841 (N_6841,N_6706,N_6760);
and U6842 (N_6842,N_6777,N_6766);
nor U6843 (N_6843,N_6774,N_6616);
or U6844 (N_6844,N_6692,N_6718);
and U6845 (N_6845,N_6687,N_6796);
nand U6846 (N_6846,N_6728,N_6699);
nand U6847 (N_6847,N_6745,N_6799);
and U6848 (N_6848,N_6638,N_6615);
nand U6849 (N_6849,N_6751,N_6669);
and U6850 (N_6850,N_6665,N_6735);
xor U6851 (N_6851,N_6734,N_6771);
xnor U6852 (N_6852,N_6695,N_6794);
or U6853 (N_6853,N_6645,N_6604);
nor U6854 (N_6854,N_6621,N_6690);
and U6855 (N_6855,N_6700,N_6647);
xnor U6856 (N_6856,N_6633,N_6661);
or U6857 (N_6857,N_6635,N_6697);
or U6858 (N_6858,N_6664,N_6701);
and U6859 (N_6859,N_6659,N_6679);
or U6860 (N_6860,N_6632,N_6742);
xnor U6861 (N_6861,N_6727,N_6743);
nor U6862 (N_6862,N_6707,N_6790);
nor U6863 (N_6863,N_6686,N_6767);
xnor U6864 (N_6864,N_6793,N_6668);
and U6865 (N_6865,N_6650,N_6675);
nor U6866 (N_6866,N_6755,N_6688);
xnor U6867 (N_6867,N_6660,N_6672);
and U6868 (N_6868,N_6611,N_6721);
nand U6869 (N_6869,N_6740,N_6641);
xnor U6870 (N_6870,N_6787,N_6762);
and U6871 (N_6871,N_6773,N_6658);
xnor U6872 (N_6872,N_6683,N_6610);
or U6873 (N_6873,N_6689,N_6730);
and U6874 (N_6874,N_6656,N_6784);
nand U6875 (N_6875,N_6684,N_6698);
nor U6876 (N_6876,N_6628,N_6654);
nand U6877 (N_6877,N_6779,N_6726);
and U6878 (N_6878,N_6682,N_6646);
or U6879 (N_6879,N_6750,N_6757);
and U6880 (N_6880,N_6636,N_6622);
xnor U6881 (N_6881,N_6676,N_6618);
nor U6882 (N_6882,N_6775,N_6788);
xor U6883 (N_6883,N_6722,N_6715);
xor U6884 (N_6884,N_6623,N_6758);
xnor U6885 (N_6885,N_6629,N_6631);
nor U6886 (N_6886,N_6763,N_6705);
nand U6887 (N_6887,N_6655,N_6637);
nand U6888 (N_6888,N_6601,N_6786);
and U6889 (N_6889,N_6666,N_6741);
nand U6890 (N_6890,N_6642,N_6708);
nor U6891 (N_6891,N_6613,N_6710);
nor U6892 (N_6892,N_6657,N_6704);
nand U6893 (N_6893,N_6674,N_6781);
nand U6894 (N_6894,N_6605,N_6703);
and U6895 (N_6895,N_6783,N_6630);
and U6896 (N_6896,N_6791,N_6693);
or U6897 (N_6897,N_6733,N_6768);
or U6898 (N_6898,N_6606,N_6747);
or U6899 (N_6899,N_6671,N_6720);
xor U6900 (N_6900,N_6666,N_6780);
or U6901 (N_6901,N_6700,N_6773);
nand U6902 (N_6902,N_6664,N_6725);
nor U6903 (N_6903,N_6662,N_6675);
nor U6904 (N_6904,N_6616,N_6629);
nor U6905 (N_6905,N_6792,N_6768);
or U6906 (N_6906,N_6617,N_6797);
nor U6907 (N_6907,N_6613,N_6615);
nor U6908 (N_6908,N_6732,N_6703);
nand U6909 (N_6909,N_6781,N_6702);
nor U6910 (N_6910,N_6657,N_6759);
nor U6911 (N_6911,N_6672,N_6621);
nand U6912 (N_6912,N_6645,N_6653);
or U6913 (N_6913,N_6795,N_6790);
and U6914 (N_6914,N_6704,N_6699);
or U6915 (N_6915,N_6627,N_6688);
xnor U6916 (N_6916,N_6623,N_6724);
nand U6917 (N_6917,N_6759,N_6720);
and U6918 (N_6918,N_6715,N_6655);
nand U6919 (N_6919,N_6655,N_6723);
nor U6920 (N_6920,N_6660,N_6624);
or U6921 (N_6921,N_6717,N_6733);
xor U6922 (N_6922,N_6692,N_6629);
and U6923 (N_6923,N_6764,N_6792);
xor U6924 (N_6924,N_6611,N_6709);
xor U6925 (N_6925,N_6748,N_6759);
or U6926 (N_6926,N_6706,N_6743);
or U6927 (N_6927,N_6706,N_6799);
xnor U6928 (N_6928,N_6753,N_6722);
nand U6929 (N_6929,N_6711,N_6642);
nor U6930 (N_6930,N_6639,N_6721);
nor U6931 (N_6931,N_6739,N_6680);
and U6932 (N_6932,N_6662,N_6699);
nand U6933 (N_6933,N_6722,N_6764);
and U6934 (N_6934,N_6734,N_6721);
or U6935 (N_6935,N_6695,N_6646);
xnor U6936 (N_6936,N_6655,N_6631);
or U6937 (N_6937,N_6648,N_6603);
xnor U6938 (N_6938,N_6694,N_6774);
xnor U6939 (N_6939,N_6715,N_6699);
nor U6940 (N_6940,N_6631,N_6644);
xor U6941 (N_6941,N_6712,N_6634);
xor U6942 (N_6942,N_6681,N_6797);
and U6943 (N_6943,N_6741,N_6639);
or U6944 (N_6944,N_6791,N_6604);
nand U6945 (N_6945,N_6649,N_6741);
xor U6946 (N_6946,N_6751,N_6673);
nand U6947 (N_6947,N_6746,N_6664);
xnor U6948 (N_6948,N_6606,N_6675);
nand U6949 (N_6949,N_6713,N_6608);
xnor U6950 (N_6950,N_6718,N_6678);
and U6951 (N_6951,N_6619,N_6669);
or U6952 (N_6952,N_6742,N_6654);
nand U6953 (N_6953,N_6727,N_6660);
or U6954 (N_6954,N_6630,N_6699);
nand U6955 (N_6955,N_6725,N_6618);
xnor U6956 (N_6956,N_6768,N_6693);
and U6957 (N_6957,N_6618,N_6748);
xnor U6958 (N_6958,N_6759,N_6732);
nor U6959 (N_6959,N_6797,N_6632);
nor U6960 (N_6960,N_6638,N_6742);
xor U6961 (N_6961,N_6740,N_6661);
nor U6962 (N_6962,N_6775,N_6604);
and U6963 (N_6963,N_6651,N_6606);
or U6964 (N_6964,N_6786,N_6724);
and U6965 (N_6965,N_6655,N_6741);
or U6966 (N_6966,N_6671,N_6783);
nand U6967 (N_6967,N_6645,N_6785);
nor U6968 (N_6968,N_6632,N_6668);
nand U6969 (N_6969,N_6609,N_6707);
or U6970 (N_6970,N_6659,N_6606);
and U6971 (N_6971,N_6719,N_6725);
and U6972 (N_6972,N_6638,N_6706);
nor U6973 (N_6973,N_6702,N_6670);
or U6974 (N_6974,N_6768,N_6694);
nand U6975 (N_6975,N_6701,N_6673);
nand U6976 (N_6976,N_6711,N_6737);
or U6977 (N_6977,N_6744,N_6743);
xor U6978 (N_6978,N_6627,N_6667);
or U6979 (N_6979,N_6603,N_6692);
xor U6980 (N_6980,N_6752,N_6623);
or U6981 (N_6981,N_6650,N_6703);
and U6982 (N_6982,N_6732,N_6742);
nand U6983 (N_6983,N_6688,N_6656);
nand U6984 (N_6984,N_6752,N_6698);
or U6985 (N_6985,N_6757,N_6690);
and U6986 (N_6986,N_6616,N_6766);
nor U6987 (N_6987,N_6793,N_6762);
or U6988 (N_6988,N_6756,N_6718);
xor U6989 (N_6989,N_6695,N_6661);
and U6990 (N_6990,N_6693,N_6633);
nand U6991 (N_6991,N_6717,N_6689);
nor U6992 (N_6992,N_6699,N_6650);
nand U6993 (N_6993,N_6776,N_6779);
nand U6994 (N_6994,N_6673,N_6715);
and U6995 (N_6995,N_6660,N_6734);
nor U6996 (N_6996,N_6791,N_6662);
xnor U6997 (N_6997,N_6775,N_6794);
and U6998 (N_6998,N_6667,N_6720);
nor U6999 (N_6999,N_6639,N_6769);
and U7000 (N_7000,N_6941,N_6851);
nor U7001 (N_7001,N_6965,N_6853);
xnor U7002 (N_7002,N_6881,N_6976);
or U7003 (N_7003,N_6835,N_6968);
nand U7004 (N_7004,N_6951,N_6989);
nand U7005 (N_7005,N_6843,N_6926);
nand U7006 (N_7006,N_6988,N_6950);
nand U7007 (N_7007,N_6856,N_6986);
and U7008 (N_7008,N_6854,N_6923);
nor U7009 (N_7009,N_6957,N_6810);
or U7010 (N_7010,N_6934,N_6836);
nor U7011 (N_7011,N_6820,N_6806);
or U7012 (N_7012,N_6939,N_6831);
nor U7013 (N_7013,N_6822,N_6917);
and U7014 (N_7014,N_6932,N_6911);
and U7015 (N_7015,N_6924,N_6945);
and U7016 (N_7016,N_6936,N_6828);
or U7017 (N_7017,N_6889,N_6969);
and U7018 (N_7018,N_6960,N_6859);
xnor U7019 (N_7019,N_6821,N_6931);
nand U7020 (N_7020,N_6882,N_6996);
or U7021 (N_7021,N_6997,N_6861);
xnor U7022 (N_7022,N_6877,N_6947);
and U7023 (N_7023,N_6834,N_6868);
xor U7024 (N_7024,N_6898,N_6993);
or U7025 (N_7025,N_6925,N_6985);
nand U7026 (N_7026,N_6816,N_6927);
xnor U7027 (N_7027,N_6921,N_6885);
xor U7028 (N_7028,N_6920,N_6837);
nand U7029 (N_7029,N_6844,N_6862);
or U7030 (N_7030,N_6866,N_6805);
nor U7031 (N_7031,N_6841,N_6894);
and U7032 (N_7032,N_6940,N_6839);
nor U7033 (N_7033,N_6896,N_6994);
nor U7034 (N_7034,N_6930,N_6987);
or U7035 (N_7035,N_6879,N_6948);
or U7036 (N_7036,N_6928,N_6966);
xnor U7037 (N_7037,N_6829,N_6801);
or U7038 (N_7038,N_6919,N_6890);
xnor U7039 (N_7039,N_6863,N_6933);
and U7040 (N_7040,N_6982,N_6971);
and U7041 (N_7041,N_6999,N_6852);
or U7042 (N_7042,N_6904,N_6963);
nand U7043 (N_7043,N_6812,N_6893);
nor U7044 (N_7044,N_6978,N_6808);
nor U7045 (N_7045,N_6880,N_6876);
or U7046 (N_7046,N_6915,N_6954);
nand U7047 (N_7047,N_6850,N_6800);
nor U7048 (N_7048,N_6938,N_6906);
nand U7049 (N_7049,N_6952,N_6891);
nand U7050 (N_7050,N_6865,N_6935);
or U7051 (N_7051,N_6897,N_6975);
xnor U7052 (N_7052,N_6870,N_6949);
nor U7053 (N_7053,N_6956,N_6809);
and U7054 (N_7054,N_6990,N_6922);
nand U7055 (N_7055,N_6973,N_6977);
or U7056 (N_7056,N_6872,N_6903);
nor U7057 (N_7057,N_6959,N_6912);
or U7058 (N_7058,N_6817,N_6895);
or U7059 (N_7059,N_6998,N_6814);
xor U7060 (N_7060,N_6842,N_6929);
or U7061 (N_7061,N_6819,N_6955);
nor U7062 (N_7062,N_6832,N_6857);
and U7063 (N_7063,N_6943,N_6979);
or U7064 (N_7064,N_6825,N_6860);
nor U7065 (N_7065,N_6937,N_6830);
nand U7066 (N_7066,N_6864,N_6995);
nor U7067 (N_7067,N_6907,N_6961);
and U7068 (N_7068,N_6807,N_6884);
nor U7069 (N_7069,N_6802,N_6840);
xor U7070 (N_7070,N_6962,N_6970);
xor U7071 (N_7071,N_6901,N_6826);
xnor U7072 (N_7072,N_6871,N_6855);
nand U7073 (N_7073,N_6823,N_6953);
or U7074 (N_7074,N_6983,N_6815);
nor U7075 (N_7075,N_6867,N_6914);
nand U7076 (N_7076,N_6883,N_6869);
xor U7077 (N_7077,N_6845,N_6902);
nand U7078 (N_7078,N_6913,N_6899);
nor U7079 (N_7079,N_6827,N_6944);
nand U7080 (N_7080,N_6813,N_6909);
xor U7081 (N_7081,N_6974,N_6803);
nand U7082 (N_7082,N_6958,N_6946);
and U7083 (N_7083,N_6804,N_6874);
or U7084 (N_7084,N_6838,N_6984);
xor U7085 (N_7085,N_6892,N_6873);
and U7086 (N_7086,N_6848,N_6886);
or U7087 (N_7087,N_6991,N_6833);
and U7088 (N_7088,N_6878,N_6964);
and U7089 (N_7089,N_6824,N_6888);
nor U7090 (N_7090,N_6910,N_6875);
or U7091 (N_7091,N_6858,N_6942);
and U7092 (N_7092,N_6981,N_6967);
nor U7093 (N_7093,N_6900,N_6905);
xor U7094 (N_7094,N_6972,N_6846);
or U7095 (N_7095,N_6918,N_6992);
or U7096 (N_7096,N_6908,N_6847);
or U7097 (N_7097,N_6849,N_6916);
nor U7098 (N_7098,N_6887,N_6811);
and U7099 (N_7099,N_6818,N_6980);
nor U7100 (N_7100,N_6893,N_6820);
or U7101 (N_7101,N_6892,N_6862);
and U7102 (N_7102,N_6903,N_6813);
nand U7103 (N_7103,N_6850,N_6924);
and U7104 (N_7104,N_6848,N_6868);
nand U7105 (N_7105,N_6811,N_6866);
xor U7106 (N_7106,N_6846,N_6952);
nor U7107 (N_7107,N_6988,N_6962);
nand U7108 (N_7108,N_6979,N_6998);
nand U7109 (N_7109,N_6957,N_6903);
nand U7110 (N_7110,N_6991,N_6905);
or U7111 (N_7111,N_6868,N_6807);
nand U7112 (N_7112,N_6925,N_6952);
xnor U7113 (N_7113,N_6834,N_6921);
or U7114 (N_7114,N_6869,N_6938);
nand U7115 (N_7115,N_6960,N_6974);
nand U7116 (N_7116,N_6818,N_6875);
nand U7117 (N_7117,N_6902,N_6978);
nor U7118 (N_7118,N_6954,N_6856);
nor U7119 (N_7119,N_6873,N_6869);
and U7120 (N_7120,N_6897,N_6881);
or U7121 (N_7121,N_6890,N_6983);
nand U7122 (N_7122,N_6922,N_6827);
nor U7123 (N_7123,N_6814,N_6833);
and U7124 (N_7124,N_6804,N_6950);
or U7125 (N_7125,N_6864,N_6913);
and U7126 (N_7126,N_6896,N_6917);
xor U7127 (N_7127,N_6801,N_6809);
nand U7128 (N_7128,N_6871,N_6908);
nor U7129 (N_7129,N_6968,N_6849);
or U7130 (N_7130,N_6947,N_6875);
xnor U7131 (N_7131,N_6930,N_6873);
nand U7132 (N_7132,N_6994,N_6842);
and U7133 (N_7133,N_6925,N_6854);
and U7134 (N_7134,N_6801,N_6905);
nor U7135 (N_7135,N_6988,N_6900);
and U7136 (N_7136,N_6853,N_6945);
nand U7137 (N_7137,N_6859,N_6835);
or U7138 (N_7138,N_6834,N_6999);
and U7139 (N_7139,N_6996,N_6991);
or U7140 (N_7140,N_6886,N_6936);
nor U7141 (N_7141,N_6967,N_6872);
and U7142 (N_7142,N_6975,N_6960);
xor U7143 (N_7143,N_6998,N_6904);
xnor U7144 (N_7144,N_6987,N_6960);
nand U7145 (N_7145,N_6945,N_6859);
or U7146 (N_7146,N_6983,N_6863);
and U7147 (N_7147,N_6999,N_6937);
xnor U7148 (N_7148,N_6999,N_6939);
xnor U7149 (N_7149,N_6828,N_6942);
and U7150 (N_7150,N_6873,N_6819);
and U7151 (N_7151,N_6830,N_6920);
nand U7152 (N_7152,N_6852,N_6874);
and U7153 (N_7153,N_6833,N_6924);
nor U7154 (N_7154,N_6907,N_6850);
or U7155 (N_7155,N_6852,N_6929);
xnor U7156 (N_7156,N_6814,N_6800);
nand U7157 (N_7157,N_6952,N_6986);
nor U7158 (N_7158,N_6856,N_6884);
or U7159 (N_7159,N_6914,N_6937);
xor U7160 (N_7160,N_6954,N_6858);
or U7161 (N_7161,N_6924,N_6820);
and U7162 (N_7162,N_6887,N_6826);
nor U7163 (N_7163,N_6934,N_6904);
nor U7164 (N_7164,N_6966,N_6956);
or U7165 (N_7165,N_6911,N_6845);
nor U7166 (N_7166,N_6837,N_6943);
nor U7167 (N_7167,N_6836,N_6857);
nand U7168 (N_7168,N_6986,N_6987);
or U7169 (N_7169,N_6932,N_6855);
and U7170 (N_7170,N_6945,N_6977);
or U7171 (N_7171,N_6988,N_6895);
or U7172 (N_7172,N_6910,N_6852);
or U7173 (N_7173,N_6809,N_6950);
nand U7174 (N_7174,N_6848,N_6909);
nand U7175 (N_7175,N_6904,N_6848);
or U7176 (N_7176,N_6999,N_6893);
nor U7177 (N_7177,N_6847,N_6832);
nand U7178 (N_7178,N_6971,N_6919);
or U7179 (N_7179,N_6967,N_6818);
xnor U7180 (N_7180,N_6857,N_6864);
or U7181 (N_7181,N_6804,N_6997);
or U7182 (N_7182,N_6947,N_6880);
nor U7183 (N_7183,N_6947,N_6823);
xnor U7184 (N_7184,N_6867,N_6812);
xnor U7185 (N_7185,N_6818,N_6968);
and U7186 (N_7186,N_6840,N_6919);
and U7187 (N_7187,N_6812,N_6965);
and U7188 (N_7188,N_6814,N_6846);
xor U7189 (N_7189,N_6858,N_6841);
xnor U7190 (N_7190,N_6937,N_6887);
nand U7191 (N_7191,N_6975,N_6943);
nor U7192 (N_7192,N_6899,N_6876);
nor U7193 (N_7193,N_6981,N_6871);
nand U7194 (N_7194,N_6872,N_6905);
xnor U7195 (N_7195,N_6873,N_6842);
or U7196 (N_7196,N_6993,N_6979);
or U7197 (N_7197,N_6905,N_6836);
nor U7198 (N_7198,N_6906,N_6842);
or U7199 (N_7199,N_6933,N_6916);
xor U7200 (N_7200,N_7193,N_7179);
or U7201 (N_7201,N_7109,N_7180);
and U7202 (N_7202,N_7049,N_7124);
nand U7203 (N_7203,N_7095,N_7198);
or U7204 (N_7204,N_7041,N_7037);
nand U7205 (N_7205,N_7188,N_7196);
and U7206 (N_7206,N_7184,N_7089);
nor U7207 (N_7207,N_7067,N_7192);
nor U7208 (N_7208,N_7068,N_7098);
or U7209 (N_7209,N_7127,N_7161);
nand U7210 (N_7210,N_7024,N_7014);
nor U7211 (N_7211,N_7149,N_7182);
nor U7212 (N_7212,N_7054,N_7141);
nor U7213 (N_7213,N_7045,N_7135);
or U7214 (N_7214,N_7131,N_7060);
xor U7215 (N_7215,N_7016,N_7186);
xnor U7216 (N_7216,N_7084,N_7197);
or U7217 (N_7217,N_7165,N_7033);
nor U7218 (N_7218,N_7071,N_7132);
nand U7219 (N_7219,N_7107,N_7072);
xnor U7220 (N_7220,N_7062,N_7001);
or U7221 (N_7221,N_7134,N_7122);
nor U7222 (N_7222,N_7085,N_7123);
and U7223 (N_7223,N_7082,N_7020);
nor U7224 (N_7224,N_7034,N_7030);
xnor U7225 (N_7225,N_7042,N_7148);
and U7226 (N_7226,N_7140,N_7046);
nor U7227 (N_7227,N_7077,N_7097);
nand U7228 (N_7228,N_7117,N_7094);
or U7229 (N_7229,N_7078,N_7119);
nor U7230 (N_7230,N_7090,N_7151);
nand U7231 (N_7231,N_7050,N_7061);
and U7232 (N_7232,N_7102,N_7137);
xnor U7233 (N_7233,N_7091,N_7063);
xnor U7234 (N_7234,N_7138,N_7006);
or U7235 (N_7235,N_7093,N_7010);
nand U7236 (N_7236,N_7076,N_7177);
nand U7237 (N_7237,N_7000,N_7155);
or U7238 (N_7238,N_7043,N_7163);
and U7239 (N_7239,N_7115,N_7057);
xor U7240 (N_7240,N_7023,N_7027);
and U7241 (N_7241,N_7136,N_7111);
or U7242 (N_7242,N_7053,N_7168);
and U7243 (N_7243,N_7189,N_7047);
or U7244 (N_7244,N_7178,N_7065);
xor U7245 (N_7245,N_7174,N_7066);
nor U7246 (N_7246,N_7081,N_7035);
nor U7247 (N_7247,N_7031,N_7160);
xnor U7248 (N_7248,N_7099,N_7157);
xor U7249 (N_7249,N_7129,N_7007);
nand U7250 (N_7250,N_7044,N_7059);
and U7251 (N_7251,N_7074,N_7086);
xor U7252 (N_7252,N_7166,N_7170);
nor U7253 (N_7253,N_7199,N_7159);
or U7254 (N_7254,N_7058,N_7012);
or U7255 (N_7255,N_7147,N_7164);
and U7256 (N_7256,N_7021,N_7187);
nand U7257 (N_7257,N_7103,N_7175);
xor U7258 (N_7258,N_7083,N_7073);
nor U7259 (N_7259,N_7185,N_7026);
and U7260 (N_7260,N_7013,N_7105);
or U7261 (N_7261,N_7079,N_7025);
nand U7262 (N_7262,N_7029,N_7088);
and U7263 (N_7263,N_7130,N_7145);
nand U7264 (N_7264,N_7018,N_7022);
nand U7265 (N_7265,N_7051,N_7154);
nor U7266 (N_7266,N_7005,N_7128);
nand U7267 (N_7267,N_7069,N_7183);
xor U7268 (N_7268,N_7101,N_7008);
nor U7269 (N_7269,N_7181,N_7144);
nor U7270 (N_7270,N_7019,N_7106);
or U7271 (N_7271,N_7104,N_7096);
nor U7272 (N_7272,N_7116,N_7191);
nand U7273 (N_7273,N_7092,N_7142);
or U7274 (N_7274,N_7120,N_7080);
nor U7275 (N_7275,N_7112,N_7133);
or U7276 (N_7276,N_7039,N_7011);
nor U7277 (N_7277,N_7056,N_7015);
nor U7278 (N_7278,N_7172,N_7004);
and U7279 (N_7279,N_7176,N_7110);
nand U7280 (N_7280,N_7195,N_7190);
xnor U7281 (N_7281,N_7113,N_7125);
nand U7282 (N_7282,N_7028,N_7064);
nand U7283 (N_7283,N_7002,N_7139);
and U7284 (N_7284,N_7153,N_7070);
and U7285 (N_7285,N_7162,N_7087);
nor U7286 (N_7286,N_7194,N_7108);
xnor U7287 (N_7287,N_7052,N_7118);
nand U7288 (N_7288,N_7167,N_7158);
xnor U7289 (N_7289,N_7150,N_7171);
and U7290 (N_7290,N_7143,N_7075);
nand U7291 (N_7291,N_7152,N_7114);
or U7292 (N_7292,N_7003,N_7169);
nand U7293 (N_7293,N_7126,N_7017);
nor U7294 (N_7294,N_7009,N_7100);
nand U7295 (N_7295,N_7032,N_7173);
xor U7296 (N_7296,N_7038,N_7040);
and U7297 (N_7297,N_7146,N_7156);
xor U7298 (N_7298,N_7121,N_7055);
nor U7299 (N_7299,N_7036,N_7048);
nor U7300 (N_7300,N_7196,N_7192);
and U7301 (N_7301,N_7117,N_7148);
xor U7302 (N_7302,N_7008,N_7083);
or U7303 (N_7303,N_7135,N_7140);
and U7304 (N_7304,N_7175,N_7162);
or U7305 (N_7305,N_7028,N_7150);
xnor U7306 (N_7306,N_7064,N_7194);
nor U7307 (N_7307,N_7176,N_7047);
or U7308 (N_7308,N_7033,N_7042);
or U7309 (N_7309,N_7149,N_7025);
or U7310 (N_7310,N_7013,N_7198);
nor U7311 (N_7311,N_7002,N_7026);
nor U7312 (N_7312,N_7132,N_7192);
nand U7313 (N_7313,N_7005,N_7159);
nor U7314 (N_7314,N_7088,N_7101);
xor U7315 (N_7315,N_7075,N_7113);
and U7316 (N_7316,N_7020,N_7036);
xor U7317 (N_7317,N_7075,N_7003);
xor U7318 (N_7318,N_7003,N_7032);
or U7319 (N_7319,N_7121,N_7149);
xnor U7320 (N_7320,N_7116,N_7076);
nor U7321 (N_7321,N_7068,N_7001);
xor U7322 (N_7322,N_7176,N_7000);
or U7323 (N_7323,N_7167,N_7046);
nor U7324 (N_7324,N_7019,N_7001);
or U7325 (N_7325,N_7017,N_7112);
xnor U7326 (N_7326,N_7160,N_7163);
nor U7327 (N_7327,N_7149,N_7177);
and U7328 (N_7328,N_7082,N_7137);
and U7329 (N_7329,N_7146,N_7071);
nand U7330 (N_7330,N_7082,N_7156);
and U7331 (N_7331,N_7015,N_7044);
and U7332 (N_7332,N_7078,N_7188);
or U7333 (N_7333,N_7147,N_7180);
and U7334 (N_7334,N_7025,N_7097);
nand U7335 (N_7335,N_7154,N_7006);
nor U7336 (N_7336,N_7057,N_7097);
nand U7337 (N_7337,N_7052,N_7079);
nand U7338 (N_7338,N_7056,N_7106);
nor U7339 (N_7339,N_7162,N_7068);
nand U7340 (N_7340,N_7056,N_7017);
or U7341 (N_7341,N_7035,N_7093);
nand U7342 (N_7342,N_7108,N_7154);
and U7343 (N_7343,N_7029,N_7180);
nor U7344 (N_7344,N_7061,N_7157);
nand U7345 (N_7345,N_7023,N_7015);
or U7346 (N_7346,N_7158,N_7138);
nand U7347 (N_7347,N_7103,N_7104);
nand U7348 (N_7348,N_7041,N_7078);
and U7349 (N_7349,N_7010,N_7059);
nand U7350 (N_7350,N_7005,N_7179);
xnor U7351 (N_7351,N_7013,N_7030);
and U7352 (N_7352,N_7182,N_7171);
or U7353 (N_7353,N_7134,N_7023);
nand U7354 (N_7354,N_7163,N_7026);
and U7355 (N_7355,N_7181,N_7115);
xnor U7356 (N_7356,N_7183,N_7148);
nor U7357 (N_7357,N_7133,N_7192);
and U7358 (N_7358,N_7069,N_7018);
nand U7359 (N_7359,N_7034,N_7019);
xnor U7360 (N_7360,N_7116,N_7133);
nor U7361 (N_7361,N_7094,N_7158);
nand U7362 (N_7362,N_7017,N_7022);
and U7363 (N_7363,N_7196,N_7071);
or U7364 (N_7364,N_7146,N_7105);
and U7365 (N_7365,N_7065,N_7086);
nand U7366 (N_7366,N_7097,N_7008);
xnor U7367 (N_7367,N_7130,N_7186);
nand U7368 (N_7368,N_7064,N_7075);
nand U7369 (N_7369,N_7175,N_7158);
nand U7370 (N_7370,N_7109,N_7112);
xor U7371 (N_7371,N_7153,N_7100);
xor U7372 (N_7372,N_7009,N_7024);
nand U7373 (N_7373,N_7096,N_7093);
xnor U7374 (N_7374,N_7110,N_7099);
or U7375 (N_7375,N_7087,N_7125);
nand U7376 (N_7376,N_7179,N_7153);
xnor U7377 (N_7377,N_7186,N_7161);
xnor U7378 (N_7378,N_7081,N_7168);
or U7379 (N_7379,N_7128,N_7133);
nand U7380 (N_7380,N_7113,N_7051);
xnor U7381 (N_7381,N_7154,N_7199);
and U7382 (N_7382,N_7015,N_7099);
nor U7383 (N_7383,N_7184,N_7033);
and U7384 (N_7384,N_7030,N_7065);
nand U7385 (N_7385,N_7097,N_7108);
and U7386 (N_7386,N_7015,N_7001);
or U7387 (N_7387,N_7011,N_7126);
nor U7388 (N_7388,N_7060,N_7129);
and U7389 (N_7389,N_7030,N_7168);
and U7390 (N_7390,N_7196,N_7077);
nor U7391 (N_7391,N_7088,N_7055);
xor U7392 (N_7392,N_7197,N_7133);
nand U7393 (N_7393,N_7142,N_7127);
or U7394 (N_7394,N_7018,N_7107);
or U7395 (N_7395,N_7172,N_7152);
and U7396 (N_7396,N_7144,N_7103);
nor U7397 (N_7397,N_7099,N_7194);
and U7398 (N_7398,N_7172,N_7023);
nand U7399 (N_7399,N_7134,N_7136);
nor U7400 (N_7400,N_7252,N_7295);
and U7401 (N_7401,N_7326,N_7369);
nand U7402 (N_7402,N_7328,N_7346);
xnor U7403 (N_7403,N_7329,N_7390);
nor U7404 (N_7404,N_7376,N_7293);
xnor U7405 (N_7405,N_7245,N_7388);
nand U7406 (N_7406,N_7363,N_7338);
or U7407 (N_7407,N_7279,N_7237);
xnor U7408 (N_7408,N_7244,N_7332);
nand U7409 (N_7409,N_7311,N_7362);
xnor U7410 (N_7410,N_7222,N_7254);
or U7411 (N_7411,N_7281,N_7273);
or U7412 (N_7412,N_7209,N_7353);
xor U7413 (N_7413,N_7305,N_7317);
or U7414 (N_7414,N_7228,N_7283);
and U7415 (N_7415,N_7345,N_7337);
nor U7416 (N_7416,N_7232,N_7284);
and U7417 (N_7417,N_7212,N_7241);
nand U7418 (N_7418,N_7218,N_7367);
and U7419 (N_7419,N_7313,N_7331);
or U7420 (N_7420,N_7334,N_7223);
xnor U7421 (N_7421,N_7253,N_7265);
xnor U7422 (N_7422,N_7202,N_7397);
nor U7423 (N_7423,N_7240,N_7392);
nand U7424 (N_7424,N_7382,N_7230);
nor U7425 (N_7425,N_7204,N_7303);
nor U7426 (N_7426,N_7231,N_7296);
xnor U7427 (N_7427,N_7300,N_7327);
nor U7428 (N_7428,N_7297,N_7221);
nand U7429 (N_7429,N_7394,N_7321);
and U7430 (N_7430,N_7272,N_7347);
xor U7431 (N_7431,N_7286,N_7319);
nor U7432 (N_7432,N_7301,N_7391);
xnor U7433 (N_7433,N_7375,N_7264);
nand U7434 (N_7434,N_7262,N_7356);
nor U7435 (N_7435,N_7280,N_7269);
xor U7436 (N_7436,N_7210,N_7277);
xor U7437 (N_7437,N_7387,N_7208);
xor U7438 (N_7438,N_7235,N_7278);
nand U7439 (N_7439,N_7217,N_7276);
xor U7440 (N_7440,N_7211,N_7372);
nor U7441 (N_7441,N_7261,N_7386);
xnor U7442 (N_7442,N_7361,N_7378);
and U7443 (N_7443,N_7294,N_7381);
nor U7444 (N_7444,N_7214,N_7370);
xnor U7445 (N_7445,N_7229,N_7312);
and U7446 (N_7446,N_7325,N_7288);
and U7447 (N_7447,N_7216,N_7355);
or U7448 (N_7448,N_7315,N_7396);
xnor U7449 (N_7449,N_7292,N_7318);
xnor U7450 (N_7450,N_7266,N_7340);
or U7451 (N_7451,N_7398,N_7291);
nor U7452 (N_7452,N_7360,N_7215);
nor U7453 (N_7453,N_7399,N_7380);
or U7454 (N_7454,N_7234,N_7383);
or U7455 (N_7455,N_7268,N_7227);
nor U7456 (N_7456,N_7351,N_7336);
or U7457 (N_7457,N_7207,N_7333);
nand U7458 (N_7458,N_7259,N_7242);
xnor U7459 (N_7459,N_7299,N_7330);
or U7460 (N_7460,N_7258,N_7274);
and U7461 (N_7461,N_7395,N_7371);
and U7462 (N_7462,N_7250,N_7343);
xnor U7463 (N_7463,N_7341,N_7309);
xnor U7464 (N_7464,N_7385,N_7200);
xor U7465 (N_7465,N_7206,N_7306);
or U7466 (N_7466,N_7335,N_7203);
nor U7467 (N_7467,N_7239,N_7352);
and U7468 (N_7468,N_7260,N_7307);
and U7469 (N_7469,N_7289,N_7320);
xor U7470 (N_7470,N_7225,N_7224);
and U7471 (N_7471,N_7287,N_7282);
nand U7472 (N_7472,N_7365,N_7249);
nor U7473 (N_7473,N_7246,N_7233);
nor U7474 (N_7474,N_7348,N_7322);
xnor U7475 (N_7475,N_7377,N_7389);
xnor U7476 (N_7476,N_7275,N_7359);
nand U7477 (N_7477,N_7310,N_7247);
or U7478 (N_7478,N_7213,N_7285);
xor U7479 (N_7479,N_7344,N_7373);
and U7480 (N_7480,N_7358,N_7350);
nor U7481 (N_7481,N_7256,N_7379);
or U7482 (N_7482,N_7238,N_7251);
and U7483 (N_7483,N_7270,N_7255);
xnor U7484 (N_7484,N_7271,N_7339);
nor U7485 (N_7485,N_7368,N_7304);
or U7486 (N_7486,N_7314,N_7384);
and U7487 (N_7487,N_7226,N_7248);
or U7488 (N_7488,N_7357,N_7267);
xor U7489 (N_7489,N_7316,N_7219);
or U7490 (N_7490,N_7298,N_7374);
xor U7491 (N_7491,N_7263,N_7201);
and U7492 (N_7492,N_7324,N_7354);
nand U7493 (N_7493,N_7323,N_7349);
xor U7494 (N_7494,N_7366,N_7302);
nand U7495 (N_7495,N_7220,N_7243);
or U7496 (N_7496,N_7257,N_7364);
and U7497 (N_7497,N_7290,N_7205);
nand U7498 (N_7498,N_7342,N_7308);
nand U7499 (N_7499,N_7393,N_7236);
and U7500 (N_7500,N_7241,N_7328);
and U7501 (N_7501,N_7240,N_7266);
nand U7502 (N_7502,N_7346,N_7266);
nor U7503 (N_7503,N_7366,N_7211);
and U7504 (N_7504,N_7310,N_7224);
nor U7505 (N_7505,N_7240,N_7309);
xnor U7506 (N_7506,N_7204,N_7247);
nand U7507 (N_7507,N_7344,N_7296);
xnor U7508 (N_7508,N_7249,N_7257);
xnor U7509 (N_7509,N_7223,N_7388);
and U7510 (N_7510,N_7260,N_7345);
nand U7511 (N_7511,N_7204,N_7219);
and U7512 (N_7512,N_7360,N_7397);
and U7513 (N_7513,N_7332,N_7273);
xor U7514 (N_7514,N_7309,N_7272);
and U7515 (N_7515,N_7255,N_7371);
xnor U7516 (N_7516,N_7312,N_7350);
or U7517 (N_7517,N_7373,N_7293);
nor U7518 (N_7518,N_7270,N_7352);
xnor U7519 (N_7519,N_7249,N_7393);
xnor U7520 (N_7520,N_7316,N_7311);
and U7521 (N_7521,N_7306,N_7376);
or U7522 (N_7522,N_7249,N_7253);
or U7523 (N_7523,N_7339,N_7290);
and U7524 (N_7524,N_7250,N_7388);
nor U7525 (N_7525,N_7389,N_7288);
or U7526 (N_7526,N_7285,N_7342);
nand U7527 (N_7527,N_7323,N_7379);
nor U7528 (N_7528,N_7281,N_7272);
xnor U7529 (N_7529,N_7386,N_7223);
or U7530 (N_7530,N_7258,N_7232);
or U7531 (N_7531,N_7372,N_7395);
or U7532 (N_7532,N_7238,N_7216);
or U7533 (N_7533,N_7224,N_7334);
nor U7534 (N_7534,N_7237,N_7206);
and U7535 (N_7535,N_7230,N_7353);
or U7536 (N_7536,N_7340,N_7315);
or U7537 (N_7537,N_7264,N_7346);
or U7538 (N_7538,N_7211,N_7391);
or U7539 (N_7539,N_7227,N_7358);
or U7540 (N_7540,N_7275,N_7396);
and U7541 (N_7541,N_7272,N_7233);
nor U7542 (N_7542,N_7353,N_7361);
nand U7543 (N_7543,N_7236,N_7251);
nor U7544 (N_7544,N_7243,N_7317);
and U7545 (N_7545,N_7364,N_7358);
and U7546 (N_7546,N_7281,N_7242);
or U7547 (N_7547,N_7287,N_7211);
xnor U7548 (N_7548,N_7314,N_7219);
nand U7549 (N_7549,N_7217,N_7393);
or U7550 (N_7550,N_7282,N_7263);
nand U7551 (N_7551,N_7240,N_7367);
xnor U7552 (N_7552,N_7264,N_7374);
xnor U7553 (N_7553,N_7282,N_7268);
xor U7554 (N_7554,N_7204,N_7353);
xor U7555 (N_7555,N_7237,N_7223);
nor U7556 (N_7556,N_7366,N_7270);
and U7557 (N_7557,N_7246,N_7358);
nor U7558 (N_7558,N_7390,N_7221);
xnor U7559 (N_7559,N_7225,N_7317);
nor U7560 (N_7560,N_7280,N_7360);
or U7561 (N_7561,N_7227,N_7365);
xor U7562 (N_7562,N_7329,N_7217);
and U7563 (N_7563,N_7334,N_7212);
xnor U7564 (N_7564,N_7338,N_7201);
or U7565 (N_7565,N_7238,N_7353);
or U7566 (N_7566,N_7242,N_7352);
nand U7567 (N_7567,N_7394,N_7287);
and U7568 (N_7568,N_7294,N_7315);
or U7569 (N_7569,N_7236,N_7216);
nor U7570 (N_7570,N_7328,N_7330);
and U7571 (N_7571,N_7339,N_7320);
xnor U7572 (N_7572,N_7310,N_7209);
or U7573 (N_7573,N_7274,N_7210);
xor U7574 (N_7574,N_7216,N_7251);
xnor U7575 (N_7575,N_7256,N_7338);
nand U7576 (N_7576,N_7236,N_7238);
and U7577 (N_7577,N_7263,N_7202);
nor U7578 (N_7578,N_7382,N_7306);
or U7579 (N_7579,N_7312,N_7385);
nand U7580 (N_7580,N_7272,N_7271);
nand U7581 (N_7581,N_7393,N_7326);
xnor U7582 (N_7582,N_7271,N_7315);
xnor U7583 (N_7583,N_7326,N_7240);
nor U7584 (N_7584,N_7308,N_7399);
nor U7585 (N_7585,N_7213,N_7293);
xnor U7586 (N_7586,N_7367,N_7368);
xnor U7587 (N_7587,N_7359,N_7292);
or U7588 (N_7588,N_7355,N_7279);
xor U7589 (N_7589,N_7365,N_7350);
or U7590 (N_7590,N_7260,N_7394);
and U7591 (N_7591,N_7221,N_7369);
nor U7592 (N_7592,N_7292,N_7273);
nand U7593 (N_7593,N_7248,N_7237);
xor U7594 (N_7594,N_7304,N_7221);
or U7595 (N_7595,N_7327,N_7373);
and U7596 (N_7596,N_7398,N_7278);
xnor U7597 (N_7597,N_7218,N_7271);
xor U7598 (N_7598,N_7394,N_7276);
xor U7599 (N_7599,N_7317,N_7266);
xnor U7600 (N_7600,N_7539,N_7470);
or U7601 (N_7601,N_7466,N_7512);
nand U7602 (N_7602,N_7422,N_7586);
or U7603 (N_7603,N_7542,N_7570);
and U7604 (N_7604,N_7562,N_7577);
nor U7605 (N_7605,N_7554,N_7482);
and U7606 (N_7606,N_7536,N_7450);
nand U7607 (N_7607,N_7434,N_7518);
nand U7608 (N_7608,N_7524,N_7533);
or U7609 (N_7609,N_7568,N_7493);
nand U7610 (N_7610,N_7495,N_7447);
nand U7611 (N_7611,N_7578,N_7448);
nor U7612 (N_7612,N_7544,N_7441);
and U7613 (N_7613,N_7436,N_7552);
or U7614 (N_7614,N_7589,N_7430);
and U7615 (N_7615,N_7445,N_7515);
xnor U7616 (N_7616,N_7432,N_7453);
nor U7617 (N_7617,N_7549,N_7507);
nor U7618 (N_7618,N_7464,N_7573);
nand U7619 (N_7619,N_7476,N_7587);
nand U7620 (N_7620,N_7560,N_7597);
nand U7621 (N_7621,N_7528,N_7474);
nor U7622 (N_7622,N_7510,N_7410);
and U7623 (N_7623,N_7460,N_7529);
or U7624 (N_7624,N_7485,N_7545);
or U7625 (N_7625,N_7576,N_7462);
and U7626 (N_7626,N_7593,N_7417);
nor U7627 (N_7627,N_7420,N_7563);
nor U7628 (N_7628,N_7402,N_7532);
nand U7629 (N_7629,N_7497,N_7550);
and U7630 (N_7630,N_7547,N_7513);
or U7631 (N_7631,N_7449,N_7592);
xor U7632 (N_7632,N_7483,N_7501);
and U7633 (N_7633,N_7456,N_7522);
nor U7634 (N_7634,N_7585,N_7454);
xnor U7635 (N_7635,N_7595,N_7408);
and U7636 (N_7636,N_7463,N_7440);
or U7637 (N_7637,N_7409,N_7411);
nor U7638 (N_7638,N_7574,N_7559);
nand U7639 (N_7639,N_7519,N_7484);
nor U7640 (N_7640,N_7413,N_7553);
nor U7641 (N_7641,N_7525,N_7492);
nor U7642 (N_7642,N_7582,N_7543);
or U7643 (N_7643,N_7433,N_7534);
xor U7644 (N_7644,N_7407,N_7516);
or U7645 (N_7645,N_7491,N_7479);
xor U7646 (N_7646,N_7455,N_7509);
nand U7647 (N_7647,N_7506,N_7467);
xor U7648 (N_7648,N_7451,N_7594);
and U7649 (N_7649,N_7469,N_7517);
nand U7650 (N_7650,N_7588,N_7425);
or U7651 (N_7651,N_7403,N_7555);
and U7652 (N_7652,N_7489,N_7500);
xnor U7653 (N_7653,N_7535,N_7527);
nor U7654 (N_7654,N_7598,N_7400);
nand U7655 (N_7655,N_7406,N_7405);
nor U7656 (N_7656,N_7514,N_7590);
nand U7657 (N_7657,N_7404,N_7546);
or U7658 (N_7658,N_7531,N_7414);
nand U7659 (N_7659,N_7478,N_7472);
nand U7660 (N_7660,N_7442,N_7591);
xnor U7661 (N_7661,N_7488,N_7438);
xnor U7662 (N_7662,N_7566,N_7538);
or U7663 (N_7663,N_7477,N_7480);
xor U7664 (N_7664,N_7557,N_7583);
and U7665 (N_7665,N_7523,N_7580);
xor U7666 (N_7666,N_7599,N_7428);
nor U7667 (N_7667,N_7426,N_7511);
or U7668 (N_7668,N_7429,N_7471);
nor U7669 (N_7669,N_7446,N_7461);
and U7670 (N_7670,N_7494,N_7558);
nor U7671 (N_7671,N_7575,N_7412);
or U7672 (N_7672,N_7490,N_7496);
or U7673 (N_7673,N_7564,N_7569);
and U7674 (N_7674,N_7526,N_7435);
nor U7675 (N_7675,N_7416,N_7502);
or U7676 (N_7676,N_7537,N_7548);
xor U7677 (N_7677,N_7581,N_7443);
nand U7678 (N_7678,N_7540,N_7505);
and U7679 (N_7679,N_7458,N_7551);
xnor U7680 (N_7680,N_7596,N_7459);
and U7681 (N_7681,N_7424,N_7475);
nor U7682 (N_7682,N_7561,N_7465);
or U7683 (N_7683,N_7423,N_7401);
and U7684 (N_7684,N_7541,N_7521);
or U7685 (N_7685,N_7503,N_7439);
nor U7686 (N_7686,N_7579,N_7571);
xnor U7687 (N_7687,N_7473,N_7486);
and U7688 (N_7688,N_7415,N_7481);
nor U7689 (N_7689,N_7437,N_7508);
nand U7690 (N_7690,N_7504,N_7567);
or U7691 (N_7691,N_7498,N_7520);
nand U7692 (N_7692,N_7444,N_7418);
and U7693 (N_7693,N_7572,N_7431);
xor U7694 (N_7694,N_7584,N_7457);
xnor U7695 (N_7695,N_7421,N_7487);
and U7696 (N_7696,N_7419,N_7499);
nand U7697 (N_7697,N_7427,N_7565);
and U7698 (N_7698,N_7530,N_7556);
nor U7699 (N_7699,N_7468,N_7452);
and U7700 (N_7700,N_7567,N_7412);
or U7701 (N_7701,N_7411,N_7408);
nand U7702 (N_7702,N_7597,N_7423);
or U7703 (N_7703,N_7484,N_7580);
and U7704 (N_7704,N_7450,N_7454);
nand U7705 (N_7705,N_7410,N_7528);
or U7706 (N_7706,N_7447,N_7429);
nand U7707 (N_7707,N_7581,N_7474);
nor U7708 (N_7708,N_7421,N_7491);
or U7709 (N_7709,N_7409,N_7553);
and U7710 (N_7710,N_7503,N_7446);
or U7711 (N_7711,N_7421,N_7554);
xnor U7712 (N_7712,N_7430,N_7417);
nand U7713 (N_7713,N_7419,N_7429);
xnor U7714 (N_7714,N_7438,N_7510);
xor U7715 (N_7715,N_7450,N_7431);
and U7716 (N_7716,N_7471,N_7548);
xor U7717 (N_7717,N_7595,N_7597);
nand U7718 (N_7718,N_7419,N_7552);
xor U7719 (N_7719,N_7499,N_7447);
or U7720 (N_7720,N_7404,N_7593);
or U7721 (N_7721,N_7416,N_7512);
nand U7722 (N_7722,N_7470,N_7535);
and U7723 (N_7723,N_7485,N_7401);
nand U7724 (N_7724,N_7594,N_7555);
nor U7725 (N_7725,N_7521,N_7450);
xnor U7726 (N_7726,N_7456,N_7520);
or U7727 (N_7727,N_7467,N_7521);
or U7728 (N_7728,N_7598,N_7504);
and U7729 (N_7729,N_7573,N_7442);
xor U7730 (N_7730,N_7524,N_7585);
nor U7731 (N_7731,N_7587,N_7456);
xor U7732 (N_7732,N_7434,N_7529);
or U7733 (N_7733,N_7546,N_7596);
or U7734 (N_7734,N_7571,N_7540);
or U7735 (N_7735,N_7589,N_7532);
xor U7736 (N_7736,N_7584,N_7558);
nor U7737 (N_7737,N_7401,N_7492);
xnor U7738 (N_7738,N_7422,N_7541);
nor U7739 (N_7739,N_7506,N_7495);
and U7740 (N_7740,N_7446,N_7501);
nor U7741 (N_7741,N_7409,N_7477);
xor U7742 (N_7742,N_7455,N_7448);
and U7743 (N_7743,N_7509,N_7495);
or U7744 (N_7744,N_7496,N_7553);
nand U7745 (N_7745,N_7407,N_7481);
xor U7746 (N_7746,N_7497,N_7493);
xnor U7747 (N_7747,N_7548,N_7549);
xnor U7748 (N_7748,N_7483,N_7587);
nor U7749 (N_7749,N_7541,N_7576);
nand U7750 (N_7750,N_7433,N_7411);
or U7751 (N_7751,N_7492,N_7580);
nor U7752 (N_7752,N_7459,N_7420);
and U7753 (N_7753,N_7546,N_7587);
or U7754 (N_7754,N_7506,N_7585);
or U7755 (N_7755,N_7557,N_7464);
xor U7756 (N_7756,N_7414,N_7404);
or U7757 (N_7757,N_7528,N_7585);
nand U7758 (N_7758,N_7507,N_7442);
nor U7759 (N_7759,N_7461,N_7423);
nand U7760 (N_7760,N_7436,N_7558);
xor U7761 (N_7761,N_7526,N_7429);
and U7762 (N_7762,N_7580,N_7443);
or U7763 (N_7763,N_7591,N_7471);
and U7764 (N_7764,N_7475,N_7588);
nand U7765 (N_7765,N_7461,N_7587);
or U7766 (N_7766,N_7571,N_7527);
or U7767 (N_7767,N_7485,N_7441);
and U7768 (N_7768,N_7428,N_7591);
or U7769 (N_7769,N_7466,N_7472);
and U7770 (N_7770,N_7585,N_7403);
nor U7771 (N_7771,N_7452,N_7429);
or U7772 (N_7772,N_7484,N_7514);
and U7773 (N_7773,N_7428,N_7552);
or U7774 (N_7774,N_7590,N_7516);
xor U7775 (N_7775,N_7559,N_7445);
xor U7776 (N_7776,N_7428,N_7454);
xor U7777 (N_7777,N_7481,N_7580);
xor U7778 (N_7778,N_7488,N_7504);
xnor U7779 (N_7779,N_7405,N_7543);
and U7780 (N_7780,N_7447,N_7564);
and U7781 (N_7781,N_7595,N_7445);
xnor U7782 (N_7782,N_7591,N_7526);
or U7783 (N_7783,N_7536,N_7472);
nand U7784 (N_7784,N_7466,N_7569);
xnor U7785 (N_7785,N_7473,N_7519);
nand U7786 (N_7786,N_7403,N_7457);
or U7787 (N_7787,N_7598,N_7413);
nor U7788 (N_7788,N_7519,N_7557);
nor U7789 (N_7789,N_7523,N_7448);
and U7790 (N_7790,N_7510,N_7411);
nor U7791 (N_7791,N_7431,N_7548);
nand U7792 (N_7792,N_7512,N_7407);
and U7793 (N_7793,N_7599,N_7505);
or U7794 (N_7794,N_7518,N_7403);
nand U7795 (N_7795,N_7582,N_7549);
nand U7796 (N_7796,N_7473,N_7447);
xnor U7797 (N_7797,N_7568,N_7428);
xor U7798 (N_7798,N_7577,N_7561);
nand U7799 (N_7799,N_7571,N_7552);
or U7800 (N_7800,N_7679,N_7762);
or U7801 (N_7801,N_7722,N_7748);
nand U7802 (N_7802,N_7646,N_7791);
and U7803 (N_7803,N_7671,N_7729);
nand U7804 (N_7804,N_7642,N_7621);
or U7805 (N_7805,N_7758,N_7647);
xor U7806 (N_7806,N_7780,N_7784);
or U7807 (N_7807,N_7604,N_7742);
nand U7808 (N_7808,N_7707,N_7640);
nand U7809 (N_7809,N_7697,N_7751);
xor U7810 (N_7810,N_7605,N_7764);
nand U7811 (N_7811,N_7656,N_7743);
nor U7812 (N_7812,N_7721,N_7714);
nor U7813 (N_7813,N_7794,N_7619);
or U7814 (N_7814,N_7644,N_7783);
and U7815 (N_7815,N_7772,N_7725);
nand U7816 (N_7816,N_7643,N_7745);
xnor U7817 (N_7817,N_7740,N_7685);
nand U7818 (N_7818,N_7688,N_7717);
and U7819 (N_7819,N_7723,N_7635);
xor U7820 (N_7820,N_7789,N_7606);
nor U7821 (N_7821,N_7645,N_7728);
and U7822 (N_7822,N_7662,N_7608);
xnor U7823 (N_7823,N_7765,N_7713);
and U7824 (N_7824,N_7797,N_7746);
and U7825 (N_7825,N_7655,N_7790);
nor U7826 (N_7826,N_7691,N_7755);
nor U7827 (N_7827,N_7613,N_7632);
xnor U7828 (N_7828,N_7630,N_7682);
nor U7829 (N_7829,N_7736,N_7607);
or U7830 (N_7830,N_7694,N_7749);
nor U7831 (N_7831,N_7704,N_7684);
and U7832 (N_7832,N_7788,N_7712);
nor U7833 (N_7833,N_7686,N_7767);
or U7834 (N_7834,N_7703,N_7770);
nand U7835 (N_7835,N_7663,N_7719);
and U7836 (N_7836,N_7711,N_7610);
xor U7837 (N_7837,N_7775,N_7733);
and U7838 (N_7838,N_7678,N_7673);
and U7839 (N_7839,N_7796,N_7744);
xnor U7840 (N_7840,N_7787,N_7638);
nor U7841 (N_7841,N_7681,N_7661);
nor U7842 (N_7842,N_7617,N_7763);
or U7843 (N_7843,N_7648,N_7739);
or U7844 (N_7844,N_7603,N_7698);
or U7845 (N_7845,N_7738,N_7750);
nor U7846 (N_7846,N_7651,N_7676);
nand U7847 (N_7847,N_7776,N_7620);
or U7848 (N_7848,N_7727,N_7702);
nand U7849 (N_7849,N_7761,N_7675);
xnor U7850 (N_7850,N_7677,N_7654);
xnor U7851 (N_7851,N_7668,N_7799);
xor U7852 (N_7852,N_7768,N_7705);
nand U7853 (N_7853,N_7720,N_7641);
nand U7854 (N_7854,N_7609,N_7771);
xnor U7855 (N_7855,N_7618,N_7759);
xnor U7856 (N_7856,N_7756,N_7693);
or U7857 (N_7857,N_7670,N_7760);
xor U7858 (N_7858,N_7669,N_7634);
xor U7859 (N_7859,N_7664,N_7601);
or U7860 (N_7860,N_7600,N_7735);
and U7861 (N_7861,N_7696,N_7622);
nor U7862 (N_7862,N_7710,N_7773);
xor U7863 (N_7863,N_7701,N_7753);
nor U7864 (N_7864,N_7674,N_7629);
nor U7865 (N_7865,N_7631,N_7659);
nor U7866 (N_7866,N_7737,N_7666);
nand U7867 (N_7867,N_7726,N_7611);
nor U7868 (N_7868,N_7754,N_7602);
or U7869 (N_7869,N_7724,N_7667);
nor U7870 (N_7870,N_7706,N_7769);
or U7871 (N_7871,N_7653,N_7782);
or U7872 (N_7872,N_7615,N_7625);
and U7873 (N_7873,N_7699,N_7792);
nor U7874 (N_7874,N_7779,N_7660);
or U7875 (N_7875,N_7716,N_7777);
nand U7876 (N_7876,N_7626,N_7757);
nor U7877 (N_7877,N_7612,N_7683);
or U7878 (N_7878,N_7623,N_7627);
xor U7879 (N_7879,N_7628,N_7734);
nand U7880 (N_7880,N_7731,N_7639);
and U7881 (N_7881,N_7774,N_7690);
and U7882 (N_7882,N_7657,N_7730);
and U7883 (N_7883,N_7700,N_7650);
nand U7884 (N_7884,N_7658,N_7793);
xor U7885 (N_7885,N_7718,N_7616);
nor U7886 (N_7886,N_7778,N_7692);
nor U7887 (N_7887,N_7732,N_7614);
nand U7888 (N_7888,N_7785,N_7747);
and U7889 (N_7889,N_7665,N_7680);
nand U7890 (N_7890,N_7689,N_7708);
or U7891 (N_7891,N_7795,N_7786);
and U7892 (N_7892,N_7637,N_7649);
xor U7893 (N_7893,N_7636,N_7741);
nor U7894 (N_7894,N_7715,N_7709);
or U7895 (N_7895,N_7695,N_7652);
and U7896 (N_7896,N_7798,N_7752);
nor U7897 (N_7897,N_7672,N_7766);
nor U7898 (N_7898,N_7781,N_7633);
and U7899 (N_7899,N_7687,N_7624);
nand U7900 (N_7900,N_7786,N_7729);
nor U7901 (N_7901,N_7604,N_7766);
xnor U7902 (N_7902,N_7645,N_7754);
xor U7903 (N_7903,N_7685,N_7667);
and U7904 (N_7904,N_7646,N_7686);
xor U7905 (N_7905,N_7705,N_7767);
nor U7906 (N_7906,N_7612,N_7624);
and U7907 (N_7907,N_7775,N_7660);
nor U7908 (N_7908,N_7609,N_7678);
xnor U7909 (N_7909,N_7710,N_7737);
nand U7910 (N_7910,N_7643,N_7736);
nand U7911 (N_7911,N_7649,N_7645);
nor U7912 (N_7912,N_7739,N_7612);
and U7913 (N_7913,N_7630,N_7661);
and U7914 (N_7914,N_7794,N_7669);
nor U7915 (N_7915,N_7740,N_7748);
nor U7916 (N_7916,N_7658,N_7669);
xor U7917 (N_7917,N_7656,N_7701);
nand U7918 (N_7918,N_7791,N_7635);
and U7919 (N_7919,N_7746,N_7716);
xnor U7920 (N_7920,N_7788,N_7640);
xor U7921 (N_7921,N_7709,N_7785);
nor U7922 (N_7922,N_7725,N_7775);
or U7923 (N_7923,N_7713,N_7683);
or U7924 (N_7924,N_7757,N_7702);
and U7925 (N_7925,N_7797,N_7674);
and U7926 (N_7926,N_7744,N_7729);
or U7927 (N_7927,N_7709,N_7795);
and U7928 (N_7928,N_7731,N_7749);
or U7929 (N_7929,N_7658,N_7767);
nand U7930 (N_7930,N_7654,N_7754);
nand U7931 (N_7931,N_7654,N_7780);
or U7932 (N_7932,N_7607,N_7610);
nor U7933 (N_7933,N_7720,N_7699);
nor U7934 (N_7934,N_7733,N_7747);
and U7935 (N_7935,N_7794,N_7684);
and U7936 (N_7936,N_7792,N_7751);
and U7937 (N_7937,N_7745,N_7684);
nand U7938 (N_7938,N_7665,N_7613);
xnor U7939 (N_7939,N_7798,N_7688);
xor U7940 (N_7940,N_7679,N_7741);
nand U7941 (N_7941,N_7650,N_7662);
xnor U7942 (N_7942,N_7758,N_7628);
or U7943 (N_7943,N_7757,N_7779);
and U7944 (N_7944,N_7707,N_7616);
nand U7945 (N_7945,N_7605,N_7676);
nand U7946 (N_7946,N_7645,N_7656);
and U7947 (N_7947,N_7717,N_7635);
nor U7948 (N_7948,N_7616,N_7627);
xnor U7949 (N_7949,N_7624,N_7617);
nand U7950 (N_7950,N_7699,N_7671);
or U7951 (N_7951,N_7702,N_7796);
xnor U7952 (N_7952,N_7740,N_7727);
nand U7953 (N_7953,N_7723,N_7775);
xnor U7954 (N_7954,N_7683,N_7761);
or U7955 (N_7955,N_7650,N_7718);
and U7956 (N_7956,N_7693,N_7720);
nor U7957 (N_7957,N_7674,N_7683);
nand U7958 (N_7958,N_7675,N_7732);
nand U7959 (N_7959,N_7728,N_7626);
nor U7960 (N_7960,N_7608,N_7657);
nand U7961 (N_7961,N_7795,N_7622);
nand U7962 (N_7962,N_7719,N_7642);
and U7963 (N_7963,N_7745,N_7698);
or U7964 (N_7964,N_7643,N_7650);
nand U7965 (N_7965,N_7704,N_7645);
xnor U7966 (N_7966,N_7713,N_7778);
and U7967 (N_7967,N_7680,N_7663);
or U7968 (N_7968,N_7626,N_7700);
or U7969 (N_7969,N_7660,N_7680);
nor U7970 (N_7970,N_7731,N_7720);
nand U7971 (N_7971,N_7771,N_7755);
or U7972 (N_7972,N_7715,N_7747);
or U7973 (N_7973,N_7721,N_7666);
and U7974 (N_7974,N_7628,N_7765);
nor U7975 (N_7975,N_7677,N_7675);
or U7976 (N_7976,N_7745,N_7717);
nor U7977 (N_7977,N_7725,N_7628);
nor U7978 (N_7978,N_7790,N_7607);
and U7979 (N_7979,N_7619,N_7646);
or U7980 (N_7980,N_7776,N_7628);
nand U7981 (N_7981,N_7711,N_7783);
or U7982 (N_7982,N_7798,N_7675);
nor U7983 (N_7983,N_7724,N_7793);
and U7984 (N_7984,N_7691,N_7762);
and U7985 (N_7985,N_7775,N_7680);
and U7986 (N_7986,N_7644,N_7755);
nor U7987 (N_7987,N_7650,N_7633);
nand U7988 (N_7988,N_7626,N_7742);
and U7989 (N_7989,N_7613,N_7766);
and U7990 (N_7990,N_7743,N_7651);
xnor U7991 (N_7991,N_7640,N_7708);
or U7992 (N_7992,N_7766,N_7706);
and U7993 (N_7993,N_7777,N_7787);
or U7994 (N_7994,N_7714,N_7635);
or U7995 (N_7995,N_7664,N_7680);
nand U7996 (N_7996,N_7683,N_7601);
nand U7997 (N_7997,N_7702,N_7772);
xnor U7998 (N_7998,N_7623,N_7687);
and U7999 (N_7999,N_7665,N_7626);
nor U8000 (N_8000,N_7915,N_7893);
and U8001 (N_8001,N_7933,N_7963);
and U8002 (N_8002,N_7871,N_7803);
nand U8003 (N_8003,N_7868,N_7802);
xor U8004 (N_8004,N_7907,N_7946);
and U8005 (N_8005,N_7926,N_7991);
or U8006 (N_8006,N_7845,N_7984);
and U8007 (N_8007,N_7920,N_7913);
or U8008 (N_8008,N_7858,N_7807);
nor U8009 (N_8009,N_7954,N_7885);
xnor U8010 (N_8010,N_7844,N_7904);
xnor U8011 (N_8011,N_7959,N_7874);
or U8012 (N_8012,N_7834,N_7811);
or U8013 (N_8013,N_7970,N_7960);
nor U8014 (N_8014,N_7979,N_7843);
and U8015 (N_8015,N_7875,N_7804);
xnor U8016 (N_8016,N_7905,N_7941);
and U8017 (N_8017,N_7854,N_7829);
nand U8018 (N_8018,N_7892,N_7869);
nand U8019 (N_8019,N_7997,N_7870);
xnor U8020 (N_8020,N_7852,N_7899);
nand U8021 (N_8021,N_7987,N_7925);
nor U8022 (N_8022,N_7894,N_7949);
nor U8023 (N_8023,N_7832,N_7932);
and U8024 (N_8024,N_7873,N_7888);
nand U8025 (N_8025,N_7918,N_7817);
and U8026 (N_8026,N_7988,N_7867);
or U8027 (N_8027,N_7831,N_7883);
nor U8028 (N_8028,N_7989,N_7996);
nand U8029 (N_8029,N_7897,N_7839);
and U8030 (N_8030,N_7809,N_7850);
nand U8031 (N_8031,N_7805,N_7895);
and U8032 (N_8032,N_7848,N_7981);
nand U8033 (N_8033,N_7815,N_7808);
or U8034 (N_8034,N_7940,N_7825);
nor U8035 (N_8035,N_7964,N_7967);
nor U8036 (N_8036,N_7813,N_7990);
nor U8037 (N_8037,N_7857,N_7966);
or U8038 (N_8038,N_7955,N_7865);
xnor U8039 (N_8039,N_7821,N_7900);
and U8040 (N_8040,N_7911,N_7968);
nor U8041 (N_8041,N_7812,N_7923);
nand U8042 (N_8042,N_7945,N_7800);
nor U8043 (N_8043,N_7898,N_7863);
and U8044 (N_8044,N_7950,N_7826);
nor U8045 (N_8045,N_7801,N_7971);
nand U8046 (N_8046,N_7973,N_7806);
or U8047 (N_8047,N_7994,N_7962);
nor U8048 (N_8048,N_7992,N_7939);
nor U8049 (N_8049,N_7935,N_7881);
nand U8050 (N_8050,N_7929,N_7853);
or U8051 (N_8051,N_7847,N_7878);
nor U8052 (N_8052,N_7951,N_7956);
nor U8053 (N_8053,N_7995,N_7903);
and U8054 (N_8054,N_7879,N_7977);
nand U8055 (N_8055,N_7985,N_7891);
nor U8056 (N_8056,N_7934,N_7846);
and U8057 (N_8057,N_7969,N_7928);
nand U8058 (N_8058,N_7910,N_7818);
or U8059 (N_8059,N_7972,N_7835);
nor U8060 (N_8060,N_7982,N_7974);
xnor U8061 (N_8061,N_7872,N_7849);
xor U8062 (N_8062,N_7855,N_7828);
nand U8063 (N_8063,N_7830,N_7851);
and U8064 (N_8064,N_7986,N_7975);
or U8065 (N_8065,N_7842,N_7993);
nor U8066 (N_8066,N_7957,N_7917);
xnor U8067 (N_8067,N_7944,N_7983);
or U8068 (N_8068,N_7833,N_7901);
and U8069 (N_8069,N_7876,N_7936);
nor U8070 (N_8070,N_7823,N_7998);
and U8071 (N_8071,N_7930,N_7884);
nor U8072 (N_8072,N_7942,N_7916);
nand U8073 (N_8073,N_7919,N_7860);
xor U8074 (N_8074,N_7827,N_7877);
nand U8075 (N_8075,N_7927,N_7864);
xor U8076 (N_8076,N_7837,N_7906);
and U8077 (N_8077,N_7948,N_7822);
and U8078 (N_8078,N_7965,N_7943);
nand U8079 (N_8079,N_7947,N_7938);
nand U8080 (N_8080,N_7882,N_7931);
and U8081 (N_8081,N_7980,N_7838);
xor U8082 (N_8082,N_7922,N_7810);
nand U8083 (N_8083,N_7889,N_7937);
and U8084 (N_8084,N_7958,N_7924);
or U8085 (N_8085,N_7909,N_7921);
and U8086 (N_8086,N_7914,N_7912);
xnor U8087 (N_8087,N_7976,N_7880);
and U8088 (N_8088,N_7896,N_7861);
and U8089 (N_8089,N_7859,N_7814);
and U8090 (N_8090,N_7816,N_7820);
xnor U8091 (N_8091,N_7952,N_7887);
nor U8092 (N_8092,N_7902,N_7908);
xnor U8093 (N_8093,N_7836,N_7856);
and U8094 (N_8094,N_7886,N_7824);
nor U8095 (N_8095,N_7978,N_7819);
or U8096 (N_8096,N_7999,N_7862);
nor U8097 (N_8097,N_7953,N_7840);
nand U8098 (N_8098,N_7841,N_7961);
xnor U8099 (N_8099,N_7866,N_7890);
xnor U8100 (N_8100,N_7916,N_7878);
nor U8101 (N_8101,N_7918,N_7847);
and U8102 (N_8102,N_7938,N_7832);
nor U8103 (N_8103,N_7998,N_7852);
xor U8104 (N_8104,N_7804,N_7887);
and U8105 (N_8105,N_7966,N_7827);
xor U8106 (N_8106,N_7982,N_7847);
nand U8107 (N_8107,N_7911,N_7973);
or U8108 (N_8108,N_7836,N_7917);
nand U8109 (N_8109,N_7993,N_7976);
nand U8110 (N_8110,N_7848,N_7993);
and U8111 (N_8111,N_7928,N_7958);
nand U8112 (N_8112,N_7988,N_7821);
or U8113 (N_8113,N_7899,N_7942);
and U8114 (N_8114,N_7932,N_7960);
nor U8115 (N_8115,N_7899,N_7997);
nor U8116 (N_8116,N_7912,N_7802);
xor U8117 (N_8117,N_7990,N_7833);
xor U8118 (N_8118,N_7929,N_7917);
or U8119 (N_8119,N_7869,N_7945);
or U8120 (N_8120,N_7976,N_7932);
nand U8121 (N_8121,N_7975,N_7842);
xor U8122 (N_8122,N_7965,N_7967);
xnor U8123 (N_8123,N_7819,N_7887);
and U8124 (N_8124,N_7883,N_7920);
or U8125 (N_8125,N_7876,N_7942);
or U8126 (N_8126,N_7919,N_7964);
or U8127 (N_8127,N_7952,N_7847);
and U8128 (N_8128,N_7908,N_7879);
or U8129 (N_8129,N_7918,N_7856);
nor U8130 (N_8130,N_7907,N_7942);
or U8131 (N_8131,N_7823,N_7966);
xor U8132 (N_8132,N_7976,N_7980);
xor U8133 (N_8133,N_7807,N_7985);
and U8134 (N_8134,N_7897,N_7828);
xnor U8135 (N_8135,N_7942,N_7901);
nand U8136 (N_8136,N_7834,N_7965);
xnor U8137 (N_8137,N_7982,N_7812);
xor U8138 (N_8138,N_7872,N_7839);
nor U8139 (N_8139,N_7867,N_7881);
nor U8140 (N_8140,N_7997,N_7961);
xnor U8141 (N_8141,N_7828,N_7884);
nor U8142 (N_8142,N_7846,N_7918);
xor U8143 (N_8143,N_7950,N_7892);
nor U8144 (N_8144,N_7853,N_7825);
nor U8145 (N_8145,N_7816,N_7953);
xnor U8146 (N_8146,N_7880,N_7808);
or U8147 (N_8147,N_7804,N_7815);
and U8148 (N_8148,N_7956,N_7969);
nor U8149 (N_8149,N_7951,N_7896);
nand U8150 (N_8150,N_7899,N_7894);
xnor U8151 (N_8151,N_7815,N_7826);
nor U8152 (N_8152,N_7800,N_7919);
or U8153 (N_8153,N_7856,N_7909);
or U8154 (N_8154,N_7998,N_7832);
and U8155 (N_8155,N_7802,N_7800);
and U8156 (N_8156,N_7870,N_7827);
xor U8157 (N_8157,N_7989,N_7848);
nand U8158 (N_8158,N_7898,N_7937);
nand U8159 (N_8159,N_7983,N_7943);
and U8160 (N_8160,N_7997,N_7933);
xnor U8161 (N_8161,N_7958,N_7988);
nor U8162 (N_8162,N_7925,N_7842);
and U8163 (N_8163,N_7906,N_7845);
xnor U8164 (N_8164,N_7805,N_7916);
nor U8165 (N_8165,N_7999,N_7986);
or U8166 (N_8166,N_7964,N_7925);
or U8167 (N_8167,N_7998,N_7919);
nor U8168 (N_8168,N_7821,N_7878);
and U8169 (N_8169,N_7853,N_7972);
nor U8170 (N_8170,N_7996,N_7880);
xnor U8171 (N_8171,N_7978,N_7859);
xnor U8172 (N_8172,N_7919,N_7906);
xor U8173 (N_8173,N_7936,N_7860);
nor U8174 (N_8174,N_7980,N_7859);
nor U8175 (N_8175,N_7806,N_7816);
xnor U8176 (N_8176,N_7868,N_7980);
and U8177 (N_8177,N_7818,N_7886);
or U8178 (N_8178,N_7830,N_7906);
nand U8179 (N_8179,N_7800,N_7924);
nand U8180 (N_8180,N_7877,N_7954);
and U8181 (N_8181,N_7889,N_7814);
nor U8182 (N_8182,N_7999,N_7996);
nand U8183 (N_8183,N_7849,N_7938);
or U8184 (N_8184,N_7905,N_7830);
and U8185 (N_8185,N_7873,N_7953);
nor U8186 (N_8186,N_7850,N_7848);
xor U8187 (N_8187,N_7930,N_7815);
nand U8188 (N_8188,N_7970,N_7848);
and U8189 (N_8189,N_7877,N_7861);
nor U8190 (N_8190,N_7878,N_7897);
nand U8191 (N_8191,N_7827,N_7894);
nor U8192 (N_8192,N_7824,N_7816);
or U8193 (N_8193,N_7919,N_7929);
nand U8194 (N_8194,N_7893,N_7829);
xnor U8195 (N_8195,N_7971,N_7802);
nor U8196 (N_8196,N_7911,N_7962);
nand U8197 (N_8197,N_7909,N_7998);
or U8198 (N_8198,N_7931,N_7927);
xnor U8199 (N_8199,N_7989,N_7890);
nor U8200 (N_8200,N_8013,N_8053);
or U8201 (N_8201,N_8178,N_8080);
xor U8202 (N_8202,N_8078,N_8012);
nand U8203 (N_8203,N_8158,N_8063);
xor U8204 (N_8204,N_8108,N_8129);
nor U8205 (N_8205,N_8003,N_8015);
nand U8206 (N_8206,N_8137,N_8112);
xor U8207 (N_8207,N_8054,N_8011);
or U8208 (N_8208,N_8002,N_8185);
xor U8209 (N_8209,N_8183,N_8181);
and U8210 (N_8210,N_8096,N_8136);
xnor U8211 (N_8211,N_8088,N_8143);
nand U8212 (N_8212,N_8024,N_8121);
and U8213 (N_8213,N_8120,N_8174);
and U8214 (N_8214,N_8028,N_8043);
and U8215 (N_8215,N_8031,N_8020);
nand U8216 (N_8216,N_8072,N_8066);
xor U8217 (N_8217,N_8099,N_8170);
and U8218 (N_8218,N_8191,N_8032);
xnor U8219 (N_8219,N_8139,N_8172);
nand U8220 (N_8220,N_8073,N_8154);
xnor U8221 (N_8221,N_8070,N_8189);
nand U8222 (N_8222,N_8091,N_8165);
nor U8223 (N_8223,N_8153,N_8017);
or U8224 (N_8224,N_8087,N_8106);
nor U8225 (N_8225,N_8037,N_8075);
and U8226 (N_8226,N_8167,N_8155);
and U8227 (N_8227,N_8022,N_8009);
nor U8228 (N_8228,N_8023,N_8140);
nand U8229 (N_8229,N_8190,N_8152);
or U8230 (N_8230,N_8019,N_8138);
nor U8231 (N_8231,N_8109,N_8094);
and U8232 (N_8232,N_8194,N_8085);
nor U8233 (N_8233,N_8059,N_8175);
nor U8234 (N_8234,N_8064,N_8057);
nor U8235 (N_8235,N_8030,N_8156);
nand U8236 (N_8236,N_8142,N_8097);
xnor U8237 (N_8237,N_8164,N_8042);
xnor U8238 (N_8238,N_8065,N_8114);
or U8239 (N_8239,N_8104,N_8103);
xnor U8240 (N_8240,N_8192,N_8118);
and U8241 (N_8241,N_8068,N_8025);
or U8242 (N_8242,N_8117,N_8010);
or U8243 (N_8243,N_8145,N_8000);
nor U8244 (N_8244,N_8041,N_8199);
nor U8245 (N_8245,N_8149,N_8071);
or U8246 (N_8246,N_8034,N_8007);
nand U8247 (N_8247,N_8004,N_8040);
nand U8248 (N_8248,N_8069,N_8067);
and U8249 (N_8249,N_8079,N_8131);
nor U8250 (N_8250,N_8123,N_8049);
nor U8251 (N_8251,N_8127,N_8027);
nor U8252 (N_8252,N_8074,N_8083);
nand U8253 (N_8253,N_8081,N_8005);
xor U8254 (N_8254,N_8124,N_8111);
xor U8255 (N_8255,N_8026,N_8001);
nor U8256 (N_8256,N_8193,N_8048);
and U8257 (N_8257,N_8058,N_8134);
and U8258 (N_8258,N_8126,N_8018);
nor U8259 (N_8259,N_8052,N_8198);
or U8260 (N_8260,N_8029,N_8107);
and U8261 (N_8261,N_8051,N_8162);
xnor U8262 (N_8262,N_8035,N_8195);
nand U8263 (N_8263,N_8014,N_8077);
and U8264 (N_8264,N_8092,N_8100);
or U8265 (N_8265,N_8182,N_8116);
or U8266 (N_8266,N_8179,N_8050);
xnor U8267 (N_8267,N_8146,N_8062);
or U8268 (N_8268,N_8036,N_8188);
nand U8269 (N_8269,N_8060,N_8044);
or U8270 (N_8270,N_8006,N_8095);
nor U8271 (N_8271,N_8122,N_8102);
nand U8272 (N_8272,N_8047,N_8082);
xor U8273 (N_8273,N_8151,N_8105);
or U8274 (N_8274,N_8086,N_8061);
or U8275 (N_8275,N_8159,N_8144);
nor U8276 (N_8276,N_8135,N_8157);
nor U8277 (N_8277,N_8115,N_8177);
nand U8278 (N_8278,N_8110,N_8176);
and U8279 (N_8279,N_8141,N_8113);
nor U8280 (N_8280,N_8090,N_8197);
or U8281 (N_8281,N_8125,N_8171);
xnor U8282 (N_8282,N_8008,N_8130);
nor U8283 (N_8283,N_8147,N_8148);
nor U8284 (N_8284,N_8098,N_8016);
or U8285 (N_8285,N_8045,N_8119);
nand U8286 (N_8286,N_8101,N_8089);
and U8287 (N_8287,N_8021,N_8173);
nor U8288 (N_8288,N_8133,N_8180);
nand U8289 (N_8289,N_8055,N_8128);
or U8290 (N_8290,N_8160,N_8038);
nand U8291 (N_8291,N_8161,N_8163);
xnor U8292 (N_8292,N_8168,N_8166);
and U8293 (N_8293,N_8093,N_8150);
and U8294 (N_8294,N_8046,N_8186);
nand U8295 (N_8295,N_8184,N_8039);
nand U8296 (N_8296,N_8033,N_8187);
nor U8297 (N_8297,N_8056,N_8132);
nand U8298 (N_8298,N_8076,N_8084);
nand U8299 (N_8299,N_8169,N_8196);
xor U8300 (N_8300,N_8072,N_8050);
nor U8301 (N_8301,N_8044,N_8131);
nor U8302 (N_8302,N_8011,N_8146);
nor U8303 (N_8303,N_8016,N_8165);
or U8304 (N_8304,N_8016,N_8176);
and U8305 (N_8305,N_8189,N_8075);
xnor U8306 (N_8306,N_8141,N_8094);
xnor U8307 (N_8307,N_8104,N_8102);
xnor U8308 (N_8308,N_8057,N_8091);
xnor U8309 (N_8309,N_8181,N_8051);
or U8310 (N_8310,N_8185,N_8141);
xnor U8311 (N_8311,N_8173,N_8099);
or U8312 (N_8312,N_8054,N_8100);
or U8313 (N_8313,N_8005,N_8118);
and U8314 (N_8314,N_8017,N_8032);
nor U8315 (N_8315,N_8136,N_8192);
or U8316 (N_8316,N_8123,N_8108);
or U8317 (N_8317,N_8017,N_8159);
nor U8318 (N_8318,N_8135,N_8016);
and U8319 (N_8319,N_8161,N_8008);
nand U8320 (N_8320,N_8079,N_8086);
nand U8321 (N_8321,N_8083,N_8042);
and U8322 (N_8322,N_8008,N_8164);
and U8323 (N_8323,N_8009,N_8159);
or U8324 (N_8324,N_8041,N_8099);
or U8325 (N_8325,N_8070,N_8041);
or U8326 (N_8326,N_8149,N_8056);
nand U8327 (N_8327,N_8014,N_8071);
or U8328 (N_8328,N_8066,N_8123);
nand U8329 (N_8329,N_8099,N_8096);
or U8330 (N_8330,N_8077,N_8150);
or U8331 (N_8331,N_8097,N_8006);
nor U8332 (N_8332,N_8183,N_8146);
or U8333 (N_8333,N_8171,N_8159);
or U8334 (N_8334,N_8060,N_8090);
and U8335 (N_8335,N_8104,N_8147);
or U8336 (N_8336,N_8069,N_8108);
xnor U8337 (N_8337,N_8012,N_8063);
or U8338 (N_8338,N_8177,N_8142);
xor U8339 (N_8339,N_8036,N_8097);
and U8340 (N_8340,N_8194,N_8179);
nor U8341 (N_8341,N_8143,N_8060);
xor U8342 (N_8342,N_8088,N_8172);
nor U8343 (N_8343,N_8040,N_8045);
and U8344 (N_8344,N_8112,N_8058);
nand U8345 (N_8345,N_8005,N_8096);
or U8346 (N_8346,N_8176,N_8069);
nor U8347 (N_8347,N_8072,N_8176);
xnor U8348 (N_8348,N_8042,N_8100);
and U8349 (N_8349,N_8060,N_8174);
or U8350 (N_8350,N_8176,N_8174);
nand U8351 (N_8351,N_8106,N_8119);
nor U8352 (N_8352,N_8138,N_8147);
nor U8353 (N_8353,N_8048,N_8078);
xnor U8354 (N_8354,N_8007,N_8061);
nand U8355 (N_8355,N_8078,N_8070);
and U8356 (N_8356,N_8040,N_8056);
nor U8357 (N_8357,N_8132,N_8169);
nor U8358 (N_8358,N_8068,N_8164);
nand U8359 (N_8359,N_8011,N_8042);
and U8360 (N_8360,N_8195,N_8126);
or U8361 (N_8361,N_8174,N_8077);
nand U8362 (N_8362,N_8115,N_8109);
or U8363 (N_8363,N_8105,N_8152);
nor U8364 (N_8364,N_8148,N_8045);
nand U8365 (N_8365,N_8033,N_8079);
xnor U8366 (N_8366,N_8112,N_8153);
xnor U8367 (N_8367,N_8031,N_8186);
nand U8368 (N_8368,N_8029,N_8059);
or U8369 (N_8369,N_8198,N_8150);
and U8370 (N_8370,N_8059,N_8128);
and U8371 (N_8371,N_8043,N_8130);
nand U8372 (N_8372,N_8040,N_8185);
xor U8373 (N_8373,N_8011,N_8162);
or U8374 (N_8374,N_8065,N_8140);
xnor U8375 (N_8375,N_8011,N_8097);
or U8376 (N_8376,N_8166,N_8025);
nand U8377 (N_8377,N_8038,N_8173);
xnor U8378 (N_8378,N_8150,N_8065);
or U8379 (N_8379,N_8162,N_8158);
xnor U8380 (N_8380,N_8006,N_8150);
xnor U8381 (N_8381,N_8177,N_8015);
and U8382 (N_8382,N_8075,N_8047);
nor U8383 (N_8383,N_8034,N_8013);
nor U8384 (N_8384,N_8085,N_8172);
and U8385 (N_8385,N_8102,N_8160);
and U8386 (N_8386,N_8011,N_8044);
and U8387 (N_8387,N_8112,N_8174);
xnor U8388 (N_8388,N_8016,N_8004);
nand U8389 (N_8389,N_8167,N_8097);
nor U8390 (N_8390,N_8022,N_8139);
or U8391 (N_8391,N_8183,N_8073);
xor U8392 (N_8392,N_8010,N_8161);
or U8393 (N_8393,N_8196,N_8170);
and U8394 (N_8394,N_8029,N_8193);
and U8395 (N_8395,N_8133,N_8009);
nor U8396 (N_8396,N_8006,N_8059);
and U8397 (N_8397,N_8064,N_8033);
nor U8398 (N_8398,N_8127,N_8167);
or U8399 (N_8399,N_8140,N_8194);
or U8400 (N_8400,N_8204,N_8331);
xnor U8401 (N_8401,N_8303,N_8394);
or U8402 (N_8402,N_8320,N_8342);
xnor U8403 (N_8403,N_8212,N_8211);
nand U8404 (N_8404,N_8379,N_8338);
and U8405 (N_8405,N_8213,N_8265);
or U8406 (N_8406,N_8356,N_8294);
nor U8407 (N_8407,N_8366,N_8393);
nand U8408 (N_8408,N_8364,N_8375);
nor U8409 (N_8409,N_8362,N_8226);
nor U8410 (N_8410,N_8233,N_8273);
nor U8411 (N_8411,N_8377,N_8234);
xnor U8412 (N_8412,N_8327,N_8282);
or U8413 (N_8413,N_8229,N_8321);
and U8414 (N_8414,N_8360,N_8358);
or U8415 (N_8415,N_8355,N_8259);
and U8416 (N_8416,N_8383,N_8354);
nand U8417 (N_8417,N_8260,N_8373);
nor U8418 (N_8418,N_8337,N_8242);
nor U8419 (N_8419,N_8370,N_8371);
xnor U8420 (N_8420,N_8230,N_8349);
and U8421 (N_8421,N_8253,N_8220);
or U8422 (N_8422,N_8288,N_8339);
nand U8423 (N_8423,N_8317,N_8348);
and U8424 (N_8424,N_8397,N_8219);
nand U8425 (N_8425,N_8332,N_8315);
and U8426 (N_8426,N_8232,N_8243);
or U8427 (N_8427,N_8334,N_8382);
xnor U8428 (N_8428,N_8245,N_8306);
xor U8429 (N_8429,N_8389,N_8399);
and U8430 (N_8430,N_8308,N_8277);
nor U8431 (N_8431,N_8262,N_8311);
nor U8432 (N_8432,N_8202,N_8221);
or U8433 (N_8433,N_8372,N_8323);
or U8434 (N_8434,N_8256,N_8322);
nor U8435 (N_8435,N_8392,N_8298);
nand U8436 (N_8436,N_8240,N_8286);
or U8437 (N_8437,N_8398,N_8254);
nand U8438 (N_8438,N_8266,N_8390);
nand U8439 (N_8439,N_8289,N_8316);
or U8440 (N_8440,N_8335,N_8200);
xnor U8441 (N_8441,N_8310,N_8210);
nor U8442 (N_8442,N_8385,N_8350);
xor U8443 (N_8443,N_8380,N_8209);
and U8444 (N_8444,N_8257,N_8279);
nor U8445 (N_8445,N_8329,N_8274);
nand U8446 (N_8446,N_8280,N_8312);
nor U8447 (N_8447,N_8261,N_8341);
or U8448 (N_8448,N_8395,N_8227);
xnor U8449 (N_8449,N_8248,N_8363);
xor U8450 (N_8450,N_8307,N_8263);
or U8451 (N_8451,N_8344,N_8214);
nand U8452 (N_8452,N_8340,N_8386);
or U8453 (N_8453,N_8206,N_8384);
nor U8454 (N_8454,N_8369,N_8302);
or U8455 (N_8455,N_8275,N_8376);
and U8456 (N_8456,N_8276,N_8281);
or U8457 (N_8457,N_8207,N_8374);
xor U8458 (N_8458,N_8391,N_8328);
or U8459 (N_8459,N_8283,N_8300);
nand U8460 (N_8460,N_8319,N_8353);
nand U8461 (N_8461,N_8333,N_8290);
xor U8462 (N_8462,N_8351,N_8228);
and U8463 (N_8463,N_8292,N_8225);
xor U8464 (N_8464,N_8301,N_8357);
nor U8465 (N_8465,N_8359,N_8267);
xor U8466 (N_8466,N_8347,N_8330);
or U8467 (N_8467,N_8381,N_8205);
nand U8468 (N_8468,N_8203,N_8318);
xnor U8469 (N_8469,N_8296,N_8241);
nand U8470 (N_8470,N_8324,N_8304);
and U8471 (N_8471,N_8217,N_8268);
or U8472 (N_8472,N_8251,N_8222);
xor U8473 (N_8473,N_8326,N_8365);
nand U8474 (N_8474,N_8325,N_8287);
or U8475 (N_8475,N_8343,N_8271);
or U8476 (N_8476,N_8352,N_8272);
nand U8477 (N_8477,N_8238,N_8378);
nand U8478 (N_8478,N_8224,N_8249);
nand U8479 (N_8479,N_8309,N_8305);
or U8480 (N_8480,N_8247,N_8278);
nor U8481 (N_8481,N_8255,N_8361);
nand U8482 (N_8482,N_8336,N_8269);
xor U8483 (N_8483,N_8246,N_8216);
nor U8484 (N_8484,N_8231,N_8218);
and U8485 (N_8485,N_8208,N_8285);
nor U8486 (N_8486,N_8368,N_8258);
and U8487 (N_8487,N_8314,N_8284);
or U8488 (N_8488,N_8244,N_8201);
xor U8489 (N_8489,N_8388,N_8346);
and U8490 (N_8490,N_8235,N_8291);
nand U8491 (N_8491,N_8345,N_8270);
nor U8492 (N_8492,N_8396,N_8299);
or U8493 (N_8493,N_8293,N_8215);
nor U8494 (N_8494,N_8367,N_8295);
nand U8495 (N_8495,N_8236,N_8237);
or U8496 (N_8496,N_8387,N_8223);
xnor U8497 (N_8497,N_8313,N_8252);
xor U8498 (N_8498,N_8264,N_8297);
nor U8499 (N_8499,N_8239,N_8250);
nand U8500 (N_8500,N_8248,N_8310);
and U8501 (N_8501,N_8236,N_8396);
nand U8502 (N_8502,N_8270,N_8243);
xor U8503 (N_8503,N_8229,N_8295);
nor U8504 (N_8504,N_8261,N_8258);
nand U8505 (N_8505,N_8234,N_8379);
xnor U8506 (N_8506,N_8268,N_8293);
nand U8507 (N_8507,N_8238,N_8335);
or U8508 (N_8508,N_8221,N_8378);
xor U8509 (N_8509,N_8234,N_8228);
xnor U8510 (N_8510,N_8287,N_8396);
nand U8511 (N_8511,N_8222,N_8263);
and U8512 (N_8512,N_8327,N_8225);
nor U8513 (N_8513,N_8392,N_8383);
and U8514 (N_8514,N_8388,N_8253);
xor U8515 (N_8515,N_8361,N_8221);
and U8516 (N_8516,N_8227,N_8284);
or U8517 (N_8517,N_8287,N_8394);
nand U8518 (N_8518,N_8325,N_8369);
nor U8519 (N_8519,N_8251,N_8333);
nor U8520 (N_8520,N_8347,N_8221);
nor U8521 (N_8521,N_8357,N_8298);
or U8522 (N_8522,N_8367,N_8360);
nand U8523 (N_8523,N_8299,N_8211);
nor U8524 (N_8524,N_8232,N_8223);
nand U8525 (N_8525,N_8354,N_8297);
nor U8526 (N_8526,N_8239,N_8289);
and U8527 (N_8527,N_8384,N_8217);
xor U8528 (N_8528,N_8362,N_8283);
and U8529 (N_8529,N_8365,N_8214);
nor U8530 (N_8530,N_8347,N_8271);
xnor U8531 (N_8531,N_8334,N_8389);
xor U8532 (N_8532,N_8288,N_8221);
xnor U8533 (N_8533,N_8329,N_8312);
nand U8534 (N_8534,N_8206,N_8389);
or U8535 (N_8535,N_8396,N_8342);
and U8536 (N_8536,N_8310,N_8257);
xor U8537 (N_8537,N_8227,N_8241);
nor U8538 (N_8538,N_8282,N_8356);
and U8539 (N_8539,N_8252,N_8202);
xor U8540 (N_8540,N_8255,N_8270);
xor U8541 (N_8541,N_8226,N_8344);
and U8542 (N_8542,N_8268,N_8338);
nor U8543 (N_8543,N_8281,N_8370);
and U8544 (N_8544,N_8217,N_8201);
and U8545 (N_8545,N_8279,N_8302);
nand U8546 (N_8546,N_8388,N_8267);
and U8547 (N_8547,N_8277,N_8234);
nand U8548 (N_8548,N_8224,N_8274);
xor U8549 (N_8549,N_8383,N_8319);
nor U8550 (N_8550,N_8385,N_8223);
and U8551 (N_8551,N_8305,N_8230);
nor U8552 (N_8552,N_8335,N_8225);
nor U8553 (N_8553,N_8281,N_8349);
and U8554 (N_8554,N_8240,N_8372);
xnor U8555 (N_8555,N_8205,N_8256);
nand U8556 (N_8556,N_8259,N_8368);
nor U8557 (N_8557,N_8373,N_8380);
xnor U8558 (N_8558,N_8328,N_8317);
nand U8559 (N_8559,N_8231,N_8201);
and U8560 (N_8560,N_8396,N_8341);
nand U8561 (N_8561,N_8252,N_8293);
nand U8562 (N_8562,N_8322,N_8376);
and U8563 (N_8563,N_8395,N_8397);
and U8564 (N_8564,N_8206,N_8326);
nand U8565 (N_8565,N_8356,N_8343);
nor U8566 (N_8566,N_8376,N_8285);
nor U8567 (N_8567,N_8323,N_8294);
or U8568 (N_8568,N_8231,N_8320);
xor U8569 (N_8569,N_8341,N_8297);
xor U8570 (N_8570,N_8338,N_8363);
nor U8571 (N_8571,N_8292,N_8231);
xor U8572 (N_8572,N_8248,N_8309);
nor U8573 (N_8573,N_8361,N_8384);
or U8574 (N_8574,N_8367,N_8395);
nand U8575 (N_8575,N_8394,N_8263);
nor U8576 (N_8576,N_8223,N_8337);
or U8577 (N_8577,N_8309,N_8205);
xor U8578 (N_8578,N_8257,N_8300);
nor U8579 (N_8579,N_8333,N_8266);
nor U8580 (N_8580,N_8370,N_8245);
or U8581 (N_8581,N_8354,N_8386);
and U8582 (N_8582,N_8263,N_8395);
or U8583 (N_8583,N_8221,N_8286);
or U8584 (N_8584,N_8295,N_8376);
xnor U8585 (N_8585,N_8346,N_8231);
and U8586 (N_8586,N_8203,N_8224);
xor U8587 (N_8587,N_8297,N_8249);
nand U8588 (N_8588,N_8323,N_8213);
or U8589 (N_8589,N_8383,N_8251);
xnor U8590 (N_8590,N_8298,N_8207);
xnor U8591 (N_8591,N_8296,N_8228);
xor U8592 (N_8592,N_8260,N_8302);
nor U8593 (N_8593,N_8375,N_8246);
and U8594 (N_8594,N_8213,N_8356);
or U8595 (N_8595,N_8234,N_8301);
nand U8596 (N_8596,N_8340,N_8325);
xor U8597 (N_8597,N_8373,N_8246);
xnor U8598 (N_8598,N_8259,N_8215);
nor U8599 (N_8599,N_8299,N_8290);
nand U8600 (N_8600,N_8528,N_8418);
xor U8601 (N_8601,N_8488,N_8499);
or U8602 (N_8602,N_8578,N_8535);
and U8603 (N_8603,N_8425,N_8401);
and U8604 (N_8604,N_8458,N_8447);
nor U8605 (N_8605,N_8482,N_8438);
or U8606 (N_8606,N_8465,N_8455);
nor U8607 (N_8607,N_8520,N_8506);
or U8608 (N_8608,N_8597,N_8584);
nor U8609 (N_8609,N_8534,N_8453);
nor U8610 (N_8610,N_8441,N_8531);
xnor U8611 (N_8611,N_8514,N_8537);
or U8612 (N_8612,N_8460,N_8496);
nand U8613 (N_8613,N_8513,N_8443);
nor U8614 (N_8614,N_8463,N_8477);
and U8615 (N_8615,N_8495,N_8414);
nand U8616 (N_8616,N_8544,N_8437);
xor U8617 (N_8617,N_8571,N_8554);
nor U8618 (N_8618,N_8574,N_8423);
or U8619 (N_8619,N_8536,N_8567);
nor U8620 (N_8620,N_8510,N_8481);
or U8621 (N_8621,N_8468,N_8442);
nand U8622 (N_8622,N_8586,N_8466);
nor U8623 (N_8623,N_8493,N_8553);
or U8624 (N_8624,N_8511,N_8433);
nand U8625 (N_8625,N_8491,N_8426);
nor U8626 (N_8626,N_8522,N_8518);
or U8627 (N_8627,N_8552,N_8568);
xnor U8628 (N_8628,N_8570,N_8408);
xnor U8629 (N_8629,N_8489,N_8421);
xor U8630 (N_8630,N_8596,N_8427);
and U8631 (N_8631,N_8525,N_8583);
or U8632 (N_8632,N_8530,N_8572);
nor U8633 (N_8633,N_8475,N_8588);
or U8634 (N_8634,N_8539,N_8573);
or U8635 (N_8635,N_8532,N_8478);
nand U8636 (N_8636,N_8565,N_8472);
or U8637 (N_8637,N_8557,N_8436);
nor U8638 (N_8638,N_8529,N_8402);
and U8639 (N_8639,N_8448,N_8400);
xor U8640 (N_8640,N_8521,N_8480);
and U8641 (N_8641,N_8487,N_8435);
and U8642 (N_8642,N_8439,N_8484);
xnor U8643 (N_8643,N_8424,N_8420);
nor U8644 (N_8644,N_8416,N_8541);
xnor U8645 (N_8645,N_8549,N_8562);
or U8646 (N_8646,N_8497,N_8474);
nand U8647 (N_8647,N_8490,N_8500);
nand U8648 (N_8648,N_8569,N_8575);
nor U8649 (N_8649,N_8551,N_8459);
and U8650 (N_8650,N_8403,N_8413);
or U8651 (N_8651,N_8446,N_8503);
nor U8652 (N_8652,N_8547,N_8450);
xnor U8653 (N_8653,N_8440,N_8467);
and U8654 (N_8654,N_8594,N_8599);
xnor U8655 (N_8655,N_8422,N_8409);
xor U8656 (N_8656,N_8563,N_8451);
or U8657 (N_8657,N_8498,N_8581);
or U8658 (N_8658,N_8429,N_8431);
or U8659 (N_8659,N_8464,N_8545);
nor U8660 (N_8660,N_8566,N_8558);
and U8661 (N_8661,N_8504,N_8579);
or U8662 (N_8662,N_8598,N_8419);
nor U8663 (N_8663,N_8515,N_8457);
nor U8664 (N_8664,N_8494,N_8434);
and U8665 (N_8665,N_8492,N_8417);
xor U8666 (N_8666,N_8509,N_8471);
and U8667 (N_8667,N_8592,N_8404);
xor U8668 (N_8668,N_8526,N_8516);
nand U8669 (N_8669,N_8512,N_8406);
and U8670 (N_8670,N_8508,N_8502);
nor U8671 (N_8671,N_8543,N_8428);
nand U8672 (N_8672,N_8542,N_8527);
nand U8673 (N_8673,N_8476,N_8410);
and U8674 (N_8674,N_8593,N_8462);
nor U8675 (N_8675,N_8561,N_8589);
and U8676 (N_8676,N_8449,N_8590);
nor U8677 (N_8677,N_8540,N_8585);
or U8678 (N_8678,N_8454,N_8412);
nor U8679 (N_8679,N_8483,N_8555);
or U8680 (N_8680,N_8444,N_8548);
xnor U8681 (N_8681,N_8445,N_8486);
and U8682 (N_8682,N_8538,N_8576);
nor U8683 (N_8683,N_8524,N_8411);
nor U8684 (N_8684,N_8577,N_8591);
nand U8685 (N_8685,N_8533,N_8517);
or U8686 (N_8686,N_8505,N_8479);
xor U8687 (N_8687,N_8519,N_8550);
or U8688 (N_8688,N_8582,N_8485);
and U8689 (N_8689,N_8415,N_8580);
nand U8690 (N_8690,N_8469,N_8432);
xor U8691 (N_8691,N_8523,N_8405);
and U8692 (N_8692,N_8564,N_8407);
and U8693 (N_8693,N_8470,N_8456);
nand U8694 (N_8694,N_8546,N_8452);
or U8695 (N_8695,N_8595,N_8507);
nand U8696 (N_8696,N_8560,N_8559);
nor U8697 (N_8697,N_8473,N_8430);
nand U8698 (N_8698,N_8587,N_8556);
or U8699 (N_8699,N_8461,N_8501);
xnor U8700 (N_8700,N_8577,N_8438);
and U8701 (N_8701,N_8567,N_8496);
xnor U8702 (N_8702,N_8592,N_8511);
and U8703 (N_8703,N_8571,N_8555);
or U8704 (N_8704,N_8563,N_8432);
and U8705 (N_8705,N_8569,N_8598);
nand U8706 (N_8706,N_8464,N_8419);
nor U8707 (N_8707,N_8484,N_8522);
nor U8708 (N_8708,N_8547,N_8466);
or U8709 (N_8709,N_8569,N_8538);
nor U8710 (N_8710,N_8411,N_8481);
nor U8711 (N_8711,N_8575,N_8592);
or U8712 (N_8712,N_8486,N_8586);
nor U8713 (N_8713,N_8495,N_8591);
and U8714 (N_8714,N_8584,N_8498);
nor U8715 (N_8715,N_8452,N_8489);
nor U8716 (N_8716,N_8590,N_8595);
xnor U8717 (N_8717,N_8565,N_8594);
or U8718 (N_8718,N_8489,N_8544);
nand U8719 (N_8719,N_8501,N_8439);
xnor U8720 (N_8720,N_8450,N_8528);
xor U8721 (N_8721,N_8407,N_8527);
and U8722 (N_8722,N_8408,N_8556);
nand U8723 (N_8723,N_8479,N_8546);
nand U8724 (N_8724,N_8506,N_8530);
or U8725 (N_8725,N_8581,N_8585);
nor U8726 (N_8726,N_8574,N_8490);
nand U8727 (N_8727,N_8581,N_8555);
nor U8728 (N_8728,N_8502,N_8459);
or U8729 (N_8729,N_8556,N_8433);
or U8730 (N_8730,N_8446,N_8468);
nand U8731 (N_8731,N_8457,N_8480);
and U8732 (N_8732,N_8566,N_8418);
nor U8733 (N_8733,N_8506,N_8449);
or U8734 (N_8734,N_8481,N_8577);
nor U8735 (N_8735,N_8472,N_8416);
xor U8736 (N_8736,N_8560,N_8586);
nor U8737 (N_8737,N_8555,N_8547);
and U8738 (N_8738,N_8401,N_8506);
or U8739 (N_8739,N_8584,N_8406);
and U8740 (N_8740,N_8472,N_8539);
xor U8741 (N_8741,N_8548,N_8586);
and U8742 (N_8742,N_8474,N_8463);
or U8743 (N_8743,N_8425,N_8408);
xnor U8744 (N_8744,N_8562,N_8494);
nand U8745 (N_8745,N_8579,N_8599);
or U8746 (N_8746,N_8506,N_8498);
and U8747 (N_8747,N_8502,N_8473);
xor U8748 (N_8748,N_8467,N_8569);
nor U8749 (N_8749,N_8404,N_8532);
or U8750 (N_8750,N_8560,N_8485);
nor U8751 (N_8751,N_8421,N_8486);
and U8752 (N_8752,N_8549,N_8469);
xnor U8753 (N_8753,N_8410,N_8589);
nand U8754 (N_8754,N_8491,N_8503);
xnor U8755 (N_8755,N_8506,N_8599);
xnor U8756 (N_8756,N_8540,N_8537);
nor U8757 (N_8757,N_8516,N_8521);
and U8758 (N_8758,N_8521,N_8451);
or U8759 (N_8759,N_8440,N_8575);
or U8760 (N_8760,N_8477,N_8565);
or U8761 (N_8761,N_8509,N_8598);
nand U8762 (N_8762,N_8486,N_8583);
nor U8763 (N_8763,N_8561,N_8494);
nand U8764 (N_8764,N_8573,N_8564);
and U8765 (N_8765,N_8593,N_8586);
nand U8766 (N_8766,N_8425,N_8522);
nand U8767 (N_8767,N_8485,N_8597);
xnor U8768 (N_8768,N_8505,N_8410);
nor U8769 (N_8769,N_8458,N_8555);
xor U8770 (N_8770,N_8460,N_8424);
and U8771 (N_8771,N_8576,N_8544);
or U8772 (N_8772,N_8498,N_8418);
nor U8773 (N_8773,N_8528,N_8535);
nor U8774 (N_8774,N_8417,N_8499);
nor U8775 (N_8775,N_8576,N_8426);
nand U8776 (N_8776,N_8492,N_8580);
xnor U8777 (N_8777,N_8439,N_8558);
nor U8778 (N_8778,N_8595,N_8562);
and U8779 (N_8779,N_8503,N_8598);
and U8780 (N_8780,N_8492,N_8463);
nor U8781 (N_8781,N_8551,N_8575);
and U8782 (N_8782,N_8537,N_8456);
nor U8783 (N_8783,N_8438,N_8465);
nor U8784 (N_8784,N_8486,N_8590);
xnor U8785 (N_8785,N_8516,N_8499);
nand U8786 (N_8786,N_8571,N_8499);
xnor U8787 (N_8787,N_8466,N_8460);
or U8788 (N_8788,N_8454,N_8578);
and U8789 (N_8789,N_8468,N_8560);
xnor U8790 (N_8790,N_8434,N_8485);
xnor U8791 (N_8791,N_8503,N_8531);
nand U8792 (N_8792,N_8444,N_8447);
or U8793 (N_8793,N_8483,N_8560);
nor U8794 (N_8794,N_8435,N_8400);
or U8795 (N_8795,N_8506,N_8544);
xor U8796 (N_8796,N_8566,N_8432);
and U8797 (N_8797,N_8476,N_8413);
xor U8798 (N_8798,N_8583,N_8418);
nor U8799 (N_8799,N_8421,N_8474);
nor U8800 (N_8800,N_8694,N_8615);
nand U8801 (N_8801,N_8720,N_8673);
or U8802 (N_8802,N_8701,N_8622);
nand U8803 (N_8803,N_8659,N_8786);
nor U8804 (N_8804,N_8736,N_8671);
or U8805 (N_8805,N_8698,N_8658);
nor U8806 (N_8806,N_8771,N_8756);
xnor U8807 (N_8807,N_8687,N_8683);
and U8808 (N_8808,N_8682,N_8775);
or U8809 (N_8809,N_8722,N_8649);
and U8810 (N_8810,N_8782,N_8778);
nor U8811 (N_8811,N_8734,N_8623);
nand U8812 (N_8812,N_8797,N_8679);
xnor U8813 (N_8813,N_8634,N_8670);
nand U8814 (N_8814,N_8616,N_8706);
nand U8815 (N_8815,N_8761,N_8688);
or U8816 (N_8816,N_8702,N_8703);
nand U8817 (N_8817,N_8638,N_8785);
nor U8818 (N_8818,N_8799,N_8677);
nor U8819 (N_8819,N_8727,N_8793);
and U8820 (N_8820,N_8691,N_8626);
and U8821 (N_8821,N_8686,N_8795);
nand U8822 (N_8822,N_8729,N_8610);
xnor U8823 (N_8823,N_8710,N_8781);
xnor U8824 (N_8824,N_8625,N_8768);
or U8825 (N_8825,N_8796,N_8743);
nand U8826 (N_8826,N_8642,N_8730);
or U8827 (N_8827,N_8618,N_8752);
nor U8828 (N_8828,N_8779,N_8725);
xor U8829 (N_8829,N_8663,N_8675);
xor U8830 (N_8830,N_8654,N_8708);
nor U8831 (N_8831,N_8717,N_8619);
nor U8832 (N_8832,N_8628,N_8646);
nand U8833 (N_8833,N_8762,N_8664);
or U8834 (N_8834,N_8630,N_8763);
and U8835 (N_8835,N_8769,N_8652);
or U8836 (N_8836,N_8693,N_8780);
xor U8837 (N_8837,N_8680,N_8755);
and U8838 (N_8838,N_8738,N_8731);
nand U8839 (N_8839,N_8635,N_8637);
nor U8840 (N_8840,N_8747,N_8739);
or U8841 (N_8841,N_8745,N_8772);
xor U8842 (N_8842,N_8653,N_8712);
or U8843 (N_8843,N_8620,N_8631);
xnor U8844 (N_8844,N_8651,N_8790);
and U8845 (N_8845,N_8629,N_8645);
nor U8846 (N_8846,N_8794,N_8666);
and U8847 (N_8847,N_8751,N_8723);
or U8848 (N_8848,N_8711,N_8692);
nor U8849 (N_8849,N_8647,N_8789);
and U8850 (N_8850,N_8719,N_8737);
or U8851 (N_8851,N_8784,N_8661);
nor U8852 (N_8852,N_8697,N_8648);
or U8853 (N_8853,N_8765,N_8740);
nand U8854 (N_8854,N_8650,N_8792);
nor U8855 (N_8855,N_8760,N_8684);
nor U8856 (N_8856,N_8709,N_8728);
or U8857 (N_8857,N_8716,N_8608);
and U8858 (N_8858,N_8639,N_8660);
nand U8859 (N_8859,N_8643,N_8668);
xor U8860 (N_8860,N_8685,N_8735);
nor U8861 (N_8861,N_8633,N_8700);
and U8862 (N_8862,N_8766,N_8721);
or U8863 (N_8863,N_8602,N_8605);
and U8864 (N_8864,N_8627,N_8678);
nand U8865 (N_8865,N_8732,N_8665);
and U8866 (N_8866,N_8770,N_8746);
nor U8867 (N_8867,N_8641,N_8798);
nor U8868 (N_8868,N_8669,N_8607);
or U8869 (N_8869,N_8742,N_8715);
or U8870 (N_8870,N_8611,N_8676);
nand U8871 (N_8871,N_8773,N_8764);
and U8872 (N_8872,N_8750,N_8690);
nand U8873 (N_8873,N_8724,N_8674);
nand U8874 (N_8874,N_8704,N_8655);
or U8875 (N_8875,N_8600,N_8718);
or U8876 (N_8876,N_8714,N_8656);
nor U8877 (N_8877,N_8681,N_8733);
or U8878 (N_8878,N_8689,N_8744);
nor U8879 (N_8879,N_8696,N_8753);
xnor U8880 (N_8880,N_8644,N_8614);
or U8881 (N_8881,N_8713,N_8672);
nand U8882 (N_8882,N_8632,N_8636);
xnor U8883 (N_8883,N_8707,N_8624);
nor U8884 (N_8884,N_8667,N_8787);
and U8885 (N_8885,N_8606,N_8695);
nand U8886 (N_8886,N_8604,N_8754);
and U8887 (N_8887,N_8776,N_8783);
or U8888 (N_8888,N_8777,N_8774);
xnor U8889 (N_8889,N_8640,N_8617);
and U8890 (N_8890,N_8741,N_8612);
nand U8891 (N_8891,N_8657,N_8699);
nor U8892 (N_8892,N_8621,N_8757);
or U8893 (N_8893,N_8613,N_8767);
xnor U8894 (N_8894,N_8791,N_8609);
and U8895 (N_8895,N_8603,N_8759);
and U8896 (N_8896,N_8662,N_8758);
nand U8897 (N_8897,N_8749,N_8705);
xor U8898 (N_8898,N_8788,N_8748);
nor U8899 (N_8899,N_8601,N_8726);
nor U8900 (N_8900,N_8791,N_8615);
xnor U8901 (N_8901,N_8750,N_8756);
xor U8902 (N_8902,N_8668,N_8670);
nor U8903 (N_8903,N_8784,N_8791);
nor U8904 (N_8904,N_8730,N_8766);
and U8905 (N_8905,N_8720,N_8696);
xnor U8906 (N_8906,N_8678,N_8700);
nor U8907 (N_8907,N_8616,N_8746);
nand U8908 (N_8908,N_8748,N_8694);
nor U8909 (N_8909,N_8697,N_8610);
and U8910 (N_8910,N_8611,N_8743);
or U8911 (N_8911,N_8606,N_8603);
and U8912 (N_8912,N_8745,N_8716);
and U8913 (N_8913,N_8659,N_8616);
xor U8914 (N_8914,N_8603,N_8746);
or U8915 (N_8915,N_8754,N_8673);
nand U8916 (N_8916,N_8723,N_8703);
and U8917 (N_8917,N_8638,N_8782);
nor U8918 (N_8918,N_8662,N_8615);
nor U8919 (N_8919,N_8678,N_8669);
nor U8920 (N_8920,N_8724,N_8763);
xor U8921 (N_8921,N_8704,N_8612);
nor U8922 (N_8922,N_8682,N_8727);
nor U8923 (N_8923,N_8679,N_8795);
or U8924 (N_8924,N_8625,N_8715);
nand U8925 (N_8925,N_8799,N_8601);
nand U8926 (N_8926,N_8702,N_8775);
nor U8927 (N_8927,N_8743,N_8643);
xor U8928 (N_8928,N_8734,N_8783);
nand U8929 (N_8929,N_8705,N_8776);
xnor U8930 (N_8930,N_8730,N_8667);
or U8931 (N_8931,N_8666,N_8604);
xnor U8932 (N_8932,N_8653,N_8664);
and U8933 (N_8933,N_8786,N_8799);
and U8934 (N_8934,N_8648,N_8763);
and U8935 (N_8935,N_8721,N_8765);
nand U8936 (N_8936,N_8608,N_8710);
nor U8937 (N_8937,N_8641,N_8757);
or U8938 (N_8938,N_8706,N_8665);
or U8939 (N_8939,N_8751,N_8620);
xnor U8940 (N_8940,N_8628,N_8796);
nor U8941 (N_8941,N_8633,N_8755);
nor U8942 (N_8942,N_8789,N_8772);
xor U8943 (N_8943,N_8695,N_8649);
nand U8944 (N_8944,N_8684,N_8776);
nor U8945 (N_8945,N_8680,N_8690);
xor U8946 (N_8946,N_8738,N_8641);
and U8947 (N_8947,N_8681,N_8621);
nor U8948 (N_8948,N_8750,N_8681);
xnor U8949 (N_8949,N_8738,N_8670);
nand U8950 (N_8950,N_8698,N_8669);
nor U8951 (N_8951,N_8619,N_8625);
xnor U8952 (N_8952,N_8748,N_8729);
nor U8953 (N_8953,N_8750,N_8687);
xnor U8954 (N_8954,N_8686,N_8646);
or U8955 (N_8955,N_8655,N_8690);
or U8956 (N_8956,N_8640,N_8616);
nor U8957 (N_8957,N_8695,N_8774);
xnor U8958 (N_8958,N_8657,N_8765);
nor U8959 (N_8959,N_8708,N_8748);
xor U8960 (N_8960,N_8672,N_8649);
and U8961 (N_8961,N_8713,N_8761);
and U8962 (N_8962,N_8716,N_8770);
and U8963 (N_8963,N_8672,N_8780);
xor U8964 (N_8964,N_8697,N_8618);
and U8965 (N_8965,N_8630,N_8679);
and U8966 (N_8966,N_8796,N_8757);
nor U8967 (N_8967,N_8773,N_8742);
or U8968 (N_8968,N_8665,N_8707);
xor U8969 (N_8969,N_8647,N_8646);
nand U8970 (N_8970,N_8688,N_8617);
nor U8971 (N_8971,N_8780,N_8729);
or U8972 (N_8972,N_8702,N_8701);
and U8973 (N_8973,N_8615,N_8669);
and U8974 (N_8974,N_8741,N_8676);
and U8975 (N_8975,N_8644,N_8792);
or U8976 (N_8976,N_8676,N_8672);
xnor U8977 (N_8977,N_8650,N_8689);
xor U8978 (N_8978,N_8702,N_8708);
nand U8979 (N_8979,N_8713,N_8773);
or U8980 (N_8980,N_8793,N_8775);
and U8981 (N_8981,N_8623,N_8646);
nand U8982 (N_8982,N_8687,N_8629);
nor U8983 (N_8983,N_8710,N_8639);
nor U8984 (N_8984,N_8715,N_8707);
and U8985 (N_8985,N_8654,N_8661);
xor U8986 (N_8986,N_8746,N_8776);
and U8987 (N_8987,N_8683,N_8606);
or U8988 (N_8988,N_8766,N_8752);
nand U8989 (N_8989,N_8794,N_8608);
and U8990 (N_8990,N_8738,N_8780);
nand U8991 (N_8991,N_8773,N_8651);
and U8992 (N_8992,N_8633,N_8754);
nand U8993 (N_8993,N_8791,N_8638);
nor U8994 (N_8994,N_8621,N_8703);
nor U8995 (N_8995,N_8602,N_8600);
and U8996 (N_8996,N_8751,N_8750);
nor U8997 (N_8997,N_8741,N_8644);
nor U8998 (N_8998,N_8740,N_8745);
or U8999 (N_8999,N_8709,N_8784);
nor U9000 (N_9000,N_8985,N_8887);
nor U9001 (N_9001,N_8841,N_8810);
nor U9002 (N_9002,N_8988,N_8839);
nor U9003 (N_9003,N_8967,N_8901);
nor U9004 (N_9004,N_8924,N_8999);
xor U9005 (N_9005,N_8979,N_8838);
or U9006 (N_9006,N_8906,N_8806);
and U9007 (N_9007,N_8889,N_8963);
or U9008 (N_9008,N_8960,N_8868);
and U9009 (N_9009,N_8909,N_8933);
nand U9010 (N_9010,N_8923,N_8872);
xor U9011 (N_9011,N_8832,N_8824);
nand U9012 (N_9012,N_8875,N_8890);
nor U9013 (N_9013,N_8958,N_8986);
xor U9014 (N_9014,N_8990,N_8918);
nand U9015 (N_9015,N_8934,N_8917);
nor U9016 (N_9016,N_8829,N_8910);
and U9017 (N_9017,N_8926,N_8807);
nor U9018 (N_9018,N_8930,N_8809);
nand U9019 (N_9019,N_8850,N_8965);
nand U9020 (N_9020,N_8995,N_8982);
xnor U9021 (N_9021,N_8880,N_8959);
nand U9022 (N_9022,N_8849,N_8856);
and U9023 (N_9023,N_8828,N_8882);
or U9024 (N_9024,N_8870,N_8914);
nand U9025 (N_9025,N_8896,N_8976);
xor U9026 (N_9026,N_8840,N_8885);
nor U9027 (N_9027,N_8892,N_8980);
xor U9028 (N_9028,N_8966,N_8867);
and U9029 (N_9029,N_8862,N_8821);
and U9030 (N_9030,N_8983,N_8811);
and U9031 (N_9031,N_8836,N_8851);
and U9032 (N_9032,N_8864,N_8897);
nor U9033 (N_9033,N_8931,N_8935);
xnor U9034 (N_9034,N_8820,N_8928);
nand U9035 (N_9035,N_8808,N_8816);
or U9036 (N_9036,N_8804,N_8920);
and U9037 (N_9037,N_8945,N_8873);
nand U9038 (N_9038,N_8978,N_8805);
nor U9039 (N_9039,N_8812,N_8912);
and U9040 (N_9040,N_8908,N_8992);
and U9041 (N_9041,N_8888,N_8863);
nand U9042 (N_9042,N_8940,N_8859);
nor U9043 (N_9043,N_8852,N_8943);
and U9044 (N_9044,N_8941,N_8922);
nand U9045 (N_9045,N_8830,N_8837);
or U9046 (N_9046,N_8884,N_8953);
nor U9047 (N_9047,N_8989,N_8815);
and U9048 (N_9048,N_8952,N_8956);
and U9049 (N_9049,N_8822,N_8916);
and U9050 (N_9050,N_8871,N_8913);
or U9051 (N_9051,N_8942,N_8893);
nand U9052 (N_9052,N_8899,N_8843);
or U9053 (N_9053,N_8987,N_8919);
nand U9054 (N_9054,N_8938,N_8950);
nand U9055 (N_9055,N_8968,N_8904);
xnor U9056 (N_9056,N_8925,N_8939);
and U9057 (N_9057,N_8819,N_8845);
nor U9058 (N_9058,N_8984,N_8858);
xnor U9059 (N_9059,N_8846,N_8835);
or U9060 (N_9060,N_8854,N_8895);
nor U9061 (N_9061,N_8996,N_8844);
and U9062 (N_9062,N_8977,N_8962);
xor U9063 (N_9063,N_8801,N_8818);
nand U9064 (N_9064,N_8961,N_8827);
xor U9065 (N_9065,N_8833,N_8877);
xor U9066 (N_9066,N_8951,N_8997);
or U9067 (N_9067,N_8921,N_8937);
and U9068 (N_9068,N_8927,N_8876);
or U9069 (N_9069,N_8879,N_8936);
and U9070 (N_9070,N_8869,N_8878);
and U9071 (N_9071,N_8883,N_8803);
nand U9072 (N_9072,N_8954,N_8813);
xnor U9073 (N_9073,N_8861,N_8911);
nor U9074 (N_9074,N_8975,N_8855);
nor U9075 (N_9075,N_8907,N_8847);
xnor U9076 (N_9076,N_8971,N_8857);
nor U9077 (N_9077,N_8974,N_8949);
and U9078 (N_9078,N_8957,N_8881);
xor U9079 (N_9079,N_8955,N_8970);
nand U9080 (N_9080,N_8826,N_8973);
nand U9081 (N_9081,N_8831,N_8866);
nor U9082 (N_9082,N_8814,N_8817);
nand U9083 (N_9083,N_8946,N_8894);
nand U9084 (N_9084,N_8964,N_8860);
nor U9085 (N_9085,N_8834,N_8991);
xor U9086 (N_9086,N_8825,N_8891);
or U9087 (N_9087,N_8993,N_8929);
xnor U9088 (N_9088,N_8981,N_8853);
and U9089 (N_9089,N_8994,N_8948);
nand U9090 (N_9090,N_8898,N_8902);
nor U9091 (N_9091,N_8842,N_8947);
or U9092 (N_9092,N_8932,N_8865);
and U9093 (N_9093,N_8903,N_8944);
nor U9094 (N_9094,N_8874,N_8800);
xor U9095 (N_9095,N_8972,N_8886);
or U9096 (N_9096,N_8848,N_8998);
nand U9097 (N_9097,N_8900,N_8915);
nand U9098 (N_9098,N_8802,N_8969);
and U9099 (N_9099,N_8905,N_8823);
nand U9100 (N_9100,N_8953,N_8892);
or U9101 (N_9101,N_8891,N_8878);
nor U9102 (N_9102,N_8939,N_8952);
nand U9103 (N_9103,N_8943,N_8840);
nor U9104 (N_9104,N_8961,N_8971);
xor U9105 (N_9105,N_8875,N_8831);
xnor U9106 (N_9106,N_8826,N_8904);
or U9107 (N_9107,N_8976,N_8977);
and U9108 (N_9108,N_8903,N_8986);
and U9109 (N_9109,N_8894,N_8841);
nand U9110 (N_9110,N_8841,N_8825);
nand U9111 (N_9111,N_8902,N_8852);
xnor U9112 (N_9112,N_8894,N_8881);
nor U9113 (N_9113,N_8952,N_8876);
nand U9114 (N_9114,N_8928,N_8890);
xor U9115 (N_9115,N_8929,N_8856);
and U9116 (N_9116,N_8921,N_8840);
nor U9117 (N_9117,N_8829,N_8964);
nand U9118 (N_9118,N_8826,N_8832);
xnor U9119 (N_9119,N_8895,N_8996);
and U9120 (N_9120,N_8886,N_8942);
and U9121 (N_9121,N_8947,N_8893);
and U9122 (N_9122,N_8838,N_8963);
xor U9123 (N_9123,N_8940,N_8861);
nor U9124 (N_9124,N_8967,N_8915);
nand U9125 (N_9125,N_8835,N_8843);
or U9126 (N_9126,N_8810,N_8809);
nand U9127 (N_9127,N_8800,N_8864);
nor U9128 (N_9128,N_8917,N_8979);
nor U9129 (N_9129,N_8831,N_8995);
xnor U9130 (N_9130,N_8935,N_8925);
nand U9131 (N_9131,N_8913,N_8847);
nor U9132 (N_9132,N_8992,N_8978);
or U9133 (N_9133,N_8814,N_8956);
nand U9134 (N_9134,N_8987,N_8850);
and U9135 (N_9135,N_8860,N_8946);
nor U9136 (N_9136,N_8991,N_8907);
or U9137 (N_9137,N_8925,N_8877);
and U9138 (N_9138,N_8931,N_8819);
and U9139 (N_9139,N_8989,N_8810);
or U9140 (N_9140,N_8944,N_8858);
xnor U9141 (N_9141,N_8855,N_8955);
and U9142 (N_9142,N_8899,N_8906);
and U9143 (N_9143,N_8929,N_8813);
nand U9144 (N_9144,N_8859,N_8974);
nor U9145 (N_9145,N_8947,N_8939);
nor U9146 (N_9146,N_8971,N_8953);
nand U9147 (N_9147,N_8876,N_8892);
and U9148 (N_9148,N_8845,N_8803);
nor U9149 (N_9149,N_8857,N_8898);
and U9150 (N_9150,N_8910,N_8947);
nand U9151 (N_9151,N_8835,N_8985);
nand U9152 (N_9152,N_8826,N_8962);
or U9153 (N_9153,N_8800,N_8901);
xor U9154 (N_9154,N_8907,N_8901);
xor U9155 (N_9155,N_8950,N_8940);
nor U9156 (N_9156,N_8870,N_8939);
or U9157 (N_9157,N_8842,N_8968);
or U9158 (N_9158,N_8810,N_8896);
or U9159 (N_9159,N_8937,N_8952);
and U9160 (N_9160,N_8920,N_8965);
nand U9161 (N_9161,N_8893,N_8987);
nor U9162 (N_9162,N_8807,N_8850);
xor U9163 (N_9163,N_8814,N_8886);
or U9164 (N_9164,N_8802,N_8870);
or U9165 (N_9165,N_8950,N_8936);
or U9166 (N_9166,N_8893,N_8925);
and U9167 (N_9167,N_8954,N_8917);
nor U9168 (N_9168,N_8949,N_8925);
and U9169 (N_9169,N_8987,N_8870);
and U9170 (N_9170,N_8970,N_8817);
xor U9171 (N_9171,N_8820,N_8864);
or U9172 (N_9172,N_8909,N_8946);
xor U9173 (N_9173,N_8990,N_8992);
or U9174 (N_9174,N_8946,N_8886);
and U9175 (N_9175,N_8955,N_8895);
nor U9176 (N_9176,N_8997,N_8801);
and U9177 (N_9177,N_8955,N_8917);
or U9178 (N_9178,N_8972,N_8914);
xor U9179 (N_9179,N_8966,N_8833);
and U9180 (N_9180,N_8816,N_8888);
nand U9181 (N_9181,N_8931,N_8845);
xor U9182 (N_9182,N_8829,N_8859);
and U9183 (N_9183,N_8971,N_8842);
nor U9184 (N_9184,N_8834,N_8952);
and U9185 (N_9185,N_8960,N_8969);
and U9186 (N_9186,N_8956,N_8804);
xor U9187 (N_9187,N_8964,N_8891);
nor U9188 (N_9188,N_8861,N_8883);
nand U9189 (N_9189,N_8823,N_8952);
xor U9190 (N_9190,N_8923,N_8880);
nand U9191 (N_9191,N_8951,N_8864);
xor U9192 (N_9192,N_8818,N_8823);
nand U9193 (N_9193,N_8867,N_8826);
xnor U9194 (N_9194,N_8916,N_8950);
nand U9195 (N_9195,N_8885,N_8989);
nor U9196 (N_9196,N_8916,N_8921);
nor U9197 (N_9197,N_8869,N_8838);
xnor U9198 (N_9198,N_8926,N_8975);
or U9199 (N_9199,N_8947,N_8997);
or U9200 (N_9200,N_9154,N_9073);
or U9201 (N_9201,N_9165,N_9130);
nand U9202 (N_9202,N_9182,N_9134);
nand U9203 (N_9203,N_9009,N_9033);
or U9204 (N_9204,N_9172,N_9138);
xnor U9205 (N_9205,N_9026,N_9099);
nand U9206 (N_9206,N_9075,N_9044);
xor U9207 (N_9207,N_9055,N_9108);
xnor U9208 (N_9208,N_9120,N_9091);
and U9209 (N_9209,N_9006,N_9093);
nand U9210 (N_9210,N_9052,N_9066);
xnor U9211 (N_9211,N_9089,N_9077);
nor U9212 (N_9212,N_9084,N_9079);
nor U9213 (N_9213,N_9169,N_9005);
and U9214 (N_9214,N_9048,N_9156);
xor U9215 (N_9215,N_9114,N_9060);
and U9216 (N_9216,N_9147,N_9041);
and U9217 (N_9217,N_9106,N_9150);
nand U9218 (N_9218,N_9000,N_9162);
nor U9219 (N_9219,N_9187,N_9196);
and U9220 (N_9220,N_9125,N_9057);
nor U9221 (N_9221,N_9034,N_9110);
xor U9222 (N_9222,N_9019,N_9148);
and U9223 (N_9223,N_9047,N_9132);
or U9224 (N_9224,N_9159,N_9070);
nor U9225 (N_9225,N_9139,N_9039);
nand U9226 (N_9226,N_9163,N_9180);
and U9227 (N_9227,N_9010,N_9038);
and U9228 (N_9228,N_9144,N_9197);
nor U9229 (N_9229,N_9017,N_9140);
xnor U9230 (N_9230,N_9141,N_9068);
nor U9231 (N_9231,N_9015,N_9049);
and U9232 (N_9232,N_9043,N_9118);
and U9233 (N_9233,N_9104,N_9067);
xnor U9234 (N_9234,N_9097,N_9087);
xnor U9235 (N_9235,N_9136,N_9167);
xnor U9236 (N_9236,N_9014,N_9123);
or U9237 (N_9237,N_9124,N_9025);
xor U9238 (N_9238,N_9058,N_9088);
nand U9239 (N_9239,N_9086,N_9184);
nand U9240 (N_9240,N_9186,N_9090);
and U9241 (N_9241,N_9064,N_9032);
and U9242 (N_9242,N_9135,N_9107);
and U9243 (N_9243,N_9189,N_9050);
and U9244 (N_9244,N_9011,N_9193);
or U9245 (N_9245,N_9171,N_9027);
xor U9246 (N_9246,N_9013,N_9179);
and U9247 (N_9247,N_9028,N_9096);
and U9248 (N_9248,N_9071,N_9054);
and U9249 (N_9249,N_9022,N_9115);
xnor U9250 (N_9250,N_9183,N_9149);
nand U9251 (N_9251,N_9185,N_9080);
xnor U9252 (N_9252,N_9194,N_9101);
or U9253 (N_9253,N_9188,N_9031);
or U9254 (N_9254,N_9024,N_9155);
and U9255 (N_9255,N_9190,N_9012);
and U9256 (N_9256,N_9176,N_9004);
nor U9257 (N_9257,N_9046,N_9145);
or U9258 (N_9258,N_9094,N_9195);
xnor U9259 (N_9259,N_9131,N_9152);
nor U9260 (N_9260,N_9113,N_9092);
or U9261 (N_9261,N_9018,N_9042);
nor U9262 (N_9262,N_9158,N_9174);
nand U9263 (N_9263,N_9157,N_9095);
nand U9264 (N_9264,N_9061,N_9081);
nand U9265 (N_9265,N_9128,N_9051);
and U9266 (N_9266,N_9122,N_9102);
or U9267 (N_9267,N_9007,N_9030);
and U9268 (N_9268,N_9117,N_9127);
xor U9269 (N_9269,N_9173,N_9069);
and U9270 (N_9270,N_9137,N_9199);
and U9271 (N_9271,N_9008,N_9072);
and U9272 (N_9272,N_9062,N_9164);
xor U9273 (N_9273,N_9181,N_9074);
nand U9274 (N_9274,N_9035,N_9161);
and U9275 (N_9275,N_9037,N_9001);
nor U9276 (N_9276,N_9021,N_9020);
xor U9277 (N_9277,N_9059,N_9191);
nor U9278 (N_9278,N_9003,N_9111);
or U9279 (N_9279,N_9029,N_9168);
nor U9280 (N_9280,N_9129,N_9198);
nand U9281 (N_9281,N_9177,N_9166);
or U9282 (N_9282,N_9100,N_9119);
or U9283 (N_9283,N_9170,N_9023);
and U9284 (N_9284,N_9103,N_9056);
and U9285 (N_9285,N_9133,N_9040);
nor U9286 (N_9286,N_9082,N_9002);
and U9287 (N_9287,N_9146,N_9078);
and U9288 (N_9288,N_9085,N_9016);
xor U9289 (N_9289,N_9076,N_9116);
nor U9290 (N_9290,N_9126,N_9045);
nor U9291 (N_9291,N_9192,N_9143);
and U9292 (N_9292,N_9083,N_9121);
xor U9293 (N_9293,N_9109,N_9063);
and U9294 (N_9294,N_9053,N_9142);
or U9295 (N_9295,N_9151,N_9098);
and U9296 (N_9296,N_9175,N_9065);
nor U9297 (N_9297,N_9112,N_9178);
nand U9298 (N_9298,N_9105,N_9153);
xor U9299 (N_9299,N_9160,N_9036);
nor U9300 (N_9300,N_9071,N_9093);
and U9301 (N_9301,N_9096,N_9080);
or U9302 (N_9302,N_9036,N_9116);
or U9303 (N_9303,N_9077,N_9154);
nor U9304 (N_9304,N_9186,N_9089);
nor U9305 (N_9305,N_9089,N_9125);
xor U9306 (N_9306,N_9103,N_9198);
xor U9307 (N_9307,N_9021,N_9061);
xnor U9308 (N_9308,N_9041,N_9054);
xnor U9309 (N_9309,N_9139,N_9011);
xor U9310 (N_9310,N_9052,N_9139);
or U9311 (N_9311,N_9140,N_9053);
nand U9312 (N_9312,N_9105,N_9142);
xor U9313 (N_9313,N_9184,N_9059);
or U9314 (N_9314,N_9097,N_9049);
and U9315 (N_9315,N_9038,N_9144);
nor U9316 (N_9316,N_9066,N_9126);
nand U9317 (N_9317,N_9105,N_9081);
or U9318 (N_9318,N_9118,N_9079);
nand U9319 (N_9319,N_9151,N_9101);
nor U9320 (N_9320,N_9099,N_9167);
or U9321 (N_9321,N_9080,N_9000);
or U9322 (N_9322,N_9037,N_9150);
nand U9323 (N_9323,N_9045,N_9129);
nand U9324 (N_9324,N_9042,N_9079);
nor U9325 (N_9325,N_9081,N_9037);
nand U9326 (N_9326,N_9185,N_9038);
xor U9327 (N_9327,N_9010,N_9026);
xor U9328 (N_9328,N_9036,N_9042);
and U9329 (N_9329,N_9071,N_9187);
nor U9330 (N_9330,N_9176,N_9141);
or U9331 (N_9331,N_9054,N_9040);
and U9332 (N_9332,N_9030,N_9153);
nor U9333 (N_9333,N_9038,N_9177);
nor U9334 (N_9334,N_9154,N_9132);
nand U9335 (N_9335,N_9188,N_9126);
or U9336 (N_9336,N_9100,N_9143);
nor U9337 (N_9337,N_9028,N_9180);
nor U9338 (N_9338,N_9138,N_9143);
or U9339 (N_9339,N_9149,N_9031);
and U9340 (N_9340,N_9178,N_9034);
or U9341 (N_9341,N_9139,N_9111);
and U9342 (N_9342,N_9101,N_9133);
xnor U9343 (N_9343,N_9089,N_9002);
or U9344 (N_9344,N_9022,N_9101);
nor U9345 (N_9345,N_9160,N_9109);
nand U9346 (N_9346,N_9181,N_9020);
or U9347 (N_9347,N_9027,N_9013);
xor U9348 (N_9348,N_9064,N_9192);
xnor U9349 (N_9349,N_9161,N_9151);
nand U9350 (N_9350,N_9083,N_9149);
and U9351 (N_9351,N_9110,N_9160);
nand U9352 (N_9352,N_9118,N_9084);
or U9353 (N_9353,N_9019,N_9177);
xnor U9354 (N_9354,N_9163,N_9198);
and U9355 (N_9355,N_9025,N_9162);
xnor U9356 (N_9356,N_9176,N_9168);
nand U9357 (N_9357,N_9019,N_9195);
nor U9358 (N_9358,N_9054,N_9051);
nor U9359 (N_9359,N_9169,N_9137);
nor U9360 (N_9360,N_9034,N_9108);
or U9361 (N_9361,N_9034,N_9039);
nor U9362 (N_9362,N_9001,N_9023);
or U9363 (N_9363,N_9184,N_9065);
xnor U9364 (N_9364,N_9079,N_9134);
xnor U9365 (N_9365,N_9011,N_9053);
nand U9366 (N_9366,N_9064,N_9198);
xnor U9367 (N_9367,N_9145,N_9095);
xnor U9368 (N_9368,N_9075,N_9176);
and U9369 (N_9369,N_9069,N_9018);
and U9370 (N_9370,N_9191,N_9136);
nor U9371 (N_9371,N_9095,N_9057);
and U9372 (N_9372,N_9035,N_9114);
nor U9373 (N_9373,N_9133,N_9038);
and U9374 (N_9374,N_9150,N_9071);
nor U9375 (N_9375,N_9058,N_9062);
xnor U9376 (N_9376,N_9013,N_9084);
and U9377 (N_9377,N_9071,N_9091);
xor U9378 (N_9378,N_9108,N_9046);
nand U9379 (N_9379,N_9138,N_9025);
and U9380 (N_9380,N_9039,N_9178);
or U9381 (N_9381,N_9162,N_9182);
nor U9382 (N_9382,N_9066,N_9057);
or U9383 (N_9383,N_9040,N_9192);
or U9384 (N_9384,N_9128,N_9137);
or U9385 (N_9385,N_9145,N_9125);
xor U9386 (N_9386,N_9147,N_9189);
or U9387 (N_9387,N_9151,N_9033);
or U9388 (N_9388,N_9188,N_9067);
and U9389 (N_9389,N_9013,N_9021);
or U9390 (N_9390,N_9068,N_9197);
and U9391 (N_9391,N_9171,N_9161);
and U9392 (N_9392,N_9172,N_9001);
and U9393 (N_9393,N_9003,N_9167);
nor U9394 (N_9394,N_9057,N_9111);
nor U9395 (N_9395,N_9178,N_9118);
or U9396 (N_9396,N_9114,N_9126);
nor U9397 (N_9397,N_9137,N_9000);
nand U9398 (N_9398,N_9151,N_9140);
or U9399 (N_9399,N_9178,N_9144);
and U9400 (N_9400,N_9274,N_9288);
nor U9401 (N_9401,N_9250,N_9323);
and U9402 (N_9402,N_9310,N_9233);
and U9403 (N_9403,N_9253,N_9211);
and U9404 (N_9404,N_9258,N_9383);
or U9405 (N_9405,N_9388,N_9257);
xor U9406 (N_9406,N_9237,N_9393);
nor U9407 (N_9407,N_9295,N_9366);
nor U9408 (N_9408,N_9372,N_9395);
or U9409 (N_9409,N_9337,N_9209);
and U9410 (N_9410,N_9389,N_9362);
or U9411 (N_9411,N_9227,N_9304);
xor U9412 (N_9412,N_9268,N_9208);
and U9413 (N_9413,N_9203,N_9215);
or U9414 (N_9414,N_9297,N_9207);
and U9415 (N_9415,N_9391,N_9213);
nand U9416 (N_9416,N_9262,N_9272);
nand U9417 (N_9417,N_9394,N_9280);
nand U9418 (N_9418,N_9277,N_9273);
xor U9419 (N_9419,N_9222,N_9200);
nand U9420 (N_9420,N_9303,N_9336);
nor U9421 (N_9421,N_9333,N_9229);
nor U9422 (N_9422,N_9326,N_9344);
nand U9423 (N_9423,N_9263,N_9279);
nor U9424 (N_9424,N_9380,N_9248);
xor U9425 (N_9425,N_9236,N_9278);
or U9426 (N_9426,N_9351,N_9354);
nand U9427 (N_9427,N_9330,N_9361);
or U9428 (N_9428,N_9242,N_9316);
nor U9429 (N_9429,N_9212,N_9398);
nand U9430 (N_9430,N_9382,N_9217);
and U9431 (N_9431,N_9219,N_9264);
xnor U9432 (N_9432,N_9235,N_9343);
and U9433 (N_9433,N_9376,N_9218);
nor U9434 (N_9434,N_9340,N_9284);
and U9435 (N_9435,N_9232,N_9285);
nor U9436 (N_9436,N_9271,N_9359);
xor U9437 (N_9437,N_9311,N_9346);
and U9438 (N_9438,N_9320,N_9313);
and U9439 (N_9439,N_9319,N_9345);
nor U9440 (N_9440,N_9228,N_9234);
xor U9441 (N_9441,N_9378,N_9334);
xnor U9442 (N_9442,N_9292,N_9287);
and U9443 (N_9443,N_9358,N_9363);
nand U9444 (N_9444,N_9241,N_9387);
xnor U9445 (N_9445,N_9305,N_9275);
nand U9446 (N_9446,N_9399,N_9254);
nor U9447 (N_9447,N_9259,N_9375);
or U9448 (N_9448,N_9360,N_9296);
nor U9449 (N_9449,N_9281,N_9314);
and U9450 (N_9450,N_9243,N_9249);
or U9451 (N_9451,N_9283,N_9377);
or U9452 (N_9452,N_9353,N_9201);
nand U9453 (N_9453,N_9214,N_9202);
xor U9454 (N_9454,N_9379,N_9269);
nand U9455 (N_9455,N_9260,N_9276);
or U9456 (N_9456,N_9369,N_9325);
nand U9457 (N_9457,N_9289,N_9392);
or U9458 (N_9458,N_9230,N_9307);
xnor U9459 (N_9459,N_9328,N_9396);
nand U9460 (N_9460,N_9204,N_9327);
or U9461 (N_9461,N_9347,N_9338);
xnor U9462 (N_9462,N_9322,N_9348);
xor U9463 (N_9463,N_9384,N_9373);
and U9464 (N_9464,N_9371,N_9205);
nand U9465 (N_9465,N_9298,N_9370);
and U9466 (N_9466,N_9365,N_9231);
nand U9467 (N_9467,N_9390,N_9270);
xnor U9468 (N_9468,N_9357,N_9252);
and U9469 (N_9469,N_9266,N_9282);
xnor U9470 (N_9470,N_9240,N_9397);
and U9471 (N_9471,N_9341,N_9317);
and U9472 (N_9472,N_9300,N_9315);
xnor U9473 (N_9473,N_9256,N_9342);
xnor U9474 (N_9474,N_9339,N_9245);
and U9475 (N_9475,N_9301,N_9220);
xnor U9476 (N_9476,N_9381,N_9309);
nor U9477 (N_9477,N_9244,N_9291);
xor U9478 (N_9478,N_9216,N_9294);
or U9479 (N_9479,N_9368,N_9299);
nand U9480 (N_9480,N_9265,N_9221);
nor U9481 (N_9481,N_9386,N_9318);
nand U9482 (N_9482,N_9210,N_9261);
xor U9483 (N_9483,N_9251,N_9356);
and U9484 (N_9484,N_9329,N_9239);
or U9485 (N_9485,N_9324,N_9331);
nor U9486 (N_9486,N_9247,N_9352);
nor U9487 (N_9487,N_9374,N_9238);
and U9488 (N_9488,N_9302,N_9286);
and U9489 (N_9489,N_9355,N_9364);
and U9490 (N_9490,N_9226,N_9246);
or U9491 (N_9491,N_9290,N_9335);
nand U9492 (N_9492,N_9223,N_9332);
and U9493 (N_9493,N_9206,N_9306);
nand U9494 (N_9494,N_9293,N_9349);
or U9495 (N_9495,N_9308,N_9385);
or U9496 (N_9496,N_9224,N_9321);
nor U9497 (N_9497,N_9367,N_9312);
nand U9498 (N_9498,N_9350,N_9267);
or U9499 (N_9499,N_9255,N_9225);
nor U9500 (N_9500,N_9239,N_9343);
nand U9501 (N_9501,N_9260,N_9364);
nand U9502 (N_9502,N_9235,N_9267);
and U9503 (N_9503,N_9294,N_9234);
xor U9504 (N_9504,N_9347,N_9222);
nand U9505 (N_9505,N_9204,N_9328);
nand U9506 (N_9506,N_9223,N_9306);
xor U9507 (N_9507,N_9227,N_9317);
xor U9508 (N_9508,N_9337,N_9267);
nand U9509 (N_9509,N_9286,N_9383);
xnor U9510 (N_9510,N_9269,N_9206);
nor U9511 (N_9511,N_9373,N_9274);
and U9512 (N_9512,N_9384,N_9357);
nor U9513 (N_9513,N_9214,N_9306);
nand U9514 (N_9514,N_9282,N_9231);
nand U9515 (N_9515,N_9374,N_9293);
xor U9516 (N_9516,N_9247,N_9330);
nand U9517 (N_9517,N_9274,N_9201);
and U9518 (N_9518,N_9303,N_9359);
and U9519 (N_9519,N_9308,N_9375);
and U9520 (N_9520,N_9312,N_9311);
and U9521 (N_9521,N_9305,N_9372);
nand U9522 (N_9522,N_9217,N_9279);
or U9523 (N_9523,N_9371,N_9356);
nand U9524 (N_9524,N_9205,N_9325);
and U9525 (N_9525,N_9365,N_9281);
or U9526 (N_9526,N_9228,N_9292);
and U9527 (N_9527,N_9289,N_9364);
nor U9528 (N_9528,N_9304,N_9305);
nor U9529 (N_9529,N_9319,N_9296);
nand U9530 (N_9530,N_9255,N_9328);
xnor U9531 (N_9531,N_9353,N_9228);
or U9532 (N_9532,N_9372,N_9247);
xor U9533 (N_9533,N_9263,N_9208);
and U9534 (N_9534,N_9390,N_9298);
nand U9535 (N_9535,N_9275,N_9328);
nand U9536 (N_9536,N_9348,N_9387);
nor U9537 (N_9537,N_9335,N_9358);
nand U9538 (N_9538,N_9379,N_9323);
nand U9539 (N_9539,N_9392,N_9269);
nor U9540 (N_9540,N_9253,N_9204);
nor U9541 (N_9541,N_9329,N_9211);
xnor U9542 (N_9542,N_9325,N_9375);
xnor U9543 (N_9543,N_9267,N_9368);
or U9544 (N_9544,N_9229,N_9327);
nor U9545 (N_9545,N_9290,N_9379);
or U9546 (N_9546,N_9260,N_9288);
and U9547 (N_9547,N_9337,N_9273);
and U9548 (N_9548,N_9287,N_9367);
or U9549 (N_9549,N_9268,N_9260);
or U9550 (N_9550,N_9342,N_9212);
or U9551 (N_9551,N_9267,N_9285);
nand U9552 (N_9552,N_9269,N_9238);
nand U9553 (N_9553,N_9326,N_9373);
nor U9554 (N_9554,N_9342,N_9353);
and U9555 (N_9555,N_9227,N_9309);
and U9556 (N_9556,N_9317,N_9360);
xnor U9557 (N_9557,N_9297,N_9265);
or U9558 (N_9558,N_9365,N_9264);
nand U9559 (N_9559,N_9213,N_9275);
xor U9560 (N_9560,N_9373,N_9259);
and U9561 (N_9561,N_9233,N_9356);
nand U9562 (N_9562,N_9321,N_9228);
and U9563 (N_9563,N_9262,N_9365);
xnor U9564 (N_9564,N_9234,N_9364);
or U9565 (N_9565,N_9361,N_9224);
nand U9566 (N_9566,N_9225,N_9362);
or U9567 (N_9567,N_9322,N_9390);
nand U9568 (N_9568,N_9333,N_9314);
nor U9569 (N_9569,N_9277,N_9240);
xor U9570 (N_9570,N_9369,N_9269);
xor U9571 (N_9571,N_9209,N_9228);
or U9572 (N_9572,N_9305,N_9399);
nor U9573 (N_9573,N_9203,N_9396);
xnor U9574 (N_9574,N_9251,N_9218);
xor U9575 (N_9575,N_9303,N_9238);
xnor U9576 (N_9576,N_9278,N_9224);
and U9577 (N_9577,N_9325,N_9338);
xor U9578 (N_9578,N_9352,N_9234);
nand U9579 (N_9579,N_9342,N_9221);
or U9580 (N_9580,N_9255,N_9229);
nand U9581 (N_9581,N_9271,N_9251);
and U9582 (N_9582,N_9279,N_9366);
xor U9583 (N_9583,N_9306,N_9312);
or U9584 (N_9584,N_9278,N_9357);
nor U9585 (N_9585,N_9325,N_9384);
or U9586 (N_9586,N_9297,N_9204);
or U9587 (N_9587,N_9232,N_9387);
and U9588 (N_9588,N_9214,N_9319);
nand U9589 (N_9589,N_9290,N_9361);
and U9590 (N_9590,N_9254,N_9382);
and U9591 (N_9591,N_9303,N_9271);
and U9592 (N_9592,N_9395,N_9251);
or U9593 (N_9593,N_9201,N_9365);
or U9594 (N_9594,N_9204,N_9247);
xor U9595 (N_9595,N_9264,N_9380);
and U9596 (N_9596,N_9271,N_9365);
xor U9597 (N_9597,N_9305,N_9325);
xor U9598 (N_9598,N_9361,N_9357);
or U9599 (N_9599,N_9291,N_9225);
nand U9600 (N_9600,N_9482,N_9454);
nand U9601 (N_9601,N_9502,N_9446);
nand U9602 (N_9602,N_9452,N_9453);
and U9603 (N_9603,N_9546,N_9518);
and U9604 (N_9604,N_9536,N_9577);
or U9605 (N_9605,N_9443,N_9411);
or U9606 (N_9606,N_9417,N_9590);
and U9607 (N_9607,N_9582,N_9495);
or U9608 (N_9608,N_9553,N_9477);
and U9609 (N_9609,N_9519,N_9409);
or U9610 (N_9610,N_9493,N_9548);
nand U9611 (N_9611,N_9424,N_9592);
xor U9612 (N_9612,N_9562,N_9526);
xor U9613 (N_9613,N_9494,N_9403);
nand U9614 (N_9614,N_9539,N_9547);
nand U9615 (N_9615,N_9401,N_9437);
xnor U9616 (N_9616,N_9529,N_9460);
and U9617 (N_9617,N_9595,N_9523);
or U9618 (N_9618,N_9457,N_9551);
and U9619 (N_9619,N_9400,N_9447);
xnor U9620 (N_9620,N_9418,N_9578);
xnor U9621 (N_9621,N_9522,N_9444);
nand U9622 (N_9622,N_9583,N_9517);
nor U9623 (N_9623,N_9571,N_9497);
xor U9624 (N_9624,N_9581,N_9542);
xor U9625 (N_9625,N_9511,N_9570);
nand U9626 (N_9626,N_9507,N_9534);
nand U9627 (N_9627,N_9568,N_9514);
and U9628 (N_9628,N_9470,N_9540);
and U9629 (N_9629,N_9586,N_9580);
and U9630 (N_9630,N_9427,N_9475);
and U9631 (N_9631,N_9550,N_9420);
or U9632 (N_9632,N_9563,N_9589);
and U9633 (N_9633,N_9594,N_9467);
or U9634 (N_9634,N_9431,N_9573);
and U9635 (N_9635,N_9596,N_9532);
nor U9636 (N_9636,N_9565,N_9512);
and U9637 (N_9637,N_9543,N_9561);
nand U9638 (N_9638,N_9406,N_9572);
or U9639 (N_9639,N_9433,N_9435);
or U9640 (N_9640,N_9516,N_9483);
and U9641 (N_9641,N_9429,N_9496);
nand U9642 (N_9642,N_9432,N_9498);
xnor U9643 (N_9643,N_9584,N_9405);
xnor U9644 (N_9644,N_9436,N_9557);
and U9645 (N_9645,N_9566,N_9415);
or U9646 (N_9646,N_9485,N_9520);
or U9647 (N_9647,N_9416,N_9500);
xnor U9648 (N_9648,N_9504,N_9412);
nor U9649 (N_9649,N_9556,N_9449);
or U9650 (N_9650,N_9492,N_9455);
xor U9651 (N_9651,N_9544,N_9419);
or U9652 (N_9652,N_9445,N_9508);
and U9653 (N_9653,N_9591,N_9588);
and U9654 (N_9654,N_9459,N_9468);
nand U9655 (N_9655,N_9422,N_9471);
or U9656 (N_9656,N_9491,N_9486);
or U9657 (N_9657,N_9509,N_9527);
and U9658 (N_9658,N_9441,N_9567);
nor U9659 (N_9659,N_9421,N_9537);
or U9660 (N_9660,N_9404,N_9456);
nor U9661 (N_9661,N_9465,N_9458);
xor U9662 (N_9662,N_9521,N_9484);
nand U9663 (N_9663,N_9531,N_9479);
or U9664 (N_9664,N_9451,N_9525);
or U9665 (N_9665,N_9515,N_9464);
nor U9666 (N_9666,N_9593,N_9473);
nor U9667 (N_9667,N_9513,N_9438);
nor U9668 (N_9668,N_9423,N_9439);
nor U9669 (N_9669,N_9474,N_9425);
xor U9670 (N_9670,N_9599,N_9476);
nand U9671 (N_9671,N_9524,N_9488);
nand U9672 (N_9672,N_9501,N_9559);
or U9673 (N_9673,N_9541,N_9469);
xnor U9674 (N_9674,N_9413,N_9598);
nor U9675 (N_9675,N_9450,N_9410);
nand U9676 (N_9676,N_9530,N_9461);
or U9677 (N_9677,N_9408,N_9558);
or U9678 (N_9678,N_9549,N_9402);
nor U9679 (N_9679,N_9472,N_9574);
nand U9680 (N_9680,N_9587,N_9487);
or U9681 (N_9681,N_9585,N_9407);
nand U9682 (N_9682,N_9576,N_9538);
and U9683 (N_9683,N_9597,N_9463);
nor U9684 (N_9684,N_9466,N_9428);
and U9685 (N_9685,N_9569,N_9506);
nand U9686 (N_9686,N_9554,N_9448);
nor U9687 (N_9687,N_9560,N_9535);
xnor U9688 (N_9688,N_9579,N_9564);
xnor U9689 (N_9689,N_9426,N_9462);
and U9690 (N_9690,N_9533,N_9430);
and U9691 (N_9691,N_9434,N_9480);
nor U9692 (N_9692,N_9575,N_9440);
or U9693 (N_9693,N_9552,N_9505);
xnor U9694 (N_9694,N_9442,N_9545);
nand U9695 (N_9695,N_9490,N_9510);
or U9696 (N_9696,N_9528,N_9478);
nor U9697 (N_9697,N_9503,N_9414);
nand U9698 (N_9698,N_9489,N_9481);
and U9699 (N_9699,N_9499,N_9555);
and U9700 (N_9700,N_9434,N_9597);
nor U9701 (N_9701,N_9576,N_9519);
and U9702 (N_9702,N_9530,N_9562);
nand U9703 (N_9703,N_9578,N_9554);
or U9704 (N_9704,N_9523,N_9418);
and U9705 (N_9705,N_9579,N_9522);
and U9706 (N_9706,N_9554,N_9537);
and U9707 (N_9707,N_9463,N_9536);
nor U9708 (N_9708,N_9562,N_9461);
xor U9709 (N_9709,N_9586,N_9456);
or U9710 (N_9710,N_9520,N_9466);
nand U9711 (N_9711,N_9429,N_9564);
and U9712 (N_9712,N_9464,N_9412);
and U9713 (N_9713,N_9422,N_9495);
nand U9714 (N_9714,N_9542,N_9408);
and U9715 (N_9715,N_9502,N_9467);
nor U9716 (N_9716,N_9539,N_9418);
xor U9717 (N_9717,N_9410,N_9477);
xor U9718 (N_9718,N_9512,N_9437);
and U9719 (N_9719,N_9419,N_9475);
nor U9720 (N_9720,N_9506,N_9489);
nand U9721 (N_9721,N_9511,N_9584);
nor U9722 (N_9722,N_9408,N_9434);
xor U9723 (N_9723,N_9556,N_9474);
nand U9724 (N_9724,N_9446,N_9577);
nand U9725 (N_9725,N_9555,N_9436);
nand U9726 (N_9726,N_9598,N_9593);
xor U9727 (N_9727,N_9425,N_9415);
xnor U9728 (N_9728,N_9449,N_9568);
nand U9729 (N_9729,N_9413,N_9497);
or U9730 (N_9730,N_9477,N_9552);
nand U9731 (N_9731,N_9442,N_9466);
nand U9732 (N_9732,N_9527,N_9456);
nand U9733 (N_9733,N_9503,N_9472);
and U9734 (N_9734,N_9451,N_9555);
nand U9735 (N_9735,N_9565,N_9460);
nand U9736 (N_9736,N_9472,N_9488);
xnor U9737 (N_9737,N_9464,N_9416);
or U9738 (N_9738,N_9421,N_9592);
nand U9739 (N_9739,N_9432,N_9504);
nor U9740 (N_9740,N_9531,N_9482);
xnor U9741 (N_9741,N_9577,N_9594);
or U9742 (N_9742,N_9443,N_9428);
xor U9743 (N_9743,N_9567,N_9440);
xnor U9744 (N_9744,N_9441,N_9427);
nor U9745 (N_9745,N_9541,N_9404);
or U9746 (N_9746,N_9581,N_9577);
nand U9747 (N_9747,N_9579,N_9523);
and U9748 (N_9748,N_9486,N_9460);
and U9749 (N_9749,N_9498,N_9416);
nor U9750 (N_9750,N_9433,N_9444);
nor U9751 (N_9751,N_9548,N_9407);
and U9752 (N_9752,N_9454,N_9446);
nand U9753 (N_9753,N_9500,N_9571);
nand U9754 (N_9754,N_9451,N_9478);
nor U9755 (N_9755,N_9556,N_9582);
or U9756 (N_9756,N_9485,N_9570);
xnor U9757 (N_9757,N_9570,N_9462);
and U9758 (N_9758,N_9478,N_9539);
or U9759 (N_9759,N_9542,N_9566);
and U9760 (N_9760,N_9446,N_9540);
nor U9761 (N_9761,N_9497,N_9519);
nand U9762 (N_9762,N_9468,N_9506);
nor U9763 (N_9763,N_9423,N_9526);
nand U9764 (N_9764,N_9420,N_9527);
xnor U9765 (N_9765,N_9470,N_9579);
and U9766 (N_9766,N_9430,N_9546);
xor U9767 (N_9767,N_9540,N_9415);
nor U9768 (N_9768,N_9556,N_9491);
or U9769 (N_9769,N_9402,N_9481);
nand U9770 (N_9770,N_9404,N_9565);
and U9771 (N_9771,N_9579,N_9547);
nor U9772 (N_9772,N_9590,N_9560);
or U9773 (N_9773,N_9561,N_9412);
nor U9774 (N_9774,N_9405,N_9478);
or U9775 (N_9775,N_9432,N_9462);
or U9776 (N_9776,N_9500,N_9529);
or U9777 (N_9777,N_9428,N_9419);
nand U9778 (N_9778,N_9563,N_9461);
or U9779 (N_9779,N_9549,N_9586);
xor U9780 (N_9780,N_9519,N_9405);
nand U9781 (N_9781,N_9442,N_9539);
or U9782 (N_9782,N_9537,N_9523);
xnor U9783 (N_9783,N_9577,N_9588);
xnor U9784 (N_9784,N_9569,N_9433);
and U9785 (N_9785,N_9533,N_9406);
xnor U9786 (N_9786,N_9449,N_9435);
nand U9787 (N_9787,N_9594,N_9549);
nand U9788 (N_9788,N_9593,N_9592);
nand U9789 (N_9789,N_9423,N_9552);
xor U9790 (N_9790,N_9583,N_9527);
nand U9791 (N_9791,N_9423,N_9553);
nand U9792 (N_9792,N_9413,N_9544);
nand U9793 (N_9793,N_9435,N_9438);
or U9794 (N_9794,N_9400,N_9490);
xor U9795 (N_9795,N_9413,N_9587);
xor U9796 (N_9796,N_9552,N_9459);
nor U9797 (N_9797,N_9421,N_9515);
nand U9798 (N_9798,N_9542,N_9489);
and U9799 (N_9799,N_9464,N_9549);
xnor U9800 (N_9800,N_9778,N_9667);
or U9801 (N_9801,N_9691,N_9685);
or U9802 (N_9802,N_9744,N_9791);
nor U9803 (N_9803,N_9713,N_9776);
or U9804 (N_9804,N_9754,N_9792);
nand U9805 (N_9805,N_9647,N_9747);
xnor U9806 (N_9806,N_9733,N_9614);
and U9807 (N_9807,N_9675,N_9687);
nor U9808 (N_9808,N_9704,N_9686);
xor U9809 (N_9809,N_9777,N_9746);
or U9810 (N_9810,N_9728,N_9715);
and U9811 (N_9811,N_9659,N_9620);
nand U9812 (N_9812,N_9642,N_9796);
or U9813 (N_9813,N_9718,N_9677);
nand U9814 (N_9814,N_9722,N_9767);
or U9815 (N_9815,N_9775,N_9731);
and U9816 (N_9816,N_9708,N_9768);
xnor U9817 (N_9817,N_9612,N_9751);
and U9818 (N_9818,N_9764,N_9712);
nor U9819 (N_9819,N_9700,N_9748);
xor U9820 (N_9820,N_9716,N_9649);
or U9821 (N_9821,N_9672,N_9654);
nand U9822 (N_9822,N_9624,N_9782);
and U9823 (N_9823,N_9710,N_9779);
xnor U9824 (N_9824,N_9636,N_9780);
or U9825 (N_9825,N_9735,N_9656);
xor U9826 (N_9826,N_9641,N_9798);
or U9827 (N_9827,N_9671,N_9772);
or U9828 (N_9828,N_9734,N_9678);
or U9829 (N_9829,N_9695,N_9773);
and U9830 (N_9830,N_9669,N_9635);
nor U9831 (N_9831,N_9762,N_9757);
or U9832 (N_9832,N_9799,N_9707);
and U9833 (N_9833,N_9766,N_9615);
or U9834 (N_9834,N_9787,N_9692);
xor U9835 (N_9835,N_9632,N_9725);
nor U9836 (N_9836,N_9771,N_9627);
and U9837 (N_9837,N_9730,N_9786);
and U9838 (N_9838,N_9797,N_9702);
and U9839 (N_9839,N_9619,N_9626);
nand U9840 (N_9840,N_9664,N_9770);
or U9841 (N_9841,N_9660,N_9701);
xnor U9842 (N_9842,N_9658,N_9765);
xor U9843 (N_9843,N_9613,N_9753);
nand U9844 (N_9844,N_9737,N_9655);
and U9845 (N_9845,N_9629,N_9645);
and U9846 (N_9846,N_9682,N_9750);
xnor U9847 (N_9847,N_9650,N_9665);
or U9848 (N_9848,N_9604,N_9607);
nor U9849 (N_9849,N_9657,N_9760);
and U9850 (N_9850,N_9758,N_9668);
or U9851 (N_9851,N_9745,N_9783);
nand U9852 (N_9852,N_9699,N_9674);
nand U9853 (N_9853,N_9774,N_9652);
xnor U9854 (N_9854,N_9644,N_9690);
and U9855 (N_9855,N_9601,N_9633);
and U9856 (N_9856,N_9653,N_9638);
and U9857 (N_9857,N_9663,N_9666);
and U9858 (N_9858,N_9742,N_9739);
and U9859 (N_9859,N_9609,N_9698);
xnor U9860 (N_9860,N_9784,N_9679);
nand U9861 (N_9861,N_9608,N_9683);
nor U9862 (N_9862,N_9617,N_9661);
nor U9863 (N_9863,N_9714,N_9749);
nand U9864 (N_9864,N_9711,N_9673);
and U9865 (N_9865,N_9606,N_9769);
xnor U9866 (N_9866,N_9724,N_9696);
or U9867 (N_9867,N_9684,N_9706);
xor U9868 (N_9868,N_9732,N_9621);
nor U9869 (N_9869,N_9648,N_9729);
nor U9870 (N_9870,N_9788,N_9662);
nor U9871 (N_9871,N_9727,N_9651);
and U9872 (N_9872,N_9605,N_9631);
nor U9873 (N_9873,N_9743,N_9600);
or U9874 (N_9874,N_9640,N_9759);
nand U9875 (N_9875,N_9622,N_9736);
nand U9876 (N_9876,N_9625,N_9602);
and U9877 (N_9877,N_9793,N_9785);
xor U9878 (N_9878,N_9639,N_9789);
or U9879 (N_9879,N_9681,N_9738);
or U9880 (N_9880,N_9670,N_9705);
xnor U9881 (N_9881,N_9623,N_9721);
or U9882 (N_9882,N_9741,N_9740);
or U9883 (N_9883,N_9697,N_9781);
nor U9884 (N_9884,N_9703,N_9763);
and U9885 (N_9885,N_9628,N_9616);
nor U9886 (N_9886,N_9795,N_9611);
xnor U9887 (N_9887,N_9755,N_9761);
or U9888 (N_9888,N_9680,N_9694);
nor U9889 (N_9889,N_9618,N_9603);
nor U9890 (N_9890,N_9693,N_9717);
nand U9891 (N_9891,N_9794,N_9610);
xor U9892 (N_9892,N_9752,N_9676);
nor U9893 (N_9893,N_9688,N_9723);
or U9894 (N_9894,N_9720,N_9646);
or U9895 (N_9895,N_9689,N_9790);
or U9896 (N_9896,N_9643,N_9634);
and U9897 (N_9897,N_9756,N_9709);
or U9898 (N_9898,N_9630,N_9726);
or U9899 (N_9899,N_9637,N_9719);
xnor U9900 (N_9900,N_9627,N_9675);
and U9901 (N_9901,N_9787,N_9661);
xor U9902 (N_9902,N_9790,N_9711);
or U9903 (N_9903,N_9684,N_9711);
xnor U9904 (N_9904,N_9770,N_9622);
and U9905 (N_9905,N_9644,N_9701);
or U9906 (N_9906,N_9778,N_9616);
nor U9907 (N_9907,N_9763,N_9778);
or U9908 (N_9908,N_9733,N_9696);
nand U9909 (N_9909,N_9765,N_9638);
or U9910 (N_9910,N_9614,N_9717);
or U9911 (N_9911,N_9751,N_9631);
nand U9912 (N_9912,N_9762,N_9642);
and U9913 (N_9913,N_9753,N_9796);
or U9914 (N_9914,N_9659,N_9661);
or U9915 (N_9915,N_9715,N_9606);
nand U9916 (N_9916,N_9678,N_9722);
xor U9917 (N_9917,N_9761,N_9743);
nor U9918 (N_9918,N_9622,N_9691);
and U9919 (N_9919,N_9691,N_9695);
nand U9920 (N_9920,N_9642,N_9790);
xnor U9921 (N_9921,N_9754,N_9623);
nor U9922 (N_9922,N_9741,N_9636);
and U9923 (N_9923,N_9751,N_9790);
or U9924 (N_9924,N_9639,N_9758);
and U9925 (N_9925,N_9740,N_9756);
or U9926 (N_9926,N_9765,N_9785);
and U9927 (N_9927,N_9663,N_9676);
or U9928 (N_9928,N_9670,N_9735);
and U9929 (N_9929,N_9736,N_9767);
nor U9930 (N_9930,N_9670,N_9687);
or U9931 (N_9931,N_9747,N_9650);
and U9932 (N_9932,N_9697,N_9794);
and U9933 (N_9933,N_9671,N_9642);
xnor U9934 (N_9934,N_9779,N_9632);
xor U9935 (N_9935,N_9718,N_9727);
nor U9936 (N_9936,N_9697,N_9620);
nand U9937 (N_9937,N_9643,N_9694);
nand U9938 (N_9938,N_9670,N_9723);
and U9939 (N_9939,N_9617,N_9612);
nor U9940 (N_9940,N_9785,N_9796);
or U9941 (N_9941,N_9697,N_9708);
xor U9942 (N_9942,N_9675,N_9692);
xor U9943 (N_9943,N_9661,N_9605);
nand U9944 (N_9944,N_9724,N_9723);
or U9945 (N_9945,N_9722,N_9642);
xnor U9946 (N_9946,N_9661,N_9604);
nor U9947 (N_9947,N_9746,N_9723);
or U9948 (N_9948,N_9684,N_9695);
xnor U9949 (N_9949,N_9723,N_9645);
and U9950 (N_9950,N_9706,N_9758);
nor U9951 (N_9951,N_9790,N_9733);
and U9952 (N_9952,N_9665,N_9718);
and U9953 (N_9953,N_9748,N_9765);
or U9954 (N_9954,N_9738,N_9730);
and U9955 (N_9955,N_9693,N_9600);
nor U9956 (N_9956,N_9674,N_9668);
xnor U9957 (N_9957,N_9618,N_9613);
or U9958 (N_9958,N_9632,N_9665);
nand U9959 (N_9959,N_9799,N_9640);
nand U9960 (N_9960,N_9676,N_9766);
or U9961 (N_9961,N_9631,N_9760);
xor U9962 (N_9962,N_9739,N_9679);
xor U9963 (N_9963,N_9784,N_9668);
xor U9964 (N_9964,N_9630,N_9696);
and U9965 (N_9965,N_9704,N_9635);
and U9966 (N_9966,N_9768,N_9652);
nand U9967 (N_9967,N_9734,N_9649);
or U9968 (N_9968,N_9748,N_9644);
and U9969 (N_9969,N_9639,N_9667);
nand U9970 (N_9970,N_9673,N_9758);
or U9971 (N_9971,N_9687,N_9610);
nor U9972 (N_9972,N_9676,N_9797);
and U9973 (N_9973,N_9634,N_9742);
xnor U9974 (N_9974,N_9736,N_9626);
nand U9975 (N_9975,N_9732,N_9619);
nand U9976 (N_9976,N_9788,N_9606);
nor U9977 (N_9977,N_9796,N_9776);
xor U9978 (N_9978,N_9790,N_9702);
nor U9979 (N_9979,N_9631,N_9601);
nand U9980 (N_9980,N_9628,N_9666);
xor U9981 (N_9981,N_9647,N_9671);
nor U9982 (N_9982,N_9661,N_9715);
or U9983 (N_9983,N_9766,N_9643);
and U9984 (N_9984,N_9786,N_9667);
or U9985 (N_9985,N_9640,N_9723);
nand U9986 (N_9986,N_9755,N_9764);
or U9987 (N_9987,N_9752,N_9624);
or U9988 (N_9988,N_9631,N_9654);
xnor U9989 (N_9989,N_9748,N_9648);
nor U9990 (N_9990,N_9751,N_9618);
or U9991 (N_9991,N_9660,N_9608);
nand U9992 (N_9992,N_9746,N_9750);
nand U9993 (N_9993,N_9603,N_9738);
and U9994 (N_9994,N_9683,N_9704);
and U9995 (N_9995,N_9703,N_9691);
nand U9996 (N_9996,N_9667,N_9737);
nor U9997 (N_9997,N_9646,N_9718);
and U9998 (N_9998,N_9662,N_9742);
xnor U9999 (N_9999,N_9762,N_9740);
or UO_0 (O_0,N_9867,N_9930);
nor UO_1 (O_1,N_9936,N_9971);
and UO_2 (O_2,N_9833,N_9803);
nand UO_3 (O_3,N_9885,N_9922);
nand UO_4 (O_4,N_9850,N_9828);
xnor UO_5 (O_5,N_9906,N_9880);
nand UO_6 (O_6,N_9998,N_9871);
xnor UO_7 (O_7,N_9895,N_9877);
xnor UO_8 (O_8,N_9851,N_9921);
and UO_9 (O_9,N_9980,N_9959);
nand UO_10 (O_10,N_9802,N_9947);
nor UO_11 (O_11,N_9812,N_9960);
xor UO_12 (O_12,N_9809,N_9990);
and UO_13 (O_13,N_9985,N_9887);
and UO_14 (O_14,N_9932,N_9912);
or UO_15 (O_15,N_9934,N_9909);
xor UO_16 (O_16,N_9962,N_9869);
or UO_17 (O_17,N_9911,N_9857);
nand UO_18 (O_18,N_9879,N_9847);
nor UO_19 (O_19,N_9839,N_9993);
xnor UO_20 (O_20,N_9891,N_9899);
and UO_21 (O_21,N_9863,N_9830);
nor UO_22 (O_22,N_9870,N_9928);
xnor UO_23 (O_23,N_9840,N_9996);
nand UO_24 (O_24,N_9817,N_9826);
nor UO_25 (O_25,N_9935,N_9991);
xnor UO_26 (O_26,N_9805,N_9968);
nand UO_27 (O_27,N_9836,N_9868);
or UO_28 (O_28,N_9919,N_9908);
or UO_29 (O_29,N_9982,N_9862);
nand UO_30 (O_30,N_9858,N_9981);
or UO_31 (O_31,N_9964,N_9856);
nor UO_32 (O_32,N_9986,N_9855);
xor UO_33 (O_33,N_9854,N_9929);
nand UO_34 (O_34,N_9910,N_9952);
nor UO_35 (O_35,N_9907,N_9810);
xnor UO_36 (O_36,N_9835,N_9811);
nand UO_37 (O_37,N_9973,N_9834);
xor UO_38 (O_38,N_9997,N_9951);
xnor UO_39 (O_39,N_9937,N_9963);
xor UO_40 (O_40,N_9859,N_9975);
or UO_41 (O_41,N_9864,N_9902);
xnor UO_42 (O_42,N_9894,N_9820);
or UO_43 (O_43,N_9819,N_9804);
xor UO_44 (O_44,N_9976,N_9886);
or UO_45 (O_45,N_9970,N_9942);
nor UO_46 (O_46,N_9861,N_9961);
or UO_47 (O_47,N_9876,N_9829);
or UO_48 (O_48,N_9845,N_9989);
or UO_49 (O_49,N_9925,N_9949);
nand UO_50 (O_50,N_9977,N_9875);
xor UO_51 (O_51,N_9822,N_9866);
or UO_52 (O_52,N_9821,N_9939);
xnor UO_53 (O_53,N_9837,N_9865);
or UO_54 (O_54,N_9943,N_9883);
nand UO_55 (O_55,N_9815,N_9843);
nand UO_56 (O_56,N_9846,N_9941);
and UO_57 (O_57,N_9882,N_9860);
nand UO_58 (O_58,N_9931,N_9966);
nand UO_59 (O_59,N_9974,N_9901);
or UO_60 (O_60,N_9965,N_9923);
nor UO_61 (O_61,N_9889,N_9916);
nor UO_62 (O_62,N_9946,N_9983);
xor UO_63 (O_63,N_9823,N_9915);
and UO_64 (O_64,N_9994,N_9806);
nor UO_65 (O_65,N_9853,N_9944);
nand UO_66 (O_66,N_9933,N_9918);
nand UO_67 (O_67,N_9953,N_9967);
or UO_68 (O_68,N_9954,N_9992);
or UO_69 (O_69,N_9984,N_9898);
nor UO_70 (O_70,N_9844,N_9948);
nor UO_71 (O_71,N_9999,N_9813);
and UO_72 (O_72,N_9800,N_9940);
nor UO_73 (O_73,N_9957,N_9878);
nand UO_74 (O_74,N_9874,N_9824);
nor UO_75 (O_75,N_9841,N_9924);
nor UO_76 (O_76,N_9888,N_9913);
or UO_77 (O_77,N_9927,N_9988);
nand UO_78 (O_78,N_9827,N_9920);
nor UO_79 (O_79,N_9938,N_9842);
xor UO_80 (O_80,N_9905,N_9979);
or UO_81 (O_81,N_9872,N_9903);
or UO_82 (O_82,N_9917,N_9890);
xnor UO_83 (O_83,N_9848,N_9852);
nand UO_84 (O_84,N_9893,N_9897);
nor UO_85 (O_85,N_9900,N_9816);
nand UO_86 (O_86,N_9896,N_9950);
or UO_87 (O_87,N_9825,N_9801);
or UO_88 (O_88,N_9884,N_9892);
and UO_89 (O_89,N_9978,N_9987);
and UO_90 (O_90,N_9814,N_9838);
or UO_91 (O_91,N_9958,N_9831);
nand UO_92 (O_92,N_9832,N_9881);
nor UO_93 (O_93,N_9849,N_9873);
nor UO_94 (O_94,N_9904,N_9955);
and UO_95 (O_95,N_9995,N_9926);
xor UO_96 (O_96,N_9818,N_9969);
or UO_97 (O_97,N_9956,N_9945);
nor UO_98 (O_98,N_9972,N_9914);
or UO_99 (O_99,N_9807,N_9808);
nand UO_100 (O_100,N_9887,N_9828);
or UO_101 (O_101,N_9904,N_9927);
nand UO_102 (O_102,N_9967,N_9870);
or UO_103 (O_103,N_9971,N_9800);
nand UO_104 (O_104,N_9855,N_9807);
xor UO_105 (O_105,N_9911,N_9993);
and UO_106 (O_106,N_9830,N_9904);
and UO_107 (O_107,N_9866,N_9881);
nor UO_108 (O_108,N_9887,N_9912);
xor UO_109 (O_109,N_9824,N_9916);
nand UO_110 (O_110,N_9972,N_9885);
and UO_111 (O_111,N_9808,N_9852);
or UO_112 (O_112,N_9819,N_9933);
nand UO_113 (O_113,N_9809,N_9846);
or UO_114 (O_114,N_9877,N_9907);
nor UO_115 (O_115,N_9856,N_9998);
or UO_116 (O_116,N_9859,N_9911);
nand UO_117 (O_117,N_9998,N_9863);
nor UO_118 (O_118,N_9822,N_9844);
and UO_119 (O_119,N_9847,N_9943);
and UO_120 (O_120,N_9956,N_9811);
and UO_121 (O_121,N_9810,N_9880);
nand UO_122 (O_122,N_9956,N_9971);
and UO_123 (O_123,N_9965,N_9883);
nand UO_124 (O_124,N_9822,N_9927);
nor UO_125 (O_125,N_9994,N_9990);
or UO_126 (O_126,N_9995,N_9929);
nor UO_127 (O_127,N_9847,N_9856);
or UO_128 (O_128,N_9880,N_9948);
or UO_129 (O_129,N_9833,N_9934);
and UO_130 (O_130,N_9959,N_9873);
nand UO_131 (O_131,N_9920,N_9935);
or UO_132 (O_132,N_9840,N_9815);
nor UO_133 (O_133,N_9911,N_9974);
or UO_134 (O_134,N_9974,N_9828);
and UO_135 (O_135,N_9970,N_9922);
nand UO_136 (O_136,N_9823,N_9863);
nor UO_137 (O_137,N_9866,N_9972);
xor UO_138 (O_138,N_9935,N_9831);
nor UO_139 (O_139,N_9897,N_9914);
xnor UO_140 (O_140,N_9887,N_9816);
xor UO_141 (O_141,N_9876,N_9826);
or UO_142 (O_142,N_9918,N_9915);
and UO_143 (O_143,N_9997,N_9908);
nor UO_144 (O_144,N_9905,N_9909);
nor UO_145 (O_145,N_9955,N_9939);
nor UO_146 (O_146,N_9930,N_9956);
nor UO_147 (O_147,N_9988,N_9982);
xor UO_148 (O_148,N_9862,N_9901);
or UO_149 (O_149,N_9847,N_9832);
nor UO_150 (O_150,N_9896,N_9863);
nand UO_151 (O_151,N_9958,N_9822);
xor UO_152 (O_152,N_9914,N_9861);
nand UO_153 (O_153,N_9892,N_9807);
nand UO_154 (O_154,N_9802,N_9912);
nand UO_155 (O_155,N_9923,N_9906);
or UO_156 (O_156,N_9917,N_9840);
xnor UO_157 (O_157,N_9857,N_9949);
nor UO_158 (O_158,N_9824,N_9808);
nor UO_159 (O_159,N_9820,N_9926);
and UO_160 (O_160,N_9987,N_9923);
nor UO_161 (O_161,N_9860,N_9996);
nor UO_162 (O_162,N_9995,N_9834);
or UO_163 (O_163,N_9949,N_9897);
and UO_164 (O_164,N_9818,N_9868);
nor UO_165 (O_165,N_9939,N_9820);
and UO_166 (O_166,N_9861,N_9876);
or UO_167 (O_167,N_9958,N_9933);
xor UO_168 (O_168,N_9907,N_9974);
or UO_169 (O_169,N_9923,N_9851);
and UO_170 (O_170,N_9915,N_9891);
or UO_171 (O_171,N_9956,N_9914);
nand UO_172 (O_172,N_9833,N_9844);
or UO_173 (O_173,N_9970,N_9907);
xnor UO_174 (O_174,N_9914,N_9976);
nand UO_175 (O_175,N_9850,N_9976);
or UO_176 (O_176,N_9894,N_9973);
nor UO_177 (O_177,N_9876,N_9897);
xnor UO_178 (O_178,N_9952,N_9997);
nand UO_179 (O_179,N_9819,N_9963);
nand UO_180 (O_180,N_9859,N_9891);
nand UO_181 (O_181,N_9949,N_9800);
or UO_182 (O_182,N_9801,N_9806);
nand UO_183 (O_183,N_9821,N_9857);
and UO_184 (O_184,N_9874,N_9944);
xor UO_185 (O_185,N_9800,N_9937);
nand UO_186 (O_186,N_9989,N_9954);
or UO_187 (O_187,N_9963,N_9887);
nor UO_188 (O_188,N_9980,N_9944);
or UO_189 (O_189,N_9841,N_9878);
xnor UO_190 (O_190,N_9943,N_9822);
nand UO_191 (O_191,N_9996,N_9810);
nand UO_192 (O_192,N_9878,N_9938);
nand UO_193 (O_193,N_9936,N_9900);
nor UO_194 (O_194,N_9923,N_9857);
or UO_195 (O_195,N_9902,N_9900);
and UO_196 (O_196,N_9960,N_9883);
and UO_197 (O_197,N_9892,N_9980);
and UO_198 (O_198,N_9883,N_9817);
or UO_199 (O_199,N_9940,N_9966);
xor UO_200 (O_200,N_9927,N_9861);
nor UO_201 (O_201,N_9807,N_9806);
nor UO_202 (O_202,N_9985,N_9916);
or UO_203 (O_203,N_9994,N_9825);
and UO_204 (O_204,N_9821,N_9844);
and UO_205 (O_205,N_9895,N_9823);
or UO_206 (O_206,N_9957,N_9814);
or UO_207 (O_207,N_9861,N_9805);
or UO_208 (O_208,N_9821,N_9979);
xor UO_209 (O_209,N_9869,N_9978);
xnor UO_210 (O_210,N_9899,N_9999);
or UO_211 (O_211,N_9875,N_9854);
xnor UO_212 (O_212,N_9808,N_9880);
nor UO_213 (O_213,N_9986,N_9964);
or UO_214 (O_214,N_9918,N_9862);
or UO_215 (O_215,N_9893,N_9877);
nand UO_216 (O_216,N_9942,N_9999);
nand UO_217 (O_217,N_9891,N_9842);
and UO_218 (O_218,N_9996,N_9902);
and UO_219 (O_219,N_9814,N_9850);
xor UO_220 (O_220,N_9847,N_9985);
or UO_221 (O_221,N_9860,N_9981);
and UO_222 (O_222,N_9863,N_9862);
and UO_223 (O_223,N_9945,N_9821);
and UO_224 (O_224,N_9945,N_9834);
nand UO_225 (O_225,N_9968,N_9845);
nor UO_226 (O_226,N_9826,N_9928);
or UO_227 (O_227,N_9883,N_9916);
nand UO_228 (O_228,N_9815,N_9803);
nor UO_229 (O_229,N_9893,N_9915);
or UO_230 (O_230,N_9983,N_9947);
nand UO_231 (O_231,N_9886,N_9804);
xnor UO_232 (O_232,N_9867,N_9847);
xor UO_233 (O_233,N_9864,N_9913);
xnor UO_234 (O_234,N_9867,N_9895);
nand UO_235 (O_235,N_9937,N_9811);
or UO_236 (O_236,N_9999,N_9938);
nor UO_237 (O_237,N_9830,N_9846);
and UO_238 (O_238,N_9922,N_9898);
nand UO_239 (O_239,N_9903,N_9818);
and UO_240 (O_240,N_9933,N_9886);
or UO_241 (O_241,N_9978,N_9972);
nand UO_242 (O_242,N_9842,N_9845);
nand UO_243 (O_243,N_9851,N_9896);
nor UO_244 (O_244,N_9851,N_9828);
nand UO_245 (O_245,N_9915,N_9924);
nand UO_246 (O_246,N_9928,N_9988);
and UO_247 (O_247,N_9877,N_9865);
xnor UO_248 (O_248,N_9880,N_9855);
nor UO_249 (O_249,N_9836,N_9960);
nand UO_250 (O_250,N_9842,N_9961);
xnor UO_251 (O_251,N_9972,N_9812);
xnor UO_252 (O_252,N_9859,N_9840);
and UO_253 (O_253,N_9849,N_9960);
nand UO_254 (O_254,N_9838,N_9856);
nand UO_255 (O_255,N_9869,N_9853);
or UO_256 (O_256,N_9915,N_9933);
nor UO_257 (O_257,N_9867,N_9912);
xor UO_258 (O_258,N_9831,N_9967);
nor UO_259 (O_259,N_9948,N_9995);
nand UO_260 (O_260,N_9925,N_9903);
and UO_261 (O_261,N_9830,N_9970);
xnor UO_262 (O_262,N_9939,N_9886);
nor UO_263 (O_263,N_9817,N_9930);
and UO_264 (O_264,N_9986,N_9807);
nor UO_265 (O_265,N_9951,N_9974);
nand UO_266 (O_266,N_9994,N_9931);
and UO_267 (O_267,N_9825,N_9870);
or UO_268 (O_268,N_9815,N_9995);
xnor UO_269 (O_269,N_9803,N_9813);
or UO_270 (O_270,N_9840,N_9909);
or UO_271 (O_271,N_9803,N_9912);
nand UO_272 (O_272,N_9807,N_9976);
xnor UO_273 (O_273,N_9917,N_9893);
xnor UO_274 (O_274,N_9985,N_9807);
xnor UO_275 (O_275,N_9878,N_9813);
and UO_276 (O_276,N_9969,N_9850);
or UO_277 (O_277,N_9970,N_9855);
nand UO_278 (O_278,N_9911,N_9810);
and UO_279 (O_279,N_9927,N_9913);
nand UO_280 (O_280,N_9841,N_9990);
and UO_281 (O_281,N_9998,N_9847);
and UO_282 (O_282,N_9900,N_9806);
xnor UO_283 (O_283,N_9895,N_9990);
or UO_284 (O_284,N_9944,N_9838);
nand UO_285 (O_285,N_9945,N_9927);
nand UO_286 (O_286,N_9840,N_9941);
or UO_287 (O_287,N_9802,N_9918);
or UO_288 (O_288,N_9878,N_9988);
and UO_289 (O_289,N_9980,N_9916);
and UO_290 (O_290,N_9877,N_9894);
or UO_291 (O_291,N_9941,N_9967);
xnor UO_292 (O_292,N_9995,N_9890);
nor UO_293 (O_293,N_9962,N_9986);
nand UO_294 (O_294,N_9960,N_9998);
nand UO_295 (O_295,N_9862,N_9845);
xor UO_296 (O_296,N_9967,N_9971);
nor UO_297 (O_297,N_9902,N_9923);
nand UO_298 (O_298,N_9990,N_9853);
xor UO_299 (O_299,N_9888,N_9810);
xor UO_300 (O_300,N_9829,N_9933);
or UO_301 (O_301,N_9890,N_9994);
and UO_302 (O_302,N_9815,N_9997);
or UO_303 (O_303,N_9979,N_9988);
xor UO_304 (O_304,N_9804,N_9902);
nand UO_305 (O_305,N_9920,N_9936);
nand UO_306 (O_306,N_9893,N_9883);
or UO_307 (O_307,N_9838,N_9854);
and UO_308 (O_308,N_9964,N_9962);
xor UO_309 (O_309,N_9827,N_9948);
and UO_310 (O_310,N_9866,N_9908);
or UO_311 (O_311,N_9947,N_9810);
nor UO_312 (O_312,N_9952,N_9844);
nor UO_313 (O_313,N_9894,N_9872);
nand UO_314 (O_314,N_9848,N_9800);
nand UO_315 (O_315,N_9971,N_9889);
or UO_316 (O_316,N_9902,N_9824);
nor UO_317 (O_317,N_9869,N_9917);
nor UO_318 (O_318,N_9834,N_9882);
nor UO_319 (O_319,N_9816,N_9851);
and UO_320 (O_320,N_9865,N_9843);
or UO_321 (O_321,N_9915,N_9909);
xor UO_322 (O_322,N_9965,N_9897);
or UO_323 (O_323,N_9981,N_9896);
or UO_324 (O_324,N_9935,N_9990);
xnor UO_325 (O_325,N_9881,N_9985);
xnor UO_326 (O_326,N_9936,N_9959);
nand UO_327 (O_327,N_9858,N_9841);
and UO_328 (O_328,N_9938,N_9943);
and UO_329 (O_329,N_9841,N_9965);
xor UO_330 (O_330,N_9868,N_9821);
or UO_331 (O_331,N_9941,N_9977);
nor UO_332 (O_332,N_9801,N_9927);
and UO_333 (O_333,N_9880,N_9827);
nand UO_334 (O_334,N_9948,N_9845);
xor UO_335 (O_335,N_9841,N_9928);
xnor UO_336 (O_336,N_9851,N_9847);
and UO_337 (O_337,N_9836,N_9970);
nand UO_338 (O_338,N_9917,N_9921);
and UO_339 (O_339,N_9901,N_9831);
and UO_340 (O_340,N_9967,N_9991);
nand UO_341 (O_341,N_9880,N_9963);
or UO_342 (O_342,N_9942,N_9819);
nand UO_343 (O_343,N_9903,N_9908);
xnor UO_344 (O_344,N_9879,N_9978);
and UO_345 (O_345,N_9992,N_9985);
xnor UO_346 (O_346,N_9940,N_9841);
xnor UO_347 (O_347,N_9842,N_9833);
xnor UO_348 (O_348,N_9967,N_9888);
nor UO_349 (O_349,N_9806,N_9870);
nor UO_350 (O_350,N_9842,N_9974);
xnor UO_351 (O_351,N_9824,N_9884);
nor UO_352 (O_352,N_9991,N_9862);
and UO_353 (O_353,N_9998,N_9818);
nand UO_354 (O_354,N_9897,N_9919);
nor UO_355 (O_355,N_9932,N_9964);
or UO_356 (O_356,N_9889,N_9952);
nor UO_357 (O_357,N_9824,N_9843);
xor UO_358 (O_358,N_9863,N_9831);
and UO_359 (O_359,N_9884,N_9986);
nor UO_360 (O_360,N_9996,N_9845);
and UO_361 (O_361,N_9889,N_9905);
nor UO_362 (O_362,N_9924,N_9869);
and UO_363 (O_363,N_9801,N_9947);
and UO_364 (O_364,N_9918,N_9844);
nor UO_365 (O_365,N_9938,N_9954);
nor UO_366 (O_366,N_9883,N_9990);
nand UO_367 (O_367,N_9840,N_9858);
and UO_368 (O_368,N_9962,N_9865);
or UO_369 (O_369,N_9945,N_9932);
nor UO_370 (O_370,N_9922,N_9996);
nand UO_371 (O_371,N_9891,N_9818);
or UO_372 (O_372,N_9810,N_9910);
or UO_373 (O_373,N_9932,N_9911);
nor UO_374 (O_374,N_9917,N_9968);
or UO_375 (O_375,N_9818,N_9846);
nor UO_376 (O_376,N_9990,N_9810);
nor UO_377 (O_377,N_9954,N_9854);
and UO_378 (O_378,N_9817,N_9990);
and UO_379 (O_379,N_9970,N_9971);
xor UO_380 (O_380,N_9895,N_9850);
nand UO_381 (O_381,N_9955,N_9862);
or UO_382 (O_382,N_9996,N_9862);
or UO_383 (O_383,N_9831,N_9914);
or UO_384 (O_384,N_9982,N_9803);
nand UO_385 (O_385,N_9994,N_9851);
nor UO_386 (O_386,N_9837,N_9871);
nor UO_387 (O_387,N_9822,N_9846);
nand UO_388 (O_388,N_9940,N_9858);
xnor UO_389 (O_389,N_9886,N_9967);
nor UO_390 (O_390,N_9975,N_9990);
xnor UO_391 (O_391,N_9873,N_9856);
xnor UO_392 (O_392,N_9819,N_9801);
nand UO_393 (O_393,N_9925,N_9937);
or UO_394 (O_394,N_9932,N_9904);
xnor UO_395 (O_395,N_9923,N_9936);
nand UO_396 (O_396,N_9985,N_9871);
nor UO_397 (O_397,N_9858,N_9867);
or UO_398 (O_398,N_9955,N_9922);
or UO_399 (O_399,N_9900,N_9910);
xor UO_400 (O_400,N_9925,N_9915);
xnor UO_401 (O_401,N_9839,N_9991);
nor UO_402 (O_402,N_9851,N_9973);
nand UO_403 (O_403,N_9879,N_9882);
and UO_404 (O_404,N_9891,N_9908);
nand UO_405 (O_405,N_9973,N_9858);
nand UO_406 (O_406,N_9834,N_9850);
and UO_407 (O_407,N_9994,N_9966);
or UO_408 (O_408,N_9884,N_9929);
and UO_409 (O_409,N_9897,N_9827);
nand UO_410 (O_410,N_9855,N_9898);
and UO_411 (O_411,N_9951,N_9890);
and UO_412 (O_412,N_9953,N_9860);
nor UO_413 (O_413,N_9957,N_9964);
or UO_414 (O_414,N_9940,N_9946);
or UO_415 (O_415,N_9955,N_9832);
nand UO_416 (O_416,N_9837,N_9985);
nor UO_417 (O_417,N_9986,N_9823);
nand UO_418 (O_418,N_9841,N_9916);
xnor UO_419 (O_419,N_9928,N_9881);
xor UO_420 (O_420,N_9838,N_9915);
or UO_421 (O_421,N_9963,N_9869);
and UO_422 (O_422,N_9801,N_9945);
nor UO_423 (O_423,N_9857,N_9886);
nand UO_424 (O_424,N_9811,N_9948);
or UO_425 (O_425,N_9867,N_9836);
nor UO_426 (O_426,N_9956,N_9909);
and UO_427 (O_427,N_9846,N_9927);
xnor UO_428 (O_428,N_9893,N_9821);
nand UO_429 (O_429,N_9869,N_9952);
or UO_430 (O_430,N_9968,N_9974);
nor UO_431 (O_431,N_9919,N_9947);
and UO_432 (O_432,N_9836,N_9907);
nor UO_433 (O_433,N_9859,N_9848);
nor UO_434 (O_434,N_9980,N_9895);
or UO_435 (O_435,N_9854,N_9836);
or UO_436 (O_436,N_9908,N_9935);
and UO_437 (O_437,N_9965,N_9815);
nand UO_438 (O_438,N_9867,N_9871);
or UO_439 (O_439,N_9880,N_9874);
nor UO_440 (O_440,N_9873,N_9948);
xor UO_441 (O_441,N_9817,N_9914);
and UO_442 (O_442,N_9826,N_9894);
xor UO_443 (O_443,N_9948,N_9896);
or UO_444 (O_444,N_9811,N_9806);
and UO_445 (O_445,N_9817,N_9961);
nor UO_446 (O_446,N_9824,N_9994);
nor UO_447 (O_447,N_9995,N_9899);
or UO_448 (O_448,N_9804,N_9973);
nor UO_449 (O_449,N_9940,N_9825);
or UO_450 (O_450,N_9979,N_9820);
xor UO_451 (O_451,N_9975,N_9804);
xor UO_452 (O_452,N_9894,N_9908);
or UO_453 (O_453,N_9916,N_9964);
nor UO_454 (O_454,N_9865,N_9801);
and UO_455 (O_455,N_9822,N_9869);
or UO_456 (O_456,N_9987,N_9939);
and UO_457 (O_457,N_9876,N_9816);
and UO_458 (O_458,N_9969,N_9978);
and UO_459 (O_459,N_9896,N_9971);
nand UO_460 (O_460,N_9960,N_9928);
nor UO_461 (O_461,N_9801,N_9908);
nor UO_462 (O_462,N_9866,N_9905);
nor UO_463 (O_463,N_9901,N_9986);
and UO_464 (O_464,N_9917,N_9879);
nand UO_465 (O_465,N_9859,N_9872);
xnor UO_466 (O_466,N_9900,N_9808);
or UO_467 (O_467,N_9934,N_9876);
and UO_468 (O_468,N_9939,N_9816);
and UO_469 (O_469,N_9830,N_9984);
nand UO_470 (O_470,N_9978,N_9974);
nand UO_471 (O_471,N_9976,N_9942);
xor UO_472 (O_472,N_9954,N_9940);
nor UO_473 (O_473,N_9906,N_9856);
or UO_474 (O_474,N_9908,N_9879);
or UO_475 (O_475,N_9993,N_9801);
and UO_476 (O_476,N_9904,N_9940);
nor UO_477 (O_477,N_9865,N_9933);
or UO_478 (O_478,N_9894,N_9800);
xor UO_479 (O_479,N_9963,N_9873);
and UO_480 (O_480,N_9948,N_9831);
or UO_481 (O_481,N_9874,N_9847);
nand UO_482 (O_482,N_9973,N_9811);
or UO_483 (O_483,N_9809,N_9810);
nor UO_484 (O_484,N_9867,N_9954);
xnor UO_485 (O_485,N_9984,N_9925);
xor UO_486 (O_486,N_9833,N_9917);
nor UO_487 (O_487,N_9944,N_9818);
nor UO_488 (O_488,N_9908,N_9960);
nor UO_489 (O_489,N_9867,N_9827);
nand UO_490 (O_490,N_9862,N_9827);
and UO_491 (O_491,N_9874,N_9940);
nand UO_492 (O_492,N_9916,N_9870);
or UO_493 (O_493,N_9890,N_9954);
nor UO_494 (O_494,N_9912,N_9954);
nor UO_495 (O_495,N_9839,N_9876);
and UO_496 (O_496,N_9888,N_9998);
nand UO_497 (O_497,N_9982,N_9871);
nand UO_498 (O_498,N_9843,N_9801);
xor UO_499 (O_499,N_9987,N_9999);
or UO_500 (O_500,N_9924,N_9902);
and UO_501 (O_501,N_9843,N_9827);
nor UO_502 (O_502,N_9927,N_9812);
nand UO_503 (O_503,N_9800,N_9850);
nand UO_504 (O_504,N_9973,N_9842);
or UO_505 (O_505,N_9997,N_9864);
and UO_506 (O_506,N_9875,N_9957);
and UO_507 (O_507,N_9925,N_9959);
and UO_508 (O_508,N_9942,N_9916);
xor UO_509 (O_509,N_9857,N_9829);
xor UO_510 (O_510,N_9811,N_9995);
nand UO_511 (O_511,N_9927,N_9939);
and UO_512 (O_512,N_9897,N_9988);
or UO_513 (O_513,N_9854,N_9879);
xnor UO_514 (O_514,N_9884,N_9979);
nand UO_515 (O_515,N_9930,N_9849);
and UO_516 (O_516,N_9922,N_9939);
or UO_517 (O_517,N_9819,N_9995);
or UO_518 (O_518,N_9809,N_9823);
or UO_519 (O_519,N_9874,N_9813);
or UO_520 (O_520,N_9979,N_9986);
or UO_521 (O_521,N_9845,N_9920);
and UO_522 (O_522,N_9977,N_9866);
nand UO_523 (O_523,N_9987,N_9808);
and UO_524 (O_524,N_9815,N_9936);
nor UO_525 (O_525,N_9872,N_9949);
and UO_526 (O_526,N_9806,N_9966);
xor UO_527 (O_527,N_9864,N_9852);
nor UO_528 (O_528,N_9851,N_9854);
nor UO_529 (O_529,N_9841,N_9842);
or UO_530 (O_530,N_9850,N_9979);
or UO_531 (O_531,N_9936,N_9874);
nand UO_532 (O_532,N_9864,N_9929);
nand UO_533 (O_533,N_9941,N_9852);
nor UO_534 (O_534,N_9950,N_9875);
and UO_535 (O_535,N_9810,N_9987);
xnor UO_536 (O_536,N_9829,N_9926);
or UO_537 (O_537,N_9853,N_9803);
xnor UO_538 (O_538,N_9956,N_9980);
nor UO_539 (O_539,N_9803,N_9821);
nand UO_540 (O_540,N_9952,N_9974);
xor UO_541 (O_541,N_9867,N_9803);
nor UO_542 (O_542,N_9956,N_9868);
and UO_543 (O_543,N_9831,N_9828);
xor UO_544 (O_544,N_9976,N_9868);
and UO_545 (O_545,N_9972,N_9951);
xor UO_546 (O_546,N_9999,N_9956);
and UO_547 (O_547,N_9982,N_9932);
xor UO_548 (O_548,N_9822,N_9826);
or UO_549 (O_549,N_9984,N_9958);
or UO_550 (O_550,N_9891,N_9934);
nor UO_551 (O_551,N_9863,N_9857);
nor UO_552 (O_552,N_9820,N_9971);
nand UO_553 (O_553,N_9920,N_9811);
nand UO_554 (O_554,N_9818,N_9833);
or UO_555 (O_555,N_9834,N_9807);
nor UO_556 (O_556,N_9966,N_9853);
or UO_557 (O_557,N_9904,N_9910);
or UO_558 (O_558,N_9860,N_9888);
nand UO_559 (O_559,N_9805,N_9904);
xor UO_560 (O_560,N_9809,N_9987);
or UO_561 (O_561,N_9807,N_9805);
nor UO_562 (O_562,N_9983,N_9813);
nor UO_563 (O_563,N_9895,N_9938);
xnor UO_564 (O_564,N_9902,N_9999);
nor UO_565 (O_565,N_9830,N_9801);
or UO_566 (O_566,N_9972,N_9877);
and UO_567 (O_567,N_9959,N_9864);
nor UO_568 (O_568,N_9898,N_9963);
or UO_569 (O_569,N_9943,N_9826);
or UO_570 (O_570,N_9860,N_9906);
nor UO_571 (O_571,N_9889,N_9823);
nor UO_572 (O_572,N_9979,N_9990);
nor UO_573 (O_573,N_9909,N_9837);
xnor UO_574 (O_574,N_9947,N_9844);
and UO_575 (O_575,N_9894,N_9823);
xor UO_576 (O_576,N_9951,N_9858);
and UO_577 (O_577,N_9841,N_9978);
nor UO_578 (O_578,N_9853,N_9884);
or UO_579 (O_579,N_9891,N_9968);
and UO_580 (O_580,N_9812,N_9983);
nor UO_581 (O_581,N_9857,N_9991);
nand UO_582 (O_582,N_9826,N_9882);
or UO_583 (O_583,N_9930,N_9836);
and UO_584 (O_584,N_9846,N_9917);
nand UO_585 (O_585,N_9865,N_9849);
nand UO_586 (O_586,N_9838,N_9855);
and UO_587 (O_587,N_9950,N_9851);
or UO_588 (O_588,N_9805,N_9813);
nand UO_589 (O_589,N_9911,N_9847);
nor UO_590 (O_590,N_9810,N_9864);
nor UO_591 (O_591,N_9998,N_9989);
nand UO_592 (O_592,N_9904,N_9882);
nand UO_593 (O_593,N_9886,N_9850);
or UO_594 (O_594,N_9902,N_9827);
xor UO_595 (O_595,N_9931,N_9924);
or UO_596 (O_596,N_9943,N_9959);
or UO_597 (O_597,N_9971,N_9976);
xnor UO_598 (O_598,N_9925,N_9857);
and UO_599 (O_599,N_9929,N_9827);
and UO_600 (O_600,N_9990,N_9876);
or UO_601 (O_601,N_9887,N_9861);
and UO_602 (O_602,N_9964,N_9985);
xor UO_603 (O_603,N_9827,N_9851);
or UO_604 (O_604,N_9936,N_9934);
and UO_605 (O_605,N_9970,N_9990);
xor UO_606 (O_606,N_9821,N_9892);
nor UO_607 (O_607,N_9931,N_9800);
xor UO_608 (O_608,N_9894,N_9864);
nand UO_609 (O_609,N_9941,N_9974);
or UO_610 (O_610,N_9994,N_9929);
and UO_611 (O_611,N_9967,N_9892);
xnor UO_612 (O_612,N_9976,N_9887);
and UO_613 (O_613,N_9943,N_9937);
nor UO_614 (O_614,N_9908,N_9945);
nor UO_615 (O_615,N_9983,N_9927);
and UO_616 (O_616,N_9973,N_9927);
xnor UO_617 (O_617,N_9811,N_9933);
xnor UO_618 (O_618,N_9998,N_9858);
and UO_619 (O_619,N_9938,N_9951);
xnor UO_620 (O_620,N_9824,N_9992);
or UO_621 (O_621,N_9956,N_9819);
or UO_622 (O_622,N_9910,N_9891);
nor UO_623 (O_623,N_9900,N_9973);
nand UO_624 (O_624,N_9895,N_9966);
and UO_625 (O_625,N_9947,N_9879);
nand UO_626 (O_626,N_9824,N_9820);
nor UO_627 (O_627,N_9938,N_9991);
nand UO_628 (O_628,N_9976,N_9845);
nand UO_629 (O_629,N_9955,N_9911);
nor UO_630 (O_630,N_9848,N_9897);
xnor UO_631 (O_631,N_9993,N_9828);
nor UO_632 (O_632,N_9866,N_9917);
or UO_633 (O_633,N_9945,N_9992);
nand UO_634 (O_634,N_9986,N_9818);
nor UO_635 (O_635,N_9858,N_9835);
xnor UO_636 (O_636,N_9812,N_9918);
or UO_637 (O_637,N_9976,N_9899);
or UO_638 (O_638,N_9892,N_9957);
xnor UO_639 (O_639,N_9912,N_9901);
xor UO_640 (O_640,N_9942,N_9918);
or UO_641 (O_641,N_9810,N_9955);
nor UO_642 (O_642,N_9954,N_9963);
nor UO_643 (O_643,N_9935,N_9867);
nand UO_644 (O_644,N_9992,N_9858);
and UO_645 (O_645,N_9984,N_9903);
and UO_646 (O_646,N_9992,N_9860);
or UO_647 (O_647,N_9800,N_9966);
nor UO_648 (O_648,N_9813,N_9812);
xnor UO_649 (O_649,N_9852,N_9861);
nor UO_650 (O_650,N_9934,N_9894);
and UO_651 (O_651,N_9922,N_9843);
nor UO_652 (O_652,N_9845,N_9890);
or UO_653 (O_653,N_9859,N_9869);
xor UO_654 (O_654,N_9889,N_9933);
xnor UO_655 (O_655,N_9815,N_9904);
xor UO_656 (O_656,N_9917,N_9830);
or UO_657 (O_657,N_9884,N_9913);
nor UO_658 (O_658,N_9804,N_9917);
or UO_659 (O_659,N_9944,N_9827);
xor UO_660 (O_660,N_9945,N_9981);
or UO_661 (O_661,N_9816,N_9927);
and UO_662 (O_662,N_9861,N_9899);
and UO_663 (O_663,N_9834,N_9804);
nor UO_664 (O_664,N_9928,N_9955);
xnor UO_665 (O_665,N_9923,N_9911);
nand UO_666 (O_666,N_9912,N_9835);
and UO_667 (O_667,N_9874,N_9907);
nand UO_668 (O_668,N_9996,N_9982);
or UO_669 (O_669,N_9860,N_9853);
nand UO_670 (O_670,N_9934,N_9943);
xnor UO_671 (O_671,N_9852,N_9895);
or UO_672 (O_672,N_9831,N_9817);
or UO_673 (O_673,N_9828,N_9973);
xor UO_674 (O_674,N_9945,N_9931);
or UO_675 (O_675,N_9800,N_9868);
and UO_676 (O_676,N_9809,N_9822);
or UO_677 (O_677,N_9802,N_9843);
xnor UO_678 (O_678,N_9829,N_9998);
nand UO_679 (O_679,N_9814,N_9833);
xor UO_680 (O_680,N_9885,N_9811);
nand UO_681 (O_681,N_9873,N_9920);
and UO_682 (O_682,N_9957,N_9871);
nand UO_683 (O_683,N_9895,N_9869);
nand UO_684 (O_684,N_9862,N_9984);
xor UO_685 (O_685,N_9877,N_9954);
nor UO_686 (O_686,N_9805,N_9958);
nor UO_687 (O_687,N_9935,N_9978);
nand UO_688 (O_688,N_9881,N_9972);
or UO_689 (O_689,N_9820,N_9909);
xnor UO_690 (O_690,N_9804,N_9986);
and UO_691 (O_691,N_9980,N_9850);
and UO_692 (O_692,N_9839,N_9851);
nor UO_693 (O_693,N_9857,N_9831);
and UO_694 (O_694,N_9979,N_9828);
nand UO_695 (O_695,N_9878,N_9923);
and UO_696 (O_696,N_9973,N_9802);
xnor UO_697 (O_697,N_9805,N_9917);
nor UO_698 (O_698,N_9898,N_9900);
or UO_699 (O_699,N_9878,N_9822);
nor UO_700 (O_700,N_9821,N_9863);
xor UO_701 (O_701,N_9815,N_9821);
xor UO_702 (O_702,N_9988,N_9814);
nand UO_703 (O_703,N_9843,N_9805);
nand UO_704 (O_704,N_9873,N_9923);
nand UO_705 (O_705,N_9811,N_9987);
and UO_706 (O_706,N_9908,N_9816);
xnor UO_707 (O_707,N_9879,N_9841);
nand UO_708 (O_708,N_9993,N_9977);
nand UO_709 (O_709,N_9811,N_9823);
xnor UO_710 (O_710,N_9955,N_9960);
nor UO_711 (O_711,N_9873,N_9993);
nor UO_712 (O_712,N_9936,N_9835);
xnor UO_713 (O_713,N_9948,N_9889);
xnor UO_714 (O_714,N_9968,N_9875);
nor UO_715 (O_715,N_9917,N_9847);
nand UO_716 (O_716,N_9889,N_9827);
and UO_717 (O_717,N_9984,N_9808);
and UO_718 (O_718,N_9928,N_9885);
nand UO_719 (O_719,N_9892,N_9944);
or UO_720 (O_720,N_9819,N_9978);
and UO_721 (O_721,N_9906,N_9837);
nand UO_722 (O_722,N_9870,N_9830);
or UO_723 (O_723,N_9921,N_9952);
or UO_724 (O_724,N_9852,N_9837);
nor UO_725 (O_725,N_9850,N_9935);
xnor UO_726 (O_726,N_9904,N_9880);
nand UO_727 (O_727,N_9840,N_9818);
nor UO_728 (O_728,N_9824,N_9868);
and UO_729 (O_729,N_9832,N_9928);
nand UO_730 (O_730,N_9985,N_9979);
nand UO_731 (O_731,N_9886,N_9896);
and UO_732 (O_732,N_9982,N_9844);
nor UO_733 (O_733,N_9935,N_9906);
xnor UO_734 (O_734,N_9998,N_9834);
nand UO_735 (O_735,N_9892,N_9940);
and UO_736 (O_736,N_9965,N_9825);
and UO_737 (O_737,N_9941,N_9975);
nand UO_738 (O_738,N_9927,N_9976);
xor UO_739 (O_739,N_9844,N_9985);
nand UO_740 (O_740,N_9939,N_9943);
xor UO_741 (O_741,N_9971,N_9838);
xnor UO_742 (O_742,N_9968,N_9922);
nor UO_743 (O_743,N_9874,N_9867);
nand UO_744 (O_744,N_9839,N_9826);
and UO_745 (O_745,N_9991,N_9920);
nor UO_746 (O_746,N_9944,N_9933);
or UO_747 (O_747,N_9980,N_9879);
or UO_748 (O_748,N_9864,N_9915);
xnor UO_749 (O_749,N_9967,N_9934);
nor UO_750 (O_750,N_9871,N_9922);
or UO_751 (O_751,N_9944,N_9843);
and UO_752 (O_752,N_9855,N_9865);
or UO_753 (O_753,N_9974,N_9904);
xnor UO_754 (O_754,N_9957,N_9984);
xnor UO_755 (O_755,N_9954,N_9802);
and UO_756 (O_756,N_9956,N_9822);
nand UO_757 (O_757,N_9831,N_9978);
or UO_758 (O_758,N_9819,N_9967);
nand UO_759 (O_759,N_9960,N_9918);
nor UO_760 (O_760,N_9850,N_9965);
nor UO_761 (O_761,N_9810,N_9946);
nand UO_762 (O_762,N_9807,N_9909);
or UO_763 (O_763,N_9905,N_9975);
nand UO_764 (O_764,N_9820,N_9945);
nor UO_765 (O_765,N_9808,N_9862);
xor UO_766 (O_766,N_9810,N_9902);
and UO_767 (O_767,N_9828,N_9950);
nor UO_768 (O_768,N_9822,N_9904);
nand UO_769 (O_769,N_9927,N_9982);
nor UO_770 (O_770,N_9858,N_9928);
or UO_771 (O_771,N_9869,N_9817);
nand UO_772 (O_772,N_9993,N_9956);
and UO_773 (O_773,N_9815,N_9890);
and UO_774 (O_774,N_9835,N_9915);
or UO_775 (O_775,N_9959,N_9971);
or UO_776 (O_776,N_9932,N_9943);
or UO_777 (O_777,N_9991,N_9849);
nand UO_778 (O_778,N_9988,N_9895);
xor UO_779 (O_779,N_9930,N_9900);
nor UO_780 (O_780,N_9935,N_9938);
xnor UO_781 (O_781,N_9876,N_9989);
xor UO_782 (O_782,N_9943,N_9833);
nor UO_783 (O_783,N_9867,N_9885);
and UO_784 (O_784,N_9942,N_9963);
nand UO_785 (O_785,N_9832,N_9878);
xnor UO_786 (O_786,N_9978,N_9821);
and UO_787 (O_787,N_9888,N_9992);
nand UO_788 (O_788,N_9812,N_9945);
or UO_789 (O_789,N_9983,N_9992);
nor UO_790 (O_790,N_9927,N_9857);
and UO_791 (O_791,N_9886,N_9876);
nor UO_792 (O_792,N_9824,N_9882);
nand UO_793 (O_793,N_9997,N_9974);
and UO_794 (O_794,N_9944,N_9837);
or UO_795 (O_795,N_9986,N_9816);
nor UO_796 (O_796,N_9883,N_9969);
xor UO_797 (O_797,N_9851,N_9834);
and UO_798 (O_798,N_9800,N_9805);
and UO_799 (O_799,N_9992,N_9901);
or UO_800 (O_800,N_9869,N_9819);
nand UO_801 (O_801,N_9829,N_9997);
or UO_802 (O_802,N_9867,N_9891);
xnor UO_803 (O_803,N_9874,N_9892);
nor UO_804 (O_804,N_9812,N_9944);
or UO_805 (O_805,N_9837,N_9815);
or UO_806 (O_806,N_9858,N_9988);
or UO_807 (O_807,N_9965,N_9898);
or UO_808 (O_808,N_9832,N_9888);
nor UO_809 (O_809,N_9847,N_9863);
xor UO_810 (O_810,N_9884,N_9901);
and UO_811 (O_811,N_9801,N_9803);
xor UO_812 (O_812,N_9810,N_9960);
and UO_813 (O_813,N_9856,N_9898);
and UO_814 (O_814,N_9889,N_9856);
or UO_815 (O_815,N_9829,N_9868);
nor UO_816 (O_816,N_9949,N_9915);
and UO_817 (O_817,N_9919,N_9956);
nand UO_818 (O_818,N_9972,N_9949);
nor UO_819 (O_819,N_9813,N_9922);
and UO_820 (O_820,N_9934,N_9826);
xnor UO_821 (O_821,N_9843,N_9904);
xor UO_822 (O_822,N_9839,N_9972);
and UO_823 (O_823,N_9840,N_9834);
nor UO_824 (O_824,N_9875,N_9949);
nor UO_825 (O_825,N_9807,N_9960);
nor UO_826 (O_826,N_9854,N_9815);
xnor UO_827 (O_827,N_9837,N_9922);
and UO_828 (O_828,N_9946,N_9899);
and UO_829 (O_829,N_9836,N_9811);
or UO_830 (O_830,N_9976,N_9834);
nor UO_831 (O_831,N_9822,N_9937);
nor UO_832 (O_832,N_9865,N_9800);
nand UO_833 (O_833,N_9980,N_9989);
and UO_834 (O_834,N_9805,N_9970);
or UO_835 (O_835,N_9992,N_9887);
nor UO_836 (O_836,N_9996,N_9941);
xnor UO_837 (O_837,N_9921,N_9819);
nor UO_838 (O_838,N_9964,N_9891);
xor UO_839 (O_839,N_9974,N_9994);
nand UO_840 (O_840,N_9886,N_9934);
nand UO_841 (O_841,N_9947,N_9881);
or UO_842 (O_842,N_9865,N_9825);
nand UO_843 (O_843,N_9840,N_9845);
and UO_844 (O_844,N_9923,N_9909);
or UO_845 (O_845,N_9995,N_9938);
nor UO_846 (O_846,N_9970,N_9827);
xnor UO_847 (O_847,N_9855,N_9856);
nor UO_848 (O_848,N_9821,N_9941);
nor UO_849 (O_849,N_9911,N_9812);
and UO_850 (O_850,N_9839,N_9829);
or UO_851 (O_851,N_9859,N_9935);
xor UO_852 (O_852,N_9841,N_9890);
and UO_853 (O_853,N_9983,N_9909);
xnor UO_854 (O_854,N_9811,N_9805);
xnor UO_855 (O_855,N_9824,N_9947);
or UO_856 (O_856,N_9995,N_9893);
nand UO_857 (O_857,N_9960,N_9871);
nand UO_858 (O_858,N_9941,N_9823);
nor UO_859 (O_859,N_9976,N_9821);
or UO_860 (O_860,N_9808,N_9980);
and UO_861 (O_861,N_9869,N_9905);
xnor UO_862 (O_862,N_9955,N_9820);
xnor UO_863 (O_863,N_9972,N_9925);
and UO_864 (O_864,N_9964,N_9863);
xnor UO_865 (O_865,N_9916,N_9933);
xor UO_866 (O_866,N_9834,N_9910);
nor UO_867 (O_867,N_9815,N_9842);
nor UO_868 (O_868,N_9892,N_9878);
and UO_869 (O_869,N_9884,N_9972);
or UO_870 (O_870,N_9815,N_9874);
xnor UO_871 (O_871,N_9994,N_9949);
nor UO_872 (O_872,N_9833,N_9806);
or UO_873 (O_873,N_9885,N_9816);
nor UO_874 (O_874,N_9832,N_9963);
and UO_875 (O_875,N_9877,N_9920);
xor UO_876 (O_876,N_9861,N_9827);
and UO_877 (O_877,N_9923,N_9900);
xor UO_878 (O_878,N_9965,N_9888);
or UO_879 (O_879,N_9800,N_9861);
or UO_880 (O_880,N_9942,N_9962);
or UO_881 (O_881,N_9950,N_9835);
and UO_882 (O_882,N_9998,N_9852);
nor UO_883 (O_883,N_9973,N_9800);
and UO_884 (O_884,N_9980,N_9890);
xor UO_885 (O_885,N_9926,N_9982);
and UO_886 (O_886,N_9885,N_9924);
xnor UO_887 (O_887,N_9800,N_9804);
or UO_888 (O_888,N_9851,N_9858);
or UO_889 (O_889,N_9835,N_9991);
nor UO_890 (O_890,N_9983,N_9826);
xnor UO_891 (O_891,N_9882,N_9867);
or UO_892 (O_892,N_9830,N_9853);
or UO_893 (O_893,N_9854,N_9959);
xnor UO_894 (O_894,N_9826,N_9850);
xor UO_895 (O_895,N_9872,N_9857);
xnor UO_896 (O_896,N_9977,N_9932);
xor UO_897 (O_897,N_9975,N_9945);
or UO_898 (O_898,N_9827,N_9963);
nor UO_899 (O_899,N_9978,N_9851);
or UO_900 (O_900,N_9844,N_9980);
and UO_901 (O_901,N_9988,N_9830);
and UO_902 (O_902,N_9881,N_9921);
xnor UO_903 (O_903,N_9947,N_9892);
and UO_904 (O_904,N_9844,N_9857);
nand UO_905 (O_905,N_9871,N_9971);
nor UO_906 (O_906,N_9879,N_9909);
xor UO_907 (O_907,N_9955,N_9898);
nor UO_908 (O_908,N_9962,N_9834);
nor UO_909 (O_909,N_9826,N_9831);
and UO_910 (O_910,N_9865,N_9974);
and UO_911 (O_911,N_9809,N_9923);
or UO_912 (O_912,N_9897,N_9894);
nor UO_913 (O_913,N_9909,N_9951);
xnor UO_914 (O_914,N_9949,N_9923);
nand UO_915 (O_915,N_9819,N_9861);
nor UO_916 (O_916,N_9945,N_9828);
xor UO_917 (O_917,N_9871,N_9900);
nor UO_918 (O_918,N_9942,N_9997);
nand UO_919 (O_919,N_9837,N_9910);
xor UO_920 (O_920,N_9894,N_9997);
nand UO_921 (O_921,N_9936,N_9943);
nor UO_922 (O_922,N_9959,N_9900);
nand UO_923 (O_923,N_9850,N_9978);
nand UO_924 (O_924,N_9936,N_9877);
nor UO_925 (O_925,N_9821,N_9874);
xnor UO_926 (O_926,N_9846,N_9998);
and UO_927 (O_927,N_9965,N_9979);
xor UO_928 (O_928,N_9955,N_9982);
or UO_929 (O_929,N_9815,N_9846);
nor UO_930 (O_930,N_9979,N_9849);
nor UO_931 (O_931,N_9877,N_9960);
nor UO_932 (O_932,N_9967,N_9827);
nand UO_933 (O_933,N_9831,N_9910);
nand UO_934 (O_934,N_9962,N_9911);
nor UO_935 (O_935,N_9958,N_9995);
nand UO_936 (O_936,N_9824,N_9978);
nand UO_937 (O_937,N_9913,N_9956);
or UO_938 (O_938,N_9912,N_9922);
or UO_939 (O_939,N_9810,N_9954);
nand UO_940 (O_940,N_9975,N_9818);
nor UO_941 (O_941,N_9836,N_9952);
and UO_942 (O_942,N_9868,N_9863);
nor UO_943 (O_943,N_9901,N_9816);
nand UO_944 (O_944,N_9996,N_9995);
xnor UO_945 (O_945,N_9830,N_9800);
or UO_946 (O_946,N_9850,N_9977);
and UO_947 (O_947,N_9896,N_9902);
and UO_948 (O_948,N_9946,N_9862);
xor UO_949 (O_949,N_9864,N_9887);
or UO_950 (O_950,N_9962,N_9900);
and UO_951 (O_951,N_9913,N_9871);
xor UO_952 (O_952,N_9828,N_9929);
or UO_953 (O_953,N_9880,N_9840);
nand UO_954 (O_954,N_9948,N_9988);
or UO_955 (O_955,N_9981,N_9837);
and UO_956 (O_956,N_9921,N_9937);
nor UO_957 (O_957,N_9983,N_9824);
and UO_958 (O_958,N_9869,N_9984);
nor UO_959 (O_959,N_9965,N_9856);
or UO_960 (O_960,N_9978,N_9839);
nor UO_961 (O_961,N_9871,N_9861);
nor UO_962 (O_962,N_9939,N_9813);
nor UO_963 (O_963,N_9858,N_9881);
or UO_964 (O_964,N_9980,N_9983);
xor UO_965 (O_965,N_9920,N_9870);
xor UO_966 (O_966,N_9867,N_9826);
and UO_967 (O_967,N_9987,N_9955);
nor UO_968 (O_968,N_9903,N_9933);
or UO_969 (O_969,N_9964,N_9845);
and UO_970 (O_970,N_9811,N_9821);
or UO_971 (O_971,N_9847,N_9944);
nor UO_972 (O_972,N_9925,N_9953);
or UO_973 (O_973,N_9822,N_9953);
xnor UO_974 (O_974,N_9810,N_9972);
and UO_975 (O_975,N_9877,N_9970);
or UO_976 (O_976,N_9826,N_9975);
xor UO_977 (O_977,N_9963,N_9950);
xor UO_978 (O_978,N_9892,N_9971);
xor UO_979 (O_979,N_9833,N_9849);
and UO_980 (O_980,N_9931,N_9934);
or UO_981 (O_981,N_9974,N_9817);
or UO_982 (O_982,N_9868,N_9944);
xor UO_983 (O_983,N_9853,N_9859);
xor UO_984 (O_984,N_9906,N_9989);
and UO_985 (O_985,N_9817,N_9810);
nor UO_986 (O_986,N_9955,N_9927);
nand UO_987 (O_987,N_9966,N_9838);
xnor UO_988 (O_988,N_9920,N_9862);
nor UO_989 (O_989,N_9814,N_9851);
or UO_990 (O_990,N_9904,N_9930);
or UO_991 (O_991,N_9822,N_9831);
nand UO_992 (O_992,N_9876,N_9985);
or UO_993 (O_993,N_9831,N_9816);
xnor UO_994 (O_994,N_9981,N_9842);
nor UO_995 (O_995,N_9915,N_9928);
and UO_996 (O_996,N_9814,N_9839);
nor UO_997 (O_997,N_9837,N_9845);
nor UO_998 (O_998,N_9863,N_9897);
xor UO_999 (O_999,N_9963,N_9927);
nand UO_1000 (O_1000,N_9847,N_9834);
nor UO_1001 (O_1001,N_9957,N_9940);
and UO_1002 (O_1002,N_9858,N_9960);
and UO_1003 (O_1003,N_9882,N_9917);
xor UO_1004 (O_1004,N_9863,N_9829);
or UO_1005 (O_1005,N_9823,N_9862);
xnor UO_1006 (O_1006,N_9910,N_9842);
nor UO_1007 (O_1007,N_9804,N_9983);
or UO_1008 (O_1008,N_9954,N_9845);
nor UO_1009 (O_1009,N_9982,N_9952);
and UO_1010 (O_1010,N_9949,N_9855);
and UO_1011 (O_1011,N_9952,N_9833);
nor UO_1012 (O_1012,N_9976,N_9980);
nor UO_1013 (O_1013,N_9829,N_9840);
xnor UO_1014 (O_1014,N_9901,N_9970);
xor UO_1015 (O_1015,N_9890,N_9901);
nor UO_1016 (O_1016,N_9885,N_9881);
or UO_1017 (O_1017,N_9959,N_9985);
nor UO_1018 (O_1018,N_9894,N_9857);
or UO_1019 (O_1019,N_9813,N_9992);
xnor UO_1020 (O_1020,N_9852,N_9818);
nor UO_1021 (O_1021,N_9815,N_9822);
nor UO_1022 (O_1022,N_9917,N_9863);
xor UO_1023 (O_1023,N_9984,N_9998);
xor UO_1024 (O_1024,N_9865,N_9816);
and UO_1025 (O_1025,N_9901,N_9887);
or UO_1026 (O_1026,N_9864,N_9931);
nor UO_1027 (O_1027,N_9838,N_9925);
nor UO_1028 (O_1028,N_9939,N_9877);
xnor UO_1029 (O_1029,N_9963,N_9825);
xor UO_1030 (O_1030,N_9902,N_9872);
nand UO_1031 (O_1031,N_9809,N_9885);
nor UO_1032 (O_1032,N_9893,N_9840);
xor UO_1033 (O_1033,N_9988,N_9822);
nor UO_1034 (O_1034,N_9940,N_9882);
and UO_1035 (O_1035,N_9997,N_9989);
nor UO_1036 (O_1036,N_9854,N_9867);
nor UO_1037 (O_1037,N_9957,N_9830);
and UO_1038 (O_1038,N_9991,N_9919);
nor UO_1039 (O_1039,N_9824,N_9910);
and UO_1040 (O_1040,N_9827,N_9803);
xor UO_1041 (O_1041,N_9979,N_9904);
nor UO_1042 (O_1042,N_9853,N_9948);
xor UO_1043 (O_1043,N_9897,N_9957);
or UO_1044 (O_1044,N_9884,N_9828);
xnor UO_1045 (O_1045,N_9939,N_9885);
xnor UO_1046 (O_1046,N_9932,N_9808);
xor UO_1047 (O_1047,N_9948,N_9970);
xor UO_1048 (O_1048,N_9960,N_9881);
xnor UO_1049 (O_1049,N_9921,N_9823);
xnor UO_1050 (O_1050,N_9833,N_9857);
or UO_1051 (O_1051,N_9870,N_9896);
nor UO_1052 (O_1052,N_9958,N_9876);
xnor UO_1053 (O_1053,N_9939,N_9833);
xor UO_1054 (O_1054,N_9982,N_9913);
and UO_1055 (O_1055,N_9879,N_9843);
or UO_1056 (O_1056,N_9993,N_9930);
nand UO_1057 (O_1057,N_9820,N_9948);
xnor UO_1058 (O_1058,N_9945,N_9985);
and UO_1059 (O_1059,N_9906,N_9926);
or UO_1060 (O_1060,N_9935,N_9942);
xnor UO_1061 (O_1061,N_9803,N_9986);
and UO_1062 (O_1062,N_9812,N_9878);
and UO_1063 (O_1063,N_9850,N_9961);
nor UO_1064 (O_1064,N_9861,N_9971);
nor UO_1065 (O_1065,N_9944,N_9815);
nand UO_1066 (O_1066,N_9941,N_9859);
and UO_1067 (O_1067,N_9991,N_9992);
or UO_1068 (O_1068,N_9986,N_9908);
or UO_1069 (O_1069,N_9926,N_9884);
xnor UO_1070 (O_1070,N_9937,N_9869);
xnor UO_1071 (O_1071,N_9937,N_9984);
nand UO_1072 (O_1072,N_9922,N_9989);
nand UO_1073 (O_1073,N_9862,N_9932);
xor UO_1074 (O_1074,N_9932,N_9965);
and UO_1075 (O_1075,N_9969,N_9965);
nor UO_1076 (O_1076,N_9977,N_9812);
nand UO_1077 (O_1077,N_9912,N_9991);
nor UO_1078 (O_1078,N_9839,N_9952);
nand UO_1079 (O_1079,N_9829,N_9909);
nor UO_1080 (O_1080,N_9882,N_9800);
xor UO_1081 (O_1081,N_9826,N_9965);
and UO_1082 (O_1082,N_9991,N_9852);
and UO_1083 (O_1083,N_9965,N_9966);
nor UO_1084 (O_1084,N_9868,N_9856);
and UO_1085 (O_1085,N_9942,N_9839);
nor UO_1086 (O_1086,N_9907,N_9911);
or UO_1087 (O_1087,N_9990,N_9825);
and UO_1088 (O_1088,N_9879,N_9894);
nor UO_1089 (O_1089,N_9866,N_9875);
nand UO_1090 (O_1090,N_9887,N_9808);
xnor UO_1091 (O_1091,N_9883,N_9994);
nand UO_1092 (O_1092,N_9839,N_9929);
or UO_1093 (O_1093,N_9940,N_9846);
or UO_1094 (O_1094,N_9933,N_9948);
and UO_1095 (O_1095,N_9900,N_9820);
or UO_1096 (O_1096,N_9901,N_9927);
or UO_1097 (O_1097,N_9851,N_9933);
and UO_1098 (O_1098,N_9926,N_9815);
or UO_1099 (O_1099,N_9967,N_9994);
or UO_1100 (O_1100,N_9800,N_9808);
xor UO_1101 (O_1101,N_9962,N_9826);
nand UO_1102 (O_1102,N_9833,N_9839);
xor UO_1103 (O_1103,N_9862,N_9980);
nand UO_1104 (O_1104,N_9872,N_9882);
or UO_1105 (O_1105,N_9927,N_9993);
or UO_1106 (O_1106,N_9888,N_9829);
nor UO_1107 (O_1107,N_9959,N_9806);
nor UO_1108 (O_1108,N_9819,N_9901);
xnor UO_1109 (O_1109,N_9898,N_9867);
or UO_1110 (O_1110,N_9916,N_9860);
nor UO_1111 (O_1111,N_9952,N_9868);
xor UO_1112 (O_1112,N_9941,N_9825);
or UO_1113 (O_1113,N_9837,N_9802);
and UO_1114 (O_1114,N_9964,N_9970);
nand UO_1115 (O_1115,N_9853,N_9976);
or UO_1116 (O_1116,N_9848,N_9960);
nor UO_1117 (O_1117,N_9927,N_9806);
or UO_1118 (O_1118,N_9820,N_9805);
and UO_1119 (O_1119,N_9802,N_9823);
or UO_1120 (O_1120,N_9817,N_9877);
xor UO_1121 (O_1121,N_9886,N_9825);
nand UO_1122 (O_1122,N_9907,N_9992);
nor UO_1123 (O_1123,N_9802,N_9835);
nor UO_1124 (O_1124,N_9968,N_9984);
and UO_1125 (O_1125,N_9861,N_9915);
nor UO_1126 (O_1126,N_9924,N_9886);
and UO_1127 (O_1127,N_9834,N_9845);
xnor UO_1128 (O_1128,N_9865,N_9845);
or UO_1129 (O_1129,N_9952,N_9966);
or UO_1130 (O_1130,N_9945,N_9939);
nor UO_1131 (O_1131,N_9915,N_9892);
nor UO_1132 (O_1132,N_9903,N_9800);
or UO_1133 (O_1133,N_9814,N_9846);
or UO_1134 (O_1134,N_9884,N_9994);
or UO_1135 (O_1135,N_9955,N_9962);
nor UO_1136 (O_1136,N_9982,N_9861);
nand UO_1137 (O_1137,N_9902,N_9964);
and UO_1138 (O_1138,N_9860,N_9995);
or UO_1139 (O_1139,N_9952,N_9864);
xnor UO_1140 (O_1140,N_9812,N_9981);
nand UO_1141 (O_1141,N_9806,N_9983);
and UO_1142 (O_1142,N_9988,N_9851);
nor UO_1143 (O_1143,N_9951,N_9925);
and UO_1144 (O_1144,N_9993,N_9940);
and UO_1145 (O_1145,N_9916,N_9848);
nand UO_1146 (O_1146,N_9934,N_9800);
xor UO_1147 (O_1147,N_9876,N_9851);
or UO_1148 (O_1148,N_9832,N_9855);
xnor UO_1149 (O_1149,N_9845,N_9861);
and UO_1150 (O_1150,N_9957,N_9965);
nor UO_1151 (O_1151,N_9896,N_9881);
nor UO_1152 (O_1152,N_9980,N_9971);
nor UO_1153 (O_1153,N_9982,N_9877);
nor UO_1154 (O_1154,N_9924,N_9909);
and UO_1155 (O_1155,N_9836,N_9846);
xnor UO_1156 (O_1156,N_9834,N_9892);
xnor UO_1157 (O_1157,N_9933,N_9961);
nand UO_1158 (O_1158,N_9963,N_9806);
xor UO_1159 (O_1159,N_9828,N_9913);
nor UO_1160 (O_1160,N_9915,N_9969);
and UO_1161 (O_1161,N_9856,N_9905);
nor UO_1162 (O_1162,N_9897,N_9986);
or UO_1163 (O_1163,N_9984,N_9946);
xnor UO_1164 (O_1164,N_9829,N_9965);
or UO_1165 (O_1165,N_9837,N_9952);
nor UO_1166 (O_1166,N_9926,N_9949);
xor UO_1167 (O_1167,N_9861,N_9942);
nand UO_1168 (O_1168,N_9839,N_9878);
nor UO_1169 (O_1169,N_9971,N_9822);
xnor UO_1170 (O_1170,N_9865,N_9883);
nor UO_1171 (O_1171,N_9823,N_9829);
nand UO_1172 (O_1172,N_9848,N_9907);
nand UO_1173 (O_1173,N_9979,N_9951);
nor UO_1174 (O_1174,N_9807,N_9932);
and UO_1175 (O_1175,N_9960,N_9927);
or UO_1176 (O_1176,N_9987,N_9969);
nand UO_1177 (O_1177,N_9918,N_9881);
nand UO_1178 (O_1178,N_9948,N_9931);
and UO_1179 (O_1179,N_9935,N_9963);
and UO_1180 (O_1180,N_9887,N_9957);
nand UO_1181 (O_1181,N_9940,N_9943);
or UO_1182 (O_1182,N_9974,N_9888);
nand UO_1183 (O_1183,N_9891,N_9959);
and UO_1184 (O_1184,N_9884,N_9875);
nand UO_1185 (O_1185,N_9895,N_9849);
xnor UO_1186 (O_1186,N_9976,N_9923);
xnor UO_1187 (O_1187,N_9955,N_9926);
xor UO_1188 (O_1188,N_9907,N_9990);
xor UO_1189 (O_1189,N_9895,N_9836);
xor UO_1190 (O_1190,N_9953,N_9944);
nand UO_1191 (O_1191,N_9821,N_9956);
xor UO_1192 (O_1192,N_9880,N_9822);
or UO_1193 (O_1193,N_9822,N_9928);
nor UO_1194 (O_1194,N_9847,N_9875);
or UO_1195 (O_1195,N_9991,N_9930);
nand UO_1196 (O_1196,N_9877,N_9989);
nand UO_1197 (O_1197,N_9923,N_9951);
xor UO_1198 (O_1198,N_9840,N_9987);
or UO_1199 (O_1199,N_9842,N_9889);
nand UO_1200 (O_1200,N_9983,N_9856);
nor UO_1201 (O_1201,N_9984,N_9836);
nand UO_1202 (O_1202,N_9853,N_9817);
xnor UO_1203 (O_1203,N_9855,N_9972);
nand UO_1204 (O_1204,N_9969,N_9974);
xnor UO_1205 (O_1205,N_9819,N_9954);
xor UO_1206 (O_1206,N_9987,N_9874);
nor UO_1207 (O_1207,N_9935,N_9997);
nand UO_1208 (O_1208,N_9977,N_9898);
nor UO_1209 (O_1209,N_9902,N_9850);
nor UO_1210 (O_1210,N_9889,N_9909);
nor UO_1211 (O_1211,N_9855,N_9952);
nor UO_1212 (O_1212,N_9959,N_9916);
and UO_1213 (O_1213,N_9965,N_9967);
nand UO_1214 (O_1214,N_9887,N_9989);
or UO_1215 (O_1215,N_9915,N_9983);
nor UO_1216 (O_1216,N_9841,N_9836);
or UO_1217 (O_1217,N_9911,N_9965);
and UO_1218 (O_1218,N_9832,N_9892);
nor UO_1219 (O_1219,N_9877,N_9854);
and UO_1220 (O_1220,N_9944,N_9813);
nand UO_1221 (O_1221,N_9815,N_9953);
and UO_1222 (O_1222,N_9887,N_9872);
or UO_1223 (O_1223,N_9898,N_9815);
or UO_1224 (O_1224,N_9859,N_9874);
or UO_1225 (O_1225,N_9839,N_9842);
and UO_1226 (O_1226,N_9988,N_9944);
and UO_1227 (O_1227,N_9952,N_9819);
and UO_1228 (O_1228,N_9928,N_9923);
and UO_1229 (O_1229,N_9967,N_9899);
and UO_1230 (O_1230,N_9806,N_9907);
nor UO_1231 (O_1231,N_9871,N_9818);
and UO_1232 (O_1232,N_9944,N_9889);
nand UO_1233 (O_1233,N_9967,N_9915);
nand UO_1234 (O_1234,N_9970,N_9821);
xnor UO_1235 (O_1235,N_9931,N_9903);
or UO_1236 (O_1236,N_9963,N_9802);
and UO_1237 (O_1237,N_9854,N_9888);
nand UO_1238 (O_1238,N_9815,N_9839);
nand UO_1239 (O_1239,N_9883,N_9907);
xnor UO_1240 (O_1240,N_9959,N_9998);
and UO_1241 (O_1241,N_9823,N_9997);
or UO_1242 (O_1242,N_9910,N_9821);
xnor UO_1243 (O_1243,N_9975,N_9802);
nand UO_1244 (O_1244,N_9802,N_9913);
xnor UO_1245 (O_1245,N_9817,N_9932);
nor UO_1246 (O_1246,N_9954,N_9863);
or UO_1247 (O_1247,N_9877,N_9927);
xnor UO_1248 (O_1248,N_9834,N_9936);
nand UO_1249 (O_1249,N_9970,N_9958);
nor UO_1250 (O_1250,N_9984,N_9840);
and UO_1251 (O_1251,N_9992,N_9820);
or UO_1252 (O_1252,N_9879,N_9940);
nand UO_1253 (O_1253,N_9883,N_9821);
nor UO_1254 (O_1254,N_9965,N_9867);
and UO_1255 (O_1255,N_9842,N_9894);
xor UO_1256 (O_1256,N_9819,N_9868);
nand UO_1257 (O_1257,N_9833,N_9836);
nand UO_1258 (O_1258,N_9872,N_9936);
nand UO_1259 (O_1259,N_9912,N_9997);
nor UO_1260 (O_1260,N_9851,N_9856);
xnor UO_1261 (O_1261,N_9819,N_9865);
and UO_1262 (O_1262,N_9886,N_9897);
nor UO_1263 (O_1263,N_9829,N_9973);
nand UO_1264 (O_1264,N_9905,N_9817);
or UO_1265 (O_1265,N_9876,N_9942);
nand UO_1266 (O_1266,N_9972,N_9963);
nor UO_1267 (O_1267,N_9852,N_9985);
xor UO_1268 (O_1268,N_9978,N_9956);
nor UO_1269 (O_1269,N_9843,N_9978);
nor UO_1270 (O_1270,N_9825,N_9804);
nor UO_1271 (O_1271,N_9942,N_9830);
or UO_1272 (O_1272,N_9993,N_9823);
xor UO_1273 (O_1273,N_9887,N_9983);
nand UO_1274 (O_1274,N_9862,N_9811);
nand UO_1275 (O_1275,N_9842,N_9927);
and UO_1276 (O_1276,N_9949,N_9985);
nand UO_1277 (O_1277,N_9962,N_9980);
nand UO_1278 (O_1278,N_9803,N_9901);
nand UO_1279 (O_1279,N_9952,N_9825);
and UO_1280 (O_1280,N_9941,N_9898);
and UO_1281 (O_1281,N_9814,N_9860);
xnor UO_1282 (O_1282,N_9873,N_9922);
nand UO_1283 (O_1283,N_9800,N_9819);
or UO_1284 (O_1284,N_9927,N_9954);
xnor UO_1285 (O_1285,N_9802,N_9939);
or UO_1286 (O_1286,N_9991,N_9975);
or UO_1287 (O_1287,N_9909,N_9987);
nor UO_1288 (O_1288,N_9854,N_9917);
xnor UO_1289 (O_1289,N_9971,N_9909);
or UO_1290 (O_1290,N_9911,N_9890);
and UO_1291 (O_1291,N_9933,N_9972);
or UO_1292 (O_1292,N_9871,N_9996);
or UO_1293 (O_1293,N_9996,N_9998);
nor UO_1294 (O_1294,N_9943,N_9806);
and UO_1295 (O_1295,N_9909,N_9846);
nand UO_1296 (O_1296,N_9815,N_9921);
nand UO_1297 (O_1297,N_9882,N_9950);
nand UO_1298 (O_1298,N_9803,N_9862);
nor UO_1299 (O_1299,N_9914,N_9848);
nand UO_1300 (O_1300,N_9815,N_9915);
xnor UO_1301 (O_1301,N_9887,N_9814);
nor UO_1302 (O_1302,N_9989,N_9986);
nand UO_1303 (O_1303,N_9809,N_9956);
or UO_1304 (O_1304,N_9849,N_9884);
xnor UO_1305 (O_1305,N_9993,N_9943);
or UO_1306 (O_1306,N_9839,N_9973);
or UO_1307 (O_1307,N_9995,N_9921);
and UO_1308 (O_1308,N_9974,N_9988);
or UO_1309 (O_1309,N_9900,N_9977);
nor UO_1310 (O_1310,N_9935,N_9879);
nand UO_1311 (O_1311,N_9848,N_9812);
xor UO_1312 (O_1312,N_9954,N_9844);
nor UO_1313 (O_1313,N_9827,N_9813);
and UO_1314 (O_1314,N_9869,N_9856);
xor UO_1315 (O_1315,N_9834,N_9982);
nor UO_1316 (O_1316,N_9953,N_9843);
xnor UO_1317 (O_1317,N_9875,N_9931);
and UO_1318 (O_1318,N_9803,N_9883);
or UO_1319 (O_1319,N_9993,N_9854);
nor UO_1320 (O_1320,N_9877,N_9884);
or UO_1321 (O_1321,N_9911,N_9915);
xor UO_1322 (O_1322,N_9847,N_9953);
xor UO_1323 (O_1323,N_9973,N_9997);
nand UO_1324 (O_1324,N_9918,N_9818);
xnor UO_1325 (O_1325,N_9891,N_9914);
and UO_1326 (O_1326,N_9887,N_9817);
xor UO_1327 (O_1327,N_9883,N_9810);
or UO_1328 (O_1328,N_9992,N_9923);
and UO_1329 (O_1329,N_9858,N_9885);
and UO_1330 (O_1330,N_9845,N_9826);
nor UO_1331 (O_1331,N_9819,N_9919);
or UO_1332 (O_1332,N_9992,N_9948);
xnor UO_1333 (O_1333,N_9838,N_9865);
or UO_1334 (O_1334,N_9837,N_9936);
and UO_1335 (O_1335,N_9916,N_9910);
xnor UO_1336 (O_1336,N_9907,N_9903);
nor UO_1337 (O_1337,N_9983,N_9855);
nor UO_1338 (O_1338,N_9884,N_9991);
nand UO_1339 (O_1339,N_9957,N_9898);
and UO_1340 (O_1340,N_9960,N_9894);
xnor UO_1341 (O_1341,N_9849,N_9971);
nor UO_1342 (O_1342,N_9978,N_9979);
xor UO_1343 (O_1343,N_9941,N_9906);
xor UO_1344 (O_1344,N_9847,N_9868);
nor UO_1345 (O_1345,N_9812,N_9805);
nor UO_1346 (O_1346,N_9848,N_9880);
and UO_1347 (O_1347,N_9923,N_9993);
and UO_1348 (O_1348,N_9851,N_9900);
and UO_1349 (O_1349,N_9956,N_9870);
nand UO_1350 (O_1350,N_9821,N_9875);
or UO_1351 (O_1351,N_9969,N_9941);
or UO_1352 (O_1352,N_9881,N_9963);
nand UO_1353 (O_1353,N_9809,N_9815);
or UO_1354 (O_1354,N_9869,N_9804);
nor UO_1355 (O_1355,N_9857,N_9956);
xnor UO_1356 (O_1356,N_9880,N_9836);
xor UO_1357 (O_1357,N_9847,N_9840);
nand UO_1358 (O_1358,N_9829,N_9981);
or UO_1359 (O_1359,N_9956,N_9925);
nand UO_1360 (O_1360,N_9933,N_9896);
nand UO_1361 (O_1361,N_9890,N_9971);
or UO_1362 (O_1362,N_9828,N_9808);
and UO_1363 (O_1363,N_9916,N_9802);
nand UO_1364 (O_1364,N_9953,N_9948);
xnor UO_1365 (O_1365,N_9859,N_9962);
or UO_1366 (O_1366,N_9986,N_9844);
and UO_1367 (O_1367,N_9982,N_9978);
and UO_1368 (O_1368,N_9976,N_9989);
and UO_1369 (O_1369,N_9972,N_9918);
nor UO_1370 (O_1370,N_9822,N_9865);
or UO_1371 (O_1371,N_9907,N_9825);
xnor UO_1372 (O_1372,N_9984,N_9848);
nand UO_1373 (O_1373,N_9845,N_9839);
or UO_1374 (O_1374,N_9932,N_9963);
nor UO_1375 (O_1375,N_9966,N_9995);
nor UO_1376 (O_1376,N_9879,N_9888);
and UO_1377 (O_1377,N_9887,N_9824);
or UO_1378 (O_1378,N_9827,N_9888);
or UO_1379 (O_1379,N_9844,N_9945);
and UO_1380 (O_1380,N_9871,N_9986);
xnor UO_1381 (O_1381,N_9877,N_9869);
and UO_1382 (O_1382,N_9866,N_9883);
or UO_1383 (O_1383,N_9976,N_9935);
or UO_1384 (O_1384,N_9990,N_9800);
nand UO_1385 (O_1385,N_9830,N_9959);
xor UO_1386 (O_1386,N_9807,N_9906);
and UO_1387 (O_1387,N_9924,N_9899);
nor UO_1388 (O_1388,N_9925,N_9955);
or UO_1389 (O_1389,N_9997,N_9868);
and UO_1390 (O_1390,N_9842,N_9904);
nand UO_1391 (O_1391,N_9809,N_9854);
nand UO_1392 (O_1392,N_9990,N_9806);
and UO_1393 (O_1393,N_9846,N_9997);
or UO_1394 (O_1394,N_9807,N_9812);
and UO_1395 (O_1395,N_9914,N_9827);
nand UO_1396 (O_1396,N_9816,N_9871);
and UO_1397 (O_1397,N_9916,N_9937);
nor UO_1398 (O_1398,N_9889,N_9939);
or UO_1399 (O_1399,N_9878,N_9925);
nor UO_1400 (O_1400,N_9938,N_9812);
or UO_1401 (O_1401,N_9936,N_9930);
or UO_1402 (O_1402,N_9802,N_9964);
and UO_1403 (O_1403,N_9846,N_9837);
or UO_1404 (O_1404,N_9931,N_9851);
or UO_1405 (O_1405,N_9878,N_9931);
nor UO_1406 (O_1406,N_9869,N_9929);
or UO_1407 (O_1407,N_9834,N_9889);
nor UO_1408 (O_1408,N_9986,N_9899);
nor UO_1409 (O_1409,N_9971,N_9880);
nor UO_1410 (O_1410,N_9940,N_9998);
xor UO_1411 (O_1411,N_9861,N_9825);
or UO_1412 (O_1412,N_9964,N_9903);
nand UO_1413 (O_1413,N_9909,N_9996);
nand UO_1414 (O_1414,N_9874,N_9971);
xnor UO_1415 (O_1415,N_9827,N_9826);
or UO_1416 (O_1416,N_9949,N_9896);
or UO_1417 (O_1417,N_9877,N_9998);
nor UO_1418 (O_1418,N_9996,N_9938);
nand UO_1419 (O_1419,N_9980,N_9863);
or UO_1420 (O_1420,N_9939,N_9801);
nor UO_1421 (O_1421,N_9983,N_9995);
and UO_1422 (O_1422,N_9901,N_9929);
or UO_1423 (O_1423,N_9977,N_9984);
nor UO_1424 (O_1424,N_9992,N_9962);
xnor UO_1425 (O_1425,N_9968,N_9829);
nand UO_1426 (O_1426,N_9970,N_9866);
xor UO_1427 (O_1427,N_9814,N_9868);
nand UO_1428 (O_1428,N_9916,N_9868);
or UO_1429 (O_1429,N_9906,N_9839);
nor UO_1430 (O_1430,N_9800,N_9972);
or UO_1431 (O_1431,N_9963,N_9965);
nand UO_1432 (O_1432,N_9928,N_9936);
nor UO_1433 (O_1433,N_9853,N_9805);
and UO_1434 (O_1434,N_9817,N_9960);
nand UO_1435 (O_1435,N_9880,N_9919);
nand UO_1436 (O_1436,N_9998,N_9925);
nor UO_1437 (O_1437,N_9967,N_9851);
nor UO_1438 (O_1438,N_9875,N_9806);
nor UO_1439 (O_1439,N_9832,N_9929);
nand UO_1440 (O_1440,N_9963,N_9860);
nor UO_1441 (O_1441,N_9971,N_9846);
nand UO_1442 (O_1442,N_9830,N_9836);
nand UO_1443 (O_1443,N_9819,N_9913);
or UO_1444 (O_1444,N_9908,N_9896);
nor UO_1445 (O_1445,N_9884,N_9998);
or UO_1446 (O_1446,N_9972,N_9917);
and UO_1447 (O_1447,N_9958,N_9971);
nor UO_1448 (O_1448,N_9938,N_9898);
and UO_1449 (O_1449,N_9822,N_9840);
nand UO_1450 (O_1450,N_9865,N_9995);
nand UO_1451 (O_1451,N_9829,N_9887);
and UO_1452 (O_1452,N_9802,N_9815);
and UO_1453 (O_1453,N_9924,N_9917);
and UO_1454 (O_1454,N_9978,N_9910);
nand UO_1455 (O_1455,N_9802,N_9991);
nor UO_1456 (O_1456,N_9830,N_9833);
nor UO_1457 (O_1457,N_9811,N_9906);
or UO_1458 (O_1458,N_9933,N_9882);
xnor UO_1459 (O_1459,N_9883,N_9837);
nand UO_1460 (O_1460,N_9859,N_9961);
nor UO_1461 (O_1461,N_9881,N_9823);
or UO_1462 (O_1462,N_9978,N_9872);
xor UO_1463 (O_1463,N_9902,N_9949);
xnor UO_1464 (O_1464,N_9847,N_9873);
nand UO_1465 (O_1465,N_9820,N_9982);
and UO_1466 (O_1466,N_9935,N_9987);
nor UO_1467 (O_1467,N_9920,N_9882);
xor UO_1468 (O_1468,N_9834,N_9832);
and UO_1469 (O_1469,N_9809,N_9948);
nand UO_1470 (O_1470,N_9882,N_9907);
and UO_1471 (O_1471,N_9988,N_9802);
and UO_1472 (O_1472,N_9885,N_9864);
nand UO_1473 (O_1473,N_9952,N_9854);
nand UO_1474 (O_1474,N_9860,N_9969);
and UO_1475 (O_1475,N_9929,N_9904);
and UO_1476 (O_1476,N_9826,N_9823);
nand UO_1477 (O_1477,N_9957,N_9879);
nor UO_1478 (O_1478,N_9959,N_9946);
nor UO_1479 (O_1479,N_9878,N_9954);
nor UO_1480 (O_1480,N_9838,N_9994);
or UO_1481 (O_1481,N_9928,N_9939);
nor UO_1482 (O_1482,N_9826,N_9906);
nor UO_1483 (O_1483,N_9873,N_9905);
or UO_1484 (O_1484,N_9900,N_9852);
and UO_1485 (O_1485,N_9808,N_9888);
nand UO_1486 (O_1486,N_9992,N_9822);
and UO_1487 (O_1487,N_9960,N_9852);
nor UO_1488 (O_1488,N_9940,N_9814);
xnor UO_1489 (O_1489,N_9816,N_9868);
nand UO_1490 (O_1490,N_9883,N_9891);
nor UO_1491 (O_1491,N_9907,N_9950);
nor UO_1492 (O_1492,N_9932,N_9974);
xnor UO_1493 (O_1493,N_9849,N_9811);
and UO_1494 (O_1494,N_9956,N_9955);
nor UO_1495 (O_1495,N_9879,N_9856);
xnor UO_1496 (O_1496,N_9808,N_9952);
and UO_1497 (O_1497,N_9961,N_9857);
xnor UO_1498 (O_1498,N_9942,N_9930);
nor UO_1499 (O_1499,N_9878,N_9860);
endmodule