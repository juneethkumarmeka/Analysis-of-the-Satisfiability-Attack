module basic_1500_15000_2000_5_levels_5xor_6(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999;
nor U0 (N_0,In_262,In_284);
nor U1 (N_1,In_888,In_803);
nor U2 (N_2,In_1403,In_940);
nand U3 (N_3,In_1494,In_1363);
nand U4 (N_4,In_781,In_267);
nand U5 (N_5,In_424,In_372);
nand U6 (N_6,In_1488,In_810);
nor U7 (N_7,In_165,In_646);
xnor U8 (N_8,In_708,In_1423);
xnor U9 (N_9,In_840,In_1306);
nand U10 (N_10,In_623,In_1260);
nor U11 (N_11,In_186,In_1320);
nand U12 (N_12,In_239,In_880);
or U13 (N_13,In_35,In_220);
nand U14 (N_14,In_151,In_1169);
nand U15 (N_15,In_271,In_1181);
or U16 (N_16,In_159,In_75);
nor U17 (N_17,In_1120,In_396);
nand U18 (N_18,In_1060,In_535);
or U19 (N_19,In_336,In_672);
nor U20 (N_20,In_81,In_1454);
xnor U21 (N_21,In_668,In_691);
nand U22 (N_22,In_453,In_867);
xnor U23 (N_23,In_1287,In_62);
nor U24 (N_24,In_210,In_1221);
nand U25 (N_25,In_1416,In_748);
and U26 (N_26,In_789,In_847);
nand U27 (N_27,In_1244,In_285);
xor U28 (N_28,In_507,In_371);
nor U29 (N_29,In_700,In_1319);
xor U30 (N_30,In_809,In_1490);
and U31 (N_31,In_856,In_1439);
nor U32 (N_32,In_964,In_169);
nand U33 (N_33,In_138,In_1185);
nand U34 (N_34,In_811,In_823);
xor U35 (N_35,In_370,In_1214);
xnor U36 (N_36,In_1083,In_294);
or U37 (N_37,In_497,In_1467);
nand U38 (N_38,In_554,In_243);
nor U39 (N_39,In_697,In_1112);
nand U40 (N_40,In_530,In_1441);
nand U41 (N_41,In_500,In_1015);
and U42 (N_42,In_1312,In_1497);
nor U43 (N_43,In_449,In_914);
or U44 (N_44,In_322,In_1030);
nand U45 (N_45,In_757,In_956);
or U46 (N_46,In_1462,In_1346);
and U47 (N_47,In_1027,In_911);
xnor U48 (N_48,In_1482,In_233);
nor U49 (N_49,In_894,In_406);
and U50 (N_50,In_1449,In_192);
and U51 (N_51,In_181,In_1079);
or U52 (N_52,In_1066,In_475);
or U53 (N_53,In_1407,In_806);
nand U54 (N_54,In_799,In_896);
and U55 (N_55,In_1379,In_1308);
or U56 (N_56,In_47,In_716);
xnor U57 (N_57,In_144,In_1086);
or U58 (N_58,In_218,In_1450);
nand U59 (N_59,In_69,In_1149);
and U60 (N_60,In_528,In_767);
or U61 (N_61,In_1394,In_320);
and U62 (N_62,In_1213,In_1303);
nand U63 (N_63,In_32,In_899);
xor U64 (N_64,In_1396,In_986);
nor U65 (N_65,In_877,In_93);
xnor U66 (N_66,In_1242,In_1433);
and U67 (N_67,In_216,In_714);
nor U68 (N_68,In_681,In_139);
nand U69 (N_69,In_978,In_965);
nor U70 (N_70,In_288,In_584);
nor U71 (N_71,In_1452,In_934);
nand U72 (N_72,In_146,In_1270);
nor U73 (N_73,In_683,In_1418);
nor U74 (N_74,In_121,In_437);
or U75 (N_75,In_1437,In_70);
or U76 (N_76,In_1434,In_1387);
or U77 (N_77,In_1177,In_1345);
or U78 (N_78,In_1298,In_743);
or U79 (N_79,In_798,In_24);
or U80 (N_80,In_1330,In_727);
and U81 (N_81,In_868,In_351);
nand U82 (N_82,In_593,In_524);
nand U83 (N_83,In_1128,In_452);
and U84 (N_84,In_126,In_689);
or U85 (N_85,In_1348,In_1077);
nor U86 (N_86,In_555,In_1126);
and U87 (N_87,In_585,In_650);
and U88 (N_88,In_1420,In_342);
or U89 (N_89,In_416,In_1310);
or U90 (N_90,In_95,In_28);
or U91 (N_91,In_758,In_183);
and U92 (N_92,In_1406,In_252);
or U93 (N_93,In_393,In_445);
nand U94 (N_94,In_1174,In_1248);
or U95 (N_95,In_785,In_1036);
nor U96 (N_96,In_621,In_208);
nand U97 (N_97,In_821,In_369);
nor U98 (N_98,In_1487,In_704);
nand U99 (N_99,In_1230,In_1273);
nor U100 (N_100,In_227,In_615);
nand U101 (N_101,In_16,In_1121);
or U102 (N_102,In_802,In_468);
nand U103 (N_103,In_1135,In_979);
nor U104 (N_104,In_251,In_383);
nor U105 (N_105,In_1068,In_925);
nand U106 (N_106,In_1334,In_924);
or U107 (N_107,In_235,In_1087);
nor U108 (N_108,In_1047,In_29);
nor U109 (N_109,In_1477,In_588);
nor U110 (N_110,In_1080,In_1251);
and U111 (N_111,In_1305,In_326);
nand U112 (N_112,In_1329,In_901);
or U113 (N_113,In_747,In_1479);
and U114 (N_114,In_1007,In_734);
nor U115 (N_115,In_102,In_594);
or U116 (N_116,In_913,In_1082);
xnor U117 (N_117,In_41,In_3);
or U118 (N_118,In_973,In_1391);
xor U119 (N_119,In_203,In_1096);
or U120 (N_120,In_495,In_985);
nand U121 (N_121,In_611,In_1313);
nand U122 (N_122,In_1364,In_1057);
and U123 (N_123,In_639,In_1026);
or U124 (N_124,In_1259,In_654);
or U125 (N_125,In_223,In_130);
nor U126 (N_126,In_1010,In_1347);
or U127 (N_127,In_381,In_1119);
xnor U128 (N_128,In_548,In_179);
and U129 (N_129,In_110,In_1219);
nand U130 (N_130,In_1243,In_676);
and U131 (N_131,In_824,In_1037);
nand U132 (N_132,In_596,In_932);
nor U133 (N_133,In_553,In_78);
xor U134 (N_134,In_349,In_509);
xor U135 (N_135,In_49,In_1034);
and U136 (N_136,In_470,In_744);
nor U137 (N_137,In_241,In_402);
or U138 (N_138,In_287,In_1);
nand U139 (N_139,In_88,In_1333);
nand U140 (N_140,In_679,In_263);
nand U141 (N_141,In_1155,In_1438);
and U142 (N_142,In_695,In_960);
or U143 (N_143,In_972,In_1466);
and U144 (N_144,In_951,In_68);
and U145 (N_145,In_450,In_542);
xor U146 (N_146,In_1207,In_1088);
nand U147 (N_147,In_995,In_219);
and U148 (N_148,In_1032,In_997);
xor U149 (N_149,In_257,In_387);
nand U150 (N_150,In_1343,In_600);
or U151 (N_151,In_214,In_664);
nand U152 (N_152,In_1218,In_941);
nor U153 (N_153,In_753,In_1326);
nand U154 (N_154,In_247,In_11);
or U155 (N_155,In_544,In_439);
nand U156 (N_156,In_1415,In_1474);
nor U157 (N_157,In_1033,In_1237);
and U158 (N_158,In_1171,In_1295);
or U159 (N_159,In_1304,In_816);
nor U160 (N_160,In_782,In_927);
xor U161 (N_161,In_1231,In_647);
or U162 (N_162,In_1226,In_1435);
xnor U163 (N_163,In_1451,In_1341);
nor U164 (N_164,In_549,In_1388);
nand U165 (N_165,In_278,In_663);
or U166 (N_166,In_626,In_1063);
nor U167 (N_167,In_55,In_486);
or U168 (N_168,In_903,In_461);
nor U169 (N_169,In_390,In_155);
nor U170 (N_170,In_1156,In_1208);
nor U171 (N_171,In_1397,In_754);
nand U172 (N_172,In_1035,In_717);
nand U173 (N_173,In_112,In_1110);
and U174 (N_174,In_887,In_261);
nand U175 (N_175,In_916,In_1378);
xor U176 (N_176,In_526,In_198);
nand U177 (N_177,In_234,In_1151);
and U178 (N_178,In_1311,In_1492);
or U179 (N_179,In_813,In_1323);
or U180 (N_180,In_1301,In_898);
and U181 (N_181,In_355,In_379);
or U182 (N_182,In_1062,In_786);
and U183 (N_183,In_23,In_516);
and U184 (N_184,In_1045,In_1205);
nor U185 (N_185,In_1276,In_187);
nand U186 (N_186,In_632,In_231);
nor U187 (N_187,In_236,In_1113);
or U188 (N_188,In_213,In_204);
or U189 (N_189,In_737,In_161);
nand U190 (N_190,In_10,In_482);
nor U191 (N_191,In_1475,In_414);
or U192 (N_192,In_1458,In_850);
or U193 (N_193,In_1202,In_1483);
and U194 (N_194,In_1382,In_1085);
and U195 (N_195,In_1132,In_1227);
or U196 (N_196,In_597,In_920);
nor U197 (N_197,In_558,In_1131);
nor U198 (N_198,In_1054,In_642);
xnor U199 (N_199,In_303,In_970);
and U200 (N_200,In_795,In_1089);
and U201 (N_201,In_619,In_1162);
or U202 (N_202,In_1336,In_709);
or U203 (N_203,In_624,In_641);
nor U204 (N_204,In_463,In_1495);
and U205 (N_205,In_72,In_556);
and U206 (N_206,In_996,In_1408);
xnor U207 (N_207,In_504,In_300);
and U208 (N_208,In_1142,In_760);
nand U209 (N_209,In_483,In_1101);
nor U210 (N_210,In_1405,In_680);
or U211 (N_211,In_1014,In_959);
nor U212 (N_212,In_428,In_9);
nand U213 (N_213,In_1193,In_1017);
nand U214 (N_214,In_602,In_25);
or U215 (N_215,In_1203,In_567);
and U216 (N_216,In_926,In_852);
nor U217 (N_217,In_419,In_61);
xor U218 (N_218,In_968,In_741);
nor U219 (N_219,In_104,In_890);
nand U220 (N_220,In_1052,In_148);
nand U221 (N_221,In_1152,In_464);
nand U222 (N_222,In_407,In_1414);
or U223 (N_223,In_22,In_409);
nand U224 (N_224,In_1165,In_79);
and U225 (N_225,In_851,In_1258);
or U226 (N_226,In_839,In_1028);
nand U227 (N_227,In_1350,In_701);
or U228 (N_228,In_1109,In_527);
or U229 (N_229,In_1296,In_1404);
xnor U230 (N_230,In_1232,In_1241);
and U231 (N_231,In_1040,In_368);
or U232 (N_232,In_137,In_57);
nand U233 (N_233,In_324,In_736);
and U234 (N_234,In_1029,In_65);
nand U235 (N_235,In_1108,In_343);
nand U236 (N_236,In_822,In_974);
nor U237 (N_237,In_882,In_1375);
and U238 (N_238,In_846,In_91);
nand U239 (N_239,In_961,In_1164);
xnor U240 (N_240,In_15,In_1234);
nor U241 (N_241,In_976,In_853);
or U242 (N_242,In_992,In_1023);
or U243 (N_243,In_1012,In_173);
xnor U244 (N_244,In_1153,In_1344);
nor U245 (N_245,In_832,In_1116);
or U246 (N_246,In_481,In_780);
or U247 (N_247,In_60,In_1421);
xnor U248 (N_248,In_636,In_922);
nand U249 (N_249,In_1018,In_1170);
nor U250 (N_250,In_106,In_429);
nor U251 (N_251,In_457,In_931);
and U252 (N_252,In_671,In_1257);
and U253 (N_253,In_707,In_1496);
xnor U254 (N_254,In_128,In_533);
nand U255 (N_255,In_455,In_761);
nand U256 (N_256,In_1356,In_1184);
nor U257 (N_257,In_589,In_167);
and U258 (N_258,In_1465,In_990);
nor U259 (N_259,In_603,In_1011);
nand U260 (N_260,In_84,In_119);
nand U261 (N_261,In_1392,In_6);
nor U262 (N_262,In_788,In_296);
nand U263 (N_263,In_784,In_1129);
and U264 (N_264,In_675,In_1127);
nand U265 (N_265,In_1078,In_515);
and U266 (N_266,In_238,In_592);
nand U267 (N_267,In_1288,In_583);
or U268 (N_268,In_207,In_1100);
nand U269 (N_269,In_354,In_797);
nand U270 (N_270,In_723,In_694);
nor U271 (N_271,In_87,In_1154);
nand U272 (N_272,In_562,In_1051);
and U273 (N_273,In_1118,In_529);
nor U274 (N_274,In_982,In_1443);
and U275 (N_275,In_967,In_268);
nand U276 (N_276,In_1064,In_1491);
or U277 (N_277,In_933,In_977);
nand U278 (N_278,In_177,In_90);
nand U279 (N_279,In_519,In_1025);
nor U280 (N_280,In_472,In_386);
nand U281 (N_281,In_388,In_521);
nand U282 (N_282,In_40,In_855);
xnor U283 (N_283,In_330,In_667);
nor U284 (N_284,In_1283,In_1267);
and U285 (N_285,In_447,In_4);
or U286 (N_286,In_1215,In_835);
xor U287 (N_287,In_1265,In_45);
and U288 (N_288,In_1206,In_886);
or U289 (N_289,In_1448,In_1370);
or U290 (N_290,In_318,In_185);
nand U291 (N_291,In_752,In_643);
xor U292 (N_292,In_1291,In_1365);
nor U293 (N_293,In_991,In_392);
or U294 (N_294,In_196,In_958);
and U295 (N_295,In_969,In_150);
or U296 (N_296,In_836,In_872);
nor U297 (N_297,In_659,In_1289);
xnor U298 (N_298,In_1331,In_328);
nor U299 (N_299,In_1210,In_1447);
nand U300 (N_300,In_848,In_158);
nor U301 (N_301,In_50,In_564);
or U302 (N_302,In_696,In_1285);
or U303 (N_303,In_232,In_735);
nand U304 (N_304,In_281,In_1358);
xnor U305 (N_305,In_279,In_817);
and U306 (N_306,In_590,In_156);
nand U307 (N_307,In_1061,In_496);
and U308 (N_308,In_1098,In_474);
nand U309 (N_309,In_952,In_77);
or U310 (N_310,In_1481,In_1468);
and U311 (N_311,In_885,In_1194);
or U312 (N_312,In_269,In_1361);
nor U313 (N_313,In_776,In_456);
nor U314 (N_314,In_99,In_249);
nor U315 (N_315,In_963,In_938);
xnor U316 (N_316,In_365,In_508);
xor U317 (N_317,In_1280,In_1383);
nand U318 (N_318,In_522,In_1233);
and U319 (N_319,In_307,In_100);
or U320 (N_320,In_259,In_282);
or U321 (N_321,In_773,In_669);
and U322 (N_322,In_164,In_598);
and U323 (N_323,In_1107,In_1297);
nor U324 (N_324,In_1317,In_484);
and U325 (N_325,In_1158,In_895);
and U326 (N_326,In_1250,In_465);
nor U327 (N_327,In_630,In_143);
and U328 (N_328,In_1190,In_1048);
and U329 (N_329,In_1453,In_154);
or U330 (N_330,In_384,In_892);
nand U331 (N_331,In_266,In_820);
and U332 (N_332,In_140,In_1381);
xor U333 (N_333,In_467,In_702);
or U334 (N_334,In_59,In_1053);
or U335 (N_335,In_473,In_658);
nor U336 (N_336,In_1003,In_692);
and U337 (N_337,In_244,In_339);
and U338 (N_338,In_153,In_131);
nor U339 (N_339,In_107,In_604);
nand U340 (N_340,In_693,In_201);
or U341 (N_341,In_113,In_1180);
nand U342 (N_342,In_572,In_966);
xor U343 (N_343,In_907,In_870);
or U344 (N_344,In_1430,In_631);
nor U345 (N_345,In_340,In_628);
and U346 (N_346,In_730,In_101);
or U347 (N_347,In_194,In_518);
xnor U348 (N_348,In_265,In_510);
nor U349 (N_349,In_713,In_1161);
and U350 (N_350,In_1115,In_206);
or U351 (N_351,In_1476,In_1167);
or U352 (N_352,In_420,In_1266);
nand U353 (N_353,In_1103,In_897);
and U354 (N_354,In_353,In_812);
nor U355 (N_355,In_804,In_649);
or U356 (N_356,In_489,In_135);
xor U357 (N_357,In_1472,In_842);
and U358 (N_358,In_1102,In_711);
nor U359 (N_359,In_532,In_175);
nor U360 (N_360,In_1369,In_7);
or U361 (N_361,In_1125,In_1354);
or U362 (N_362,In_557,In_491);
and U363 (N_363,In_385,In_1293);
or U364 (N_364,In_613,In_1236);
nand U365 (N_365,In_831,In_579);
nor U366 (N_366,In_1046,In_1140);
nor U367 (N_367,In_601,In_124);
and U368 (N_368,In_1145,In_605);
nand U369 (N_369,In_272,In_994);
nand U370 (N_370,In_1412,In_415);
and U371 (N_371,In_666,In_1067);
and U372 (N_372,In_792,In_1039);
nor U373 (N_373,In_117,In_405);
and U374 (N_374,In_577,In_85);
or U375 (N_375,In_791,In_860);
or U376 (N_376,In_1262,In_205);
or U377 (N_377,In_1009,In_1385);
or U378 (N_378,In_1016,In_536);
nor U379 (N_379,In_1264,In_180);
or U380 (N_380,In_344,In_308);
xnor U381 (N_381,In_346,In_1372);
or U382 (N_382,In_1020,In_480);
or U383 (N_383,In_722,In_721);
xor U384 (N_384,In_1031,In_1278);
and U385 (N_385,In_1389,In_248);
or U386 (N_386,In_255,In_1008);
nand U387 (N_387,In_844,In_302);
nand U388 (N_388,In_550,In_616);
nand U389 (N_389,In_923,In_298);
nand U390 (N_390,In_1058,In_999);
nand U391 (N_391,In_1198,In_634);
and U392 (N_392,In_1073,In_1359);
nand U393 (N_393,In_541,In_929);
or U394 (N_394,In_1091,In_1252);
and U395 (N_395,In_1228,In_1186);
nand U396 (N_396,In_200,In_942);
nand U397 (N_397,In_1001,In_289);
nor U398 (N_398,In_622,In_525);
nor U399 (N_399,In_937,In_477);
nor U400 (N_400,In_418,In_382);
nor U401 (N_401,In_750,In_685);
nor U402 (N_402,In_580,In_1124);
nor U403 (N_403,In_1486,In_1484);
nor U404 (N_404,In_193,In_987);
nor U405 (N_405,In_1272,In_984);
or U406 (N_406,In_690,In_1444);
nand U407 (N_407,In_1390,In_170);
and U408 (N_408,In_1282,In_221);
and U409 (N_409,In_17,In_1106);
or U410 (N_410,In_38,In_808);
nor U411 (N_411,In_655,In_1093);
and U412 (N_412,In_1290,In_1411);
and U413 (N_413,In_152,In_830);
nor U414 (N_414,In_48,In_1144);
nor U415 (N_415,In_404,In_1179);
or U416 (N_416,In_618,In_715);
or U417 (N_417,In_998,In_794);
or U418 (N_418,In_1263,In_316);
nor U419 (N_419,In_228,In_774);
or U420 (N_420,In_947,In_438);
nand U421 (N_421,In_58,In_1137);
nor U422 (N_422,In_408,In_86);
and U423 (N_423,In_242,In_865);
or U424 (N_424,In_367,In_1188);
or U425 (N_425,In_825,In_26);
nand U426 (N_426,In_779,In_1070);
or U427 (N_427,In_653,In_134);
xnor U428 (N_428,In_313,In_762);
xor U429 (N_429,In_46,In_1445);
nor U430 (N_430,In_195,In_1211);
or U431 (N_431,In_710,In_625);
xor U432 (N_432,In_96,In_432);
nand U433 (N_433,In_571,In_291);
or U434 (N_434,In_1410,In_845);
nand U435 (N_435,In_1299,In_534);
or U436 (N_436,In_1173,In_738);
nor U437 (N_437,In_391,In_191);
nand U438 (N_438,In_1292,In_512);
or U439 (N_439,In_801,In_904);
nand U440 (N_440,In_426,In_43);
or U441 (N_441,In_361,In_157);
nand U442 (N_442,In_768,In_930);
or U443 (N_443,In_394,In_494);
or U444 (N_444,In_66,In_1401);
or U445 (N_445,In_502,In_260);
nand U446 (N_446,In_380,In_657);
nor U447 (N_447,In_436,In_487);
nand U448 (N_448,In_523,In_1338);
or U449 (N_449,In_1090,In_1143);
and U450 (N_450,In_1327,In_610);
and U451 (N_451,In_1376,In_423);
or U452 (N_452,In_314,In_1166);
nor U453 (N_453,In_335,In_20);
and U454 (N_454,In_172,In_398);
nand U455 (N_455,In_975,In_1335);
and U456 (N_456,In_787,In_162);
nor U457 (N_457,In_168,In_576);
nand U458 (N_458,In_103,In_292);
nor U459 (N_459,In_1328,In_1300);
or U460 (N_460,In_678,In_935);
nor U461 (N_461,In_1440,In_1013);
and U462 (N_462,In_902,In_127);
nor U463 (N_463,In_401,In_1357);
and U464 (N_464,In_1360,In_211);
nand U465 (N_465,In_725,In_569);
and U466 (N_466,In_828,In_74);
nor U467 (N_467,In_347,In_1340);
nand U468 (N_468,In_1480,In_256);
and U469 (N_469,In_364,In_76);
xnor U470 (N_470,In_270,In_63);
xor U471 (N_471,In_304,In_1470);
or U472 (N_472,In_1240,In_1247);
and U473 (N_473,In_1111,In_1302);
nand U474 (N_474,In_80,In_764);
nor U475 (N_475,In_1307,In_814);
nand U476 (N_476,In_315,In_720);
nor U477 (N_477,In_478,In_319);
nand U478 (N_478,In_297,In_1038);
or U479 (N_479,In_869,In_425);
nor U480 (N_480,In_83,In_943);
xnor U481 (N_481,In_366,In_1367);
or U482 (N_482,In_769,In_1196);
and U483 (N_483,In_740,In_51);
or U484 (N_484,In_413,In_566);
nor U485 (N_485,In_751,In_105);
xnor U486 (N_486,In_706,In_1192);
xor U487 (N_487,In_1429,In_332);
or U488 (N_488,In_705,In_833);
nand U489 (N_489,In_673,In_19);
nor U490 (N_490,In_1209,In_909);
nand U491 (N_491,In_499,In_862);
nor U492 (N_492,In_399,In_1284);
and U493 (N_493,In_1351,In_133);
or U494 (N_494,In_444,In_1099);
or U495 (N_495,In_333,In_893);
and U496 (N_496,In_854,In_1374);
nor U497 (N_497,In_18,In_863);
nor U498 (N_498,In_250,In_1183);
nor U499 (N_499,In_608,In_1493);
nor U500 (N_500,In_182,In_640);
nor U501 (N_501,In_1021,In_1402);
and U502 (N_502,In_859,In_337);
or U503 (N_503,In_226,In_800);
nand U504 (N_504,In_1222,In_638);
and U505 (N_505,In_276,In_498);
nand U506 (N_506,In_1160,In_217);
and U507 (N_507,In_501,In_1148);
nor U508 (N_508,In_145,In_581);
nor U509 (N_509,In_389,In_570);
or U510 (N_510,In_511,In_699);
or U511 (N_511,In_980,In_1104);
nor U512 (N_512,In_34,In_724);
nand U513 (N_513,In_1473,In_873);
and U514 (N_514,In_560,In_1332);
nor U515 (N_515,In_136,In_957);
nor U516 (N_516,In_687,In_1220);
nor U517 (N_517,In_772,In_1373);
xnor U518 (N_518,In_363,In_42);
nor U519 (N_519,In_540,In_1176);
nand U520 (N_520,In_188,In_190);
and U521 (N_521,In_442,In_1498);
nand U522 (N_522,In_954,In_275);
nand U523 (N_523,In_1446,In_645);
and U524 (N_524,In_1212,In_749);
or U525 (N_525,In_1134,In_73);
or U526 (N_526,In_1094,In_1428);
nor U527 (N_527,In_375,In_237);
and U528 (N_528,In_1239,In_612);
or U529 (N_529,In_1342,In_1425);
nor U530 (N_530,In_686,In_240);
xnor U531 (N_531,In_397,In_635);
or U532 (N_532,In_866,In_614);
and U533 (N_533,In_1413,In_1175);
nor U534 (N_534,In_174,In_321);
nor U535 (N_535,In_21,In_900);
nand U536 (N_536,In_1024,In_841);
xnor U537 (N_537,In_563,In_1076);
and U538 (N_538,In_476,In_1150);
nor U539 (N_539,In_1294,In_759);
or U540 (N_540,In_125,In_1172);
or U541 (N_541,In_258,In_629);
nor U542 (N_542,In_1271,In_1200);
or U543 (N_543,In_224,In_1136);
xor U544 (N_544,In_1349,In_908);
nor U545 (N_545,In_312,In_732);
and U546 (N_546,In_264,In_1041);
or U547 (N_547,In_503,In_1380);
xnor U548 (N_548,In_905,In_441);
nand U549 (N_549,In_412,In_729);
or U550 (N_550,In_988,In_637);
and U551 (N_551,In_1274,In_765);
nor U552 (N_552,In_141,In_12);
xnor U553 (N_553,In_1217,In_559);
xnor U554 (N_554,In_123,In_871);
nor U555 (N_555,In_466,In_1059);
nand U556 (N_556,In_771,In_1424);
nor U557 (N_557,In_325,In_1235);
nand U558 (N_558,In_1355,In_981);
nor U559 (N_559,In_178,In_568);
and U560 (N_560,In_493,In_652);
xor U561 (N_561,In_921,In_807);
or U562 (N_562,In_492,In_1147);
nand U563 (N_563,In_458,In_362);
and U564 (N_564,In_745,In_334);
nor U565 (N_565,In_1269,In_688);
nor U566 (N_566,In_197,In_827);
nand U567 (N_567,In_962,In_1163);
nor U568 (N_568,In_587,In_94);
nand U569 (N_569,In_485,In_1309);
nand U570 (N_570,In_858,In_971);
xnor U571 (N_571,In_1256,In_33);
nor U572 (N_572,In_936,In_1075);
nand U573 (N_573,In_617,In_395);
nor U574 (N_574,In_620,In_1318);
and U575 (N_575,In_718,In_698);
xor U576 (N_576,In_1314,In_818);
and U577 (N_577,In_1069,In_273);
nor U578 (N_578,In_864,In_1225);
nand U579 (N_579,In_1105,In_1187);
nor U580 (N_580,In_1261,In_1049);
nor U581 (N_581,In_1464,In_82);
nand U582 (N_582,In_883,In_815);
nand U583 (N_583,In_1055,In_728);
and U584 (N_584,In_775,In_1224);
nor U585 (N_585,In_849,In_586);
or U586 (N_586,In_254,In_513);
and U587 (N_587,In_1182,In_338);
nand U588 (N_588,In_1006,In_1419);
nor U589 (N_589,In_1072,In_27);
nand U590 (N_590,In_1138,In_403);
or U591 (N_591,In_1386,In_1253);
or U592 (N_592,In_199,In_843);
or U593 (N_593,In_537,In_1114);
and U594 (N_594,In_1000,In_5);
nor U595 (N_595,In_1268,In_881);
nor U596 (N_596,In_884,In_948);
nor U597 (N_597,In_430,In_551);
nand U598 (N_598,In_245,In_64);
and U599 (N_599,In_1489,In_944);
nand U600 (N_600,In_1427,In_546);
nand U601 (N_601,In_1461,In_1229);
nor U602 (N_602,In_111,In_277);
or U603 (N_603,In_230,In_306);
nand U604 (N_604,In_376,In_1195);
nand U605 (N_605,In_606,In_607);
nand U606 (N_606,In_1399,In_1325);
or U607 (N_607,In_1071,In_609);
or U608 (N_608,In_1442,In_1281);
or U609 (N_609,In_661,In_1322);
nand U610 (N_610,In_796,In_1084);
or U611 (N_611,In_1395,In_939);
nor U612 (N_612,In_1157,In_946);
or U613 (N_613,In_1478,In_451);
nand U614 (N_614,In_54,In_1499);
or U615 (N_615,In_684,In_129);
nor U616 (N_616,In_1426,In_746);
and U617 (N_617,In_310,In_1216);
nor U618 (N_618,In_417,In_479);
xor U619 (N_619,In_30,In_1081);
or U620 (N_620,In_1277,In_89);
or U621 (N_621,In_591,In_360);
nor U622 (N_622,In_1485,In_1042);
or U623 (N_623,In_599,In_1074);
or U624 (N_624,In_644,In_1050);
or U625 (N_625,In_506,In_949);
or U626 (N_626,In_280,In_552);
nor U627 (N_627,In_331,In_374);
nand U628 (N_628,In_53,In_674);
or U629 (N_629,In_52,In_1422);
nor U630 (N_630,In_574,In_1366);
or U631 (N_631,In_13,In_1398);
or U632 (N_632,In_919,In_1191);
or U633 (N_633,In_443,In_726);
nor U634 (N_634,In_373,In_1159);
xnor U635 (N_635,In_1122,In_448);
and U636 (N_636,In_2,In_1005);
nand U637 (N_637,In_575,In_215);
or U638 (N_638,In_915,In_878);
and U639 (N_639,In_132,In_766);
or U640 (N_640,In_793,In_202);
or U641 (N_641,In_37,In_1409);
and U642 (N_642,In_819,In_56);
and U643 (N_643,In_359,In_1431);
nor U644 (N_644,In_1255,In_1460);
xor U645 (N_645,In_875,In_648);
nand U646 (N_646,In_1197,In_538);
or U647 (N_647,In_1393,In_756);
nand U648 (N_648,In_834,In_517);
nand U649 (N_649,In_345,In_97);
xnor U650 (N_650,In_1436,In_212);
or U651 (N_651,In_400,In_378);
nor U652 (N_652,In_431,In_1362);
or U653 (N_653,In_783,In_184);
or U654 (N_654,In_1238,In_283);
and U655 (N_655,In_1459,In_719);
and U656 (N_656,In_350,In_545);
or U657 (N_657,In_171,In_1275);
nor U658 (N_658,In_891,In_301);
nor U659 (N_659,In_329,In_918);
or U660 (N_660,In_829,In_953);
nor U661 (N_661,In_1321,In_116);
or U662 (N_662,In_703,In_147);
nor U663 (N_663,In_286,In_149);
and U664 (N_664,In_677,In_454);
or U665 (N_665,In_98,In_462);
nor U666 (N_666,In_656,In_1384);
nor U667 (N_667,In_118,In_1417);
and U668 (N_668,In_44,In_876);
nand U669 (N_669,In_160,In_323);
nor U670 (N_670,In_410,In_293);
nand U671 (N_671,In_471,In_573);
and U672 (N_672,In_912,In_950);
or U673 (N_673,In_460,In_427);
nor U674 (N_674,In_1178,In_488);
nor U675 (N_675,In_1469,In_356);
and U676 (N_676,In_627,In_739);
and U677 (N_677,In_1043,In_857);
and U678 (N_678,In_561,In_1371);
nor U679 (N_679,In_1002,In_163);
and U680 (N_680,In_440,In_1246);
or U681 (N_681,In_1400,In_446);
xnor U682 (N_682,In_122,In_1456);
and U683 (N_683,In_861,In_421);
nor U684 (N_684,In_1368,In_67);
or U685 (N_685,In_299,In_514);
nor U686 (N_686,In_1019,In_327);
nor U687 (N_687,In_578,In_377);
and U688 (N_688,In_176,In_1056);
and U689 (N_689,In_108,In_805);
nor U690 (N_690,In_0,In_879);
or U691 (N_691,In_1168,In_435);
nor U692 (N_692,In_92,In_712);
and U693 (N_693,In_229,In_928);
nor U694 (N_694,In_1189,In_305);
and U695 (N_695,In_341,In_910);
nor U696 (N_696,In_352,In_1204);
or U697 (N_697,In_777,In_955);
nor U698 (N_698,In_31,In_838);
and U699 (N_699,In_71,In_582);
nor U700 (N_700,In_837,In_731);
nor U701 (N_701,In_36,In_295);
nand U702 (N_702,In_778,In_742);
or U703 (N_703,In_1095,In_1455);
nand U704 (N_704,In_531,In_1223);
or U705 (N_705,In_993,In_1141);
nand U706 (N_706,In_189,In_209);
nor U707 (N_707,In_1324,In_1117);
or U708 (N_708,In_790,In_1432);
nor U709 (N_709,In_433,In_1199);
nor U710 (N_710,In_633,In_670);
nand U711 (N_711,In_1130,In_109);
nor U712 (N_712,In_505,In_1146);
or U713 (N_713,In_945,In_1353);
nor U714 (N_714,In_290,In_1471);
nor U715 (N_715,In_1254,In_763);
nand U716 (N_716,In_889,In_874);
nor U717 (N_717,In_983,In_1316);
and U718 (N_718,In_253,In_1201);
nand U719 (N_719,In_115,In_246);
or U720 (N_720,In_1377,In_1139);
or U721 (N_721,In_651,In_8);
nor U722 (N_722,In_1022,In_733);
xor U723 (N_723,In_411,In_142);
and U724 (N_724,In_422,In_114);
or U725 (N_725,In_317,In_490);
nand U726 (N_726,In_459,In_660);
xnor U727 (N_727,In_120,In_989);
or U728 (N_728,In_906,In_682);
or U729 (N_729,In_348,In_665);
and U730 (N_730,In_1133,In_39);
nor U731 (N_731,In_917,In_1337);
xnor U732 (N_732,In_520,In_595);
nand U733 (N_733,In_274,In_1065);
and U734 (N_734,In_14,In_1004);
nor U735 (N_735,In_826,In_311);
nor U736 (N_736,In_662,In_222);
nor U737 (N_737,In_469,In_1097);
and U738 (N_738,In_166,In_309);
and U739 (N_739,In_543,In_755);
or U740 (N_740,In_225,In_1249);
and U741 (N_741,In_1123,In_1339);
nand U742 (N_742,In_1245,In_1463);
nor U743 (N_743,In_770,In_539);
and U744 (N_744,In_357,In_565);
or U745 (N_745,In_1279,In_1457);
nor U746 (N_746,In_1352,In_1044);
or U747 (N_747,In_547,In_434);
and U748 (N_748,In_1315,In_358);
nand U749 (N_749,In_1286,In_1092);
xor U750 (N_750,In_190,In_1088);
nand U751 (N_751,In_733,In_892);
and U752 (N_752,In_363,In_432);
or U753 (N_753,In_1256,In_304);
and U754 (N_754,In_1460,In_1459);
xnor U755 (N_755,In_266,In_2);
and U756 (N_756,In_1480,In_994);
or U757 (N_757,In_900,In_1450);
nor U758 (N_758,In_1014,In_675);
and U759 (N_759,In_134,In_89);
xor U760 (N_760,In_739,In_780);
or U761 (N_761,In_1458,In_567);
nor U762 (N_762,In_692,In_1333);
or U763 (N_763,In_990,In_803);
and U764 (N_764,In_260,In_108);
or U765 (N_765,In_19,In_546);
xnor U766 (N_766,In_435,In_841);
and U767 (N_767,In_985,In_480);
and U768 (N_768,In_1371,In_1460);
nand U769 (N_769,In_833,In_10);
nand U770 (N_770,In_1432,In_1346);
and U771 (N_771,In_887,In_706);
xnor U772 (N_772,In_789,In_1041);
nand U773 (N_773,In_895,In_589);
nor U774 (N_774,In_421,In_931);
xor U775 (N_775,In_1326,In_963);
and U776 (N_776,In_1260,In_1407);
nor U777 (N_777,In_389,In_900);
or U778 (N_778,In_1188,In_1316);
nor U779 (N_779,In_1203,In_717);
nand U780 (N_780,In_338,In_975);
nor U781 (N_781,In_1334,In_940);
nand U782 (N_782,In_850,In_478);
nor U783 (N_783,In_1119,In_1474);
nand U784 (N_784,In_1326,In_154);
nand U785 (N_785,In_22,In_741);
nor U786 (N_786,In_1310,In_507);
or U787 (N_787,In_1060,In_989);
nor U788 (N_788,In_321,In_12);
nand U789 (N_789,In_241,In_149);
nand U790 (N_790,In_614,In_1102);
or U791 (N_791,In_1446,In_1012);
xor U792 (N_792,In_27,In_1342);
nand U793 (N_793,In_683,In_799);
or U794 (N_794,In_979,In_911);
or U795 (N_795,In_184,In_1136);
or U796 (N_796,In_638,In_1161);
and U797 (N_797,In_170,In_1198);
nor U798 (N_798,In_183,In_1259);
and U799 (N_799,In_795,In_424);
xor U800 (N_800,In_1068,In_350);
nor U801 (N_801,In_262,In_958);
or U802 (N_802,In_1137,In_708);
and U803 (N_803,In_345,In_680);
nand U804 (N_804,In_308,In_35);
and U805 (N_805,In_885,In_599);
nand U806 (N_806,In_805,In_1110);
nand U807 (N_807,In_551,In_1366);
nand U808 (N_808,In_499,In_920);
nand U809 (N_809,In_807,In_1254);
and U810 (N_810,In_181,In_839);
and U811 (N_811,In_1166,In_1192);
or U812 (N_812,In_1309,In_378);
and U813 (N_813,In_1109,In_1360);
xnor U814 (N_814,In_736,In_1447);
and U815 (N_815,In_208,In_343);
nand U816 (N_816,In_637,In_1131);
nand U817 (N_817,In_1054,In_1123);
or U818 (N_818,In_1470,In_158);
nor U819 (N_819,In_1082,In_402);
and U820 (N_820,In_1351,In_381);
nand U821 (N_821,In_1167,In_1022);
or U822 (N_822,In_526,In_727);
and U823 (N_823,In_939,In_1308);
xnor U824 (N_824,In_1081,In_849);
nand U825 (N_825,In_1015,In_1102);
nand U826 (N_826,In_62,In_1142);
or U827 (N_827,In_883,In_1229);
nand U828 (N_828,In_1283,In_648);
and U829 (N_829,In_561,In_813);
or U830 (N_830,In_282,In_511);
xor U831 (N_831,In_1181,In_625);
or U832 (N_832,In_994,In_301);
nand U833 (N_833,In_1075,In_182);
nand U834 (N_834,In_327,In_1280);
xnor U835 (N_835,In_604,In_1280);
nand U836 (N_836,In_341,In_450);
nand U837 (N_837,In_188,In_416);
nand U838 (N_838,In_1342,In_657);
nor U839 (N_839,In_169,In_1222);
nand U840 (N_840,In_146,In_230);
xor U841 (N_841,In_299,In_546);
nor U842 (N_842,In_627,In_159);
nand U843 (N_843,In_1325,In_1013);
or U844 (N_844,In_831,In_208);
nand U845 (N_845,In_988,In_1143);
nand U846 (N_846,In_1359,In_1433);
nand U847 (N_847,In_844,In_43);
and U848 (N_848,In_930,In_1248);
nor U849 (N_849,In_291,In_1433);
nor U850 (N_850,In_51,In_879);
or U851 (N_851,In_325,In_567);
nor U852 (N_852,In_183,In_1497);
and U853 (N_853,In_477,In_1103);
or U854 (N_854,In_788,In_928);
or U855 (N_855,In_1470,In_1029);
nand U856 (N_856,In_905,In_26);
nor U857 (N_857,In_806,In_1399);
xor U858 (N_858,In_1387,In_557);
and U859 (N_859,In_1329,In_133);
or U860 (N_860,In_10,In_355);
xor U861 (N_861,In_335,In_683);
nand U862 (N_862,In_1302,In_1164);
and U863 (N_863,In_738,In_772);
or U864 (N_864,In_434,In_601);
or U865 (N_865,In_305,In_1132);
and U866 (N_866,In_975,In_28);
and U867 (N_867,In_36,In_944);
nor U868 (N_868,In_209,In_1268);
nand U869 (N_869,In_427,In_1430);
and U870 (N_870,In_1318,In_709);
and U871 (N_871,In_295,In_0);
nor U872 (N_872,In_687,In_280);
and U873 (N_873,In_832,In_1042);
and U874 (N_874,In_290,In_1196);
and U875 (N_875,In_875,In_304);
nor U876 (N_876,In_817,In_740);
and U877 (N_877,In_735,In_870);
or U878 (N_878,In_447,In_276);
xor U879 (N_879,In_968,In_828);
nand U880 (N_880,In_983,In_296);
or U881 (N_881,In_345,In_486);
or U882 (N_882,In_390,In_280);
nand U883 (N_883,In_891,In_878);
or U884 (N_884,In_730,In_536);
and U885 (N_885,In_821,In_31);
nand U886 (N_886,In_510,In_1440);
nand U887 (N_887,In_722,In_1229);
or U888 (N_888,In_1342,In_242);
nor U889 (N_889,In_783,In_655);
or U890 (N_890,In_306,In_969);
nand U891 (N_891,In_1423,In_302);
and U892 (N_892,In_433,In_673);
or U893 (N_893,In_631,In_368);
nor U894 (N_894,In_71,In_1152);
or U895 (N_895,In_100,In_240);
or U896 (N_896,In_68,In_1441);
nand U897 (N_897,In_7,In_1332);
xor U898 (N_898,In_1007,In_414);
nand U899 (N_899,In_162,In_1288);
nand U900 (N_900,In_1182,In_385);
nand U901 (N_901,In_1358,In_1299);
and U902 (N_902,In_530,In_1074);
nor U903 (N_903,In_682,In_1096);
nor U904 (N_904,In_889,In_1454);
nand U905 (N_905,In_1458,In_156);
or U906 (N_906,In_377,In_712);
or U907 (N_907,In_184,In_967);
xor U908 (N_908,In_590,In_707);
xor U909 (N_909,In_200,In_133);
and U910 (N_910,In_1203,In_158);
or U911 (N_911,In_777,In_706);
and U912 (N_912,In_228,In_240);
nor U913 (N_913,In_1129,In_454);
or U914 (N_914,In_203,In_633);
nor U915 (N_915,In_833,In_1406);
or U916 (N_916,In_9,In_547);
or U917 (N_917,In_759,In_259);
or U918 (N_918,In_1141,In_810);
nand U919 (N_919,In_1405,In_1426);
nand U920 (N_920,In_701,In_1023);
and U921 (N_921,In_937,In_1110);
nor U922 (N_922,In_156,In_309);
and U923 (N_923,In_136,In_1138);
nand U924 (N_924,In_333,In_241);
and U925 (N_925,In_801,In_708);
nor U926 (N_926,In_1358,In_1060);
or U927 (N_927,In_1100,In_1108);
nand U928 (N_928,In_908,In_947);
or U929 (N_929,In_656,In_573);
nand U930 (N_930,In_366,In_170);
or U931 (N_931,In_747,In_1331);
or U932 (N_932,In_448,In_1126);
xor U933 (N_933,In_1227,In_1162);
nor U934 (N_934,In_1143,In_744);
nor U935 (N_935,In_787,In_985);
nor U936 (N_936,In_1118,In_1304);
or U937 (N_937,In_703,In_605);
and U938 (N_938,In_972,In_1108);
or U939 (N_939,In_523,In_1405);
or U940 (N_940,In_29,In_1257);
xor U941 (N_941,In_70,In_971);
or U942 (N_942,In_818,In_1470);
and U943 (N_943,In_1334,In_328);
and U944 (N_944,In_1164,In_1208);
and U945 (N_945,In_452,In_667);
or U946 (N_946,In_868,In_244);
nand U947 (N_947,In_1361,In_859);
and U948 (N_948,In_1409,In_462);
and U949 (N_949,In_1288,In_188);
xnor U950 (N_950,In_157,In_1307);
or U951 (N_951,In_983,In_25);
xnor U952 (N_952,In_551,In_360);
nand U953 (N_953,In_1490,In_1066);
or U954 (N_954,In_1338,In_918);
nand U955 (N_955,In_45,In_1447);
nor U956 (N_956,In_916,In_1309);
and U957 (N_957,In_280,In_1241);
xnor U958 (N_958,In_1484,In_415);
or U959 (N_959,In_455,In_1354);
xnor U960 (N_960,In_232,In_1353);
or U961 (N_961,In_874,In_532);
and U962 (N_962,In_933,In_819);
and U963 (N_963,In_1125,In_105);
or U964 (N_964,In_1307,In_278);
nand U965 (N_965,In_292,In_1385);
nand U966 (N_966,In_1338,In_1316);
xor U967 (N_967,In_538,In_687);
or U968 (N_968,In_1498,In_915);
or U969 (N_969,In_226,In_1077);
or U970 (N_970,In_198,In_1140);
xnor U971 (N_971,In_761,In_142);
or U972 (N_972,In_1039,In_753);
and U973 (N_973,In_363,In_63);
nand U974 (N_974,In_1264,In_1136);
nor U975 (N_975,In_699,In_287);
and U976 (N_976,In_581,In_291);
and U977 (N_977,In_939,In_602);
and U978 (N_978,In_1345,In_262);
and U979 (N_979,In_19,In_48);
nand U980 (N_980,In_1162,In_100);
and U981 (N_981,In_566,In_1441);
or U982 (N_982,In_94,In_36);
nand U983 (N_983,In_1252,In_159);
or U984 (N_984,In_431,In_496);
or U985 (N_985,In_255,In_231);
nor U986 (N_986,In_1206,In_746);
and U987 (N_987,In_644,In_895);
and U988 (N_988,In_1069,In_1190);
nand U989 (N_989,In_194,In_508);
or U990 (N_990,In_1495,In_459);
and U991 (N_991,In_747,In_199);
and U992 (N_992,In_65,In_226);
or U993 (N_993,In_207,In_566);
or U994 (N_994,In_824,In_933);
nor U995 (N_995,In_770,In_492);
nand U996 (N_996,In_922,In_967);
xnor U997 (N_997,In_600,In_889);
and U998 (N_998,In_60,In_1356);
or U999 (N_999,In_236,In_419);
nand U1000 (N_1000,In_1433,In_343);
or U1001 (N_1001,In_809,In_740);
nor U1002 (N_1002,In_323,In_899);
and U1003 (N_1003,In_566,In_43);
and U1004 (N_1004,In_1139,In_1417);
and U1005 (N_1005,In_960,In_1176);
xor U1006 (N_1006,In_614,In_1407);
and U1007 (N_1007,In_460,In_270);
or U1008 (N_1008,In_884,In_393);
or U1009 (N_1009,In_1368,In_512);
nand U1010 (N_1010,In_112,In_800);
nand U1011 (N_1011,In_562,In_954);
nor U1012 (N_1012,In_725,In_45);
and U1013 (N_1013,In_580,In_1402);
nand U1014 (N_1014,In_864,In_391);
and U1015 (N_1015,In_535,In_74);
or U1016 (N_1016,In_227,In_1228);
nor U1017 (N_1017,In_877,In_271);
or U1018 (N_1018,In_51,In_663);
and U1019 (N_1019,In_203,In_907);
nand U1020 (N_1020,In_479,In_1079);
nor U1021 (N_1021,In_1236,In_448);
or U1022 (N_1022,In_1447,In_191);
nand U1023 (N_1023,In_1154,In_1238);
and U1024 (N_1024,In_873,In_696);
or U1025 (N_1025,In_502,In_377);
nor U1026 (N_1026,In_1094,In_327);
nand U1027 (N_1027,In_1363,In_1269);
nor U1028 (N_1028,In_784,In_1170);
or U1029 (N_1029,In_1266,In_113);
or U1030 (N_1030,In_1253,In_868);
or U1031 (N_1031,In_296,In_1009);
nor U1032 (N_1032,In_718,In_628);
nand U1033 (N_1033,In_272,In_971);
nand U1034 (N_1034,In_777,In_3);
or U1035 (N_1035,In_592,In_10);
or U1036 (N_1036,In_680,In_586);
and U1037 (N_1037,In_238,In_922);
and U1038 (N_1038,In_29,In_354);
and U1039 (N_1039,In_1271,In_1100);
and U1040 (N_1040,In_1451,In_1298);
nor U1041 (N_1041,In_889,In_673);
xnor U1042 (N_1042,In_596,In_1361);
and U1043 (N_1043,In_768,In_865);
nor U1044 (N_1044,In_994,In_852);
nor U1045 (N_1045,In_799,In_765);
or U1046 (N_1046,In_266,In_38);
and U1047 (N_1047,In_140,In_136);
nand U1048 (N_1048,In_812,In_1484);
nor U1049 (N_1049,In_1349,In_1031);
and U1050 (N_1050,In_856,In_489);
and U1051 (N_1051,In_385,In_1112);
or U1052 (N_1052,In_1499,In_1207);
and U1053 (N_1053,In_678,In_1489);
nand U1054 (N_1054,In_904,In_775);
nand U1055 (N_1055,In_591,In_154);
or U1056 (N_1056,In_618,In_587);
and U1057 (N_1057,In_1342,In_860);
and U1058 (N_1058,In_60,In_1453);
nand U1059 (N_1059,In_1379,In_386);
or U1060 (N_1060,In_156,In_1434);
nor U1061 (N_1061,In_199,In_418);
or U1062 (N_1062,In_972,In_29);
nor U1063 (N_1063,In_63,In_534);
nor U1064 (N_1064,In_1008,In_822);
or U1065 (N_1065,In_1357,In_36);
and U1066 (N_1066,In_814,In_1200);
nand U1067 (N_1067,In_1135,In_679);
or U1068 (N_1068,In_1269,In_273);
nand U1069 (N_1069,In_504,In_1065);
nand U1070 (N_1070,In_724,In_339);
nor U1071 (N_1071,In_133,In_1376);
or U1072 (N_1072,In_741,In_282);
xnor U1073 (N_1073,In_1333,In_659);
and U1074 (N_1074,In_236,In_576);
xnor U1075 (N_1075,In_47,In_532);
nand U1076 (N_1076,In_948,In_331);
and U1077 (N_1077,In_522,In_201);
xnor U1078 (N_1078,In_842,In_386);
xor U1079 (N_1079,In_298,In_1042);
or U1080 (N_1080,In_621,In_1294);
or U1081 (N_1081,In_1424,In_1417);
and U1082 (N_1082,In_1272,In_617);
or U1083 (N_1083,In_1376,In_260);
or U1084 (N_1084,In_383,In_1412);
or U1085 (N_1085,In_572,In_628);
nand U1086 (N_1086,In_1233,In_143);
and U1087 (N_1087,In_1298,In_1326);
nand U1088 (N_1088,In_308,In_946);
nand U1089 (N_1089,In_1490,In_953);
nand U1090 (N_1090,In_382,In_302);
and U1091 (N_1091,In_889,In_726);
or U1092 (N_1092,In_1306,In_78);
and U1093 (N_1093,In_758,In_630);
xor U1094 (N_1094,In_249,In_1442);
nor U1095 (N_1095,In_82,In_83);
nand U1096 (N_1096,In_1041,In_614);
and U1097 (N_1097,In_913,In_968);
and U1098 (N_1098,In_349,In_705);
and U1099 (N_1099,In_33,In_1129);
xnor U1100 (N_1100,In_921,In_690);
and U1101 (N_1101,In_1301,In_587);
nand U1102 (N_1102,In_1092,In_1415);
xnor U1103 (N_1103,In_1295,In_119);
nor U1104 (N_1104,In_1209,In_341);
or U1105 (N_1105,In_278,In_1483);
nand U1106 (N_1106,In_356,In_60);
nand U1107 (N_1107,In_1238,In_525);
or U1108 (N_1108,In_1445,In_979);
nor U1109 (N_1109,In_69,In_1044);
and U1110 (N_1110,In_1004,In_1293);
and U1111 (N_1111,In_76,In_783);
and U1112 (N_1112,In_718,In_1470);
or U1113 (N_1113,In_1313,In_273);
nand U1114 (N_1114,In_302,In_100);
and U1115 (N_1115,In_839,In_586);
nand U1116 (N_1116,In_127,In_25);
nand U1117 (N_1117,In_798,In_865);
or U1118 (N_1118,In_522,In_438);
and U1119 (N_1119,In_869,In_1472);
and U1120 (N_1120,In_374,In_130);
nand U1121 (N_1121,In_81,In_1144);
xor U1122 (N_1122,In_276,In_93);
nand U1123 (N_1123,In_1336,In_526);
or U1124 (N_1124,In_1491,In_1302);
nand U1125 (N_1125,In_150,In_814);
nand U1126 (N_1126,In_1413,In_582);
nand U1127 (N_1127,In_1364,In_283);
or U1128 (N_1128,In_505,In_320);
or U1129 (N_1129,In_1420,In_913);
nor U1130 (N_1130,In_1074,In_514);
or U1131 (N_1131,In_472,In_541);
nor U1132 (N_1132,In_739,In_806);
nand U1133 (N_1133,In_1132,In_1006);
nand U1134 (N_1134,In_135,In_28);
or U1135 (N_1135,In_79,In_1071);
nand U1136 (N_1136,In_9,In_81);
nand U1137 (N_1137,In_191,In_156);
or U1138 (N_1138,In_757,In_227);
or U1139 (N_1139,In_490,In_1004);
or U1140 (N_1140,In_853,In_518);
and U1141 (N_1141,In_1331,In_804);
nand U1142 (N_1142,In_1081,In_218);
nor U1143 (N_1143,In_240,In_1335);
or U1144 (N_1144,In_882,In_94);
and U1145 (N_1145,In_423,In_291);
or U1146 (N_1146,In_328,In_809);
xor U1147 (N_1147,In_1496,In_1105);
nor U1148 (N_1148,In_1375,In_1159);
or U1149 (N_1149,In_897,In_547);
xnor U1150 (N_1150,In_883,In_704);
and U1151 (N_1151,In_1117,In_114);
nand U1152 (N_1152,In_1372,In_1354);
nor U1153 (N_1153,In_1212,In_1374);
nand U1154 (N_1154,In_118,In_321);
nand U1155 (N_1155,In_157,In_715);
and U1156 (N_1156,In_1179,In_525);
and U1157 (N_1157,In_712,In_547);
nand U1158 (N_1158,In_1072,In_713);
xnor U1159 (N_1159,In_310,In_846);
nor U1160 (N_1160,In_1082,In_182);
or U1161 (N_1161,In_1121,In_309);
nor U1162 (N_1162,In_675,In_1054);
xor U1163 (N_1163,In_821,In_1064);
or U1164 (N_1164,In_30,In_718);
nor U1165 (N_1165,In_39,In_613);
and U1166 (N_1166,In_302,In_942);
and U1167 (N_1167,In_483,In_1425);
nand U1168 (N_1168,In_827,In_700);
nand U1169 (N_1169,In_257,In_1357);
and U1170 (N_1170,In_1098,In_1199);
or U1171 (N_1171,In_1316,In_1147);
nor U1172 (N_1172,In_161,In_1150);
and U1173 (N_1173,In_1210,In_869);
and U1174 (N_1174,In_1488,In_1459);
or U1175 (N_1175,In_1488,In_1291);
nor U1176 (N_1176,In_658,In_1338);
xnor U1177 (N_1177,In_900,In_1130);
and U1178 (N_1178,In_3,In_1245);
and U1179 (N_1179,In_83,In_330);
nor U1180 (N_1180,In_544,In_538);
and U1181 (N_1181,In_1336,In_684);
nor U1182 (N_1182,In_235,In_601);
nor U1183 (N_1183,In_820,In_551);
nor U1184 (N_1184,In_1478,In_993);
and U1185 (N_1185,In_318,In_1066);
nor U1186 (N_1186,In_1381,In_792);
xnor U1187 (N_1187,In_663,In_184);
nand U1188 (N_1188,In_121,In_1264);
or U1189 (N_1189,In_807,In_342);
nor U1190 (N_1190,In_805,In_1386);
nor U1191 (N_1191,In_611,In_420);
nor U1192 (N_1192,In_668,In_154);
nor U1193 (N_1193,In_1429,In_736);
nand U1194 (N_1194,In_621,In_1215);
nand U1195 (N_1195,In_1497,In_569);
or U1196 (N_1196,In_245,In_947);
nand U1197 (N_1197,In_27,In_899);
nand U1198 (N_1198,In_1003,In_1056);
and U1199 (N_1199,In_293,In_458);
and U1200 (N_1200,In_415,In_269);
nor U1201 (N_1201,In_452,In_1383);
or U1202 (N_1202,In_423,In_767);
nand U1203 (N_1203,In_90,In_466);
or U1204 (N_1204,In_416,In_1070);
nand U1205 (N_1205,In_453,In_661);
and U1206 (N_1206,In_688,In_499);
nand U1207 (N_1207,In_996,In_417);
and U1208 (N_1208,In_1178,In_260);
or U1209 (N_1209,In_664,In_442);
or U1210 (N_1210,In_1378,In_655);
and U1211 (N_1211,In_366,In_1016);
nand U1212 (N_1212,In_1236,In_882);
and U1213 (N_1213,In_756,In_710);
nor U1214 (N_1214,In_341,In_1249);
nor U1215 (N_1215,In_1001,In_302);
and U1216 (N_1216,In_773,In_105);
nand U1217 (N_1217,In_174,In_349);
nand U1218 (N_1218,In_1148,In_1354);
nor U1219 (N_1219,In_526,In_1140);
nand U1220 (N_1220,In_813,In_1244);
and U1221 (N_1221,In_1042,In_1070);
or U1222 (N_1222,In_620,In_760);
or U1223 (N_1223,In_834,In_1028);
nand U1224 (N_1224,In_1285,In_677);
and U1225 (N_1225,In_145,In_537);
xnor U1226 (N_1226,In_350,In_629);
nand U1227 (N_1227,In_677,In_685);
nand U1228 (N_1228,In_674,In_187);
nor U1229 (N_1229,In_199,In_728);
nor U1230 (N_1230,In_1066,In_377);
xnor U1231 (N_1231,In_1023,In_354);
and U1232 (N_1232,In_1441,In_431);
nor U1233 (N_1233,In_777,In_313);
nor U1234 (N_1234,In_686,In_1400);
nand U1235 (N_1235,In_1355,In_832);
nand U1236 (N_1236,In_353,In_536);
nor U1237 (N_1237,In_668,In_1438);
nand U1238 (N_1238,In_337,In_688);
nand U1239 (N_1239,In_1188,In_238);
and U1240 (N_1240,In_943,In_149);
nor U1241 (N_1241,In_1404,In_541);
or U1242 (N_1242,In_1128,In_1024);
nor U1243 (N_1243,In_1454,In_660);
nor U1244 (N_1244,In_262,In_36);
nor U1245 (N_1245,In_296,In_1046);
or U1246 (N_1246,In_1437,In_1272);
xor U1247 (N_1247,In_690,In_1063);
or U1248 (N_1248,In_575,In_996);
nand U1249 (N_1249,In_1218,In_162);
or U1250 (N_1250,In_450,In_43);
nor U1251 (N_1251,In_534,In_632);
or U1252 (N_1252,In_1340,In_289);
nor U1253 (N_1253,In_1454,In_242);
nand U1254 (N_1254,In_1103,In_346);
xnor U1255 (N_1255,In_607,In_729);
or U1256 (N_1256,In_516,In_67);
xnor U1257 (N_1257,In_1144,In_499);
or U1258 (N_1258,In_190,In_1275);
and U1259 (N_1259,In_539,In_768);
nor U1260 (N_1260,In_17,In_601);
or U1261 (N_1261,In_1355,In_215);
or U1262 (N_1262,In_252,In_741);
nand U1263 (N_1263,In_578,In_1317);
or U1264 (N_1264,In_633,In_863);
nor U1265 (N_1265,In_163,In_918);
xnor U1266 (N_1266,In_1316,In_769);
or U1267 (N_1267,In_446,In_1451);
xnor U1268 (N_1268,In_1327,In_4);
nor U1269 (N_1269,In_583,In_225);
nor U1270 (N_1270,In_439,In_968);
and U1271 (N_1271,In_804,In_857);
nor U1272 (N_1272,In_1079,In_1176);
or U1273 (N_1273,In_52,In_531);
nor U1274 (N_1274,In_802,In_1244);
or U1275 (N_1275,In_933,In_1276);
or U1276 (N_1276,In_1456,In_1202);
nor U1277 (N_1277,In_561,In_1097);
nor U1278 (N_1278,In_876,In_907);
and U1279 (N_1279,In_467,In_889);
nor U1280 (N_1280,In_359,In_1285);
nand U1281 (N_1281,In_591,In_165);
and U1282 (N_1282,In_1042,In_464);
nor U1283 (N_1283,In_344,In_490);
nor U1284 (N_1284,In_778,In_1196);
nor U1285 (N_1285,In_508,In_1141);
nand U1286 (N_1286,In_651,In_1276);
xor U1287 (N_1287,In_253,In_884);
nor U1288 (N_1288,In_1138,In_285);
nor U1289 (N_1289,In_1321,In_943);
or U1290 (N_1290,In_630,In_1111);
or U1291 (N_1291,In_636,In_934);
nand U1292 (N_1292,In_1432,In_1453);
xor U1293 (N_1293,In_925,In_1416);
xnor U1294 (N_1294,In_392,In_368);
nand U1295 (N_1295,In_450,In_733);
nand U1296 (N_1296,In_196,In_1461);
nor U1297 (N_1297,In_129,In_1128);
and U1298 (N_1298,In_71,In_773);
and U1299 (N_1299,In_535,In_945);
or U1300 (N_1300,In_106,In_1010);
nand U1301 (N_1301,In_944,In_940);
or U1302 (N_1302,In_1272,In_1339);
nor U1303 (N_1303,In_824,In_735);
xor U1304 (N_1304,In_775,In_957);
or U1305 (N_1305,In_1147,In_1180);
and U1306 (N_1306,In_121,In_1246);
or U1307 (N_1307,In_17,In_406);
nand U1308 (N_1308,In_1129,In_857);
or U1309 (N_1309,In_462,In_1114);
or U1310 (N_1310,In_701,In_1348);
and U1311 (N_1311,In_1416,In_152);
and U1312 (N_1312,In_1208,In_1393);
nor U1313 (N_1313,In_1444,In_379);
nor U1314 (N_1314,In_396,In_988);
nand U1315 (N_1315,In_21,In_1049);
nand U1316 (N_1316,In_119,In_1019);
nor U1317 (N_1317,In_922,In_25);
nor U1318 (N_1318,In_433,In_1350);
nand U1319 (N_1319,In_641,In_680);
nor U1320 (N_1320,In_191,In_110);
or U1321 (N_1321,In_542,In_203);
xnor U1322 (N_1322,In_1069,In_214);
nand U1323 (N_1323,In_634,In_442);
and U1324 (N_1324,In_23,In_1301);
xor U1325 (N_1325,In_360,In_795);
and U1326 (N_1326,In_1417,In_412);
and U1327 (N_1327,In_1095,In_926);
nand U1328 (N_1328,In_384,In_38);
nor U1329 (N_1329,In_616,In_323);
and U1330 (N_1330,In_136,In_57);
or U1331 (N_1331,In_162,In_1432);
or U1332 (N_1332,In_141,In_521);
nand U1333 (N_1333,In_469,In_100);
nand U1334 (N_1334,In_942,In_1439);
xnor U1335 (N_1335,In_1457,In_522);
and U1336 (N_1336,In_587,In_1265);
and U1337 (N_1337,In_547,In_685);
and U1338 (N_1338,In_678,In_515);
nor U1339 (N_1339,In_246,In_589);
nor U1340 (N_1340,In_1080,In_615);
xor U1341 (N_1341,In_1343,In_1077);
nand U1342 (N_1342,In_1410,In_982);
and U1343 (N_1343,In_292,In_597);
xnor U1344 (N_1344,In_1038,In_931);
or U1345 (N_1345,In_1117,In_215);
or U1346 (N_1346,In_1403,In_1016);
and U1347 (N_1347,In_1110,In_683);
nor U1348 (N_1348,In_743,In_493);
and U1349 (N_1349,In_1044,In_413);
xor U1350 (N_1350,In_1173,In_290);
xor U1351 (N_1351,In_1040,In_754);
and U1352 (N_1352,In_464,In_1379);
nor U1353 (N_1353,In_1465,In_1327);
or U1354 (N_1354,In_815,In_1027);
nor U1355 (N_1355,In_425,In_796);
and U1356 (N_1356,In_1157,In_92);
and U1357 (N_1357,In_422,In_48);
nor U1358 (N_1358,In_960,In_15);
and U1359 (N_1359,In_742,In_1283);
or U1360 (N_1360,In_624,In_539);
or U1361 (N_1361,In_733,In_465);
or U1362 (N_1362,In_596,In_1341);
or U1363 (N_1363,In_794,In_629);
or U1364 (N_1364,In_691,In_749);
and U1365 (N_1365,In_395,In_1069);
nand U1366 (N_1366,In_1247,In_1191);
nand U1367 (N_1367,In_336,In_687);
nor U1368 (N_1368,In_1380,In_1239);
or U1369 (N_1369,In_991,In_454);
and U1370 (N_1370,In_277,In_1314);
or U1371 (N_1371,In_1187,In_1329);
and U1372 (N_1372,In_679,In_949);
nor U1373 (N_1373,In_505,In_917);
or U1374 (N_1374,In_1342,In_774);
and U1375 (N_1375,In_727,In_903);
and U1376 (N_1376,In_1216,In_472);
nor U1377 (N_1377,In_903,In_1234);
nand U1378 (N_1378,In_1404,In_736);
or U1379 (N_1379,In_1184,In_903);
or U1380 (N_1380,In_1249,In_1268);
nor U1381 (N_1381,In_24,In_806);
nand U1382 (N_1382,In_1183,In_770);
and U1383 (N_1383,In_456,In_452);
nand U1384 (N_1384,In_1279,In_395);
nand U1385 (N_1385,In_1233,In_756);
xnor U1386 (N_1386,In_1182,In_864);
nand U1387 (N_1387,In_506,In_224);
or U1388 (N_1388,In_241,In_1330);
and U1389 (N_1389,In_1049,In_12);
nand U1390 (N_1390,In_682,In_101);
nand U1391 (N_1391,In_1438,In_455);
nand U1392 (N_1392,In_1305,In_1461);
nand U1393 (N_1393,In_596,In_852);
or U1394 (N_1394,In_1010,In_883);
or U1395 (N_1395,In_543,In_22);
or U1396 (N_1396,In_1376,In_1474);
xor U1397 (N_1397,In_1379,In_745);
or U1398 (N_1398,In_1278,In_241);
nor U1399 (N_1399,In_910,In_321);
xnor U1400 (N_1400,In_1092,In_1356);
nand U1401 (N_1401,In_838,In_9);
or U1402 (N_1402,In_855,In_256);
nand U1403 (N_1403,In_275,In_330);
nand U1404 (N_1404,In_989,In_139);
nor U1405 (N_1405,In_1330,In_1084);
and U1406 (N_1406,In_874,In_301);
nor U1407 (N_1407,In_1439,In_1009);
and U1408 (N_1408,In_830,In_321);
nand U1409 (N_1409,In_9,In_1430);
or U1410 (N_1410,In_157,In_1194);
nor U1411 (N_1411,In_482,In_428);
or U1412 (N_1412,In_1430,In_1492);
nor U1413 (N_1413,In_196,In_580);
and U1414 (N_1414,In_1223,In_958);
nor U1415 (N_1415,In_1121,In_477);
or U1416 (N_1416,In_533,In_591);
and U1417 (N_1417,In_266,In_1464);
nand U1418 (N_1418,In_799,In_425);
or U1419 (N_1419,In_1458,In_267);
xor U1420 (N_1420,In_193,In_972);
and U1421 (N_1421,In_602,In_1235);
nor U1422 (N_1422,In_170,In_1140);
and U1423 (N_1423,In_112,In_464);
xor U1424 (N_1424,In_150,In_944);
nand U1425 (N_1425,In_1303,In_104);
and U1426 (N_1426,In_1225,In_1036);
or U1427 (N_1427,In_668,In_60);
xnor U1428 (N_1428,In_1400,In_156);
or U1429 (N_1429,In_726,In_1244);
nor U1430 (N_1430,In_358,In_960);
nor U1431 (N_1431,In_1034,In_313);
nand U1432 (N_1432,In_219,In_858);
nor U1433 (N_1433,In_910,In_691);
or U1434 (N_1434,In_823,In_920);
and U1435 (N_1435,In_565,In_1073);
nor U1436 (N_1436,In_1409,In_531);
nand U1437 (N_1437,In_627,In_98);
nand U1438 (N_1438,In_124,In_1369);
or U1439 (N_1439,In_237,In_912);
nor U1440 (N_1440,In_1165,In_554);
or U1441 (N_1441,In_95,In_499);
and U1442 (N_1442,In_835,In_298);
nand U1443 (N_1443,In_1283,In_412);
nor U1444 (N_1444,In_202,In_279);
and U1445 (N_1445,In_665,In_566);
or U1446 (N_1446,In_1205,In_1438);
nand U1447 (N_1447,In_1126,In_451);
xor U1448 (N_1448,In_651,In_426);
nor U1449 (N_1449,In_1009,In_1199);
or U1450 (N_1450,In_561,In_264);
nand U1451 (N_1451,In_1032,In_271);
or U1452 (N_1452,In_358,In_621);
or U1453 (N_1453,In_341,In_1065);
xor U1454 (N_1454,In_295,In_338);
nor U1455 (N_1455,In_823,In_721);
xor U1456 (N_1456,In_421,In_601);
and U1457 (N_1457,In_1114,In_111);
or U1458 (N_1458,In_358,In_981);
and U1459 (N_1459,In_329,In_1310);
and U1460 (N_1460,In_1495,In_82);
nand U1461 (N_1461,In_905,In_275);
and U1462 (N_1462,In_1318,In_714);
nand U1463 (N_1463,In_1405,In_577);
nand U1464 (N_1464,In_34,In_48);
and U1465 (N_1465,In_76,In_871);
nor U1466 (N_1466,In_1286,In_329);
and U1467 (N_1467,In_185,In_282);
or U1468 (N_1468,In_783,In_785);
or U1469 (N_1469,In_924,In_210);
and U1470 (N_1470,In_18,In_262);
nand U1471 (N_1471,In_290,In_574);
and U1472 (N_1472,In_1427,In_176);
nand U1473 (N_1473,In_249,In_88);
and U1474 (N_1474,In_256,In_789);
nor U1475 (N_1475,In_85,In_283);
xnor U1476 (N_1476,In_1207,In_1121);
xor U1477 (N_1477,In_880,In_1390);
nor U1478 (N_1478,In_900,In_656);
xor U1479 (N_1479,In_347,In_818);
or U1480 (N_1480,In_235,In_746);
and U1481 (N_1481,In_1235,In_1141);
or U1482 (N_1482,In_911,In_671);
nand U1483 (N_1483,In_1420,In_138);
nand U1484 (N_1484,In_595,In_635);
nand U1485 (N_1485,In_33,In_1291);
and U1486 (N_1486,In_447,In_1047);
xnor U1487 (N_1487,In_437,In_527);
nand U1488 (N_1488,In_202,In_10);
and U1489 (N_1489,In_998,In_943);
nor U1490 (N_1490,In_530,In_515);
and U1491 (N_1491,In_207,In_233);
or U1492 (N_1492,In_1445,In_163);
xnor U1493 (N_1493,In_125,In_448);
or U1494 (N_1494,In_1450,In_468);
nand U1495 (N_1495,In_278,In_1455);
nor U1496 (N_1496,In_1210,In_627);
nand U1497 (N_1497,In_537,In_1194);
and U1498 (N_1498,In_848,In_1485);
nand U1499 (N_1499,In_678,In_777);
xnor U1500 (N_1500,In_1076,In_196);
xnor U1501 (N_1501,In_1009,In_1303);
nand U1502 (N_1502,In_297,In_490);
xor U1503 (N_1503,In_273,In_1144);
and U1504 (N_1504,In_1145,In_1012);
nand U1505 (N_1505,In_385,In_48);
nor U1506 (N_1506,In_1205,In_1287);
nor U1507 (N_1507,In_1240,In_1433);
nand U1508 (N_1508,In_1368,In_118);
nor U1509 (N_1509,In_418,In_1324);
nor U1510 (N_1510,In_1229,In_1317);
xnor U1511 (N_1511,In_1413,In_474);
nand U1512 (N_1512,In_123,In_190);
nor U1513 (N_1513,In_1376,In_283);
nand U1514 (N_1514,In_219,In_438);
or U1515 (N_1515,In_884,In_1292);
and U1516 (N_1516,In_1368,In_409);
or U1517 (N_1517,In_1032,In_1348);
nand U1518 (N_1518,In_593,In_43);
nand U1519 (N_1519,In_213,In_1312);
or U1520 (N_1520,In_663,In_987);
nand U1521 (N_1521,In_1007,In_713);
xor U1522 (N_1522,In_1277,In_912);
nand U1523 (N_1523,In_1049,In_59);
nand U1524 (N_1524,In_125,In_1128);
xor U1525 (N_1525,In_366,In_1285);
nand U1526 (N_1526,In_253,In_1175);
and U1527 (N_1527,In_1386,In_1007);
nor U1528 (N_1528,In_953,In_1367);
or U1529 (N_1529,In_1395,In_355);
nand U1530 (N_1530,In_925,In_600);
xor U1531 (N_1531,In_1356,In_70);
nand U1532 (N_1532,In_523,In_752);
nand U1533 (N_1533,In_1317,In_193);
and U1534 (N_1534,In_845,In_654);
nor U1535 (N_1535,In_325,In_1247);
and U1536 (N_1536,In_583,In_1324);
nor U1537 (N_1537,In_150,In_1213);
nor U1538 (N_1538,In_173,In_1199);
and U1539 (N_1539,In_784,In_706);
or U1540 (N_1540,In_1017,In_904);
nor U1541 (N_1541,In_389,In_1201);
and U1542 (N_1542,In_519,In_1053);
nand U1543 (N_1543,In_531,In_1144);
nand U1544 (N_1544,In_1025,In_1080);
and U1545 (N_1545,In_460,In_1189);
xor U1546 (N_1546,In_1172,In_1320);
or U1547 (N_1547,In_1182,In_41);
nor U1548 (N_1548,In_81,In_1271);
nand U1549 (N_1549,In_169,In_538);
and U1550 (N_1550,In_850,In_206);
nand U1551 (N_1551,In_238,In_466);
and U1552 (N_1552,In_26,In_379);
or U1553 (N_1553,In_584,In_388);
xor U1554 (N_1554,In_947,In_1455);
or U1555 (N_1555,In_1440,In_877);
nand U1556 (N_1556,In_728,In_1322);
and U1557 (N_1557,In_1379,In_433);
xnor U1558 (N_1558,In_754,In_574);
xor U1559 (N_1559,In_616,In_1105);
xor U1560 (N_1560,In_672,In_995);
nor U1561 (N_1561,In_135,In_6);
xnor U1562 (N_1562,In_1012,In_47);
nand U1563 (N_1563,In_1099,In_40);
nor U1564 (N_1564,In_807,In_821);
or U1565 (N_1565,In_1494,In_1459);
nor U1566 (N_1566,In_742,In_834);
or U1567 (N_1567,In_1443,In_1142);
nor U1568 (N_1568,In_1098,In_137);
nor U1569 (N_1569,In_478,In_1201);
or U1570 (N_1570,In_504,In_640);
nor U1571 (N_1571,In_1450,In_71);
nand U1572 (N_1572,In_1103,In_115);
nor U1573 (N_1573,In_1203,In_1116);
nor U1574 (N_1574,In_1043,In_1486);
nand U1575 (N_1575,In_975,In_903);
or U1576 (N_1576,In_1097,In_1155);
xor U1577 (N_1577,In_663,In_1418);
and U1578 (N_1578,In_42,In_1003);
or U1579 (N_1579,In_965,In_924);
nand U1580 (N_1580,In_1251,In_1261);
xor U1581 (N_1581,In_410,In_1075);
and U1582 (N_1582,In_1458,In_105);
nand U1583 (N_1583,In_1497,In_1461);
nor U1584 (N_1584,In_1487,In_1414);
and U1585 (N_1585,In_928,In_562);
and U1586 (N_1586,In_469,In_1111);
or U1587 (N_1587,In_367,In_993);
nor U1588 (N_1588,In_6,In_471);
or U1589 (N_1589,In_614,In_736);
or U1590 (N_1590,In_536,In_1131);
nor U1591 (N_1591,In_459,In_1022);
nand U1592 (N_1592,In_1123,In_1070);
nand U1593 (N_1593,In_625,In_126);
nand U1594 (N_1594,In_1477,In_667);
nand U1595 (N_1595,In_641,In_1288);
or U1596 (N_1596,In_790,In_276);
nor U1597 (N_1597,In_192,In_280);
and U1598 (N_1598,In_1108,In_1186);
nand U1599 (N_1599,In_77,In_607);
nand U1600 (N_1600,In_102,In_7);
or U1601 (N_1601,In_983,In_1164);
nor U1602 (N_1602,In_1244,In_450);
nand U1603 (N_1603,In_1496,In_304);
xnor U1604 (N_1604,In_1064,In_527);
or U1605 (N_1605,In_301,In_1046);
nand U1606 (N_1606,In_1041,In_831);
nand U1607 (N_1607,In_452,In_118);
nor U1608 (N_1608,In_336,In_660);
or U1609 (N_1609,In_592,In_700);
nand U1610 (N_1610,In_111,In_704);
nand U1611 (N_1611,In_117,In_1399);
or U1612 (N_1612,In_216,In_1133);
xor U1613 (N_1613,In_98,In_884);
nand U1614 (N_1614,In_1435,In_508);
nor U1615 (N_1615,In_1476,In_855);
xnor U1616 (N_1616,In_1357,In_1456);
or U1617 (N_1617,In_654,In_331);
nor U1618 (N_1618,In_1239,In_961);
xor U1619 (N_1619,In_483,In_572);
and U1620 (N_1620,In_1120,In_706);
nor U1621 (N_1621,In_1175,In_167);
nor U1622 (N_1622,In_852,In_50);
and U1623 (N_1623,In_1435,In_723);
xnor U1624 (N_1624,In_1052,In_237);
and U1625 (N_1625,In_72,In_591);
xnor U1626 (N_1626,In_390,In_672);
or U1627 (N_1627,In_1175,In_1417);
and U1628 (N_1628,In_398,In_623);
nand U1629 (N_1629,In_414,In_1205);
and U1630 (N_1630,In_1442,In_9);
nand U1631 (N_1631,In_770,In_710);
nor U1632 (N_1632,In_1297,In_616);
nand U1633 (N_1633,In_153,In_45);
nand U1634 (N_1634,In_28,In_544);
nand U1635 (N_1635,In_1100,In_1000);
nand U1636 (N_1636,In_635,In_1348);
and U1637 (N_1637,In_1176,In_323);
nand U1638 (N_1638,In_1057,In_1029);
nand U1639 (N_1639,In_1361,In_600);
xor U1640 (N_1640,In_187,In_605);
and U1641 (N_1641,In_1310,In_562);
or U1642 (N_1642,In_38,In_631);
xnor U1643 (N_1643,In_794,In_1470);
or U1644 (N_1644,In_1106,In_379);
xor U1645 (N_1645,In_678,In_215);
nor U1646 (N_1646,In_1354,In_971);
or U1647 (N_1647,In_700,In_573);
nor U1648 (N_1648,In_92,In_293);
nand U1649 (N_1649,In_720,In_748);
and U1650 (N_1650,In_381,In_1183);
nor U1651 (N_1651,In_769,In_877);
or U1652 (N_1652,In_71,In_1122);
or U1653 (N_1653,In_215,In_457);
nand U1654 (N_1654,In_903,In_1243);
nand U1655 (N_1655,In_457,In_96);
and U1656 (N_1656,In_16,In_1443);
and U1657 (N_1657,In_1271,In_851);
nand U1658 (N_1658,In_447,In_274);
and U1659 (N_1659,In_821,In_554);
nand U1660 (N_1660,In_1061,In_444);
and U1661 (N_1661,In_1067,In_1043);
nand U1662 (N_1662,In_107,In_884);
and U1663 (N_1663,In_890,In_653);
nand U1664 (N_1664,In_1486,In_824);
and U1665 (N_1665,In_108,In_983);
and U1666 (N_1666,In_645,In_1096);
xor U1667 (N_1667,In_1,In_764);
and U1668 (N_1668,In_1156,In_1363);
or U1669 (N_1669,In_52,In_560);
or U1670 (N_1670,In_1454,In_475);
nor U1671 (N_1671,In_661,In_698);
and U1672 (N_1672,In_763,In_722);
nand U1673 (N_1673,In_81,In_900);
nor U1674 (N_1674,In_1316,In_1344);
nor U1675 (N_1675,In_720,In_1276);
and U1676 (N_1676,In_13,In_869);
nor U1677 (N_1677,In_417,In_595);
and U1678 (N_1678,In_553,In_1372);
and U1679 (N_1679,In_362,In_1366);
xor U1680 (N_1680,In_343,In_438);
and U1681 (N_1681,In_390,In_149);
or U1682 (N_1682,In_1182,In_445);
nand U1683 (N_1683,In_913,In_100);
nand U1684 (N_1684,In_717,In_537);
and U1685 (N_1685,In_878,In_1439);
or U1686 (N_1686,In_725,In_481);
or U1687 (N_1687,In_1149,In_690);
nor U1688 (N_1688,In_1382,In_1012);
or U1689 (N_1689,In_511,In_1215);
nand U1690 (N_1690,In_259,In_1419);
and U1691 (N_1691,In_656,In_961);
and U1692 (N_1692,In_1269,In_249);
and U1693 (N_1693,In_978,In_1209);
nand U1694 (N_1694,In_701,In_378);
and U1695 (N_1695,In_358,In_133);
and U1696 (N_1696,In_183,In_136);
and U1697 (N_1697,In_1092,In_1123);
nor U1698 (N_1698,In_521,In_924);
and U1699 (N_1699,In_1108,In_449);
nand U1700 (N_1700,In_904,In_1202);
xnor U1701 (N_1701,In_13,In_880);
xnor U1702 (N_1702,In_248,In_547);
nand U1703 (N_1703,In_333,In_878);
and U1704 (N_1704,In_913,In_423);
and U1705 (N_1705,In_1144,In_1035);
or U1706 (N_1706,In_950,In_1058);
and U1707 (N_1707,In_713,In_33);
xnor U1708 (N_1708,In_535,In_1260);
or U1709 (N_1709,In_95,In_915);
nor U1710 (N_1710,In_466,In_375);
nand U1711 (N_1711,In_993,In_1100);
and U1712 (N_1712,In_949,In_933);
nor U1713 (N_1713,In_1387,In_13);
or U1714 (N_1714,In_590,In_1462);
nor U1715 (N_1715,In_333,In_1022);
or U1716 (N_1716,In_38,In_1003);
or U1717 (N_1717,In_1140,In_1451);
nor U1718 (N_1718,In_466,In_44);
xor U1719 (N_1719,In_269,In_839);
nand U1720 (N_1720,In_3,In_980);
nand U1721 (N_1721,In_668,In_1168);
nor U1722 (N_1722,In_486,In_677);
and U1723 (N_1723,In_1035,In_307);
or U1724 (N_1724,In_787,In_73);
nor U1725 (N_1725,In_1337,In_1008);
or U1726 (N_1726,In_568,In_1256);
nand U1727 (N_1727,In_244,In_848);
and U1728 (N_1728,In_687,In_243);
or U1729 (N_1729,In_1150,In_244);
xnor U1730 (N_1730,In_841,In_537);
and U1731 (N_1731,In_754,In_1171);
and U1732 (N_1732,In_1157,In_570);
or U1733 (N_1733,In_997,In_1324);
and U1734 (N_1734,In_720,In_1025);
nor U1735 (N_1735,In_1283,In_1322);
and U1736 (N_1736,In_999,In_542);
nor U1737 (N_1737,In_1035,In_1086);
and U1738 (N_1738,In_152,In_606);
and U1739 (N_1739,In_452,In_48);
nor U1740 (N_1740,In_559,In_210);
nand U1741 (N_1741,In_123,In_1364);
nor U1742 (N_1742,In_329,In_817);
and U1743 (N_1743,In_298,In_573);
or U1744 (N_1744,In_1367,In_372);
or U1745 (N_1745,In_1111,In_1142);
or U1746 (N_1746,In_674,In_915);
and U1747 (N_1747,In_762,In_730);
nor U1748 (N_1748,In_216,In_1376);
nand U1749 (N_1749,In_1449,In_850);
and U1750 (N_1750,In_562,In_1001);
and U1751 (N_1751,In_1015,In_89);
nand U1752 (N_1752,In_746,In_1315);
and U1753 (N_1753,In_623,In_476);
nand U1754 (N_1754,In_1410,In_811);
nand U1755 (N_1755,In_1253,In_1398);
and U1756 (N_1756,In_275,In_1111);
nand U1757 (N_1757,In_492,In_944);
or U1758 (N_1758,In_208,In_883);
nor U1759 (N_1759,In_1474,In_1160);
nor U1760 (N_1760,In_1444,In_1365);
nand U1761 (N_1761,In_1201,In_1455);
or U1762 (N_1762,In_537,In_824);
xnor U1763 (N_1763,In_1246,In_879);
or U1764 (N_1764,In_1120,In_779);
nand U1765 (N_1765,In_718,In_564);
and U1766 (N_1766,In_786,In_623);
and U1767 (N_1767,In_209,In_736);
or U1768 (N_1768,In_1227,In_476);
nand U1769 (N_1769,In_816,In_1373);
and U1770 (N_1770,In_702,In_272);
nand U1771 (N_1771,In_133,In_946);
or U1772 (N_1772,In_689,In_1066);
or U1773 (N_1773,In_966,In_655);
nor U1774 (N_1774,In_1344,In_524);
or U1775 (N_1775,In_1449,In_1045);
or U1776 (N_1776,In_898,In_1144);
nor U1777 (N_1777,In_545,In_943);
nand U1778 (N_1778,In_1048,In_1096);
and U1779 (N_1779,In_274,In_1350);
nor U1780 (N_1780,In_549,In_711);
nor U1781 (N_1781,In_45,In_1321);
and U1782 (N_1782,In_158,In_859);
nor U1783 (N_1783,In_1267,In_1263);
nor U1784 (N_1784,In_279,In_1065);
and U1785 (N_1785,In_1314,In_1373);
nand U1786 (N_1786,In_255,In_1402);
xnor U1787 (N_1787,In_262,In_1163);
or U1788 (N_1788,In_862,In_890);
nor U1789 (N_1789,In_901,In_226);
nor U1790 (N_1790,In_937,In_1018);
and U1791 (N_1791,In_5,In_517);
and U1792 (N_1792,In_711,In_1096);
nor U1793 (N_1793,In_1308,In_210);
nand U1794 (N_1794,In_310,In_87);
and U1795 (N_1795,In_577,In_695);
nand U1796 (N_1796,In_1244,In_1196);
nor U1797 (N_1797,In_396,In_156);
and U1798 (N_1798,In_270,In_435);
and U1799 (N_1799,In_505,In_97);
and U1800 (N_1800,In_169,In_1482);
nand U1801 (N_1801,In_826,In_234);
and U1802 (N_1802,In_919,In_1363);
nor U1803 (N_1803,In_388,In_519);
nor U1804 (N_1804,In_232,In_10);
nand U1805 (N_1805,In_1477,In_274);
nand U1806 (N_1806,In_1346,In_985);
or U1807 (N_1807,In_319,In_331);
or U1808 (N_1808,In_439,In_480);
nand U1809 (N_1809,In_717,In_81);
or U1810 (N_1810,In_1087,In_449);
nand U1811 (N_1811,In_108,In_1484);
and U1812 (N_1812,In_916,In_1466);
or U1813 (N_1813,In_692,In_1014);
nand U1814 (N_1814,In_743,In_317);
or U1815 (N_1815,In_8,In_1361);
nor U1816 (N_1816,In_1382,In_787);
nand U1817 (N_1817,In_607,In_1081);
nor U1818 (N_1818,In_205,In_210);
and U1819 (N_1819,In_963,In_515);
nor U1820 (N_1820,In_1211,In_45);
and U1821 (N_1821,In_1300,In_1486);
and U1822 (N_1822,In_977,In_700);
and U1823 (N_1823,In_77,In_318);
or U1824 (N_1824,In_1144,In_164);
xor U1825 (N_1825,In_30,In_482);
nor U1826 (N_1826,In_356,In_1100);
and U1827 (N_1827,In_1171,In_1221);
nand U1828 (N_1828,In_568,In_64);
xor U1829 (N_1829,In_236,In_76);
and U1830 (N_1830,In_664,In_425);
nand U1831 (N_1831,In_856,In_415);
xor U1832 (N_1832,In_1075,In_1260);
xnor U1833 (N_1833,In_520,In_166);
nor U1834 (N_1834,In_1002,In_510);
xnor U1835 (N_1835,In_79,In_1398);
nand U1836 (N_1836,In_1406,In_469);
xor U1837 (N_1837,In_449,In_1003);
nor U1838 (N_1838,In_75,In_873);
xnor U1839 (N_1839,In_401,In_1494);
nor U1840 (N_1840,In_1412,In_29);
nand U1841 (N_1841,In_604,In_724);
or U1842 (N_1842,In_102,In_243);
and U1843 (N_1843,In_1136,In_1482);
or U1844 (N_1844,In_299,In_347);
nand U1845 (N_1845,In_85,In_684);
and U1846 (N_1846,In_477,In_1231);
or U1847 (N_1847,In_1431,In_1424);
nor U1848 (N_1848,In_1083,In_967);
or U1849 (N_1849,In_590,In_1104);
or U1850 (N_1850,In_122,In_1365);
or U1851 (N_1851,In_1086,In_364);
nand U1852 (N_1852,In_280,In_243);
xor U1853 (N_1853,In_1382,In_36);
or U1854 (N_1854,In_850,In_1418);
and U1855 (N_1855,In_592,In_1390);
xor U1856 (N_1856,In_27,In_878);
xor U1857 (N_1857,In_266,In_1395);
and U1858 (N_1858,In_507,In_250);
nand U1859 (N_1859,In_83,In_1344);
nand U1860 (N_1860,In_71,In_575);
or U1861 (N_1861,In_54,In_126);
nor U1862 (N_1862,In_235,In_388);
nor U1863 (N_1863,In_204,In_1008);
nor U1864 (N_1864,In_470,In_26);
xor U1865 (N_1865,In_1230,In_416);
and U1866 (N_1866,In_1062,In_1180);
and U1867 (N_1867,In_33,In_510);
and U1868 (N_1868,In_496,In_250);
xor U1869 (N_1869,In_755,In_1);
nor U1870 (N_1870,In_573,In_714);
or U1871 (N_1871,In_396,In_1037);
or U1872 (N_1872,In_141,In_517);
nor U1873 (N_1873,In_1177,In_59);
and U1874 (N_1874,In_1398,In_553);
and U1875 (N_1875,In_108,In_1291);
nor U1876 (N_1876,In_367,In_462);
nor U1877 (N_1877,In_496,In_1121);
or U1878 (N_1878,In_671,In_1350);
nand U1879 (N_1879,In_697,In_1395);
xor U1880 (N_1880,In_912,In_855);
and U1881 (N_1881,In_233,In_1069);
and U1882 (N_1882,In_1245,In_338);
and U1883 (N_1883,In_510,In_1443);
nand U1884 (N_1884,In_1210,In_398);
or U1885 (N_1885,In_1375,In_1463);
or U1886 (N_1886,In_167,In_259);
nor U1887 (N_1887,In_417,In_186);
and U1888 (N_1888,In_882,In_243);
nor U1889 (N_1889,In_773,In_364);
nor U1890 (N_1890,In_1059,In_1176);
nand U1891 (N_1891,In_581,In_1459);
or U1892 (N_1892,In_1372,In_1105);
or U1893 (N_1893,In_362,In_1196);
or U1894 (N_1894,In_486,In_866);
nand U1895 (N_1895,In_33,In_458);
nand U1896 (N_1896,In_1370,In_270);
nand U1897 (N_1897,In_1117,In_1161);
nand U1898 (N_1898,In_1278,In_223);
and U1899 (N_1899,In_666,In_1148);
nand U1900 (N_1900,In_475,In_1011);
and U1901 (N_1901,In_18,In_1284);
or U1902 (N_1902,In_953,In_229);
and U1903 (N_1903,In_912,In_1319);
nor U1904 (N_1904,In_488,In_700);
and U1905 (N_1905,In_394,In_916);
nand U1906 (N_1906,In_1402,In_413);
nor U1907 (N_1907,In_847,In_697);
or U1908 (N_1908,In_381,In_761);
or U1909 (N_1909,In_1327,In_222);
or U1910 (N_1910,In_956,In_1044);
xor U1911 (N_1911,In_336,In_846);
nor U1912 (N_1912,In_661,In_459);
or U1913 (N_1913,In_717,In_482);
xnor U1914 (N_1914,In_1028,In_554);
or U1915 (N_1915,In_426,In_729);
nand U1916 (N_1916,In_1013,In_88);
nor U1917 (N_1917,In_547,In_844);
and U1918 (N_1918,In_360,In_926);
nand U1919 (N_1919,In_949,In_26);
nor U1920 (N_1920,In_670,In_180);
and U1921 (N_1921,In_317,In_953);
nor U1922 (N_1922,In_916,In_395);
or U1923 (N_1923,In_1239,In_78);
nand U1924 (N_1924,In_610,In_559);
or U1925 (N_1925,In_45,In_602);
xor U1926 (N_1926,In_1048,In_191);
nor U1927 (N_1927,In_313,In_637);
and U1928 (N_1928,In_535,In_1120);
nand U1929 (N_1929,In_553,In_1330);
or U1930 (N_1930,In_23,In_483);
or U1931 (N_1931,In_903,In_1380);
nor U1932 (N_1932,In_417,In_75);
nor U1933 (N_1933,In_487,In_1327);
nand U1934 (N_1934,In_1316,In_460);
nor U1935 (N_1935,In_712,In_1472);
or U1936 (N_1936,In_881,In_110);
or U1937 (N_1937,In_1321,In_1215);
nand U1938 (N_1938,In_1168,In_916);
nor U1939 (N_1939,In_1444,In_515);
nor U1940 (N_1940,In_662,In_396);
nor U1941 (N_1941,In_1371,In_178);
or U1942 (N_1942,In_895,In_1177);
and U1943 (N_1943,In_1314,In_1412);
nor U1944 (N_1944,In_65,In_481);
or U1945 (N_1945,In_1496,In_1358);
nor U1946 (N_1946,In_576,In_308);
or U1947 (N_1947,In_150,In_546);
xnor U1948 (N_1948,In_148,In_922);
nor U1949 (N_1949,In_387,In_192);
nand U1950 (N_1950,In_1048,In_501);
nor U1951 (N_1951,In_1367,In_70);
nor U1952 (N_1952,In_1129,In_1391);
or U1953 (N_1953,In_175,In_311);
xor U1954 (N_1954,In_421,In_481);
or U1955 (N_1955,In_1146,In_1001);
nor U1956 (N_1956,In_891,In_1268);
nand U1957 (N_1957,In_555,In_716);
and U1958 (N_1958,In_1049,In_22);
xor U1959 (N_1959,In_1426,In_1061);
and U1960 (N_1960,In_1298,In_17);
and U1961 (N_1961,In_786,In_328);
or U1962 (N_1962,In_506,In_336);
and U1963 (N_1963,In_406,In_422);
or U1964 (N_1964,In_678,In_1463);
or U1965 (N_1965,In_728,In_664);
xor U1966 (N_1966,In_96,In_275);
nand U1967 (N_1967,In_568,In_326);
and U1968 (N_1968,In_411,In_721);
nor U1969 (N_1969,In_142,In_1224);
and U1970 (N_1970,In_1010,In_205);
and U1971 (N_1971,In_1096,In_171);
nand U1972 (N_1972,In_1377,In_1044);
nor U1973 (N_1973,In_231,In_737);
or U1974 (N_1974,In_692,In_989);
nand U1975 (N_1975,In_336,In_436);
and U1976 (N_1976,In_78,In_208);
or U1977 (N_1977,In_1469,In_844);
and U1978 (N_1978,In_28,In_269);
xor U1979 (N_1979,In_45,In_1369);
nand U1980 (N_1980,In_786,In_65);
nor U1981 (N_1981,In_61,In_149);
xnor U1982 (N_1982,In_1121,In_768);
or U1983 (N_1983,In_834,In_1254);
nor U1984 (N_1984,In_116,In_504);
and U1985 (N_1985,In_1267,In_633);
nand U1986 (N_1986,In_868,In_269);
or U1987 (N_1987,In_802,In_48);
and U1988 (N_1988,In_608,In_273);
nand U1989 (N_1989,In_403,In_477);
nand U1990 (N_1990,In_1326,In_248);
xor U1991 (N_1991,In_629,In_1401);
or U1992 (N_1992,In_1103,In_875);
or U1993 (N_1993,In_877,In_1195);
xnor U1994 (N_1994,In_192,In_410);
or U1995 (N_1995,In_516,In_1206);
nor U1996 (N_1996,In_1468,In_469);
nand U1997 (N_1997,In_1064,In_1076);
xor U1998 (N_1998,In_1231,In_454);
or U1999 (N_1999,In_723,In_719);
nor U2000 (N_2000,In_613,In_742);
nand U2001 (N_2001,In_654,In_202);
and U2002 (N_2002,In_205,In_531);
xor U2003 (N_2003,In_303,In_338);
nor U2004 (N_2004,In_350,In_249);
nand U2005 (N_2005,In_1064,In_1080);
and U2006 (N_2006,In_307,In_603);
xor U2007 (N_2007,In_1026,In_1390);
nand U2008 (N_2008,In_771,In_84);
xnor U2009 (N_2009,In_1353,In_354);
nor U2010 (N_2010,In_796,In_1044);
or U2011 (N_2011,In_785,In_587);
or U2012 (N_2012,In_203,In_1047);
or U2013 (N_2013,In_873,In_133);
xnor U2014 (N_2014,In_238,In_1309);
or U2015 (N_2015,In_899,In_1201);
nand U2016 (N_2016,In_391,In_1348);
or U2017 (N_2017,In_567,In_1234);
and U2018 (N_2018,In_758,In_877);
nor U2019 (N_2019,In_1293,In_139);
and U2020 (N_2020,In_64,In_44);
nor U2021 (N_2021,In_634,In_655);
and U2022 (N_2022,In_633,In_692);
nor U2023 (N_2023,In_506,In_1417);
and U2024 (N_2024,In_248,In_132);
or U2025 (N_2025,In_385,In_267);
nand U2026 (N_2026,In_87,In_1104);
xor U2027 (N_2027,In_1027,In_1356);
xnor U2028 (N_2028,In_338,In_748);
nand U2029 (N_2029,In_27,In_1111);
and U2030 (N_2030,In_896,In_696);
or U2031 (N_2031,In_784,In_1205);
nand U2032 (N_2032,In_674,In_1223);
nor U2033 (N_2033,In_30,In_578);
or U2034 (N_2034,In_846,In_381);
and U2035 (N_2035,In_1143,In_851);
or U2036 (N_2036,In_149,In_931);
and U2037 (N_2037,In_794,In_651);
and U2038 (N_2038,In_1166,In_540);
nor U2039 (N_2039,In_1049,In_349);
or U2040 (N_2040,In_940,In_1165);
xnor U2041 (N_2041,In_729,In_645);
or U2042 (N_2042,In_1459,In_175);
nand U2043 (N_2043,In_1417,In_13);
nor U2044 (N_2044,In_907,In_74);
nand U2045 (N_2045,In_1254,In_543);
nor U2046 (N_2046,In_81,In_1107);
or U2047 (N_2047,In_685,In_1070);
nor U2048 (N_2048,In_418,In_1257);
nand U2049 (N_2049,In_646,In_1031);
nor U2050 (N_2050,In_424,In_830);
nor U2051 (N_2051,In_785,In_319);
nand U2052 (N_2052,In_697,In_1241);
and U2053 (N_2053,In_1205,In_238);
nor U2054 (N_2054,In_291,In_1187);
nor U2055 (N_2055,In_1091,In_1347);
or U2056 (N_2056,In_860,In_803);
nand U2057 (N_2057,In_287,In_299);
nor U2058 (N_2058,In_423,In_1255);
nor U2059 (N_2059,In_930,In_166);
nand U2060 (N_2060,In_303,In_916);
nand U2061 (N_2061,In_251,In_832);
nor U2062 (N_2062,In_1027,In_162);
nor U2063 (N_2063,In_1043,In_1243);
nor U2064 (N_2064,In_698,In_394);
or U2065 (N_2065,In_164,In_87);
xnor U2066 (N_2066,In_189,In_75);
and U2067 (N_2067,In_1041,In_845);
and U2068 (N_2068,In_1099,In_896);
or U2069 (N_2069,In_982,In_610);
nand U2070 (N_2070,In_79,In_444);
and U2071 (N_2071,In_784,In_1378);
or U2072 (N_2072,In_316,In_254);
nor U2073 (N_2073,In_447,In_1069);
nor U2074 (N_2074,In_179,In_222);
or U2075 (N_2075,In_774,In_854);
nand U2076 (N_2076,In_1321,In_1247);
and U2077 (N_2077,In_322,In_975);
or U2078 (N_2078,In_1448,In_41);
xnor U2079 (N_2079,In_107,In_298);
nand U2080 (N_2080,In_546,In_1225);
or U2081 (N_2081,In_534,In_999);
xor U2082 (N_2082,In_1426,In_1127);
nor U2083 (N_2083,In_690,In_1168);
xnor U2084 (N_2084,In_958,In_112);
or U2085 (N_2085,In_695,In_1215);
nand U2086 (N_2086,In_1062,In_625);
nor U2087 (N_2087,In_1007,In_187);
or U2088 (N_2088,In_826,In_308);
nor U2089 (N_2089,In_660,In_1244);
and U2090 (N_2090,In_448,In_235);
or U2091 (N_2091,In_762,In_928);
xnor U2092 (N_2092,In_1375,In_435);
xnor U2093 (N_2093,In_176,In_842);
nor U2094 (N_2094,In_498,In_1115);
nor U2095 (N_2095,In_1023,In_388);
or U2096 (N_2096,In_680,In_1477);
nand U2097 (N_2097,In_205,In_337);
xnor U2098 (N_2098,In_1013,In_842);
and U2099 (N_2099,In_1159,In_12);
or U2100 (N_2100,In_1492,In_644);
or U2101 (N_2101,In_218,In_1470);
or U2102 (N_2102,In_1277,In_1107);
nand U2103 (N_2103,In_1390,In_162);
nand U2104 (N_2104,In_769,In_789);
or U2105 (N_2105,In_545,In_1207);
nand U2106 (N_2106,In_726,In_667);
and U2107 (N_2107,In_758,In_1322);
nand U2108 (N_2108,In_116,In_346);
or U2109 (N_2109,In_950,In_358);
nand U2110 (N_2110,In_1007,In_1267);
and U2111 (N_2111,In_1066,In_271);
nand U2112 (N_2112,In_488,In_810);
nor U2113 (N_2113,In_440,In_142);
and U2114 (N_2114,In_95,In_319);
and U2115 (N_2115,In_613,In_1379);
or U2116 (N_2116,In_931,In_338);
and U2117 (N_2117,In_615,In_33);
nand U2118 (N_2118,In_36,In_117);
and U2119 (N_2119,In_889,In_1112);
nor U2120 (N_2120,In_580,In_253);
nor U2121 (N_2121,In_1288,In_857);
or U2122 (N_2122,In_114,In_1050);
nor U2123 (N_2123,In_1342,In_37);
and U2124 (N_2124,In_107,In_721);
or U2125 (N_2125,In_448,In_1331);
xor U2126 (N_2126,In_782,In_199);
nor U2127 (N_2127,In_803,In_23);
nor U2128 (N_2128,In_603,In_362);
and U2129 (N_2129,In_46,In_1071);
xnor U2130 (N_2130,In_960,In_1217);
and U2131 (N_2131,In_924,In_306);
or U2132 (N_2132,In_1218,In_636);
and U2133 (N_2133,In_19,In_153);
nor U2134 (N_2134,In_400,In_1217);
and U2135 (N_2135,In_13,In_204);
and U2136 (N_2136,In_1022,In_69);
nor U2137 (N_2137,In_224,In_1429);
and U2138 (N_2138,In_1147,In_1349);
xnor U2139 (N_2139,In_897,In_369);
nand U2140 (N_2140,In_1123,In_973);
nor U2141 (N_2141,In_1424,In_1085);
and U2142 (N_2142,In_386,In_259);
or U2143 (N_2143,In_1112,In_491);
nand U2144 (N_2144,In_1016,In_1129);
nor U2145 (N_2145,In_506,In_667);
or U2146 (N_2146,In_968,In_558);
nand U2147 (N_2147,In_736,In_1181);
and U2148 (N_2148,In_1226,In_370);
nor U2149 (N_2149,In_1466,In_973);
and U2150 (N_2150,In_982,In_209);
nand U2151 (N_2151,In_678,In_1213);
and U2152 (N_2152,In_247,In_294);
nor U2153 (N_2153,In_1109,In_630);
and U2154 (N_2154,In_1490,In_170);
nor U2155 (N_2155,In_501,In_1491);
or U2156 (N_2156,In_534,In_798);
nor U2157 (N_2157,In_1033,In_1471);
nor U2158 (N_2158,In_1228,In_425);
nand U2159 (N_2159,In_1475,In_145);
or U2160 (N_2160,In_753,In_904);
and U2161 (N_2161,In_267,In_228);
or U2162 (N_2162,In_1075,In_987);
nor U2163 (N_2163,In_1197,In_1336);
xor U2164 (N_2164,In_334,In_835);
nor U2165 (N_2165,In_723,In_751);
or U2166 (N_2166,In_523,In_736);
or U2167 (N_2167,In_716,In_683);
nand U2168 (N_2168,In_554,In_1477);
or U2169 (N_2169,In_516,In_798);
or U2170 (N_2170,In_523,In_726);
xnor U2171 (N_2171,In_1466,In_790);
or U2172 (N_2172,In_254,In_1344);
nor U2173 (N_2173,In_537,In_808);
and U2174 (N_2174,In_1016,In_349);
and U2175 (N_2175,In_1225,In_468);
nand U2176 (N_2176,In_1455,In_1155);
nor U2177 (N_2177,In_899,In_550);
nand U2178 (N_2178,In_1291,In_142);
nor U2179 (N_2179,In_722,In_714);
or U2180 (N_2180,In_851,In_313);
and U2181 (N_2181,In_1437,In_89);
or U2182 (N_2182,In_348,In_1021);
and U2183 (N_2183,In_392,In_631);
and U2184 (N_2184,In_1206,In_611);
nor U2185 (N_2185,In_293,In_320);
or U2186 (N_2186,In_309,In_1454);
nand U2187 (N_2187,In_836,In_1479);
nor U2188 (N_2188,In_132,In_920);
nand U2189 (N_2189,In_810,In_841);
nor U2190 (N_2190,In_4,In_693);
nor U2191 (N_2191,In_1007,In_446);
xnor U2192 (N_2192,In_870,In_166);
xor U2193 (N_2193,In_610,In_145);
nand U2194 (N_2194,In_1172,In_850);
nand U2195 (N_2195,In_435,In_1026);
nand U2196 (N_2196,In_1031,In_384);
xor U2197 (N_2197,In_8,In_300);
nor U2198 (N_2198,In_495,In_893);
and U2199 (N_2199,In_1470,In_705);
xor U2200 (N_2200,In_136,In_639);
nor U2201 (N_2201,In_337,In_1003);
nor U2202 (N_2202,In_97,In_320);
xnor U2203 (N_2203,In_50,In_1380);
xor U2204 (N_2204,In_1442,In_1065);
or U2205 (N_2205,In_1348,In_842);
or U2206 (N_2206,In_1051,In_327);
or U2207 (N_2207,In_111,In_1291);
nand U2208 (N_2208,In_1227,In_649);
or U2209 (N_2209,In_324,In_1048);
or U2210 (N_2210,In_812,In_29);
or U2211 (N_2211,In_1224,In_1044);
nand U2212 (N_2212,In_644,In_725);
nor U2213 (N_2213,In_688,In_72);
or U2214 (N_2214,In_885,In_975);
and U2215 (N_2215,In_1177,In_768);
nand U2216 (N_2216,In_1396,In_14);
nand U2217 (N_2217,In_11,In_882);
nor U2218 (N_2218,In_550,In_1344);
nor U2219 (N_2219,In_820,In_587);
nand U2220 (N_2220,In_92,In_833);
nor U2221 (N_2221,In_486,In_307);
nor U2222 (N_2222,In_1056,In_1345);
xor U2223 (N_2223,In_273,In_261);
nor U2224 (N_2224,In_191,In_572);
xnor U2225 (N_2225,In_848,In_1159);
and U2226 (N_2226,In_1213,In_463);
and U2227 (N_2227,In_460,In_91);
nor U2228 (N_2228,In_888,In_1240);
or U2229 (N_2229,In_1465,In_1263);
or U2230 (N_2230,In_1298,In_351);
nor U2231 (N_2231,In_464,In_1320);
or U2232 (N_2232,In_801,In_50);
nor U2233 (N_2233,In_860,In_1004);
nor U2234 (N_2234,In_114,In_621);
and U2235 (N_2235,In_1383,In_206);
and U2236 (N_2236,In_119,In_583);
nor U2237 (N_2237,In_1101,In_933);
or U2238 (N_2238,In_490,In_486);
xnor U2239 (N_2239,In_323,In_142);
nand U2240 (N_2240,In_92,In_581);
or U2241 (N_2241,In_675,In_211);
or U2242 (N_2242,In_1089,In_569);
nor U2243 (N_2243,In_1114,In_165);
and U2244 (N_2244,In_1499,In_265);
nand U2245 (N_2245,In_1215,In_972);
nor U2246 (N_2246,In_1062,In_1303);
or U2247 (N_2247,In_900,In_1116);
nand U2248 (N_2248,In_1411,In_1016);
or U2249 (N_2249,In_237,In_221);
nand U2250 (N_2250,In_835,In_917);
and U2251 (N_2251,In_25,In_374);
xor U2252 (N_2252,In_1215,In_338);
nor U2253 (N_2253,In_399,In_1063);
xor U2254 (N_2254,In_1193,In_643);
nand U2255 (N_2255,In_1276,In_1079);
nor U2256 (N_2256,In_1114,In_1180);
and U2257 (N_2257,In_1485,In_769);
or U2258 (N_2258,In_472,In_920);
nand U2259 (N_2259,In_779,In_62);
nand U2260 (N_2260,In_920,In_1313);
and U2261 (N_2261,In_641,In_294);
nand U2262 (N_2262,In_597,In_1293);
nand U2263 (N_2263,In_1131,In_795);
nor U2264 (N_2264,In_814,In_417);
or U2265 (N_2265,In_1266,In_922);
nor U2266 (N_2266,In_4,In_1336);
nand U2267 (N_2267,In_1261,In_128);
and U2268 (N_2268,In_1423,In_629);
xor U2269 (N_2269,In_295,In_859);
nor U2270 (N_2270,In_660,In_694);
nor U2271 (N_2271,In_720,In_202);
nand U2272 (N_2272,In_126,In_517);
and U2273 (N_2273,In_1491,In_840);
or U2274 (N_2274,In_1445,In_603);
and U2275 (N_2275,In_271,In_1442);
and U2276 (N_2276,In_1320,In_1304);
and U2277 (N_2277,In_810,In_648);
or U2278 (N_2278,In_820,In_1206);
nand U2279 (N_2279,In_310,In_828);
and U2280 (N_2280,In_1245,In_1299);
nor U2281 (N_2281,In_250,In_1129);
and U2282 (N_2282,In_1406,In_1384);
nor U2283 (N_2283,In_1033,In_309);
nor U2284 (N_2284,In_575,In_1021);
or U2285 (N_2285,In_574,In_576);
and U2286 (N_2286,In_672,In_1428);
or U2287 (N_2287,In_1464,In_858);
and U2288 (N_2288,In_893,In_275);
xnor U2289 (N_2289,In_405,In_878);
and U2290 (N_2290,In_1056,In_434);
and U2291 (N_2291,In_84,In_732);
or U2292 (N_2292,In_1372,In_1065);
xor U2293 (N_2293,In_1296,In_665);
nand U2294 (N_2294,In_1460,In_992);
and U2295 (N_2295,In_1073,In_1216);
nor U2296 (N_2296,In_1298,In_1213);
or U2297 (N_2297,In_49,In_1032);
and U2298 (N_2298,In_554,In_1479);
nand U2299 (N_2299,In_244,In_1395);
nand U2300 (N_2300,In_1470,In_442);
and U2301 (N_2301,In_227,In_709);
or U2302 (N_2302,In_1064,In_109);
nor U2303 (N_2303,In_1443,In_968);
nand U2304 (N_2304,In_449,In_1370);
and U2305 (N_2305,In_1092,In_959);
and U2306 (N_2306,In_1204,In_211);
or U2307 (N_2307,In_1005,In_178);
nor U2308 (N_2308,In_1304,In_1204);
nor U2309 (N_2309,In_327,In_565);
nor U2310 (N_2310,In_1136,In_838);
nor U2311 (N_2311,In_120,In_1453);
nor U2312 (N_2312,In_1280,In_1471);
and U2313 (N_2313,In_1117,In_1341);
xor U2314 (N_2314,In_738,In_861);
nand U2315 (N_2315,In_798,In_711);
nand U2316 (N_2316,In_711,In_572);
and U2317 (N_2317,In_203,In_147);
nand U2318 (N_2318,In_464,In_685);
or U2319 (N_2319,In_358,In_1122);
or U2320 (N_2320,In_663,In_200);
nor U2321 (N_2321,In_685,In_1173);
nand U2322 (N_2322,In_561,In_1176);
nand U2323 (N_2323,In_843,In_177);
nor U2324 (N_2324,In_557,In_221);
nor U2325 (N_2325,In_459,In_1066);
and U2326 (N_2326,In_8,In_1308);
nand U2327 (N_2327,In_834,In_588);
nand U2328 (N_2328,In_105,In_689);
nor U2329 (N_2329,In_148,In_327);
and U2330 (N_2330,In_405,In_994);
nand U2331 (N_2331,In_995,In_1247);
nor U2332 (N_2332,In_673,In_1497);
and U2333 (N_2333,In_355,In_484);
nand U2334 (N_2334,In_150,In_292);
or U2335 (N_2335,In_529,In_30);
or U2336 (N_2336,In_299,In_1315);
or U2337 (N_2337,In_1411,In_958);
xor U2338 (N_2338,In_732,In_508);
or U2339 (N_2339,In_1098,In_696);
nor U2340 (N_2340,In_550,In_523);
or U2341 (N_2341,In_727,In_827);
nor U2342 (N_2342,In_1465,In_1224);
nor U2343 (N_2343,In_1215,In_70);
or U2344 (N_2344,In_403,In_1441);
or U2345 (N_2345,In_947,In_473);
nand U2346 (N_2346,In_279,In_775);
and U2347 (N_2347,In_1004,In_412);
and U2348 (N_2348,In_491,In_1316);
and U2349 (N_2349,In_1100,In_185);
xnor U2350 (N_2350,In_1496,In_1474);
or U2351 (N_2351,In_53,In_168);
xnor U2352 (N_2352,In_1237,In_625);
nand U2353 (N_2353,In_1140,In_1074);
nand U2354 (N_2354,In_1098,In_384);
or U2355 (N_2355,In_40,In_57);
or U2356 (N_2356,In_22,In_316);
nor U2357 (N_2357,In_1410,In_1455);
nor U2358 (N_2358,In_637,In_531);
and U2359 (N_2359,In_1364,In_758);
or U2360 (N_2360,In_371,In_958);
and U2361 (N_2361,In_551,In_718);
nor U2362 (N_2362,In_1340,In_598);
nor U2363 (N_2363,In_901,In_65);
or U2364 (N_2364,In_446,In_826);
nor U2365 (N_2365,In_797,In_1384);
nor U2366 (N_2366,In_1344,In_1121);
nor U2367 (N_2367,In_1331,In_1082);
or U2368 (N_2368,In_660,In_1220);
nor U2369 (N_2369,In_18,In_62);
or U2370 (N_2370,In_1150,In_1344);
nand U2371 (N_2371,In_509,In_1063);
nand U2372 (N_2372,In_1026,In_1415);
xor U2373 (N_2373,In_241,In_125);
or U2374 (N_2374,In_1290,In_466);
xor U2375 (N_2375,In_644,In_1002);
and U2376 (N_2376,In_266,In_953);
nand U2377 (N_2377,In_1181,In_1071);
or U2378 (N_2378,In_523,In_1279);
nand U2379 (N_2379,In_581,In_1041);
nor U2380 (N_2380,In_815,In_300);
nor U2381 (N_2381,In_632,In_1227);
or U2382 (N_2382,In_114,In_681);
nand U2383 (N_2383,In_966,In_113);
nand U2384 (N_2384,In_612,In_541);
and U2385 (N_2385,In_225,In_268);
nand U2386 (N_2386,In_657,In_1087);
nand U2387 (N_2387,In_1392,In_418);
xor U2388 (N_2388,In_214,In_419);
nor U2389 (N_2389,In_92,In_1415);
nand U2390 (N_2390,In_851,In_168);
nor U2391 (N_2391,In_889,In_850);
nor U2392 (N_2392,In_633,In_718);
or U2393 (N_2393,In_1444,In_530);
nor U2394 (N_2394,In_1250,In_63);
nand U2395 (N_2395,In_217,In_995);
or U2396 (N_2396,In_370,In_1189);
and U2397 (N_2397,In_1253,In_307);
nand U2398 (N_2398,In_590,In_207);
and U2399 (N_2399,In_427,In_1452);
xnor U2400 (N_2400,In_500,In_1360);
or U2401 (N_2401,In_696,In_263);
nor U2402 (N_2402,In_292,In_1455);
or U2403 (N_2403,In_128,In_101);
or U2404 (N_2404,In_745,In_628);
and U2405 (N_2405,In_41,In_171);
nor U2406 (N_2406,In_118,In_1006);
and U2407 (N_2407,In_531,In_1181);
and U2408 (N_2408,In_536,In_408);
or U2409 (N_2409,In_1174,In_806);
and U2410 (N_2410,In_812,In_942);
or U2411 (N_2411,In_168,In_1064);
nand U2412 (N_2412,In_627,In_1110);
or U2413 (N_2413,In_698,In_208);
and U2414 (N_2414,In_1401,In_568);
or U2415 (N_2415,In_901,In_853);
nand U2416 (N_2416,In_1239,In_670);
nor U2417 (N_2417,In_1227,In_597);
nor U2418 (N_2418,In_635,In_1109);
nand U2419 (N_2419,In_500,In_796);
or U2420 (N_2420,In_297,In_545);
nor U2421 (N_2421,In_1056,In_1253);
and U2422 (N_2422,In_625,In_1117);
nor U2423 (N_2423,In_321,In_1285);
and U2424 (N_2424,In_863,In_383);
nand U2425 (N_2425,In_1034,In_1067);
nand U2426 (N_2426,In_788,In_345);
and U2427 (N_2427,In_487,In_494);
or U2428 (N_2428,In_703,In_261);
and U2429 (N_2429,In_456,In_1300);
nand U2430 (N_2430,In_678,In_1079);
and U2431 (N_2431,In_1256,In_667);
nand U2432 (N_2432,In_1037,In_779);
and U2433 (N_2433,In_14,In_445);
nor U2434 (N_2434,In_929,In_968);
nand U2435 (N_2435,In_235,In_330);
or U2436 (N_2436,In_517,In_434);
and U2437 (N_2437,In_1446,In_872);
and U2438 (N_2438,In_1444,In_68);
nor U2439 (N_2439,In_1252,In_222);
or U2440 (N_2440,In_857,In_513);
or U2441 (N_2441,In_1047,In_735);
nor U2442 (N_2442,In_1249,In_1364);
nor U2443 (N_2443,In_505,In_1133);
and U2444 (N_2444,In_1297,In_293);
and U2445 (N_2445,In_1469,In_803);
and U2446 (N_2446,In_288,In_136);
nor U2447 (N_2447,In_1010,In_889);
and U2448 (N_2448,In_991,In_923);
or U2449 (N_2449,In_1474,In_1181);
and U2450 (N_2450,In_1077,In_1280);
xor U2451 (N_2451,In_433,In_513);
nor U2452 (N_2452,In_1363,In_1287);
nor U2453 (N_2453,In_723,In_648);
nor U2454 (N_2454,In_1130,In_576);
nand U2455 (N_2455,In_345,In_60);
nand U2456 (N_2456,In_901,In_210);
or U2457 (N_2457,In_1075,In_290);
or U2458 (N_2458,In_933,In_768);
or U2459 (N_2459,In_866,In_365);
and U2460 (N_2460,In_1136,In_450);
nor U2461 (N_2461,In_583,In_1211);
nor U2462 (N_2462,In_791,In_632);
nor U2463 (N_2463,In_830,In_746);
nand U2464 (N_2464,In_509,In_201);
nor U2465 (N_2465,In_436,In_1204);
or U2466 (N_2466,In_127,In_1438);
or U2467 (N_2467,In_1481,In_52);
xor U2468 (N_2468,In_1005,In_1160);
or U2469 (N_2469,In_878,In_981);
and U2470 (N_2470,In_1183,In_1193);
or U2471 (N_2471,In_222,In_1296);
or U2472 (N_2472,In_375,In_523);
nor U2473 (N_2473,In_505,In_1386);
or U2474 (N_2474,In_1324,In_309);
xnor U2475 (N_2475,In_1433,In_706);
and U2476 (N_2476,In_214,In_112);
or U2477 (N_2477,In_698,In_1218);
and U2478 (N_2478,In_1211,In_1134);
and U2479 (N_2479,In_576,In_1438);
nand U2480 (N_2480,In_491,In_52);
nor U2481 (N_2481,In_1096,In_944);
xor U2482 (N_2482,In_683,In_663);
or U2483 (N_2483,In_1468,In_5);
nand U2484 (N_2484,In_749,In_1255);
nand U2485 (N_2485,In_1151,In_665);
nor U2486 (N_2486,In_658,In_39);
nand U2487 (N_2487,In_1460,In_191);
nor U2488 (N_2488,In_1374,In_237);
nand U2489 (N_2489,In_163,In_169);
and U2490 (N_2490,In_736,In_1025);
or U2491 (N_2491,In_1217,In_1197);
nor U2492 (N_2492,In_876,In_1443);
nor U2493 (N_2493,In_1112,In_1122);
nand U2494 (N_2494,In_1443,In_210);
or U2495 (N_2495,In_8,In_1453);
and U2496 (N_2496,In_585,In_863);
nand U2497 (N_2497,In_238,In_50);
nor U2498 (N_2498,In_1465,In_694);
xor U2499 (N_2499,In_1266,In_860);
or U2500 (N_2500,In_629,In_734);
nor U2501 (N_2501,In_1043,In_199);
xor U2502 (N_2502,In_670,In_1097);
and U2503 (N_2503,In_417,In_855);
or U2504 (N_2504,In_849,In_898);
nor U2505 (N_2505,In_1410,In_73);
or U2506 (N_2506,In_866,In_76);
or U2507 (N_2507,In_923,In_206);
xnor U2508 (N_2508,In_3,In_491);
xor U2509 (N_2509,In_103,In_228);
or U2510 (N_2510,In_683,In_1222);
and U2511 (N_2511,In_811,In_1073);
nor U2512 (N_2512,In_659,In_1440);
xor U2513 (N_2513,In_522,In_1058);
nand U2514 (N_2514,In_637,In_3);
nor U2515 (N_2515,In_1276,In_26);
or U2516 (N_2516,In_717,In_722);
and U2517 (N_2517,In_309,In_1101);
or U2518 (N_2518,In_1363,In_509);
or U2519 (N_2519,In_1096,In_53);
nor U2520 (N_2520,In_1166,In_389);
xor U2521 (N_2521,In_1357,In_838);
or U2522 (N_2522,In_879,In_1463);
nand U2523 (N_2523,In_477,In_1189);
or U2524 (N_2524,In_570,In_1396);
nand U2525 (N_2525,In_55,In_1198);
or U2526 (N_2526,In_602,In_407);
nand U2527 (N_2527,In_1153,In_1150);
nand U2528 (N_2528,In_1335,In_1473);
nor U2529 (N_2529,In_654,In_684);
or U2530 (N_2530,In_449,In_124);
nor U2531 (N_2531,In_1304,In_443);
nand U2532 (N_2532,In_1376,In_212);
nand U2533 (N_2533,In_935,In_523);
nand U2534 (N_2534,In_79,In_8);
and U2535 (N_2535,In_992,In_697);
or U2536 (N_2536,In_476,In_812);
nand U2537 (N_2537,In_1479,In_172);
and U2538 (N_2538,In_1101,In_398);
or U2539 (N_2539,In_1099,In_606);
xnor U2540 (N_2540,In_324,In_1046);
or U2541 (N_2541,In_1461,In_1348);
and U2542 (N_2542,In_672,In_637);
xnor U2543 (N_2543,In_1089,In_166);
and U2544 (N_2544,In_198,In_962);
or U2545 (N_2545,In_1486,In_658);
or U2546 (N_2546,In_732,In_28);
nand U2547 (N_2547,In_488,In_1067);
xor U2548 (N_2548,In_1141,In_1457);
nor U2549 (N_2549,In_622,In_432);
and U2550 (N_2550,In_738,In_919);
or U2551 (N_2551,In_833,In_1241);
or U2552 (N_2552,In_923,In_757);
xor U2553 (N_2553,In_934,In_1173);
and U2554 (N_2554,In_860,In_460);
or U2555 (N_2555,In_1152,In_1379);
nand U2556 (N_2556,In_632,In_789);
or U2557 (N_2557,In_388,In_59);
or U2558 (N_2558,In_595,In_88);
nand U2559 (N_2559,In_126,In_1312);
and U2560 (N_2560,In_1100,In_1437);
xor U2561 (N_2561,In_362,In_1195);
nor U2562 (N_2562,In_738,In_276);
nand U2563 (N_2563,In_209,In_1353);
and U2564 (N_2564,In_49,In_1018);
nor U2565 (N_2565,In_819,In_570);
nand U2566 (N_2566,In_20,In_4);
nand U2567 (N_2567,In_796,In_301);
nor U2568 (N_2568,In_1405,In_1206);
or U2569 (N_2569,In_539,In_63);
or U2570 (N_2570,In_269,In_763);
or U2571 (N_2571,In_535,In_1301);
nor U2572 (N_2572,In_1095,In_423);
nand U2573 (N_2573,In_1313,In_817);
nor U2574 (N_2574,In_1319,In_292);
or U2575 (N_2575,In_716,In_979);
or U2576 (N_2576,In_765,In_1132);
and U2577 (N_2577,In_1010,In_1258);
nor U2578 (N_2578,In_1448,In_126);
nor U2579 (N_2579,In_325,In_440);
xnor U2580 (N_2580,In_477,In_1083);
nor U2581 (N_2581,In_676,In_899);
nand U2582 (N_2582,In_217,In_462);
and U2583 (N_2583,In_926,In_349);
nand U2584 (N_2584,In_546,In_833);
nor U2585 (N_2585,In_420,In_430);
or U2586 (N_2586,In_596,In_269);
nor U2587 (N_2587,In_1194,In_400);
and U2588 (N_2588,In_357,In_1191);
and U2589 (N_2589,In_537,In_367);
xor U2590 (N_2590,In_1297,In_350);
nor U2591 (N_2591,In_1383,In_445);
and U2592 (N_2592,In_670,In_1449);
or U2593 (N_2593,In_1003,In_115);
nor U2594 (N_2594,In_691,In_1334);
and U2595 (N_2595,In_1009,In_1490);
nor U2596 (N_2596,In_831,In_1424);
and U2597 (N_2597,In_714,In_1350);
and U2598 (N_2598,In_374,In_1277);
or U2599 (N_2599,In_1309,In_242);
and U2600 (N_2600,In_1016,In_489);
xnor U2601 (N_2601,In_52,In_60);
or U2602 (N_2602,In_706,In_1047);
or U2603 (N_2603,In_727,In_1105);
nor U2604 (N_2604,In_364,In_242);
and U2605 (N_2605,In_1118,In_407);
or U2606 (N_2606,In_984,In_1390);
nor U2607 (N_2607,In_63,In_631);
nor U2608 (N_2608,In_815,In_802);
and U2609 (N_2609,In_693,In_240);
or U2610 (N_2610,In_1056,In_1310);
or U2611 (N_2611,In_1017,In_652);
or U2612 (N_2612,In_387,In_531);
nand U2613 (N_2613,In_337,In_929);
and U2614 (N_2614,In_233,In_744);
and U2615 (N_2615,In_517,In_930);
or U2616 (N_2616,In_676,In_705);
nand U2617 (N_2617,In_99,In_631);
and U2618 (N_2618,In_308,In_1472);
or U2619 (N_2619,In_499,In_279);
nand U2620 (N_2620,In_494,In_147);
and U2621 (N_2621,In_1059,In_1012);
nor U2622 (N_2622,In_4,In_615);
nor U2623 (N_2623,In_1195,In_869);
nor U2624 (N_2624,In_988,In_904);
and U2625 (N_2625,In_688,In_754);
xnor U2626 (N_2626,In_484,In_1350);
nand U2627 (N_2627,In_1085,In_810);
nor U2628 (N_2628,In_1089,In_1252);
nand U2629 (N_2629,In_443,In_342);
xnor U2630 (N_2630,In_31,In_201);
and U2631 (N_2631,In_305,In_672);
nand U2632 (N_2632,In_1259,In_1306);
or U2633 (N_2633,In_200,In_1368);
nand U2634 (N_2634,In_465,In_870);
nand U2635 (N_2635,In_622,In_1445);
and U2636 (N_2636,In_905,In_646);
nand U2637 (N_2637,In_774,In_741);
xor U2638 (N_2638,In_1308,In_1139);
and U2639 (N_2639,In_777,In_939);
nor U2640 (N_2640,In_991,In_1312);
nor U2641 (N_2641,In_1408,In_920);
and U2642 (N_2642,In_899,In_975);
xor U2643 (N_2643,In_671,In_581);
nand U2644 (N_2644,In_970,In_135);
or U2645 (N_2645,In_226,In_128);
nor U2646 (N_2646,In_477,In_904);
and U2647 (N_2647,In_1214,In_1107);
or U2648 (N_2648,In_387,In_1411);
or U2649 (N_2649,In_60,In_260);
xor U2650 (N_2650,In_1130,In_313);
and U2651 (N_2651,In_898,In_1031);
or U2652 (N_2652,In_1322,In_69);
xor U2653 (N_2653,In_379,In_737);
nor U2654 (N_2654,In_950,In_1397);
nand U2655 (N_2655,In_858,In_736);
or U2656 (N_2656,In_127,In_384);
nand U2657 (N_2657,In_209,In_837);
nor U2658 (N_2658,In_1061,In_490);
or U2659 (N_2659,In_24,In_972);
xor U2660 (N_2660,In_754,In_16);
and U2661 (N_2661,In_1266,In_1059);
nand U2662 (N_2662,In_895,In_704);
or U2663 (N_2663,In_1002,In_1429);
xnor U2664 (N_2664,In_1247,In_836);
nor U2665 (N_2665,In_1384,In_887);
nor U2666 (N_2666,In_139,In_1329);
nor U2667 (N_2667,In_387,In_1275);
nor U2668 (N_2668,In_779,In_186);
nor U2669 (N_2669,In_791,In_357);
and U2670 (N_2670,In_1196,In_1124);
nor U2671 (N_2671,In_778,In_15);
and U2672 (N_2672,In_1415,In_388);
or U2673 (N_2673,In_1387,In_267);
and U2674 (N_2674,In_620,In_975);
and U2675 (N_2675,In_832,In_512);
xor U2676 (N_2676,In_105,In_60);
or U2677 (N_2677,In_215,In_930);
xnor U2678 (N_2678,In_1354,In_848);
xnor U2679 (N_2679,In_974,In_15);
nand U2680 (N_2680,In_175,In_1355);
or U2681 (N_2681,In_1427,In_468);
or U2682 (N_2682,In_1019,In_78);
nand U2683 (N_2683,In_1438,In_40);
and U2684 (N_2684,In_1047,In_809);
xnor U2685 (N_2685,In_1273,In_344);
nor U2686 (N_2686,In_1388,In_875);
and U2687 (N_2687,In_982,In_33);
nor U2688 (N_2688,In_928,In_466);
xor U2689 (N_2689,In_23,In_308);
or U2690 (N_2690,In_1390,In_73);
or U2691 (N_2691,In_161,In_1155);
or U2692 (N_2692,In_1147,In_379);
nor U2693 (N_2693,In_1208,In_870);
or U2694 (N_2694,In_25,In_819);
or U2695 (N_2695,In_912,In_405);
xnor U2696 (N_2696,In_1424,In_1174);
xor U2697 (N_2697,In_944,In_687);
or U2698 (N_2698,In_1118,In_821);
and U2699 (N_2699,In_667,In_1315);
nor U2700 (N_2700,In_1186,In_520);
nor U2701 (N_2701,In_1392,In_144);
nor U2702 (N_2702,In_115,In_578);
or U2703 (N_2703,In_871,In_592);
or U2704 (N_2704,In_809,In_214);
nand U2705 (N_2705,In_1424,In_544);
nor U2706 (N_2706,In_1408,In_778);
or U2707 (N_2707,In_182,In_607);
and U2708 (N_2708,In_1042,In_693);
xor U2709 (N_2709,In_1025,In_23);
nand U2710 (N_2710,In_862,In_1425);
xor U2711 (N_2711,In_222,In_900);
and U2712 (N_2712,In_617,In_1056);
nor U2713 (N_2713,In_1342,In_1126);
nand U2714 (N_2714,In_840,In_208);
nor U2715 (N_2715,In_607,In_988);
and U2716 (N_2716,In_1099,In_372);
or U2717 (N_2717,In_691,In_275);
and U2718 (N_2718,In_160,In_36);
or U2719 (N_2719,In_741,In_1281);
nor U2720 (N_2720,In_170,In_1437);
nor U2721 (N_2721,In_708,In_838);
xor U2722 (N_2722,In_1372,In_587);
nand U2723 (N_2723,In_1223,In_498);
nor U2724 (N_2724,In_761,In_809);
nor U2725 (N_2725,In_1284,In_222);
nor U2726 (N_2726,In_188,In_901);
or U2727 (N_2727,In_1446,In_607);
or U2728 (N_2728,In_883,In_683);
and U2729 (N_2729,In_104,In_1064);
nand U2730 (N_2730,In_390,In_1034);
nand U2731 (N_2731,In_120,In_1156);
or U2732 (N_2732,In_84,In_127);
nand U2733 (N_2733,In_799,In_925);
nor U2734 (N_2734,In_536,In_1118);
or U2735 (N_2735,In_692,In_32);
nor U2736 (N_2736,In_587,In_980);
or U2737 (N_2737,In_940,In_404);
nor U2738 (N_2738,In_1425,In_924);
nor U2739 (N_2739,In_429,In_261);
and U2740 (N_2740,In_1360,In_346);
or U2741 (N_2741,In_615,In_1223);
or U2742 (N_2742,In_446,In_796);
nand U2743 (N_2743,In_139,In_320);
nand U2744 (N_2744,In_1303,In_774);
nor U2745 (N_2745,In_117,In_150);
nor U2746 (N_2746,In_808,In_497);
nor U2747 (N_2747,In_928,In_313);
nor U2748 (N_2748,In_32,In_248);
nor U2749 (N_2749,In_994,In_1396);
nand U2750 (N_2750,In_823,In_1138);
and U2751 (N_2751,In_125,In_114);
nor U2752 (N_2752,In_417,In_728);
and U2753 (N_2753,In_659,In_1373);
nand U2754 (N_2754,In_1425,In_1365);
nand U2755 (N_2755,In_1099,In_1041);
or U2756 (N_2756,In_272,In_859);
nor U2757 (N_2757,In_928,In_1195);
nor U2758 (N_2758,In_169,In_1258);
nand U2759 (N_2759,In_828,In_98);
nand U2760 (N_2760,In_1380,In_1002);
or U2761 (N_2761,In_942,In_675);
and U2762 (N_2762,In_573,In_1039);
nor U2763 (N_2763,In_74,In_1460);
and U2764 (N_2764,In_831,In_1279);
nand U2765 (N_2765,In_177,In_189);
or U2766 (N_2766,In_1046,In_876);
or U2767 (N_2767,In_1307,In_843);
and U2768 (N_2768,In_1341,In_59);
nand U2769 (N_2769,In_1229,In_991);
and U2770 (N_2770,In_383,In_790);
and U2771 (N_2771,In_978,In_1097);
and U2772 (N_2772,In_775,In_1128);
xnor U2773 (N_2773,In_665,In_457);
nor U2774 (N_2774,In_603,In_1029);
or U2775 (N_2775,In_447,In_536);
and U2776 (N_2776,In_106,In_100);
nand U2777 (N_2777,In_1284,In_1234);
nor U2778 (N_2778,In_23,In_951);
nor U2779 (N_2779,In_612,In_1430);
or U2780 (N_2780,In_101,In_728);
nor U2781 (N_2781,In_1214,In_1260);
nand U2782 (N_2782,In_549,In_1108);
and U2783 (N_2783,In_1193,In_571);
nand U2784 (N_2784,In_72,In_1163);
or U2785 (N_2785,In_523,In_629);
and U2786 (N_2786,In_593,In_799);
nor U2787 (N_2787,In_1359,In_536);
nor U2788 (N_2788,In_784,In_876);
nand U2789 (N_2789,In_925,In_433);
or U2790 (N_2790,In_470,In_441);
or U2791 (N_2791,In_300,In_1461);
or U2792 (N_2792,In_436,In_46);
or U2793 (N_2793,In_1451,In_299);
nor U2794 (N_2794,In_866,In_956);
and U2795 (N_2795,In_742,In_1311);
xor U2796 (N_2796,In_1331,In_1390);
or U2797 (N_2797,In_455,In_1009);
and U2798 (N_2798,In_893,In_1340);
nand U2799 (N_2799,In_117,In_333);
nand U2800 (N_2800,In_666,In_207);
nor U2801 (N_2801,In_1487,In_980);
nand U2802 (N_2802,In_509,In_367);
nand U2803 (N_2803,In_806,In_121);
nand U2804 (N_2804,In_1161,In_146);
xnor U2805 (N_2805,In_175,In_1083);
and U2806 (N_2806,In_1182,In_261);
and U2807 (N_2807,In_586,In_1357);
nor U2808 (N_2808,In_590,In_277);
or U2809 (N_2809,In_31,In_723);
xor U2810 (N_2810,In_99,In_1368);
nand U2811 (N_2811,In_942,In_736);
xor U2812 (N_2812,In_735,In_869);
nand U2813 (N_2813,In_128,In_529);
nand U2814 (N_2814,In_613,In_1422);
nor U2815 (N_2815,In_937,In_897);
nand U2816 (N_2816,In_60,In_176);
nor U2817 (N_2817,In_400,In_1129);
nor U2818 (N_2818,In_1316,In_1009);
nand U2819 (N_2819,In_866,In_401);
or U2820 (N_2820,In_1359,In_1171);
nand U2821 (N_2821,In_1486,In_1362);
nor U2822 (N_2822,In_1113,In_715);
nor U2823 (N_2823,In_1183,In_234);
nand U2824 (N_2824,In_181,In_783);
and U2825 (N_2825,In_630,In_426);
nand U2826 (N_2826,In_1256,In_652);
nand U2827 (N_2827,In_28,In_103);
nand U2828 (N_2828,In_634,In_857);
nand U2829 (N_2829,In_284,In_437);
nor U2830 (N_2830,In_565,In_20);
nor U2831 (N_2831,In_344,In_1143);
or U2832 (N_2832,In_30,In_1499);
nand U2833 (N_2833,In_604,In_929);
or U2834 (N_2834,In_1058,In_736);
nand U2835 (N_2835,In_552,In_204);
nand U2836 (N_2836,In_68,In_455);
nand U2837 (N_2837,In_1418,In_610);
and U2838 (N_2838,In_181,In_1216);
and U2839 (N_2839,In_625,In_437);
nor U2840 (N_2840,In_298,In_1099);
or U2841 (N_2841,In_113,In_1278);
or U2842 (N_2842,In_1475,In_1392);
xnor U2843 (N_2843,In_827,In_992);
nand U2844 (N_2844,In_630,In_604);
nand U2845 (N_2845,In_1158,In_1429);
nor U2846 (N_2846,In_1159,In_1366);
nand U2847 (N_2847,In_1039,In_62);
and U2848 (N_2848,In_1310,In_1248);
and U2849 (N_2849,In_253,In_1492);
nor U2850 (N_2850,In_920,In_923);
and U2851 (N_2851,In_496,In_450);
nand U2852 (N_2852,In_481,In_1046);
xnor U2853 (N_2853,In_203,In_815);
or U2854 (N_2854,In_1346,In_1393);
nand U2855 (N_2855,In_1089,In_107);
or U2856 (N_2856,In_842,In_779);
and U2857 (N_2857,In_174,In_919);
nand U2858 (N_2858,In_1268,In_272);
nor U2859 (N_2859,In_1034,In_226);
and U2860 (N_2860,In_336,In_463);
nor U2861 (N_2861,In_957,In_712);
nand U2862 (N_2862,In_1410,In_1351);
and U2863 (N_2863,In_106,In_1367);
xor U2864 (N_2864,In_672,In_750);
or U2865 (N_2865,In_820,In_724);
nor U2866 (N_2866,In_881,In_778);
or U2867 (N_2867,In_216,In_864);
and U2868 (N_2868,In_450,In_71);
and U2869 (N_2869,In_16,In_866);
xnor U2870 (N_2870,In_673,In_392);
nor U2871 (N_2871,In_1381,In_28);
xnor U2872 (N_2872,In_1141,In_966);
or U2873 (N_2873,In_564,In_389);
nand U2874 (N_2874,In_367,In_744);
or U2875 (N_2875,In_1172,In_218);
nand U2876 (N_2876,In_1475,In_1188);
nand U2877 (N_2877,In_1276,In_923);
nor U2878 (N_2878,In_611,In_81);
or U2879 (N_2879,In_1061,In_1237);
nand U2880 (N_2880,In_574,In_295);
nor U2881 (N_2881,In_1346,In_1259);
or U2882 (N_2882,In_1177,In_1480);
and U2883 (N_2883,In_1276,In_1460);
and U2884 (N_2884,In_1245,In_1348);
xor U2885 (N_2885,In_703,In_420);
xnor U2886 (N_2886,In_952,In_1330);
nand U2887 (N_2887,In_606,In_631);
nand U2888 (N_2888,In_505,In_763);
nor U2889 (N_2889,In_537,In_276);
nor U2890 (N_2890,In_924,In_787);
nor U2891 (N_2891,In_983,In_1495);
or U2892 (N_2892,In_253,In_298);
nand U2893 (N_2893,In_648,In_523);
nor U2894 (N_2894,In_198,In_1304);
xnor U2895 (N_2895,In_217,In_1086);
nor U2896 (N_2896,In_17,In_361);
or U2897 (N_2897,In_1129,In_1101);
or U2898 (N_2898,In_347,In_621);
nor U2899 (N_2899,In_7,In_1431);
nor U2900 (N_2900,In_1367,In_1226);
and U2901 (N_2901,In_530,In_338);
nand U2902 (N_2902,In_1247,In_812);
nor U2903 (N_2903,In_1199,In_698);
and U2904 (N_2904,In_1447,In_788);
and U2905 (N_2905,In_1065,In_188);
nor U2906 (N_2906,In_556,In_198);
nor U2907 (N_2907,In_633,In_1214);
or U2908 (N_2908,In_820,In_1047);
xor U2909 (N_2909,In_1441,In_787);
and U2910 (N_2910,In_5,In_1214);
and U2911 (N_2911,In_852,In_391);
nor U2912 (N_2912,In_239,In_382);
and U2913 (N_2913,In_1306,In_1468);
and U2914 (N_2914,In_695,In_466);
nor U2915 (N_2915,In_618,In_700);
nand U2916 (N_2916,In_498,In_195);
nor U2917 (N_2917,In_492,In_859);
nand U2918 (N_2918,In_1195,In_1496);
and U2919 (N_2919,In_1310,In_267);
or U2920 (N_2920,In_986,In_541);
or U2921 (N_2921,In_1237,In_326);
xnor U2922 (N_2922,In_742,In_727);
nand U2923 (N_2923,In_1187,In_946);
nand U2924 (N_2924,In_1122,In_1471);
xor U2925 (N_2925,In_156,In_679);
or U2926 (N_2926,In_1401,In_493);
nor U2927 (N_2927,In_1086,In_1311);
nor U2928 (N_2928,In_428,In_16);
nor U2929 (N_2929,In_1346,In_668);
and U2930 (N_2930,In_1358,In_83);
nand U2931 (N_2931,In_105,In_1116);
and U2932 (N_2932,In_1338,In_1001);
nor U2933 (N_2933,In_184,In_697);
xor U2934 (N_2934,In_1165,In_661);
and U2935 (N_2935,In_591,In_65);
or U2936 (N_2936,In_955,In_1357);
or U2937 (N_2937,In_635,In_604);
or U2938 (N_2938,In_145,In_941);
or U2939 (N_2939,In_849,In_769);
nand U2940 (N_2940,In_643,In_254);
or U2941 (N_2941,In_1124,In_1101);
nand U2942 (N_2942,In_5,In_110);
nand U2943 (N_2943,In_529,In_1148);
or U2944 (N_2944,In_1034,In_427);
nand U2945 (N_2945,In_1141,In_840);
or U2946 (N_2946,In_977,In_478);
nor U2947 (N_2947,In_1350,In_542);
and U2948 (N_2948,In_189,In_1149);
nand U2949 (N_2949,In_783,In_199);
nand U2950 (N_2950,In_102,In_1117);
xor U2951 (N_2951,In_252,In_86);
xor U2952 (N_2952,In_700,In_505);
or U2953 (N_2953,In_948,In_1086);
nor U2954 (N_2954,In_267,In_1093);
or U2955 (N_2955,In_493,In_1075);
nand U2956 (N_2956,In_301,In_1038);
nand U2957 (N_2957,In_737,In_1496);
nand U2958 (N_2958,In_883,In_1462);
nand U2959 (N_2959,In_901,In_1423);
nor U2960 (N_2960,In_1145,In_1401);
or U2961 (N_2961,In_1318,In_158);
nand U2962 (N_2962,In_543,In_526);
nor U2963 (N_2963,In_1343,In_751);
and U2964 (N_2964,In_146,In_817);
or U2965 (N_2965,In_1110,In_1036);
xnor U2966 (N_2966,In_1194,In_756);
or U2967 (N_2967,In_1013,In_1315);
nand U2968 (N_2968,In_553,In_1093);
nor U2969 (N_2969,In_1403,In_1052);
and U2970 (N_2970,In_749,In_613);
nand U2971 (N_2971,In_551,In_353);
and U2972 (N_2972,In_175,In_569);
nor U2973 (N_2973,In_1068,In_259);
nor U2974 (N_2974,In_1496,In_1480);
nand U2975 (N_2975,In_731,In_464);
and U2976 (N_2976,In_853,In_58);
and U2977 (N_2977,In_1493,In_181);
xnor U2978 (N_2978,In_319,In_114);
xor U2979 (N_2979,In_787,In_971);
and U2980 (N_2980,In_1207,In_1170);
xor U2981 (N_2981,In_1185,In_1201);
and U2982 (N_2982,In_1303,In_470);
nand U2983 (N_2983,In_809,In_1319);
and U2984 (N_2984,In_351,In_1016);
or U2985 (N_2985,In_1271,In_1453);
nor U2986 (N_2986,In_1279,In_1217);
nand U2987 (N_2987,In_1327,In_1329);
xor U2988 (N_2988,In_1240,In_1043);
nor U2989 (N_2989,In_324,In_1435);
nand U2990 (N_2990,In_375,In_702);
nand U2991 (N_2991,In_1488,In_770);
or U2992 (N_2992,In_187,In_1014);
or U2993 (N_2993,In_983,In_1484);
or U2994 (N_2994,In_1126,In_1127);
xnor U2995 (N_2995,In_233,In_918);
nand U2996 (N_2996,In_1107,In_1390);
and U2997 (N_2997,In_818,In_1207);
and U2998 (N_2998,In_1357,In_1217);
nor U2999 (N_2999,In_543,In_1008);
nor U3000 (N_3000,N_2537,N_2803);
nand U3001 (N_3001,N_2364,N_2098);
xnor U3002 (N_3002,N_362,N_1218);
nor U3003 (N_3003,N_1973,N_719);
nand U3004 (N_3004,N_1528,N_1696);
nor U3005 (N_3005,N_1548,N_2448);
or U3006 (N_3006,N_499,N_1034);
nand U3007 (N_3007,N_30,N_1748);
nor U3008 (N_3008,N_1722,N_2682);
and U3009 (N_3009,N_1462,N_1094);
or U3010 (N_3010,N_1603,N_2414);
nand U3011 (N_3011,N_2193,N_330);
nor U3012 (N_3012,N_883,N_574);
and U3013 (N_3013,N_960,N_1683);
xnor U3014 (N_3014,N_1820,N_346);
and U3015 (N_3015,N_132,N_934);
or U3016 (N_3016,N_1488,N_1285);
xnor U3017 (N_3017,N_494,N_2099);
or U3018 (N_3018,N_1172,N_1938);
nand U3019 (N_3019,N_995,N_2360);
and U3020 (N_3020,N_2436,N_2766);
nor U3021 (N_3021,N_2369,N_2569);
nor U3022 (N_3022,N_2928,N_2594);
or U3023 (N_3023,N_546,N_1658);
nand U3024 (N_3024,N_789,N_43);
xor U3025 (N_3025,N_1768,N_1644);
nor U3026 (N_3026,N_54,N_882);
nand U3027 (N_3027,N_416,N_2015);
and U3028 (N_3028,N_2916,N_561);
nor U3029 (N_3029,N_87,N_2684);
and U3030 (N_3030,N_1984,N_2900);
nand U3031 (N_3031,N_1915,N_1381);
and U3032 (N_3032,N_1982,N_1123);
xor U3033 (N_3033,N_1415,N_981);
nor U3034 (N_3034,N_1663,N_1229);
and U3035 (N_3035,N_2323,N_472);
or U3036 (N_3036,N_1519,N_2996);
nand U3037 (N_3037,N_2646,N_2069);
xor U3038 (N_3038,N_2267,N_484);
or U3039 (N_3039,N_535,N_1131);
nor U3040 (N_3040,N_1595,N_2999);
or U3041 (N_3041,N_1120,N_699);
nand U3042 (N_3042,N_2269,N_1135);
or U3043 (N_3043,N_1787,N_197);
and U3044 (N_3044,N_2093,N_1894);
nand U3045 (N_3045,N_1966,N_800);
nor U3046 (N_3046,N_1088,N_856);
xor U3047 (N_3047,N_2903,N_33);
nand U3048 (N_3048,N_493,N_1236);
nor U3049 (N_3049,N_614,N_1186);
and U3050 (N_3050,N_1056,N_1671);
nand U3051 (N_3051,N_101,N_2725);
nor U3052 (N_3052,N_1864,N_77);
and U3053 (N_3053,N_2678,N_2019);
and U3054 (N_3054,N_2089,N_319);
nand U3055 (N_3055,N_1339,N_837);
nor U3056 (N_3056,N_1275,N_1495);
nand U3057 (N_3057,N_2181,N_2653);
and U3058 (N_3058,N_2250,N_918);
nand U3059 (N_3059,N_2525,N_978);
nand U3060 (N_3060,N_2681,N_2306);
nand U3061 (N_3061,N_1446,N_154);
nor U3062 (N_3062,N_858,N_1622);
nand U3063 (N_3063,N_1659,N_1070);
or U3064 (N_3064,N_1,N_1393);
nand U3065 (N_3065,N_2590,N_2246);
or U3066 (N_3066,N_1932,N_2844);
and U3067 (N_3067,N_10,N_66);
nor U3068 (N_3068,N_1771,N_2856);
nor U3069 (N_3069,N_720,N_185);
xor U3070 (N_3070,N_2187,N_620);
or U3071 (N_3071,N_1277,N_1247);
nor U3072 (N_3072,N_1078,N_2483);
nand U3073 (N_3073,N_2162,N_756);
and U3074 (N_3074,N_2200,N_1109);
or U3075 (N_3075,N_223,N_1505);
xor U3076 (N_3076,N_2373,N_152);
xor U3077 (N_3077,N_2127,N_1125);
nand U3078 (N_3078,N_806,N_1767);
nand U3079 (N_3079,N_2042,N_255);
or U3080 (N_3080,N_1053,N_1835);
and U3081 (N_3081,N_2126,N_64);
nor U3082 (N_3082,N_2888,N_277);
nand U3083 (N_3083,N_2602,N_2346);
nor U3084 (N_3084,N_2396,N_1266);
nand U3085 (N_3085,N_1292,N_977);
nor U3086 (N_3086,N_2493,N_1886);
nor U3087 (N_3087,N_1399,N_1029);
and U3088 (N_3088,N_2988,N_1838);
nor U3089 (N_3089,N_2268,N_860);
or U3090 (N_3090,N_287,N_2011);
xor U3091 (N_3091,N_322,N_318);
nand U3092 (N_3092,N_1589,N_2733);
nor U3093 (N_3093,N_1591,N_2121);
or U3094 (N_3094,N_2545,N_137);
xnor U3095 (N_3095,N_529,N_704);
or U3096 (N_3096,N_969,N_1279);
nand U3097 (N_3097,N_1686,N_1005);
or U3098 (N_3098,N_183,N_964);
and U3099 (N_3099,N_486,N_1171);
nand U3100 (N_3100,N_1910,N_2224);
nand U3101 (N_3101,N_1583,N_2066);
and U3102 (N_3102,N_2980,N_1956);
nand U3103 (N_3103,N_2951,N_79);
xnor U3104 (N_3104,N_2878,N_376);
or U3105 (N_3105,N_1244,N_1240);
or U3106 (N_3106,N_2519,N_1269);
nor U3107 (N_3107,N_1342,N_2206);
and U3108 (N_3108,N_1365,N_2673);
and U3109 (N_3109,N_2391,N_2057);
nand U3110 (N_3110,N_1300,N_2022);
nand U3111 (N_3111,N_109,N_2504);
nor U3112 (N_3112,N_448,N_742);
or U3113 (N_3113,N_524,N_2741);
or U3114 (N_3114,N_2430,N_1032);
and U3115 (N_3115,N_1968,N_686);
and U3116 (N_3116,N_2570,N_2552);
nor U3117 (N_3117,N_1732,N_1922);
xnor U3118 (N_3118,N_2593,N_1202);
or U3119 (N_3119,N_2070,N_1931);
xor U3120 (N_3120,N_2686,N_804);
or U3121 (N_3121,N_2804,N_1112);
and U3122 (N_3122,N_1978,N_2397);
or U3123 (N_3123,N_611,N_1550);
xnor U3124 (N_3124,N_1570,N_1454);
or U3125 (N_3125,N_955,N_2122);
nand U3126 (N_3126,N_42,N_2288);
or U3127 (N_3127,N_2751,N_823);
and U3128 (N_3128,N_24,N_413);
or U3129 (N_3129,N_2103,N_1116);
xor U3130 (N_3130,N_1627,N_2600);
and U3131 (N_3131,N_1345,N_2447);
nor U3132 (N_3132,N_2025,N_452);
and U3133 (N_3133,N_2734,N_1332);
nand U3134 (N_3134,N_666,N_1535);
nor U3135 (N_3135,N_2439,N_1189);
nand U3136 (N_3136,N_1650,N_2182);
nand U3137 (N_3137,N_7,N_1261);
and U3138 (N_3138,N_631,N_1118);
or U3139 (N_3139,N_1753,N_1974);
and U3140 (N_3140,N_296,N_1106);
nand U3141 (N_3141,N_573,N_503);
and U3142 (N_3142,N_2562,N_1308);
nor U3143 (N_3143,N_145,N_1513);
nor U3144 (N_3144,N_2976,N_2925);
or U3145 (N_3145,N_623,N_2072);
nand U3146 (N_3146,N_2960,N_831);
xnor U3147 (N_3147,N_1062,N_2514);
and U3148 (N_3148,N_644,N_1940);
and U3149 (N_3149,N_2505,N_2754);
nor U3150 (N_3150,N_1882,N_2050);
and U3151 (N_3151,N_972,N_495);
or U3152 (N_3152,N_2843,N_830);
nand U3153 (N_3153,N_1044,N_779);
nand U3154 (N_3154,N_1039,N_2502);
nor U3155 (N_3155,N_95,N_568);
nand U3156 (N_3156,N_437,N_2654);
or U3157 (N_3157,N_2732,N_327);
nor U3158 (N_3158,N_117,N_1201);
or U3159 (N_3159,N_2131,N_2938);
or U3160 (N_3160,N_533,N_1992);
or U3161 (N_3161,N_526,N_570);
nand U3162 (N_3162,N_2293,N_2995);
nor U3163 (N_3163,N_1432,N_1874);
nand U3164 (N_3164,N_721,N_2290);
and U3165 (N_3165,N_712,N_2252);
and U3166 (N_3166,N_1544,N_500);
and U3167 (N_3167,N_1316,N_1442);
nand U3168 (N_3168,N_1810,N_1074);
or U3169 (N_3169,N_557,N_1414);
and U3170 (N_3170,N_1936,N_194);
xnor U3171 (N_3171,N_1440,N_1404);
nand U3172 (N_3172,N_1605,N_868);
xor U3173 (N_3173,N_1610,N_1108);
or U3174 (N_3174,N_656,N_1041);
or U3175 (N_3175,N_1167,N_1000);
and U3176 (N_3176,N_2120,N_82);
nand U3177 (N_3177,N_1181,N_348);
nor U3178 (N_3178,N_2344,N_1560);
or U3179 (N_3179,N_1649,N_1666);
xor U3180 (N_3180,N_1707,N_737);
xor U3181 (N_3181,N_740,N_1871);
nand U3182 (N_3182,N_2768,N_2541);
nor U3183 (N_3183,N_1066,N_2286);
or U3184 (N_3184,N_1177,N_2076);
nor U3185 (N_3185,N_2518,N_1290);
and U3186 (N_3186,N_57,N_177);
nand U3187 (N_3187,N_2532,N_2220);
xnor U3188 (N_3188,N_2873,N_1929);
xor U3189 (N_3189,N_2917,N_547);
nand U3190 (N_3190,N_106,N_1493);
or U3191 (N_3191,N_358,N_807);
and U3192 (N_3192,N_2125,N_605);
and U3193 (N_3193,N_371,N_1766);
and U3194 (N_3194,N_1776,N_1945);
nand U3195 (N_3195,N_1369,N_896);
nand U3196 (N_3196,N_2990,N_1312);
nor U3197 (N_3197,N_86,N_253);
or U3198 (N_3198,N_2535,N_2141);
and U3199 (N_3199,N_312,N_1380);
and U3200 (N_3200,N_1188,N_1789);
xnor U3201 (N_3201,N_399,N_2491);
xor U3202 (N_3202,N_239,N_67);
nor U3203 (N_3203,N_2728,N_2589);
nand U3204 (N_3204,N_554,N_1654);
nor U3205 (N_3205,N_1738,N_2598);
nand U3206 (N_3206,N_1010,N_2939);
and U3207 (N_3207,N_1356,N_2891);
or U3208 (N_3208,N_1750,N_141);
nand U3209 (N_3209,N_744,N_1711);
nand U3210 (N_3210,N_369,N_1001);
nand U3211 (N_3211,N_2607,N_626);
nand U3212 (N_3212,N_1567,N_150);
nand U3213 (N_3213,N_1107,N_116);
and U3214 (N_3214,N_462,N_938);
nor U3215 (N_3215,N_1427,N_1853);
xor U3216 (N_3216,N_1652,N_361);
nor U3217 (N_3217,N_2394,N_1788);
and U3218 (N_3218,N_460,N_2672);
and U3219 (N_3219,N_1095,N_26);
nor U3220 (N_3220,N_1258,N_1971);
and U3221 (N_3221,N_665,N_1815);
nand U3222 (N_3222,N_2329,N_295);
or U3223 (N_3223,N_1273,N_13);
and U3224 (N_3224,N_1504,N_1217);
and U3225 (N_3225,N_270,N_2029);
xor U3226 (N_3226,N_687,N_1139);
and U3227 (N_3227,N_2544,N_39);
or U3228 (N_3228,N_507,N_1555);
nor U3229 (N_3229,N_2304,N_1297);
xor U3230 (N_3230,N_2998,N_2561);
xor U3231 (N_3231,N_2802,N_181);
nand U3232 (N_3232,N_2566,N_2223);
nor U3233 (N_3233,N_1304,N_1720);
xnor U3234 (N_3234,N_506,N_192);
nor U3235 (N_3235,N_2437,N_373);
and U3236 (N_3236,N_2415,N_1411);
or U3237 (N_3237,N_316,N_2467);
or U3238 (N_3238,N_966,N_1621);
and U3239 (N_3239,N_638,N_1930);
xor U3240 (N_3240,N_2641,N_786);
xnor U3241 (N_3241,N_35,N_1645);
and U3242 (N_3242,N_388,N_1322);
nand U3243 (N_3243,N_846,N_12);
nor U3244 (N_3244,N_2282,N_1180);
nand U3245 (N_3245,N_1872,N_2339);
xnor U3246 (N_3246,N_228,N_286);
nor U3247 (N_3247,N_2595,N_1698);
and U3248 (N_3248,N_2817,N_2406);
or U3249 (N_3249,N_1841,N_27);
nand U3250 (N_3250,N_889,N_368);
nor U3251 (N_3251,N_2738,N_2934);
and U3252 (N_3252,N_1408,N_1885);
nand U3253 (N_3253,N_1140,N_625);
nor U3254 (N_3254,N_2210,N_2845);
and U3255 (N_3255,N_2533,N_2813);
nand U3256 (N_3256,N_232,N_2006);
and U3257 (N_3257,N_1298,N_1418);
or U3258 (N_3258,N_1975,N_1642);
nand U3259 (N_3259,N_2407,N_748);
nor U3260 (N_3260,N_1455,N_52);
and U3261 (N_3261,N_1026,N_2706);
and U3262 (N_3262,N_1330,N_2184);
xor U3263 (N_3263,N_0,N_465);
nor U3264 (N_3264,N_2096,N_124);
and U3265 (N_3265,N_2107,N_2978);
nand U3266 (N_3266,N_1684,N_191);
and U3267 (N_3267,N_1749,N_2579);
nand U3268 (N_3268,N_1863,N_336);
nand U3269 (N_3269,N_2331,N_2771);
nor U3270 (N_3270,N_887,N_715);
and U3271 (N_3271,N_2135,N_994);
and U3272 (N_3272,N_2826,N_2059);
nand U3273 (N_3273,N_76,N_1407);
or U3274 (N_3274,N_1335,N_1469);
nand U3275 (N_3275,N_2580,N_2972);
and U3276 (N_3276,N_2388,N_2667);
nor U3277 (N_3277,N_2823,N_479);
or U3278 (N_3278,N_1822,N_387);
and U3279 (N_3279,N_2547,N_759);
nand U3280 (N_3280,N_2991,N_927);
nor U3281 (N_3281,N_1508,N_2134);
and U3282 (N_3282,N_2597,N_1134);
and U3283 (N_3283,N_1199,N_1710);
or U3284 (N_3284,N_2425,N_2866);
or U3285 (N_3285,N_2529,N_2379);
nor U3286 (N_3286,N_1705,N_1367);
and U3287 (N_3287,N_653,N_2772);
nor U3288 (N_3288,N_751,N_2175);
nor U3289 (N_3289,N_2926,N_2719);
and U3290 (N_3290,N_634,N_1182);
or U3291 (N_3291,N_902,N_1348);
and U3292 (N_3292,N_32,N_2523);
xnor U3293 (N_3293,N_645,N_1828);
nor U3294 (N_3294,N_401,N_2168);
and U3295 (N_3295,N_212,N_1307);
or U3296 (N_3296,N_2305,N_37);
and U3297 (N_3297,N_947,N_2016);
or U3298 (N_3298,N_671,N_1487);
nor U3299 (N_3299,N_491,N_2639);
or U3300 (N_3300,N_637,N_1558);
xnor U3301 (N_3301,N_1250,N_1856);
nor U3302 (N_3302,N_1206,N_224);
xnor U3303 (N_3303,N_1092,N_2992);
nand U3304 (N_3304,N_2136,N_690);
xnor U3305 (N_3305,N_394,N_1374);
and U3306 (N_3306,N_2703,N_1607);
nor U3307 (N_3307,N_724,N_867);
or U3308 (N_3308,N_2695,N_222);
xnor U3309 (N_3309,N_1214,N_1800);
or U3310 (N_3310,N_1124,N_848);
and U3311 (N_3311,N_1260,N_2962);
and U3312 (N_3312,N_488,N_1081);
nor U3313 (N_3313,N_2730,N_1594);
nor U3314 (N_3314,N_2221,N_153);
xnor U3315 (N_3315,N_2188,N_600);
nor U3316 (N_3316,N_1765,N_1475);
or U3317 (N_3317,N_8,N_1902);
nor U3318 (N_3318,N_905,N_1173);
and U3319 (N_3319,N_1772,N_1803);
nor U3320 (N_3320,N_1278,N_958);
xnor U3321 (N_3321,N_1251,N_1055);
or U3322 (N_3322,N_113,N_207);
nand U3323 (N_3323,N_767,N_734);
nand U3324 (N_3324,N_703,N_2838);
and U3325 (N_3325,N_1063,N_937);
nand U3326 (N_3326,N_2337,N_236);
or U3327 (N_3327,N_1581,N_2281);
and U3328 (N_3328,N_1879,N_241);
or U3329 (N_3329,N_1373,N_2446);
and U3330 (N_3330,N_2117,N_1104);
xnor U3331 (N_3331,N_446,N_2499);
nor U3332 (N_3332,N_1067,N_1018);
nand U3333 (N_3333,N_2231,N_2465);
nor U3334 (N_3334,N_1518,N_195);
nand U3335 (N_3335,N_1352,N_2612);
nor U3336 (N_3336,N_1631,N_2746);
nand U3337 (N_3337,N_2133,N_107);
and U3338 (N_3338,N_741,N_1023);
or U3339 (N_3339,N_1629,N_1540);
or U3340 (N_3340,N_2749,N_2124);
and U3341 (N_3341,N_1386,N_2827);
xor U3342 (N_3342,N_2949,N_962);
xor U3343 (N_3343,N_2160,N_2553);
nand U3344 (N_3344,N_60,N_1573);
xnor U3345 (N_3345,N_1498,N_2756);
and U3346 (N_3346,N_2457,N_2509);
xor U3347 (N_3347,N_2086,N_916);
or U3348 (N_3348,N_451,N_63);
nor U3349 (N_3349,N_1951,N_2222);
or U3350 (N_3350,N_372,N_925);
or U3351 (N_3351,N_1576,N_2779);
nand U3352 (N_3352,N_636,N_2435);
or U3353 (N_3353,N_426,N_337);
nor U3354 (N_3354,N_843,N_254);
nand U3355 (N_3355,N_1525,N_2936);
and U3356 (N_3356,N_44,N_1080);
nor U3357 (N_3357,N_799,N_2979);
nor U3358 (N_3358,N_1578,N_1150);
and U3359 (N_3359,N_1861,N_1831);
nor U3360 (N_3360,N_2717,N_335);
or U3361 (N_3361,N_884,N_1472);
nor U3362 (N_3362,N_1618,N_2084);
and U3363 (N_3363,N_2104,N_1675);
xnor U3364 (N_3364,N_2575,N_445);
or U3365 (N_3365,N_338,N_68);
or U3366 (N_3366,N_2488,N_542);
and U3367 (N_3367,N_2020,N_293);
nand U3368 (N_3368,N_617,N_1769);
and U3369 (N_3369,N_819,N_615);
nor U3370 (N_3370,N_2877,N_257);
xnor U3371 (N_3371,N_1632,N_2894);
and U3372 (N_3372,N_467,N_1762);
and U3373 (N_3373,N_1877,N_2308);
nand U3374 (N_3374,N_853,N_2530);
or U3375 (N_3375,N_2883,N_1763);
nor U3376 (N_3376,N_2538,N_709);
and U3377 (N_3377,N_1281,N_1406);
and U3378 (N_3378,N_1702,N_377);
nand U3379 (N_3379,N_2138,N_289);
nor U3380 (N_3380,N_2325,N_1834);
or U3381 (N_3381,N_504,N_72);
nor U3382 (N_3382,N_2359,N_1382);
nand U3383 (N_3383,N_1985,N_200);
and U3384 (N_3384,N_171,N_360);
or U3385 (N_3385,N_2413,N_581);
nand U3386 (N_3386,N_359,N_1895);
nand U3387 (N_3387,N_1817,N_2558);
or U3388 (N_3388,N_1635,N_332);
nor U3389 (N_3389,N_2034,N_2164);
nand U3390 (N_3390,N_383,N_1204);
or U3391 (N_3391,N_1816,N_872);
nand U3392 (N_3392,N_201,N_2898);
nor U3393 (N_3393,N_263,N_461);
nand U3394 (N_3394,N_607,N_2235);
and U3395 (N_3395,N_1448,N_539);
nor U3396 (N_3396,N_2197,N_1859);
and U3397 (N_3397,N_757,N_833);
or U3398 (N_3398,N_2309,N_1999);
or U3399 (N_3399,N_2140,N_412);
and U3400 (N_3400,N_817,N_1830);
or U3401 (N_3401,N_1630,N_1137);
and U3402 (N_3402,N_1007,N_1624);
nand U3403 (N_3403,N_411,N_2062);
nand U3404 (N_3404,N_402,N_2820);
and U3405 (N_3405,N_1031,N_2791);
nand U3406 (N_3406,N_237,N_2777);
nand U3407 (N_3407,N_400,N_1203);
nor U3408 (N_3408,N_2808,N_2555);
nand U3409 (N_3409,N_2361,N_2053);
or U3410 (N_3410,N_2243,N_1572);
nor U3411 (N_3411,N_1741,N_1101);
or U3412 (N_3412,N_2317,N_180);
nand U3413 (N_3413,N_2985,N_1935);
and U3414 (N_3414,N_1794,N_1643);
or U3415 (N_3415,N_1954,N_2257);
xor U3416 (N_3416,N_1138,N_2387);
nand U3417 (N_3417,N_159,N_697);
nor U3418 (N_3418,N_1383,N_1176);
or U3419 (N_3419,N_1503,N_549);
or U3420 (N_3420,N_1646,N_822);
nand U3421 (N_3421,N_1328,N_99);
nand U3422 (N_3422,N_1371,N_2662);
nand U3423 (N_3423,N_1235,N_1678);
and U3424 (N_3424,N_523,N_2186);
and U3425 (N_3425,N_341,N_1227);
nor U3426 (N_3426,N_1990,N_588);
or U3427 (N_3427,N_84,N_249);
nand U3428 (N_3428,N_1347,N_120);
or U3429 (N_3429,N_2276,N_753);
or U3430 (N_3430,N_1084,N_49);
or U3431 (N_3431,N_2986,N_2351);
or U3432 (N_3432,N_1293,N_2192);
nand U3433 (N_3433,N_1042,N_1028);
or U3434 (N_3434,N_424,N_892);
nand U3435 (N_3435,N_477,N_2409);
nor U3436 (N_3436,N_1554,N_2279);
nor U3437 (N_3437,N_1502,N_2849);
or U3438 (N_3438,N_172,N_652);
xnor U3439 (N_3439,N_2484,N_1708);
nand U3440 (N_3440,N_2776,N_766);
nand U3441 (N_3441,N_1784,N_1832);
nand U3442 (N_3442,N_1358,N_1739);
nor U3443 (N_3443,N_2386,N_1802);
and U3444 (N_3444,N_604,N_182);
nor U3445 (N_3445,N_711,N_4);
nand U3446 (N_3446,N_1998,N_2482);
nand U3447 (N_3447,N_2567,N_1878);
nand U3448 (N_3448,N_2831,N_2842);
nor U3449 (N_3449,N_325,N_752);
xor U3450 (N_3450,N_1590,N_1845);
nor U3451 (N_3451,N_971,N_1993);
or U3452 (N_3452,N_926,N_442);
nand U3453 (N_3453,N_2068,N_1436);
nand U3454 (N_3454,N_351,N_2886);
or U3455 (N_3455,N_1953,N_2863);
and U3456 (N_3456,N_2799,N_672);
nand U3457 (N_3457,N_725,N_2479);
and U3458 (N_3458,N_355,N_2423);
nor U3459 (N_3459,N_1958,N_2081);
or U3460 (N_3460,N_2013,N_2237);
nand U3461 (N_3461,N_5,N_456);
or U3462 (N_3462,N_2274,N_1695);
nor U3463 (N_3463,N_2630,N_1515);
or U3464 (N_3464,N_935,N_1333);
nand U3465 (N_3465,N_2485,N_2753);
or U3466 (N_3466,N_545,N_1485);
nand U3467 (N_3467,N_1372,N_793);
and U3468 (N_3468,N_1674,N_2345);
nand U3469 (N_3469,N_345,N_62);
and U3470 (N_3470,N_414,N_1030);
and U3471 (N_3471,N_1865,N_429);
or U3472 (N_3472,N_464,N_2764);
nor U3473 (N_3473,N_901,N_1396);
and U3474 (N_3474,N_447,N_2623);
nor U3475 (N_3475,N_242,N_2710);
nor U3476 (N_3476,N_61,N_877);
xor U3477 (N_3477,N_1559,N_1798);
and U3478 (N_3478,N_1410,N_659);
nand U3479 (N_3479,N_2240,N_468);
or U3480 (N_3480,N_354,N_189);
nor U3481 (N_3481,N_2869,N_2649);
nand U3482 (N_3482,N_1919,N_1779);
nand U3483 (N_3483,N_489,N_407);
or U3484 (N_3484,N_968,N_1146);
nor U3485 (N_3485,N_755,N_214);
nor U3486 (N_3486,N_531,N_1526);
or U3487 (N_3487,N_432,N_2651);
xnor U3488 (N_3488,N_2578,N_1395);
nor U3489 (N_3489,N_2289,N_566);
nand U3490 (N_3490,N_1780,N_924);
or U3491 (N_3491,N_646,N_2955);
and U3492 (N_3492,N_2952,N_1239);
and U3493 (N_3493,N_2794,N_2384);
nand U3494 (N_3494,N_1989,N_1191);
and U3495 (N_3495,N_532,N_749);
and U3496 (N_3496,N_1634,N_2789);
xor U3497 (N_3497,N_1976,N_459);
nor U3498 (N_3498,N_326,N_990);
nor U3499 (N_3499,N_2114,N_1424);
nand U3500 (N_3500,N_1737,N_434);
nor U3501 (N_3501,N_1565,N_385);
or U3502 (N_3502,N_1987,N_1689);
nand U3503 (N_3503,N_2196,N_2411);
and U3504 (N_3504,N_2620,N_624);
or U3505 (N_3505,N_320,N_1574);
and U3506 (N_3506,N_198,N_2729);
nand U3507 (N_3507,N_123,N_2676);
nor U3508 (N_3508,N_1362,N_122);
and U3509 (N_3509,N_1097,N_2724);
and U3510 (N_3510,N_1013,N_25);
or U3511 (N_3511,N_2680,N_2643);
and U3512 (N_3512,N_119,N_2356);
or U3513 (N_3513,N_2543,N_929);
xnor U3514 (N_3514,N_2713,N_2981);
nand U3515 (N_3515,N_1584,N_2003);
nand U3516 (N_3516,N_2051,N_231);
nor U3517 (N_3517,N_785,N_1256);
xnor U3518 (N_3518,N_1620,N_2592);
xor U3519 (N_3519,N_2868,N_1099);
and U3520 (N_3520,N_89,N_1349);
nand U3521 (N_3521,N_1161,N_1703);
and U3522 (N_3522,N_1341,N_1272);
or U3523 (N_3523,N_2683,N_2613);
and U3524 (N_3524,N_777,N_1045);
xnor U3525 (N_3525,N_851,N_1785);
nor U3526 (N_3526,N_2721,N_1152);
nor U3527 (N_3527,N_1814,N_1318);
or U3528 (N_3528,N_1669,N_80);
nand U3529 (N_3529,N_520,N_583);
and U3530 (N_3530,N_2615,N_2441);
nand U3531 (N_3531,N_900,N_2238);
nand U3532 (N_3532,N_2392,N_2860);
nor U3533 (N_3533,N_746,N_2450);
xnor U3534 (N_3534,N_379,N_1527);
nor U3535 (N_3535,N_2704,N_1450);
or U3536 (N_3536,N_1154,N_112);
or U3537 (N_3537,N_342,N_28);
nand U3538 (N_3538,N_1433,N_1280);
xnor U3539 (N_3539,N_2258,N_959);
and U3540 (N_3540,N_658,N_2702);
and U3541 (N_3541,N_146,N_515);
or U3542 (N_3542,N_2534,N_2452);
or U3543 (N_3543,N_985,N_1126);
and U3544 (N_3544,N_2554,N_2716);
nor U3545 (N_3545,N_2012,N_772);
or U3546 (N_3546,N_2942,N_2442);
nand U3547 (N_3547,N_939,N_2747);
nor U3548 (N_3548,N_808,N_2165);
or U3549 (N_3549,N_2966,N_745);
nor U3550 (N_3550,N_1059,N_2318);
or U3551 (N_3551,N_2468,N_758);
nand U3552 (N_3552,N_2014,N_1166);
nand U3553 (N_3553,N_2655,N_2097);
or U3554 (N_3554,N_2248,N_74);
and U3555 (N_3555,N_1764,N_1419);
nand U3556 (N_3556,N_2967,N_364);
and U3557 (N_3557,N_2032,N_1065);
or U3558 (N_3558,N_244,N_2583);
nor U3559 (N_3559,N_2506,N_1456);
or U3560 (N_3560,N_2262,N_1778);
nor U3561 (N_3561,N_1806,N_2422);
or U3562 (N_3562,N_268,N_1541);
nand U3563 (N_3563,N_2179,N_629);
nor U3564 (N_3564,N_2692,N_2984);
nor U3565 (N_3565,N_2233,N_1334);
nor U3566 (N_3566,N_1378,N_1071);
nor U3567 (N_3567,N_1494,N_1795);
xnor U3568 (N_3568,N_2513,N_852);
xor U3569 (N_3569,N_650,N_578);
and U3570 (N_3570,N_1579,N_791);
nand U3571 (N_3571,N_248,N_2077);
and U3572 (N_3572,N_2424,N_1797);
nor U3573 (N_3573,N_693,N_315);
nand U3574 (N_3574,N_2375,N_419);
nand U3575 (N_3575,N_682,N_2618);
and U3576 (N_3576,N_85,N_2320);
and U3577 (N_3577,N_1183,N_541);
xnor U3578 (N_3578,N_961,N_544);
nor U3579 (N_3579,N_1761,N_1473);
and U3580 (N_3580,N_841,N_353);
and U3581 (N_3581,N_912,N_2975);
nand U3582 (N_3582,N_2516,N_1662);
or U3583 (N_3583,N_2092,N_2377);
nor U3584 (N_3584,N_384,N_630);
xor U3585 (N_3585,N_2918,N_2451);
nor U3586 (N_3586,N_498,N_1443);
xor U3587 (N_3587,N_70,N_2294);
and U3588 (N_3588,N_1903,N_2065);
xnor U3589 (N_3589,N_1257,N_2818);
nor U3590 (N_3590,N_874,N_1869);
or U3591 (N_3591,N_2074,N_1486);
nor U3592 (N_3592,N_2774,N_2964);
or U3593 (N_3593,N_280,N_2696);
nor U3594 (N_3594,N_999,N_2390);
nor U3595 (N_3595,N_864,N_747);
nand U3596 (N_3596,N_138,N_1892);
nand U3597 (N_3597,N_475,N_125);
and U3598 (N_3598,N_2584,N_603);
nor U3599 (N_3599,N_2189,N_569);
and U3600 (N_3600,N_2171,N_1151);
nand U3601 (N_3601,N_1452,N_675);
or U3602 (N_3602,N_2218,N_2697);
and U3603 (N_3603,N_2227,N_2775);
nor U3604 (N_3604,N_1027,N_1587);
or U3605 (N_3605,N_2347,N_651);
nand U3606 (N_3606,N_156,N_2909);
nor U3607 (N_3607,N_1996,N_2271);
nor U3608 (N_3608,N_482,N_1640);
or U3609 (N_3609,N_606,N_1270);
xor U3610 (N_3610,N_1453,N_1346);
and U3611 (N_3611,N_1611,N_1016);
nand U3612 (N_3612,N_2549,N_1353);
and U3613 (N_3613,N_2930,N_2087);
nand U3614 (N_3614,N_2517,N_100);
nor U3615 (N_3615,N_2083,N_1401);
or U3616 (N_3616,N_949,N_2969);
and U3617 (N_3617,N_22,N_441);
nor U3618 (N_3618,N_798,N_2904);
and U3619 (N_3619,N_763,N_1008);
nand U3620 (N_3620,N_2163,N_1117);
nor U3621 (N_3621,N_688,N_1950);
nor U3622 (N_3622,N_2113,N_2207);
nor U3623 (N_3623,N_1685,N_1466);
nand U3624 (N_3624,N_2151,N_2790);
or U3625 (N_3625,N_1102,N_1967);
nand U3626 (N_3626,N_2058,N_2847);
xor U3627 (N_3627,N_1416,N_1420);
and U3628 (N_3628,N_1986,N_1076);
and U3629 (N_3629,N_736,N_2209);
nor U3630 (N_3630,N_2670,N_2486);
or U3631 (N_3631,N_375,N_2144);
or U3632 (N_3632,N_1090,N_580);
and U3633 (N_3633,N_679,N_667);
and U3634 (N_3634,N_648,N_1907);
nand U3635 (N_3635,N_1604,N_1972);
and U3636 (N_3636,N_1661,N_2507);
or U3637 (N_3637,N_2228,N_669);
or U3638 (N_3638,N_1746,N_444);
and U3639 (N_3639,N_2203,N_1890);
and U3640 (N_3640,N_2172,N_2599);
and U3641 (N_3641,N_75,N_1673);
nand U3642 (N_3642,N_1221,N_418);
or U3643 (N_3643,N_1344,N_559);
or U3644 (N_3644,N_1870,N_1912);
and U3645 (N_3645,N_2822,N_815);
and U3646 (N_3646,N_1873,N_382);
nor U3647 (N_3647,N_596,N_2694);
xor U3648 (N_3648,N_584,N_1509);
and U3649 (N_3649,N_2326,N_726);
or U3650 (N_3650,N_694,N_1712);
nand U3651 (N_3651,N_760,N_139);
and U3652 (N_3652,N_2819,N_1301);
and U3653 (N_3653,N_91,N_2005);
and U3654 (N_3654,N_458,N_743);
xor U3655 (N_3655,N_1849,N_2474);
nor U3656 (N_3656,N_890,N_1262);
or U3657 (N_3657,N_2371,N_1465);
or U3658 (N_3658,N_2854,N_811);
and U3659 (N_3659,N_144,N_1299);
and U3660 (N_3660,N_1207,N_1477);
or U3661 (N_3661,N_210,N_943);
and U3662 (N_3662,N_2994,N_2522);
nand U3663 (N_3663,N_536,N_1639);
and U3664 (N_3664,N_2935,N_940);
nand U3665 (N_3665,N_1024,N_954);
nor U3666 (N_3666,N_1208,N_2382);
nor U3667 (N_3667,N_1875,N_1813);
or U3668 (N_3668,N_2914,N_344);
nand U3669 (N_3669,N_2418,N_2758);
and U3670 (N_3670,N_1243,N_2079);
xor U3671 (N_3671,N_417,N_2433);
nor U3672 (N_3672,N_945,N_1128);
or U3673 (N_3673,N_850,N_1781);
nand U3674 (N_3674,N_2496,N_835);
nor U3675 (N_3675,N_1467,N_262);
nor U3676 (N_3676,N_2283,N_1887);
nand U3677 (N_3677,N_1682,N_2581);
or U3678 (N_3678,N_2811,N_1949);
xor U3679 (N_3679,N_436,N_2902);
and U3680 (N_3680,N_1035,N_1918);
nand U3681 (N_3681,N_2071,N_1038);
and U3682 (N_3682,N_2557,N_2266);
or U3683 (N_3683,N_1384,N_1242);
and U3684 (N_3684,N_2536,N_2782);
nand U3685 (N_3685,N_2078,N_1791);
or U3686 (N_3686,N_1848,N_894);
nand U3687 (N_3687,N_2082,N_1343);
nor U3688 (N_3688,N_983,N_750);
nor U3689 (N_3689,N_2156,N_1687);
nand U3690 (N_3690,N_660,N_1286);
nor U3691 (N_3691,N_1656,N_1808);
and U3692 (N_3692,N_1178,N_1435);
nand U3693 (N_3693,N_1324,N_754);
and U3694 (N_3694,N_517,N_2405);
or U3695 (N_3695,N_505,N_1799);
and U3696 (N_3696,N_2021,N_548);
nor U3697 (N_3697,N_147,N_16);
and U3698 (N_3698,N_673,N_1734);
or U3699 (N_3699,N_2761,N_1553);
and U3700 (N_3700,N_235,N_2417);
nor U3701 (N_3701,N_2829,N_2341);
and U3702 (N_3702,N_1997,N_622);
nor U3703 (N_3703,N_788,N_2577);
or U3704 (N_3704,N_1534,N_920);
nand U3705 (N_3705,N_2314,N_1231);
nor U3706 (N_3706,N_1364,N_1153);
and U3707 (N_3707,N_6,N_169);
nor U3708 (N_3708,N_641,N_732);
and U3709 (N_3709,N_457,N_133);
or U3710 (N_3710,N_1759,N_1664);
and U3711 (N_3711,N_142,N_2132);
nand U3712 (N_3712,N_2629,N_2261);
and U3713 (N_3713,N_1264,N_2920);
nor U3714 (N_3714,N_1484,N_1385);
and U3715 (N_3715,N_2478,N_427);
nand U3716 (N_3716,N_1002,N_2357);
and U3717 (N_3717,N_328,N_2275);
nand U3718 (N_3718,N_56,N_771);
and U3719 (N_3719,N_508,N_2893);
xor U3720 (N_3720,N_1185,N_2797);
nor U3721 (N_3721,N_2915,N_1969);
xor U3722 (N_3722,N_1020,N_1121);
nand U3723 (N_3723,N_1376,N_1524);
nor U3724 (N_3724,N_2674,N_870);
xnor U3725 (N_3725,N_2565,N_1397);
nor U3726 (N_3726,N_2851,N_2383);
xor U3727 (N_3727,N_431,N_2865);
nor U3728 (N_3728,N_1294,N_313);
and U3729 (N_3729,N_922,N_409);
or U3730 (N_3730,N_982,N_655);
or U3731 (N_3731,N_2740,N_691);
nor U3732 (N_3732,N_553,N_790);
xor U3733 (N_3733,N_2462,N_2426);
nor U3734 (N_3734,N_1198,N_1926);
nor U3735 (N_3735,N_2296,N_421);
nor U3736 (N_3736,N_2010,N_633);
or U3737 (N_3737,N_2458,N_1866);
nand U3738 (N_3738,N_143,N_363);
nor U3739 (N_3739,N_2061,N_696);
or U3740 (N_3740,N_1036,N_2752);
nor U3741 (N_3741,N_1599,N_577);
and U3742 (N_3742,N_1568,N_1085);
nor U3743 (N_3743,N_126,N_1563);
nor U3744 (N_3744,N_582,N_2463);
nor U3745 (N_3745,N_1619,N_2225);
nand U3746 (N_3746,N_104,N_1716);
nor U3747 (N_3747,N_1069,N_820);
nor U3748 (N_3748,N_234,N_2365);
nand U3749 (N_3749,N_1255,N_2118);
nor U3750 (N_3750,N_2748,N_2033);
nand U3751 (N_3751,N_2576,N_2470);
nor U3752 (N_3752,N_1704,N_1867);
nand U3753 (N_3753,N_609,N_1388);
or U3754 (N_3754,N_509,N_1223);
nand U3755 (N_3755,N_863,N_2568);
nand U3756 (N_3756,N_881,N_538);
nand U3757 (N_3757,N_1829,N_575);
nand U3758 (N_3758,N_818,N_1860);
nor U3759 (N_3759,N_2300,N_2945);
nor U3760 (N_3760,N_2299,N_435);
or U3761 (N_3761,N_2977,N_2353);
nor U3762 (N_3762,N_2897,N_1246);
xnor U3763 (N_3763,N_1615,N_1981);
nand U3764 (N_3764,N_1359,N_591);
nor U3765 (N_3765,N_1311,N_967);
nand U3766 (N_3766,N_105,N_2190);
nor U3767 (N_3767,N_1252,N_1211);
nor U3768 (N_3768,N_1715,N_689);
nor U3769 (N_3769,N_2786,N_2636);
or U3770 (N_3770,N_1284,N_58);
and U3771 (N_3771,N_2848,N_1403);
nor U3772 (N_3772,N_2770,N_738);
nand U3773 (N_3773,N_378,N_306);
and U3774 (N_3774,N_2471,N_2205);
nand U3775 (N_3775,N_393,N_802);
or U3776 (N_3776,N_951,N_1925);
or U3777 (N_3777,N_1811,N_706);
and U3778 (N_3778,N_2531,N_2185);
nor U3779 (N_3779,N_1168,N_2687);
nand U3780 (N_3780,N_1520,N_440);
and U3781 (N_3781,N_2219,N_1850);
or U3782 (N_3782,N_1147,N_2401);
xor U3783 (N_3783,N_2378,N_2723);
and U3784 (N_3784,N_1616,N_1754);
nor U3785 (N_3785,N_1786,N_2879);
nand U3786 (N_3786,N_2473,N_1271);
nor U3787 (N_3787,N_1303,N_184);
and U3788 (N_3788,N_1060,N_1220);
nand U3789 (N_3789,N_768,N_2511);
and U3790 (N_3790,N_1457,N_2948);
nor U3791 (N_3791,N_1009,N_857);
and U3792 (N_3792,N_866,N_1672);
nor U3793 (N_3793,N_240,N_1539);
and U3794 (N_3794,N_783,N_795);
and U3795 (N_3795,N_2675,N_1556);
nand U3796 (N_3796,N_1970,N_643);
nand U3797 (N_3797,N_2363,N_875);
or U3798 (N_3798,N_1500,N_29);
or U3799 (N_3799,N_1184,N_1824);
nand U3800 (N_3800,N_963,N_2204);
xor U3801 (N_3801,N_1598,N_1751);
nor U3802 (N_3802,N_781,N_1638);
xor U3803 (N_3803,N_1868,N_1468);
nand U3804 (N_3804,N_1052,N_991);
nor U3805 (N_3805,N_1441,N_2709);
nor U3806 (N_3806,N_2727,N_965);
and U3807 (N_3807,N_907,N_1331);
xnor U3808 (N_3808,N_1533,N_193);
and U3809 (N_3809,N_1577,N_593);
nand U3810 (N_3810,N_1019,N_1697);
or U3811 (N_3811,N_2973,N_2342);
nand U3812 (N_3812,N_1725,N_2229);
or U3813 (N_3813,N_1637,N_1901);
nor U3814 (N_3814,N_175,N_1900);
nor U3815 (N_3815,N_73,N_1254);
and U3816 (N_3816,N_1155,N_2521);
nor U3817 (N_3817,N_2040,N_632);
nand U3818 (N_3818,N_408,N_2816);
or U3819 (N_3819,N_2399,N_1537);
nand U3820 (N_3820,N_168,N_1792);
nor U3821 (N_3821,N_1142,N_627);
nand U3822 (N_3822,N_2635,N_1351);
and U3823 (N_3823,N_1602,N_233);
or U3824 (N_3824,N_1437,N_812);
and U3825 (N_3825,N_2929,N_1267);
xor U3826 (N_3826,N_845,N_1305);
nor U3827 (N_3827,N_2169,N_365);
xnor U3828 (N_3828,N_2152,N_2119);
and U3829 (N_3829,N_2957,N_824);
or U3830 (N_3830,N_1309,N_1523);
nand U3831 (N_3831,N_899,N_2677);
nand U3832 (N_3832,N_1636,N_23);
or U3833 (N_3833,N_1226,N_343);
and U3834 (N_3834,N_1159,N_2459);
nand U3835 (N_3835,N_2622,N_2604);
nand U3836 (N_3836,N_765,N_1400);
nand U3837 (N_3837,N_1948,N_256);
or U3838 (N_3838,N_2621,N_1782);
and U3839 (N_3839,N_2472,N_278);
and U3840 (N_3840,N_680,N_903);
or U3841 (N_3841,N_997,N_976);
and U3842 (N_3842,N_2693,N_1050);
nand U3843 (N_3843,N_1490,N_34);
xnor U3844 (N_3844,N_2142,N_2381);
nor U3845 (N_3845,N_40,N_71);
and U3846 (N_3846,N_1670,N_1077);
xor U3847 (N_3847,N_2094,N_1422);
nor U3848 (N_3848,N_2336,N_778);
or U3849 (N_3849,N_367,N_2416);
or U3850 (N_3850,N_187,N_832);
xor U3851 (N_3851,N_269,N_1586);
nand U3852 (N_3852,N_1210,N_1105);
or U3853 (N_3853,N_69,N_885);
xnor U3854 (N_3854,N_516,N_1906);
nor U3855 (N_3855,N_2881,N_1793);
xor U3856 (N_3856,N_1004,N_1897);
nor U3857 (N_3857,N_1947,N_2055);
or U3858 (N_3858,N_130,N_2603);
and U3859 (N_3859,N_2657,N_2788);
nand U3860 (N_3860,N_2688,N_1601);
nor U3861 (N_3861,N_118,N_1338);
xor U3862 (N_3862,N_511,N_911);
and U3863 (N_3863,N_1883,N_2023);
or U3864 (N_3864,N_514,N_1549);
xnor U3865 (N_3865,N_1807,N_1825);
nor U3866 (N_3866,N_942,N_1818);
nand U3867 (N_3867,N_1086,N_211);
nand U3868 (N_3868,N_1083,N_2112);
and U3869 (N_3869,N_2431,N_1288);
and U3870 (N_3870,N_510,N_2792);
nand U3871 (N_3871,N_1655,N_1562);
nor U3872 (N_3872,N_157,N_2906);
xor U3873 (N_3873,N_1566,N_988);
or U3874 (N_3874,N_1546,N_463);
and U3875 (N_3875,N_1580,N_2759);
or U3876 (N_3876,N_1628,N_764);
nand U3877 (N_3877,N_1233,N_707);
and U3878 (N_3878,N_2111,N_2846);
and U3879 (N_3879,N_1145,N_1115);
nand U3880 (N_3880,N_1743,N_917);
nor U3881 (N_3881,N_1633,N_797);
nand U3882 (N_3882,N_904,N_2492);
nor U3883 (N_3883,N_1413,N_490);
and U3884 (N_3884,N_809,N_3);
and U3885 (N_3885,N_1224,N_2661);
nand U3886 (N_3886,N_2480,N_1329);
nor U3887 (N_3887,N_2787,N_2054);
nand U3888 (N_3888,N_2625,N_642);
nand U3889 (N_3889,N_2208,N_2285);
or U3890 (N_3890,N_2202,N_2095);
and U3891 (N_3891,N_340,N_2783);
or U3892 (N_3892,N_1858,N_1724);
and U3893 (N_3893,N_1552,N_1719);
xor U3894 (N_3894,N_2571,N_470);
and U3895 (N_3895,N_433,N_2429);
and U3896 (N_3896,N_108,N_392);
or U3897 (N_3897,N_1162,N_2679);
xnor U3898 (N_3898,N_941,N_2340);
nand U3899 (N_3899,N_979,N_1165);
and U3900 (N_3900,N_1360,N_933);
nand U3901 (N_3901,N_2582,N_1677);
nor U3902 (N_3902,N_928,N_1496);
nand U3903 (N_3903,N_2495,N_2376);
xnor U3904 (N_3904,N_2259,N_2292);
xor U3905 (N_3905,N_1709,N_1068);
xnor U3906 (N_3906,N_2180,N_1114);
or U3907 (N_3907,N_1449,N_552);
and U3908 (N_3908,N_333,N_1511);
or U3909 (N_3909,N_1458,N_1313);
and U3910 (N_3910,N_2272,N_1375);
and U3911 (N_3911,N_285,N_1043);
and U3912 (N_3912,N_478,N_272);
nor U3913 (N_3913,N_1363,N_2230);
or U3914 (N_3914,N_1193,N_227);
nand U3915 (N_3915,N_220,N_1891);
nor U3916 (N_3916,N_2735,N_579);
nor U3917 (N_3917,N_2212,N_2956);
nand U3918 (N_3918,N_2737,N_663);
nand U3919 (N_3919,N_597,N_1175);
and U3920 (N_3920,N_2444,N_2368);
nand U3921 (N_3921,N_1190,N_275);
nor U3922 (N_3922,N_1679,N_1200);
nor U3923 (N_3923,N_1585,N_1718);
nor U3924 (N_3924,N_1075,N_1073);
and U3925 (N_3925,N_2921,N_908);
or U3926 (N_3926,N_2239,N_1370);
nand U3927 (N_3927,N_761,N_1464);
nand U3928 (N_3928,N_1072,N_1690);
and U3929 (N_3929,N_2793,N_2587);
nor U3930 (N_3930,N_895,N_2366);
nor U3931 (N_3931,N_1946,N_2830);
nor U3932 (N_3932,N_2380,N_2264);
nand U3933 (N_3933,N_391,N_2004);
nor U3934 (N_3934,N_2198,N_2039);
nand U3935 (N_3935,N_2800,N_980);
or U3936 (N_3936,N_2085,N_310);
nand U3937 (N_3937,N_813,N_1194);
xnor U3938 (N_3938,N_2950,N_2750);
and U3939 (N_3939,N_1648,N_2664);
and U3940 (N_3940,N_1357,N_136);
nand U3941 (N_3941,N_2027,N_2247);
nand U3942 (N_3942,N_309,N_2338);
nand U3943 (N_3943,N_2049,N_2993);
or U3944 (N_3944,N_1265,N_1366);
xor U3945 (N_3945,N_970,N_2217);
nor U3946 (N_3946,N_2159,N_2350);
and U3947 (N_3947,N_1170,N_2241);
or U3948 (N_3948,N_662,N_2617);
and U3949 (N_3949,N_876,N_2890);
xor U3950 (N_3950,N_891,N_290);
and U3951 (N_3951,N_1700,N_2147);
and U3952 (N_3952,N_731,N_297);
nand U3953 (N_3953,N_47,N_1744);
or U3954 (N_3954,N_2880,N_1390);
or U3955 (N_3955,N_1592,N_2691);
and U3956 (N_3956,N_1840,N_381);
nand U3957 (N_3957,N_2923,N_2475);
nand U3958 (N_3958,N_865,N_2214);
nor U3959 (N_3959,N_301,N_1532);
and U3960 (N_3960,N_998,N_1653);
nor U3961 (N_3961,N_261,N_716);
xnor U3962 (N_3962,N_2550,N_555);
nor U3963 (N_3963,N_1003,N_1319);
nor U3964 (N_3964,N_2707,N_1699);
nor U3965 (N_3965,N_2002,N_93);
nor U3966 (N_3966,N_1268,N_1021);
nand U3967 (N_3967,N_1529,N_174);
and U3968 (N_3968,N_274,N_2968);
and U3969 (N_3969,N_2510,N_1314);
nand U3970 (N_3970,N_2895,N_1756);
and U3971 (N_3971,N_993,N_1514);
nand U3972 (N_3972,N_1727,N_2718);
nor U3973 (N_3973,N_1310,N_2174);
or U3974 (N_3974,N_810,N_1321);
nor U3975 (N_3975,N_1491,N_1735);
or U3976 (N_3976,N_502,N_173);
nand U3977 (N_3977,N_551,N_1144);
nor U3978 (N_3978,N_2963,N_2959);
xor U3979 (N_3979,N_2303,N_718);
and U3980 (N_3980,N_1157,N_714);
nor U3981 (N_3981,N_1983,N_871);
or U3982 (N_3982,N_1569,N_1924);
or U3983 (N_3983,N_2226,N_2524);
nor U3984 (N_3984,N_1447,N_247);
or U3985 (N_3985,N_560,N_1510);
and U3986 (N_3986,N_1354,N_2280);
nand U3987 (N_3987,N_1821,N_291);
and U3988 (N_3988,N_2500,N_2037);
or U3989 (N_3989,N_674,N_1196);
nor U3990 (N_3990,N_880,N_1480);
nor U3991 (N_3991,N_2855,N_2298);
nand U3992 (N_3992,N_2526,N_2933);
nand U3993 (N_3993,N_1361,N_1098);
nand U3994 (N_3994,N_2627,N_838);
xnor U3995 (N_3995,N_1606,N_2512);
nand U3996 (N_3996,N_453,N_1225);
or U3997 (N_3997,N_683,N_331);
or U3998 (N_3998,N_1048,N_2658);
xor U3999 (N_3999,N_2105,N_708);
nand U4000 (N_4000,N_661,N_483);
and U4001 (N_4001,N_1942,N_1755);
nand U4002 (N_4002,N_794,N_2438);
nand U4003 (N_4003,N_307,N_1582);
xnor U4004 (N_4004,N_1736,N_2316);
or U4005 (N_4005,N_18,N_2857);
and U4006 (N_4006,N_2440,N_640);
nand U4007 (N_4007,N_53,N_449);
nand U4008 (N_4008,N_46,N_92);
or U4009 (N_4009,N_1091,N_1729);
or U4010 (N_4010,N_1158,N_861);
nand U4011 (N_4011,N_2982,N_110);
nand U4012 (N_4012,N_2763,N_395);
nand U4013 (N_4013,N_203,N_543);
xor U4014 (N_4014,N_595,N_1921);
and U4015 (N_4015,N_2385,N_1474);
and U4016 (N_4016,N_1368,N_2319);
nor U4017 (N_4017,N_2689,N_1960);
and U4018 (N_4018,N_305,N_2765);
or U4019 (N_4019,N_522,N_1439);
xnor U4020 (N_4020,N_1757,N_97);
or U4021 (N_4021,N_2080,N_1481);
nor U4022 (N_4022,N_2953,N_2637);
xor U4023 (N_4023,N_519,N_2736);
and U4024 (N_4024,N_2943,N_728);
nand U4025 (N_4025,N_1597,N_1497);
or U4026 (N_4026,N_2874,N_2876);
xnor U4027 (N_4027,N_1564,N_1479);
and U4028 (N_4028,N_2158,N_2404);
and U4029 (N_4029,N_571,N_2726);
and U4030 (N_4030,N_914,N_205);
nor U4031 (N_4031,N_590,N_2882);
and U4032 (N_4032,N_1614,N_2315);
and U4033 (N_4033,N_1289,N_21);
or U4034 (N_4034,N_2542,N_827);
nand U4035 (N_4035,N_2912,N_1082);
nand U4036 (N_4036,N_730,N_1017);
or U4037 (N_4037,N_2757,N_2334);
and U4038 (N_4038,N_1444,N_1489);
nor U4039 (N_4039,N_2278,N_1543);
or U4040 (N_4040,N_485,N_685);
and U4041 (N_4041,N_1963,N_2412);
nor U4042 (N_4042,N_1111,N_2028);
nand U4043 (N_4043,N_647,N_2596);
nand U4044 (N_4044,N_1941,N_398);
or U4045 (N_4045,N_2302,N_773);
nor U4046 (N_4046,N_2139,N_1693);
nand U4047 (N_4047,N_1745,N_2989);
or U4048 (N_4048,N_1337,N_2176);
and U4049 (N_4049,N_2145,N_2780);
nor U4050 (N_4050,N_2311,N_844);
and U4051 (N_4051,N_2971,N_2410);
or U4052 (N_4052,N_225,N_1291);
nor U4053 (N_4053,N_1096,N_1681);
nor U4054 (N_4054,N_1394,N_2199);
and U4055 (N_4055,N_2913,N_534);
or U4056 (N_4056,N_525,N_352);
nor U4057 (N_4057,N_1451,N_1049);
xnor U4058 (N_4058,N_1423,N_415);
nand U4059 (N_4059,N_2714,N_321);
nor U4060 (N_4060,N_1742,N_102);
or U4061 (N_4061,N_1688,N_1323);
nor U4062 (N_4062,N_1747,N_1773);
or U4063 (N_4063,N_204,N_2236);
nor U4064 (N_4064,N_1833,N_2644);
and U4065 (N_4065,N_2563,N_1847);
and U4066 (N_4066,N_284,N_2432);
and U4067 (N_4067,N_1517,N_1665);
nand U4068 (N_4068,N_1842,N_386);
nand U4069 (N_4069,N_213,N_425);
nor U4070 (N_4070,N_2798,N_2234);
xor U4071 (N_4071,N_956,N_2195);
nor U4072 (N_4072,N_2091,N_422);
nor U4073 (N_4073,N_243,N_2632);
or U4074 (N_4074,N_267,N_1542);
and U4075 (N_4075,N_19,N_2924);
and U4076 (N_4076,N_2265,N_2944);
or U4077 (N_4077,N_208,N_769);
nand U4078 (N_4078,N_2249,N_2708);
or U4079 (N_4079,N_527,N_2313);
or U4080 (N_4080,N_471,N_898);
nand U4081 (N_4081,N_1022,N_739);
and U4082 (N_4082,N_2251,N_1964);
or U4083 (N_4083,N_469,N_723);
xnor U4084 (N_4084,N_2454,N_2101);
nor U4085 (N_4085,N_1857,N_2946);
nor U4086 (N_4086,N_2374,N_910);
nor U4087 (N_4087,N_2564,N_2324);
or U4088 (N_4088,N_380,N_2744);
xnor U4089 (N_4089,N_2872,N_1823);
nor U4090 (N_4090,N_513,N_1775);
nand U4091 (N_4091,N_292,N_1731);
or U4092 (N_4092,N_221,N_975);
nand U4093 (N_4093,N_893,N_2024);
xor U4094 (N_4094,N_20,N_1862);
and U4095 (N_4095,N_2348,N_2332);
nor U4096 (N_4096,N_2453,N_1506);
or U4097 (N_4097,N_155,N_1812);
and U4098 (N_4098,N_229,N_1507);
or U4099 (N_4099,N_2393,N_403);
or U4100 (N_4100,N_1136,N_1127);
or U4101 (N_4101,N_1995,N_814);
xor U4102 (N_4102,N_2821,N_2528);
or U4103 (N_4103,N_1315,N_1459);
nand U4104 (N_4104,N_2810,N_347);
nand U4105 (N_4105,N_1898,N_2408);
nand U4106 (N_4106,N_466,N_599);
nor U4107 (N_4107,N_311,N_2666);
nand U4108 (N_4108,N_2665,N_1701);
and U4109 (N_4109,N_932,N_2041);
and U4110 (N_4110,N_238,N_2889);
nand U4111 (N_4111,N_2398,N_654);
nand U4112 (N_4112,N_1899,N_888);
or U4113 (N_4113,N_873,N_1844);
nor U4114 (N_4114,N_2035,N_2270);
or U4115 (N_4115,N_2887,N_1046);
nor U4116 (N_4116,N_1914,N_1927);
nand U4117 (N_4117,N_2987,N_668);
nor U4118 (N_4118,N_2551,N_2850);
nand U4119 (N_4119,N_2428,N_1051);
nor U4120 (N_4120,N_300,N_821);
nor U4121 (N_4121,N_1991,N_2026);
and U4122 (N_4122,N_1740,N_2489);
nand U4123 (N_4123,N_2245,N_2712);
xor U4124 (N_4124,N_834,N_2008);
and U4125 (N_4125,N_2460,N_1839);
and U4126 (N_4126,N_847,N_567);
or U4127 (N_4127,N_98,N_1248);
nor U4128 (N_4128,N_2685,N_48);
and U4129 (N_4129,N_2905,N_2161);
nor U4130 (N_4130,N_664,N_1325);
nor U4131 (N_4131,N_2585,N_59);
xnor U4132 (N_4132,N_792,N_2403);
nand U4133 (N_4133,N_2153,N_2781);
and U4134 (N_4134,N_2908,N_2853);
nand U4135 (N_4135,N_602,N_2400);
xnor U4136 (N_4136,N_878,N_1192);
nor U4137 (N_4137,N_1600,N_1905);
xor U4138 (N_4138,N_684,N_2745);
nand U4139 (N_4139,N_1959,N_1179);
and U4140 (N_4140,N_1276,N_265);
xnor U4141 (N_4141,N_2067,N_283);
nor U4142 (N_4142,N_1143,N_1530);
xor U4143 (N_4143,N_1012,N_1726);
nand U4144 (N_4144,N_2116,N_2742);
and U4145 (N_4145,N_148,N_2109);
or U4146 (N_4146,N_705,N_610);
nand U4147 (N_4147,N_1796,N_2601);
and U4148 (N_4148,N_2166,N_796);
or U4149 (N_4149,N_2885,N_389);
or U4150 (N_4150,N_2352,N_2146);
nand U4151 (N_4151,N_1160,N_45);
or U4152 (N_4152,N_1195,N_2660);
xnor U4153 (N_4153,N_2864,N_1463);
nor U4154 (N_4154,N_2,N_1025);
nor U4155 (N_4155,N_849,N_692);
and U4156 (N_4156,N_2631,N_1213);
and U4157 (N_4157,N_1881,N_1937);
and U4158 (N_4158,N_2242,N_2932);
nor U4159 (N_4159,N_487,N_2036);
or U4160 (N_4160,N_1230,N_842);
nor U4161 (N_4161,N_1212,N_2297);
and U4162 (N_4162,N_323,N_2260);
or U4163 (N_4163,N_374,N_613);
nand U4164 (N_4164,N_2191,N_2836);
nor U4165 (N_4165,N_1557,N_405);
nand U4166 (N_4166,N_1222,N_2961);
nand U4167 (N_4167,N_317,N_2031);
or U4168 (N_4168,N_127,N_576);
or U4169 (N_4169,N_565,N_1612);
or U4170 (N_4170,N_2867,N_1909);
and U4171 (N_4171,N_2648,N_2640);
and U4172 (N_4172,N_1499,N_103);
xor U4173 (N_4173,N_1805,N_2001);
or U4174 (N_4174,N_202,N_2044);
and U4175 (N_4175,N_2038,N_2177);
nor U4176 (N_4176,N_2481,N_701);
or U4177 (N_4177,N_1461,N_1089);
nor U4178 (N_4178,N_639,N_294);
xnor U4179 (N_4179,N_2150,N_111);
and U4180 (N_4180,N_2154,N_1391);
nor U4181 (N_4181,N_1596,N_1752);
and U4182 (N_4182,N_2045,N_1377);
or U4183 (N_4183,N_1274,N_616);
nor U4184 (N_4184,N_530,N_2626);
or U4185 (N_4185,N_1431,N_51);
xnor U4186 (N_4186,N_2043,N_1660);
and U4187 (N_4187,N_215,N_2896);
and U4188 (N_4188,N_1547,N_2769);
and U4189 (N_4189,N_594,N_564);
and U4190 (N_4190,N_2633,N_2477);
nor U4191 (N_4191,N_1110,N_230);
nor U4192 (N_4192,N_782,N_2875);
nand U4193 (N_4193,N_2834,N_2157);
nor U4194 (N_4194,N_2841,N_1680);
nor U4195 (N_4195,N_2443,N_2108);
nand U4196 (N_4196,N_2958,N_1545);
nand U4197 (N_4197,N_209,N_2650);
xor U4198 (N_4198,N_2255,N_9);
nand U4199 (N_4199,N_357,N_2559);
and U4200 (N_4200,N_619,N_2090);
nand U4201 (N_4201,N_2647,N_2354);
nand U4202 (N_4202,N_199,N_492);
and U4203 (N_4203,N_1952,N_1421);
nor U4204 (N_4204,N_1169,N_1888);
and U4205 (N_4205,N_273,N_1040);
nor U4206 (N_4206,N_2123,N_2455);
and U4207 (N_4207,N_2652,N_149);
nor U4208 (N_4208,N_1148,N_324);
xor U4209 (N_4209,N_801,N_1355);
and U4210 (N_4210,N_1728,N_1476);
nand U4211 (N_4211,N_2690,N_2983);
or U4212 (N_4212,N_2515,N_1249);
and U4213 (N_4213,N_1774,N_2253);
or U4214 (N_4214,N_2048,N_886);
and U4215 (N_4215,N_537,N_1852);
or U4216 (N_4216,N_936,N_2700);
and U4217 (N_4217,N_2149,N_1714);
and U4218 (N_4218,N_592,N_1445);
nor U4219 (N_4219,N_281,N_1425);
nor U4220 (N_4220,N_2508,N_1047);
nor U4221 (N_4221,N_2698,N_131);
or U4222 (N_4222,N_1238,N_2586);
and U4223 (N_4223,N_1282,N_1187);
nor U4224 (N_4224,N_1531,N_670);
nor U4225 (N_4225,N_1011,N_135);
xnor U4226 (N_4226,N_2137,N_41);
xnor U4227 (N_4227,N_776,N_1721);
xor U4228 (N_4228,N_2427,N_2420);
or U4229 (N_4229,N_2609,N_931);
and U4230 (N_4230,N_953,N_190);
nand U4231 (N_4231,N_2858,N_1575);
nor U4232 (N_4232,N_1536,N_2919);
nand U4233 (N_4233,N_2619,N_2333);
and U4234 (N_4234,N_2419,N_36);
or U4235 (N_4235,N_2560,N_423);
nand U4236 (N_4236,N_1561,N_563);
nor U4237 (N_4237,N_512,N_2178);
nor U4238 (N_4238,N_2892,N_2931);
nand U4239 (N_4239,N_1326,N_840);
xor U4240 (N_4240,N_2572,N_2464);
nand U4241 (N_4241,N_1283,N_2490);
and U4242 (N_4242,N_1327,N_404);
and U4243 (N_4243,N_1593,N_94);
xor U4244 (N_4244,N_428,N_2273);
nand U4245 (N_4245,N_158,N_2642);
or U4246 (N_4246,N_2839,N_140);
or U4247 (N_4247,N_2018,N_2611);
nand U4248 (N_4248,N_948,N_1336);
or U4249 (N_4249,N_2824,N_2614);
nor U4250 (N_4250,N_2720,N_1317);
nor U4251 (N_4251,N_2434,N_288);
and U4252 (N_4252,N_1809,N_957);
nand U4253 (N_4253,N_481,N_1492);
and U4254 (N_4254,N_2295,N_2130);
and U4255 (N_4255,N_2194,N_2367);
and U4256 (N_4256,N_2389,N_2671);
nor U4257 (N_4257,N_1512,N_2901);
and U4258 (N_4258,N_196,N_1087);
and U4259 (N_4259,N_869,N_2922);
and U4260 (N_4260,N_2461,N_219);
nand U4261 (N_4261,N_2840,N_635);
nand U4262 (N_4262,N_862,N_2767);
and U4263 (N_4263,N_1855,N_2307);
or U4264 (N_4264,N_2656,N_618);
nand U4265 (N_4265,N_2000,N_356);
and U4266 (N_4266,N_217,N_1237);
nand U4267 (N_4267,N_2349,N_1130);
or U4268 (N_4268,N_1100,N_420);
xor U4269 (N_4269,N_2073,N_2476);
nor U4270 (N_4270,N_2705,N_1920);
xor U4271 (N_4271,N_266,N_780);
and U4272 (N_4272,N_1692,N_2884);
and U4273 (N_4273,N_370,N_1015);
xnor U4274 (N_4274,N_2616,N_805);
nand U4275 (N_4275,N_1893,N_930);
nor U4276 (N_4276,N_15,N_717);
nor U4277 (N_4277,N_1733,N_677);
and U4278 (N_4278,N_2539,N_2910);
or U4279 (N_4279,N_2927,N_2456);
or U4280 (N_4280,N_829,N_598);
and U4281 (N_4281,N_38,N_1826);
and U4282 (N_4282,N_2773,N_1876);
xnor U4283 (N_4283,N_839,N_1896);
or U4284 (N_4284,N_83,N_1837);
and U4285 (N_4285,N_2743,N_2064);
or U4286 (N_4286,N_81,N_1061);
nor U4287 (N_4287,N_2762,N_987);
xnor U4288 (N_4288,N_2201,N_2321);
and U4289 (N_4289,N_859,N_161);
nand U4290 (N_4290,N_170,N_298);
and U4291 (N_4291,N_1783,N_1259);
nand U4292 (N_4292,N_698,N_2701);
nor U4293 (N_4293,N_349,N_14);
nor U4294 (N_4294,N_2312,N_774);
nor U4295 (N_4295,N_2825,N_31);
or U4296 (N_4296,N_702,N_2659);
or U4297 (N_4297,N_722,N_410);
nand U4298 (N_4298,N_1884,N_1241);
or U4299 (N_4299,N_129,N_1917);
nor U4300 (N_4300,N_2947,N_2449);
and U4301 (N_4301,N_803,N_2859);
and U4302 (N_4302,N_2605,N_1691);
and U4303 (N_4303,N_2128,N_2143);
nor U4304 (N_4304,N_1164,N_2244);
xnor U4305 (N_4305,N_909,N_1295);
xor U4306 (N_4306,N_1482,N_681);
and U4307 (N_4307,N_1340,N_676);
or U4308 (N_4308,N_450,N_1717);
nor U4309 (N_4309,N_299,N_919);
or U4310 (N_4310,N_2739,N_1478);
nand U4311 (N_4311,N_115,N_334);
nor U4312 (N_4312,N_2801,N_2466);
nand U4313 (N_4313,N_1889,N_946);
nand U4314 (N_4314,N_2833,N_186);
nand U4315 (N_4315,N_2256,N_1851);
xor U4316 (N_4316,N_1521,N_1880);
or U4317 (N_4317,N_2501,N_915);
xor U4318 (N_4318,N_430,N_572);
or U4319 (N_4319,N_1263,N_1430);
or U4320 (N_4320,N_1854,N_2497);
or U4321 (N_4321,N_282,N_1409);
and U4322 (N_4322,N_1215,N_2556);
and U4323 (N_4323,N_913,N_2870);
nand U4324 (N_4324,N_1006,N_2911);
nand U4325 (N_4325,N_188,N_1980);
or U4326 (N_4326,N_2548,N_339);
xnor U4327 (N_4327,N_826,N_952);
nand U4328 (N_4328,N_1429,N_2591);
or U4329 (N_4329,N_2628,N_2715);
nor U4330 (N_4330,N_906,N_1387);
and U4331 (N_4331,N_2731,N_2102);
nand U4332 (N_4332,N_2805,N_2815);
or U4333 (N_4333,N_787,N_1944);
nor U4334 (N_4334,N_1079,N_825);
and U4335 (N_4335,N_2634,N_1296);
or U4336 (N_4336,N_556,N_151);
and U4337 (N_4337,N_2277,N_1934);
or U4338 (N_4338,N_1965,N_2965);
and U4339 (N_4339,N_496,N_2807);
nor U4340 (N_4340,N_562,N_2362);
and U4341 (N_4341,N_2760,N_2060);
and U4342 (N_4342,N_2494,N_518);
nand U4343 (N_4343,N_1129,N_1471);
nand U4344 (N_4344,N_986,N_1571);
and U4345 (N_4345,N_50,N_1209);
and U4346 (N_4346,N_879,N_1228);
nand U4347 (N_4347,N_1174,N_2907);
and U4348 (N_4348,N_176,N_1667);
or U4349 (N_4349,N_2796,N_1623);
nor U4350 (N_4350,N_2009,N_246);
and U4351 (N_4351,N_996,N_2785);
nand U4352 (N_4352,N_974,N_2421);
xor U4353 (N_4353,N_1588,N_2007);
nor U4354 (N_4354,N_55,N_1417);
nor U4355 (N_4355,N_2503,N_2487);
or U4356 (N_4356,N_528,N_302);
nor U4357 (N_4357,N_1804,N_396);
nor U4358 (N_4358,N_264,N_735);
and U4359 (N_4359,N_1846,N_166);
nor U4360 (N_4360,N_2167,N_2610);
and U4361 (N_4361,N_1119,N_733);
nor U4362 (N_4362,N_167,N_1163);
nand U4363 (N_4363,N_1149,N_1961);
and U4364 (N_4364,N_897,N_816);
or U4365 (N_4365,N_271,N_178);
nand U4366 (N_4366,N_2291,N_1613);
or U4367 (N_4367,N_1625,N_1197);
nor U4368 (N_4368,N_2335,N_279);
nand U4369 (N_4369,N_473,N_2937);
nand U4370 (N_4370,N_2155,N_304);
or U4371 (N_4371,N_2263,N_700);
and U4372 (N_4372,N_1904,N_2835);
or U4373 (N_4373,N_2624,N_455);
or U4374 (N_4374,N_1908,N_1760);
nand U4375 (N_4375,N_589,N_1668);
and U4376 (N_4376,N_1609,N_2355);
and U4377 (N_4377,N_1676,N_2520);
or U4378 (N_4378,N_2871,N_2017);
or U4379 (N_4379,N_2173,N_2899);
nor U4380 (N_4380,N_727,N_1014);
nor U4381 (N_4381,N_216,N_1253);
nand U4382 (N_4382,N_501,N_2301);
nor U4383 (N_4383,N_855,N_251);
nor U4384 (N_4384,N_1245,N_2711);
and U4385 (N_4385,N_163,N_1113);
or U4386 (N_4386,N_1470,N_1234);
or U4387 (N_4387,N_1943,N_2328);
or U4388 (N_4388,N_2370,N_2638);
nor U4389 (N_4389,N_2402,N_1977);
xor U4390 (N_4390,N_1306,N_1122);
and U4391 (N_4391,N_1522,N_2310);
or U4392 (N_4392,N_252,N_206);
or U4393 (N_4393,N_390,N_1836);
nand U4394 (N_4394,N_762,N_1438);
nor U4395 (N_4395,N_1483,N_923);
or U4396 (N_4396,N_397,N_1058);
nand U4397 (N_4397,N_1979,N_1132);
and U4398 (N_4398,N_944,N_1916);
nand U4399 (N_4399,N_2941,N_989);
or U4400 (N_4400,N_474,N_2100);
or U4401 (N_4401,N_1955,N_1054);
or U4402 (N_4402,N_973,N_621);
or U4403 (N_4403,N_1398,N_2046);
nand U4404 (N_4404,N_276,N_558);
xnor U4405 (N_4405,N_2052,N_1617);
nand U4406 (N_4406,N_90,N_2075);
nand U4407 (N_4407,N_1933,N_1608);
or U4408 (N_4408,N_2211,N_1706);
nor U4409 (N_4409,N_329,N_2215);
and U4410 (N_4410,N_2110,N_2216);
or U4411 (N_4411,N_121,N_2148);
xnor U4412 (N_4412,N_11,N_2358);
nor U4413 (N_4413,N_2254,N_160);
and U4414 (N_4414,N_1412,N_1379);
nand U4415 (N_4415,N_1103,N_480);
nand U4416 (N_4416,N_1302,N_2322);
nor U4417 (N_4417,N_96,N_1389);
nor U4418 (N_4418,N_65,N_350);
or U4419 (N_4419,N_1647,N_114);
or U4420 (N_4420,N_1713,N_1232);
nand U4421 (N_4421,N_1501,N_1641);
nor U4422 (N_4422,N_1913,N_1827);
nor U4423 (N_4423,N_250,N_2445);
nor U4424 (N_4424,N_1392,N_303);
and U4425 (N_4425,N_2852,N_2795);
or U4426 (N_4426,N_2755,N_2806);
and U4427 (N_4427,N_260,N_2498);
or U4428 (N_4428,N_984,N_601);
and U4429 (N_4429,N_2588,N_2974);
and U4430 (N_4430,N_1843,N_2030);
or U4431 (N_4431,N_1064,N_1819);
and U4432 (N_4432,N_226,N_1037);
or U4433 (N_4433,N_1723,N_1287);
nand U4434 (N_4434,N_2778,N_1790);
or U4435 (N_4435,N_713,N_628);
nor U4436 (N_4436,N_88,N_2287);
nand U4437 (N_4437,N_1033,N_2284);
or U4438 (N_4438,N_1551,N_2327);
and U4439 (N_4439,N_406,N_540);
xnor U4440 (N_4440,N_162,N_729);
nand U4441 (N_4441,N_2663,N_1405);
or U4442 (N_4442,N_2832,N_828);
and U4443 (N_4443,N_366,N_695);
or U4444 (N_4444,N_165,N_2606);
nand U4445 (N_4445,N_2784,N_314);
xnor U4446 (N_4446,N_2047,N_2129);
nor U4447 (N_4447,N_1994,N_497);
nor U4448 (N_4448,N_1777,N_1057);
and U4449 (N_4449,N_2343,N_608);
or U4450 (N_4450,N_1988,N_1928);
nor U4451 (N_4451,N_179,N_521);
and U4452 (N_4452,N_476,N_439);
and U4453 (N_4453,N_2527,N_2106);
xor U4454 (N_4454,N_2573,N_2954);
or U4455 (N_4455,N_1205,N_1770);
and U4456 (N_4456,N_245,N_2469);
and U4457 (N_4457,N_164,N_1320);
nand U4458 (N_4458,N_2997,N_550);
nand U4459 (N_4459,N_2088,N_1962);
nor U4460 (N_4460,N_2809,N_1434);
and U4461 (N_4461,N_1923,N_1156);
nor U4462 (N_4462,N_2861,N_2669);
nor U4463 (N_4463,N_2395,N_2722);
and U4464 (N_4464,N_1694,N_2232);
nor U4465 (N_4465,N_2213,N_218);
nand U4466 (N_4466,N_1657,N_784);
xor U4467 (N_4467,N_2183,N_2970);
xnor U4468 (N_4468,N_2645,N_1730);
and U4469 (N_4469,N_921,N_454);
or U4470 (N_4470,N_1219,N_17);
nor U4471 (N_4471,N_2699,N_258);
nor U4472 (N_4472,N_1350,N_2837);
xor U4473 (N_4473,N_1651,N_2546);
and U4474 (N_4474,N_438,N_2540);
nor U4475 (N_4475,N_2372,N_1141);
nor U4476 (N_4476,N_657,N_1758);
or U4477 (N_4477,N_586,N_1460);
nor U4478 (N_4478,N_585,N_1428);
nor U4479 (N_4479,N_2063,N_1516);
nand U4480 (N_4480,N_1801,N_854);
nor U4481 (N_4481,N_992,N_1957);
or U4482 (N_4482,N_649,N_612);
nor U4483 (N_4483,N_128,N_2940);
nand U4484 (N_4484,N_1538,N_710);
or U4485 (N_4485,N_2828,N_2330);
nor U4486 (N_4486,N_2814,N_678);
xor U4487 (N_4487,N_1402,N_1426);
or U4488 (N_4488,N_1911,N_587);
nor U4489 (N_4489,N_2170,N_134);
and U4490 (N_4490,N_2862,N_443);
or U4491 (N_4491,N_2608,N_1626);
nor U4492 (N_4492,N_950,N_1939);
and U4493 (N_4493,N_308,N_1093);
and U4494 (N_4494,N_78,N_259);
and U4495 (N_4495,N_1133,N_2574);
or U4496 (N_4496,N_2812,N_2115);
and U4497 (N_4497,N_2056,N_775);
nand U4498 (N_4498,N_1216,N_836);
and U4499 (N_4499,N_770,N_2668);
nand U4500 (N_4500,N_1164,N_209);
nand U4501 (N_4501,N_1245,N_2200);
nor U4502 (N_4502,N_1960,N_515);
and U4503 (N_4503,N_2732,N_1268);
xor U4504 (N_4504,N_492,N_2611);
nor U4505 (N_4505,N_1810,N_1135);
nor U4506 (N_4506,N_2283,N_952);
or U4507 (N_4507,N_1444,N_1317);
nor U4508 (N_4508,N_2998,N_964);
nor U4509 (N_4509,N_869,N_938);
nor U4510 (N_4510,N_782,N_144);
or U4511 (N_4511,N_1554,N_2293);
xor U4512 (N_4512,N_51,N_2813);
or U4513 (N_4513,N_114,N_2537);
nand U4514 (N_4514,N_437,N_1930);
or U4515 (N_4515,N_1638,N_112);
or U4516 (N_4516,N_1651,N_2845);
xnor U4517 (N_4517,N_2843,N_2918);
and U4518 (N_4518,N_2266,N_2213);
and U4519 (N_4519,N_2078,N_837);
or U4520 (N_4520,N_2381,N_820);
and U4521 (N_4521,N_2360,N_1845);
and U4522 (N_4522,N_2021,N_2761);
nor U4523 (N_4523,N_2980,N_2346);
nand U4524 (N_4524,N_1008,N_117);
and U4525 (N_4525,N_1037,N_2725);
nor U4526 (N_4526,N_2874,N_2845);
xnor U4527 (N_4527,N_203,N_1000);
nor U4528 (N_4528,N_60,N_1032);
or U4529 (N_4529,N_173,N_2398);
and U4530 (N_4530,N_2975,N_567);
and U4531 (N_4531,N_576,N_592);
and U4532 (N_4532,N_201,N_1375);
nor U4533 (N_4533,N_2547,N_1300);
and U4534 (N_4534,N_617,N_2456);
nand U4535 (N_4535,N_2703,N_2820);
or U4536 (N_4536,N_825,N_108);
and U4537 (N_4537,N_2472,N_2774);
nand U4538 (N_4538,N_911,N_174);
nand U4539 (N_4539,N_45,N_317);
xor U4540 (N_4540,N_1624,N_2835);
nand U4541 (N_4541,N_1531,N_1634);
nor U4542 (N_4542,N_2273,N_2503);
and U4543 (N_4543,N_586,N_1127);
or U4544 (N_4544,N_2549,N_1907);
and U4545 (N_4545,N_385,N_1443);
and U4546 (N_4546,N_298,N_2718);
nand U4547 (N_4547,N_2853,N_2433);
or U4548 (N_4548,N_2352,N_1730);
and U4549 (N_4549,N_416,N_2641);
nand U4550 (N_4550,N_2104,N_2259);
and U4551 (N_4551,N_2024,N_1594);
nor U4552 (N_4552,N_1793,N_1933);
nand U4553 (N_4553,N_1149,N_1751);
and U4554 (N_4554,N_1506,N_2408);
nor U4555 (N_4555,N_2640,N_672);
or U4556 (N_4556,N_1075,N_2212);
nor U4557 (N_4557,N_507,N_2643);
nand U4558 (N_4558,N_868,N_1876);
and U4559 (N_4559,N_2194,N_2916);
nand U4560 (N_4560,N_1295,N_1223);
and U4561 (N_4561,N_628,N_778);
and U4562 (N_4562,N_453,N_2193);
nand U4563 (N_4563,N_1669,N_1144);
nor U4564 (N_4564,N_44,N_1939);
xor U4565 (N_4565,N_7,N_1386);
xor U4566 (N_4566,N_2256,N_210);
nand U4567 (N_4567,N_2682,N_2165);
and U4568 (N_4568,N_1153,N_276);
or U4569 (N_4569,N_2158,N_2899);
or U4570 (N_4570,N_226,N_1909);
and U4571 (N_4571,N_985,N_1570);
or U4572 (N_4572,N_2634,N_1185);
and U4573 (N_4573,N_543,N_2410);
nor U4574 (N_4574,N_347,N_654);
and U4575 (N_4575,N_221,N_915);
nand U4576 (N_4576,N_1403,N_2892);
and U4577 (N_4577,N_1334,N_961);
xnor U4578 (N_4578,N_2385,N_1439);
nand U4579 (N_4579,N_1102,N_2645);
xor U4580 (N_4580,N_1520,N_124);
or U4581 (N_4581,N_2769,N_1956);
nor U4582 (N_4582,N_389,N_1942);
nand U4583 (N_4583,N_1339,N_2629);
nand U4584 (N_4584,N_320,N_618);
and U4585 (N_4585,N_1356,N_141);
or U4586 (N_4586,N_1418,N_2391);
nand U4587 (N_4587,N_721,N_1463);
or U4588 (N_4588,N_2439,N_1741);
nor U4589 (N_4589,N_614,N_1280);
nor U4590 (N_4590,N_182,N_96);
and U4591 (N_4591,N_1517,N_2049);
or U4592 (N_4592,N_839,N_1453);
nor U4593 (N_4593,N_1246,N_228);
nor U4594 (N_4594,N_2644,N_1059);
nand U4595 (N_4595,N_2512,N_1632);
nor U4596 (N_4596,N_673,N_2862);
and U4597 (N_4597,N_459,N_2271);
nor U4598 (N_4598,N_348,N_2233);
xor U4599 (N_4599,N_2052,N_2863);
or U4600 (N_4600,N_2902,N_62);
or U4601 (N_4601,N_2952,N_562);
nand U4602 (N_4602,N_2352,N_2855);
or U4603 (N_4603,N_182,N_738);
nand U4604 (N_4604,N_707,N_1822);
nor U4605 (N_4605,N_307,N_2089);
or U4606 (N_4606,N_1126,N_2523);
nand U4607 (N_4607,N_778,N_2470);
or U4608 (N_4608,N_1456,N_1007);
or U4609 (N_4609,N_1935,N_1484);
nand U4610 (N_4610,N_2058,N_484);
nand U4611 (N_4611,N_95,N_1480);
xor U4612 (N_4612,N_1669,N_513);
or U4613 (N_4613,N_1708,N_922);
or U4614 (N_4614,N_1398,N_2243);
or U4615 (N_4615,N_1244,N_1622);
or U4616 (N_4616,N_783,N_1548);
xnor U4617 (N_4617,N_1953,N_1355);
xor U4618 (N_4618,N_279,N_326);
nor U4619 (N_4619,N_11,N_2450);
nand U4620 (N_4620,N_2121,N_1275);
or U4621 (N_4621,N_403,N_130);
nor U4622 (N_4622,N_16,N_1344);
or U4623 (N_4623,N_2417,N_2987);
and U4624 (N_4624,N_877,N_203);
nor U4625 (N_4625,N_456,N_2724);
or U4626 (N_4626,N_775,N_402);
nor U4627 (N_4627,N_2578,N_1773);
nand U4628 (N_4628,N_480,N_1409);
and U4629 (N_4629,N_275,N_2201);
nand U4630 (N_4630,N_1892,N_1681);
nand U4631 (N_4631,N_2432,N_2265);
and U4632 (N_4632,N_95,N_1075);
and U4633 (N_4633,N_517,N_1768);
nand U4634 (N_4634,N_164,N_697);
and U4635 (N_4635,N_2220,N_2173);
and U4636 (N_4636,N_2527,N_1039);
xnor U4637 (N_4637,N_2418,N_1546);
and U4638 (N_4638,N_1135,N_709);
xnor U4639 (N_4639,N_259,N_1916);
nand U4640 (N_4640,N_1168,N_1880);
and U4641 (N_4641,N_724,N_881);
nand U4642 (N_4642,N_1828,N_1080);
nor U4643 (N_4643,N_2740,N_1754);
or U4644 (N_4644,N_59,N_2321);
nand U4645 (N_4645,N_1891,N_604);
or U4646 (N_4646,N_147,N_2681);
and U4647 (N_4647,N_2005,N_1315);
or U4648 (N_4648,N_1467,N_236);
or U4649 (N_4649,N_2258,N_2351);
and U4650 (N_4650,N_2512,N_312);
or U4651 (N_4651,N_2662,N_999);
nand U4652 (N_4652,N_2062,N_1892);
nand U4653 (N_4653,N_26,N_2890);
nor U4654 (N_4654,N_1198,N_1441);
nand U4655 (N_4655,N_1811,N_2758);
or U4656 (N_4656,N_2663,N_1964);
and U4657 (N_4657,N_1487,N_1155);
and U4658 (N_4658,N_2647,N_1000);
nand U4659 (N_4659,N_168,N_1141);
or U4660 (N_4660,N_2436,N_1932);
nand U4661 (N_4661,N_1718,N_1855);
xnor U4662 (N_4662,N_2694,N_1965);
nand U4663 (N_4663,N_853,N_1782);
nand U4664 (N_4664,N_1005,N_2289);
xor U4665 (N_4665,N_210,N_1115);
nand U4666 (N_4666,N_900,N_637);
nor U4667 (N_4667,N_669,N_262);
nor U4668 (N_4668,N_2458,N_1851);
and U4669 (N_4669,N_649,N_1318);
and U4670 (N_4670,N_548,N_1493);
xor U4671 (N_4671,N_1506,N_2560);
nor U4672 (N_4672,N_2302,N_1441);
nand U4673 (N_4673,N_2901,N_1816);
and U4674 (N_4674,N_568,N_1894);
nor U4675 (N_4675,N_1230,N_2189);
xor U4676 (N_4676,N_1296,N_1857);
nor U4677 (N_4677,N_1881,N_2467);
or U4678 (N_4678,N_1442,N_517);
xnor U4679 (N_4679,N_2689,N_1138);
or U4680 (N_4680,N_976,N_1503);
or U4681 (N_4681,N_1703,N_733);
and U4682 (N_4682,N_79,N_2822);
and U4683 (N_4683,N_2302,N_489);
nand U4684 (N_4684,N_1317,N_151);
and U4685 (N_4685,N_529,N_2228);
and U4686 (N_4686,N_392,N_980);
and U4687 (N_4687,N_1235,N_309);
and U4688 (N_4688,N_180,N_1281);
nor U4689 (N_4689,N_1616,N_2604);
nand U4690 (N_4690,N_2550,N_1461);
or U4691 (N_4691,N_1179,N_104);
and U4692 (N_4692,N_2100,N_556);
nand U4693 (N_4693,N_2391,N_2906);
and U4694 (N_4694,N_2140,N_2553);
nor U4695 (N_4695,N_2360,N_382);
nand U4696 (N_4696,N_2572,N_97);
xnor U4697 (N_4697,N_1433,N_570);
nor U4698 (N_4698,N_1129,N_907);
and U4699 (N_4699,N_982,N_455);
nand U4700 (N_4700,N_1036,N_187);
nor U4701 (N_4701,N_1246,N_2274);
nor U4702 (N_4702,N_2842,N_2878);
nor U4703 (N_4703,N_2356,N_1549);
nand U4704 (N_4704,N_1894,N_373);
nor U4705 (N_4705,N_2892,N_1553);
nand U4706 (N_4706,N_845,N_269);
nor U4707 (N_4707,N_165,N_1251);
and U4708 (N_4708,N_1214,N_2817);
and U4709 (N_4709,N_347,N_63);
or U4710 (N_4710,N_557,N_92);
xnor U4711 (N_4711,N_362,N_1421);
xnor U4712 (N_4712,N_1301,N_2518);
and U4713 (N_4713,N_830,N_2180);
xnor U4714 (N_4714,N_362,N_480);
xnor U4715 (N_4715,N_635,N_1375);
and U4716 (N_4716,N_1967,N_1385);
nor U4717 (N_4717,N_1137,N_1981);
or U4718 (N_4718,N_85,N_917);
nand U4719 (N_4719,N_1299,N_93);
xnor U4720 (N_4720,N_238,N_1520);
and U4721 (N_4721,N_1419,N_950);
or U4722 (N_4722,N_1002,N_1978);
nor U4723 (N_4723,N_321,N_457);
or U4724 (N_4724,N_989,N_127);
or U4725 (N_4725,N_1110,N_2256);
or U4726 (N_4726,N_1745,N_2819);
and U4727 (N_4727,N_2608,N_2649);
and U4728 (N_4728,N_2255,N_1103);
and U4729 (N_4729,N_805,N_671);
or U4730 (N_4730,N_1215,N_654);
or U4731 (N_4731,N_2895,N_790);
nor U4732 (N_4732,N_2381,N_303);
and U4733 (N_4733,N_1563,N_2416);
nand U4734 (N_4734,N_772,N_2766);
xnor U4735 (N_4735,N_1960,N_882);
and U4736 (N_4736,N_2479,N_214);
and U4737 (N_4737,N_1113,N_1158);
nor U4738 (N_4738,N_1682,N_2927);
or U4739 (N_4739,N_961,N_1040);
and U4740 (N_4740,N_92,N_1905);
and U4741 (N_4741,N_2634,N_2584);
nor U4742 (N_4742,N_2367,N_616);
or U4743 (N_4743,N_2129,N_1844);
nor U4744 (N_4744,N_1039,N_2104);
or U4745 (N_4745,N_150,N_2759);
nand U4746 (N_4746,N_352,N_1757);
nor U4747 (N_4747,N_1648,N_1802);
nand U4748 (N_4748,N_2385,N_2279);
nand U4749 (N_4749,N_889,N_2145);
and U4750 (N_4750,N_921,N_97);
nand U4751 (N_4751,N_1372,N_1514);
nor U4752 (N_4752,N_1405,N_2348);
or U4753 (N_4753,N_1927,N_1338);
or U4754 (N_4754,N_2736,N_2926);
or U4755 (N_4755,N_2851,N_2143);
xor U4756 (N_4756,N_2032,N_2892);
or U4757 (N_4757,N_509,N_2372);
or U4758 (N_4758,N_2988,N_1804);
nor U4759 (N_4759,N_1661,N_1683);
nand U4760 (N_4760,N_1417,N_2415);
or U4761 (N_4761,N_725,N_1651);
nand U4762 (N_4762,N_1370,N_2703);
nand U4763 (N_4763,N_2769,N_2604);
nand U4764 (N_4764,N_2645,N_1441);
or U4765 (N_4765,N_2499,N_2661);
nand U4766 (N_4766,N_960,N_1501);
nor U4767 (N_4767,N_59,N_2608);
and U4768 (N_4768,N_2038,N_349);
or U4769 (N_4769,N_376,N_2596);
or U4770 (N_4770,N_1108,N_1387);
and U4771 (N_4771,N_361,N_1128);
or U4772 (N_4772,N_2735,N_2165);
and U4773 (N_4773,N_691,N_118);
xnor U4774 (N_4774,N_1363,N_2861);
or U4775 (N_4775,N_2345,N_868);
or U4776 (N_4776,N_1341,N_492);
nor U4777 (N_4777,N_2093,N_1577);
and U4778 (N_4778,N_1771,N_2982);
nor U4779 (N_4779,N_2330,N_1024);
xor U4780 (N_4780,N_2653,N_2067);
nor U4781 (N_4781,N_2262,N_2108);
and U4782 (N_4782,N_1738,N_1279);
xor U4783 (N_4783,N_175,N_550);
nor U4784 (N_4784,N_2080,N_1999);
nand U4785 (N_4785,N_2876,N_2596);
nor U4786 (N_4786,N_1928,N_2045);
or U4787 (N_4787,N_2193,N_2757);
or U4788 (N_4788,N_2479,N_1774);
and U4789 (N_4789,N_310,N_1578);
nor U4790 (N_4790,N_2795,N_792);
or U4791 (N_4791,N_1053,N_1952);
and U4792 (N_4792,N_0,N_2181);
nor U4793 (N_4793,N_1288,N_2942);
nand U4794 (N_4794,N_284,N_1324);
nor U4795 (N_4795,N_1778,N_371);
nand U4796 (N_4796,N_1674,N_624);
nor U4797 (N_4797,N_780,N_746);
nor U4798 (N_4798,N_227,N_752);
nor U4799 (N_4799,N_755,N_516);
or U4800 (N_4800,N_693,N_2372);
nor U4801 (N_4801,N_868,N_1923);
and U4802 (N_4802,N_137,N_2904);
or U4803 (N_4803,N_293,N_1456);
and U4804 (N_4804,N_2913,N_756);
or U4805 (N_4805,N_2432,N_1855);
and U4806 (N_4806,N_1341,N_2575);
nand U4807 (N_4807,N_1530,N_458);
and U4808 (N_4808,N_397,N_684);
or U4809 (N_4809,N_320,N_1946);
nor U4810 (N_4810,N_2425,N_2495);
or U4811 (N_4811,N_2240,N_2455);
nor U4812 (N_4812,N_648,N_679);
nor U4813 (N_4813,N_1612,N_158);
nand U4814 (N_4814,N_2254,N_829);
nor U4815 (N_4815,N_2631,N_2968);
or U4816 (N_4816,N_926,N_178);
and U4817 (N_4817,N_2137,N_2151);
nor U4818 (N_4818,N_679,N_2074);
nand U4819 (N_4819,N_447,N_249);
nor U4820 (N_4820,N_1339,N_13);
nor U4821 (N_4821,N_2671,N_190);
or U4822 (N_4822,N_2400,N_2183);
or U4823 (N_4823,N_2640,N_938);
xnor U4824 (N_4824,N_2043,N_2614);
xor U4825 (N_4825,N_511,N_2112);
or U4826 (N_4826,N_1696,N_1527);
or U4827 (N_4827,N_2531,N_903);
nor U4828 (N_4828,N_824,N_127);
nand U4829 (N_4829,N_2186,N_1084);
and U4830 (N_4830,N_2294,N_581);
nor U4831 (N_4831,N_2547,N_2443);
nand U4832 (N_4832,N_232,N_324);
or U4833 (N_4833,N_257,N_2826);
and U4834 (N_4834,N_2853,N_1741);
nand U4835 (N_4835,N_2768,N_2659);
or U4836 (N_4836,N_291,N_2376);
xor U4837 (N_4837,N_232,N_897);
and U4838 (N_4838,N_2294,N_1968);
nor U4839 (N_4839,N_421,N_1448);
nor U4840 (N_4840,N_1983,N_1296);
nand U4841 (N_4841,N_2897,N_335);
nor U4842 (N_4842,N_178,N_2186);
nand U4843 (N_4843,N_1965,N_1458);
or U4844 (N_4844,N_1880,N_2885);
nand U4845 (N_4845,N_556,N_2936);
xnor U4846 (N_4846,N_2749,N_1182);
nor U4847 (N_4847,N_137,N_2993);
nor U4848 (N_4848,N_2805,N_2528);
nand U4849 (N_4849,N_275,N_1843);
nor U4850 (N_4850,N_657,N_195);
and U4851 (N_4851,N_435,N_661);
nor U4852 (N_4852,N_2345,N_1358);
and U4853 (N_4853,N_1821,N_2757);
nor U4854 (N_4854,N_2309,N_1225);
or U4855 (N_4855,N_1426,N_75);
and U4856 (N_4856,N_2674,N_1400);
and U4857 (N_4857,N_1013,N_168);
xor U4858 (N_4858,N_1396,N_755);
nor U4859 (N_4859,N_2030,N_583);
or U4860 (N_4860,N_169,N_467);
nand U4861 (N_4861,N_2573,N_2560);
nand U4862 (N_4862,N_1030,N_1540);
or U4863 (N_4863,N_2452,N_527);
nor U4864 (N_4864,N_584,N_1209);
nor U4865 (N_4865,N_1924,N_885);
nand U4866 (N_4866,N_2697,N_1167);
or U4867 (N_4867,N_2971,N_1411);
nor U4868 (N_4868,N_856,N_926);
nor U4869 (N_4869,N_2287,N_1099);
and U4870 (N_4870,N_2917,N_2675);
nor U4871 (N_4871,N_702,N_2995);
nor U4872 (N_4872,N_912,N_2301);
nand U4873 (N_4873,N_1873,N_2374);
or U4874 (N_4874,N_173,N_2707);
or U4875 (N_4875,N_1882,N_1196);
xnor U4876 (N_4876,N_1802,N_1636);
and U4877 (N_4877,N_2923,N_2007);
or U4878 (N_4878,N_2411,N_2366);
and U4879 (N_4879,N_2734,N_1062);
or U4880 (N_4880,N_2043,N_92);
or U4881 (N_4881,N_2551,N_1766);
nand U4882 (N_4882,N_1782,N_2078);
xor U4883 (N_4883,N_1813,N_1704);
and U4884 (N_4884,N_1556,N_2432);
or U4885 (N_4885,N_1597,N_2914);
nand U4886 (N_4886,N_2489,N_2643);
or U4887 (N_4887,N_2185,N_813);
nor U4888 (N_4888,N_1281,N_1808);
nor U4889 (N_4889,N_58,N_1484);
nand U4890 (N_4890,N_2365,N_850);
and U4891 (N_4891,N_1199,N_2952);
nand U4892 (N_4892,N_987,N_806);
nor U4893 (N_4893,N_1788,N_2136);
and U4894 (N_4894,N_1105,N_646);
xnor U4895 (N_4895,N_1734,N_1393);
or U4896 (N_4896,N_2192,N_1832);
xnor U4897 (N_4897,N_1321,N_2131);
and U4898 (N_4898,N_220,N_843);
nand U4899 (N_4899,N_79,N_2689);
or U4900 (N_4900,N_1291,N_594);
or U4901 (N_4901,N_2882,N_1678);
or U4902 (N_4902,N_2959,N_432);
xnor U4903 (N_4903,N_1397,N_2797);
and U4904 (N_4904,N_32,N_897);
and U4905 (N_4905,N_2024,N_1116);
nand U4906 (N_4906,N_2082,N_2258);
and U4907 (N_4907,N_2183,N_511);
xor U4908 (N_4908,N_2007,N_562);
nor U4909 (N_4909,N_545,N_319);
nand U4910 (N_4910,N_241,N_2408);
nor U4911 (N_4911,N_2633,N_1733);
nor U4912 (N_4912,N_2851,N_2931);
or U4913 (N_4913,N_909,N_2080);
xnor U4914 (N_4914,N_2630,N_1011);
or U4915 (N_4915,N_590,N_2603);
nand U4916 (N_4916,N_1176,N_77);
and U4917 (N_4917,N_2918,N_2473);
and U4918 (N_4918,N_1102,N_515);
nor U4919 (N_4919,N_1540,N_2460);
and U4920 (N_4920,N_1247,N_308);
and U4921 (N_4921,N_1109,N_360);
or U4922 (N_4922,N_480,N_1907);
nor U4923 (N_4923,N_208,N_1961);
nand U4924 (N_4924,N_935,N_109);
xnor U4925 (N_4925,N_1634,N_1152);
nor U4926 (N_4926,N_2536,N_1738);
or U4927 (N_4927,N_2627,N_1840);
nand U4928 (N_4928,N_384,N_2018);
and U4929 (N_4929,N_1213,N_1708);
and U4930 (N_4930,N_637,N_2888);
xor U4931 (N_4931,N_203,N_926);
nor U4932 (N_4932,N_1610,N_897);
and U4933 (N_4933,N_1407,N_640);
nor U4934 (N_4934,N_2425,N_2050);
nand U4935 (N_4935,N_2196,N_113);
nor U4936 (N_4936,N_589,N_2874);
nor U4937 (N_4937,N_1956,N_2636);
or U4938 (N_4938,N_2082,N_2127);
and U4939 (N_4939,N_1615,N_1543);
nor U4940 (N_4940,N_2032,N_1413);
xor U4941 (N_4941,N_648,N_2628);
or U4942 (N_4942,N_2969,N_1175);
nand U4943 (N_4943,N_66,N_438);
nor U4944 (N_4944,N_1893,N_1224);
or U4945 (N_4945,N_425,N_2124);
or U4946 (N_4946,N_451,N_542);
or U4947 (N_4947,N_652,N_77);
nand U4948 (N_4948,N_699,N_2892);
nand U4949 (N_4949,N_502,N_30);
xnor U4950 (N_4950,N_1621,N_684);
and U4951 (N_4951,N_1005,N_75);
nor U4952 (N_4952,N_1209,N_1308);
nor U4953 (N_4953,N_2264,N_912);
nand U4954 (N_4954,N_2329,N_1386);
nor U4955 (N_4955,N_1822,N_100);
nor U4956 (N_4956,N_983,N_1001);
nor U4957 (N_4957,N_416,N_2133);
nor U4958 (N_4958,N_1355,N_1168);
and U4959 (N_4959,N_631,N_825);
or U4960 (N_4960,N_1091,N_663);
or U4961 (N_4961,N_2307,N_1637);
and U4962 (N_4962,N_382,N_670);
or U4963 (N_4963,N_1206,N_2423);
or U4964 (N_4964,N_2143,N_2448);
nor U4965 (N_4965,N_2317,N_943);
or U4966 (N_4966,N_348,N_2223);
or U4967 (N_4967,N_2312,N_803);
and U4968 (N_4968,N_1464,N_547);
nand U4969 (N_4969,N_1152,N_2646);
nand U4970 (N_4970,N_379,N_939);
nor U4971 (N_4971,N_1028,N_1927);
nor U4972 (N_4972,N_517,N_996);
or U4973 (N_4973,N_1539,N_1146);
xor U4974 (N_4974,N_1070,N_2485);
or U4975 (N_4975,N_707,N_2933);
nor U4976 (N_4976,N_85,N_2649);
nor U4977 (N_4977,N_1940,N_1138);
and U4978 (N_4978,N_1384,N_1173);
and U4979 (N_4979,N_614,N_1519);
or U4980 (N_4980,N_2504,N_1101);
or U4981 (N_4981,N_226,N_1669);
and U4982 (N_4982,N_2979,N_42);
nor U4983 (N_4983,N_356,N_631);
xor U4984 (N_4984,N_511,N_2951);
and U4985 (N_4985,N_333,N_2009);
or U4986 (N_4986,N_2673,N_1907);
xor U4987 (N_4987,N_1343,N_2946);
nand U4988 (N_4988,N_2106,N_1186);
xor U4989 (N_4989,N_22,N_835);
nor U4990 (N_4990,N_2303,N_206);
and U4991 (N_4991,N_250,N_1546);
or U4992 (N_4992,N_79,N_1503);
nand U4993 (N_4993,N_992,N_943);
nand U4994 (N_4994,N_2784,N_491);
nor U4995 (N_4995,N_69,N_1798);
nand U4996 (N_4996,N_1861,N_663);
and U4997 (N_4997,N_1856,N_2470);
nor U4998 (N_4998,N_1286,N_2247);
nand U4999 (N_4999,N_2920,N_1282);
nand U5000 (N_5000,N_151,N_1098);
nor U5001 (N_5001,N_2226,N_1785);
nand U5002 (N_5002,N_1441,N_1508);
or U5003 (N_5003,N_1091,N_91);
nor U5004 (N_5004,N_2597,N_1206);
or U5005 (N_5005,N_1292,N_801);
nand U5006 (N_5006,N_1894,N_537);
or U5007 (N_5007,N_863,N_2585);
nor U5008 (N_5008,N_287,N_290);
or U5009 (N_5009,N_1488,N_2441);
xor U5010 (N_5010,N_341,N_2963);
or U5011 (N_5011,N_185,N_2404);
or U5012 (N_5012,N_1936,N_1483);
and U5013 (N_5013,N_333,N_1711);
and U5014 (N_5014,N_2063,N_2525);
and U5015 (N_5015,N_1017,N_2780);
and U5016 (N_5016,N_752,N_719);
or U5017 (N_5017,N_905,N_123);
xnor U5018 (N_5018,N_365,N_2974);
or U5019 (N_5019,N_992,N_1747);
nand U5020 (N_5020,N_1870,N_1790);
xnor U5021 (N_5021,N_1832,N_620);
and U5022 (N_5022,N_748,N_1254);
nand U5023 (N_5023,N_2258,N_2992);
nor U5024 (N_5024,N_2303,N_1776);
and U5025 (N_5025,N_821,N_946);
and U5026 (N_5026,N_1196,N_167);
nor U5027 (N_5027,N_297,N_2936);
nand U5028 (N_5028,N_2598,N_2339);
nor U5029 (N_5029,N_108,N_1701);
nand U5030 (N_5030,N_869,N_2206);
nor U5031 (N_5031,N_1551,N_617);
xnor U5032 (N_5032,N_548,N_2656);
nand U5033 (N_5033,N_2696,N_2857);
nand U5034 (N_5034,N_529,N_812);
nand U5035 (N_5035,N_1387,N_2340);
or U5036 (N_5036,N_2626,N_293);
nor U5037 (N_5037,N_379,N_2463);
or U5038 (N_5038,N_1437,N_1294);
or U5039 (N_5039,N_1516,N_1631);
nor U5040 (N_5040,N_976,N_2058);
and U5041 (N_5041,N_2502,N_1255);
nor U5042 (N_5042,N_1719,N_610);
nand U5043 (N_5043,N_1472,N_1604);
nand U5044 (N_5044,N_2642,N_991);
nor U5045 (N_5045,N_1150,N_832);
and U5046 (N_5046,N_1467,N_447);
nor U5047 (N_5047,N_1392,N_69);
nor U5048 (N_5048,N_2638,N_2527);
nand U5049 (N_5049,N_1462,N_1070);
or U5050 (N_5050,N_1816,N_2101);
nand U5051 (N_5051,N_2001,N_1260);
nand U5052 (N_5052,N_2811,N_2526);
nor U5053 (N_5053,N_165,N_520);
nor U5054 (N_5054,N_2156,N_2382);
nor U5055 (N_5055,N_2711,N_1034);
nand U5056 (N_5056,N_2695,N_2797);
or U5057 (N_5057,N_725,N_742);
or U5058 (N_5058,N_652,N_2048);
nand U5059 (N_5059,N_2886,N_1634);
nor U5060 (N_5060,N_1768,N_427);
and U5061 (N_5061,N_761,N_706);
or U5062 (N_5062,N_199,N_2451);
or U5063 (N_5063,N_1541,N_976);
or U5064 (N_5064,N_2014,N_1833);
or U5065 (N_5065,N_478,N_185);
or U5066 (N_5066,N_1012,N_1423);
and U5067 (N_5067,N_24,N_311);
nand U5068 (N_5068,N_101,N_516);
or U5069 (N_5069,N_1063,N_136);
and U5070 (N_5070,N_2082,N_602);
and U5071 (N_5071,N_696,N_1709);
nor U5072 (N_5072,N_52,N_2953);
or U5073 (N_5073,N_1256,N_1243);
nor U5074 (N_5074,N_1229,N_1767);
and U5075 (N_5075,N_2451,N_1379);
or U5076 (N_5076,N_2235,N_118);
and U5077 (N_5077,N_2294,N_1179);
nor U5078 (N_5078,N_67,N_318);
nor U5079 (N_5079,N_702,N_2172);
nor U5080 (N_5080,N_961,N_862);
nor U5081 (N_5081,N_1337,N_2712);
and U5082 (N_5082,N_2510,N_2057);
nand U5083 (N_5083,N_2306,N_64);
xnor U5084 (N_5084,N_279,N_2825);
and U5085 (N_5085,N_443,N_2882);
or U5086 (N_5086,N_2978,N_2240);
xor U5087 (N_5087,N_1919,N_1224);
nand U5088 (N_5088,N_1574,N_1305);
nor U5089 (N_5089,N_1929,N_1367);
and U5090 (N_5090,N_2058,N_526);
nor U5091 (N_5091,N_2836,N_2402);
or U5092 (N_5092,N_1761,N_1866);
xnor U5093 (N_5093,N_2049,N_577);
nor U5094 (N_5094,N_1021,N_1474);
xnor U5095 (N_5095,N_2994,N_1674);
and U5096 (N_5096,N_1620,N_1117);
nand U5097 (N_5097,N_664,N_2730);
xnor U5098 (N_5098,N_1873,N_2676);
and U5099 (N_5099,N_1925,N_2509);
nor U5100 (N_5100,N_1515,N_1090);
nand U5101 (N_5101,N_2226,N_921);
nand U5102 (N_5102,N_2607,N_2168);
nor U5103 (N_5103,N_2858,N_35);
nor U5104 (N_5104,N_1389,N_624);
nor U5105 (N_5105,N_2557,N_141);
nand U5106 (N_5106,N_1006,N_1468);
and U5107 (N_5107,N_266,N_514);
nor U5108 (N_5108,N_861,N_1365);
or U5109 (N_5109,N_167,N_1083);
nor U5110 (N_5110,N_1706,N_2270);
nor U5111 (N_5111,N_1441,N_1303);
nand U5112 (N_5112,N_2262,N_2560);
nand U5113 (N_5113,N_2662,N_2851);
or U5114 (N_5114,N_563,N_2471);
nor U5115 (N_5115,N_1292,N_1205);
or U5116 (N_5116,N_82,N_2098);
nor U5117 (N_5117,N_1440,N_2289);
nand U5118 (N_5118,N_153,N_1983);
or U5119 (N_5119,N_2351,N_2309);
or U5120 (N_5120,N_1155,N_1491);
nor U5121 (N_5121,N_2550,N_1973);
xor U5122 (N_5122,N_60,N_1064);
nor U5123 (N_5123,N_1221,N_2515);
xor U5124 (N_5124,N_1468,N_2488);
and U5125 (N_5125,N_1113,N_2677);
and U5126 (N_5126,N_2101,N_2662);
nor U5127 (N_5127,N_485,N_2184);
nor U5128 (N_5128,N_1181,N_476);
and U5129 (N_5129,N_1768,N_1565);
and U5130 (N_5130,N_1774,N_1165);
and U5131 (N_5131,N_2138,N_1965);
nor U5132 (N_5132,N_1621,N_1260);
xnor U5133 (N_5133,N_1702,N_2133);
nand U5134 (N_5134,N_2312,N_478);
and U5135 (N_5135,N_1504,N_2286);
and U5136 (N_5136,N_2488,N_1944);
nand U5137 (N_5137,N_1382,N_2498);
nand U5138 (N_5138,N_2813,N_455);
or U5139 (N_5139,N_866,N_2621);
nor U5140 (N_5140,N_2472,N_1865);
and U5141 (N_5141,N_866,N_1738);
nor U5142 (N_5142,N_259,N_2419);
xnor U5143 (N_5143,N_2000,N_2315);
nor U5144 (N_5144,N_133,N_788);
and U5145 (N_5145,N_1090,N_865);
nor U5146 (N_5146,N_970,N_2139);
nand U5147 (N_5147,N_1948,N_2488);
or U5148 (N_5148,N_2388,N_2749);
nor U5149 (N_5149,N_332,N_2201);
nor U5150 (N_5150,N_770,N_433);
nand U5151 (N_5151,N_742,N_789);
or U5152 (N_5152,N_60,N_1620);
or U5153 (N_5153,N_1521,N_1559);
and U5154 (N_5154,N_1849,N_1185);
xor U5155 (N_5155,N_583,N_1720);
nand U5156 (N_5156,N_603,N_550);
nor U5157 (N_5157,N_1832,N_286);
or U5158 (N_5158,N_2800,N_369);
and U5159 (N_5159,N_175,N_835);
nand U5160 (N_5160,N_1080,N_29);
or U5161 (N_5161,N_2346,N_675);
xor U5162 (N_5162,N_142,N_29);
nand U5163 (N_5163,N_1873,N_1680);
and U5164 (N_5164,N_2932,N_613);
and U5165 (N_5165,N_16,N_2451);
nor U5166 (N_5166,N_1661,N_2092);
and U5167 (N_5167,N_756,N_1114);
nor U5168 (N_5168,N_763,N_1569);
or U5169 (N_5169,N_901,N_754);
or U5170 (N_5170,N_1624,N_945);
nand U5171 (N_5171,N_230,N_2599);
xnor U5172 (N_5172,N_2093,N_1071);
nor U5173 (N_5173,N_2956,N_1248);
or U5174 (N_5174,N_760,N_1525);
and U5175 (N_5175,N_2706,N_1666);
nand U5176 (N_5176,N_2752,N_84);
nor U5177 (N_5177,N_1151,N_2062);
nand U5178 (N_5178,N_2240,N_330);
nand U5179 (N_5179,N_2642,N_2898);
nand U5180 (N_5180,N_1290,N_426);
nand U5181 (N_5181,N_2084,N_2352);
and U5182 (N_5182,N_2148,N_245);
and U5183 (N_5183,N_1073,N_79);
nor U5184 (N_5184,N_946,N_1601);
or U5185 (N_5185,N_1850,N_487);
nor U5186 (N_5186,N_2227,N_199);
and U5187 (N_5187,N_1450,N_1668);
nor U5188 (N_5188,N_665,N_2835);
nand U5189 (N_5189,N_1160,N_1761);
nand U5190 (N_5190,N_1351,N_2268);
or U5191 (N_5191,N_763,N_170);
and U5192 (N_5192,N_2639,N_2000);
nand U5193 (N_5193,N_451,N_2600);
or U5194 (N_5194,N_2436,N_2181);
or U5195 (N_5195,N_2517,N_2467);
nand U5196 (N_5196,N_1592,N_2805);
and U5197 (N_5197,N_2287,N_1353);
or U5198 (N_5198,N_967,N_1839);
nor U5199 (N_5199,N_2171,N_954);
nand U5200 (N_5200,N_35,N_642);
and U5201 (N_5201,N_2331,N_551);
and U5202 (N_5202,N_2945,N_1260);
nor U5203 (N_5203,N_118,N_693);
nand U5204 (N_5204,N_979,N_1042);
nand U5205 (N_5205,N_2892,N_2116);
nand U5206 (N_5206,N_498,N_2361);
and U5207 (N_5207,N_1940,N_2441);
or U5208 (N_5208,N_1334,N_1948);
nor U5209 (N_5209,N_2730,N_15);
and U5210 (N_5210,N_2250,N_212);
xnor U5211 (N_5211,N_921,N_1112);
or U5212 (N_5212,N_2348,N_2179);
and U5213 (N_5213,N_376,N_2916);
nor U5214 (N_5214,N_1981,N_1603);
nand U5215 (N_5215,N_1971,N_98);
and U5216 (N_5216,N_23,N_363);
nor U5217 (N_5217,N_2245,N_2190);
or U5218 (N_5218,N_2509,N_1388);
nand U5219 (N_5219,N_126,N_1937);
or U5220 (N_5220,N_1082,N_2273);
or U5221 (N_5221,N_1177,N_2660);
nand U5222 (N_5222,N_1312,N_2129);
nor U5223 (N_5223,N_1482,N_1712);
nor U5224 (N_5224,N_2022,N_118);
nor U5225 (N_5225,N_1721,N_1860);
nand U5226 (N_5226,N_2957,N_2062);
or U5227 (N_5227,N_2904,N_1516);
nor U5228 (N_5228,N_2450,N_385);
nand U5229 (N_5229,N_2274,N_2603);
or U5230 (N_5230,N_2525,N_197);
nor U5231 (N_5231,N_599,N_2471);
nand U5232 (N_5232,N_876,N_1083);
nor U5233 (N_5233,N_1647,N_472);
and U5234 (N_5234,N_2464,N_95);
nor U5235 (N_5235,N_1451,N_2960);
and U5236 (N_5236,N_2137,N_331);
nor U5237 (N_5237,N_1242,N_2629);
or U5238 (N_5238,N_1136,N_1281);
or U5239 (N_5239,N_1193,N_1737);
nor U5240 (N_5240,N_2056,N_224);
nand U5241 (N_5241,N_1170,N_597);
nor U5242 (N_5242,N_118,N_2584);
nor U5243 (N_5243,N_1731,N_2189);
nand U5244 (N_5244,N_138,N_2834);
xor U5245 (N_5245,N_2634,N_491);
or U5246 (N_5246,N_1440,N_2255);
nor U5247 (N_5247,N_2200,N_2698);
nand U5248 (N_5248,N_1465,N_1797);
and U5249 (N_5249,N_979,N_2291);
and U5250 (N_5250,N_2480,N_2988);
nor U5251 (N_5251,N_2507,N_1582);
or U5252 (N_5252,N_203,N_816);
nor U5253 (N_5253,N_2106,N_872);
nand U5254 (N_5254,N_2737,N_2149);
or U5255 (N_5255,N_1402,N_995);
or U5256 (N_5256,N_2395,N_2758);
nor U5257 (N_5257,N_986,N_2073);
nor U5258 (N_5258,N_1486,N_1762);
nand U5259 (N_5259,N_2227,N_481);
or U5260 (N_5260,N_1661,N_690);
xor U5261 (N_5261,N_2206,N_1100);
nand U5262 (N_5262,N_2205,N_1513);
nand U5263 (N_5263,N_1364,N_1315);
or U5264 (N_5264,N_1810,N_1218);
or U5265 (N_5265,N_2000,N_860);
and U5266 (N_5266,N_2052,N_799);
and U5267 (N_5267,N_110,N_46);
and U5268 (N_5268,N_302,N_2033);
nand U5269 (N_5269,N_752,N_2414);
or U5270 (N_5270,N_2670,N_93);
xnor U5271 (N_5271,N_154,N_2891);
and U5272 (N_5272,N_1606,N_426);
nand U5273 (N_5273,N_634,N_1610);
and U5274 (N_5274,N_1342,N_2178);
nor U5275 (N_5275,N_94,N_705);
nand U5276 (N_5276,N_2459,N_875);
and U5277 (N_5277,N_1537,N_1973);
nand U5278 (N_5278,N_801,N_2059);
nand U5279 (N_5279,N_1766,N_835);
or U5280 (N_5280,N_768,N_379);
xnor U5281 (N_5281,N_747,N_2025);
and U5282 (N_5282,N_2783,N_1209);
or U5283 (N_5283,N_281,N_2430);
and U5284 (N_5284,N_131,N_2596);
nor U5285 (N_5285,N_2676,N_1676);
or U5286 (N_5286,N_2968,N_1693);
nor U5287 (N_5287,N_2471,N_2681);
or U5288 (N_5288,N_2393,N_749);
or U5289 (N_5289,N_1831,N_948);
and U5290 (N_5290,N_2743,N_1642);
nand U5291 (N_5291,N_2888,N_49);
and U5292 (N_5292,N_474,N_2921);
nand U5293 (N_5293,N_2929,N_134);
and U5294 (N_5294,N_1099,N_2480);
nor U5295 (N_5295,N_860,N_1582);
nand U5296 (N_5296,N_1318,N_728);
and U5297 (N_5297,N_2495,N_706);
xnor U5298 (N_5298,N_68,N_648);
xor U5299 (N_5299,N_1507,N_696);
and U5300 (N_5300,N_2245,N_237);
nand U5301 (N_5301,N_2622,N_43);
nor U5302 (N_5302,N_1615,N_2539);
nor U5303 (N_5303,N_440,N_121);
nor U5304 (N_5304,N_873,N_503);
nor U5305 (N_5305,N_508,N_1290);
nor U5306 (N_5306,N_2940,N_70);
xor U5307 (N_5307,N_1402,N_2321);
nor U5308 (N_5308,N_2068,N_908);
or U5309 (N_5309,N_881,N_1265);
nor U5310 (N_5310,N_1287,N_2330);
nor U5311 (N_5311,N_1407,N_723);
or U5312 (N_5312,N_1929,N_124);
and U5313 (N_5313,N_1714,N_2900);
or U5314 (N_5314,N_1575,N_284);
nand U5315 (N_5315,N_187,N_795);
or U5316 (N_5316,N_1728,N_2795);
or U5317 (N_5317,N_2958,N_686);
nor U5318 (N_5318,N_2986,N_1894);
nand U5319 (N_5319,N_2066,N_2650);
xnor U5320 (N_5320,N_2671,N_1506);
nor U5321 (N_5321,N_1133,N_123);
or U5322 (N_5322,N_2780,N_2010);
and U5323 (N_5323,N_366,N_1370);
or U5324 (N_5324,N_2273,N_1490);
nor U5325 (N_5325,N_2649,N_1793);
nor U5326 (N_5326,N_1532,N_2007);
or U5327 (N_5327,N_1561,N_1543);
nor U5328 (N_5328,N_2049,N_610);
and U5329 (N_5329,N_1241,N_2091);
or U5330 (N_5330,N_2384,N_1534);
or U5331 (N_5331,N_1925,N_1477);
xor U5332 (N_5332,N_854,N_2998);
nor U5333 (N_5333,N_1603,N_1997);
xnor U5334 (N_5334,N_1402,N_1844);
or U5335 (N_5335,N_2842,N_2222);
nand U5336 (N_5336,N_2527,N_141);
or U5337 (N_5337,N_1053,N_2674);
and U5338 (N_5338,N_1890,N_2299);
xor U5339 (N_5339,N_1197,N_1209);
and U5340 (N_5340,N_293,N_2462);
and U5341 (N_5341,N_134,N_1919);
nand U5342 (N_5342,N_1401,N_1716);
nor U5343 (N_5343,N_2974,N_1754);
nor U5344 (N_5344,N_2208,N_49);
nor U5345 (N_5345,N_753,N_2273);
and U5346 (N_5346,N_1728,N_1502);
nand U5347 (N_5347,N_209,N_322);
or U5348 (N_5348,N_2315,N_2783);
nor U5349 (N_5349,N_583,N_458);
or U5350 (N_5350,N_2685,N_2868);
or U5351 (N_5351,N_552,N_2286);
or U5352 (N_5352,N_2931,N_2252);
or U5353 (N_5353,N_2739,N_2497);
nand U5354 (N_5354,N_1776,N_1966);
or U5355 (N_5355,N_1774,N_2247);
nor U5356 (N_5356,N_1580,N_724);
or U5357 (N_5357,N_2919,N_2815);
or U5358 (N_5358,N_535,N_741);
nor U5359 (N_5359,N_2243,N_2576);
or U5360 (N_5360,N_2082,N_401);
and U5361 (N_5361,N_1528,N_628);
or U5362 (N_5362,N_2742,N_1924);
nand U5363 (N_5363,N_2042,N_2398);
or U5364 (N_5364,N_1413,N_838);
and U5365 (N_5365,N_783,N_1882);
nand U5366 (N_5366,N_1439,N_1281);
xnor U5367 (N_5367,N_954,N_239);
and U5368 (N_5368,N_447,N_779);
or U5369 (N_5369,N_1829,N_323);
and U5370 (N_5370,N_1863,N_716);
or U5371 (N_5371,N_1009,N_2610);
and U5372 (N_5372,N_161,N_2887);
nor U5373 (N_5373,N_370,N_1790);
nor U5374 (N_5374,N_830,N_1060);
or U5375 (N_5375,N_1065,N_2440);
nor U5376 (N_5376,N_1730,N_927);
and U5377 (N_5377,N_1112,N_1932);
and U5378 (N_5378,N_1577,N_743);
or U5379 (N_5379,N_1496,N_1522);
and U5380 (N_5380,N_1473,N_1479);
nand U5381 (N_5381,N_1430,N_2400);
nor U5382 (N_5382,N_961,N_877);
xnor U5383 (N_5383,N_2982,N_2706);
or U5384 (N_5384,N_783,N_1428);
and U5385 (N_5385,N_1026,N_802);
nor U5386 (N_5386,N_2137,N_1264);
and U5387 (N_5387,N_1764,N_2002);
xor U5388 (N_5388,N_1373,N_103);
nor U5389 (N_5389,N_1982,N_248);
or U5390 (N_5390,N_515,N_2068);
or U5391 (N_5391,N_1048,N_836);
and U5392 (N_5392,N_1201,N_865);
and U5393 (N_5393,N_529,N_766);
nor U5394 (N_5394,N_41,N_1870);
and U5395 (N_5395,N_2782,N_2908);
nor U5396 (N_5396,N_352,N_1663);
or U5397 (N_5397,N_2314,N_2033);
or U5398 (N_5398,N_1886,N_683);
and U5399 (N_5399,N_2019,N_589);
or U5400 (N_5400,N_742,N_2399);
and U5401 (N_5401,N_2652,N_1823);
nor U5402 (N_5402,N_2962,N_1535);
and U5403 (N_5403,N_1593,N_1723);
nand U5404 (N_5404,N_1211,N_1809);
and U5405 (N_5405,N_628,N_675);
and U5406 (N_5406,N_795,N_1980);
and U5407 (N_5407,N_1000,N_2396);
or U5408 (N_5408,N_2506,N_2429);
nor U5409 (N_5409,N_2768,N_1265);
nor U5410 (N_5410,N_20,N_2761);
nand U5411 (N_5411,N_105,N_2785);
or U5412 (N_5412,N_1767,N_1601);
xnor U5413 (N_5413,N_1683,N_2290);
nor U5414 (N_5414,N_1336,N_2412);
nor U5415 (N_5415,N_886,N_1946);
nor U5416 (N_5416,N_1280,N_272);
nor U5417 (N_5417,N_1390,N_18);
and U5418 (N_5418,N_941,N_1003);
or U5419 (N_5419,N_2006,N_2712);
and U5420 (N_5420,N_2891,N_1711);
or U5421 (N_5421,N_2111,N_1176);
nand U5422 (N_5422,N_281,N_111);
or U5423 (N_5423,N_1693,N_2595);
or U5424 (N_5424,N_858,N_908);
xor U5425 (N_5425,N_2390,N_2272);
nand U5426 (N_5426,N_2517,N_2402);
nor U5427 (N_5427,N_28,N_1195);
or U5428 (N_5428,N_2601,N_2885);
or U5429 (N_5429,N_2928,N_1854);
nor U5430 (N_5430,N_2751,N_2927);
and U5431 (N_5431,N_2469,N_1329);
or U5432 (N_5432,N_1203,N_2177);
nor U5433 (N_5433,N_1562,N_260);
xor U5434 (N_5434,N_943,N_1551);
nand U5435 (N_5435,N_1042,N_1360);
xor U5436 (N_5436,N_206,N_191);
nor U5437 (N_5437,N_1939,N_478);
or U5438 (N_5438,N_2583,N_1338);
nor U5439 (N_5439,N_1131,N_1314);
and U5440 (N_5440,N_2351,N_2172);
nor U5441 (N_5441,N_2168,N_2041);
and U5442 (N_5442,N_1066,N_704);
nand U5443 (N_5443,N_2036,N_2819);
and U5444 (N_5444,N_361,N_2408);
nand U5445 (N_5445,N_2400,N_2035);
or U5446 (N_5446,N_51,N_1747);
or U5447 (N_5447,N_2259,N_1102);
and U5448 (N_5448,N_1663,N_2565);
nand U5449 (N_5449,N_877,N_2240);
nand U5450 (N_5450,N_1765,N_520);
and U5451 (N_5451,N_737,N_939);
xnor U5452 (N_5452,N_2054,N_1415);
and U5453 (N_5453,N_2528,N_2271);
nand U5454 (N_5454,N_2053,N_647);
and U5455 (N_5455,N_1661,N_2294);
nand U5456 (N_5456,N_37,N_1490);
and U5457 (N_5457,N_1173,N_2217);
nand U5458 (N_5458,N_1542,N_206);
or U5459 (N_5459,N_903,N_529);
and U5460 (N_5460,N_797,N_2939);
nand U5461 (N_5461,N_2111,N_1796);
nand U5462 (N_5462,N_984,N_840);
and U5463 (N_5463,N_744,N_758);
xor U5464 (N_5464,N_181,N_257);
and U5465 (N_5465,N_1487,N_657);
nand U5466 (N_5466,N_2282,N_1042);
or U5467 (N_5467,N_1305,N_1645);
nor U5468 (N_5468,N_1972,N_2398);
nand U5469 (N_5469,N_766,N_540);
and U5470 (N_5470,N_433,N_391);
or U5471 (N_5471,N_1048,N_552);
nand U5472 (N_5472,N_2259,N_232);
or U5473 (N_5473,N_926,N_200);
and U5474 (N_5474,N_692,N_608);
xor U5475 (N_5475,N_713,N_2224);
or U5476 (N_5476,N_2612,N_607);
and U5477 (N_5477,N_2234,N_1203);
xor U5478 (N_5478,N_1828,N_2866);
and U5479 (N_5479,N_481,N_644);
xnor U5480 (N_5480,N_1608,N_2757);
and U5481 (N_5481,N_1245,N_2737);
or U5482 (N_5482,N_930,N_262);
and U5483 (N_5483,N_2868,N_1862);
and U5484 (N_5484,N_2022,N_2263);
and U5485 (N_5485,N_205,N_2709);
nand U5486 (N_5486,N_1616,N_2704);
nor U5487 (N_5487,N_1239,N_1305);
nor U5488 (N_5488,N_2476,N_1680);
or U5489 (N_5489,N_2821,N_1376);
and U5490 (N_5490,N_1607,N_1221);
nor U5491 (N_5491,N_2036,N_1478);
nor U5492 (N_5492,N_513,N_2468);
and U5493 (N_5493,N_1876,N_965);
and U5494 (N_5494,N_771,N_2608);
xor U5495 (N_5495,N_644,N_192);
and U5496 (N_5496,N_2684,N_2609);
or U5497 (N_5497,N_2291,N_40);
or U5498 (N_5498,N_1388,N_2716);
nand U5499 (N_5499,N_1404,N_684);
and U5500 (N_5500,N_2976,N_1654);
xnor U5501 (N_5501,N_2432,N_1266);
nor U5502 (N_5502,N_1834,N_484);
xnor U5503 (N_5503,N_66,N_255);
or U5504 (N_5504,N_1340,N_472);
and U5505 (N_5505,N_1816,N_1616);
or U5506 (N_5506,N_962,N_2728);
or U5507 (N_5507,N_2231,N_1449);
xor U5508 (N_5508,N_2657,N_1340);
nor U5509 (N_5509,N_98,N_1012);
and U5510 (N_5510,N_2412,N_2383);
xor U5511 (N_5511,N_1041,N_1729);
nor U5512 (N_5512,N_800,N_701);
nand U5513 (N_5513,N_2277,N_2066);
nand U5514 (N_5514,N_770,N_721);
nand U5515 (N_5515,N_648,N_2229);
and U5516 (N_5516,N_1905,N_2198);
and U5517 (N_5517,N_934,N_768);
nand U5518 (N_5518,N_952,N_1929);
and U5519 (N_5519,N_531,N_2145);
and U5520 (N_5520,N_64,N_2551);
or U5521 (N_5521,N_1457,N_2732);
or U5522 (N_5522,N_1928,N_394);
nor U5523 (N_5523,N_2847,N_794);
or U5524 (N_5524,N_417,N_2452);
or U5525 (N_5525,N_785,N_1659);
nand U5526 (N_5526,N_1332,N_2913);
or U5527 (N_5527,N_2737,N_685);
and U5528 (N_5528,N_90,N_2980);
xnor U5529 (N_5529,N_1576,N_1040);
and U5530 (N_5530,N_214,N_334);
nand U5531 (N_5531,N_1714,N_78);
and U5532 (N_5532,N_1689,N_2270);
nand U5533 (N_5533,N_385,N_2812);
nand U5534 (N_5534,N_717,N_907);
and U5535 (N_5535,N_1518,N_2350);
or U5536 (N_5536,N_295,N_2428);
nand U5537 (N_5537,N_2558,N_2690);
nand U5538 (N_5538,N_1117,N_2486);
nor U5539 (N_5539,N_1320,N_1110);
or U5540 (N_5540,N_1051,N_777);
xnor U5541 (N_5541,N_2455,N_168);
nand U5542 (N_5542,N_1068,N_673);
nand U5543 (N_5543,N_240,N_2698);
and U5544 (N_5544,N_623,N_1512);
nand U5545 (N_5545,N_717,N_2584);
nand U5546 (N_5546,N_625,N_2629);
and U5547 (N_5547,N_23,N_1558);
or U5548 (N_5548,N_706,N_1840);
and U5549 (N_5549,N_1760,N_2726);
nor U5550 (N_5550,N_1844,N_2201);
nor U5551 (N_5551,N_997,N_2749);
nor U5552 (N_5552,N_543,N_2869);
nor U5553 (N_5553,N_675,N_1678);
and U5554 (N_5554,N_2484,N_945);
or U5555 (N_5555,N_1846,N_2526);
and U5556 (N_5556,N_573,N_1558);
nor U5557 (N_5557,N_1684,N_114);
or U5558 (N_5558,N_1453,N_192);
xnor U5559 (N_5559,N_1242,N_2258);
or U5560 (N_5560,N_2177,N_2003);
or U5561 (N_5561,N_49,N_1634);
nor U5562 (N_5562,N_899,N_737);
or U5563 (N_5563,N_220,N_1883);
nand U5564 (N_5564,N_1375,N_1995);
xor U5565 (N_5565,N_2991,N_647);
nand U5566 (N_5566,N_1620,N_2184);
nand U5567 (N_5567,N_1120,N_2055);
and U5568 (N_5568,N_269,N_1468);
or U5569 (N_5569,N_385,N_1270);
nand U5570 (N_5570,N_902,N_579);
or U5571 (N_5571,N_85,N_930);
nand U5572 (N_5572,N_647,N_1161);
or U5573 (N_5573,N_1741,N_1333);
nand U5574 (N_5574,N_199,N_1340);
nor U5575 (N_5575,N_354,N_683);
nor U5576 (N_5576,N_2143,N_940);
or U5577 (N_5577,N_283,N_2716);
and U5578 (N_5578,N_2056,N_648);
nor U5579 (N_5579,N_1917,N_2048);
nor U5580 (N_5580,N_665,N_505);
nand U5581 (N_5581,N_1050,N_2490);
and U5582 (N_5582,N_2023,N_2764);
or U5583 (N_5583,N_1298,N_699);
and U5584 (N_5584,N_2271,N_2279);
nor U5585 (N_5585,N_186,N_1525);
or U5586 (N_5586,N_93,N_2891);
or U5587 (N_5587,N_2022,N_976);
nand U5588 (N_5588,N_118,N_2608);
or U5589 (N_5589,N_107,N_809);
or U5590 (N_5590,N_1054,N_672);
and U5591 (N_5591,N_1517,N_2431);
nor U5592 (N_5592,N_283,N_2742);
and U5593 (N_5593,N_1217,N_831);
or U5594 (N_5594,N_2268,N_2119);
nor U5595 (N_5595,N_2549,N_1083);
and U5596 (N_5596,N_364,N_1925);
and U5597 (N_5597,N_13,N_2666);
nand U5598 (N_5598,N_706,N_698);
and U5599 (N_5599,N_591,N_218);
nor U5600 (N_5600,N_2506,N_2207);
nand U5601 (N_5601,N_2111,N_531);
nand U5602 (N_5602,N_727,N_1091);
and U5603 (N_5603,N_1478,N_1141);
nor U5604 (N_5604,N_2228,N_991);
nor U5605 (N_5605,N_213,N_1137);
nand U5606 (N_5606,N_2493,N_494);
or U5607 (N_5607,N_1923,N_1851);
and U5608 (N_5608,N_642,N_1262);
nand U5609 (N_5609,N_2259,N_890);
nor U5610 (N_5610,N_2265,N_1973);
and U5611 (N_5611,N_2758,N_196);
and U5612 (N_5612,N_1430,N_956);
xnor U5613 (N_5613,N_827,N_1697);
nor U5614 (N_5614,N_1492,N_563);
and U5615 (N_5615,N_1882,N_308);
nor U5616 (N_5616,N_955,N_1613);
xnor U5617 (N_5617,N_198,N_2643);
and U5618 (N_5618,N_2885,N_34);
nor U5619 (N_5619,N_1448,N_2506);
nor U5620 (N_5620,N_359,N_2916);
nor U5621 (N_5621,N_2662,N_2340);
or U5622 (N_5622,N_32,N_2884);
nand U5623 (N_5623,N_452,N_1664);
or U5624 (N_5624,N_2438,N_2544);
and U5625 (N_5625,N_348,N_210);
nand U5626 (N_5626,N_121,N_468);
nor U5627 (N_5627,N_2307,N_840);
and U5628 (N_5628,N_1699,N_531);
xor U5629 (N_5629,N_1105,N_15);
and U5630 (N_5630,N_2818,N_678);
or U5631 (N_5631,N_2600,N_2783);
nor U5632 (N_5632,N_947,N_2942);
nand U5633 (N_5633,N_1591,N_324);
xor U5634 (N_5634,N_2463,N_2926);
nor U5635 (N_5635,N_2010,N_2454);
nand U5636 (N_5636,N_1366,N_2386);
and U5637 (N_5637,N_2203,N_937);
or U5638 (N_5638,N_2531,N_154);
or U5639 (N_5639,N_1792,N_817);
nor U5640 (N_5640,N_391,N_2940);
and U5641 (N_5641,N_820,N_1752);
xnor U5642 (N_5642,N_1461,N_159);
and U5643 (N_5643,N_1414,N_1788);
and U5644 (N_5644,N_98,N_1488);
nor U5645 (N_5645,N_2730,N_2567);
xor U5646 (N_5646,N_417,N_768);
nor U5647 (N_5647,N_670,N_1324);
or U5648 (N_5648,N_1720,N_2951);
and U5649 (N_5649,N_821,N_1652);
or U5650 (N_5650,N_539,N_1073);
xor U5651 (N_5651,N_342,N_2697);
or U5652 (N_5652,N_497,N_93);
nor U5653 (N_5653,N_2889,N_1590);
or U5654 (N_5654,N_1206,N_1489);
and U5655 (N_5655,N_2939,N_1118);
nand U5656 (N_5656,N_1567,N_1091);
or U5657 (N_5657,N_1365,N_403);
xnor U5658 (N_5658,N_1434,N_2241);
or U5659 (N_5659,N_554,N_774);
nand U5660 (N_5660,N_2825,N_1310);
or U5661 (N_5661,N_670,N_416);
nor U5662 (N_5662,N_105,N_2576);
nor U5663 (N_5663,N_2898,N_1640);
or U5664 (N_5664,N_98,N_2636);
nand U5665 (N_5665,N_1984,N_553);
xnor U5666 (N_5666,N_2242,N_1331);
xnor U5667 (N_5667,N_2904,N_810);
nand U5668 (N_5668,N_393,N_2716);
nand U5669 (N_5669,N_1238,N_2933);
nor U5670 (N_5670,N_861,N_1686);
or U5671 (N_5671,N_2979,N_2800);
and U5672 (N_5672,N_2880,N_340);
xor U5673 (N_5673,N_1121,N_56);
and U5674 (N_5674,N_1122,N_524);
nor U5675 (N_5675,N_2291,N_1109);
and U5676 (N_5676,N_252,N_2734);
nand U5677 (N_5677,N_2208,N_1641);
and U5678 (N_5678,N_2498,N_139);
and U5679 (N_5679,N_2439,N_1742);
and U5680 (N_5680,N_947,N_2505);
xnor U5681 (N_5681,N_2251,N_886);
nor U5682 (N_5682,N_2061,N_398);
or U5683 (N_5683,N_2519,N_450);
and U5684 (N_5684,N_802,N_2845);
or U5685 (N_5685,N_2084,N_1840);
or U5686 (N_5686,N_356,N_725);
xnor U5687 (N_5687,N_2069,N_2609);
and U5688 (N_5688,N_229,N_760);
and U5689 (N_5689,N_227,N_1077);
and U5690 (N_5690,N_169,N_352);
and U5691 (N_5691,N_1821,N_2558);
or U5692 (N_5692,N_128,N_336);
or U5693 (N_5693,N_1416,N_130);
nand U5694 (N_5694,N_246,N_975);
or U5695 (N_5695,N_2036,N_1389);
nor U5696 (N_5696,N_1156,N_2945);
xor U5697 (N_5697,N_2028,N_965);
nor U5698 (N_5698,N_319,N_1236);
xor U5699 (N_5699,N_2609,N_1266);
nor U5700 (N_5700,N_2499,N_1185);
nor U5701 (N_5701,N_2362,N_2864);
or U5702 (N_5702,N_1346,N_757);
or U5703 (N_5703,N_70,N_2850);
or U5704 (N_5704,N_1962,N_407);
and U5705 (N_5705,N_2204,N_2025);
and U5706 (N_5706,N_988,N_2973);
xor U5707 (N_5707,N_1736,N_747);
xnor U5708 (N_5708,N_1224,N_741);
nand U5709 (N_5709,N_280,N_1950);
nor U5710 (N_5710,N_1682,N_161);
or U5711 (N_5711,N_1274,N_584);
or U5712 (N_5712,N_1125,N_914);
or U5713 (N_5713,N_2524,N_378);
or U5714 (N_5714,N_2262,N_832);
nor U5715 (N_5715,N_1928,N_257);
or U5716 (N_5716,N_150,N_2846);
xor U5717 (N_5717,N_1582,N_95);
nand U5718 (N_5718,N_136,N_149);
and U5719 (N_5719,N_2773,N_1957);
nor U5720 (N_5720,N_740,N_1462);
and U5721 (N_5721,N_680,N_2008);
and U5722 (N_5722,N_654,N_919);
xor U5723 (N_5723,N_2222,N_888);
nand U5724 (N_5724,N_653,N_2523);
nand U5725 (N_5725,N_2345,N_1751);
or U5726 (N_5726,N_2179,N_1503);
nand U5727 (N_5727,N_1380,N_2261);
or U5728 (N_5728,N_2536,N_1547);
or U5729 (N_5729,N_95,N_2806);
nand U5730 (N_5730,N_953,N_2539);
nand U5731 (N_5731,N_2179,N_2914);
nor U5732 (N_5732,N_2360,N_1174);
nand U5733 (N_5733,N_1769,N_1425);
xnor U5734 (N_5734,N_2742,N_393);
nor U5735 (N_5735,N_1277,N_2548);
or U5736 (N_5736,N_2747,N_1629);
and U5737 (N_5737,N_2433,N_2694);
nor U5738 (N_5738,N_2876,N_2018);
nor U5739 (N_5739,N_2192,N_2711);
xor U5740 (N_5740,N_2617,N_1076);
or U5741 (N_5741,N_6,N_1281);
and U5742 (N_5742,N_2520,N_909);
or U5743 (N_5743,N_2227,N_2989);
nor U5744 (N_5744,N_2438,N_1497);
nand U5745 (N_5745,N_124,N_383);
xor U5746 (N_5746,N_672,N_1619);
nor U5747 (N_5747,N_2430,N_1529);
or U5748 (N_5748,N_839,N_682);
xnor U5749 (N_5749,N_619,N_2843);
and U5750 (N_5750,N_591,N_1752);
and U5751 (N_5751,N_1642,N_322);
nor U5752 (N_5752,N_668,N_1876);
nor U5753 (N_5753,N_1251,N_1797);
nor U5754 (N_5754,N_2723,N_920);
or U5755 (N_5755,N_2442,N_1711);
nand U5756 (N_5756,N_1980,N_2201);
nand U5757 (N_5757,N_2674,N_998);
xnor U5758 (N_5758,N_2724,N_815);
nor U5759 (N_5759,N_2558,N_2176);
nor U5760 (N_5760,N_2764,N_33);
nand U5761 (N_5761,N_1115,N_363);
and U5762 (N_5762,N_431,N_2257);
and U5763 (N_5763,N_1307,N_2702);
nor U5764 (N_5764,N_118,N_1296);
and U5765 (N_5765,N_513,N_2061);
or U5766 (N_5766,N_2868,N_1907);
and U5767 (N_5767,N_2482,N_388);
and U5768 (N_5768,N_459,N_2471);
nand U5769 (N_5769,N_1592,N_1933);
nand U5770 (N_5770,N_2223,N_1253);
nor U5771 (N_5771,N_1418,N_2047);
xor U5772 (N_5772,N_2695,N_2826);
xor U5773 (N_5773,N_1683,N_1244);
and U5774 (N_5774,N_586,N_981);
or U5775 (N_5775,N_2921,N_139);
xor U5776 (N_5776,N_1853,N_1501);
or U5777 (N_5777,N_1109,N_781);
nand U5778 (N_5778,N_2113,N_2375);
and U5779 (N_5779,N_782,N_2685);
or U5780 (N_5780,N_2027,N_2804);
nand U5781 (N_5781,N_1988,N_1941);
or U5782 (N_5782,N_2411,N_958);
xnor U5783 (N_5783,N_1588,N_2144);
or U5784 (N_5784,N_811,N_1158);
nor U5785 (N_5785,N_1827,N_185);
nand U5786 (N_5786,N_1366,N_914);
nand U5787 (N_5787,N_1632,N_1731);
xor U5788 (N_5788,N_556,N_1831);
or U5789 (N_5789,N_2157,N_1532);
and U5790 (N_5790,N_2182,N_2994);
or U5791 (N_5791,N_319,N_2181);
nand U5792 (N_5792,N_1866,N_1611);
nand U5793 (N_5793,N_628,N_1815);
and U5794 (N_5794,N_315,N_795);
nor U5795 (N_5795,N_1437,N_668);
nor U5796 (N_5796,N_2163,N_2022);
and U5797 (N_5797,N_2575,N_811);
nand U5798 (N_5798,N_1089,N_2281);
nor U5799 (N_5799,N_2448,N_721);
nand U5800 (N_5800,N_1770,N_1501);
and U5801 (N_5801,N_2964,N_2776);
xnor U5802 (N_5802,N_1216,N_79);
or U5803 (N_5803,N_1203,N_1298);
nor U5804 (N_5804,N_1642,N_95);
nor U5805 (N_5805,N_17,N_2505);
xor U5806 (N_5806,N_612,N_2411);
nand U5807 (N_5807,N_507,N_1425);
and U5808 (N_5808,N_1831,N_2807);
nand U5809 (N_5809,N_1958,N_2608);
nor U5810 (N_5810,N_498,N_825);
nand U5811 (N_5811,N_195,N_2062);
xor U5812 (N_5812,N_2214,N_1757);
or U5813 (N_5813,N_453,N_618);
xnor U5814 (N_5814,N_2525,N_1535);
nand U5815 (N_5815,N_263,N_1685);
and U5816 (N_5816,N_549,N_2165);
xor U5817 (N_5817,N_1646,N_298);
or U5818 (N_5818,N_105,N_1228);
nor U5819 (N_5819,N_1631,N_2717);
or U5820 (N_5820,N_833,N_1206);
nor U5821 (N_5821,N_2706,N_1511);
nor U5822 (N_5822,N_1946,N_263);
nor U5823 (N_5823,N_1398,N_2134);
or U5824 (N_5824,N_945,N_2820);
and U5825 (N_5825,N_1140,N_1504);
or U5826 (N_5826,N_1055,N_837);
xor U5827 (N_5827,N_2606,N_1845);
xnor U5828 (N_5828,N_2531,N_1601);
nor U5829 (N_5829,N_17,N_1434);
nor U5830 (N_5830,N_1240,N_1698);
and U5831 (N_5831,N_863,N_150);
nor U5832 (N_5832,N_2351,N_1554);
or U5833 (N_5833,N_835,N_1870);
nand U5834 (N_5834,N_2238,N_872);
nor U5835 (N_5835,N_2939,N_860);
and U5836 (N_5836,N_1745,N_272);
or U5837 (N_5837,N_2301,N_2494);
xnor U5838 (N_5838,N_1890,N_558);
nor U5839 (N_5839,N_739,N_294);
or U5840 (N_5840,N_1118,N_382);
and U5841 (N_5841,N_2584,N_202);
nor U5842 (N_5842,N_2691,N_237);
nor U5843 (N_5843,N_2827,N_122);
nor U5844 (N_5844,N_1679,N_373);
and U5845 (N_5845,N_131,N_2945);
nor U5846 (N_5846,N_2982,N_2561);
nand U5847 (N_5847,N_1620,N_1273);
nand U5848 (N_5848,N_987,N_581);
nor U5849 (N_5849,N_2341,N_2505);
or U5850 (N_5850,N_1806,N_1136);
nor U5851 (N_5851,N_1445,N_121);
nor U5852 (N_5852,N_432,N_398);
xnor U5853 (N_5853,N_1957,N_1637);
or U5854 (N_5854,N_2402,N_22);
nand U5855 (N_5855,N_1653,N_1543);
and U5856 (N_5856,N_624,N_435);
and U5857 (N_5857,N_970,N_2696);
or U5858 (N_5858,N_486,N_316);
or U5859 (N_5859,N_1140,N_1185);
nand U5860 (N_5860,N_1445,N_2362);
and U5861 (N_5861,N_2202,N_1703);
nor U5862 (N_5862,N_917,N_1588);
nand U5863 (N_5863,N_112,N_1622);
or U5864 (N_5864,N_1964,N_980);
or U5865 (N_5865,N_665,N_2542);
nor U5866 (N_5866,N_2941,N_1128);
nand U5867 (N_5867,N_200,N_680);
nand U5868 (N_5868,N_1267,N_2126);
and U5869 (N_5869,N_2511,N_2644);
or U5870 (N_5870,N_2546,N_679);
and U5871 (N_5871,N_2702,N_93);
or U5872 (N_5872,N_2965,N_1281);
and U5873 (N_5873,N_1937,N_1723);
nor U5874 (N_5874,N_2493,N_159);
nand U5875 (N_5875,N_2956,N_1654);
xnor U5876 (N_5876,N_838,N_2234);
nand U5877 (N_5877,N_602,N_812);
nor U5878 (N_5878,N_1496,N_205);
and U5879 (N_5879,N_2940,N_1507);
nor U5880 (N_5880,N_1701,N_1847);
xor U5881 (N_5881,N_2749,N_2956);
nand U5882 (N_5882,N_646,N_2798);
and U5883 (N_5883,N_897,N_927);
xor U5884 (N_5884,N_1040,N_475);
and U5885 (N_5885,N_1627,N_1572);
xnor U5886 (N_5886,N_493,N_2180);
nor U5887 (N_5887,N_2719,N_770);
or U5888 (N_5888,N_368,N_1950);
xor U5889 (N_5889,N_1392,N_851);
nand U5890 (N_5890,N_2660,N_158);
xnor U5891 (N_5891,N_1121,N_2840);
and U5892 (N_5892,N_1217,N_1250);
nor U5893 (N_5893,N_1728,N_2580);
xor U5894 (N_5894,N_1106,N_1244);
nor U5895 (N_5895,N_474,N_2688);
or U5896 (N_5896,N_1051,N_21);
or U5897 (N_5897,N_2473,N_2440);
nand U5898 (N_5898,N_2097,N_2534);
nor U5899 (N_5899,N_1912,N_2723);
nand U5900 (N_5900,N_1082,N_2251);
nand U5901 (N_5901,N_2749,N_2086);
xor U5902 (N_5902,N_1078,N_1690);
nand U5903 (N_5903,N_1573,N_1067);
nor U5904 (N_5904,N_1756,N_490);
and U5905 (N_5905,N_1468,N_2446);
xnor U5906 (N_5906,N_1030,N_2090);
nand U5907 (N_5907,N_501,N_2913);
or U5908 (N_5908,N_10,N_1586);
nand U5909 (N_5909,N_1360,N_911);
nand U5910 (N_5910,N_2666,N_155);
and U5911 (N_5911,N_2063,N_2313);
or U5912 (N_5912,N_1157,N_2154);
nand U5913 (N_5913,N_137,N_695);
nand U5914 (N_5914,N_2363,N_2555);
nor U5915 (N_5915,N_1591,N_757);
nor U5916 (N_5916,N_1128,N_396);
and U5917 (N_5917,N_2803,N_658);
or U5918 (N_5918,N_701,N_2004);
nand U5919 (N_5919,N_174,N_1546);
and U5920 (N_5920,N_2968,N_489);
or U5921 (N_5921,N_892,N_677);
nor U5922 (N_5922,N_1506,N_315);
and U5923 (N_5923,N_1216,N_1493);
nor U5924 (N_5924,N_2042,N_2559);
and U5925 (N_5925,N_1240,N_2267);
nor U5926 (N_5926,N_2222,N_409);
nand U5927 (N_5927,N_2126,N_1646);
nand U5928 (N_5928,N_967,N_1081);
and U5929 (N_5929,N_2081,N_2335);
or U5930 (N_5930,N_1470,N_857);
or U5931 (N_5931,N_1782,N_843);
or U5932 (N_5932,N_1742,N_2121);
nand U5933 (N_5933,N_723,N_425);
or U5934 (N_5934,N_707,N_1176);
or U5935 (N_5935,N_1841,N_1546);
nand U5936 (N_5936,N_1513,N_745);
nand U5937 (N_5937,N_2390,N_587);
nand U5938 (N_5938,N_394,N_2693);
and U5939 (N_5939,N_344,N_1727);
and U5940 (N_5940,N_374,N_2550);
nand U5941 (N_5941,N_291,N_1170);
and U5942 (N_5942,N_2026,N_650);
nand U5943 (N_5943,N_1619,N_96);
or U5944 (N_5944,N_99,N_1944);
nand U5945 (N_5945,N_2175,N_2801);
and U5946 (N_5946,N_2581,N_2356);
and U5947 (N_5947,N_1502,N_1046);
nor U5948 (N_5948,N_2837,N_343);
nand U5949 (N_5949,N_235,N_340);
nor U5950 (N_5950,N_1488,N_1669);
and U5951 (N_5951,N_1114,N_736);
xor U5952 (N_5952,N_1338,N_358);
nand U5953 (N_5953,N_2636,N_1973);
nor U5954 (N_5954,N_535,N_1821);
nor U5955 (N_5955,N_2229,N_1616);
and U5956 (N_5956,N_1695,N_1320);
and U5957 (N_5957,N_1984,N_113);
nand U5958 (N_5958,N_131,N_544);
nand U5959 (N_5959,N_43,N_1785);
nor U5960 (N_5960,N_2251,N_2772);
nand U5961 (N_5961,N_2941,N_2896);
xnor U5962 (N_5962,N_2088,N_1620);
and U5963 (N_5963,N_2767,N_1088);
xnor U5964 (N_5964,N_750,N_2864);
or U5965 (N_5965,N_2063,N_2816);
and U5966 (N_5966,N_1308,N_2763);
nand U5967 (N_5967,N_1627,N_953);
nand U5968 (N_5968,N_2266,N_876);
or U5969 (N_5969,N_2569,N_711);
xor U5970 (N_5970,N_2249,N_57);
or U5971 (N_5971,N_2304,N_1849);
and U5972 (N_5972,N_455,N_2974);
xnor U5973 (N_5973,N_2365,N_633);
or U5974 (N_5974,N_2731,N_922);
nand U5975 (N_5975,N_2998,N_917);
nor U5976 (N_5976,N_20,N_2295);
nor U5977 (N_5977,N_1199,N_2666);
and U5978 (N_5978,N_2703,N_2431);
nor U5979 (N_5979,N_154,N_1303);
xor U5980 (N_5980,N_2087,N_2400);
nand U5981 (N_5981,N_1787,N_887);
or U5982 (N_5982,N_1627,N_251);
and U5983 (N_5983,N_2486,N_639);
and U5984 (N_5984,N_1074,N_2439);
or U5985 (N_5985,N_898,N_796);
nor U5986 (N_5986,N_376,N_1105);
nand U5987 (N_5987,N_1372,N_55);
nand U5988 (N_5988,N_884,N_2982);
and U5989 (N_5989,N_2960,N_1777);
and U5990 (N_5990,N_1796,N_1855);
and U5991 (N_5991,N_2400,N_2501);
nor U5992 (N_5992,N_611,N_2666);
nand U5993 (N_5993,N_2473,N_801);
or U5994 (N_5994,N_1937,N_2066);
and U5995 (N_5995,N_252,N_1318);
or U5996 (N_5996,N_1241,N_1497);
and U5997 (N_5997,N_347,N_2693);
nand U5998 (N_5998,N_1485,N_2243);
xnor U5999 (N_5999,N_1215,N_2032);
nor U6000 (N_6000,N_5876,N_4278);
or U6001 (N_6001,N_5210,N_4411);
or U6002 (N_6002,N_3593,N_4515);
or U6003 (N_6003,N_3007,N_5667);
xnor U6004 (N_6004,N_4210,N_4535);
nand U6005 (N_6005,N_5713,N_3661);
nand U6006 (N_6006,N_3194,N_5726);
or U6007 (N_6007,N_3099,N_4125);
and U6008 (N_6008,N_5441,N_4438);
nand U6009 (N_6009,N_3304,N_4156);
and U6010 (N_6010,N_3455,N_5609);
xor U6011 (N_6011,N_3765,N_5179);
nand U6012 (N_6012,N_5197,N_5243);
nor U6013 (N_6013,N_5767,N_4033);
and U6014 (N_6014,N_4476,N_5585);
and U6015 (N_6015,N_5226,N_4766);
xor U6016 (N_6016,N_4936,N_4767);
or U6017 (N_6017,N_5718,N_3047);
xor U6018 (N_6018,N_5323,N_5459);
or U6019 (N_6019,N_4858,N_3915);
xnor U6020 (N_6020,N_3408,N_4857);
xor U6021 (N_6021,N_5056,N_5989);
or U6022 (N_6022,N_3260,N_3161);
nand U6023 (N_6023,N_3750,N_3509);
or U6024 (N_6024,N_4347,N_4258);
nand U6025 (N_6025,N_3688,N_5329);
nand U6026 (N_6026,N_4869,N_4913);
nand U6027 (N_6027,N_4630,N_4626);
nand U6028 (N_6028,N_4350,N_4493);
and U6029 (N_6029,N_4245,N_5270);
and U6030 (N_6030,N_5305,N_4520);
xor U6031 (N_6031,N_5768,N_3851);
and U6032 (N_6032,N_4610,N_5065);
or U6033 (N_6033,N_5214,N_3555);
and U6034 (N_6034,N_4206,N_5551);
nand U6035 (N_6035,N_4290,N_3682);
or U6036 (N_6036,N_3764,N_3998);
and U6037 (N_6037,N_3436,N_3002);
xnor U6038 (N_6038,N_3559,N_4066);
and U6039 (N_6039,N_3320,N_3654);
or U6040 (N_6040,N_5389,N_3604);
or U6041 (N_6041,N_5165,N_4804);
and U6042 (N_6042,N_4485,N_4542);
or U6043 (N_6043,N_3423,N_4504);
nand U6044 (N_6044,N_3535,N_5310);
or U6045 (N_6045,N_3933,N_3698);
or U6046 (N_6046,N_4590,N_4802);
or U6047 (N_6047,N_4376,N_4458);
or U6048 (N_6048,N_5645,N_5028);
and U6049 (N_6049,N_5685,N_5984);
nand U6050 (N_6050,N_5793,N_5646);
and U6051 (N_6051,N_5422,N_4334);
or U6052 (N_6052,N_3967,N_3692);
nand U6053 (N_6053,N_3263,N_5172);
or U6054 (N_6054,N_3174,N_3339);
and U6055 (N_6055,N_5890,N_4046);
and U6056 (N_6056,N_4108,N_4680);
or U6057 (N_6057,N_4027,N_4712);
nand U6058 (N_6058,N_3272,N_5674);
nand U6059 (N_6059,N_4615,N_3873);
and U6060 (N_6060,N_3500,N_4216);
nand U6061 (N_6061,N_5786,N_3222);
nand U6062 (N_6062,N_5633,N_5791);
nand U6063 (N_6063,N_4600,N_4084);
and U6064 (N_6064,N_3034,N_5101);
or U6065 (N_6065,N_5190,N_3662);
nor U6066 (N_6066,N_5657,N_4616);
or U6067 (N_6067,N_3261,N_4763);
nand U6068 (N_6068,N_4259,N_5727);
or U6069 (N_6069,N_3628,N_3085);
or U6070 (N_6070,N_5591,N_4338);
and U6071 (N_6071,N_4753,N_5637);
nor U6072 (N_6072,N_4888,N_5140);
nand U6073 (N_6073,N_3783,N_3714);
nand U6074 (N_6074,N_5517,N_3429);
or U6075 (N_6075,N_4558,N_4446);
or U6076 (N_6076,N_3126,N_4381);
nor U6077 (N_6077,N_5852,N_4329);
nand U6078 (N_6078,N_3010,N_5449);
nand U6079 (N_6079,N_3273,N_4380);
nand U6080 (N_6080,N_5057,N_3317);
xor U6081 (N_6081,N_3301,N_3486);
xor U6082 (N_6082,N_5639,N_3872);
nand U6083 (N_6083,N_3288,N_5209);
nand U6084 (N_6084,N_4693,N_4544);
or U6085 (N_6085,N_3674,N_5952);
nor U6086 (N_6086,N_4647,N_4408);
nor U6087 (N_6087,N_3954,N_5135);
nor U6088 (N_6088,N_4147,N_3163);
nor U6089 (N_6089,N_3380,N_4965);
and U6090 (N_6090,N_4690,N_4636);
nand U6091 (N_6091,N_4429,N_5905);
nor U6092 (N_6092,N_4022,N_4249);
or U6093 (N_6093,N_5312,N_5180);
nand U6094 (N_6094,N_5572,N_3746);
and U6095 (N_6095,N_5029,N_4538);
nor U6096 (N_6096,N_3665,N_4586);
nor U6097 (N_6097,N_4394,N_3969);
nor U6098 (N_6098,N_4549,N_5117);
or U6099 (N_6099,N_4100,N_5898);
or U6100 (N_6100,N_5353,N_3516);
nor U6101 (N_6101,N_5799,N_4436);
or U6102 (N_6102,N_3158,N_4642);
or U6103 (N_6103,N_5332,N_5527);
nand U6104 (N_6104,N_3930,N_5297);
or U6105 (N_6105,N_5687,N_5625);
or U6106 (N_6106,N_4820,N_3697);
and U6107 (N_6107,N_4555,N_3710);
xnor U6108 (N_6108,N_5651,N_3564);
xor U6109 (N_6109,N_5245,N_4218);
or U6110 (N_6110,N_4724,N_4089);
or U6111 (N_6111,N_3849,N_4010);
nor U6112 (N_6112,N_3122,N_4410);
nand U6113 (N_6113,N_4826,N_4025);
nor U6114 (N_6114,N_5139,N_4990);
xnor U6115 (N_6115,N_5457,N_4505);
nor U6116 (N_6116,N_5322,N_4704);
nor U6117 (N_6117,N_3470,N_5066);
nor U6118 (N_6118,N_3217,N_4514);
nor U6119 (N_6119,N_4568,N_4328);
nor U6120 (N_6120,N_5397,N_4934);
nor U6121 (N_6121,N_5272,N_5155);
and U6122 (N_6122,N_3570,N_4933);
xnor U6123 (N_6123,N_3501,N_5588);
nand U6124 (N_6124,N_3229,N_4565);
nand U6125 (N_6125,N_5159,N_5684);
nand U6126 (N_6126,N_5365,N_3031);
nand U6127 (N_6127,N_3305,N_5394);
or U6128 (N_6128,N_5286,N_5881);
nor U6129 (N_6129,N_3585,N_5105);
and U6130 (N_6130,N_5529,N_4006);
or U6131 (N_6131,N_3556,N_3666);
nand U6132 (N_6132,N_3493,N_3656);
nor U6133 (N_6133,N_3601,N_4403);
and U6134 (N_6134,N_3241,N_5544);
nand U6135 (N_6135,N_3473,N_5947);
nand U6136 (N_6136,N_4839,N_3799);
or U6137 (N_6137,N_5604,N_4669);
and U6138 (N_6138,N_4134,N_5194);
or U6139 (N_6139,N_4162,N_5019);
or U6140 (N_6140,N_5508,N_4070);
xor U6141 (N_6141,N_4465,N_3647);
nand U6142 (N_6142,N_5118,N_4694);
or U6143 (N_6143,N_4998,N_5642);
and U6144 (N_6144,N_3120,N_4805);
and U6145 (N_6145,N_5002,N_3013);
and U6146 (N_6146,N_4227,N_4975);
nand U6147 (N_6147,N_5319,N_4152);
nand U6148 (N_6148,N_4676,N_3311);
xnor U6149 (N_6149,N_5149,N_5317);
xor U6150 (N_6150,N_4357,N_4614);
and U6151 (N_6151,N_5941,N_5106);
nor U6152 (N_6152,N_3676,N_3011);
nor U6153 (N_6153,N_4672,N_4984);
nand U6154 (N_6154,N_3921,N_3021);
nor U6155 (N_6155,N_5150,N_3622);
or U6156 (N_6156,N_4234,N_3964);
nand U6157 (N_6157,N_5315,N_5949);
and U6158 (N_6158,N_4199,N_4736);
or U6159 (N_6159,N_3098,N_5831);
nand U6160 (N_6160,N_4247,N_5448);
or U6161 (N_6161,N_5320,N_3822);
nor U6162 (N_6162,N_3402,N_5443);
and U6163 (N_6163,N_5933,N_5782);
or U6164 (N_6164,N_5195,N_4051);
nand U6165 (N_6165,N_4881,N_3356);
nor U6166 (N_6166,N_4194,N_4670);
or U6167 (N_6167,N_3059,N_5838);
xor U6168 (N_6168,N_3206,N_3538);
xnor U6169 (N_6169,N_4132,N_4124);
and U6170 (N_6170,N_4226,N_4917);
nand U6171 (N_6171,N_5556,N_4738);
nand U6172 (N_6172,N_3447,N_5186);
nand U6173 (N_6173,N_3431,N_4903);
nand U6174 (N_6174,N_5024,N_5212);
or U6175 (N_6175,N_4448,N_5917);
xnor U6176 (N_6176,N_5559,N_5496);
and U6177 (N_6177,N_3097,N_3815);
or U6178 (N_6178,N_5673,N_4551);
or U6179 (N_6179,N_4049,N_3258);
xnor U6180 (N_6180,N_5380,N_5271);
nor U6181 (N_6181,N_4282,N_4640);
nor U6182 (N_6182,N_4102,N_4407);
and U6183 (N_6183,N_3721,N_5452);
and U6184 (N_6184,N_3796,N_5045);
nand U6185 (N_6185,N_3411,N_3325);
and U6186 (N_6186,N_5916,N_3322);
nor U6187 (N_6187,N_5853,N_5256);
nor U6188 (N_6188,N_4479,N_5914);
nand U6189 (N_6189,N_4516,N_5951);
and U6190 (N_6190,N_4528,N_3850);
nor U6191 (N_6191,N_3882,N_4849);
nand U6192 (N_6192,N_3388,N_4176);
or U6193 (N_6193,N_4360,N_3179);
or U6194 (N_6194,N_5574,N_4629);
nor U6195 (N_6195,N_4511,N_4588);
or U6196 (N_6196,N_4644,N_3949);
or U6197 (N_6197,N_5849,N_3513);
or U6198 (N_6198,N_4868,N_4268);
nor U6199 (N_6199,N_3005,N_3956);
and U6200 (N_6200,N_4842,N_3887);
and U6201 (N_6201,N_3042,N_4293);
nand U6202 (N_6202,N_4427,N_5497);
nor U6203 (N_6203,N_4193,N_3549);
or U6204 (N_6204,N_4923,N_5541);
and U6205 (N_6205,N_3994,N_4424);
nand U6206 (N_6206,N_5418,N_4466);
nand U6207 (N_6207,N_4215,N_5971);
nand U6208 (N_6208,N_3706,N_4203);
and U6209 (N_6209,N_5828,N_3040);
and U6210 (N_6210,N_5942,N_4365);
nand U6211 (N_6211,N_5946,N_5558);
or U6212 (N_6212,N_3723,N_4821);
nand U6213 (N_6213,N_5217,N_5439);
and U6214 (N_6214,N_3345,N_4035);
nand U6215 (N_6215,N_4378,N_5668);
and U6216 (N_6216,N_5089,N_5247);
and U6217 (N_6217,N_5652,N_3597);
xor U6218 (N_6218,N_4816,N_5611);
nand U6219 (N_6219,N_4294,N_5033);
nand U6220 (N_6220,N_3858,N_3484);
or U6221 (N_6221,N_3213,N_3485);
nor U6222 (N_6222,N_5521,N_3342);
xor U6223 (N_6223,N_5754,N_4583);
or U6224 (N_6224,N_3791,N_3135);
xnor U6225 (N_6225,N_4748,N_5580);
nand U6226 (N_6226,N_3862,N_3498);
and U6227 (N_6227,N_3833,N_4951);
nand U6228 (N_6228,N_3648,N_4488);
nor U6229 (N_6229,N_4886,N_4628);
and U6230 (N_6230,N_5096,N_5265);
or U6231 (N_6231,N_4081,N_5442);
and U6232 (N_6232,N_5965,N_3543);
xnor U6233 (N_6233,N_4159,N_4937);
nand U6234 (N_6234,N_4317,N_5511);
and U6235 (N_6235,N_3449,N_4279);
xnor U6236 (N_6236,N_5489,N_4609);
xnor U6237 (N_6237,N_3175,N_5746);
nor U6238 (N_6238,N_3965,N_5880);
nor U6239 (N_6239,N_5676,N_3720);
nor U6240 (N_6240,N_3640,N_3053);
xor U6241 (N_6241,N_3468,N_5144);
nand U6242 (N_6242,N_4085,N_4418);
or U6243 (N_6243,N_5598,N_4617);
and U6244 (N_6244,N_3702,N_5552);
or U6245 (N_6245,N_3909,N_5338);
nor U6246 (N_6246,N_3772,N_4580);
and U6247 (N_6247,N_4569,N_5086);
or U6248 (N_6248,N_4495,N_4456);
and U6249 (N_6249,N_4652,N_4737);
nor U6250 (N_6250,N_3458,N_3871);
nand U6251 (N_6251,N_4540,N_5249);
nand U6252 (N_6252,N_4506,N_5691);
nand U6253 (N_6253,N_3557,N_4143);
or U6254 (N_6254,N_4797,N_3739);
or U6255 (N_6255,N_5675,N_4856);
and U6256 (N_6256,N_3530,N_5376);
nor U6257 (N_6257,N_3707,N_3992);
nor U6258 (N_6258,N_3172,N_3568);
or U6259 (N_6259,N_4808,N_5069);
nor U6260 (N_6260,N_5013,N_3550);
nor U6261 (N_6261,N_5901,N_4047);
nand U6262 (N_6262,N_5863,N_3963);
nor U6263 (N_6263,N_5520,N_4061);
nor U6264 (N_6264,N_4760,N_4899);
and U6265 (N_6265,N_4799,N_3296);
nor U6266 (N_6266,N_4341,N_5557);
or U6267 (N_6267,N_3925,N_4235);
or U6268 (N_6268,N_3582,N_5824);
and U6269 (N_6269,N_5549,N_5886);
nor U6270 (N_6270,N_4167,N_3962);
xnor U6271 (N_6271,N_5475,N_5395);
nor U6272 (N_6272,N_4008,N_3328);
and U6273 (N_6273,N_5769,N_5950);
and U6274 (N_6274,N_4757,N_4426);
and U6275 (N_6275,N_3542,N_5386);
xnor U6276 (N_6276,N_4281,N_5283);
and U6277 (N_6277,N_4324,N_5367);
nor U6278 (N_6278,N_3924,N_3511);
and U6279 (N_6279,N_3074,N_5648);
or U6280 (N_6280,N_3495,N_5083);
nand U6281 (N_6281,N_4959,N_4525);
nand U6282 (N_6282,N_5498,N_5641);
or U6283 (N_6283,N_5114,N_4011);
nand U6284 (N_6284,N_4725,N_4039);
and U6285 (N_6285,N_4920,N_3983);
or U6286 (N_6286,N_5023,N_5973);
nand U6287 (N_6287,N_4289,N_5597);
and U6288 (N_6288,N_5766,N_4579);
xor U6289 (N_6289,N_4063,N_4322);
or U6290 (N_6290,N_4020,N_4863);
or U6291 (N_6291,N_5396,N_5430);
nor U6292 (N_6292,N_5783,N_3294);
or U6293 (N_6293,N_3270,N_4607);
or U6294 (N_6294,N_4859,N_4140);
nand U6295 (N_6295,N_5470,N_3806);
nand U6296 (N_6296,N_5358,N_4337);
and U6297 (N_6297,N_5918,N_4860);
or U6298 (N_6298,N_5739,N_4393);
nand U6299 (N_6299,N_5812,N_5343);
and U6300 (N_6300,N_3978,N_5382);
nand U6301 (N_6301,N_4599,N_3818);
nand U6302 (N_6302,N_4911,N_3912);
or U6303 (N_6303,N_4603,N_5492);
xnor U6304 (N_6304,N_3279,N_3156);
or U6305 (N_6305,N_3425,N_5036);
and U6306 (N_6306,N_4929,N_5887);
and U6307 (N_6307,N_5129,N_5522);
or U6308 (N_6308,N_5502,N_4741);
and U6309 (N_6309,N_3607,N_5910);
nor U6310 (N_6310,N_5125,N_3732);
and U6311 (N_6311,N_3981,N_3087);
nor U6312 (N_6312,N_5299,N_5653);
nor U6313 (N_6313,N_4300,N_3396);
or U6314 (N_6314,N_4185,N_5590);
nand U6315 (N_6315,N_4878,N_5578);
and U6316 (N_6316,N_5935,N_4349);
nor U6317 (N_6317,N_4751,N_4562);
nand U6318 (N_6318,N_3731,N_5224);
nor U6319 (N_6319,N_5595,N_3390);
nor U6320 (N_6320,N_4204,N_3023);
xor U6321 (N_6321,N_5432,N_4999);
xnor U6322 (N_6322,N_5316,N_4960);
and U6323 (N_6323,N_5907,N_3914);
or U6324 (N_6324,N_5716,N_3281);
and U6325 (N_6325,N_4734,N_3793);
or U6326 (N_6326,N_3885,N_3551);
or U6327 (N_6327,N_4634,N_4735);
xor U6328 (N_6328,N_3290,N_4499);
nand U6329 (N_6329,N_4405,N_3548);
xnor U6330 (N_6330,N_3341,N_3979);
or U6331 (N_6331,N_3743,N_5656);
xor U6332 (N_6332,N_3733,N_4351);
nor U6333 (N_6333,N_4284,N_3117);
and U6334 (N_6334,N_5304,N_5995);
and U6335 (N_6335,N_4703,N_4131);
nand U6336 (N_6336,N_5850,N_3326);
and U6337 (N_6337,N_5012,N_3957);
and U6338 (N_6338,N_3465,N_3366);
nand U6339 (N_6339,N_3381,N_5364);
and U6340 (N_6340,N_3028,N_4833);
nand U6341 (N_6341,N_5906,N_5514);
or U6342 (N_6342,N_4087,N_5373);
or U6343 (N_6343,N_3738,N_5875);
and U6344 (N_6344,N_4015,N_3859);
or U6345 (N_6345,N_3460,N_5576);
nand U6346 (N_6346,N_4158,N_4356);
xor U6347 (N_6347,N_4401,N_4487);
xnor U6348 (N_6348,N_5710,N_3330);
nand U6349 (N_6349,N_5415,N_4971);
or U6350 (N_6350,N_3173,N_5006);
and U6351 (N_6351,N_5908,N_4315);
nand U6352 (N_6352,N_3997,N_3609);
and U6353 (N_6353,N_5613,N_4439);
or U6354 (N_6354,N_5825,N_4449);
nand U6355 (N_6355,N_4497,N_3119);
and U6356 (N_6356,N_3908,N_3920);
nand U6357 (N_6357,N_4745,N_4930);
and U6358 (N_6358,N_4539,N_5251);
nand U6359 (N_6359,N_5963,N_5119);
nor U6360 (N_6360,N_3589,N_3846);
nand U6361 (N_6361,N_5870,N_3505);
or U6362 (N_6362,N_3183,N_4658);
nor U6363 (N_6363,N_5943,N_5133);
or U6364 (N_6364,N_5919,N_4252);
nand U6365 (N_6365,N_4208,N_4001);
and U6366 (N_6366,N_5131,N_5605);
and U6367 (N_6367,N_4945,N_4453);
nor U6368 (N_6368,N_5998,N_3427);
nor U6369 (N_6369,N_4082,N_4653);
and U6370 (N_6370,N_3623,N_5110);
nor U6371 (N_6371,N_3980,N_4581);
and U6372 (N_6372,N_4175,N_4601);
nand U6373 (N_6373,N_4837,N_3192);
nor U6374 (N_6374,N_3186,N_3030);
or U6375 (N_6375,N_5287,N_5956);
xor U6376 (N_6376,N_4952,N_5669);
and U6377 (N_6377,N_5344,N_4801);
or U6378 (N_6378,N_5438,N_4942);
nor U6379 (N_6379,N_3147,N_4787);
and U6380 (N_6380,N_3138,N_5911);
nand U6381 (N_6381,N_3986,N_4645);
or U6382 (N_6382,N_4437,N_5662);
nand U6383 (N_6383,N_4762,N_3160);
or U6384 (N_6384,N_4433,N_3324);
nor U6385 (N_6385,N_4094,N_3629);
or U6386 (N_6386,N_3901,N_5567);
nor U6387 (N_6387,N_5084,N_5242);
nor U6388 (N_6388,N_4872,N_3378);
nand U6389 (N_6389,N_4815,N_3718);
or U6390 (N_6390,N_5606,N_5680);
and U6391 (N_6391,N_3142,N_5072);
xor U6392 (N_6392,N_5034,N_4898);
nor U6393 (N_6393,N_5787,N_3347);
and U6394 (N_6394,N_4988,N_3233);
nor U6395 (N_6395,N_5506,N_3752);
and U6396 (N_6396,N_5339,N_5264);
xnor U6397 (N_6397,N_5371,N_4314);
nor U6398 (N_6398,N_3266,N_3941);
nor U6399 (N_6399,N_3779,N_4385);
or U6400 (N_6400,N_5399,N_3004);
or U6401 (N_6401,N_5839,N_3159);
nand U6402 (N_6402,N_5706,N_3017);
and U6403 (N_6403,N_3265,N_3152);
nor U6404 (N_6404,N_4973,N_5533);
nand U6405 (N_6405,N_3070,N_3045);
nand U6406 (N_6406,N_5760,N_4689);
and U6407 (N_6407,N_4931,N_5695);
or U6408 (N_6408,N_3019,N_4240);
nand U6409 (N_6409,N_3937,N_5189);
or U6410 (N_6410,N_3014,N_3536);
nor U6411 (N_6411,N_5733,N_4250);
nand U6412 (N_6412,N_3856,N_3695);
nor U6413 (N_6413,N_3323,N_5173);
or U6414 (N_6414,N_3776,N_5904);
xnor U6415 (N_6415,N_3284,N_5672);
xor U6416 (N_6416,N_3828,N_3510);
xor U6417 (N_6417,N_4639,N_4423);
nand U6418 (N_6418,N_4596,N_5524);
and U6419 (N_6419,N_4486,N_4744);
and U6420 (N_6420,N_5416,N_4894);
and U6421 (N_6421,N_5670,N_3988);
nand U6422 (N_6422,N_5335,N_5705);
or U6423 (N_6423,N_3065,N_4313);
nor U6424 (N_6424,N_3749,N_4391);
nor U6425 (N_6425,N_4148,N_4072);
xnor U6426 (N_6426,N_4026,N_4416);
nor U6427 (N_6427,N_4662,N_5143);
nand U6428 (N_6428,N_5883,N_5134);
nor U6429 (N_6429,N_3939,N_3006);
and U6430 (N_6430,N_5252,N_4963);
nand U6431 (N_6431,N_3679,N_3176);
nand U6432 (N_6432,N_5445,N_5798);
xor U6433 (N_6433,N_4865,N_5184);
and U6434 (N_6434,N_3015,N_5781);
and U6435 (N_6435,N_3811,N_3235);
xnor U6436 (N_6436,N_5509,N_4727);
nand U6437 (N_6437,N_4432,N_5618);
or U6438 (N_6438,N_3376,N_3391);
or U6439 (N_6439,N_4993,N_3781);
nor U6440 (N_6440,N_3035,N_3625);
nor U6441 (N_6441,N_4442,N_5778);
nand U6442 (N_6442,N_3121,N_3141);
nor U6443 (N_6443,N_4678,N_5814);
and U6444 (N_6444,N_4382,N_5679);
or U6445 (N_6445,N_5121,N_3221);
xor U6446 (N_6446,N_5811,N_4257);
or U6447 (N_6447,N_4320,N_3337);
nor U6448 (N_6448,N_4854,N_3927);
nand U6449 (N_6449,N_3309,N_3993);
xnor U6450 (N_6450,N_4556,N_3075);
or U6451 (N_6451,N_3621,N_3614);
or U6452 (N_6452,N_5630,N_4074);
xor U6453 (N_6453,N_5277,N_3515);
nand U6454 (N_6454,N_3095,N_4052);
nor U6455 (N_6455,N_3123,N_5161);
and U6456 (N_6456,N_4968,N_3802);
xnor U6457 (N_6457,N_3918,N_4981);
or U6458 (N_6458,N_4280,N_4253);
nor U6459 (N_6459,N_5753,N_4333);
nor U6460 (N_6460,N_4564,N_4827);
nand U6461 (N_6461,N_3533,N_3073);
nand U6462 (N_6462,N_4205,N_4950);
or U6463 (N_6463,N_5806,N_5239);
nor U6464 (N_6464,N_5145,N_4572);
and U6465 (N_6465,N_5342,N_3712);
xor U6466 (N_6466,N_5490,N_5017);
or U6467 (N_6467,N_5861,N_4062);
nand U6468 (N_6468,N_4631,N_4896);
or U6469 (N_6469,N_4790,N_4113);
and U6470 (N_6470,N_5234,N_4375);
xnor U6471 (N_6471,N_4450,N_3643);
nor U6472 (N_6472,N_4657,N_4261);
or U6473 (N_6473,N_3024,N_5259);
nor U6474 (N_6474,N_5388,N_3422);
nand U6475 (N_6475,N_3630,N_3365);
nor U6476 (N_6476,N_3291,N_5848);
nand U6477 (N_6477,N_4217,N_3816);
nand U6478 (N_6478,N_5219,N_3693);
nand U6479 (N_6479,N_3775,N_5537);
nor U6480 (N_6480,N_4552,N_3478);
or U6481 (N_6481,N_4780,N_4602);
nor U6482 (N_6482,N_5078,N_4832);
xnor U6483 (N_6483,N_3219,N_4743);
or U6484 (N_6484,N_5743,N_5756);
or U6485 (N_6485,N_4587,N_4608);
and U6486 (N_6486,N_4720,N_3448);
and U6487 (N_6487,N_5202,N_4604);
nand U6488 (N_6488,N_5157,N_3048);
nor U6489 (N_6489,N_5921,N_4784);
or U6490 (N_6490,N_4096,N_5465);
nand U6491 (N_6491,N_5289,N_3757);
nor U6492 (N_6492,N_5628,N_4422);
and U6493 (N_6493,N_3758,N_3225);
and U6494 (N_6494,N_4431,N_5041);
nand U6495 (N_6495,N_4793,N_4454);
nor U6496 (N_6496,N_5022,N_5295);
and U6497 (N_6497,N_5579,N_5154);
and U6498 (N_6498,N_4301,N_4684);
or U6499 (N_6499,N_5420,N_4164);
or U6500 (N_6500,N_3467,N_5187);
and U6501 (N_6501,N_4272,N_3606);
and U6502 (N_6502,N_4835,N_4445);
or U6503 (N_6503,N_3490,N_3267);
and U6504 (N_6504,N_5594,N_5405);
and U6505 (N_6505,N_5977,N_3973);
and U6506 (N_6506,N_5858,N_3360);
and U6507 (N_6507,N_5513,N_4718);
nand U6508 (N_6508,N_4028,N_3287);
nor U6509 (N_6509,N_5414,N_3841);
or U6510 (N_6510,N_3727,N_5532);
or U6511 (N_6511,N_3306,N_4949);
xor U6512 (N_6512,N_5638,N_4110);
nand U6513 (N_6513,N_5764,N_4153);
nor U6514 (N_6514,N_3384,N_5775);
or U6515 (N_6515,N_3991,N_4387);
and U6516 (N_6516,N_3504,N_4541);
nor U6517 (N_6517,N_3385,N_4870);
and U6518 (N_6518,N_3237,N_4352);
nor U6519 (N_6519,N_5737,N_3153);
and U6520 (N_6520,N_3835,N_5473);
nand U6521 (N_6521,N_5519,N_3906);
nor U6522 (N_6522,N_4633,N_3683);
and U6523 (N_6523,N_4146,N_3926);
and U6524 (N_6524,N_3708,N_5203);
nor U6525 (N_6525,N_5708,N_3343);
nand U6526 (N_6526,N_3754,N_5383);
and U6527 (N_6527,N_5030,N_3650);
nor U6528 (N_6528,N_3571,N_3910);
or U6529 (N_6529,N_4598,N_3329);
xor U6530 (N_6530,N_5829,N_3907);
xnor U6531 (N_6531,N_4764,N_5581);
nand U6532 (N_6532,N_5996,N_4907);
and U6533 (N_6533,N_4836,N_3715);
nand U6534 (N_6534,N_4032,N_5163);
nand U6535 (N_6535,N_5341,N_3608);
nor U6536 (N_6536,N_4526,N_5479);
and U6537 (N_6537,N_4478,N_5752);
xor U6538 (N_6538,N_4018,N_4248);
nand U6539 (N_6539,N_4656,N_5417);
xnor U6540 (N_6540,N_3081,N_4938);
and U6541 (N_6541,N_3327,N_3102);
and U6542 (N_6542,N_3353,N_4276);
nor U6543 (N_6543,N_5818,N_5221);
nand U6544 (N_6544,N_5491,N_3348);
and U6545 (N_6545,N_4585,N_3853);
nor U6546 (N_6546,N_3518,N_4500);
nand U6547 (N_6547,N_5974,N_5095);
nor U6548 (N_6548,N_4553,N_5360);
xor U6549 (N_6549,N_5817,N_3646);
nor U6550 (N_6550,N_3677,N_3145);
nand U6551 (N_6551,N_4021,N_4316);
or U6552 (N_6552,N_4413,N_4545);
and U6553 (N_6553,N_4823,N_5156);
and U6554 (N_6554,N_3373,N_3471);
nor U6555 (N_6555,N_3203,N_5621);
and U6556 (N_6556,N_4916,N_5816);
xor U6557 (N_6557,N_4323,N_3043);
or U6558 (N_6558,N_4775,N_5425);
and U6559 (N_6559,N_3077,N_3190);
and U6560 (N_6560,N_5777,N_4702);
nor U6561 (N_6561,N_5884,N_5333);
nor U6562 (N_6562,N_4384,N_5964);
nor U6563 (N_6563,N_4691,N_3526);
nor U6564 (N_6564,N_5027,N_5822);
and U6565 (N_6565,N_4919,N_5260);
nand U6566 (N_6566,N_4943,N_4298);
nor U6567 (N_6567,N_5525,N_4756);
and U6568 (N_6568,N_4776,N_3369);
nand U6569 (N_6569,N_4719,N_4012);
nand U6570 (N_6570,N_4447,N_4677);
nor U6571 (N_6571,N_5229,N_5719);
and U6572 (N_6572,N_3483,N_3067);
nand U6573 (N_6573,N_5619,N_4366);
or U6574 (N_6574,N_3826,N_3868);
nor U6575 (N_6575,N_3009,N_5873);
and U6576 (N_6576,N_3875,N_5855);
nor U6577 (N_6577,N_5988,N_3810);
nand U6578 (N_6578,N_3259,N_3737);
or U6579 (N_6579,N_4292,N_4575);
and U6580 (N_6580,N_5860,N_5393);
and U6581 (N_6581,N_5980,N_3293);
xor U6582 (N_6582,N_3821,N_5599);
and U6583 (N_6583,N_3845,N_4922);
nor U6584 (N_6584,N_3195,N_3139);
and U6585 (N_6585,N_5450,N_3199);
or U6586 (N_6586,N_4471,N_5000);
nor U6587 (N_6587,N_3798,N_5314);
nor U6588 (N_6588,N_5037,N_3769);
or U6589 (N_6589,N_3842,N_3745);
or U6590 (N_6590,N_3321,N_5090);
xor U6591 (N_6591,N_5300,N_4852);
or U6592 (N_6592,N_5403,N_5216);
nand U6593 (N_6593,N_5407,N_4291);
xnor U6594 (N_6594,N_4697,N_5426);
nand U6595 (N_6595,N_5324,N_3131);
nand U6596 (N_6596,N_5073,N_3522);
or U6597 (N_6597,N_4834,N_4713);
nand U6598 (N_6598,N_4961,N_5958);
or U6599 (N_6599,N_4312,N_3877);
and U6600 (N_6600,N_3935,N_5048);
nand U6601 (N_6601,N_5345,N_5035);
and U6602 (N_6602,N_3247,N_4142);
or U6603 (N_6603,N_4396,N_5120);
nor U6604 (N_6604,N_5966,N_5516);
and U6605 (N_6605,N_3426,N_5044);
and U6606 (N_6606,N_4303,N_3840);
nand U6607 (N_6607,N_3058,N_5185);
and U6608 (N_6608,N_3228,N_5944);
nand U6609 (N_6609,N_3946,N_5008);
nand U6610 (N_6610,N_4941,N_5001);
nand U6611 (N_6611,N_4367,N_4192);
or U6612 (N_6612,N_3494,N_5991);
nor U6613 (N_6613,N_4921,N_3285);
nor U6614 (N_6614,N_5985,N_3817);
nand U6615 (N_6615,N_5293,N_4758);
or U6616 (N_6616,N_3902,N_5288);
nor U6617 (N_6617,N_3371,N_5292);
and U6618 (N_6618,N_3636,N_4390);
or U6619 (N_6619,N_4980,N_3397);
nor U6620 (N_6620,N_3655,N_4696);
nand U6621 (N_6621,N_5757,N_4244);
or U6622 (N_6622,N_3162,N_5206);
nor U6623 (N_6623,N_3091,N_4174);
or U6624 (N_6624,N_4264,N_5079);
or U6625 (N_6625,N_3748,N_4307);
nor U6626 (N_6626,N_5994,N_4895);
nor U6627 (N_6627,N_4750,N_3561);
nand U6628 (N_6628,N_3704,N_4331);
and U6629 (N_6629,N_5926,N_5357);
and U6630 (N_6630,N_3245,N_5841);
nor U6631 (N_6631,N_4755,N_5447);
nand U6632 (N_6632,N_4420,N_4127);
nor U6633 (N_6633,N_4882,N_4362);
or U6634 (N_6634,N_4246,N_5620);
or U6635 (N_6635,N_4177,N_3438);
nor U6636 (N_6636,N_3524,N_4910);
nand U6637 (N_6637,N_4668,N_3632);
nor U6638 (N_6638,N_3469,N_5561);
xnor U6639 (N_6639,N_3736,N_4412);
xor U6640 (N_6640,N_5802,N_4119);
nor U6641 (N_6641,N_4891,N_3255);
nand U6642 (N_6642,N_5750,N_5128);
xnor U6643 (N_6643,N_5138,N_5751);
and U6644 (N_6644,N_4846,N_4830);
or U6645 (N_6645,N_5761,N_3916);
or U6646 (N_6646,N_4666,N_4343);
nand U6647 (N_6647,N_4905,N_5592);
and U6648 (N_6648,N_5369,N_4700);
nor U6649 (N_6649,N_3340,N_3357);
nor U6650 (N_6650,N_5531,N_4844);
nor U6651 (N_6651,N_4779,N_4778);
or U6652 (N_6652,N_4991,N_5469);
nand U6653 (N_6653,N_4809,N_5896);
and U6654 (N_6654,N_5741,N_4536);
nand U6655 (N_6655,N_3314,N_4622);
nand U6656 (N_6656,N_5493,N_3354);
or U6657 (N_6657,N_5923,N_3346);
or U6658 (N_6658,N_3419,N_3966);
nor U6659 (N_6659,N_5321,N_5031);
nand U6660 (N_6660,N_5535,N_5467);
nor U6661 (N_6661,N_3234,N_5938);
or U6662 (N_6662,N_3430,N_5480);
nand U6663 (N_6663,N_5697,N_4803);
nor U6664 (N_6664,N_5255,N_5460);
and U6665 (N_6665,N_3037,N_3479);
or U6666 (N_6666,N_3236,N_3446);
or U6667 (N_6667,N_3000,N_3392);
or U6668 (N_6668,N_4477,N_5603);
or U6669 (N_6669,N_4348,N_5801);
or U6670 (N_6670,N_3316,N_3919);
nor U6671 (N_6671,N_4223,N_4531);
xnor U6672 (N_6672,N_5250,N_3003);
and U6673 (N_6673,N_4501,N_4573);
nand U6674 (N_6674,N_4037,N_3936);
nor U6675 (N_6675,N_5454,N_5732);
and U6676 (N_6676,N_4207,N_5164);
xor U6677 (N_6677,N_4732,N_3349);
nor U6678 (N_6678,N_5647,N_5294);
nand U6679 (N_6679,N_4030,N_3128);
and U6680 (N_6680,N_4958,N_4855);
nand U6681 (N_6681,N_3942,N_4414);
nand U6682 (N_6682,N_4785,N_3773);
and U6683 (N_6683,N_4605,N_3439);
nand U6684 (N_6684,N_4649,N_4819);
nor U6685 (N_6685,N_5538,N_5510);
nor U6686 (N_6686,N_5665,N_4474);
nor U6687 (N_6687,N_5765,N_4230);
nor U6688 (N_6688,N_5810,N_3127);
and U6689 (N_6689,N_3545,N_4136);
nand U6690 (N_6690,N_3214,N_5981);
nand U6691 (N_6691,N_4997,N_3157);
and U6692 (N_6692,N_4434,N_3335);
nor U6693 (N_6693,N_3475,N_3155);
and U6694 (N_6694,N_4128,N_3572);
nand U6695 (N_6695,N_5444,N_4692);
nand U6696 (N_6696,N_4686,N_4796);
xor U6697 (N_6697,N_5181,N_3864);
xnor U6698 (N_6698,N_3900,N_5097);
nor U6699 (N_6699,N_5570,N_4288);
nor U6700 (N_6700,N_3820,N_4716);
xnor U6701 (N_6701,N_4507,N_5222);
and U6702 (N_6702,N_3808,N_3056);
and U6703 (N_6703,N_4482,N_4297);
nor U6704 (N_6704,N_4359,N_4112);
nand U6705 (N_6705,N_5960,N_5495);
nor U6706 (N_6706,N_5007,N_5807);
nand U6707 (N_6707,N_3359,N_5268);
nand U6708 (N_6708,N_3867,N_3442);
or U6709 (N_6709,N_5961,N_3338);
xor U6710 (N_6710,N_4800,N_3308);
and U6711 (N_6711,N_5362,N_3990);
nand U6712 (N_6712,N_5240,N_4457);
nor U6713 (N_6713,N_3508,N_3539);
or U6714 (N_6714,N_4954,N_4377);
or U6715 (N_6715,N_5352,N_5589);
or U6716 (N_6716,N_3188,N_5087);
nand U6717 (N_6717,N_3984,N_3763);
and U6718 (N_6718,N_3211,N_5004);
and U6719 (N_6719,N_5927,N_5115);
nor U6720 (N_6720,N_4472,N_5208);
nand U6721 (N_6721,N_5233,N_5308);
nor U6722 (N_6722,N_3735,N_4595);
or U6723 (N_6723,N_4673,N_5721);
nor U6724 (N_6724,N_3591,N_4625);
or U6725 (N_6725,N_4508,N_4956);
xnor U6726 (N_6726,N_3249,N_3230);
or U6727 (N_6727,N_5427,N_4893);
and U6728 (N_6728,N_4795,N_3534);
xnor U6729 (N_6729,N_4940,N_5957);
and U6730 (N_6730,N_3931,N_4104);
nor U6731 (N_6731,N_4632,N_3896);
or U6732 (N_6732,N_3025,N_3974);
or U6733 (N_6733,N_4527,N_4533);
nand U6734 (N_6734,N_4374,N_5658);
nand U6735 (N_6735,N_3264,N_3855);
nand U6736 (N_6736,N_5575,N_4057);
nor U6737 (N_6737,N_5654,N_3741);
or U6738 (N_6738,N_5192,N_5404);
and U6739 (N_6739,N_3269,N_3913);
and U6740 (N_6740,N_3298,N_3148);
and U6741 (N_6741,N_5327,N_4884);
and U6742 (N_6742,N_5384,N_5700);
nor U6743 (N_6743,N_4053,N_3631);
and U6744 (N_6744,N_4409,N_5872);
nand U6745 (N_6745,N_4326,N_5458);
or U6746 (N_6746,N_5248,N_5326);
and U6747 (N_6747,N_4892,N_5410);
and U6748 (N_6748,N_4731,N_4955);
nor U6749 (N_6749,N_5453,N_3399);
nor U6750 (N_6750,N_3947,N_3132);
or U6751 (N_6751,N_5276,N_3202);
or U6752 (N_6752,N_5085,N_5142);
xnor U6753 (N_6753,N_3492,N_3804);
xor U6754 (N_6754,N_5983,N_4781);
nor U6755 (N_6755,N_5177,N_3813);
and U6756 (N_6756,N_5488,N_4236);
nand U6757 (N_6757,N_4184,N_3212);
or U6758 (N_6758,N_3445,N_3989);
nor U6759 (N_6759,N_4304,N_5804);
and U6760 (N_6760,N_3064,N_5227);
nand U6761 (N_6761,N_5738,N_4023);
nor U6762 (N_6762,N_5107,N_4794);
nor U6763 (N_6763,N_3987,N_5722);
or U6764 (N_6764,N_4674,N_3443);
nor U6765 (N_6765,N_4567,N_5088);
or U6766 (N_6766,N_4679,N_3554);
or U6767 (N_6767,N_4013,N_4229);
nor U6768 (N_6768,N_4723,N_4463);
xor U6769 (N_6769,N_5631,N_5569);
or U6770 (N_6770,N_4611,N_4095);
and U6771 (N_6771,N_5232,N_5895);
and U6772 (N_6772,N_3893,N_3252);
or U6773 (N_6773,N_3982,N_4031);
or U6774 (N_6774,N_4086,N_5307);
nand U6775 (N_6775,N_3684,N_5116);
nor U6776 (N_6776,N_5723,N_3416);
and U6777 (N_6777,N_4214,N_3307);
nand U6778 (N_6778,N_4105,N_4237);
nand U6779 (N_6779,N_5355,N_5122);
nand U6780 (N_6780,N_4330,N_5146);
xor U6781 (N_6781,N_3143,N_5282);
nand U6782 (N_6782,N_4005,N_3823);
nor U6783 (N_6783,N_4850,N_5068);
and U6784 (N_6784,N_5821,N_5126);
or U6785 (N_6785,N_4262,N_3777);
xnor U6786 (N_6786,N_5925,N_4302);
nor U6787 (N_6787,N_3200,N_4876);
nand U6788 (N_6788,N_3076,N_5635);
nor U6789 (N_6789,N_3080,N_4339);
nand U6790 (N_6790,N_3953,N_4976);
nor U6791 (N_6791,N_3268,N_3525);
or U6792 (N_6792,N_3066,N_3728);
or U6793 (N_6793,N_5563,N_3929);
or U6794 (N_6794,N_3090,N_3541);
and U6795 (N_6795,N_3814,N_3637);
nand U6796 (N_6796,N_3613,N_3033);
or U6797 (N_6797,N_4233,N_4906);
nor U6798 (N_6798,N_5237,N_4470);
nor U6799 (N_6799,N_4017,N_5471);
or U6800 (N_6800,N_5484,N_5231);
nand U6801 (N_6801,N_3459,N_5846);
or U6802 (N_6802,N_3729,N_3393);
and U6803 (N_6803,N_4267,N_4749);
and U6804 (N_6804,N_5472,N_5279);
xnor U6805 (N_6805,N_3319,N_3022);
xnor U6806 (N_6806,N_3415,N_4783);
or U6807 (N_6807,N_4042,N_3639);
xor U6808 (N_6808,N_3686,N_4467);
nor U6809 (N_6809,N_5038,N_5878);
nand U6810 (N_6810,N_5823,N_3060);
and U6811 (N_6811,N_3996,N_5523);
nor U6812 (N_6812,N_3177,N_4524);
nand U6813 (N_6813,N_3472,N_3619);
and U6814 (N_6814,N_5830,N_5856);
xnor U6815 (N_6815,N_4786,N_3441);
or U6816 (N_6816,N_5770,N_4651);
nand U6817 (N_6817,N_3052,N_3497);
or U6818 (N_6818,N_5505,N_4473);
nand U6819 (N_6819,N_5568,N_3248);
nand U6820 (N_6820,N_5715,N_3362);
and U6821 (N_6821,N_5409,N_3129);
xnor U6822 (N_6822,N_4660,N_5864);
and U6823 (N_6823,N_4904,N_3350);
nor U6824 (N_6824,N_5374,N_4624);
nand U6825 (N_6825,N_4048,N_5990);
or U6826 (N_6826,N_4484,N_3620);
xnor U6827 (N_6827,N_5169,N_3332);
nor U6828 (N_6828,N_3029,N_5207);
or U6829 (N_6829,N_3794,N_4219);
xnor U6830 (N_6830,N_4211,N_3977);
and U6831 (N_6831,N_4714,N_5170);
nand U6832 (N_6832,N_5071,N_4202);
nor U6833 (N_6833,N_3961,N_4151);
xor U6834 (N_6834,N_3852,N_4225);
nand U6835 (N_6835,N_3641,N_5434);
nand U6836 (N_6836,N_3547,N_4056);
and U6837 (N_6837,N_5565,N_5451);
and U6838 (N_6838,N_3669,N_3387);
or U6839 (N_6839,N_5789,N_5888);
or U6840 (N_6840,N_4708,N_5429);
or U6841 (N_6841,N_5629,N_5840);
and U6842 (N_6842,N_4123,N_4016);
nand U6843 (N_6843,N_3124,N_3461);
and U6844 (N_6844,N_3553,N_4342);
nand U6845 (N_6845,N_5571,N_3719);
nor U6846 (N_6846,N_3227,N_3531);
or U6847 (N_6847,N_5390,N_5796);
and U6848 (N_6848,N_3573,N_3700);
nor U6849 (N_6849,N_4231,N_4242);
nand U6850 (N_6850,N_5168,N_4195);
or U6851 (N_6851,N_4141,N_5678);
nor U6852 (N_6852,N_3544,N_3761);
nor U6853 (N_6853,N_4101,N_3506);
and U6854 (N_6854,N_5061,N_5200);
or U6855 (N_6855,N_4178,N_4059);
nand U6856 (N_6856,N_4003,N_3785);
nor U6857 (N_6857,N_3154,N_5999);
and U6858 (N_6858,N_5340,N_3681);
nand U6859 (N_6859,N_3096,N_5015);
and U6860 (N_6860,N_4106,N_4318);
nor U6861 (N_6861,N_4709,N_4181);
nand U6862 (N_6862,N_4722,N_5130);
or U6863 (N_6863,N_4273,N_5969);
nor U6864 (N_6864,N_5696,N_4073);
or U6865 (N_6865,N_5431,N_3690);
or U6866 (N_6866,N_3208,N_4967);
and U6867 (N_6867,N_5067,N_3699);
nor U6868 (N_6868,N_3689,N_3895);
nand U6869 (N_6869,N_5526,N_5273);
nor U6870 (N_6870,N_3069,N_5945);
and U6871 (N_6871,N_5934,N_5986);
and U6872 (N_6872,N_4925,N_3197);
and U6873 (N_6873,N_3280,N_4650);
and U6874 (N_6874,N_3050,N_4621);
nor U6875 (N_6875,N_5940,N_3787);
or U6876 (N_6876,N_3016,N_5455);
and U6877 (N_6877,N_5869,N_4129);
or U6878 (N_6878,N_4571,N_4064);
or U6879 (N_6879,N_3955,N_5987);
xor U6880 (N_6880,N_3244,N_3193);
and U6881 (N_6881,N_5049,N_4118);
or U6882 (N_6882,N_5285,N_4460);
and U6883 (N_6883,N_5385,N_3711);
or U6884 (N_6884,N_4972,N_4740);
or U6885 (N_6885,N_5704,N_3726);
nor U6886 (N_6886,N_3903,N_5714);
or U6887 (N_6887,N_4109,N_5408);
nor U6888 (N_6888,N_5868,N_5932);
nor U6889 (N_6889,N_5924,N_5837);
or U6890 (N_6890,N_4838,N_4115);
nand U6891 (N_6891,N_5877,N_3452);
xor U6892 (N_6892,N_4388,N_5689);
nand U6893 (N_6893,N_5546,N_3598);
nand U6894 (N_6894,N_5437,N_3274);
nor U6895 (N_6895,N_3071,N_5683);
nor U6896 (N_6896,N_3036,N_5400);
or U6897 (N_6897,N_4490,N_3537);
nor U6898 (N_6898,N_4071,N_4813);
nand U6899 (N_6899,N_3832,N_3151);
or U6900 (N_6900,N_3238,N_3579);
xnor U6901 (N_6901,N_3434,N_3958);
or U6902 (N_6902,N_3231,N_4957);
and U6903 (N_6903,N_4188,N_4560);
nand U6904 (N_6904,N_5997,N_3605);
nand U6905 (N_6905,N_4861,N_5463);
or U6906 (N_6906,N_4873,N_5659);
nor U6907 (N_6907,N_5857,N_3830);
and U6908 (N_6908,N_3667,N_4627);
nand U6909 (N_6909,N_3590,N_5098);
nand U6910 (N_6910,N_3944,N_3829);
nand U6911 (N_6911,N_3724,N_4772);
xnor U6912 (N_6912,N_5003,N_3782);
nand U6913 (N_6913,N_3652,N_5461);
and U6914 (N_6914,N_4455,N_4186);
and U6915 (N_6915,N_5347,N_5843);
nand U6916 (N_6916,N_3108,N_4848);
and U6917 (N_6917,N_4811,N_5847);
nand U6918 (N_6918,N_5903,N_3580);
and U6919 (N_6919,N_4036,N_3768);
and U6920 (N_6920,N_3876,N_3051);
nor U6921 (N_6921,N_5703,N_4196);
nor U6922 (N_6922,N_3169,N_3610);
nor U6923 (N_6923,N_5892,N_5712);
nand U6924 (N_6924,N_5978,N_5176);
and U6925 (N_6925,N_4646,N_5055);
and U6926 (N_6926,N_3950,N_3612);
nand U6927 (N_6927,N_5512,N_5334);
or U6928 (N_6928,N_3026,N_4468);
or U6929 (N_6929,N_3424,N_5547);
nor U6930 (N_6930,N_4695,N_5236);
xnor U6931 (N_6931,N_3386,N_4398);
or U6932 (N_6932,N_5836,N_3812);
nor U6933 (N_6933,N_5290,N_3464);
xnor U6934 (N_6934,N_4263,N_3358);
or U6935 (N_6935,N_4275,N_5433);
or U6936 (N_6936,N_3187,N_3588);
xnor U6937 (N_6937,N_3189,N_5785);
or U6938 (N_6938,N_4509,N_3370);
nor U6939 (N_6939,N_3512,N_4114);
nand U6940 (N_6940,N_5503,N_4191);
nand U6941 (N_6941,N_4189,N_3586);
xnor U6942 (N_6942,N_4885,N_3904);
or U6943 (N_6943,N_5147,N_3196);
nor U6944 (N_6944,N_4075,N_4345);
nand U6945 (N_6945,N_5280,N_5064);
xor U6946 (N_6946,N_5891,N_4183);
and U6947 (N_6947,N_3039,N_5601);
nand U6948 (N_6948,N_5375,N_5968);
nor U6949 (N_6949,N_5359,N_4578);
and U6950 (N_6950,N_3113,N_3405);
or U6951 (N_6951,N_3055,N_3334);
or U6952 (N_6952,N_4050,N_5016);
nand U6953 (N_6953,N_4548,N_5043);
or U6954 (N_6954,N_3713,N_4769);
or U6955 (N_6955,N_5939,N_3878);
nand U6956 (N_6956,N_4667,N_4358);
or U6957 (N_6957,N_4845,N_4889);
or U6958 (N_6958,N_3800,N_5587);
or U6959 (N_6959,N_4492,N_3651);
and U6960 (N_6960,N_3529,N_5643);
or U6961 (N_6961,N_3860,N_5081);
and U6962 (N_6962,N_4287,N_5728);
nand U6963 (N_6963,N_5494,N_5141);
nor U6964 (N_6964,N_3760,N_5636);
nor U6965 (N_6965,N_4355,N_5193);
nand U6966 (N_6966,N_3658,N_3807);
nand U6967 (N_6967,N_3477,N_3635);
nand U6968 (N_6968,N_5499,N_3869);
nand U6969 (N_6969,N_3519,N_5011);
nor U6970 (N_6970,N_3642,N_4068);
and U6971 (N_6971,N_4144,N_5564);
and U6972 (N_6972,N_5099,N_4890);
or U6973 (N_6973,N_4270,N_4383);
and U6974 (N_6974,N_4761,N_4771);
nand U6975 (N_6975,N_3271,N_4659);
nor U6976 (N_6976,N_4619,N_4080);
or U6977 (N_6977,N_4117,N_3756);
nor U6978 (N_6978,N_3382,N_5476);
or U6979 (N_6979,N_4133,N_4311);
and U6980 (N_6980,N_5199,N_4901);
or U6981 (N_6981,N_5032,N_5303);
or U6982 (N_6982,N_4171,N_3948);
nor U6983 (N_6983,N_3673,N_3250);
nand U6984 (N_6984,N_3680,N_4915);
or U6985 (N_6985,N_4914,N_3615);
and U6986 (N_6986,N_3150,N_5500);
nor U6987 (N_6987,N_5440,N_5915);
xor U6988 (N_6988,N_4166,N_3368);
nor U6989 (N_6989,N_5052,N_4523);
nor U6990 (N_6990,N_4019,N_5171);
xnor U6991 (N_6991,N_4168,N_5534);
or U6992 (N_6992,N_3398,N_4090);
nand U6993 (N_6993,N_5238,N_4285);
and U6994 (N_6994,N_4875,N_4462);
nor U6995 (N_6995,N_3691,N_5776);
nand U6996 (N_6996,N_5124,N_4831);
nand U6997 (N_6997,N_5253,N_3753);
or U6998 (N_6998,N_4002,N_4768);
or U6999 (N_6999,N_3546,N_3725);
and U7000 (N_7000,N_5874,N_4847);
nor U7001 (N_7001,N_3226,N_4594);
xor U7002 (N_7002,N_3797,N_5370);
or U7003 (N_7003,N_5555,N_3999);
nor U7004 (N_7004,N_3198,N_3118);
xnor U7005 (N_7005,N_4419,N_3560);
nor U7006 (N_7006,N_4887,N_4198);
nand U7007 (N_7007,N_4654,N_3884);
and U7008 (N_7008,N_5859,N_4145);
or U7009 (N_7009,N_5566,N_5560);
nand U7010 (N_7010,N_5183,N_3375);
nand U7011 (N_7011,N_3318,N_5215);
nand U7012 (N_7012,N_4083,N_4097);
and U7013 (N_7013,N_5820,N_4179);
or U7014 (N_7014,N_3928,N_3086);
nor U7015 (N_7015,N_4613,N_4877);
nor U7016 (N_7016,N_5368,N_5325);
nor U7017 (N_7017,N_3789,N_3514);
nand U7018 (N_7018,N_3299,N_3489);
and U7019 (N_7019,N_5485,N_4648);
nand U7020 (N_7020,N_3180,N_5744);
nor U7021 (N_7021,N_4661,N_5042);
nand U7022 (N_7022,N_3352,N_4029);
xnor U7023 (N_7023,N_4004,N_5309);
nand U7024 (N_7024,N_5318,N_5167);
nand U7025 (N_7025,N_3734,N_4421);
and U7026 (N_7026,N_4295,N_5112);
and U7027 (N_7027,N_3300,N_3576);
nand U7028 (N_7028,N_4992,N_5351);
xnor U7029 (N_7029,N_5103,N_5198);
nand U7030 (N_7030,N_3110,N_3503);
xor U7031 (N_7031,N_4274,N_5100);
and U7032 (N_7032,N_4606,N_5391);
and U7033 (N_7033,N_4137,N_5688);
or U7034 (N_7034,N_4060,N_3784);
or U7035 (N_7035,N_5402,N_3282);
nand U7036 (N_7036,N_3331,N_4818);
nand U7037 (N_7037,N_3216,N_4170);
nand U7038 (N_7038,N_4190,N_3701);
nand U7039 (N_7039,N_5462,N_5539);
or U7040 (N_7040,N_3218,N_4928);
or U7041 (N_7041,N_4747,N_5005);
nand U7042 (N_7042,N_3834,N_5622);
nand U7043 (N_7043,N_4897,N_3351);
or U7044 (N_7044,N_3670,N_5540);
nand U7045 (N_7045,N_3082,N_5379);
nand U7046 (N_7046,N_3975,N_4130);
nor U7047 (N_7047,N_5815,N_3041);
nor U7048 (N_7048,N_4717,N_4909);
and U7049 (N_7049,N_5354,N_4574);
or U7050 (N_7050,N_5261,N_5763);
and U7051 (N_7051,N_5879,N_3888);
and U7052 (N_7052,N_5228,N_5466);
and U7053 (N_7053,N_4107,N_3671);
nor U7054 (N_7054,N_5731,N_5266);
or U7055 (N_7055,N_5014,N_4041);
nor U7056 (N_7056,N_5223,N_3663);
nand U7057 (N_7057,N_3809,N_4024);
nor U7058 (N_7058,N_4007,N_4683);
nand U7059 (N_7059,N_4309,N_4635);
nor U7060 (N_7060,N_4430,N_3418);
and U7061 (N_7061,N_5779,N_3134);
or U7062 (N_7062,N_3574,N_5474);
and U7063 (N_7063,N_4612,N_5518);
nor U7064 (N_7064,N_3044,N_3256);
nor U7065 (N_7065,N_3400,N_5278);
nand U7066 (N_7066,N_5797,N_4200);
nand U7067 (N_7067,N_3722,N_5735);
xnor U7068 (N_7068,N_4475,N_5428);
or U7069 (N_7069,N_5913,N_5132);
nand U7070 (N_7070,N_3242,N_4935);
nor U7071 (N_7071,N_5025,N_3709);
and U7072 (N_7072,N_3562,N_3527);
and U7073 (N_7073,N_5258,N_4519);
nand U7074 (N_7074,N_5677,N_5614);
xnor U7075 (N_7075,N_5486,N_3361);
or U7076 (N_7076,N_5976,N_3363);
or U7077 (N_7077,N_4373,N_5889);
nor U7078 (N_7078,N_4681,N_3130);
or U7079 (N_7079,N_4643,N_4389);
or U7080 (N_7080,N_3083,N_5018);
nor U7081 (N_7081,N_5794,N_4765);
or U7082 (N_7082,N_3453,N_4459);
nor U7083 (N_7083,N_4705,N_5724);
and U7084 (N_7084,N_5955,N_4451);
and U7085 (N_7085,N_4902,N_3960);
and U7086 (N_7086,N_4977,N_4428);
xor U7087 (N_7087,N_3061,N_3136);
nand U7088 (N_7088,N_3140,N_5627);
nand U7089 (N_7089,N_4126,N_4664);
or U7090 (N_7090,N_3664,N_3934);
nor U7091 (N_7091,N_3644,N_5755);
xnor U7092 (N_7092,N_5411,N_4577);
nor U7093 (N_7093,N_5772,N_4912);
and U7094 (N_7094,N_3767,N_3805);
or U7095 (N_7095,N_5740,N_5348);
or U7096 (N_7096,N_4900,N_4563);
and U7097 (N_7097,N_3407,N_3870);
nand U7098 (N_7098,N_4043,N_3454);
nand U7099 (N_7099,N_5398,N_5867);
nor U7100 (N_7100,N_4944,N_4591);
and U7101 (N_7101,N_5730,N_3355);
and U7102 (N_7102,N_5235,N_3795);
or U7103 (N_7103,N_4983,N_4169);
xnor U7104 (N_7104,N_4554,N_4685);
xnor U7105 (N_7105,N_5481,N_4792);
or U7106 (N_7106,N_5612,N_5759);
or U7107 (N_7107,N_5302,N_4546);
and U7108 (N_7108,N_3976,N_5501);
nor U7109 (N_7109,N_5366,N_4496);
nand U7110 (N_7110,N_5062,N_3032);
nand U7111 (N_7111,N_3880,N_3617);
nor U7112 (N_7112,N_3751,N_5577);
xor U7113 (N_7113,N_3945,N_5075);
or U7114 (N_7114,N_5436,N_3185);
or U7115 (N_7115,N_3740,N_5784);
nor U7116 (N_7116,N_3232,N_3432);
or U7117 (N_7117,N_4187,N_4729);
xnor U7118 (N_7118,N_3491,N_5378);
or U7119 (N_7119,N_4559,N_5553);
nor U7120 (N_7120,N_3394,N_4238);
and U7121 (N_7121,N_3224,N_4908);
and U7122 (N_7122,N_4989,N_4425);
or U7123 (N_7123,N_5021,N_3771);
or U7124 (N_7124,N_3018,N_4103);
or U7125 (N_7125,N_5967,N_3717);
or U7126 (N_7126,N_4266,N_3057);
nand U7127 (N_7127,N_5749,N_4728);
nand U7128 (N_7128,N_5616,N_4789);
or U7129 (N_7129,N_3843,N_4953);
nand U7130 (N_7130,N_3336,N_3295);
and U7131 (N_7131,N_3063,N_4710);
nor U7132 (N_7132,N_4480,N_5080);
nor U7133 (N_7133,N_3603,N_5046);
nor U7134 (N_7134,N_3788,N_5330);
xor U7135 (N_7135,N_3755,N_3857);
nor U7136 (N_7136,N_5550,N_4510);
xnor U7137 (N_7137,N_4840,N_3201);
or U7138 (N_7138,N_4557,N_4255);
nand U7139 (N_7139,N_3278,N_3220);
or U7140 (N_7140,N_3730,N_3847);
nor U7141 (N_7141,N_4399,N_3440);
nand U7142 (N_7142,N_3507,N_3634);
xor U7143 (N_7143,N_3705,N_3168);
and U7144 (N_7144,N_4489,N_5953);
and U7145 (N_7145,N_5220,N_3890);
or U7146 (N_7146,N_3747,N_3463);
nor U7147 (N_7147,N_4054,N_3466);
nor U7148 (N_7148,N_5039,N_3879);
nand U7149 (N_7149,N_3421,N_5970);
or U7150 (N_7150,N_3938,N_4862);
and U7151 (N_7151,N_3364,N_3254);
nand U7152 (N_7152,N_3520,N_3207);
nor U7153 (N_7153,N_3624,N_3532);
nor U7154 (N_7154,N_4038,N_3502);
nand U7155 (N_7155,N_5844,N_5762);
or U7156 (N_7156,N_5543,N_5182);
and U7157 (N_7157,N_3694,N_4045);
or U7158 (N_7158,N_4655,N_5634);
and U7159 (N_7159,N_4566,N_4774);
and U7160 (N_7160,N_3932,N_5922);
nand U7161 (N_7161,N_3819,N_4491);
and U7162 (N_7162,N_4529,N_3068);
and U7163 (N_7163,N_5800,N_5275);
nand U7164 (N_7164,N_3437,N_3243);
and U7165 (N_7165,N_5912,N_4116);
or U7166 (N_7166,N_4157,N_5377);
and U7167 (N_7167,N_3170,N_4395);
nand U7168 (N_7168,N_4824,N_4111);
xor U7169 (N_7169,N_5699,N_5655);
nand U7170 (N_7170,N_5050,N_4371);
or U7171 (N_7171,N_5805,N_5111);
nor U7172 (N_7172,N_3744,N_4344);
nand U7173 (N_7173,N_4069,N_3774);
nand U7174 (N_7174,N_4321,N_5929);
or U7175 (N_7175,N_4759,N_3696);
or U7176 (N_7176,N_3521,N_5127);
nor U7177 (N_7177,N_3672,N_3178);
nand U7178 (N_7178,N_3803,N_5617);
nor U7179 (N_7179,N_3584,N_3985);
or U7180 (N_7180,N_5707,N_5992);
or U7181 (N_7181,N_5792,N_5381);
or U7182 (N_7182,N_3409,N_5178);
nor U7183 (N_7183,N_3565,N_5608);
nand U7184 (N_7184,N_5504,N_4224);
or U7185 (N_7185,N_4327,N_4212);
nor U7186 (N_7186,N_5729,N_3951);
xnor U7187 (N_7187,N_4099,N_3716);
nor U7188 (N_7188,N_4363,N_3171);
xnor U7189 (N_7189,N_5218,N_5736);
and U7190 (N_7190,N_4880,N_5477);
nand U7191 (N_7191,N_3594,N_4260);
and U7192 (N_7192,N_3923,N_3970);
and U7193 (N_7193,N_4182,N_5102);
or U7194 (N_7194,N_5593,N_4483);
nand U7195 (N_7195,N_4962,N_5166);
nand U7196 (N_7196,N_5962,N_4996);
or U7197 (N_7197,N_4404,N_5842);
and U7198 (N_7198,N_4325,N_4386);
nand U7199 (N_7199,N_3836,N_4926);
and U7200 (N_7200,N_5091,N_4481);
and U7201 (N_7201,N_5483,N_3874);
nor U7202 (N_7202,N_3457,N_4770);
and U7203 (N_7203,N_3204,N_5536);
and U7204 (N_7204,N_5175,N_4706);
and U7205 (N_7205,N_5692,N_4160);
nor U7206 (N_7206,N_4721,N_5241);
nor U7207 (N_7207,N_3685,N_5213);
nor U7208 (N_7208,N_5204,N_5158);
nor U7209 (N_7209,N_3389,N_4180);
nor U7210 (N_7210,N_4570,N_4221);
nor U7211 (N_7211,N_4592,N_4978);
nand U7212 (N_7212,N_4213,N_5833);
nor U7213 (N_7213,N_3972,N_4239);
or U7214 (N_7214,N_5742,N_4671);
and U7215 (N_7215,N_3540,N_5851);
xor U7216 (N_7216,N_3778,N_5076);
nand U7217 (N_7217,N_4265,N_4979);
nand U7218 (N_7218,N_4593,N_4637);
nand U7219 (N_7219,N_4517,N_5698);
nor U7220 (N_7220,N_3854,N_5372);
and U7221 (N_7221,N_3257,N_5363);
nand U7222 (N_7222,N_4665,N_5188);
and U7223 (N_7223,N_4098,N_5392);
nor U7224 (N_7224,N_5020,N_3100);
nor U7225 (N_7225,N_5424,N_5211);
or U7226 (N_7226,N_4149,N_5900);
nand U7227 (N_7227,N_4841,N_4513);
nand U7228 (N_7228,N_3404,N_3315);
and U7229 (N_7229,N_3675,N_4452);
and U7230 (N_7230,N_4254,N_5201);
or U7231 (N_7231,N_4810,N_5600);
or U7232 (N_7232,N_5313,N_4947);
or U7233 (N_7233,N_3104,N_5311);
and U7234 (N_7234,N_4065,N_4296);
nand U7235 (N_7235,N_5040,N_5835);
nand U7236 (N_7236,N_3552,N_3088);
and U7237 (N_7237,N_3638,N_3210);
or U7238 (N_7238,N_5583,N_3759);
nor U7239 (N_7239,N_4825,N_5582);
nor U7240 (N_7240,N_4299,N_5975);
or U7241 (N_7241,N_4055,N_5717);
nor U7242 (N_7242,N_4663,N_4687);
nand U7243 (N_7243,N_3049,N_4332);
and U7244 (N_7244,N_4251,N_4970);
and U7245 (N_7245,N_3898,N_4782);
and U7246 (N_7246,N_5301,N_3144);
or U7247 (N_7247,N_3558,N_4417);
nor U7248 (N_7248,N_5487,N_3383);
nand U7249 (N_7249,N_3078,N_5406);
and U7250 (N_7250,N_3395,N_3240);
and U7251 (N_7251,N_4597,N_4310);
xor U7252 (N_7252,N_4806,N_5350);
nand U7253 (N_7253,N_3137,N_4688);
and U7254 (N_7254,N_5982,N_4461);
xnor U7255 (N_7255,N_4469,N_5748);
nor U7256 (N_7256,N_5246,N_5720);
and U7257 (N_7257,N_4305,N_5666);
nor U7258 (N_7258,N_3742,N_4150);
and U7259 (N_7259,N_4561,N_5412);
xor U7260 (N_7260,N_5530,N_4286);
and U7261 (N_7261,N_3106,N_3107);
nand U7262 (N_7262,N_4503,N_3482);
or U7263 (N_7263,N_5281,N_3837);
nand U7264 (N_7264,N_5296,N_3377);
or U7265 (N_7265,N_3146,N_4851);
xnor U7266 (N_7266,N_5507,N_5649);
or U7267 (N_7267,N_3569,N_3839);
or U7268 (N_7268,N_3886,N_4077);
and U7269 (N_7269,N_3824,N_4584);
or U7270 (N_7270,N_3109,N_3451);
and U7271 (N_7271,N_4040,N_3831);
or U7272 (N_7272,N_5774,N_4843);
and U7273 (N_7273,N_3668,N_4308);
nand U7274 (N_7274,N_3481,N_5328);
or U7275 (N_7275,N_3054,N_4623);
nor U7276 (N_7276,N_4122,N_3251);
nand U7277 (N_7277,N_5136,N_5148);
or U7278 (N_7278,N_4866,N_5902);
nor U7279 (N_7279,N_3861,N_3101);
and U7280 (N_7280,N_4512,N_3112);
and U7281 (N_7281,N_4773,N_3563);
or U7282 (N_7282,N_4867,N_4812);
or U7283 (N_7283,N_3191,N_5274);
xor U7284 (N_7284,N_3618,N_3827);
or U7285 (N_7285,N_5026,N_5160);
nor U7286 (N_7286,N_3633,N_3223);
nand U7287 (N_7287,N_4336,N_3079);
and U7288 (N_7288,N_5542,N_5361);
or U7289 (N_7289,N_3653,N_3602);
nand U7290 (N_7290,N_3038,N_5936);
nor U7291 (N_7291,N_3084,N_3367);
and U7292 (N_7292,N_3687,N_3283);
nor U7293 (N_7293,N_3046,N_5813);
xor U7294 (N_7294,N_3302,N_5725);
nor U7295 (N_7295,N_5047,N_4319);
nor U7296 (N_7296,N_3891,N_4406);
nand U7297 (N_7297,N_4173,N_5419);
and U7298 (N_7298,N_4256,N_3496);
nand U7299 (N_7299,N_5058,N_4400);
or U7300 (N_7300,N_4058,N_5899);
or U7301 (N_7301,N_4340,N_3792);
and U7302 (N_7302,N_4924,N_4985);
xnor U7303 (N_7303,N_4964,N_4009);
xnor U7304 (N_7304,N_4864,N_5153);
nor U7305 (N_7305,N_3596,N_4966);
or U7306 (N_7306,N_3027,N_5854);
xor U7307 (N_7307,N_5694,N_5413);
nor U7308 (N_7308,N_3801,N_3600);
nor U7309 (N_7309,N_5808,N_3072);
and U7310 (N_7310,N_5596,N_4822);
nand U7311 (N_7311,N_4502,N_4715);
and U7312 (N_7312,N_3379,N_5060);
and U7313 (N_7313,N_4372,N_3581);
or U7314 (N_7314,N_3480,N_5845);
and U7315 (N_7315,N_4739,N_3592);
nand U7316 (N_7316,N_4092,N_4791);
nor U7317 (N_7317,N_5893,N_4120);
or U7318 (N_7318,N_5205,N_5123);
nand U7319 (N_7319,N_5387,N_3627);
nor U7320 (N_7320,N_4698,N_3780);
nand U7321 (N_7321,N_3406,N_4155);
and U7322 (N_7322,N_5826,N_3262);
or U7323 (N_7323,N_3649,N_5650);
and U7324 (N_7324,N_5954,N_5109);
nand U7325 (N_7325,N_5928,N_4397);
xnor U7326 (N_7326,N_5196,N_4078);
or U7327 (N_7327,N_3401,N_3277);
and U7328 (N_7328,N_4014,N_5690);
or U7329 (N_7329,N_3865,N_5885);
and U7330 (N_7330,N_3253,N_5162);
and U7331 (N_7331,N_4939,N_5959);
and U7332 (N_7332,N_4354,N_4121);
nor U7333 (N_7333,N_5401,N_4547);
nor U7334 (N_7334,N_3578,N_5113);
xor U7335 (N_7335,N_3008,N_3528);
nor U7336 (N_7336,N_3286,N_3374);
nand U7337 (N_7337,N_3303,N_4370);
or U7338 (N_7338,N_4532,N_5819);
nor U7339 (N_7339,N_3165,N_5993);
and U7340 (N_7340,N_5734,N_5930);
or U7341 (N_7341,N_5771,N_5894);
nor U7342 (N_7342,N_4918,N_3566);
xnor U7343 (N_7343,N_3645,N_3790);
nand U7344 (N_7344,N_4464,N_5871);
and U7345 (N_7345,N_4034,N_4543);
nor U7346 (N_7346,N_4883,N_3001);
nand U7347 (N_7347,N_4995,N_5702);
nand U7348 (N_7348,N_4948,N_4220);
and U7349 (N_7349,N_3611,N_3372);
nand U7350 (N_7350,N_4163,N_3474);
or U7351 (N_7351,N_4283,N_4435);
xnor U7352 (N_7352,N_4682,N_3239);
xnor U7353 (N_7353,N_5262,N_3881);
and U7354 (N_7354,N_4742,N_4076);
nand U7355 (N_7355,N_4788,N_5010);
xnor U7356 (N_7356,N_3125,N_3922);
nor U7357 (N_7357,N_4443,N_3209);
nand U7358 (N_7358,N_4874,N_5795);
nand U7359 (N_7359,N_3115,N_3313);
or U7360 (N_7360,N_5701,N_4154);
and U7361 (N_7361,N_5972,N_5602);
and U7362 (N_7362,N_5862,N_3523);
and U7363 (N_7363,N_3825,N_5681);
and U7364 (N_7364,N_3310,N_5257);
nor U7365 (N_7365,N_5615,N_5077);
xor U7366 (N_7366,N_3116,N_3094);
xor U7367 (N_7367,N_3587,N_5435);
or U7368 (N_7368,N_5931,N_3275);
and U7369 (N_7369,N_4576,N_3292);
nand U7370 (N_7370,N_4135,N_5573);
or U7371 (N_7371,N_3786,N_3020);
and U7372 (N_7372,N_4277,N_4172);
or U7373 (N_7373,N_3435,N_5671);
and U7374 (N_7374,N_5284,N_4498);
and U7375 (N_7375,N_5306,N_3164);
nor U7376 (N_7376,N_5640,N_4530);
or U7377 (N_7377,N_4814,N_4752);
xnor U7378 (N_7378,N_5230,N_4730);
nor U7379 (N_7379,N_5610,N_3488);
and U7380 (N_7380,N_3093,N_5979);
nor U7381 (N_7381,N_3583,N_3167);
nor U7382 (N_7382,N_5349,N_5832);
nor U7383 (N_7383,N_3333,N_5174);
nor U7384 (N_7384,N_5827,N_3567);
or U7385 (N_7385,N_5054,N_4079);
and U7386 (N_7386,N_5336,N_4871);
nor U7387 (N_7387,N_4829,N_4369);
nand U7388 (N_7388,N_5644,N_4641);
or U7389 (N_7389,N_3105,N_4444);
nand U7390 (N_7390,N_3577,N_3414);
and U7391 (N_7391,N_4241,N_4733);
nand U7392 (N_7392,N_3659,N_3844);
nand U7393 (N_7393,N_4243,N_5070);
and U7394 (N_7394,N_5244,N_3089);
or U7395 (N_7395,N_3487,N_3897);
and U7396 (N_7396,N_5267,N_3149);
nor U7397 (N_7397,N_4798,N_5298);
nor U7398 (N_7398,N_4675,N_5920);
nor U7399 (N_7399,N_4306,N_4522);
nand U7400 (N_7400,N_3184,N_3894);
nor U7401 (N_7401,N_3657,N_5337);
or U7402 (N_7402,N_5356,N_4707);
nand U7403 (N_7403,N_3940,N_5548);
or U7404 (N_7404,N_3626,N_3866);
and U7405 (N_7405,N_3444,N_5660);
or U7406 (N_7406,N_4379,N_4161);
nor U7407 (N_7407,N_3838,N_4817);
and U7408 (N_7408,N_5269,N_5082);
or U7409 (N_7409,N_3971,N_4589);
nor U7410 (N_7410,N_3766,N_5092);
nand U7411 (N_7411,N_3111,N_5346);
nand U7412 (N_7412,N_4441,N_5152);
and U7413 (N_7413,N_3499,N_4537);
nand U7414 (N_7414,N_3312,N_5456);
xor U7415 (N_7415,N_3205,N_4346);
nand U7416 (N_7416,N_5515,N_5464);
or U7417 (N_7417,N_3412,N_3215);
or U7418 (N_7418,N_5803,N_4618);
nor U7419 (N_7419,N_5478,N_5554);
nor U7420 (N_7420,N_5151,N_5623);
or U7421 (N_7421,N_4091,N_4368);
or U7422 (N_7422,N_3899,N_5586);
nand U7423 (N_7423,N_5948,N_5423);
or U7424 (N_7424,N_4093,N_3012);
nand U7425 (N_7425,N_4982,N_3678);
nand U7426 (N_7426,N_3883,N_3917);
or U7427 (N_7427,N_5562,N_4415);
nor U7428 (N_7428,N_3456,N_3959);
nand U7429 (N_7429,N_3889,N_3420);
xnor U7430 (N_7430,N_4777,N_4699);
nor U7431 (N_7431,N_5909,N_5711);
nand U7432 (N_7432,N_5331,N_3762);
xor U7433 (N_7433,N_3417,N_5528);
and U7434 (N_7434,N_3703,N_5663);
or U7435 (N_7435,N_4582,N_3103);
nor U7436 (N_7436,N_5051,N_5263);
nand U7437 (N_7437,N_5094,N_3770);
and U7438 (N_7438,N_3462,N_4807);
xor U7439 (N_7439,N_3413,N_3595);
and U7440 (N_7440,N_4534,N_5661);
and U7441 (N_7441,N_5682,N_5937);
nor U7442 (N_7442,N_4088,N_4746);
and U7443 (N_7443,N_3344,N_3403);
xor U7444 (N_7444,N_5747,N_5607);
nand U7445 (N_7445,N_5093,N_3848);
nor U7446 (N_7446,N_3995,N_5074);
nor U7447 (N_7447,N_3114,N_4000);
nand U7448 (N_7448,N_4518,N_5468);
xnor U7449 (N_7449,N_5788,N_4932);
or U7450 (N_7450,N_5709,N_3599);
and U7451 (N_7451,N_5059,N_4228);
nor U7452 (N_7452,N_3166,N_3276);
and U7453 (N_7453,N_5773,N_4638);
and U7454 (N_7454,N_4828,N_5686);
nand U7455 (N_7455,N_4197,N_5790);
or U7456 (N_7456,N_4067,N_4201);
and U7457 (N_7457,N_5104,N_4392);
nor U7458 (N_7458,N_3905,N_3289);
or U7459 (N_7459,N_4711,N_4440);
xnor U7460 (N_7460,N_5897,N_5482);
nor U7461 (N_7461,N_3428,N_4620);
and U7462 (N_7462,N_4209,N_3181);
and U7463 (N_7463,N_4044,N_3182);
nand U7464 (N_7464,N_5632,N_3892);
nor U7465 (N_7465,N_4550,N_5745);
nand U7466 (N_7466,N_5191,N_5063);
xor U7467 (N_7467,N_5624,N_4222);
nand U7468 (N_7468,N_3410,N_3450);
and U7469 (N_7469,N_3911,N_3092);
nand U7470 (N_7470,N_5865,N_3517);
or U7471 (N_7471,N_4853,N_3943);
xnor U7472 (N_7472,N_5584,N_5626);
nor U7473 (N_7473,N_3476,N_4353);
or U7474 (N_7474,N_5882,N_5137);
or U7475 (N_7475,N_4269,N_4521);
nand U7476 (N_7476,N_4946,N_3133);
or U7477 (N_7477,N_4364,N_4986);
nand U7478 (N_7478,N_3863,N_4494);
and U7479 (N_7479,N_5108,N_5053);
nand U7480 (N_7480,N_4994,N_5758);
and U7481 (N_7481,N_4232,N_5545);
nand U7482 (N_7482,N_4271,N_4701);
or U7483 (N_7483,N_3575,N_4726);
and U7484 (N_7484,N_4361,N_5664);
or U7485 (N_7485,N_3433,N_3062);
and U7486 (N_7486,N_4974,N_5834);
nor U7487 (N_7487,N_5421,N_5780);
nand U7488 (N_7488,N_5225,N_4969);
and U7489 (N_7489,N_3968,N_4927);
nand U7490 (N_7490,N_5693,N_4402);
nand U7491 (N_7491,N_4138,N_4879);
and U7492 (N_7492,N_3660,N_5254);
nand U7493 (N_7493,N_5809,N_5291);
or U7494 (N_7494,N_3616,N_4987);
or U7495 (N_7495,N_4165,N_3952);
xnor U7496 (N_7496,N_4335,N_3297);
or U7497 (N_7497,N_4754,N_5446);
and U7498 (N_7498,N_4139,N_5866);
xnor U7499 (N_7499,N_5009,N_3246);
or U7500 (N_7500,N_3733,N_3963);
nand U7501 (N_7501,N_4241,N_3096);
nor U7502 (N_7502,N_5953,N_4795);
and U7503 (N_7503,N_3331,N_5860);
or U7504 (N_7504,N_4094,N_5802);
and U7505 (N_7505,N_3181,N_5382);
and U7506 (N_7506,N_5646,N_4192);
nor U7507 (N_7507,N_5334,N_4327);
and U7508 (N_7508,N_5776,N_5872);
nor U7509 (N_7509,N_5596,N_5552);
and U7510 (N_7510,N_3268,N_4595);
or U7511 (N_7511,N_4876,N_5304);
nor U7512 (N_7512,N_4444,N_3064);
nand U7513 (N_7513,N_5439,N_3569);
or U7514 (N_7514,N_5062,N_4078);
and U7515 (N_7515,N_5206,N_4180);
xor U7516 (N_7516,N_5937,N_5144);
nand U7517 (N_7517,N_4505,N_4946);
or U7518 (N_7518,N_3390,N_3815);
or U7519 (N_7519,N_4059,N_5519);
or U7520 (N_7520,N_4955,N_5408);
nand U7521 (N_7521,N_4117,N_4016);
nor U7522 (N_7522,N_4014,N_4510);
or U7523 (N_7523,N_5206,N_3561);
nand U7524 (N_7524,N_4902,N_4559);
xnor U7525 (N_7525,N_3310,N_4594);
nor U7526 (N_7526,N_4996,N_5759);
nor U7527 (N_7527,N_5189,N_5359);
nor U7528 (N_7528,N_4425,N_4619);
nor U7529 (N_7529,N_5214,N_5282);
xnor U7530 (N_7530,N_3390,N_5889);
or U7531 (N_7531,N_3754,N_4818);
and U7532 (N_7532,N_3573,N_4131);
nand U7533 (N_7533,N_5669,N_5063);
nor U7534 (N_7534,N_3560,N_4623);
nor U7535 (N_7535,N_4707,N_3797);
and U7536 (N_7536,N_3539,N_3567);
and U7537 (N_7537,N_3587,N_4169);
nand U7538 (N_7538,N_5774,N_4947);
xor U7539 (N_7539,N_3869,N_4861);
and U7540 (N_7540,N_4737,N_5215);
nand U7541 (N_7541,N_3455,N_5923);
nor U7542 (N_7542,N_4277,N_4173);
or U7543 (N_7543,N_4223,N_5293);
and U7544 (N_7544,N_4403,N_3521);
nor U7545 (N_7545,N_3041,N_5174);
nand U7546 (N_7546,N_3118,N_3026);
or U7547 (N_7547,N_3296,N_5917);
nand U7548 (N_7548,N_3766,N_3746);
and U7549 (N_7549,N_4573,N_3826);
or U7550 (N_7550,N_4547,N_4116);
nor U7551 (N_7551,N_3300,N_4547);
nand U7552 (N_7552,N_3070,N_4380);
and U7553 (N_7553,N_3365,N_5025);
or U7554 (N_7554,N_4955,N_4125);
xor U7555 (N_7555,N_5283,N_5630);
and U7556 (N_7556,N_3931,N_5655);
xor U7557 (N_7557,N_3116,N_3229);
or U7558 (N_7558,N_5441,N_4387);
and U7559 (N_7559,N_4597,N_4404);
and U7560 (N_7560,N_4481,N_3227);
nand U7561 (N_7561,N_4752,N_5999);
nor U7562 (N_7562,N_4272,N_3502);
or U7563 (N_7563,N_3806,N_5069);
nand U7564 (N_7564,N_5136,N_5959);
or U7565 (N_7565,N_5935,N_5442);
or U7566 (N_7566,N_4742,N_5930);
nor U7567 (N_7567,N_4480,N_4528);
and U7568 (N_7568,N_4744,N_4427);
nor U7569 (N_7569,N_4648,N_5771);
and U7570 (N_7570,N_5704,N_3960);
nor U7571 (N_7571,N_3830,N_4838);
nand U7572 (N_7572,N_3762,N_4990);
and U7573 (N_7573,N_3973,N_4503);
and U7574 (N_7574,N_4412,N_4345);
and U7575 (N_7575,N_5383,N_4427);
nand U7576 (N_7576,N_3039,N_4334);
nand U7577 (N_7577,N_4547,N_3142);
nor U7578 (N_7578,N_3899,N_5895);
and U7579 (N_7579,N_5662,N_4169);
xnor U7580 (N_7580,N_5428,N_4106);
xnor U7581 (N_7581,N_4742,N_3633);
or U7582 (N_7582,N_5571,N_5262);
nor U7583 (N_7583,N_3933,N_3374);
nor U7584 (N_7584,N_4363,N_5176);
and U7585 (N_7585,N_4852,N_5780);
and U7586 (N_7586,N_5172,N_4988);
or U7587 (N_7587,N_3151,N_4911);
xor U7588 (N_7588,N_3611,N_3750);
or U7589 (N_7589,N_4797,N_5126);
nand U7590 (N_7590,N_3506,N_4759);
nor U7591 (N_7591,N_4323,N_5596);
nor U7592 (N_7592,N_5685,N_3064);
nor U7593 (N_7593,N_5516,N_4752);
nor U7594 (N_7594,N_4808,N_5554);
nor U7595 (N_7595,N_4403,N_4164);
nor U7596 (N_7596,N_4741,N_4426);
nor U7597 (N_7597,N_5805,N_5164);
and U7598 (N_7598,N_3566,N_4230);
or U7599 (N_7599,N_3233,N_5163);
nand U7600 (N_7600,N_3977,N_4191);
and U7601 (N_7601,N_5560,N_3685);
nand U7602 (N_7602,N_4790,N_3666);
nor U7603 (N_7603,N_4068,N_3063);
xnor U7604 (N_7604,N_3631,N_3876);
and U7605 (N_7605,N_3329,N_5135);
or U7606 (N_7606,N_5509,N_4634);
nand U7607 (N_7607,N_4318,N_5597);
nor U7608 (N_7608,N_3623,N_3480);
or U7609 (N_7609,N_3266,N_5065);
and U7610 (N_7610,N_5077,N_5206);
and U7611 (N_7611,N_5140,N_3341);
nand U7612 (N_7612,N_3080,N_5520);
or U7613 (N_7613,N_3732,N_5478);
xor U7614 (N_7614,N_4099,N_3220);
and U7615 (N_7615,N_3972,N_3672);
or U7616 (N_7616,N_5766,N_3011);
or U7617 (N_7617,N_3269,N_5769);
and U7618 (N_7618,N_4217,N_5206);
nor U7619 (N_7619,N_4743,N_5885);
xor U7620 (N_7620,N_4790,N_3091);
nand U7621 (N_7621,N_4527,N_5360);
nand U7622 (N_7622,N_3114,N_4476);
nand U7623 (N_7623,N_4066,N_4793);
xnor U7624 (N_7624,N_3239,N_5703);
or U7625 (N_7625,N_4023,N_5244);
nor U7626 (N_7626,N_4862,N_3778);
nor U7627 (N_7627,N_3579,N_3401);
nor U7628 (N_7628,N_5233,N_4943);
nand U7629 (N_7629,N_5942,N_5224);
xor U7630 (N_7630,N_5276,N_3144);
nor U7631 (N_7631,N_3232,N_3833);
or U7632 (N_7632,N_3979,N_5774);
nor U7633 (N_7633,N_3229,N_3069);
nor U7634 (N_7634,N_4096,N_4921);
and U7635 (N_7635,N_4153,N_3654);
xor U7636 (N_7636,N_3744,N_3705);
and U7637 (N_7637,N_3284,N_3821);
or U7638 (N_7638,N_5742,N_3921);
nand U7639 (N_7639,N_4233,N_4534);
nand U7640 (N_7640,N_4150,N_4811);
nor U7641 (N_7641,N_3772,N_3786);
nor U7642 (N_7642,N_3979,N_3206);
and U7643 (N_7643,N_3995,N_3310);
and U7644 (N_7644,N_4330,N_3889);
xnor U7645 (N_7645,N_5299,N_5493);
or U7646 (N_7646,N_5721,N_5368);
or U7647 (N_7647,N_5410,N_4191);
or U7648 (N_7648,N_5053,N_3256);
nand U7649 (N_7649,N_4967,N_5142);
or U7650 (N_7650,N_5328,N_5074);
nor U7651 (N_7651,N_3830,N_3342);
or U7652 (N_7652,N_3748,N_3223);
and U7653 (N_7653,N_3258,N_4408);
and U7654 (N_7654,N_3615,N_5478);
and U7655 (N_7655,N_4419,N_5158);
nor U7656 (N_7656,N_4606,N_5481);
and U7657 (N_7657,N_5586,N_5297);
or U7658 (N_7658,N_5646,N_4818);
nor U7659 (N_7659,N_5523,N_5236);
nor U7660 (N_7660,N_4148,N_5546);
nor U7661 (N_7661,N_5062,N_3016);
and U7662 (N_7662,N_5106,N_5399);
or U7663 (N_7663,N_5289,N_4634);
and U7664 (N_7664,N_4243,N_3644);
nor U7665 (N_7665,N_4009,N_3085);
nand U7666 (N_7666,N_4516,N_3578);
nand U7667 (N_7667,N_3915,N_4612);
nand U7668 (N_7668,N_4586,N_4771);
or U7669 (N_7669,N_5570,N_4162);
or U7670 (N_7670,N_5885,N_5261);
xnor U7671 (N_7671,N_3027,N_4367);
or U7672 (N_7672,N_5652,N_5051);
and U7673 (N_7673,N_4227,N_4926);
nor U7674 (N_7674,N_4733,N_3794);
and U7675 (N_7675,N_4151,N_4650);
nand U7676 (N_7676,N_5139,N_5423);
xor U7677 (N_7677,N_4079,N_5779);
and U7678 (N_7678,N_5215,N_5553);
nand U7679 (N_7679,N_5775,N_5238);
xnor U7680 (N_7680,N_3282,N_4451);
and U7681 (N_7681,N_3225,N_3249);
or U7682 (N_7682,N_4363,N_3163);
nor U7683 (N_7683,N_5577,N_4482);
or U7684 (N_7684,N_4310,N_5758);
nand U7685 (N_7685,N_4031,N_3394);
xor U7686 (N_7686,N_3078,N_3980);
or U7687 (N_7687,N_3688,N_5840);
nor U7688 (N_7688,N_5218,N_5648);
or U7689 (N_7689,N_3583,N_3716);
and U7690 (N_7690,N_4882,N_4724);
and U7691 (N_7691,N_4631,N_3333);
nand U7692 (N_7692,N_5192,N_5771);
and U7693 (N_7693,N_4148,N_3987);
or U7694 (N_7694,N_5601,N_4472);
nor U7695 (N_7695,N_5968,N_3845);
nand U7696 (N_7696,N_5491,N_5819);
nor U7697 (N_7697,N_4578,N_4200);
and U7698 (N_7698,N_3297,N_4317);
nand U7699 (N_7699,N_4996,N_4419);
nand U7700 (N_7700,N_4102,N_3912);
or U7701 (N_7701,N_4854,N_3310);
nor U7702 (N_7702,N_3175,N_4247);
nor U7703 (N_7703,N_4871,N_4631);
nand U7704 (N_7704,N_3743,N_3140);
xor U7705 (N_7705,N_3006,N_3224);
and U7706 (N_7706,N_5664,N_5501);
nor U7707 (N_7707,N_3755,N_3351);
or U7708 (N_7708,N_4574,N_3011);
and U7709 (N_7709,N_5213,N_3486);
nand U7710 (N_7710,N_3738,N_4602);
nand U7711 (N_7711,N_5211,N_5032);
or U7712 (N_7712,N_5645,N_4683);
or U7713 (N_7713,N_5453,N_4888);
nor U7714 (N_7714,N_3211,N_3299);
nand U7715 (N_7715,N_5215,N_5650);
nor U7716 (N_7716,N_3902,N_4321);
and U7717 (N_7717,N_4684,N_5190);
xnor U7718 (N_7718,N_5075,N_3128);
xnor U7719 (N_7719,N_3997,N_4155);
and U7720 (N_7720,N_3056,N_5902);
and U7721 (N_7721,N_3458,N_4159);
xnor U7722 (N_7722,N_4802,N_4715);
xor U7723 (N_7723,N_4093,N_3644);
or U7724 (N_7724,N_3986,N_5703);
and U7725 (N_7725,N_5253,N_4565);
nand U7726 (N_7726,N_5087,N_3438);
or U7727 (N_7727,N_4761,N_5040);
nand U7728 (N_7728,N_3910,N_5542);
and U7729 (N_7729,N_4287,N_5350);
nand U7730 (N_7730,N_5858,N_3260);
xor U7731 (N_7731,N_3678,N_5707);
or U7732 (N_7732,N_4881,N_4719);
or U7733 (N_7733,N_5431,N_3668);
nand U7734 (N_7734,N_4548,N_5066);
nand U7735 (N_7735,N_3191,N_4081);
or U7736 (N_7736,N_4557,N_3764);
xor U7737 (N_7737,N_3649,N_3363);
and U7738 (N_7738,N_3056,N_3621);
nor U7739 (N_7739,N_4508,N_3148);
nand U7740 (N_7740,N_5714,N_3133);
or U7741 (N_7741,N_5055,N_3281);
or U7742 (N_7742,N_4976,N_3693);
or U7743 (N_7743,N_4421,N_3619);
xnor U7744 (N_7744,N_4723,N_5286);
nor U7745 (N_7745,N_5755,N_3952);
nor U7746 (N_7746,N_3316,N_4401);
nor U7747 (N_7747,N_3989,N_5991);
or U7748 (N_7748,N_4701,N_3716);
and U7749 (N_7749,N_5004,N_4011);
and U7750 (N_7750,N_5205,N_5787);
nand U7751 (N_7751,N_3065,N_5528);
nor U7752 (N_7752,N_3306,N_3322);
and U7753 (N_7753,N_4175,N_3213);
or U7754 (N_7754,N_4259,N_4897);
or U7755 (N_7755,N_3342,N_5868);
or U7756 (N_7756,N_3042,N_5614);
or U7757 (N_7757,N_3542,N_5382);
and U7758 (N_7758,N_5032,N_5750);
nand U7759 (N_7759,N_5340,N_5981);
nor U7760 (N_7760,N_4884,N_5582);
nand U7761 (N_7761,N_4911,N_3598);
or U7762 (N_7762,N_5419,N_3450);
or U7763 (N_7763,N_4678,N_5808);
nor U7764 (N_7764,N_4664,N_3698);
xnor U7765 (N_7765,N_3856,N_5383);
xnor U7766 (N_7766,N_5518,N_3676);
nand U7767 (N_7767,N_3328,N_3217);
and U7768 (N_7768,N_5036,N_4750);
nor U7769 (N_7769,N_5006,N_3368);
xnor U7770 (N_7770,N_3417,N_4711);
or U7771 (N_7771,N_3306,N_3675);
nor U7772 (N_7772,N_4799,N_3689);
and U7773 (N_7773,N_5357,N_5864);
nor U7774 (N_7774,N_3546,N_5031);
nand U7775 (N_7775,N_3469,N_3324);
xor U7776 (N_7776,N_3403,N_3327);
nor U7777 (N_7777,N_5155,N_4392);
nor U7778 (N_7778,N_3641,N_3865);
or U7779 (N_7779,N_5499,N_3794);
nor U7780 (N_7780,N_5932,N_3126);
nor U7781 (N_7781,N_4980,N_4526);
xor U7782 (N_7782,N_3761,N_5299);
nand U7783 (N_7783,N_4905,N_4104);
nand U7784 (N_7784,N_4732,N_4185);
nand U7785 (N_7785,N_4184,N_5064);
xnor U7786 (N_7786,N_3975,N_5078);
nand U7787 (N_7787,N_5087,N_4276);
and U7788 (N_7788,N_3886,N_4211);
xnor U7789 (N_7789,N_5300,N_5692);
or U7790 (N_7790,N_3542,N_4812);
nand U7791 (N_7791,N_3631,N_5537);
and U7792 (N_7792,N_3424,N_3385);
or U7793 (N_7793,N_4421,N_4216);
and U7794 (N_7794,N_4056,N_4831);
and U7795 (N_7795,N_3447,N_4838);
xor U7796 (N_7796,N_3021,N_3088);
nor U7797 (N_7797,N_5913,N_4554);
or U7798 (N_7798,N_4533,N_3363);
xnor U7799 (N_7799,N_4060,N_3732);
nand U7800 (N_7800,N_4273,N_3165);
nand U7801 (N_7801,N_5595,N_5997);
and U7802 (N_7802,N_5386,N_3463);
nor U7803 (N_7803,N_5049,N_4631);
or U7804 (N_7804,N_5520,N_4306);
nor U7805 (N_7805,N_5445,N_5775);
or U7806 (N_7806,N_3828,N_4834);
nand U7807 (N_7807,N_4289,N_5464);
or U7808 (N_7808,N_3121,N_3823);
nor U7809 (N_7809,N_3095,N_3402);
nand U7810 (N_7810,N_5542,N_5286);
nor U7811 (N_7811,N_3425,N_4852);
nor U7812 (N_7812,N_5553,N_4583);
or U7813 (N_7813,N_4373,N_3846);
nor U7814 (N_7814,N_4045,N_3002);
nand U7815 (N_7815,N_4646,N_4022);
and U7816 (N_7816,N_4306,N_5912);
or U7817 (N_7817,N_5439,N_5976);
or U7818 (N_7818,N_4848,N_5986);
xnor U7819 (N_7819,N_4699,N_5062);
and U7820 (N_7820,N_4409,N_4778);
nor U7821 (N_7821,N_3769,N_5218);
and U7822 (N_7822,N_4959,N_4551);
nor U7823 (N_7823,N_5394,N_3167);
or U7824 (N_7824,N_3562,N_4051);
xor U7825 (N_7825,N_4109,N_4598);
xnor U7826 (N_7826,N_5367,N_5442);
or U7827 (N_7827,N_4421,N_3670);
nand U7828 (N_7828,N_5571,N_4706);
nor U7829 (N_7829,N_5065,N_5247);
nor U7830 (N_7830,N_4415,N_5484);
and U7831 (N_7831,N_5987,N_3188);
xor U7832 (N_7832,N_3047,N_4600);
nand U7833 (N_7833,N_4508,N_4520);
nor U7834 (N_7834,N_3831,N_5455);
and U7835 (N_7835,N_5334,N_5865);
nor U7836 (N_7836,N_3678,N_5627);
and U7837 (N_7837,N_3385,N_5774);
and U7838 (N_7838,N_3996,N_5804);
nand U7839 (N_7839,N_4902,N_3410);
and U7840 (N_7840,N_3872,N_3492);
and U7841 (N_7841,N_4537,N_3834);
and U7842 (N_7842,N_3612,N_5006);
or U7843 (N_7843,N_4359,N_5918);
or U7844 (N_7844,N_5212,N_5020);
or U7845 (N_7845,N_4316,N_5266);
and U7846 (N_7846,N_3849,N_3052);
or U7847 (N_7847,N_4545,N_3067);
xnor U7848 (N_7848,N_5108,N_3628);
and U7849 (N_7849,N_4366,N_3713);
nand U7850 (N_7850,N_5383,N_3175);
nor U7851 (N_7851,N_5803,N_3122);
xor U7852 (N_7852,N_3306,N_4923);
or U7853 (N_7853,N_4400,N_4065);
and U7854 (N_7854,N_4170,N_4772);
xor U7855 (N_7855,N_5063,N_5255);
or U7856 (N_7856,N_3517,N_4654);
nand U7857 (N_7857,N_4678,N_5107);
nor U7858 (N_7858,N_4752,N_5305);
nor U7859 (N_7859,N_4453,N_5028);
or U7860 (N_7860,N_5826,N_4163);
and U7861 (N_7861,N_3697,N_4566);
nor U7862 (N_7862,N_3769,N_4167);
nor U7863 (N_7863,N_3149,N_5602);
nand U7864 (N_7864,N_5343,N_3322);
and U7865 (N_7865,N_3486,N_3299);
nand U7866 (N_7866,N_5455,N_3922);
or U7867 (N_7867,N_3644,N_5404);
nand U7868 (N_7868,N_3132,N_3285);
xor U7869 (N_7869,N_3611,N_4478);
and U7870 (N_7870,N_5823,N_4832);
or U7871 (N_7871,N_5208,N_5599);
nor U7872 (N_7872,N_4645,N_5623);
xnor U7873 (N_7873,N_4148,N_3433);
nor U7874 (N_7874,N_3972,N_4180);
or U7875 (N_7875,N_3155,N_5252);
or U7876 (N_7876,N_3723,N_3186);
and U7877 (N_7877,N_4988,N_4125);
or U7878 (N_7878,N_5639,N_3802);
or U7879 (N_7879,N_5539,N_3482);
nor U7880 (N_7880,N_5789,N_3281);
nor U7881 (N_7881,N_3951,N_5923);
and U7882 (N_7882,N_3292,N_3210);
and U7883 (N_7883,N_3222,N_5512);
nor U7884 (N_7884,N_4500,N_5865);
and U7885 (N_7885,N_3280,N_5503);
or U7886 (N_7886,N_4622,N_4587);
nor U7887 (N_7887,N_4407,N_3654);
nor U7888 (N_7888,N_3886,N_4413);
xnor U7889 (N_7889,N_5573,N_4943);
xor U7890 (N_7890,N_5771,N_4328);
xnor U7891 (N_7891,N_4532,N_5434);
nand U7892 (N_7892,N_3819,N_5332);
nor U7893 (N_7893,N_5795,N_5206);
nand U7894 (N_7894,N_3557,N_5479);
and U7895 (N_7895,N_4665,N_4105);
nand U7896 (N_7896,N_5542,N_5917);
and U7897 (N_7897,N_5624,N_5619);
and U7898 (N_7898,N_4968,N_3217);
xor U7899 (N_7899,N_5882,N_5304);
nor U7900 (N_7900,N_5392,N_4158);
and U7901 (N_7901,N_5088,N_5137);
and U7902 (N_7902,N_4795,N_3202);
nor U7903 (N_7903,N_5332,N_4368);
and U7904 (N_7904,N_4688,N_3797);
xor U7905 (N_7905,N_5386,N_4273);
nor U7906 (N_7906,N_5498,N_3163);
xnor U7907 (N_7907,N_4958,N_4194);
nand U7908 (N_7908,N_3710,N_3749);
or U7909 (N_7909,N_5007,N_3113);
and U7910 (N_7910,N_4041,N_3483);
nand U7911 (N_7911,N_5735,N_4235);
nor U7912 (N_7912,N_4610,N_5760);
and U7913 (N_7913,N_3758,N_4200);
nor U7914 (N_7914,N_5870,N_4762);
and U7915 (N_7915,N_5938,N_3964);
nand U7916 (N_7916,N_4533,N_3450);
or U7917 (N_7917,N_5650,N_3616);
xor U7918 (N_7918,N_4159,N_4137);
nand U7919 (N_7919,N_4399,N_3195);
nor U7920 (N_7920,N_5446,N_5934);
nand U7921 (N_7921,N_3607,N_3063);
and U7922 (N_7922,N_3010,N_5638);
xor U7923 (N_7923,N_5427,N_4681);
and U7924 (N_7924,N_5458,N_5212);
and U7925 (N_7925,N_4400,N_5469);
nor U7926 (N_7926,N_4181,N_4274);
and U7927 (N_7927,N_3234,N_4629);
nand U7928 (N_7928,N_3882,N_3714);
or U7929 (N_7929,N_5245,N_5983);
nor U7930 (N_7930,N_5632,N_5533);
and U7931 (N_7931,N_4365,N_4097);
and U7932 (N_7932,N_5280,N_4148);
nor U7933 (N_7933,N_5869,N_4708);
nor U7934 (N_7934,N_5010,N_3481);
or U7935 (N_7935,N_4616,N_5592);
nand U7936 (N_7936,N_5080,N_5622);
nand U7937 (N_7937,N_3188,N_3836);
or U7938 (N_7938,N_4945,N_3927);
or U7939 (N_7939,N_5010,N_5223);
or U7940 (N_7940,N_4252,N_3680);
or U7941 (N_7941,N_3289,N_3824);
or U7942 (N_7942,N_3307,N_5100);
and U7943 (N_7943,N_3657,N_3522);
or U7944 (N_7944,N_5566,N_4232);
nor U7945 (N_7945,N_5146,N_3401);
and U7946 (N_7946,N_3062,N_5242);
nand U7947 (N_7947,N_5509,N_4672);
nand U7948 (N_7948,N_5681,N_5911);
nand U7949 (N_7949,N_5731,N_4729);
and U7950 (N_7950,N_4154,N_5368);
or U7951 (N_7951,N_4403,N_3793);
nor U7952 (N_7952,N_5047,N_3396);
xor U7953 (N_7953,N_3281,N_4066);
nor U7954 (N_7954,N_3935,N_3429);
and U7955 (N_7955,N_5901,N_5053);
and U7956 (N_7956,N_5062,N_5605);
or U7957 (N_7957,N_3180,N_5554);
and U7958 (N_7958,N_5037,N_3876);
nand U7959 (N_7959,N_5423,N_4981);
or U7960 (N_7960,N_5125,N_5388);
or U7961 (N_7961,N_3319,N_5787);
nand U7962 (N_7962,N_3437,N_4718);
xor U7963 (N_7963,N_3358,N_4670);
or U7964 (N_7964,N_5133,N_4097);
or U7965 (N_7965,N_5678,N_5465);
nand U7966 (N_7966,N_3887,N_3799);
and U7967 (N_7967,N_3378,N_3922);
or U7968 (N_7968,N_3344,N_3335);
or U7969 (N_7969,N_5972,N_4181);
and U7970 (N_7970,N_4817,N_3635);
nand U7971 (N_7971,N_4879,N_5816);
and U7972 (N_7972,N_4007,N_3929);
nand U7973 (N_7973,N_4423,N_3851);
nand U7974 (N_7974,N_5282,N_3096);
or U7975 (N_7975,N_4614,N_3271);
or U7976 (N_7976,N_5755,N_3303);
nor U7977 (N_7977,N_3326,N_3107);
nand U7978 (N_7978,N_5352,N_5361);
nor U7979 (N_7979,N_3447,N_3059);
nor U7980 (N_7980,N_5472,N_5381);
and U7981 (N_7981,N_5126,N_5659);
nand U7982 (N_7982,N_3283,N_4121);
nand U7983 (N_7983,N_3423,N_3777);
nand U7984 (N_7984,N_5072,N_3640);
or U7985 (N_7985,N_3536,N_4734);
or U7986 (N_7986,N_4599,N_3234);
nand U7987 (N_7987,N_4156,N_5893);
nor U7988 (N_7988,N_4213,N_5807);
or U7989 (N_7989,N_5576,N_4276);
and U7990 (N_7990,N_3378,N_5977);
xor U7991 (N_7991,N_3249,N_5742);
nand U7992 (N_7992,N_3489,N_4629);
or U7993 (N_7993,N_3476,N_3455);
and U7994 (N_7994,N_3701,N_3691);
nand U7995 (N_7995,N_3064,N_3179);
nand U7996 (N_7996,N_4747,N_3817);
nor U7997 (N_7997,N_4206,N_4406);
nand U7998 (N_7998,N_5723,N_3938);
xnor U7999 (N_7999,N_5800,N_4684);
nor U8000 (N_8000,N_3698,N_5265);
nor U8001 (N_8001,N_4510,N_3311);
nand U8002 (N_8002,N_3557,N_5329);
and U8003 (N_8003,N_5095,N_5978);
or U8004 (N_8004,N_3383,N_5785);
nand U8005 (N_8005,N_5380,N_4035);
or U8006 (N_8006,N_4857,N_4986);
xnor U8007 (N_8007,N_3008,N_3786);
and U8008 (N_8008,N_4947,N_3496);
nor U8009 (N_8009,N_5751,N_3685);
and U8010 (N_8010,N_3697,N_3745);
and U8011 (N_8011,N_4199,N_4797);
nor U8012 (N_8012,N_5715,N_3987);
nor U8013 (N_8013,N_3880,N_3315);
and U8014 (N_8014,N_5437,N_4067);
nor U8015 (N_8015,N_4453,N_3142);
and U8016 (N_8016,N_3602,N_5313);
xnor U8017 (N_8017,N_5993,N_3202);
or U8018 (N_8018,N_4705,N_4977);
nor U8019 (N_8019,N_5450,N_5548);
nor U8020 (N_8020,N_5107,N_5688);
nor U8021 (N_8021,N_5534,N_4570);
nor U8022 (N_8022,N_5622,N_4159);
and U8023 (N_8023,N_3570,N_4719);
or U8024 (N_8024,N_4712,N_3615);
nor U8025 (N_8025,N_5939,N_4426);
and U8026 (N_8026,N_5222,N_3241);
nand U8027 (N_8027,N_4157,N_4012);
nor U8028 (N_8028,N_4479,N_4994);
nor U8029 (N_8029,N_5796,N_3380);
nor U8030 (N_8030,N_4565,N_3607);
or U8031 (N_8031,N_5637,N_5143);
xor U8032 (N_8032,N_5564,N_4725);
nor U8033 (N_8033,N_4986,N_5989);
nor U8034 (N_8034,N_5408,N_5507);
nor U8035 (N_8035,N_3471,N_4808);
and U8036 (N_8036,N_4896,N_3988);
and U8037 (N_8037,N_3712,N_5815);
nand U8038 (N_8038,N_4811,N_4297);
xnor U8039 (N_8039,N_4219,N_5615);
nor U8040 (N_8040,N_5764,N_4596);
nor U8041 (N_8041,N_3301,N_5518);
or U8042 (N_8042,N_5604,N_4403);
or U8043 (N_8043,N_5858,N_3925);
nand U8044 (N_8044,N_4835,N_5607);
or U8045 (N_8045,N_3200,N_4168);
or U8046 (N_8046,N_5300,N_4311);
and U8047 (N_8047,N_3817,N_3562);
and U8048 (N_8048,N_5969,N_3707);
xor U8049 (N_8049,N_5558,N_3796);
and U8050 (N_8050,N_3165,N_5388);
nand U8051 (N_8051,N_3176,N_5238);
nand U8052 (N_8052,N_5029,N_4937);
and U8053 (N_8053,N_5638,N_3816);
and U8054 (N_8054,N_4658,N_4359);
or U8055 (N_8055,N_3853,N_5602);
and U8056 (N_8056,N_5866,N_3202);
and U8057 (N_8057,N_3624,N_5829);
and U8058 (N_8058,N_4234,N_3901);
and U8059 (N_8059,N_5163,N_3744);
nand U8060 (N_8060,N_5964,N_4929);
and U8061 (N_8061,N_4144,N_3608);
xor U8062 (N_8062,N_4153,N_3202);
and U8063 (N_8063,N_4864,N_4628);
nand U8064 (N_8064,N_3191,N_4801);
or U8065 (N_8065,N_3426,N_3994);
and U8066 (N_8066,N_3187,N_3716);
nand U8067 (N_8067,N_3547,N_4580);
xnor U8068 (N_8068,N_5466,N_5004);
nand U8069 (N_8069,N_5199,N_4430);
and U8070 (N_8070,N_5632,N_5089);
or U8071 (N_8071,N_4544,N_5849);
nor U8072 (N_8072,N_5330,N_3557);
and U8073 (N_8073,N_3485,N_4268);
nand U8074 (N_8074,N_4186,N_5357);
nand U8075 (N_8075,N_4003,N_5162);
nor U8076 (N_8076,N_3638,N_5279);
nor U8077 (N_8077,N_4691,N_3207);
nand U8078 (N_8078,N_4213,N_4520);
nand U8079 (N_8079,N_4455,N_4558);
nand U8080 (N_8080,N_4731,N_5956);
nand U8081 (N_8081,N_4542,N_5504);
nand U8082 (N_8082,N_3051,N_3858);
or U8083 (N_8083,N_5451,N_3723);
nand U8084 (N_8084,N_4486,N_3864);
nand U8085 (N_8085,N_4717,N_3367);
nand U8086 (N_8086,N_3090,N_5886);
and U8087 (N_8087,N_3905,N_5899);
and U8088 (N_8088,N_4578,N_5843);
nor U8089 (N_8089,N_4178,N_4549);
and U8090 (N_8090,N_3680,N_3221);
nand U8091 (N_8091,N_3399,N_3331);
or U8092 (N_8092,N_4380,N_4268);
xnor U8093 (N_8093,N_5454,N_3773);
nor U8094 (N_8094,N_4870,N_5749);
or U8095 (N_8095,N_5923,N_5448);
nand U8096 (N_8096,N_3226,N_5326);
and U8097 (N_8097,N_5290,N_4512);
and U8098 (N_8098,N_4473,N_3192);
nor U8099 (N_8099,N_4282,N_4468);
or U8100 (N_8100,N_4975,N_3517);
nand U8101 (N_8101,N_5159,N_3938);
xnor U8102 (N_8102,N_4925,N_3826);
nor U8103 (N_8103,N_4950,N_3082);
nor U8104 (N_8104,N_3879,N_4151);
and U8105 (N_8105,N_3331,N_5402);
and U8106 (N_8106,N_4986,N_4033);
nor U8107 (N_8107,N_3890,N_3619);
or U8108 (N_8108,N_5625,N_3793);
xor U8109 (N_8109,N_5950,N_3428);
xnor U8110 (N_8110,N_3433,N_4933);
nand U8111 (N_8111,N_5722,N_5642);
xnor U8112 (N_8112,N_4158,N_4380);
and U8113 (N_8113,N_5384,N_3965);
nor U8114 (N_8114,N_4354,N_3814);
or U8115 (N_8115,N_4545,N_3984);
or U8116 (N_8116,N_3793,N_5813);
or U8117 (N_8117,N_5910,N_5738);
or U8118 (N_8118,N_4117,N_5505);
xor U8119 (N_8119,N_5188,N_3293);
or U8120 (N_8120,N_3035,N_3549);
nand U8121 (N_8121,N_5972,N_3697);
nand U8122 (N_8122,N_5013,N_5726);
and U8123 (N_8123,N_3749,N_4342);
or U8124 (N_8124,N_5856,N_3367);
or U8125 (N_8125,N_4725,N_5778);
and U8126 (N_8126,N_4950,N_5825);
nand U8127 (N_8127,N_5068,N_5555);
and U8128 (N_8128,N_4657,N_3873);
or U8129 (N_8129,N_5557,N_3077);
nand U8130 (N_8130,N_5854,N_5421);
or U8131 (N_8131,N_4800,N_4024);
or U8132 (N_8132,N_4267,N_5930);
and U8133 (N_8133,N_5080,N_4721);
nor U8134 (N_8134,N_5328,N_5213);
xnor U8135 (N_8135,N_4355,N_5844);
or U8136 (N_8136,N_4377,N_3517);
nand U8137 (N_8137,N_4075,N_5891);
nor U8138 (N_8138,N_4267,N_3812);
xor U8139 (N_8139,N_4494,N_4812);
or U8140 (N_8140,N_5520,N_3374);
nor U8141 (N_8141,N_4080,N_4584);
nor U8142 (N_8142,N_3308,N_4099);
xnor U8143 (N_8143,N_4538,N_3719);
nand U8144 (N_8144,N_4207,N_4084);
nor U8145 (N_8145,N_4804,N_3615);
nor U8146 (N_8146,N_3771,N_5547);
xnor U8147 (N_8147,N_5667,N_4466);
nor U8148 (N_8148,N_4426,N_3382);
xnor U8149 (N_8149,N_3962,N_4452);
and U8150 (N_8150,N_5012,N_5460);
nor U8151 (N_8151,N_3312,N_5554);
nand U8152 (N_8152,N_5723,N_4867);
nor U8153 (N_8153,N_3684,N_5714);
nor U8154 (N_8154,N_5064,N_3562);
xnor U8155 (N_8155,N_4150,N_4449);
nand U8156 (N_8156,N_4645,N_3533);
nand U8157 (N_8157,N_3936,N_4827);
nand U8158 (N_8158,N_3245,N_3331);
nor U8159 (N_8159,N_5614,N_4975);
or U8160 (N_8160,N_5579,N_3695);
or U8161 (N_8161,N_4270,N_4857);
xnor U8162 (N_8162,N_5658,N_4133);
and U8163 (N_8163,N_5825,N_3292);
and U8164 (N_8164,N_5432,N_3956);
nand U8165 (N_8165,N_5039,N_5448);
or U8166 (N_8166,N_5341,N_5694);
and U8167 (N_8167,N_5700,N_5862);
xor U8168 (N_8168,N_5830,N_4083);
and U8169 (N_8169,N_5774,N_5088);
and U8170 (N_8170,N_5646,N_5328);
nor U8171 (N_8171,N_3587,N_3980);
and U8172 (N_8172,N_4025,N_3560);
or U8173 (N_8173,N_4110,N_4511);
nand U8174 (N_8174,N_5988,N_3507);
nand U8175 (N_8175,N_5294,N_5733);
nor U8176 (N_8176,N_4660,N_3839);
nand U8177 (N_8177,N_5685,N_3575);
nand U8178 (N_8178,N_5431,N_4063);
and U8179 (N_8179,N_4060,N_4312);
and U8180 (N_8180,N_5305,N_5426);
and U8181 (N_8181,N_3710,N_4723);
nand U8182 (N_8182,N_4565,N_3014);
and U8183 (N_8183,N_5289,N_5718);
nor U8184 (N_8184,N_3210,N_4003);
nand U8185 (N_8185,N_3529,N_5684);
or U8186 (N_8186,N_4127,N_5545);
nand U8187 (N_8187,N_3023,N_4288);
or U8188 (N_8188,N_4011,N_5173);
nand U8189 (N_8189,N_4938,N_3490);
nand U8190 (N_8190,N_5285,N_4899);
or U8191 (N_8191,N_5428,N_3397);
nor U8192 (N_8192,N_3861,N_3269);
or U8193 (N_8193,N_3271,N_5522);
nand U8194 (N_8194,N_4083,N_4005);
or U8195 (N_8195,N_5789,N_4375);
nand U8196 (N_8196,N_5344,N_4158);
or U8197 (N_8197,N_3666,N_4378);
or U8198 (N_8198,N_3363,N_5240);
or U8199 (N_8199,N_5856,N_5376);
nand U8200 (N_8200,N_3230,N_5312);
nor U8201 (N_8201,N_4975,N_3201);
or U8202 (N_8202,N_3737,N_3628);
nand U8203 (N_8203,N_3245,N_4837);
nand U8204 (N_8204,N_4871,N_4720);
nand U8205 (N_8205,N_3813,N_5312);
nand U8206 (N_8206,N_4335,N_5635);
or U8207 (N_8207,N_3143,N_3704);
xor U8208 (N_8208,N_5175,N_5958);
nand U8209 (N_8209,N_4970,N_3049);
or U8210 (N_8210,N_5140,N_4437);
nor U8211 (N_8211,N_4738,N_3333);
nand U8212 (N_8212,N_5492,N_3424);
and U8213 (N_8213,N_4909,N_4610);
and U8214 (N_8214,N_5783,N_3781);
nand U8215 (N_8215,N_3572,N_4891);
and U8216 (N_8216,N_3874,N_5723);
xor U8217 (N_8217,N_3222,N_5736);
nor U8218 (N_8218,N_3474,N_4138);
nor U8219 (N_8219,N_5736,N_3730);
nor U8220 (N_8220,N_5316,N_4031);
and U8221 (N_8221,N_3273,N_5099);
or U8222 (N_8222,N_4162,N_3431);
or U8223 (N_8223,N_5315,N_4318);
or U8224 (N_8224,N_5262,N_5925);
and U8225 (N_8225,N_5977,N_3377);
nor U8226 (N_8226,N_3107,N_4999);
xnor U8227 (N_8227,N_5391,N_4450);
and U8228 (N_8228,N_4164,N_5621);
and U8229 (N_8229,N_5906,N_5758);
xnor U8230 (N_8230,N_3845,N_5648);
nand U8231 (N_8231,N_4546,N_3018);
nand U8232 (N_8232,N_5248,N_4452);
nor U8233 (N_8233,N_5258,N_5716);
nand U8234 (N_8234,N_4301,N_4058);
or U8235 (N_8235,N_4921,N_3191);
and U8236 (N_8236,N_3817,N_3673);
nand U8237 (N_8237,N_5285,N_4045);
nor U8238 (N_8238,N_5001,N_4358);
nor U8239 (N_8239,N_3375,N_4629);
nor U8240 (N_8240,N_3668,N_3153);
nand U8241 (N_8241,N_5639,N_3031);
xor U8242 (N_8242,N_3298,N_5549);
nand U8243 (N_8243,N_5573,N_5155);
and U8244 (N_8244,N_4468,N_5362);
and U8245 (N_8245,N_4902,N_5432);
nand U8246 (N_8246,N_3541,N_4756);
nand U8247 (N_8247,N_3170,N_4893);
and U8248 (N_8248,N_5847,N_5298);
nor U8249 (N_8249,N_3926,N_3951);
and U8250 (N_8250,N_3679,N_3851);
xnor U8251 (N_8251,N_5010,N_5030);
nand U8252 (N_8252,N_5381,N_5258);
or U8253 (N_8253,N_5167,N_5415);
nor U8254 (N_8254,N_3819,N_4036);
nand U8255 (N_8255,N_3060,N_3288);
or U8256 (N_8256,N_3312,N_4203);
nor U8257 (N_8257,N_5979,N_4042);
nor U8258 (N_8258,N_5785,N_4254);
and U8259 (N_8259,N_3320,N_4684);
or U8260 (N_8260,N_4412,N_4657);
and U8261 (N_8261,N_3267,N_4452);
or U8262 (N_8262,N_5788,N_3179);
or U8263 (N_8263,N_5343,N_5085);
and U8264 (N_8264,N_3375,N_3924);
or U8265 (N_8265,N_3937,N_4460);
nand U8266 (N_8266,N_3431,N_3532);
nor U8267 (N_8267,N_4529,N_4926);
nand U8268 (N_8268,N_3456,N_4677);
nand U8269 (N_8269,N_3157,N_5184);
nand U8270 (N_8270,N_5103,N_3389);
nor U8271 (N_8271,N_5563,N_3347);
nor U8272 (N_8272,N_5049,N_4987);
or U8273 (N_8273,N_3733,N_4563);
nand U8274 (N_8274,N_5156,N_5310);
nor U8275 (N_8275,N_4033,N_4855);
and U8276 (N_8276,N_4704,N_4673);
nand U8277 (N_8277,N_4528,N_4142);
nand U8278 (N_8278,N_3969,N_4567);
nor U8279 (N_8279,N_5104,N_3098);
or U8280 (N_8280,N_5440,N_4869);
or U8281 (N_8281,N_5232,N_4535);
nand U8282 (N_8282,N_5569,N_4802);
nor U8283 (N_8283,N_5576,N_3720);
or U8284 (N_8284,N_4015,N_3494);
xor U8285 (N_8285,N_3288,N_5678);
xnor U8286 (N_8286,N_3196,N_4174);
and U8287 (N_8287,N_3026,N_3231);
nand U8288 (N_8288,N_3784,N_3538);
nor U8289 (N_8289,N_3281,N_4074);
and U8290 (N_8290,N_5735,N_4104);
or U8291 (N_8291,N_3886,N_4774);
and U8292 (N_8292,N_3614,N_5294);
xnor U8293 (N_8293,N_5998,N_4037);
and U8294 (N_8294,N_4461,N_4843);
nand U8295 (N_8295,N_5440,N_3011);
nor U8296 (N_8296,N_5492,N_3085);
nand U8297 (N_8297,N_3182,N_4013);
nand U8298 (N_8298,N_5278,N_3331);
and U8299 (N_8299,N_3671,N_4359);
xnor U8300 (N_8300,N_5192,N_5005);
or U8301 (N_8301,N_3446,N_5266);
nor U8302 (N_8302,N_3063,N_4015);
nor U8303 (N_8303,N_4332,N_4970);
nor U8304 (N_8304,N_4137,N_4345);
or U8305 (N_8305,N_4055,N_4786);
nand U8306 (N_8306,N_5015,N_4413);
nor U8307 (N_8307,N_5674,N_5645);
xnor U8308 (N_8308,N_5718,N_5179);
nor U8309 (N_8309,N_4403,N_4790);
nand U8310 (N_8310,N_4760,N_4901);
or U8311 (N_8311,N_3390,N_3214);
or U8312 (N_8312,N_3171,N_3572);
xnor U8313 (N_8313,N_4004,N_5169);
nor U8314 (N_8314,N_5085,N_3320);
nand U8315 (N_8315,N_3088,N_3147);
nand U8316 (N_8316,N_4940,N_5984);
nor U8317 (N_8317,N_5543,N_4895);
xor U8318 (N_8318,N_4205,N_4479);
and U8319 (N_8319,N_4333,N_4231);
nand U8320 (N_8320,N_5700,N_3141);
nand U8321 (N_8321,N_5078,N_3179);
and U8322 (N_8322,N_5190,N_3276);
or U8323 (N_8323,N_4775,N_4046);
or U8324 (N_8324,N_4322,N_3668);
or U8325 (N_8325,N_3100,N_5847);
nand U8326 (N_8326,N_3338,N_5837);
or U8327 (N_8327,N_4042,N_3285);
or U8328 (N_8328,N_3705,N_3312);
xor U8329 (N_8329,N_3084,N_4469);
xor U8330 (N_8330,N_5943,N_3173);
nor U8331 (N_8331,N_3917,N_5728);
and U8332 (N_8332,N_5078,N_5620);
xnor U8333 (N_8333,N_4285,N_3163);
nor U8334 (N_8334,N_3907,N_3380);
nor U8335 (N_8335,N_4967,N_5463);
xor U8336 (N_8336,N_5724,N_3634);
nor U8337 (N_8337,N_5038,N_3452);
nor U8338 (N_8338,N_5495,N_5610);
nand U8339 (N_8339,N_4362,N_3527);
xnor U8340 (N_8340,N_3326,N_3712);
or U8341 (N_8341,N_5356,N_3640);
and U8342 (N_8342,N_5219,N_5857);
nand U8343 (N_8343,N_5944,N_3634);
or U8344 (N_8344,N_3881,N_4690);
and U8345 (N_8345,N_4910,N_5740);
and U8346 (N_8346,N_4956,N_3732);
and U8347 (N_8347,N_5951,N_5161);
and U8348 (N_8348,N_5884,N_3190);
and U8349 (N_8349,N_5215,N_5475);
nor U8350 (N_8350,N_5175,N_5403);
or U8351 (N_8351,N_3665,N_4074);
and U8352 (N_8352,N_4007,N_3327);
or U8353 (N_8353,N_5197,N_5744);
nand U8354 (N_8354,N_5023,N_5235);
nor U8355 (N_8355,N_4904,N_4455);
nand U8356 (N_8356,N_4595,N_5299);
nand U8357 (N_8357,N_5875,N_3266);
or U8358 (N_8358,N_3431,N_4772);
nor U8359 (N_8359,N_4868,N_3167);
and U8360 (N_8360,N_5965,N_4229);
nor U8361 (N_8361,N_5284,N_5911);
nand U8362 (N_8362,N_4638,N_4908);
or U8363 (N_8363,N_3060,N_4403);
or U8364 (N_8364,N_4425,N_5600);
xnor U8365 (N_8365,N_5995,N_4160);
nand U8366 (N_8366,N_3680,N_4268);
xnor U8367 (N_8367,N_5473,N_5230);
and U8368 (N_8368,N_4785,N_4775);
nand U8369 (N_8369,N_3371,N_3705);
nand U8370 (N_8370,N_3363,N_5570);
nor U8371 (N_8371,N_3146,N_3150);
nand U8372 (N_8372,N_3659,N_4674);
and U8373 (N_8373,N_5412,N_4686);
or U8374 (N_8374,N_3816,N_4427);
nor U8375 (N_8375,N_3142,N_3174);
nand U8376 (N_8376,N_4459,N_3765);
xor U8377 (N_8377,N_5383,N_4576);
nand U8378 (N_8378,N_5685,N_5433);
and U8379 (N_8379,N_3794,N_3145);
nor U8380 (N_8380,N_4788,N_4724);
nand U8381 (N_8381,N_5752,N_3061);
or U8382 (N_8382,N_5650,N_3907);
nor U8383 (N_8383,N_5975,N_4556);
and U8384 (N_8384,N_4210,N_5306);
nor U8385 (N_8385,N_5117,N_5075);
or U8386 (N_8386,N_5279,N_4134);
xnor U8387 (N_8387,N_3421,N_3182);
or U8388 (N_8388,N_3994,N_5192);
nor U8389 (N_8389,N_4084,N_4309);
nand U8390 (N_8390,N_3646,N_3554);
nand U8391 (N_8391,N_4839,N_4344);
nor U8392 (N_8392,N_3679,N_5286);
nor U8393 (N_8393,N_3072,N_5383);
nand U8394 (N_8394,N_3092,N_3203);
and U8395 (N_8395,N_4674,N_5024);
nand U8396 (N_8396,N_3617,N_3668);
or U8397 (N_8397,N_5408,N_3058);
nor U8398 (N_8398,N_4219,N_5647);
nand U8399 (N_8399,N_4772,N_4563);
nand U8400 (N_8400,N_3773,N_4445);
or U8401 (N_8401,N_5412,N_5992);
nor U8402 (N_8402,N_4963,N_5322);
and U8403 (N_8403,N_4654,N_5846);
and U8404 (N_8404,N_3845,N_3684);
nor U8405 (N_8405,N_4674,N_3761);
nand U8406 (N_8406,N_4051,N_5575);
nor U8407 (N_8407,N_3242,N_3505);
or U8408 (N_8408,N_3161,N_4434);
xnor U8409 (N_8409,N_4051,N_3956);
nand U8410 (N_8410,N_5493,N_3844);
nand U8411 (N_8411,N_4172,N_4290);
xor U8412 (N_8412,N_4423,N_5539);
and U8413 (N_8413,N_3901,N_3476);
and U8414 (N_8414,N_4773,N_4842);
and U8415 (N_8415,N_5695,N_4760);
or U8416 (N_8416,N_3951,N_5646);
and U8417 (N_8417,N_5302,N_5423);
xor U8418 (N_8418,N_4451,N_3159);
and U8419 (N_8419,N_5324,N_4921);
or U8420 (N_8420,N_4203,N_4413);
nor U8421 (N_8421,N_5432,N_3556);
or U8422 (N_8422,N_3216,N_3791);
and U8423 (N_8423,N_3015,N_5428);
nor U8424 (N_8424,N_3119,N_5586);
nand U8425 (N_8425,N_5568,N_3359);
nor U8426 (N_8426,N_5733,N_4544);
nand U8427 (N_8427,N_5398,N_5194);
xor U8428 (N_8428,N_4791,N_5393);
and U8429 (N_8429,N_4227,N_5187);
nor U8430 (N_8430,N_3646,N_5603);
or U8431 (N_8431,N_5661,N_5804);
nor U8432 (N_8432,N_5648,N_4040);
nor U8433 (N_8433,N_3134,N_4400);
xor U8434 (N_8434,N_5733,N_4550);
and U8435 (N_8435,N_5079,N_4824);
nand U8436 (N_8436,N_4871,N_4828);
nand U8437 (N_8437,N_3031,N_3838);
nor U8438 (N_8438,N_4016,N_4573);
nand U8439 (N_8439,N_3566,N_4355);
or U8440 (N_8440,N_5593,N_4380);
or U8441 (N_8441,N_4230,N_3274);
and U8442 (N_8442,N_5413,N_3389);
nor U8443 (N_8443,N_5718,N_3278);
nor U8444 (N_8444,N_5406,N_5088);
nand U8445 (N_8445,N_5569,N_4845);
or U8446 (N_8446,N_5617,N_4767);
nand U8447 (N_8447,N_4983,N_4164);
or U8448 (N_8448,N_4849,N_3312);
nand U8449 (N_8449,N_5900,N_3507);
or U8450 (N_8450,N_5552,N_4960);
xor U8451 (N_8451,N_4013,N_5097);
and U8452 (N_8452,N_5367,N_3679);
nand U8453 (N_8453,N_5062,N_3615);
nor U8454 (N_8454,N_5652,N_3788);
and U8455 (N_8455,N_4812,N_4689);
nor U8456 (N_8456,N_3073,N_3898);
nor U8457 (N_8457,N_5271,N_4846);
xnor U8458 (N_8458,N_4041,N_3272);
nand U8459 (N_8459,N_4829,N_3833);
nand U8460 (N_8460,N_5554,N_3746);
and U8461 (N_8461,N_3331,N_4693);
xor U8462 (N_8462,N_4049,N_4195);
or U8463 (N_8463,N_3494,N_4664);
xor U8464 (N_8464,N_3650,N_4135);
nand U8465 (N_8465,N_5991,N_4926);
or U8466 (N_8466,N_3807,N_5055);
and U8467 (N_8467,N_5305,N_3521);
and U8468 (N_8468,N_5570,N_4663);
and U8469 (N_8469,N_5794,N_3575);
nand U8470 (N_8470,N_5943,N_5500);
or U8471 (N_8471,N_3764,N_3849);
or U8472 (N_8472,N_5250,N_5385);
and U8473 (N_8473,N_3130,N_3131);
or U8474 (N_8474,N_4102,N_3806);
xnor U8475 (N_8475,N_3232,N_5370);
and U8476 (N_8476,N_4149,N_3820);
nand U8477 (N_8477,N_3416,N_3909);
and U8478 (N_8478,N_4662,N_4603);
xor U8479 (N_8479,N_3386,N_4208);
nand U8480 (N_8480,N_4957,N_5055);
nor U8481 (N_8481,N_4638,N_5607);
and U8482 (N_8482,N_3523,N_3802);
or U8483 (N_8483,N_4549,N_4771);
nor U8484 (N_8484,N_3865,N_4671);
nand U8485 (N_8485,N_4308,N_3174);
and U8486 (N_8486,N_5062,N_5132);
and U8487 (N_8487,N_5068,N_3111);
xor U8488 (N_8488,N_5217,N_3178);
nor U8489 (N_8489,N_4173,N_5789);
or U8490 (N_8490,N_3581,N_4315);
or U8491 (N_8491,N_3320,N_3611);
nor U8492 (N_8492,N_3464,N_4740);
or U8493 (N_8493,N_5713,N_5417);
nor U8494 (N_8494,N_5525,N_4326);
or U8495 (N_8495,N_4813,N_4879);
nand U8496 (N_8496,N_5402,N_5963);
nor U8497 (N_8497,N_3268,N_4529);
and U8498 (N_8498,N_5950,N_4423);
and U8499 (N_8499,N_5336,N_4858);
or U8500 (N_8500,N_3944,N_3351);
nor U8501 (N_8501,N_4714,N_4226);
nor U8502 (N_8502,N_3894,N_3387);
and U8503 (N_8503,N_3300,N_5763);
and U8504 (N_8504,N_5628,N_3003);
and U8505 (N_8505,N_4590,N_3701);
nand U8506 (N_8506,N_4243,N_3583);
xnor U8507 (N_8507,N_5667,N_3630);
nand U8508 (N_8508,N_4337,N_4832);
nor U8509 (N_8509,N_5990,N_4985);
nand U8510 (N_8510,N_4452,N_4679);
and U8511 (N_8511,N_5446,N_3804);
nor U8512 (N_8512,N_5020,N_4933);
nor U8513 (N_8513,N_3440,N_5994);
or U8514 (N_8514,N_4013,N_4940);
and U8515 (N_8515,N_3763,N_5260);
and U8516 (N_8516,N_5775,N_3810);
nor U8517 (N_8517,N_5248,N_4241);
and U8518 (N_8518,N_4693,N_3641);
xor U8519 (N_8519,N_3306,N_5299);
and U8520 (N_8520,N_4475,N_3804);
and U8521 (N_8521,N_5179,N_5104);
xor U8522 (N_8522,N_3953,N_3779);
or U8523 (N_8523,N_3360,N_5742);
nor U8524 (N_8524,N_3563,N_4047);
nand U8525 (N_8525,N_4575,N_5181);
xor U8526 (N_8526,N_5313,N_4155);
and U8527 (N_8527,N_3476,N_5798);
and U8528 (N_8528,N_4959,N_3313);
nand U8529 (N_8529,N_5506,N_5899);
nand U8530 (N_8530,N_3741,N_3386);
or U8531 (N_8531,N_5662,N_5689);
xnor U8532 (N_8532,N_4763,N_5527);
nand U8533 (N_8533,N_3522,N_5315);
xnor U8534 (N_8534,N_4880,N_5575);
nor U8535 (N_8535,N_5907,N_5610);
or U8536 (N_8536,N_3372,N_5371);
nand U8537 (N_8537,N_4668,N_3063);
nor U8538 (N_8538,N_3486,N_4101);
xnor U8539 (N_8539,N_3272,N_4436);
xor U8540 (N_8540,N_3879,N_4891);
or U8541 (N_8541,N_3140,N_4970);
or U8542 (N_8542,N_4217,N_4973);
or U8543 (N_8543,N_4027,N_3880);
xor U8544 (N_8544,N_3403,N_5740);
xor U8545 (N_8545,N_4705,N_4577);
and U8546 (N_8546,N_5471,N_4727);
and U8547 (N_8547,N_4404,N_5090);
and U8548 (N_8548,N_5437,N_3662);
or U8549 (N_8549,N_5374,N_3466);
nand U8550 (N_8550,N_3867,N_5633);
nor U8551 (N_8551,N_4844,N_5452);
xor U8552 (N_8552,N_3278,N_5722);
nand U8553 (N_8553,N_5567,N_4730);
and U8554 (N_8554,N_5045,N_5711);
nand U8555 (N_8555,N_3303,N_4750);
and U8556 (N_8556,N_3892,N_3731);
or U8557 (N_8557,N_5700,N_5299);
and U8558 (N_8558,N_4066,N_3357);
nor U8559 (N_8559,N_4053,N_5122);
nor U8560 (N_8560,N_4464,N_4752);
nor U8561 (N_8561,N_4269,N_4320);
nor U8562 (N_8562,N_5141,N_5104);
and U8563 (N_8563,N_3754,N_3680);
nor U8564 (N_8564,N_5883,N_4832);
and U8565 (N_8565,N_4454,N_4909);
or U8566 (N_8566,N_5181,N_3996);
and U8567 (N_8567,N_4741,N_5208);
nor U8568 (N_8568,N_4954,N_5723);
or U8569 (N_8569,N_4653,N_3790);
and U8570 (N_8570,N_4771,N_5531);
or U8571 (N_8571,N_4521,N_5103);
or U8572 (N_8572,N_3774,N_3881);
or U8573 (N_8573,N_5454,N_5924);
or U8574 (N_8574,N_3489,N_4000);
or U8575 (N_8575,N_5861,N_3058);
nand U8576 (N_8576,N_5920,N_4309);
nand U8577 (N_8577,N_5380,N_4317);
nor U8578 (N_8578,N_4367,N_5533);
or U8579 (N_8579,N_4714,N_4116);
nand U8580 (N_8580,N_3129,N_3343);
nand U8581 (N_8581,N_4712,N_3398);
xnor U8582 (N_8582,N_4238,N_3005);
nor U8583 (N_8583,N_4465,N_5221);
nor U8584 (N_8584,N_3093,N_4235);
nand U8585 (N_8585,N_5019,N_3561);
nand U8586 (N_8586,N_4805,N_4671);
or U8587 (N_8587,N_3536,N_3287);
nor U8588 (N_8588,N_4476,N_3350);
and U8589 (N_8589,N_5017,N_5538);
and U8590 (N_8590,N_3626,N_3918);
and U8591 (N_8591,N_5281,N_3539);
xnor U8592 (N_8592,N_3678,N_4379);
or U8593 (N_8593,N_4012,N_5758);
or U8594 (N_8594,N_3519,N_4275);
xnor U8595 (N_8595,N_4769,N_3526);
nand U8596 (N_8596,N_3589,N_3010);
nor U8597 (N_8597,N_3714,N_4043);
nor U8598 (N_8598,N_4708,N_5161);
or U8599 (N_8599,N_3379,N_3206);
nand U8600 (N_8600,N_5390,N_4993);
nor U8601 (N_8601,N_4543,N_4098);
nor U8602 (N_8602,N_5083,N_3276);
nor U8603 (N_8603,N_3284,N_5064);
and U8604 (N_8604,N_4997,N_3683);
nand U8605 (N_8605,N_5577,N_3186);
and U8606 (N_8606,N_5670,N_4339);
nand U8607 (N_8607,N_3380,N_4009);
and U8608 (N_8608,N_3977,N_5229);
and U8609 (N_8609,N_3686,N_5917);
nand U8610 (N_8610,N_4811,N_5504);
nand U8611 (N_8611,N_5453,N_3500);
or U8612 (N_8612,N_3903,N_5983);
nand U8613 (N_8613,N_5185,N_3508);
or U8614 (N_8614,N_4387,N_3267);
nor U8615 (N_8615,N_5025,N_3983);
nor U8616 (N_8616,N_4981,N_4949);
nand U8617 (N_8617,N_5956,N_5688);
nor U8618 (N_8618,N_3047,N_5892);
nor U8619 (N_8619,N_5099,N_4657);
and U8620 (N_8620,N_3789,N_4749);
nor U8621 (N_8621,N_3600,N_3265);
or U8622 (N_8622,N_3182,N_5858);
xnor U8623 (N_8623,N_4575,N_3664);
and U8624 (N_8624,N_3352,N_5614);
and U8625 (N_8625,N_5624,N_5863);
or U8626 (N_8626,N_5352,N_3877);
and U8627 (N_8627,N_5991,N_3275);
and U8628 (N_8628,N_5085,N_4611);
or U8629 (N_8629,N_4959,N_5745);
or U8630 (N_8630,N_5869,N_4130);
nand U8631 (N_8631,N_3044,N_4268);
nor U8632 (N_8632,N_3805,N_5644);
xor U8633 (N_8633,N_5157,N_5500);
and U8634 (N_8634,N_4606,N_5404);
xnor U8635 (N_8635,N_4763,N_5122);
and U8636 (N_8636,N_3866,N_5179);
xor U8637 (N_8637,N_3438,N_5750);
nor U8638 (N_8638,N_4352,N_3581);
or U8639 (N_8639,N_4535,N_4509);
or U8640 (N_8640,N_4628,N_4414);
nor U8641 (N_8641,N_5435,N_5858);
nor U8642 (N_8642,N_5399,N_4084);
or U8643 (N_8643,N_4944,N_3570);
and U8644 (N_8644,N_4557,N_5920);
nor U8645 (N_8645,N_5281,N_5791);
nor U8646 (N_8646,N_5280,N_3624);
and U8647 (N_8647,N_4101,N_3649);
nor U8648 (N_8648,N_5580,N_3157);
nor U8649 (N_8649,N_3617,N_3385);
nor U8650 (N_8650,N_3193,N_4468);
or U8651 (N_8651,N_4402,N_5398);
nand U8652 (N_8652,N_5414,N_3099);
xnor U8653 (N_8653,N_3027,N_5396);
or U8654 (N_8654,N_3933,N_5406);
nor U8655 (N_8655,N_3976,N_3474);
and U8656 (N_8656,N_3238,N_3702);
or U8657 (N_8657,N_4368,N_5706);
nor U8658 (N_8658,N_4353,N_5955);
and U8659 (N_8659,N_4903,N_4020);
nor U8660 (N_8660,N_5292,N_4650);
or U8661 (N_8661,N_5863,N_4837);
nand U8662 (N_8662,N_3335,N_5256);
xnor U8663 (N_8663,N_4094,N_5531);
nor U8664 (N_8664,N_5826,N_3416);
or U8665 (N_8665,N_5981,N_5647);
or U8666 (N_8666,N_4804,N_4393);
or U8667 (N_8667,N_3384,N_5992);
nor U8668 (N_8668,N_3478,N_5247);
nand U8669 (N_8669,N_3931,N_4359);
or U8670 (N_8670,N_4744,N_4524);
nand U8671 (N_8671,N_4481,N_4244);
nor U8672 (N_8672,N_4573,N_3445);
or U8673 (N_8673,N_3704,N_5262);
nand U8674 (N_8674,N_5041,N_5947);
nor U8675 (N_8675,N_5816,N_3727);
nor U8676 (N_8676,N_4425,N_5723);
nand U8677 (N_8677,N_5816,N_5123);
xnor U8678 (N_8678,N_3202,N_4928);
nand U8679 (N_8679,N_4751,N_3080);
xnor U8680 (N_8680,N_5174,N_4677);
or U8681 (N_8681,N_5974,N_3184);
nor U8682 (N_8682,N_4860,N_5188);
and U8683 (N_8683,N_3618,N_5806);
nor U8684 (N_8684,N_5919,N_5898);
or U8685 (N_8685,N_4333,N_5660);
nand U8686 (N_8686,N_4906,N_3331);
and U8687 (N_8687,N_4551,N_4731);
xnor U8688 (N_8688,N_5513,N_4400);
nand U8689 (N_8689,N_5726,N_5592);
xnor U8690 (N_8690,N_5495,N_3794);
and U8691 (N_8691,N_5072,N_4288);
xor U8692 (N_8692,N_4921,N_4141);
and U8693 (N_8693,N_5250,N_3657);
nor U8694 (N_8694,N_4344,N_4823);
and U8695 (N_8695,N_4494,N_3342);
or U8696 (N_8696,N_5339,N_3936);
and U8697 (N_8697,N_5998,N_4188);
or U8698 (N_8698,N_5853,N_4878);
and U8699 (N_8699,N_5661,N_4743);
and U8700 (N_8700,N_3373,N_4951);
and U8701 (N_8701,N_5297,N_4545);
or U8702 (N_8702,N_3937,N_4657);
nor U8703 (N_8703,N_3669,N_5416);
or U8704 (N_8704,N_3779,N_3251);
or U8705 (N_8705,N_4551,N_4850);
xor U8706 (N_8706,N_5685,N_5199);
nor U8707 (N_8707,N_3493,N_4332);
nor U8708 (N_8708,N_3702,N_5561);
nand U8709 (N_8709,N_4136,N_3998);
nand U8710 (N_8710,N_3177,N_4426);
nor U8711 (N_8711,N_5510,N_3800);
nor U8712 (N_8712,N_5147,N_4786);
and U8713 (N_8713,N_4958,N_5360);
nand U8714 (N_8714,N_5449,N_4500);
and U8715 (N_8715,N_5256,N_3508);
and U8716 (N_8716,N_3384,N_4061);
or U8717 (N_8717,N_3429,N_3460);
nor U8718 (N_8718,N_4002,N_4342);
nand U8719 (N_8719,N_3487,N_5889);
nor U8720 (N_8720,N_4855,N_4577);
and U8721 (N_8721,N_4114,N_3306);
nor U8722 (N_8722,N_5543,N_4029);
nand U8723 (N_8723,N_3562,N_5558);
and U8724 (N_8724,N_4625,N_5740);
nor U8725 (N_8725,N_4142,N_3527);
nand U8726 (N_8726,N_5750,N_4426);
nand U8727 (N_8727,N_5048,N_5982);
nor U8728 (N_8728,N_4227,N_5968);
or U8729 (N_8729,N_5612,N_3208);
nor U8730 (N_8730,N_3288,N_4355);
nand U8731 (N_8731,N_5825,N_3565);
or U8732 (N_8732,N_3596,N_5813);
nand U8733 (N_8733,N_5867,N_4061);
or U8734 (N_8734,N_5690,N_5012);
xnor U8735 (N_8735,N_5035,N_3726);
nor U8736 (N_8736,N_3572,N_5710);
nand U8737 (N_8737,N_4052,N_5114);
nand U8738 (N_8738,N_3685,N_4796);
or U8739 (N_8739,N_4413,N_4088);
xor U8740 (N_8740,N_4122,N_5940);
nand U8741 (N_8741,N_4613,N_4545);
nand U8742 (N_8742,N_3689,N_4730);
or U8743 (N_8743,N_4825,N_5497);
nand U8744 (N_8744,N_5250,N_3887);
xor U8745 (N_8745,N_3908,N_5483);
and U8746 (N_8746,N_5917,N_4926);
nor U8747 (N_8747,N_4029,N_3804);
xor U8748 (N_8748,N_3773,N_5115);
or U8749 (N_8749,N_3831,N_3433);
nand U8750 (N_8750,N_4629,N_5378);
nand U8751 (N_8751,N_4446,N_5472);
and U8752 (N_8752,N_5150,N_4841);
or U8753 (N_8753,N_5122,N_3623);
and U8754 (N_8754,N_3304,N_4032);
nand U8755 (N_8755,N_4410,N_4404);
or U8756 (N_8756,N_4999,N_3754);
or U8757 (N_8757,N_4129,N_5686);
or U8758 (N_8758,N_5411,N_3023);
xnor U8759 (N_8759,N_3708,N_5189);
or U8760 (N_8760,N_5767,N_4558);
or U8761 (N_8761,N_4772,N_3839);
and U8762 (N_8762,N_4460,N_4442);
and U8763 (N_8763,N_3543,N_5607);
nand U8764 (N_8764,N_4610,N_3025);
nand U8765 (N_8765,N_4576,N_5354);
and U8766 (N_8766,N_4676,N_5816);
or U8767 (N_8767,N_3059,N_4238);
or U8768 (N_8768,N_5878,N_5433);
or U8769 (N_8769,N_4810,N_5039);
or U8770 (N_8770,N_3916,N_3802);
nand U8771 (N_8771,N_5888,N_3855);
xnor U8772 (N_8772,N_4192,N_5598);
or U8773 (N_8773,N_5683,N_3139);
nand U8774 (N_8774,N_5647,N_3896);
and U8775 (N_8775,N_5695,N_5859);
or U8776 (N_8776,N_5155,N_3530);
and U8777 (N_8777,N_5753,N_5199);
or U8778 (N_8778,N_5408,N_3745);
and U8779 (N_8779,N_5486,N_4574);
nand U8780 (N_8780,N_4130,N_4359);
nand U8781 (N_8781,N_3021,N_4249);
nor U8782 (N_8782,N_5436,N_5601);
and U8783 (N_8783,N_4301,N_4296);
and U8784 (N_8784,N_4113,N_5010);
nand U8785 (N_8785,N_4526,N_3605);
or U8786 (N_8786,N_3967,N_3797);
or U8787 (N_8787,N_4727,N_3335);
nor U8788 (N_8788,N_5085,N_3160);
nand U8789 (N_8789,N_4168,N_5759);
nand U8790 (N_8790,N_5403,N_4842);
nand U8791 (N_8791,N_5296,N_5629);
and U8792 (N_8792,N_3360,N_4039);
nor U8793 (N_8793,N_5659,N_5170);
nand U8794 (N_8794,N_5838,N_5831);
nor U8795 (N_8795,N_5831,N_3960);
nand U8796 (N_8796,N_4900,N_5403);
nand U8797 (N_8797,N_5475,N_5746);
or U8798 (N_8798,N_4695,N_3586);
nor U8799 (N_8799,N_3491,N_5918);
nor U8800 (N_8800,N_5923,N_4361);
or U8801 (N_8801,N_5078,N_3625);
and U8802 (N_8802,N_3327,N_3267);
xnor U8803 (N_8803,N_4561,N_3075);
nand U8804 (N_8804,N_5359,N_4020);
nor U8805 (N_8805,N_4777,N_5467);
or U8806 (N_8806,N_3388,N_4366);
nor U8807 (N_8807,N_5428,N_5361);
and U8808 (N_8808,N_5919,N_3137);
and U8809 (N_8809,N_3065,N_4289);
nand U8810 (N_8810,N_5046,N_3900);
xor U8811 (N_8811,N_4111,N_5409);
nand U8812 (N_8812,N_4702,N_4739);
or U8813 (N_8813,N_5260,N_5559);
nor U8814 (N_8814,N_5401,N_3420);
nor U8815 (N_8815,N_4268,N_4983);
nor U8816 (N_8816,N_5909,N_3363);
or U8817 (N_8817,N_3945,N_5922);
and U8818 (N_8818,N_5077,N_5016);
xor U8819 (N_8819,N_3748,N_5172);
xor U8820 (N_8820,N_4328,N_3086);
and U8821 (N_8821,N_4973,N_3374);
nor U8822 (N_8822,N_4721,N_5116);
nand U8823 (N_8823,N_5149,N_4789);
nand U8824 (N_8824,N_5265,N_4248);
nand U8825 (N_8825,N_3010,N_4860);
nand U8826 (N_8826,N_4701,N_3089);
xnor U8827 (N_8827,N_3220,N_5045);
nor U8828 (N_8828,N_3971,N_4200);
or U8829 (N_8829,N_4911,N_4342);
or U8830 (N_8830,N_3274,N_4685);
nand U8831 (N_8831,N_3672,N_4050);
nand U8832 (N_8832,N_4783,N_5963);
xor U8833 (N_8833,N_3109,N_3974);
xor U8834 (N_8834,N_5909,N_4537);
and U8835 (N_8835,N_3088,N_5880);
or U8836 (N_8836,N_3322,N_4901);
xor U8837 (N_8837,N_5741,N_5823);
nor U8838 (N_8838,N_3446,N_4256);
nand U8839 (N_8839,N_3575,N_3806);
or U8840 (N_8840,N_4442,N_4081);
nor U8841 (N_8841,N_4025,N_5035);
or U8842 (N_8842,N_3863,N_4327);
xnor U8843 (N_8843,N_5832,N_3274);
nand U8844 (N_8844,N_5000,N_4514);
or U8845 (N_8845,N_5408,N_4682);
nor U8846 (N_8846,N_5177,N_5926);
and U8847 (N_8847,N_3077,N_5701);
nor U8848 (N_8848,N_4437,N_4624);
or U8849 (N_8849,N_3072,N_3493);
and U8850 (N_8850,N_3184,N_3819);
nand U8851 (N_8851,N_4042,N_5529);
nand U8852 (N_8852,N_5530,N_4240);
and U8853 (N_8853,N_5418,N_5972);
nor U8854 (N_8854,N_5536,N_3307);
or U8855 (N_8855,N_5022,N_3129);
nor U8856 (N_8856,N_5754,N_3947);
or U8857 (N_8857,N_4985,N_4368);
and U8858 (N_8858,N_5106,N_3273);
nor U8859 (N_8859,N_4004,N_5116);
nand U8860 (N_8860,N_5811,N_3675);
or U8861 (N_8861,N_4062,N_4520);
nand U8862 (N_8862,N_5283,N_4177);
nand U8863 (N_8863,N_3677,N_3076);
and U8864 (N_8864,N_5845,N_5378);
or U8865 (N_8865,N_3592,N_3351);
nand U8866 (N_8866,N_4852,N_4197);
nand U8867 (N_8867,N_4525,N_3760);
and U8868 (N_8868,N_4002,N_5397);
or U8869 (N_8869,N_4245,N_5880);
or U8870 (N_8870,N_4672,N_3686);
and U8871 (N_8871,N_4145,N_4489);
xor U8872 (N_8872,N_3568,N_4129);
nor U8873 (N_8873,N_3583,N_4249);
xnor U8874 (N_8874,N_4270,N_3618);
or U8875 (N_8875,N_5698,N_4830);
or U8876 (N_8876,N_3908,N_3603);
nand U8877 (N_8877,N_4704,N_4038);
nand U8878 (N_8878,N_4293,N_5828);
nor U8879 (N_8879,N_3099,N_4007);
nand U8880 (N_8880,N_5215,N_3431);
nand U8881 (N_8881,N_3901,N_3156);
and U8882 (N_8882,N_3850,N_3789);
nor U8883 (N_8883,N_3730,N_5860);
or U8884 (N_8884,N_5404,N_3610);
nand U8885 (N_8885,N_4256,N_5894);
nand U8886 (N_8886,N_4841,N_3877);
nor U8887 (N_8887,N_4868,N_4816);
nand U8888 (N_8888,N_5174,N_3500);
xnor U8889 (N_8889,N_4245,N_5734);
or U8890 (N_8890,N_4591,N_5486);
and U8891 (N_8891,N_5918,N_5526);
nor U8892 (N_8892,N_5063,N_5231);
nand U8893 (N_8893,N_3613,N_5328);
nand U8894 (N_8894,N_4082,N_3316);
nor U8895 (N_8895,N_5240,N_3580);
nor U8896 (N_8896,N_4511,N_5543);
nor U8897 (N_8897,N_5309,N_4440);
nor U8898 (N_8898,N_3207,N_5983);
nand U8899 (N_8899,N_4465,N_5040);
nand U8900 (N_8900,N_4040,N_3799);
and U8901 (N_8901,N_4403,N_5051);
nor U8902 (N_8902,N_5845,N_3073);
and U8903 (N_8903,N_5179,N_5429);
and U8904 (N_8904,N_3098,N_5126);
xor U8905 (N_8905,N_4522,N_4877);
nor U8906 (N_8906,N_5836,N_3129);
and U8907 (N_8907,N_4920,N_5958);
and U8908 (N_8908,N_4999,N_4456);
or U8909 (N_8909,N_3804,N_3097);
and U8910 (N_8910,N_3479,N_3653);
xor U8911 (N_8911,N_4782,N_4310);
nor U8912 (N_8912,N_3674,N_5845);
or U8913 (N_8913,N_4574,N_4949);
xnor U8914 (N_8914,N_4745,N_3372);
nand U8915 (N_8915,N_3231,N_5038);
and U8916 (N_8916,N_3366,N_4316);
nand U8917 (N_8917,N_3928,N_3071);
or U8918 (N_8918,N_3165,N_4245);
or U8919 (N_8919,N_4663,N_3663);
nand U8920 (N_8920,N_4396,N_3951);
nand U8921 (N_8921,N_3714,N_4361);
nand U8922 (N_8922,N_4959,N_4734);
nand U8923 (N_8923,N_4048,N_4182);
and U8924 (N_8924,N_3615,N_3080);
and U8925 (N_8925,N_4785,N_4763);
and U8926 (N_8926,N_3919,N_3835);
nor U8927 (N_8927,N_5901,N_4776);
or U8928 (N_8928,N_3573,N_4009);
nand U8929 (N_8929,N_4633,N_4802);
and U8930 (N_8930,N_4825,N_5011);
nand U8931 (N_8931,N_3294,N_5999);
or U8932 (N_8932,N_3931,N_3110);
and U8933 (N_8933,N_4272,N_3765);
nor U8934 (N_8934,N_3944,N_3210);
or U8935 (N_8935,N_4186,N_4610);
nor U8936 (N_8936,N_5909,N_4008);
and U8937 (N_8937,N_3318,N_5853);
or U8938 (N_8938,N_3327,N_3425);
or U8939 (N_8939,N_3296,N_4467);
or U8940 (N_8940,N_3324,N_4677);
or U8941 (N_8941,N_4142,N_4593);
xor U8942 (N_8942,N_4497,N_5192);
and U8943 (N_8943,N_4308,N_3466);
and U8944 (N_8944,N_4280,N_4585);
nor U8945 (N_8945,N_4615,N_4158);
nor U8946 (N_8946,N_5486,N_5727);
nor U8947 (N_8947,N_3684,N_4087);
and U8948 (N_8948,N_3243,N_4156);
xor U8949 (N_8949,N_4301,N_5305);
xnor U8950 (N_8950,N_5126,N_5290);
and U8951 (N_8951,N_4921,N_3426);
nand U8952 (N_8952,N_4225,N_4190);
nand U8953 (N_8953,N_3191,N_3150);
or U8954 (N_8954,N_3606,N_3477);
or U8955 (N_8955,N_4290,N_5420);
and U8956 (N_8956,N_5573,N_3885);
and U8957 (N_8957,N_5103,N_3640);
or U8958 (N_8958,N_4351,N_3250);
nand U8959 (N_8959,N_4063,N_4038);
nand U8960 (N_8960,N_3252,N_4186);
or U8961 (N_8961,N_3932,N_3626);
or U8962 (N_8962,N_3860,N_3803);
nor U8963 (N_8963,N_4925,N_5659);
nand U8964 (N_8964,N_3763,N_5717);
nand U8965 (N_8965,N_4029,N_4688);
or U8966 (N_8966,N_3211,N_3802);
nor U8967 (N_8967,N_4520,N_5417);
nor U8968 (N_8968,N_3261,N_4449);
and U8969 (N_8969,N_5998,N_4362);
and U8970 (N_8970,N_5694,N_3728);
nor U8971 (N_8971,N_4232,N_4673);
or U8972 (N_8972,N_3473,N_3325);
nand U8973 (N_8973,N_4693,N_4902);
xnor U8974 (N_8974,N_5255,N_3483);
nand U8975 (N_8975,N_4395,N_5045);
nand U8976 (N_8976,N_5387,N_4692);
or U8977 (N_8977,N_5219,N_4849);
and U8978 (N_8978,N_3138,N_5968);
nand U8979 (N_8979,N_3743,N_4756);
and U8980 (N_8980,N_5335,N_3960);
or U8981 (N_8981,N_3976,N_5161);
nor U8982 (N_8982,N_4882,N_5868);
and U8983 (N_8983,N_3661,N_4728);
and U8984 (N_8984,N_5526,N_3854);
nor U8985 (N_8985,N_4159,N_5937);
nor U8986 (N_8986,N_5636,N_5273);
nand U8987 (N_8987,N_4206,N_4509);
or U8988 (N_8988,N_4606,N_4557);
or U8989 (N_8989,N_4370,N_4701);
nand U8990 (N_8990,N_4218,N_3421);
nand U8991 (N_8991,N_3639,N_3935);
and U8992 (N_8992,N_3821,N_3085);
or U8993 (N_8993,N_4911,N_4774);
nor U8994 (N_8994,N_4247,N_5621);
nor U8995 (N_8995,N_3939,N_5482);
or U8996 (N_8996,N_4635,N_3798);
nand U8997 (N_8997,N_5901,N_4542);
nand U8998 (N_8998,N_3189,N_5490);
or U8999 (N_8999,N_4805,N_4542);
or U9000 (N_9000,N_7637,N_8474);
xor U9001 (N_9001,N_6374,N_6066);
or U9002 (N_9002,N_7909,N_7609);
and U9003 (N_9003,N_7611,N_8948);
xor U9004 (N_9004,N_8311,N_7123);
or U9005 (N_9005,N_6270,N_6562);
nor U9006 (N_9006,N_8512,N_6576);
or U9007 (N_9007,N_7107,N_6225);
nand U9008 (N_9008,N_7529,N_6676);
nand U9009 (N_9009,N_7744,N_6854);
nor U9010 (N_9010,N_7563,N_6983);
and U9011 (N_9011,N_6406,N_6951);
or U9012 (N_9012,N_7935,N_8825);
and U9013 (N_9013,N_7135,N_7568);
xnor U9014 (N_9014,N_7493,N_7495);
and U9015 (N_9015,N_8359,N_7442);
or U9016 (N_9016,N_8463,N_7371);
or U9017 (N_9017,N_6131,N_6026);
nand U9018 (N_9018,N_7031,N_8953);
nor U9019 (N_9019,N_8529,N_6319);
and U9020 (N_9020,N_8244,N_7046);
nand U9021 (N_9021,N_8853,N_6185);
and U9022 (N_9022,N_6766,N_8972);
nor U9023 (N_9023,N_8274,N_8920);
nand U9024 (N_9024,N_7116,N_6070);
nand U9025 (N_9025,N_7569,N_7004);
xor U9026 (N_9026,N_6559,N_7966);
nand U9027 (N_9027,N_8331,N_6715);
and U9028 (N_9028,N_7625,N_7772);
nor U9029 (N_9029,N_6347,N_8636);
or U9030 (N_9030,N_7931,N_8802);
nand U9031 (N_9031,N_7692,N_6060);
nor U9032 (N_9032,N_7296,N_7986);
and U9033 (N_9033,N_7267,N_7087);
or U9034 (N_9034,N_8880,N_7617);
nand U9035 (N_9035,N_6965,N_7794);
nor U9036 (N_9036,N_7205,N_7958);
nor U9037 (N_9037,N_8049,N_6310);
and U9038 (N_9038,N_8374,N_8727);
nor U9039 (N_9039,N_7142,N_7034);
nor U9040 (N_9040,N_6897,N_6710);
nand U9041 (N_9041,N_6541,N_8392);
and U9042 (N_9042,N_7300,N_6474);
and U9043 (N_9043,N_7159,N_7051);
xor U9044 (N_9044,N_6181,N_8319);
nand U9045 (N_9045,N_6111,N_6115);
and U9046 (N_9046,N_6706,N_6714);
or U9047 (N_9047,N_6915,N_6527);
nand U9048 (N_9048,N_6617,N_6738);
or U9049 (N_9049,N_8170,N_7638);
or U9050 (N_9050,N_6537,N_8764);
or U9051 (N_9051,N_8364,N_7843);
or U9052 (N_9052,N_6076,N_7012);
and U9053 (N_9053,N_6037,N_6062);
or U9054 (N_9054,N_7791,N_7539);
nor U9055 (N_9055,N_8224,N_6348);
nor U9056 (N_9056,N_7021,N_7596);
nor U9057 (N_9057,N_6450,N_6875);
nand U9058 (N_9058,N_6979,N_7374);
xnor U9059 (N_9059,N_6728,N_6466);
or U9060 (N_9060,N_6036,N_8255);
and U9061 (N_9061,N_7335,N_8423);
or U9062 (N_9062,N_8669,N_6762);
or U9063 (N_9063,N_8603,N_8234);
and U9064 (N_9064,N_6914,N_7647);
and U9065 (N_9065,N_8609,N_8232);
and U9066 (N_9066,N_8175,N_7740);
xnor U9067 (N_9067,N_8222,N_8733);
xor U9068 (N_9068,N_6521,N_8496);
and U9069 (N_9069,N_7188,N_6815);
nor U9070 (N_9070,N_7818,N_6067);
or U9071 (N_9071,N_8441,N_7122);
or U9072 (N_9072,N_8363,N_7304);
or U9073 (N_9073,N_6819,N_6910);
nor U9074 (N_9074,N_8054,N_8765);
and U9075 (N_9075,N_8469,N_7944);
xnor U9076 (N_9076,N_7349,N_8079);
or U9077 (N_9077,N_7786,N_7000);
and U9078 (N_9078,N_7472,N_7429);
and U9079 (N_9079,N_6707,N_7410);
and U9080 (N_9080,N_6152,N_6250);
and U9081 (N_9081,N_6911,N_6280);
and U9082 (N_9082,N_6969,N_6780);
and U9083 (N_9083,N_6497,N_8070);
nand U9084 (N_9084,N_8811,N_7286);
nand U9085 (N_9085,N_8554,N_7242);
nand U9086 (N_9086,N_7646,N_8347);
and U9087 (N_9087,N_6774,N_6948);
nor U9088 (N_9088,N_7910,N_6156);
nor U9089 (N_9089,N_7862,N_7392);
and U9090 (N_9090,N_7573,N_8048);
and U9091 (N_9091,N_6602,N_7126);
nor U9092 (N_9092,N_7311,N_7496);
and U9093 (N_9093,N_6653,N_8389);
nand U9094 (N_9094,N_8277,N_8318);
nor U9095 (N_9095,N_8623,N_8421);
and U9096 (N_9096,N_6256,N_8412);
nand U9097 (N_9097,N_7578,N_6960);
nor U9098 (N_9098,N_8998,N_6629);
and U9099 (N_9099,N_8295,N_6545);
nand U9100 (N_9100,N_8415,N_7247);
nand U9101 (N_9101,N_8835,N_8883);
nor U9102 (N_9102,N_7849,N_7704);
nand U9103 (N_9103,N_7831,N_6028);
nand U9104 (N_9104,N_8982,N_8522);
nor U9105 (N_9105,N_8160,N_7451);
nor U9106 (N_9106,N_8029,N_6229);
and U9107 (N_9107,N_8367,N_8176);
nor U9108 (N_9108,N_7788,N_8707);
and U9109 (N_9109,N_8622,N_6486);
and U9110 (N_9110,N_8466,N_7198);
or U9111 (N_9111,N_8887,N_7597);
or U9112 (N_9112,N_6294,N_6534);
nand U9113 (N_9113,N_7134,N_7968);
nor U9114 (N_9114,N_6320,N_6144);
and U9115 (N_9115,N_8133,N_6592);
or U9116 (N_9116,N_7945,N_7390);
or U9117 (N_9117,N_6317,N_6243);
xnor U9118 (N_9118,N_8738,N_7722);
or U9119 (N_9119,N_6913,N_6402);
xor U9120 (N_9120,N_8040,N_8111);
or U9121 (N_9121,N_6981,N_7708);
and U9122 (N_9122,N_8523,N_7081);
and U9123 (N_9123,N_6061,N_8718);
nor U9124 (N_9124,N_6956,N_6831);
and U9125 (N_9125,N_7439,N_8292);
and U9126 (N_9126,N_7640,N_6438);
and U9127 (N_9127,N_7725,N_8492);
or U9128 (N_9128,N_6560,N_7858);
nor U9129 (N_9129,N_7797,N_8071);
and U9130 (N_9130,N_7467,N_7151);
and U9131 (N_9131,N_6895,N_7867);
or U9132 (N_9132,N_6014,N_8671);
nor U9133 (N_9133,N_7995,N_8140);
xor U9134 (N_9134,N_6891,N_6380);
and U9135 (N_9135,N_8650,N_8524);
and U9136 (N_9136,N_8684,N_6172);
or U9137 (N_9137,N_7604,N_8033);
nand U9138 (N_9138,N_6069,N_7255);
nor U9139 (N_9139,N_8407,N_7693);
nand U9140 (N_9140,N_8985,N_7307);
nand U9141 (N_9141,N_8266,N_8116);
or U9142 (N_9142,N_7076,N_7068);
nor U9143 (N_9143,N_8674,N_6709);
and U9144 (N_9144,N_6868,N_8987);
and U9145 (N_9145,N_7354,N_6202);
nor U9146 (N_9146,N_6599,N_7908);
or U9147 (N_9147,N_7847,N_7431);
nand U9148 (N_9148,N_7922,N_6395);
or U9149 (N_9149,N_7803,N_6551);
and U9150 (N_9150,N_8023,N_8775);
nand U9151 (N_9151,N_7508,N_8180);
nand U9152 (N_9152,N_8283,N_8500);
nor U9153 (N_9153,N_8246,N_6323);
and U9154 (N_9154,N_6690,N_7854);
nor U9155 (N_9155,N_8997,N_7943);
nand U9156 (N_9156,N_6928,N_7887);
and U9157 (N_9157,N_7395,N_6168);
nand U9158 (N_9158,N_8344,N_7070);
nand U9159 (N_9159,N_6946,N_6845);
and U9160 (N_9160,N_6110,N_6341);
nand U9161 (N_9161,N_8369,N_6385);
nor U9162 (N_9162,N_7651,N_7372);
or U9163 (N_9163,N_6700,N_6329);
and U9164 (N_9164,N_8399,N_8753);
nor U9165 (N_9165,N_6673,N_6113);
nand U9166 (N_9166,N_7037,N_6253);
or U9167 (N_9167,N_8911,N_8627);
nor U9168 (N_9168,N_7144,N_6730);
nor U9169 (N_9169,N_7920,N_7874);
xnor U9170 (N_9170,N_6839,N_7119);
nand U9171 (N_9171,N_8156,N_8725);
nand U9172 (N_9172,N_7627,N_8453);
and U9173 (N_9173,N_7621,N_6898);
or U9174 (N_9174,N_7710,N_6887);
xor U9175 (N_9175,N_6102,N_8538);
nor U9176 (N_9176,N_7701,N_6972);
and U9177 (N_9177,N_7005,N_6099);
nand U9178 (N_9178,N_6890,N_8386);
or U9179 (N_9179,N_6638,N_7677);
and U9180 (N_9180,N_6355,N_6488);
and U9181 (N_9181,N_8205,N_6412);
xnor U9182 (N_9182,N_8947,N_8580);
and U9183 (N_9183,N_8268,N_6779);
nor U9184 (N_9184,N_7320,N_6570);
and U9185 (N_9185,N_6192,N_6727);
xnor U9186 (N_9186,N_6127,N_7518);
nor U9187 (N_9187,N_6169,N_7036);
xor U9188 (N_9188,N_8105,N_7895);
or U9189 (N_9189,N_8709,N_7891);
or U9190 (N_9190,N_7077,N_6025);
nand U9191 (N_9191,N_6574,N_8456);
nor U9192 (N_9192,N_6659,N_6975);
or U9193 (N_9193,N_6086,N_8867);
nor U9194 (N_9194,N_7662,N_7544);
or U9195 (N_9195,N_8414,N_6164);
nand U9196 (N_9196,N_6642,N_6246);
or U9197 (N_9197,N_7057,N_6342);
and U9198 (N_9198,N_7393,N_8831);
or U9199 (N_9199,N_7266,N_8759);
nor U9200 (N_9200,N_6368,N_8562);
nor U9201 (N_9201,N_7757,N_8711);
xor U9202 (N_9202,N_7750,N_8448);
and U9203 (N_9203,N_7681,N_8434);
or U9204 (N_9204,N_7301,N_8652);
and U9205 (N_9205,N_6454,N_6394);
or U9206 (N_9206,N_7288,N_6324);
and U9207 (N_9207,N_7305,N_6382);
or U9208 (N_9208,N_7700,N_7804);
and U9209 (N_9209,N_8696,N_6286);
and U9210 (N_9210,N_7089,N_6096);
xnor U9211 (N_9211,N_7167,N_6524);
nor U9212 (N_9212,N_6615,N_8132);
or U9213 (N_9213,N_6188,N_8281);
and U9214 (N_9214,N_8939,N_7822);
or U9215 (N_9215,N_8868,N_7515);
nor U9216 (N_9216,N_6487,N_6332);
nor U9217 (N_9217,N_8022,N_7033);
nor U9218 (N_9218,N_6105,N_6702);
xnor U9219 (N_9219,N_8158,N_7732);
and U9220 (N_9220,N_7618,N_7869);
nor U9221 (N_9221,N_6484,N_8698);
and U9222 (N_9222,N_6974,N_6558);
xnor U9223 (N_9223,N_7537,N_6456);
and U9224 (N_9224,N_8648,N_8061);
or U9225 (N_9225,N_8573,N_6939);
nor U9226 (N_9226,N_6589,N_8422);
xor U9227 (N_9227,N_6704,N_7685);
nor U9228 (N_9228,N_6808,N_8944);
nand U9229 (N_9229,N_7739,N_8167);
or U9230 (N_9230,N_6451,N_6107);
and U9231 (N_9231,N_7180,N_8280);
nor U9232 (N_9232,N_7904,N_8642);
nand U9233 (N_9233,N_7752,N_7222);
nor U9234 (N_9234,N_6353,N_8619);
or U9235 (N_9235,N_8537,N_6040);
or U9236 (N_9236,N_7003,N_6718);
nor U9237 (N_9237,N_8781,N_6716);
nand U9238 (N_9238,N_8613,N_6360);
nand U9239 (N_9239,N_8437,N_7616);
nor U9240 (N_9240,N_6849,N_7083);
and U9241 (N_9241,N_6518,N_6473);
nor U9242 (N_9242,N_7202,N_7237);
nand U9243 (N_9243,N_8308,N_6609);
and U9244 (N_9244,N_7094,N_8478);
nand U9245 (N_9245,N_6255,N_6556);
and U9246 (N_9246,N_7714,N_8506);
or U9247 (N_9247,N_8690,N_6407);
and U9248 (N_9248,N_6398,N_6325);
nor U9249 (N_9249,N_8772,N_7405);
nand U9250 (N_9250,N_6649,N_6482);
or U9251 (N_9251,N_8417,N_6549);
nand U9252 (N_9252,N_7868,N_6240);
and U9253 (N_9253,N_7498,N_7800);
and U9254 (N_9254,N_8035,N_8249);
nor U9255 (N_9255,N_7998,N_6747);
or U9256 (N_9256,N_8226,N_7324);
nor U9257 (N_9257,N_6145,N_6088);
nor U9258 (N_9258,N_6000,N_7989);
and U9259 (N_9259,N_7181,N_8313);
or U9260 (N_9260,N_6749,N_8429);
and U9261 (N_9261,N_7705,N_8575);
xor U9262 (N_9262,N_6616,N_6433);
nor U9263 (N_9263,N_8881,N_6300);
nor U9264 (N_9264,N_7019,N_7901);
nand U9265 (N_9265,N_8844,N_8686);
xor U9266 (N_9266,N_6532,N_6803);
nor U9267 (N_9267,N_8307,N_8872);
or U9268 (N_9268,N_6198,N_8024);
and U9269 (N_9269,N_6583,N_7303);
nand U9270 (N_9270,N_8015,N_6400);
nor U9271 (N_9271,N_7576,N_7052);
nor U9272 (N_9272,N_8726,N_8976);
and U9273 (N_9273,N_6483,N_6163);
nor U9274 (N_9274,N_8768,N_8897);
nand U9275 (N_9275,N_6798,N_8967);
nor U9276 (N_9276,N_8168,N_7548);
xor U9277 (N_9277,N_7661,N_6542);
or U9278 (N_9278,N_6778,N_6994);
nor U9279 (N_9279,N_8842,N_7587);
and U9280 (N_9280,N_6177,N_7834);
nor U9281 (N_9281,N_6947,N_8873);
nor U9282 (N_9282,N_6628,N_7355);
or U9283 (N_9283,N_7519,N_8233);
and U9284 (N_9284,N_7022,N_7907);
or U9285 (N_9285,N_6650,N_8254);
nor U9286 (N_9286,N_8957,N_7026);
or U9287 (N_9287,N_8092,N_8017);
nor U9288 (N_9288,N_7864,N_8008);
or U9289 (N_9289,N_6695,N_8321);
or U9290 (N_9290,N_7738,N_7369);
nor U9291 (N_9291,N_6162,N_6889);
or U9292 (N_9292,N_8253,N_7359);
and U9293 (N_9293,N_7105,N_6907);
or U9294 (N_9294,N_7482,N_8635);
xor U9295 (N_9295,N_6987,N_8950);
xnor U9296 (N_9296,N_8005,N_6731);
or U9297 (N_9297,N_7733,N_7447);
xnor U9298 (N_9298,N_8826,N_7509);
nor U9299 (N_9299,N_6414,N_6885);
xor U9300 (N_9300,N_7204,N_6646);
nand U9301 (N_9301,N_6752,N_7614);
nand U9302 (N_9302,N_6667,N_7201);
nor U9303 (N_9303,N_8827,N_8815);
or U9304 (N_9304,N_6800,N_8212);
and U9305 (N_9305,N_8541,N_6927);
or U9306 (N_9306,N_8425,N_8739);
nand U9307 (N_9307,N_8142,N_7659);
xnor U9308 (N_9308,N_6905,N_8191);
or U9309 (N_9309,N_6278,N_6830);
and U9310 (N_9310,N_7812,N_7913);
nor U9311 (N_9311,N_6500,N_8403);
nor U9312 (N_9312,N_8761,N_7457);
and U9313 (N_9313,N_8218,N_6684);
nor U9314 (N_9314,N_6984,N_8213);
and U9315 (N_9315,N_7902,N_8370);
and U9316 (N_9316,N_8202,N_7168);
or U9317 (N_9317,N_6813,N_6698);
nand U9318 (N_9318,N_8447,N_8964);
nor U9319 (N_9319,N_7761,N_8720);
nor U9320 (N_9320,N_6807,N_8498);
nand U9321 (N_9321,N_7063,N_6783);
or U9322 (N_9322,N_7145,N_6043);
and U9323 (N_9323,N_6477,N_6926);
nand U9324 (N_9324,N_8334,N_8539);
nand U9325 (N_9325,N_7860,N_8381);
nand U9326 (N_9326,N_8187,N_7178);
xor U9327 (N_9327,N_7555,N_6788);
nor U9328 (N_9328,N_7054,N_7279);
nand U9329 (N_9329,N_8293,N_8128);
nand U9330 (N_9330,N_8969,N_6193);
nand U9331 (N_9331,N_8892,N_8395);
nand U9332 (N_9332,N_6045,N_6242);
and U9333 (N_9333,N_7877,N_8058);
and U9334 (N_9334,N_8763,N_7631);
or U9335 (N_9335,N_8977,N_8130);
and U9336 (N_9336,N_8305,N_8662);
nor U9337 (N_9337,N_6520,N_8896);
and U9338 (N_9338,N_7602,N_7656);
or U9339 (N_9339,N_7848,N_6787);
or U9340 (N_9340,N_8596,N_8760);
nor U9341 (N_9341,N_6753,N_8545);
or U9342 (N_9342,N_8699,N_8221);
or U9343 (N_9343,N_7308,N_6266);
or U9344 (N_9344,N_8332,N_7792);
and U9345 (N_9345,N_8306,N_6670);
nor U9346 (N_9346,N_7485,N_6430);
and U9347 (N_9347,N_6178,N_8150);
or U9348 (N_9348,N_7810,N_8647);
and U9349 (N_9349,N_7483,N_7436);
xnor U9350 (N_9350,N_8960,N_7041);
or U9351 (N_9351,N_6619,N_8779);
nor U9352 (N_9352,N_8602,N_8701);
nor U9353 (N_9353,N_6781,N_6717);
nand U9354 (N_9354,N_6786,N_6767);
or U9355 (N_9355,N_8929,N_8518);
or U9356 (N_9356,N_6033,N_8558);
or U9357 (N_9357,N_7771,N_7718);
and U9358 (N_9358,N_7892,N_8258);
nand U9359 (N_9359,N_6623,N_8104);
and U9360 (N_9360,N_7673,N_7969);
nand U9361 (N_9361,N_8304,N_8080);
and U9362 (N_9362,N_8703,N_8225);
nor U9363 (N_9363,N_8161,N_7292);
or U9364 (N_9364,N_7558,N_7153);
nor U9365 (N_9365,N_8550,N_8819);
xor U9366 (N_9366,N_7861,N_8430);
and U9367 (N_9367,N_6452,N_8965);
xnor U9368 (N_9368,N_6909,N_8649);
and U9369 (N_9369,N_7253,N_8491);
and U9370 (N_9370,N_7010,N_8876);
nor U9371 (N_9371,N_6572,N_8438);
and U9372 (N_9372,N_8519,N_7776);
and U9373 (N_9373,N_8385,N_7104);
or U9374 (N_9374,N_6034,N_8816);
or U9375 (N_9375,N_7668,N_8074);
and U9376 (N_9376,N_8444,N_7608);
and U9377 (N_9377,N_6721,N_8584);
and U9378 (N_9378,N_8504,N_8617);
and U9379 (N_9379,N_6581,N_6600);
nand U9380 (N_9380,N_7574,N_7327);
xor U9381 (N_9381,N_8410,N_7873);
xnor U9382 (N_9382,N_7663,N_6460);
or U9383 (N_9383,N_8208,N_8814);
nand U9384 (N_9384,N_8455,N_7566);
and U9385 (N_9385,N_8495,N_8162);
and U9386 (N_9386,N_6298,N_6647);
xor U9387 (N_9387,N_8664,N_7851);
nand U9388 (N_9388,N_6964,N_7013);
nand U9389 (N_9389,N_6265,N_6227);
nor U9390 (N_9390,N_8078,N_8793);
nor U9391 (N_9391,N_6679,N_8296);
nand U9392 (N_9392,N_8570,N_6331);
nand U9393 (N_9393,N_7978,N_7333);
nor U9394 (N_9394,N_8184,N_6967);
or U9395 (N_9395,N_7125,N_7476);
nor U9396 (N_9396,N_7992,N_7884);
or U9397 (N_9397,N_8611,N_6594);
and U9398 (N_9398,N_8863,N_7643);
nor U9399 (N_9399,N_8644,N_6008);
and U9400 (N_9400,N_6285,N_8632);
nor U9401 (N_9401,N_6251,N_6296);
and U9402 (N_9402,N_6904,N_6259);
nor U9403 (N_9403,N_7402,N_6197);
nand U9404 (N_9404,N_6870,N_7543);
xnor U9405 (N_9405,N_6013,N_7993);
nor U9406 (N_9406,N_7127,N_8938);
nand U9407 (N_9407,N_7235,N_6569);
and U9408 (N_9408,N_7406,N_6413);
nand U9409 (N_9409,N_7503,N_7108);
nand U9410 (N_9410,N_8517,N_7918);
xnor U9411 (N_9411,N_7550,N_8204);
nand U9412 (N_9412,N_6495,N_6120);
nor U9413 (N_9413,N_8340,N_6936);
nand U9414 (N_9414,N_6306,N_8065);
or U9415 (N_9415,N_8451,N_8777);
nor U9416 (N_9416,N_6597,N_8688);
and U9417 (N_9417,N_8108,N_8153);
nor U9418 (N_9418,N_6170,N_8267);
or U9419 (N_9419,N_6201,N_8740);
and U9420 (N_9420,N_8203,N_6458);
xor U9421 (N_9421,N_7670,N_6843);
xnor U9422 (N_9422,N_8680,N_7345);
and U9423 (N_9423,N_7613,N_6392);
nor U9424 (N_9424,N_8754,N_6846);
and U9425 (N_9425,N_8245,N_6418);
and U9426 (N_9426,N_7465,N_8728);
nor U9427 (N_9427,N_7919,N_7208);
or U9428 (N_9428,N_6795,N_7844);
nor U9429 (N_9429,N_7513,N_8454);
and U9430 (N_9430,N_7678,N_7979);
nand U9431 (N_9431,N_7743,N_7997);
nor U9432 (N_9432,N_8269,N_6658);
and U9433 (N_9433,N_6632,N_7271);
nand U9434 (N_9434,N_6643,N_6158);
nor U9435 (N_9435,N_7244,N_7841);
nor U9436 (N_9436,N_7764,N_8050);
nor U9437 (N_9437,N_6094,N_6671);
and U9438 (N_9438,N_7580,N_7365);
nor U9439 (N_9439,N_8721,N_7890);
nor U9440 (N_9440,N_7541,N_6504);
and U9441 (N_9441,N_6734,N_7397);
or U9442 (N_9442,N_7455,N_7572);
and U9443 (N_9443,N_7817,N_6136);
nand U9444 (N_9444,N_6379,N_7090);
nand U9445 (N_9445,N_6509,N_8378);
or U9446 (N_9446,N_7148,N_8076);
nand U9447 (N_9447,N_8767,N_8568);
or U9448 (N_9448,N_8732,N_7002);
and U9449 (N_9449,N_8481,N_6384);
xnor U9450 (N_9450,N_8297,N_7099);
nor U9451 (N_9451,N_8067,N_6247);
or U9452 (N_9452,N_6773,N_7309);
or U9453 (N_9453,N_8634,N_6258);
nand U9454 (N_9454,N_7584,N_8633);
or U9455 (N_9455,N_7619,N_6421);
or U9456 (N_9456,N_8082,N_8241);
nand U9457 (N_9457,N_7799,N_6719);
or U9458 (N_9458,N_6239,N_8262);
or U9459 (N_9459,N_6277,N_6814);
and U9460 (N_9460,N_8118,N_6090);
nor U9461 (N_9461,N_7972,N_7575);
nand U9462 (N_9462,N_7401,N_8569);
or U9463 (N_9463,N_7236,N_7835);
xor U9464 (N_9464,N_8081,N_8196);
xnor U9465 (N_9465,N_7672,N_7226);
nand U9466 (N_9466,N_7912,N_7438);
or U9467 (N_9467,N_7071,N_8736);
nand U9468 (N_9468,N_6851,N_8322);
or U9469 (N_9469,N_6003,N_6770);
or U9470 (N_9470,N_7448,N_7006);
nand U9471 (N_9471,N_8354,N_7562);
and U9472 (N_9472,N_7163,N_8682);
nand U9473 (N_9473,N_7737,N_8930);
and U9474 (N_9474,N_8016,N_6333);
nand U9475 (N_9475,N_6917,N_6449);
nand U9476 (N_9476,N_8526,N_6584);
xnor U9477 (N_9477,N_6955,N_7629);
nor U9478 (N_9478,N_7411,N_6977);
and U9479 (N_9479,N_6661,N_7589);
xor U9480 (N_9480,N_6945,N_7106);
xor U9481 (N_9481,N_8810,N_7556);
nor U9482 (N_9482,N_8066,N_8931);
or U9483 (N_9483,N_7828,N_8801);
and U9484 (N_9484,N_7653,N_8265);
or U9485 (N_9485,N_6234,N_7377);
or U9486 (N_9486,N_6848,N_8527);
and U9487 (N_9487,N_6825,N_6287);
nand U9488 (N_9488,N_7437,N_7233);
nand U9489 (N_9489,N_6529,N_6962);
or U9490 (N_9490,N_8486,N_7598);
or U9491 (N_9491,N_6732,N_7581);
nand U9492 (N_9492,N_6055,N_6514);
nand U9493 (N_9493,N_7667,N_7155);
and U9494 (N_9494,N_7420,N_8903);
or U9495 (N_9495,N_8755,N_8937);
or U9496 (N_9496,N_6873,N_7754);
xor U9497 (N_9497,N_6057,N_6047);
xnor U9498 (N_9498,N_8147,N_6245);
nor U9499 (N_9499,N_8788,N_8420);
nor U9500 (N_9500,N_8223,N_6940);
and U9501 (N_9501,N_6303,N_8062);
xor U9502 (N_9502,N_6221,N_8207);
nand U9503 (N_9503,N_7819,N_6146);
xor U9504 (N_9504,N_8004,N_6916);
nor U9505 (N_9505,N_7446,N_7855);
and U9506 (N_9506,N_7723,N_7461);
and U9507 (N_9507,N_6988,N_6089);
or U9508 (N_9508,N_6393,N_6143);
nor U9509 (N_9509,N_6824,N_6063);
nor U9510 (N_9510,N_6388,N_8628);
nand U9511 (N_9511,N_6128,N_8771);
or U9512 (N_9512,N_7994,N_6108);
nor U9513 (N_9513,N_6547,N_7428);
nand U9514 (N_9514,N_7488,N_8194);
nor U9515 (N_9515,N_8762,N_7100);
and U9516 (N_9516,N_6244,N_8343);
xnor U9517 (N_9517,N_6992,N_6109);
nor U9518 (N_9518,N_8502,N_6624);
nor U9519 (N_9519,N_7636,N_8708);
or U9520 (N_9520,N_6376,N_8638);
or U9521 (N_9521,N_6660,N_7762);
and U9522 (N_9522,N_7338,N_8256);
and U9523 (N_9523,N_8121,N_7319);
and U9524 (N_9524,N_6723,N_8551);
nor U9525 (N_9525,N_7779,N_7095);
nand U9526 (N_9526,N_7213,N_7689);
nor U9527 (N_9527,N_7711,N_7480);
nor U9528 (N_9528,N_7312,N_6190);
or U9529 (N_9529,N_8325,N_6363);
and U9530 (N_9530,N_8483,N_7883);
nand U9531 (N_9531,N_6302,N_8019);
or U9532 (N_9532,N_7047,N_6879);
nand U9533 (N_9533,N_7223,N_6444);
nor U9534 (N_9534,N_8031,N_6035);
nand U9535 (N_9535,N_7380,N_7290);
nand U9536 (N_9536,N_6396,N_7375);
and U9537 (N_9537,N_6517,N_7875);
or U9538 (N_9538,N_6598,N_6548);
or U9539 (N_9539,N_8516,N_6339);
and U9540 (N_9540,N_7961,N_7845);
and U9541 (N_9541,N_8587,N_8068);
and U9542 (N_9542,N_6511,N_8719);
nand U9543 (N_9543,N_6351,N_8436);
or U9544 (N_9544,N_6557,N_8287);
or U9545 (N_9545,N_7680,N_7753);
nor U9546 (N_9546,N_8919,N_7284);
xnor U9547 (N_9547,N_8199,N_7326);
nor U9548 (N_9548,N_6344,N_8400);
nor U9549 (N_9549,N_6761,N_7434);
xor U9550 (N_9550,N_6015,N_6457);
nor U9551 (N_9551,N_7749,N_8095);
xor U9552 (N_9552,N_6850,N_7200);
nor U9553 (N_9553,N_8157,N_6575);
nor U9554 (N_9554,N_7024,N_8428);
or U9555 (N_9555,N_8712,N_8188);
and U9556 (N_9556,N_7853,N_8164);
and U9557 (N_9557,N_7540,N_8365);
and U9558 (N_9558,N_7798,N_8852);
nand U9559 (N_9559,N_6217,N_7612);
or U9560 (N_9560,N_6966,N_6565);
and U9561 (N_9561,N_7139,N_8115);
or U9562 (N_9562,N_6536,N_6417);
nor U9563 (N_9563,N_8449,N_8582);
xor U9564 (N_9564,N_6032,N_8694);
xor U9565 (N_9565,N_7664,N_7302);
nand U9566 (N_9566,N_7601,N_6284);
nor U9567 (N_9567,N_7229,N_6903);
nor U9568 (N_9568,N_6080,N_7674);
or U9569 (N_9569,N_6056,N_6493);
xnor U9570 (N_9570,N_7141,N_6510);
and U9571 (N_9571,N_6952,N_6337);
and U9572 (N_9572,N_7219,N_6986);
nor U9573 (N_9573,N_7975,N_8735);
and U9574 (N_9574,N_7720,N_6075);
or U9575 (N_9575,N_7881,N_7721);
nor U9576 (N_9576,N_6970,N_7830);
xor U9577 (N_9577,N_7586,N_7014);
and U9578 (N_9578,N_8171,N_8528);
and U9579 (N_9579,N_8612,N_6501);
nor U9580 (N_9580,N_8607,N_7525);
nand U9581 (N_9581,N_7399,N_7443);
or U9582 (N_9582,N_7261,N_6292);
nand U9583 (N_9583,N_6129,N_8310);
nor U9584 (N_9584,N_7517,N_6626);
or U9585 (N_9585,N_7379,N_6696);
and U9586 (N_9586,N_8484,N_6138);
nand U9587 (N_9587,N_8329,N_7507);
or U9588 (N_9588,N_8402,N_8471);
or U9589 (N_9589,N_7965,N_8705);
nor U9590 (N_9590,N_7527,N_8605);
and U9591 (N_9591,N_8678,N_7058);
nor U9592 (N_9592,N_8843,N_8567);
nand U9593 (N_9593,N_6157,N_8106);
nand U9594 (N_9594,N_6601,N_8264);
nor U9595 (N_9595,N_8794,N_6944);
nor U9596 (N_9596,N_8837,N_7336);
nor U9597 (N_9597,N_7657,N_6648);
or U9598 (N_9598,N_7929,N_7294);
or U9599 (N_9599,N_8056,N_8822);
xnor U9600 (N_9600,N_8494,N_7157);
nor U9601 (N_9601,N_6183,N_6691);
xor U9602 (N_9602,N_7536,N_7486);
nand U9603 (N_9603,N_7387,N_8909);
nor U9604 (N_9604,N_8521,N_7497);
or U9605 (N_9605,N_8510,N_8592);
nand U9606 (N_9606,N_6427,N_7277);
xor U9607 (N_9607,N_6416,N_6869);
and U9608 (N_9608,N_8501,N_8989);
nand U9609 (N_9609,N_8242,N_7759);
nor U9610 (N_9610,N_6805,N_6645);
and U9611 (N_9611,N_6499,N_6463);
nor U9612 (N_9612,N_7973,N_8756);
nand U9613 (N_9613,N_6073,N_7499);
nand U9614 (N_9614,N_8227,N_8675);
or U9615 (N_9615,N_6756,N_8722);
or U9616 (N_9616,N_8914,N_6289);
nor U9617 (N_9617,N_8806,N_8833);
and U9618 (N_9618,N_6279,N_7011);
and U9619 (N_9619,N_6561,N_6415);
nor U9620 (N_9620,N_8915,N_6448);
and U9621 (N_9621,N_7826,N_7252);
nor U9622 (N_9622,N_7020,N_8279);
nor U9623 (N_9623,N_8593,N_8139);
nand U9624 (N_9624,N_6365,N_7130);
and U9625 (N_9625,N_8263,N_7726);
or U9626 (N_9626,N_6001,N_8055);
xor U9627 (N_9627,N_7872,N_6126);
and U9628 (N_9628,N_6858,N_7194);
nor U9629 (N_9629,N_7263,N_8390);
xnor U9630 (N_9630,N_8189,N_6782);
or U9631 (N_9631,N_7214,N_7297);
nor U9632 (N_9632,N_8540,N_6853);
xnor U9633 (N_9633,N_8284,N_8503);
nor U9634 (N_9634,N_8342,N_6215);
or U9635 (N_9635,N_7983,N_6389);
and U9636 (N_9636,N_8588,N_7991);
xor U9637 (N_9637,N_8653,N_8465);
and U9638 (N_9638,N_7866,N_6429);
nor U9639 (N_9639,N_6656,N_6657);
nand U9640 (N_9640,N_8141,N_7293);
or U9641 (N_9641,N_7425,N_7694);
xor U9642 (N_9642,N_8792,N_6993);
or U9643 (N_9643,N_6685,N_6209);
and U9644 (N_9644,N_6216,N_7274);
nand U9645 (N_9645,N_8272,N_8159);
nor U9646 (N_9646,N_8467,N_7040);
or U9647 (N_9647,N_7028,N_8716);
nand U9648 (N_9648,N_8710,N_7025);
and U9649 (N_9649,N_8479,N_6604);
nand U9650 (N_9650,N_6639,N_7709);
or U9651 (N_9651,N_7963,N_8473);
and U9652 (N_9652,N_6122,N_8487);
nor U9653 (N_9653,N_6455,N_7352);
nor U9654 (N_9654,N_8734,N_6856);
nand U9655 (N_9655,N_7430,N_6662);
or U9656 (N_9656,N_8572,N_7914);
nand U9657 (N_9657,N_6124,N_6683);
or U9658 (N_9658,N_6082,N_6613);
or U9659 (N_9659,N_8791,N_7839);
nor U9660 (N_9660,N_8094,N_8770);
and U9661 (N_9661,N_7634,N_7138);
nand U9662 (N_9662,N_8052,N_8685);
or U9663 (N_9663,N_7758,N_6391);
and U9664 (N_9664,N_6857,N_8536);
or U9665 (N_9665,N_8515,N_8276);
and U9666 (N_9666,N_6573,N_8183);
nand U9667 (N_9667,N_7494,N_8884);
and U9668 (N_9668,N_7171,N_8457);
or U9669 (N_9669,N_6874,N_8514);
nor U9670 (N_9670,N_6932,N_6214);
nand U9671 (N_9671,N_7278,N_7343);
or U9672 (N_9672,N_8084,N_8626);
nand U9673 (N_9673,N_8166,N_7129);
and U9674 (N_9674,N_6065,N_6390);
nand U9675 (N_9675,N_6835,N_8145);
and U9676 (N_9676,N_6211,N_7775);
nand U9677 (N_9677,N_6316,N_8912);
xor U9678 (N_9678,N_7137,N_6352);
and U9679 (N_9679,N_7298,N_8758);
nor U9680 (N_9680,N_8275,N_6354);
nand U9681 (N_9681,N_7088,N_7730);
nand U9682 (N_9682,N_8413,N_6912);
or U9683 (N_9683,N_7955,N_8002);
or U9684 (N_9684,N_8011,N_6507);
nor U9685 (N_9685,N_6821,N_8210);
nor U9686 (N_9686,N_6464,N_8442);
nand U9687 (N_9687,N_6268,N_6797);
nand U9688 (N_9688,N_7641,N_8618);
xor U9689 (N_9689,N_6420,N_6544);
nor U9690 (N_9690,N_6768,N_6810);
or U9691 (N_9691,N_6515,N_8149);
or U9692 (N_9692,N_7250,N_6862);
nand U9693 (N_9693,N_8597,N_7269);
nand U9694 (N_9694,N_8531,N_8702);
xnor U9695 (N_9695,N_8489,N_7837);
and U9696 (N_9696,N_8862,N_6362);
or U9697 (N_9697,N_8038,N_7454);
or U9698 (N_9698,N_8746,N_7350);
and U9699 (N_9699,N_6712,N_7532);
xnor U9700 (N_9700,N_6461,N_8625);
or U9701 (N_9701,N_7784,N_7146);
nand U9702 (N_9702,N_7806,N_6585);
and U9703 (N_9703,N_8497,N_6538);
nor U9704 (N_9704,N_6104,N_8829);
nand U9705 (N_9705,N_6078,N_7334);
or U9706 (N_9706,N_7193,N_7166);
and U9707 (N_9707,N_6953,N_6989);
nand U9708 (N_9708,N_6103,N_8988);
nor U9709 (N_9709,N_7676,N_8335);
and U9710 (N_9710,N_6432,N_8173);
and U9711 (N_9711,N_7449,N_8003);
nand U9712 (N_9712,N_6997,N_7796);
or U9713 (N_9713,N_6553,N_8534);
nor U9714 (N_9714,N_7728,N_7964);
and U9715 (N_9715,N_6841,N_8252);
nor U9716 (N_9716,N_6980,N_7259);
nand U9717 (N_9717,N_7840,N_8547);
nand U9718 (N_9718,N_6689,N_6855);
nor U9719 (N_9719,N_6725,N_7546);
xnor U9720 (N_9720,N_8117,N_6777);
nor U9721 (N_9721,N_8114,N_6301);
and U9722 (N_9722,N_6005,N_6182);
and U9723 (N_9723,N_7767,N_8786);
nand U9724 (N_9724,N_7715,N_6522);
nor U9725 (N_9725,N_8294,N_7649);
nand U9726 (N_9726,N_6958,N_8462);
nand U9727 (N_9727,N_7154,N_6754);
or U9728 (N_9728,N_8615,N_7197);
or U9729 (N_9729,N_6220,N_6641);
or U9730 (N_9730,N_8382,N_8571);
or U9731 (N_9731,N_7742,N_8839);
nor U9732 (N_9732,N_6587,N_7342);
nor U9733 (N_9733,N_8847,N_7121);
or U9734 (N_9734,N_8090,N_6167);
or U9735 (N_9735,N_8574,N_6343);
nand U9736 (N_9736,N_6776,N_7489);
or U9737 (N_9737,N_8849,N_6930);
or U9738 (N_9738,N_8559,N_6346);
and U9739 (N_9739,N_6262,N_8656);
and U9740 (N_9740,N_7273,N_8433);
nor U9741 (N_9741,N_8211,N_7976);
and U9742 (N_9742,N_7169,N_8513);
nor U9743 (N_9743,N_8350,N_8888);
or U9744 (N_9744,N_8197,N_7557);
nand U9745 (N_9745,N_8661,N_8243);
nor U9746 (N_9746,N_7504,N_6176);
or U9747 (N_9747,N_7112,N_6785);
or U9748 (N_9748,N_7143,N_7475);
and U9749 (N_9749,N_8553,N_6160);
and U9750 (N_9750,N_8405,N_6410);
or U9751 (N_9751,N_7287,N_8851);
xnor U9752 (N_9752,N_8904,N_6995);
or U9753 (N_9753,N_8046,N_6434);
nand U9754 (N_9754,N_6938,N_8214);
and U9755 (N_9755,N_7825,N_6439);
nor U9756 (N_9756,N_7059,N_6607);
nor U9757 (N_9757,N_7516,N_8916);
and U9758 (N_9758,N_6155,N_6186);
nor U9759 (N_9759,N_7452,N_8352);
nor U9760 (N_9760,N_7652,N_8102);
nor U9761 (N_9761,N_8146,N_8209);
nand U9762 (N_9762,N_6327,N_7412);
or U9763 (N_9763,N_8846,N_8790);
or U9764 (N_9764,N_8778,N_7481);
or U9765 (N_9765,N_8877,N_8122);
and U9766 (N_9766,N_8542,N_8085);
or U9767 (N_9767,N_7727,N_7787);
and U9768 (N_9768,N_7654,N_7948);
nand U9769 (N_9769,N_6503,N_7522);
xnor U9770 (N_9770,N_7418,N_8543);
and U9771 (N_9771,N_6231,N_6100);
or U9772 (N_9772,N_8657,N_8371);
xor U9773 (N_9773,N_8505,N_7773);
nand U9774 (N_9774,N_6675,N_7172);
nor U9775 (N_9775,N_6184,N_8576);
nor U9776 (N_9776,N_6742,N_7785);
nor U9777 (N_9777,N_7769,N_6531);
and U9778 (N_9778,N_6526,N_7199);
nor U9779 (N_9779,N_7221,N_8042);
and U9780 (N_9780,N_6230,N_7067);
and U9781 (N_9781,N_6027,N_6322);
and U9782 (N_9782,N_6882,N_8231);
xor U9783 (N_9783,N_8072,N_8361);
or U9784 (N_9784,N_7600,N_6011);
nor U9785 (N_9785,N_8857,N_6249);
nand U9786 (N_9786,N_8186,N_7176);
xor U9787 (N_9787,N_7258,N_6840);
or U9788 (N_9788,N_6941,N_7623);
nor U9789 (N_9789,N_6282,N_6367);
nor U9790 (N_9790,N_8229,N_6338);
nor U9791 (N_9791,N_7591,N_7682);
and U9792 (N_9792,N_8235,N_8818);
nor U9793 (N_9793,N_8336,N_7366);
and U9794 (N_9794,N_7120,N_7666);
and U9795 (N_9795,N_7490,N_7023);
nand U9796 (N_9796,N_7383,N_7551);
nand U9797 (N_9797,N_6442,N_7703);
nand U9798 (N_9798,N_8995,N_8047);
and U9799 (N_9799,N_8804,N_6042);
xnor U9800 (N_9800,N_6118,N_8954);
and U9801 (N_9801,N_8871,N_7110);
nand U9802 (N_9802,N_7092,N_6528);
or U9803 (N_9803,N_7376,N_6921);
and U9804 (N_9804,N_6737,N_6077);
nor U9805 (N_9805,N_6087,N_6611);
nor U9806 (N_9806,N_8697,N_6312);
nor U9807 (N_9807,N_6588,N_7132);
nand U9808 (N_9808,N_6760,N_7526);
and U9809 (N_9809,N_6130,N_7632);
and U9810 (N_9810,N_6973,N_6012);
and U9811 (N_9811,N_6248,N_7879);
and U9812 (N_9812,N_7691,N_6153);
xnor U9813 (N_9813,N_8261,N_8119);
nor U9814 (N_9814,N_8980,N_8672);
xnor U9815 (N_9815,N_7346,N_6998);
nor U9816 (N_9816,N_8461,N_8798);
nand U9817 (N_9817,N_6345,N_6937);
or U9818 (N_9818,N_6513,N_6308);
nand U9819 (N_9819,N_7850,N_6141);
and U9820 (N_9820,N_7502,N_6792);
nand U9821 (N_9821,N_6373,N_7650);
or U9822 (N_9822,N_8906,N_7136);
and U9823 (N_9823,N_6954,N_7857);
xnor U9824 (N_9824,N_6180,N_6441);
and U9825 (N_9825,N_6894,N_8856);
and U9826 (N_9826,N_8101,N_6232);
and U9827 (N_9827,N_6943,N_8730);
nor U9828 (N_9828,N_6423,N_7639);
nand U9829 (N_9829,N_6206,N_8135);
and U9830 (N_9830,N_6713,N_7398);
nor U9831 (N_9831,N_7243,N_6375);
xnor U9832 (N_9832,N_6644,N_8000);
or U9833 (N_9833,N_6436,N_6191);
nand U9834 (N_9834,N_6485,N_8941);
or U9835 (N_9835,N_7240,N_7409);
or U9836 (N_9836,N_6092,N_6832);
nand U9837 (N_9837,N_6288,N_6405);
nand U9838 (N_9838,N_8136,N_6387);
or U9839 (N_9839,N_8341,N_7175);
xnor U9840 (N_9840,N_7882,N_7699);
and U9841 (N_9841,N_7404,N_7361);
and U9842 (N_9842,N_6081,N_8026);
or U9843 (N_9843,N_8643,N_6566);
or U9844 (N_9844,N_7949,N_6804);
xor U9845 (N_9845,N_6654,N_8799);
nand U9846 (N_9846,N_8206,N_6408);
nor U9847 (N_9847,N_7330,N_7140);
and U9848 (N_9848,N_8940,N_6844);
xor U9849 (N_9849,N_7947,N_6399);
and U9850 (N_9850,N_8803,N_7310);
nand U9851 (N_9851,N_7487,N_6674);
and U9852 (N_9852,N_8789,N_6235);
nand U9853 (N_9853,N_7113,N_6755);
nand U9854 (N_9854,N_8219,N_8458);
and U9855 (N_9855,N_8103,N_6411);
xor U9856 (N_9856,N_6525,N_7885);
and U9857 (N_9857,N_6672,N_7934);
and U9858 (N_9858,N_8408,N_7216);
nor U9859 (N_9859,N_7833,N_7615);
nor U9860 (N_9860,N_7315,N_7389);
nor U9861 (N_9861,N_7001,N_6445);
or U9862 (N_9862,N_8113,N_6051);
nand U9863 (N_9863,N_6490,N_7042);
nand U9864 (N_9864,N_6996,N_6884);
nor U9865 (N_9865,N_7774,N_6881);
nand U9866 (N_9866,N_7426,N_6959);
or U9867 (N_9867,N_7938,N_6133);
and U9868 (N_9868,N_6729,N_6563);
and U9869 (N_9869,N_8096,N_7805);
nor U9870 (N_9870,N_8009,N_7789);
nand U9871 (N_9871,N_8230,N_7283);
xnor U9872 (N_9872,N_8169,N_7808);
nor U9873 (N_9873,N_7756,N_6226);
and U9874 (N_9874,N_8805,N_6634);
xnor U9875 (N_9875,N_8560,N_8704);
or U9876 (N_9876,N_7765,N_8286);
or U9877 (N_9877,N_7950,N_6336);
nor U9878 (N_9878,N_7238,N_6018);
or U9879 (N_9879,N_6739,N_7545);
nand U9880 (N_9880,N_8366,N_6652);
nand U9881 (N_9881,N_7053,N_6590);
or U9882 (N_9882,N_6409,N_6687);
nand U9883 (N_9883,N_6637,N_7523);
nor U9884 (N_9884,N_8742,N_8098);
xor U9885 (N_9885,N_7746,N_6359);
nand U9886 (N_9886,N_7091,N_8404);
nand U9887 (N_9887,N_8556,N_8780);
nor U9888 (N_9888,N_7821,N_8776);
and U9889 (N_9889,N_8715,N_7606);
nor U9890 (N_9890,N_6318,N_6991);
or U9891 (N_9891,N_7988,N_8259);
or U9892 (N_9892,N_6020,N_8745);
nor U9893 (N_9893,N_8958,N_7635);
and U9894 (N_9894,N_8476,N_7039);
nor U9895 (N_9895,N_6435,N_7876);
or U9896 (N_9896,N_8181,N_6233);
or U9897 (N_9897,N_8564,N_6758);
nor U9898 (N_9898,N_7741,N_7367);
and U9899 (N_9899,N_7427,N_6971);
or U9900 (N_9900,N_8557,N_8426);
nor U9901 (N_9901,N_7050,N_6358);
and U9902 (N_9902,N_6048,N_7880);
nor U9903 (N_9903,N_8817,N_6125);
and U9904 (N_9904,N_6159,N_7593);
nand U9905 (N_9905,N_6829,N_6871);
nand U9906 (N_9906,N_6241,N_7160);
nor U9907 (N_9907,N_7690,N_8824);
or U9908 (N_9908,N_7567,N_6578);
or U9909 (N_9909,N_7272,N_6591);
nand U9910 (N_9910,N_7337,N_6404);
nand U9911 (N_9911,N_6794,N_7655);
and U9912 (N_9912,N_8629,N_6505);
and U9913 (N_9913,N_6764,N_6765);
or U9914 (N_9914,N_7124,N_8975);
nor U9915 (N_9915,N_6957,N_8750);
or U9916 (N_9916,N_8446,N_6533);
nand U9917 (N_9917,N_6044,N_6009);
nand U9918 (N_9918,N_7974,N_8773);
nand U9919 (N_9919,N_6364,N_8320);
and U9920 (N_9920,N_6860,N_8309);
or U9921 (N_9921,N_7524,N_7378);
or U9922 (N_9922,N_8874,N_7903);
nand U9923 (N_9923,N_7801,N_7109);
xor U9924 (N_9924,N_6582,N_6074);
nand U9925 (N_9925,N_7341,N_7583);
nor U9926 (N_9926,N_7466,N_8379);
and U9927 (N_9927,N_6963,N_8894);
and U9928 (N_9928,N_7441,N_7928);
xor U9929 (N_9929,N_6837,N_8291);
or U9930 (N_9930,N_8637,N_7463);
nand U9931 (N_9931,N_6212,N_8700);
nor U9932 (N_9932,N_7814,N_7980);
or U9933 (N_9933,N_6799,N_8018);
nand U9934 (N_9934,N_8854,N_7453);
nand U9935 (N_9935,N_7414,N_7971);
and U9936 (N_9936,N_6772,N_8144);
xor U9937 (N_9937,N_7048,N_8163);
nor U9938 (N_9938,N_7147,N_7018);
nand U9939 (N_9939,N_7984,N_8377);
nand U9940 (N_9940,N_7424,N_7260);
or U9941 (N_9941,N_8796,N_6007);
and U9942 (N_9942,N_7585,N_7642);
xor U9943 (N_9943,N_7203,N_8848);
or U9944 (N_9944,N_8477,N_8178);
or U9945 (N_9945,N_8565,N_6635);
nand U9946 (N_9946,N_6424,N_6471);
nor U9947 (N_9947,N_7942,N_6978);
and U9948 (N_9948,N_6204,N_6274);
nor U9949 (N_9949,N_6023,N_8655);
or U9950 (N_9950,N_6942,N_7582);
or U9951 (N_9951,N_6476,N_7603);
and U9952 (N_9952,N_8383,N_8899);
or U9953 (N_9953,N_7027,N_8864);
and U9954 (N_9954,N_8391,N_6622);
nor U9955 (N_9955,N_6834,N_7400);
nand U9956 (N_9956,N_8782,N_8288);
and U9957 (N_9957,N_6254,N_8946);
nor U9958 (N_9958,N_7712,N_7074);
nand U9959 (N_9959,N_6950,N_8236);
and U9960 (N_9960,N_7923,N_6029);
nand U9961 (N_9961,N_6481,N_8177);
nand U9962 (N_9962,N_8744,N_6309);
and U9963 (N_9963,N_8999,N_8396);
or U9964 (N_9964,N_8646,N_6237);
nor U9965 (N_9965,N_6478,N_8670);
nor U9966 (N_9966,N_6150,N_7838);
nor U9967 (N_9967,N_7008,N_7492);
or U9968 (N_9968,N_8841,N_8861);
and U9969 (N_9969,N_8290,N_8271);
nor U9970 (N_9970,N_8051,N_6612);
or U9971 (N_9971,N_7695,N_6006);
or U9972 (N_9972,N_7444,N_7684);
and U9973 (N_9973,N_8807,N_6543);
or U9974 (N_9974,N_7688,N_8007);
or U9975 (N_9975,N_6608,N_8360);
or U9976 (N_9976,N_6929,N_6677);
nor U9977 (N_9977,N_7118,N_7531);
and U9978 (N_9978,N_6678,N_7501);
nor U9979 (N_9979,N_6793,N_7594);
xor U9980 (N_9980,N_6017,N_8419);
xnor U9981 (N_9981,N_6666,N_8440);
nor U9982 (N_9982,N_7055,N_8398);
xor U9983 (N_9983,N_8936,N_7658);
nor U9984 (N_9984,N_8651,N_7815);
nand U9985 (N_9985,N_7770,N_8257);
or U9986 (N_9986,N_6864,N_8640);
or U9987 (N_9987,N_8751,N_7030);
nand U9988 (N_9988,N_8384,N_7227);
nand U9989 (N_9989,N_7212,N_6260);
and U9990 (N_9990,N_6796,N_8301);
xnor U9991 (N_9991,N_6817,N_8053);
nand U9992 (N_9992,N_6836,N_6516);
nand U9993 (N_9993,N_8375,N_7114);
nand U9994 (N_9994,N_7007,N_6189);
or U9995 (N_9995,N_7348,N_8346);
and U9996 (N_9996,N_7035,N_7386);
or U9997 (N_9997,N_7097,N_6498);
nor U9998 (N_9998,N_7225,N_8834);
nor U9999 (N_9999,N_7458,N_6272);
nor U10000 (N_10000,N_7435,N_6833);
nor U10001 (N_10001,N_8689,N_8148);
xnor U10002 (N_10002,N_7510,N_7588);
and U10003 (N_10003,N_8706,N_7161);
or U10004 (N_10004,N_8185,N_8902);
nor U10005 (N_10005,N_6550,N_7820);
or U10006 (N_10006,N_6275,N_6366);
and U10007 (N_10007,N_6985,N_7385);
nor U10008 (N_10008,N_6861,N_6084);
nor U10009 (N_10009,N_6085,N_8809);
and U10010 (N_10010,N_8228,N_6703);
nor U10011 (N_10011,N_6923,N_8097);
nand U10012 (N_10012,N_7713,N_6403);
or U10013 (N_10013,N_7029,N_8994);
or U10014 (N_10014,N_6596,N_8769);
or U10015 (N_10015,N_8654,N_8195);
or U10016 (N_10016,N_8749,N_8993);
nand U10017 (N_10017,N_7898,N_6052);
or U10018 (N_10018,N_8435,N_8507);
and U10019 (N_10019,N_7932,N_6446);
nand U10020 (N_10020,N_8757,N_7795);
nor U10021 (N_10021,N_6640,N_6470);
nand U10022 (N_10022,N_8488,N_7170);
and U10023 (N_10023,N_6740,N_8681);
nor U10024 (N_10024,N_7421,N_7060);
nand U10025 (N_10025,N_6072,N_6419);
nand U10026 (N_10026,N_8339,N_8220);
nor U10027 (N_10027,N_7595,N_6098);
nor U10028 (N_10028,N_6314,N_6004);
and U10029 (N_10029,N_7571,N_8499);
nand U10030 (N_10030,N_6489,N_7930);
and U10031 (N_10031,N_7456,N_8933);
and U10032 (N_10032,N_6437,N_6205);
nor U10033 (N_10033,N_7911,N_6443);
nand U10034 (N_10034,N_7671,N_7939);
nor U10035 (N_10035,N_7878,N_8387);
or U10036 (N_10036,N_7364,N_6492);
nor U10037 (N_10037,N_8450,N_6222);
and U10038 (N_10038,N_8891,N_7846);
nand U10039 (N_10039,N_8795,N_7078);
nand U10040 (N_10040,N_8351,N_8154);
and U10041 (N_10041,N_8464,N_6166);
nand U10042 (N_10042,N_8193,N_8692);
nand U10043 (N_10043,N_6822,N_8358);
and U10044 (N_10044,N_7533,N_7232);
nor U10045 (N_10045,N_8468,N_8182);
xor U10046 (N_10046,N_7479,N_6802);
and U10047 (N_10047,N_8687,N_6290);
or U10048 (N_10048,N_6593,N_7084);
nand U10049 (N_10049,N_6886,N_8598);
or U10050 (N_10050,N_8544,N_8693);
xor U10051 (N_10051,N_6236,N_7570);
xor U10052 (N_10052,N_7245,N_7462);
and U10053 (N_10053,N_7368,N_8979);
nor U10054 (N_10054,N_8239,N_7745);
or U10055 (N_10055,N_6101,N_7813);
nand U10056 (N_10056,N_7633,N_7256);
nor U10057 (N_10057,N_7072,N_7445);
nand U10058 (N_10058,N_8659,N_6523);
nor U10059 (N_10059,N_7339,N_8138);
or U10060 (N_10060,N_6428,N_6826);
nor U10061 (N_10061,N_6295,N_8900);
nand U10062 (N_10062,N_7164,N_7719);
nor U10063 (N_10063,N_7781,N_7870);
and U10064 (N_10064,N_6665,N_8578);
or U10065 (N_10065,N_8143,N_8418);
or U10066 (N_10066,N_8589,N_8362);
nor U10067 (N_10067,N_7131,N_8594);
nor U10068 (N_10068,N_6883,N_8091);
or U10069 (N_10069,N_8955,N_7344);
nand U10070 (N_10070,N_7177,N_8723);
nand U10071 (N_10071,N_8151,N_6920);
nand U10072 (N_10072,N_8923,N_7897);
nand U10073 (N_10073,N_7317,N_6827);
or U10074 (N_10074,N_8520,N_6811);
or U10075 (N_10075,N_8737,N_7117);
nor U10076 (N_10076,N_7889,N_6906);
and U10077 (N_10077,N_7313,N_7206);
nand U10078 (N_10078,N_7065,N_8073);
or U10079 (N_10079,N_8482,N_6631);
or U10080 (N_10080,N_8409,N_7906);
nand U10081 (N_10081,N_6539,N_7275);
and U10082 (N_10082,N_7936,N_7156);
and U10083 (N_10083,N_6603,N_6828);
and U10084 (N_10084,N_7281,N_6271);
or U10085 (N_10085,N_6195,N_8439);
nand U10086 (N_10086,N_7231,N_6267);
nand U10087 (N_10087,N_6350,N_7009);
nor U10088 (N_10088,N_6031,N_6083);
nor U10089 (N_10089,N_8882,N_6744);
or U10090 (N_10090,N_6918,N_7511);
or U10091 (N_10091,N_8289,N_8961);
and U10092 (N_10092,N_8898,N_7182);
or U10093 (N_10093,N_8952,N_7554);
and U10094 (N_10094,N_7249,N_8963);
nand U10095 (N_10095,N_7622,N_7832);
nor U10096 (N_10096,N_7605,N_6174);
nand U10097 (N_10097,N_6142,N_8866);
and U10098 (N_10098,N_6806,N_8198);
or U10099 (N_10099,N_8006,N_8679);
and U10100 (N_10100,N_7940,N_7686);
or U10101 (N_10101,N_6194,N_8317);
nor U10102 (N_10102,N_6580,N_7763);
and U10103 (N_10103,N_6876,N_6554);
nor U10104 (N_10104,N_8431,N_8585);
or U10105 (N_10105,N_8555,N_8641);
nand U10106 (N_10106,N_8673,N_7577);
nor U10107 (N_10107,N_8459,N_6269);
nand U10108 (N_10108,N_8905,N_8368);
nand U10109 (N_10109,N_7391,N_8012);
nand U10110 (N_10110,N_6605,N_8566);
and U10111 (N_10111,N_8724,N_8237);
or U10112 (N_10112,N_7747,N_8610);
nor U10113 (N_10113,N_6019,N_6315);
xnor U10114 (N_10114,N_7464,N_6546);
xnor U10115 (N_10115,N_8986,N_6931);
nand U10116 (N_10116,N_7915,N_8608);
or U10117 (N_10117,N_7079,N_6305);
nand U10118 (N_10118,N_8838,N_8624);
or U10119 (N_10119,N_6053,N_8840);
nor U10120 (N_10120,N_7717,N_7859);
nand U10121 (N_10121,N_7624,N_7626);
nand U10122 (N_10122,N_7607,N_7473);
nand U10123 (N_10123,N_7888,N_8337);
nand U10124 (N_10124,N_8910,N_6620);
nor U10125 (N_10125,N_6506,N_8134);
or U10126 (N_10126,N_6175,N_6757);
or U10127 (N_10127,N_7937,N_7956);
and U10128 (N_10128,N_8971,N_8666);
nor U10129 (N_10129,N_7234,N_6307);
nand U10130 (N_10130,N_7417,N_8251);
nand U10131 (N_10131,N_8943,N_7085);
xor U10132 (N_10132,N_7173,N_6187);
and U10133 (N_10133,N_7899,N_6697);
xor U10134 (N_10134,N_8621,N_8731);
nand U10135 (N_10135,N_7702,N_6555);
nand U10136 (N_10136,N_8406,N_6132);
or U10137 (N_10137,N_7280,N_6711);
nand U10138 (N_10138,N_6745,N_8028);
or U10139 (N_10139,N_6467,N_8044);
and U10140 (N_10140,N_8932,N_7239);
or U10141 (N_10141,N_8394,N_6480);
and U10142 (N_10142,N_6902,N_8059);
or U10143 (N_10143,N_6693,N_6263);
nand U10144 (N_10144,N_8083,N_8926);
and U10145 (N_10145,N_8922,N_8300);
or U10146 (N_10146,N_6208,N_7679);
and U10147 (N_10147,N_6093,N_8345);
nand U10148 (N_10148,N_8112,N_7043);
xnor U10149 (N_10149,N_6257,N_8676);
and U10150 (N_10150,N_7470,N_7564);
nor U10151 (N_10151,N_7306,N_6680);
nand U10152 (N_10152,N_7953,N_7542);
nor U10153 (N_10153,N_6502,N_6933);
or U10154 (N_10154,N_7735,N_6335);
or U10155 (N_10155,N_8616,N_7505);
nor U10156 (N_10156,N_7093,N_6261);
and U10157 (N_10157,N_7921,N_8027);
and U10158 (N_10158,N_7264,N_7299);
and U10159 (N_10159,N_7793,N_8355);
nand U10160 (N_10160,N_7056,N_7357);
nand U10161 (N_10161,N_7230,N_8472);
nor U10162 (N_10162,N_6039,N_7802);
or U10163 (N_10163,N_6577,N_8859);
nand U10164 (N_10164,N_8797,N_7610);
and U10165 (N_10165,N_6699,N_7329);
or U10166 (N_10166,N_7665,N_6790);
or U10167 (N_10167,N_6982,N_8338);
and U10168 (N_10168,N_6741,N_6378);
and U10169 (N_10169,N_6812,N_8927);
or U10170 (N_10170,N_8869,N_6769);
and U10171 (N_10171,N_8107,N_8683);
nand U10172 (N_10172,N_6022,N_7925);
and U10173 (N_10173,N_7413,N_7069);
or U10174 (N_10174,N_7836,N_6147);
nand U10175 (N_10175,N_7927,N_7331);
and U10176 (N_10176,N_7896,N_8099);
nor U10177 (N_10177,N_6686,N_7561);
xor U10178 (N_10178,N_8323,N_6961);
and U10179 (N_10179,N_7015,N_8021);
xor U10180 (N_10180,N_7323,N_6041);
or U10181 (N_10181,N_6054,N_8064);
nand U10182 (N_10182,N_6148,N_7760);
and U10183 (N_10183,N_6692,N_7044);
or U10184 (N_10184,N_6361,N_7748);
nor U10185 (N_10185,N_8120,N_7460);
nor U10186 (N_10186,N_6664,N_7724);
or U10187 (N_10187,N_7960,N_7373);
or U10188 (N_10188,N_7254,N_6114);
nor U10189 (N_10189,N_7276,N_6050);
xnor U10190 (N_10190,N_8127,N_8966);
or U10191 (N_10191,N_7152,N_7215);
nor U10192 (N_10192,N_7422,N_7827);
nor U10193 (N_10193,N_7285,N_7262);
nor U10194 (N_10194,N_7073,N_8956);
or U10195 (N_10195,N_8152,N_8045);
and U10196 (N_10196,N_7477,N_8326);
or U10197 (N_10197,N_6508,N_7967);
or U10198 (N_10198,N_8509,N_8663);
or U10199 (N_10199,N_8388,N_6877);
nor U10200 (N_10200,N_8879,N_8299);
nor U10201 (N_10201,N_6370,N_7061);
or U10202 (N_10202,N_8925,N_7865);
nand U10203 (N_10203,N_7534,N_7982);
and U10204 (N_10204,N_8100,N_8713);
and U10205 (N_10205,N_6681,N_6422);
nor U10206 (N_10206,N_6154,N_8075);
and U10207 (N_10207,N_6273,N_8460);
or U10208 (N_10208,N_7736,N_7318);
or U10209 (N_10209,N_8645,N_7210);
nand U10210 (N_10210,N_8129,N_8591);
xor U10211 (N_10211,N_6465,N_8179);
xnor U10212 (N_10212,N_7959,N_8908);
nor U10213 (N_10213,N_6809,N_8787);
and U10214 (N_10214,N_7648,N_6763);
or U10215 (N_10215,N_6880,N_8123);
or U10216 (N_10216,N_6381,N_8774);
and U10217 (N_10217,N_7824,N_7957);
and U10218 (N_10218,N_7491,N_6722);
nor U10219 (N_10219,N_6893,N_7098);
nor U10220 (N_10220,N_7474,N_8741);
nand U10221 (N_10221,N_8001,N_6801);
xor U10222 (N_10222,N_7016,N_6281);
nand U10223 (N_10223,N_6161,N_7755);
xor U10224 (N_10224,N_6586,N_8324);
nand U10225 (N_10225,N_6459,N_8784);
or U10226 (N_10226,N_6818,N_8032);
nand U10227 (N_10227,N_7241,N_7970);
and U10228 (N_10228,N_7538,N_6224);
or U10229 (N_10229,N_6552,N_8533);
nand U10230 (N_10230,N_8200,N_8747);
and U10231 (N_10231,N_7500,N_7321);
and U10232 (N_10232,N_8668,N_8089);
nand U10233 (N_10233,N_7433,N_8800);
nor U10234 (N_10234,N_8093,N_7856);
xnor U10235 (N_10235,N_7416,N_8270);
or U10236 (N_10236,N_7547,N_7158);
xor U10237 (N_10237,N_6888,N_7228);
nor U10238 (N_10238,N_6668,N_6369);
and U10239 (N_10239,N_6922,N_6633);
nor U10240 (N_10240,N_7316,N_7917);
or U10241 (N_10241,N_8945,N_8014);
or U10242 (N_10242,N_8137,N_8552);
or U10243 (N_10243,N_6540,N_7924);
and U10244 (N_10244,N_6383,N_6068);
and U10245 (N_10245,N_7049,N_6016);
xor U10246 (N_10246,N_7450,N_7987);
and U10247 (N_10247,N_7218,N_7592);
nand U10248 (N_10248,N_7660,N_8907);
and U10249 (N_10249,N_6173,N_7268);
or U10250 (N_10250,N_7469,N_7382);
nor U10251 (N_10251,N_6401,N_6651);
nor U10252 (N_10252,N_6878,N_8984);
nand U10253 (N_10253,N_6377,N_8695);
and U10254 (N_10254,N_6137,N_7149);
nand U10255 (N_10255,N_6567,N_7282);
and U10256 (N_10256,N_8878,N_7528);
nand U10257 (N_10257,N_8549,N_8088);
xnor U10258 (N_10258,N_7751,N_8667);
and U10259 (N_10259,N_8865,N_8314);
or U10260 (N_10260,N_7353,N_6530);
nand U10261 (N_10261,N_8996,N_6200);
and U10262 (N_10262,N_7314,N_8416);
nor U10263 (N_10263,N_6059,N_7871);
or U10264 (N_10264,N_8397,N_8298);
and U10265 (N_10265,N_6171,N_6472);
xor U10266 (N_10266,N_7347,N_7407);
nor U10267 (N_10267,N_8970,N_6117);
nand U10268 (N_10268,N_8192,N_7362);
or U10269 (N_10269,N_7716,N_8037);
or U10270 (N_10270,N_7115,N_7408);
and U10271 (N_10271,N_6708,N_6976);
and U10272 (N_10272,N_8983,N_8962);
nor U10273 (N_10273,N_8850,N_8981);
or U10274 (N_10274,N_6736,N_7521);
nor U10275 (N_10275,N_7209,N_7066);
xor U10276 (N_10276,N_6863,N_8490);
and U10277 (N_10277,N_6203,N_8470);
nor U10278 (N_10278,N_6621,N_7777);
or U10279 (N_10279,N_7514,N_6123);
and U10280 (N_10280,N_7985,N_7565);
or U10281 (N_10281,N_8057,N_8485);
and U10282 (N_10282,N_7207,N_7423);
and U10283 (N_10283,N_7192,N_7289);
or U10284 (N_10284,N_7220,N_7811);
nand U10285 (N_10285,N_7133,N_8978);
or U10286 (N_10286,N_6116,N_8595);
nand U10287 (N_10287,N_6097,N_6823);
xor U10288 (N_10288,N_8312,N_7478);
or U10289 (N_10289,N_6326,N_6775);
and U10290 (N_10290,N_8579,N_7780);
nand U10291 (N_10291,N_8034,N_8830);
nand U10292 (N_10292,N_6535,N_8316);
and U10293 (N_10293,N_6330,N_8583);
nor U10294 (N_10294,N_7644,N_6630);
nand U10295 (N_10295,N_6218,N_8563);
and U10296 (N_10296,N_6397,N_7893);
nor U10297 (N_10297,N_8677,N_7190);
nor U10298 (N_10298,N_6999,N_8427);
and U10299 (N_10299,N_8216,N_7549);
nor U10300 (N_10300,N_6024,N_8348);
nor U10301 (N_10301,N_8752,N_8886);
nor U10302 (N_10302,N_6199,N_8125);
nor U10303 (N_10303,N_8303,N_8658);
xnor U10304 (N_10304,N_7186,N_6694);
nand U10305 (N_10305,N_6228,N_7829);
xor U10306 (N_10306,N_8828,N_6919);
or U10307 (N_10307,N_8250,N_6372);
nor U10308 (N_10308,N_7075,N_7697);
or U10309 (N_10309,N_7403,N_8660);
and U10310 (N_10310,N_8921,N_7863);
nand U10311 (N_10311,N_7729,N_7954);
and U10312 (N_10312,N_6426,N_8561);
or U10313 (N_10313,N_6610,N_8060);
nor U10314 (N_10314,N_7916,N_7363);
nand U10315 (N_10315,N_7459,N_7816);
nand U10316 (N_10316,N_6371,N_6606);
nor U10317 (N_10317,N_7946,N_7905);
xnor U10318 (N_10318,N_6002,N_8285);
or U10319 (N_10319,N_8639,N_7045);
nor U10320 (N_10320,N_8036,N_8821);
nor U10321 (N_10321,N_7687,N_6759);
nor U10322 (N_10322,N_7384,N_7706);
nand U10323 (N_10323,N_8951,N_6038);
nand U10324 (N_10324,N_6496,N_8041);
nor U10325 (N_10325,N_6304,N_6820);
nand U10326 (N_10326,N_6663,N_6058);
xor U10327 (N_10327,N_7196,N_7111);
or U10328 (N_10328,N_7270,N_7894);
and U10329 (N_10329,N_8901,N_6896);
and U10330 (N_10330,N_6568,N_7224);
nand U10331 (N_10331,N_8577,N_7080);
nand U10332 (N_10332,N_8480,N_7265);
or U10333 (N_10333,N_7096,N_7419);
nor U10334 (N_10334,N_8917,N_7933);
or U10335 (N_10335,N_8601,N_7211);
or U10336 (N_10336,N_6842,N_6791);
nor U10337 (N_10337,N_8586,N_8895);
nand U10338 (N_10338,N_6724,N_7941);
nand U10339 (N_10339,N_6297,N_7328);
nor U10340 (N_10340,N_6571,N_8087);
nor U10341 (N_10341,N_6701,N_8600);
nor U10342 (N_10342,N_6151,N_6743);
nor U10343 (N_10343,N_6750,N_6140);
nand U10344 (N_10344,N_8353,N_6682);
xnor U10345 (N_10345,N_7102,N_7064);
xnor U10346 (N_10346,N_7332,N_7977);
nand U10347 (N_10347,N_6771,N_8875);
and U10348 (N_10348,N_8535,N_8959);
or U10349 (N_10349,N_8248,N_8942);
and U10350 (N_10350,N_8124,N_8278);
nand U10351 (N_10351,N_7322,N_6095);
nand U10352 (N_10352,N_6135,N_6010);
and U10353 (N_10353,N_6134,N_6866);
nor U10354 (N_10354,N_8109,N_7340);
or U10355 (N_10355,N_6934,N_8445);
nand U10356 (N_10356,N_7257,N_6223);
xnor U10357 (N_10357,N_7351,N_7358);
xnor U10358 (N_10358,N_8893,N_6924);
nand U10359 (N_10359,N_8172,N_6139);
or U10360 (N_10360,N_6210,N_7484);
nor U10361 (N_10361,N_7599,N_7951);
xnor U10362 (N_10362,N_6321,N_8913);
nor U10363 (N_10363,N_7038,N_6021);
or U10364 (N_10364,N_8532,N_6112);
and U10365 (N_10365,N_7579,N_8990);
or U10366 (N_10366,N_6627,N_8928);
nand U10367 (N_10367,N_6726,N_6564);
or U10368 (N_10368,N_8748,N_8010);
and U10369 (N_10369,N_8548,N_6935);
or U10370 (N_10370,N_7990,N_7530);
and U10371 (N_10371,N_8620,N_8845);
and U10372 (N_10372,N_6179,N_6313);
nor U10373 (N_10373,N_8992,N_6908);
nand U10374 (N_10374,N_8393,N_8631);
nor U10375 (N_10375,N_8025,N_7778);
nand U10376 (N_10376,N_7248,N_8380);
nand U10377 (N_10377,N_6852,N_8174);
or U10378 (N_10378,N_8870,N_6349);
and U10379 (N_10379,N_7766,N_7809);
or U10380 (N_10380,N_8247,N_6046);
nor U10381 (N_10381,N_8860,N_8766);
nand U10382 (N_10382,N_8260,N_8858);
nand U10383 (N_10383,N_8424,N_6064);
and U10384 (N_10384,N_7731,N_8201);
and U10385 (N_10385,N_7590,N_6328);
nor U10386 (N_10386,N_6688,N_6900);
nor U10387 (N_10387,N_7370,N_7734);
and U10388 (N_10388,N_7981,N_7512);
or U10389 (N_10389,N_8606,N_6614);
and U10390 (N_10390,N_8717,N_8918);
or U10391 (N_10391,N_8238,N_6276);
nor U10392 (N_10392,N_6735,N_8855);
and U10393 (N_10393,N_8714,N_7325);
or U10394 (N_10394,N_8511,N_8889);
and U10395 (N_10395,N_8273,N_6990);
nand U10396 (N_10396,N_7183,N_7886);
nand U10397 (N_10397,N_7086,N_7432);
or U10398 (N_10398,N_8812,N_8327);
xnor U10399 (N_10399,N_6299,N_6469);
xnor U10400 (N_10400,N_8302,N_6968);
xor U10401 (N_10401,N_7807,N_7101);
or U10402 (N_10402,N_7535,N_8131);
nand U10403 (N_10403,N_8493,N_7174);
nor U10404 (N_10404,N_6847,N_6121);
and U10405 (N_10405,N_7082,N_6106);
nand U10406 (N_10406,N_7128,N_8546);
or U10407 (N_10407,N_8401,N_6751);
and U10408 (N_10408,N_6899,N_6293);
nand U10409 (N_10409,N_6119,N_8729);
and U10410 (N_10410,N_8813,N_8443);
nand U10411 (N_10411,N_8452,N_6049);
nor U10412 (N_10412,N_8630,N_7952);
xnor U10413 (N_10413,N_7630,N_7356);
and U10414 (N_10414,N_8820,N_8691);
and U10415 (N_10415,N_7768,N_8890);
nor U10416 (N_10416,N_7553,N_7783);
xor U10417 (N_10417,N_8282,N_6475);
nand U10418 (N_10418,N_7628,N_8614);
xor U10419 (N_10419,N_8373,N_7707);
nand U10420 (N_10420,N_6865,N_8968);
nand U10421 (N_10421,N_6655,N_6196);
or U10422 (N_10422,N_8885,N_8785);
and U10423 (N_10423,N_8039,N_7103);
nor U10424 (N_10424,N_6431,N_6030);
nor U10425 (N_10425,N_8349,N_8043);
nor U10426 (N_10426,N_6468,N_8974);
xor U10427 (N_10427,N_7295,N_6213);
and U10428 (N_10428,N_6091,N_6334);
nand U10429 (N_10429,N_7852,N_7996);
or U10430 (N_10430,N_7782,N_8086);
xor U10431 (N_10431,N_7471,N_8808);
xnor U10432 (N_10432,N_8330,N_6816);
and U10433 (N_10433,N_7552,N_7396);
and U10434 (N_10434,N_6165,N_8935);
nor U10435 (N_10435,N_6838,N_6071);
and U10436 (N_10436,N_8432,N_6925);
xnor U10437 (N_10437,N_6238,N_8743);
and U10438 (N_10438,N_6892,N_6462);
nand U10439 (N_10439,N_7150,N_7187);
xor U10440 (N_10440,N_7900,N_6512);
nand U10441 (N_10441,N_8165,N_6283);
and U10442 (N_10442,N_7620,N_7191);
nand U10443 (N_10443,N_6901,N_7440);
or U10444 (N_10444,N_6494,N_6519);
or U10445 (N_10445,N_8949,N_6625);
nor U10446 (N_10446,N_6264,N_6357);
nor U10447 (N_10447,N_6784,N_6748);
nor U10448 (N_10448,N_7675,N_6252);
or U10449 (N_10449,N_8973,N_6636);
or U10450 (N_10450,N_7017,N_8581);
or U10451 (N_10451,N_8991,N_7645);
or U10452 (N_10452,N_6720,N_6491);
and U10453 (N_10453,N_8110,N_8217);
nand U10454 (N_10454,N_8376,N_6579);
nand U10455 (N_10455,N_8315,N_8836);
nand U10456 (N_10456,N_7189,N_8155);
or U10457 (N_10457,N_7506,N_7388);
and U10458 (N_10458,N_8372,N_8013);
nand U10459 (N_10459,N_6479,N_6447);
or U10460 (N_10460,N_7559,N_8783);
nor U10461 (N_10461,N_6386,N_8924);
nand U10462 (N_10462,N_6207,N_8590);
or U10463 (N_10463,N_7683,N_6425);
or U10464 (N_10464,N_7468,N_7032);
nor U10465 (N_10465,N_7669,N_8530);
nor U10466 (N_10466,N_7842,N_7823);
nor U10467 (N_10467,N_7179,N_8599);
xor U10468 (N_10468,N_7790,N_8823);
or U10469 (N_10469,N_7962,N_7062);
nand U10470 (N_10470,N_7217,N_7415);
nand U10471 (N_10471,N_7520,N_8020);
nand U10472 (N_10472,N_6079,N_6149);
or U10473 (N_10473,N_7246,N_7926);
nor U10474 (N_10474,N_8240,N_8077);
nor U10475 (N_10475,N_7696,N_6859);
nor U10476 (N_10476,N_8333,N_7184);
xor U10477 (N_10477,N_6311,N_6872);
and U10478 (N_10478,N_7560,N_6867);
xnor U10479 (N_10479,N_6356,N_8357);
nand U10480 (N_10480,N_7381,N_8215);
xor U10481 (N_10481,N_6733,N_8475);
and U10482 (N_10482,N_8525,N_6746);
xnor U10483 (N_10483,N_8328,N_7291);
xnor U10484 (N_10484,N_6291,N_7360);
nor U10485 (N_10485,N_6618,N_8069);
or U10486 (N_10486,N_8508,N_7185);
xor U10487 (N_10487,N_7999,N_6949);
xnor U10488 (N_10488,N_7195,N_8665);
or U10489 (N_10489,N_8126,N_8030);
and U10490 (N_10490,N_6789,N_6595);
and U10491 (N_10491,N_8832,N_8604);
nor U10492 (N_10492,N_8356,N_7394);
nor U10493 (N_10493,N_7162,N_6453);
and U10494 (N_10494,N_8934,N_7165);
nand U10495 (N_10495,N_8063,N_6669);
and U10496 (N_10496,N_6219,N_6705);
or U10497 (N_10497,N_6340,N_8190);
and U10498 (N_10498,N_7251,N_6440);
or U10499 (N_10499,N_8411,N_7698);
nor U10500 (N_10500,N_6760,N_8841);
nor U10501 (N_10501,N_6149,N_8044);
nand U10502 (N_10502,N_6766,N_7117);
nor U10503 (N_10503,N_8616,N_7088);
nor U10504 (N_10504,N_8236,N_6023);
and U10505 (N_10505,N_8881,N_7255);
nor U10506 (N_10506,N_8040,N_7234);
nand U10507 (N_10507,N_6207,N_7760);
nor U10508 (N_10508,N_6622,N_8706);
xor U10509 (N_10509,N_8789,N_8520);
nor U10510 (N_10510,N_6926,N_6957);
and U10511 (N_10511,N_8568,N_8127);
and U10512 (N_10512,N_6102,N_6059);
or U10513 (N_10513,N_7045,N_6145);
nand U10514 (N_10514,N_7598,N_6360);
nand U10515 (N_10515,N_8907,N_8656);
or U10516 (N_10516,N_6769,N_7304);
nand U10517 (N_10517,N_6865,N_6582);
and U10518 (N_10518,N_8773,N_8939);
or U10519 (N_10519,N_8285,N_7115);
and U10520 (N_10520,N_7624,N_8869);
nor U10521 (N_10521,N_6252,N_6199);
nor U10522 (N_10522,N_6655,N_7654);
and U10523 (N_10523,N_8082,N_8910);
or U10524 (N_10524,N_7648,N_8209);
or U10525 (N_10525,N_7485,N_6306);
nor U10526 (N_10526,N_6562,N_8067);
and U10527 (N_10527,N_7248,N_8189);
or U10528 (N_10528,N_8963,N_8621);
nor U10529 (N_10529,N_8779,N_8180);
and U10530 (N_10530,N_6602,N_6502);
nor U10531 (N_10531,N_6263,N_6258);
nor U10532 (N_10532,N_8775,N_8150);
or U10533 (N_10533,N_7100,N_8289);
nand U10534 (N_10534,N_8586,N_7858);
nor U10535 (N_10535,N_8172,N_6389);
or U10536 (N_10536,N_7801,N_8452);
and U10537 (N_10537,N_6760,N_8390);
nor U10538 (N_10538,N_6916,N_7860);
or U10539 (N_10539,N_8594,N_7309);
or U10540 (N_10540,N_8508,N_6755);
nand U10541 (N_10541,N_8830,N_7185);
or U10542 (N_10542,N_8947,N_8329);
and U10543 (N_10543,N_7254,N_8264);
xor U10544 (N_10544,N_7785,N_8731);
and U10545 (N_10545,N_7404,N_6927);
nand U10546 (N_10546,N_8307,N_6211);
and U10547 (N_10547,N_8600,N_6865);
and U10548 (N_10548,N_6877,N_7131);
and U10549 (N_10549,N_8226,N_7798);
nor U10550 (N_10550,N_6170,N_8510);
and U10551 (N_10551,N_8044,N_7292);
and U10552 (N_10552,N_8964,N_8415);
and U10553 (N_10553,N_6585,N_6427);
or U10554 (N_10554,N_8454,N_6797);
and U10555 (N_10555,N_8571,N_7587);
and U10556 (N_10556,N_7738,N_7811);
nand U10557 (N_10557,N_7295,N_8457);
nor U10558 (N_10558,N_7080,N_6678);
xor U10559 (N_10559,N_7542,N_6210);
and U10560 (N_10560,N_6152,N_6619);
and U10561 (N_10561,N_8093,N_7678);
nor U10562 (N_10562,N_7116,N_7732);
or U10563 (N_10563,N_8760,N_8790);
xnor U10564 (N_10564,N_7008,N_8307);
nand U10565 (N_10565,N_7457,N_7190);
nor U10566 (N_10566,N_8504,N_7517);
and U10567 (N_10567,N_6719,N_8522);
or U10568 (N_10568,N_7889,N_6622);
or U10569 (N_10569,N_6846,N_8345);
nor U10570 (N_10570,N_7837,N_8430);
or U10571 (N_10571,N_7182,N_8295);
nor U10572 (N_10572,N_7020,N_6662);
nor U10573 (N_10573,N_6156,N_7707);
nand U10574 (N_10574,N_8424,N_8457);
nand U10575 (N_10575,N_8754,N_8006);
and U10576 (N_10576,N_8471,N_7256);
nand U10577 (N_10577,N_7637,N_7924);
and U10578 (N_10578,N_7259,N_6480);
xor U10579 (N_10579,N_7799,N_8183);
nand U10580 (N_10580,N_6250,N_7639);
nand U10581 (N_10581,N_8078,N_7948);
nor U10582 (N_10582,N_8039,N_7092);
and U10583 (N_10583,N_7288,N_7717);
nand U10584 (N_10584,N_8156,N_7873);
nand U10585 (N_10585,N_7562,N_8675);
nor U10586 (N_10586,N_6825,N_6661);
xor U10587 (N_10587,N_8735,N_8800);
and U10588 (N_10588,N_6378,N_6059);
nand U10589 (N_10589,N_8405,N_7403);
and U10590 (N_10590,N_8190,N_8199);
nor U10591 (N_10591,N_6250,N_7418);
and U10592 (N_10592,N_6664,N_8921);
xor U10593 (N_10593,N_7918,N_7557);
xnor U10594 (N_10594,N_6840,N_8632);
or U10595 (N_10595,N_7590,N_6174);
or U10596 (N_10596,N_8375,N_7998);
or U10597 (N_10597,N_6021,N_7839);
or U10598 (N_10598,N_8643,N_8324);
xor U10599 (N_10599,N_7828,N_6188);
and U10600 (N_10600,N_8069,N_7242);
or U10601 (N_10601,N_6710,N_7284);
nor U10602 (N_10602,N_6611,N_8845);
and U10603 (N_10603,N_7246,N_6230);
nand U10604 (N_10604,N_7508,N_6353);
nand U10605 (N_10605,N_8666,N_8301);
and U10606 (N_10606,N_6026,N_8517);
and U10607 (N_10607,N_7735,N_7432);
nand U10608 (N_10608,N_6841,N_7441);
or U10609 (N_10609,N_7443,N_7768);
and U10610 (N_10610,N_6024,N_8529);
and U10611 (N_10611,N_8636,N_8114);
nor U10612 (N_10612,N_8241,N_7409);
and U10613 (N_10613,N_6380,N_8493);
and U10614 (N_10614,N_7938,N_8230);
nor U10615 (N_10615,N_7487,N_7539);
or U10616 (N_10616,N_6990,N_6577);
nand U10617 (N_10617,N_8280,N_6761);
and U10618 (N_10618,N_7236,N_8274);
or U10619 (N_10619,N_6505,N_8428);
nand U10620 (N_10620,N_8925,N_6126);
or U10621 (N_10621,N_7001,N_7250);
or U10622 (N_10622,N_6426,N_8850);
or U10623 (N_10623,N_8911,N_6463);
nor U10624 (N_10624,N_8964,N_8180);
nor U10625 (N_10625,N_8554,N_6492);
nand U10626 (N_10626,N_6113,N_8651);
nor U10627 (N_10627,N_7673,N_8262);
xnor U10628 (N_10628,N_7464,N_7731);
nor U10629 (N_10629,N_6541,N_8780);
and U10630 (N_10630,N_6395,N_7975);
nand U10631 (N_10631,N_6215,N_8491);
and U10632 (N_10632,N_8611,N_7558);
nor U10633 (N_10633,N_7543,N_7021);
or U10634 (N_10634,N_8855,N_7125);
nand U10635 (N_10635,N_8699,N_8728);
nand U10636 (N_10636,N_8473,N_6911);
or U10637 (N_10637,N_8855,N_7613);
nand U10638 (N_10638,N_6861,N_8122);
nor U10639 (N_10639,N_8738,N_8565);
nand U10640 (N_10640,N_6165,N_6048);
nor U10641 (N_10641,N_6860,N_8696);
nor U10642 (N_10642,N_6091,N_7114);
or U10643 (N_10643,N_7780,N_6432);
xor U10644 (N_10644,N_8820,N_8951);
and U10645 (N_10645,N_7505,N_8088);
or U10646 (N_10646,N_6043,N_8028);
xor U10647 (N_10647,N_6666,N_8172);
or U10648 (N_10648,N_8357,N_7232);
nand U10649 (N_10649,N_6395,N_7414);
xor U10650 (N_10650,N_6341,N_8570);
nand U10651 (N_10651,N_6164,N_8662);
and U10652 (N_10652,N_6097,N_7393);
nor U10653 (N_10653,N_6750,N_6475);
and U10654 (N_10654,N_6157,N_8441);
and U10655 (N_10655,N_7155,N_8152);
or U10656 (N_10656,N_8718,N_8846);
nor U10657 (N_10657,N_6356,N_6851);
or U10658 (N_10658,N_6492,N_6652);
and U10659 (N_10659,N_8800,N_6517);
or U10660 (N_10660,N_6162,N_6786);
xor U10661 (N_10661,N_7710,N_8276);
nor U10662 (N_10662,N_8601,N_7800);
nand U10663 (N_10663,N_7558,N_7841);
and U10664 (N_10664,N_6140,N_7541);
nor U10665 (N_10665,N_6395,N_7025);
nand U10666 (N_10666,N_7617,N_7852);
and U10667 (N_10667,N_7389,N_6461);
xor U10668 (N_10668,N_8742,N_7373);
nor U10669 (N_10669,N_6282,N_7012);
nand U10670 (N_10670,N_6576,N_6850);
and U10671 (N_10671,N_8181,N_8797);
or U10672 (N_10672,N_7130,N_6181);
nand U10673 (N_10673,N_6080,N_6688);
xor U10674 (N_10674,N_8401,N_6669);
nor U10675 (N_10675,N_7865,N_6047);
nor U10676 (N_10676,N_6698,N_8632);
or U10677 (N_10677,N_7867,N_7669);
and U10678 (N_10678,N_8373,N_6251);
nor U10679 (N_10679,N_7495,N_7779);
or U10680 (N_10680,N_7810,N_7534);
nand U10681 (N_10681,N_6722,N_8671);
or U10682 (N_10682,N_8867,N_7808);
nor U10683 (N_10683,N_7384,N_8274);
nor U10684 (N_10684,N_6346,N_6604);
and U10685 (N_10685,N_6028,N_8479);
nor U10686 (N_10686,N_7381,N_7280);
nor U10687 (N_10687,N_8256,N_8366);
nor U10688 (N_10688,N_6588,N_7996);
or U10689 (N_10689,N_6693,N_8506);
nand U10690 (N_10690,N_8865,N_7042);
nand U10691 (N_10691,N_7828,N_7287);
nor U10692 (N_10692,N_8895,N_6072);
xor U10693 (N_10693,N_7058,N_6977);
or U10694 (N_10694,N_7619,N_7275);
or U10695 (N_10695,N_8284,N_6259);
and U10696 (N_10696,N_6188,N_6902);
xnor U10697 (N_10697,N_7021,N_8826);
nor U10698 (N_10698,N_6691,N_6866);
xnor U10699 (N_10699,N_7467,N_8030);
nand U10700 (N_10700,N_8970,N_6052);
nor U10701 (N_10701,N_6118,N_7624);
nand U10702 (N_10702,N_6088,N_6477);
or U10703 (N_10703,N_8160,N_8352);
nand U10704 (N_10704,N_6686,N_7268);
or U10705 (N_10705,N_8069,N_8446);
or U10706 (N_10706,N_7115,N_6926);
nor U10707 (N_10707,N_8423,N_7676);
and U10708 (N_10708,N_8339,N_7403);
and U10709 (N_10709,N_8192,N_7003);
nand U10710 (N_10710,N_7111,N_6381);
nand U10711 (N_10711,N_7425,N_8260);
nor U10712 (N_10712,N_7712,N_8660);
nor U10713 (N_10713,N_7219,N_6955);
or U10714 (N_10714,N_8992,N_7647);
nor U10715 (N_10715,N_6149,N_6433);
nor U10716 (N_10716,N_6011,N_6579);
or U10717 (N_10717,N_7493,N_8427);
xor U10718 (N_10718,N_7928,N_8986);
xor U10719 (N_10719,N_6203,N_6871);
nor U10720 (N_10720,N_8809,N_7252);
nor U10721 (N_10721,N_6965,N_6579);
nand U10722 (N_10722,N_6853,N_7343);
or U10723 (N_10723,N_6552,N_8683);
or U10724 (N_10724,N_7953,N_6690);
or U10725 (N_10725,N_8756,N_8045);
xnor U10726 (N_10726,N_6408,N_6808);
or U10727 (N_10727,N_6850,N_7883);
and U10728 (N_10728,N_8022,N_6474);
xor U10729 (N_10729,N_6196,N_7324);
and U10730 (N_10730,N_7918,N_6976);
nor U10731 (N_10731,N_6137,N_6138);
nand U10732 (N_10732,N_6991,N_7747);
nor U10733 (N_10733,N_8499,N_8267);
xnor U10734 (N_10734,N_7367,N_6635);
and U10735 (N_10735,N_8868,N_8720);
and U10736 (N_10736,N_7673,N_6065);
and U10737 (N_10737,N_8877,N_7761);
xor U10738 (N_10738,N_6737,N_7068);
or U10739 (N_10739,N_7600,N_7513);
nand U10740 (N_10740,N_7099,N_6713);
nand U10741 (N_10741,N_6516,N_7654);
nand U10742 (N_10742,N_8643,N_6530);
and U10743 (N_10743,N_7932,N_8301);
xnor U10744 (N_10744,N_7781,N_8836);
or U10745 (N_10745,N_6165,N_6132);
or U10746 (N_10746,N_6788,N_7739);
or U10747 (N_10747,N_6019,N_8849);
or U10748 (N_10748,N_8339,N_8287);
nor U10749 (N_10749,N_8976,N_7444);
nor U10750 (N_10750,N_6608,N_6942);
nor U10751 (N_10751,N_7008,N_6255);
xor U10752 (N_10752,N_8978,N_6757);
xor U10753 (N_10753,N_6368,N_6370);
or U10754 (N_10754,N_7693,N_6276);
xnor U10755 (N_10755,N_6595,N_7954);
nor U10756 (N_10756,N_6096,N_6500);
and U10757 (N_10757,N_6381,N_7224);
nor U10758 (N_10758,N_6996,N_6881);
or U10759 (N_10759,N_8835,N_8991);
and U10760 (N_10760,N_6617,N_8645);
nor U10761 (N_10761,N_6610,N_6896);
nand U10762 (N_10762,N_7816,N_7202);
nor U10763 (N_10763,N_6174,N_8676);
xor U10764 (N_10764,N_6665,N_6568);
or U10765 (N_10765,N_6203,N_7920);
and U10766 (N_10766,N_8158,N_8234);
nor U10767 (N_10767,N_7559,N_8368);
nor U10768 (N_10768,N_7863,N_8504);
or U10769 (N_10769,N_8531,N_6855);
or U10770 (N_10770,N_8190,N_8985);
nor U10771 (N_10771,N_6444,N_8031);
nand U10772 (N_10772,N_6208,N_6744);
or U10773 (N_10773,N_7350,N_8516);
or U10774 (N_10774,N_7766,N_8845);
or U10775 (N_10775,N_8588,N_6910);
xor U10776 (N_10776,N_8303,N_7111);
nor U10777 (N_10777,N_8283,N_8180);
and U10778 (N_10778,N_8266,N_6857);
or U10779 (N_10779,N_8995,N_6257);
or U10780 (N_10780,N_7953,N_6464);
nor U10781 (N_10781,N_6878,N_7495);
or U10782 (N_10782,N_6318,N_8235);
nor U10783 (N_10783,N_8360,N_6267);
and U10784 (N_10784,N_6627,N_7470);
and U10785 (N_10785,N_8051,N_7517);
and U10786 (N_10786,N_6836,N_6696);
and U10787 (N_10787,N_6798,N_6725);
nor U10788 (N_10788,N_6321,N_8450);
and U10789 (N_10789,N_6213,N_6726);
nand U10790 (N_10790,N_6617,N_8592);
or U10791 (N_10791,N_8166,N_8590);
and U10792 (N_10792,N_8695,N_6886);
nand U10793 (N_10793,N_7366,N_8527);
nor U10794 (N_10794,N_6858,N_8301);
and U10795 (N_10795,N_8285,N_6550);
nand U10796 (N_10796,N_8362,N_7585);
or U10797 (N_10797,N_8415,N_6803);
nand U10798 (N_10798,N_6346,N_7878);
and U10799 (N_10799,N_6528,N_7946);
or U10800 (N_10800,N_6377,N_7344);
or U10801 (N_10801,N_8499,N_6433);
nor U10802 (N_10802,N_7599,N_8555);
and U10803 (N_10803,N_7072,N_7278);
nor U10804 (N_10804,N_6002,N_7067);
nand U10805 (N_10805,N_8361,N_7126);
or U10806 (N_10806,N_6859,N_6974);
or U10807 (N_10807,N_6988,N_6412);
nor U10808 (N_10808,N_8509,N_6497);
xnor U10809 (N_10809,N_7297,N_8298);
or U10810 (N_10810,N_7381,N_8902);
or U10811 (N_10811,N_6341,N_6925);
or U10812 (N_10812,N_7232,N_8002);
and U10813 (N_10813,N_7780,N_6659);
nand U10814 (N_10814,N_7553,N_8090);
nor U10815 (N_10815,N_6201,N_6389);
and U10816 (N_10816,N_6040,N_7975);
and U10817 (N_10817,N_7393,N_8269);
nor U10818 (N_10818,N_6815,N_7773);
nand U10819 (N_10819,N_6901,N_6909);
and U10820 (N_10820,N_6265,N_8489);
nor U10821 (N_10821,N_6018,N_7905);
nand U10822 (N_10822,N_8495,N_6801);
nor U10823 (N_10823,N_7375,N_6915);
or U10824 (N_10824,N_8752,N_8250);
nor U10825 (N_10825,N_8017,N_7465);
nand U10826 (N_10826,N_7450,N_6024);
nor U10827 (N_10827,N_7570,N_8390);
nand U10828 (N_10828,N_6540,N_7493);
and U10829 (N_10829,N_7408,N_6835);
nor U10830 (N_10830,N_7381,N_8738);
or U10831 (N_10831,N_6281,N_6047);
and U10832 (N_10832,N_7360,N_7469);
nand U10833 (N_10833,N_8316,N_8067);
and U10834 (N_10834,N_7176,N_7343);
xnor U10835 (N_10835,N_6990,N_6893);
and U10836 (N_10836,N_8101,N_8650);
nor U10837 (N_10837,N_8361,N_6216);
nand U10838 (N_10838,N_8512,N_6098);
and U10839 (N_10839,N_6515,N_7206);
nor U10840 (N_10840,N_7936,N_8047);
or U10841 (N_10841,N_7606,N_8145);
nor U10842 (N_10842,N_6210,N_6875);
xor U10843 (N_10843,N_7839,N_8905);
or U10844 (N_10844,N_6280,N_6667);
nor U10845 (N_10845,N_6124,N_8491);
nor U10846 (N_10846,N_7291,N_6660);
nor U10847 (N_10847,N_6594,N_8130);
nor U10848 (N_10848,N_6393,N_8599);
and U10849 (N_10849,N_6874,N_6167);
nand U10850 (N_10850,N_7836,N_8764);
nand U10851 (N_10851,N_6535,N_7081);
nand U10852 (N_10852,N_6644,N_6075);
xnor U10853 (N_10853,N_8148,N_8829);
nand U10854 (N_10854,N_8547,N_6261);
nor U10855 (N_10855,N_7062,N_6221);
xnor U10856 (N_10856,N_7302,N_7841);
nor U10857 (N_10857,N_7378,N_7937);
or U10858 (N_10858,N_7572,N_7707);
nand U10859 (N_10859,N_8813,N_6826);
xor U10860 (N_10860,N_7172,N_7242);
nand U10861 (N_10861,N_7878,N_7002);
nand U10862 (N_10862,N_7154,N_7577);
nand U10863 (N_10863,N_7201,N_8860);
or U10864 (N_10864,N_7529,N_7499);
nand U10865 (N_10865,N_8847,N_7948);
and U10866 (N_10866,N_8060,N_7776);
nor U10867 (N_10867,N_6339,N_7788);
and U10868 (N_10868,N_6422,N_7664);
and U10869 (N_10869,N_7346,N_6081);
or U10870 (N_10870,N_8431,N_8036);
and U10871 (N_10871,N_7393,N_6191);
nand U10872 (N_10872,N_7043,N_8612);
nand U10873 (N_10873,N_7040,N_6104);
nand U10874 (N_10874,N_8895,N_7478);
xor U10875 (N_10875,N_8268,N_7864);
nor U10876 (N_10876,N_7249,N_6499);
or U10877 (N_10877,N_8627,N_8625);
and U10878 (N_10878,N_7936,N_6846);
nand U10879 (N_10879,N_8136,N_8928);
nand U10880 (N_10880,N_7310,N_6903);
and U10881 (N_10881,N_7635,N_7497);
and U10882 (N_10882,N_6566,N_7901);
nand U10883 (N_10883,N_8541,N_8431);
nor U10884 (N_10884,N_8177,N_7828);
and U10885 (N_10885,N_6236,N_7431);
xnor U10886 (N_10886,N_6421,N_8732);
and U10887 (N_10887,N_7497,N_6217);
and U10888 (N_10888,N_8480,N_7931);
nand U10889 (N_10889,N_6826,N_8181);
or U10890 (N_10890,N_7049,N_6178);
xor U10891 (N_10891,N_8958,N_6477);
or U10892 (N_10892,N_6629,N_7979);
and U10893 (N_10893,N_8961,N_7477);
and U10894 (N_10894,N_7476,N_7722);
xnor U10895 (N_10895,N_7015,N_7284);
xor U10896 (N_10896,N_6978,N_7863);
nand U10897 (N_10897,N_7570,N_8169);
and U10898 (N_10898,N_6948,N_6086);
and U10899 (N_10899,N_7041,N_8531);
xor U10900 (N_10900,N_7139,N_7348);
or U10901 (N_10901,N_6748,N_6198);
nand U10902 (N_10902,N_6146,N_8885);
xnor U10903 (N_10903,N_8840,N_8493);
nand U10904 (N_10904,N_7449,N_6125);
nor U10905 (N_10905,N_6269,N_7210);
or U10906 (N_10906,N_7006,N_8934);
and U10907 (N_10907,N_7965,N_7248);
nand U10908 (N_10908,N_8060,N_6422);
nor U10909 (N_10909,N_6276,N_8716);
nor U10910 (N_10910,N_8505,N_6765);
nand U10911 (N_10911,N_8834,N_8587);
nor U10912 (N_10912,N_7356,N_8539);
or U10913 (N_10913,N_8790,N_8074);
and U10914 (N_10914,N_7940,N_7749);
nand U10915 (N_10915,N_7422,N_7219);
nand U10916 (N_10916,N_8437,N_7269);
nor U10917 (N_10917,N_7824,N_8266);
and U10918 (N_10918,N_6847,N_7530);
nor U10919 (N_10919,N_6019,N_7563);
or U10920 (N_10920,N_7419,N_7486);
nand U10921 (N_10921,N_7603,N_8412);
xnor U10922 (N_10922,N_8543,N_6415);
nand U10923 (N_10923,N_7489,N_6560);
xor U10924 (N_10924,N_6059,N_8022);
nor U10925 (N_10925,N_7025,N_6174);
nor U10926 (N_10926,N_7288,N_6772);
and U10927 (N_10927,N_8736,N_8634);
nor U10928 (N_10928,N_7744,N_7054);
xnor U10929 (N_10929,N_8455,N_6777);
nor U10930 (N_10930,N_8259,N_8450);
nor U10931 (N_10931,N_6353,N_6996);
or U10932 (N_10932,N_8216,N_8047);
or U10933 (N_10933,N_7778,N_7238);
and U10934 (N_10934,N_7243,N_7200);
nand U10935 (N_10935,N_7198,N_6550);
and U10936 (N_10936,N_7000,N_8715);
nor U10937 (N_10937,N_6848,N_6923);
or U10938 (N_10938,N_8271,N_7783);
nor U10939 (N_10939,N_8026,N_8303);
and U10940 (N_10940,N_7297,N_8670);
nor U10941 (N_10941,N_6611,N_6093);
and U10942 (N_10942,N_7355,N_6255);
or U10943 (N_10943,N_7599,N_7276);
and U10944 (N_10944,N_6812,N_7087);
nand U10945 (N_10945,N_7740,N_8843);
or U10946 (N_10946,N_8730,N_8073);
or U10947 (N_10947,N_7273,N_7336);
and U10948 (N_10948,N_6955,N_6208);
or U10949 (N_10949,N_6683,N_8129);
or U10950 (N_10950,N_7305,N_8834);
or U10951 (N_10951,N_6610,N_7865);
or U10952 (N_10952,N_7452,N_6640);
or U10953 (N_10953,N_8606,N_6488);
or U10954 (N_10954,N_8200,N_7036);
or U10955 (N_10955,N_7043,N_7908);
nand U10956 (N_10956,N_6263,N_8827);
and U10957 (N_10957,N_6358,N_8015);
or U10958 (N_10958,N_6976,N_7947);
nor U10959 (N_10959,N_6965,N_7292);
and U10960 (N_10960,N_8599,N_6002);
or U10961 (N_10961,N_6365,N_6015);
nand U10962 (N_10962,N_7672,N_7664);
nor U10963 (N_10963,N_8760,N_7379);
and U10964 (N_10964,N_6124,N_7535);
and U10965 (N_10965,N_6835,N_6672);
nor U10966 (N_10966,N_7013,N_8732);
nor U10967 (N_10967,N_7364,N_6701);
or U10968 (N_10968,N_8269,N_6388);
nor U10969 (N_10969,N_6738,N_8424);
nand U10970 (N_10970,N_8630,N_7558);
nand U10971 (N_10971,N_6070,N_7266);
or U10972 (N_10972,N_7081,N_6133);
or U10973 (N_10973,N_8307,N_7749);
nor U10974 (N_10974,N_7578,N_8624);
nor U10975 (N_10975,N_6607,N_7936);
or U10976 (N_10976,N_7196,N_8578);
or U10977 (N_10977,N_7406,N_8621);
or U10978 (N_10978,N_8062,N_6923);
xor U10979 (N_10979,N_7076,N_8640);
nand U10980 (N_10980,N_6497,N_6627);
nor U10981 (N_10981,N_8628,N_8626);
or U10982 (N_10982,N_6232,N_7703);
nor U10983 (N_10983,N_8328,N_6747);
xnor U10984 (N_10984,N_7787,N_6940);
nor U10985 (N_10985,N_7268,N_8318);
and U10986 (N_10986,N_7988,N_6821);
and U10987 (N_10987,N_6365,N_8080);
or U10988 (N_10988,N_8235,N_7978);
or U10989 (N_10989,N_7086,N_6691);
xor U10990 (N_10990,N_6940,N_8254);
nand U10991 (N_10991,N_6956,N_6487);
nor U10992 (N_10992,N_6970,N_8995);
or U10993 (N_10993,N_7529,N_8098);
nor U10994 (N_10994,N_8109,N_8799);
nor U10995 (N_10995,N_8532,N_7068);
nand U10996 (N_10996,N_6899,N_8843);
xor U10997 (N_10997,N_8474,N_6696);
and U10998 (N_10998,N_6550,N_6022);
and U10999 (N_10999,N_8702,N_6998);
nand U11000 (N_11000,N_8859,N_7048);
and U11001 (N_11001,N_6538,N_6754);
and U11002 (N_11002,N_7040,N_7673);
and U11003 (N_11003,N_6198,N_6942);
or U11004 (N_11004,N_6389,N_7235);
xnor U11005 (N_11005,N_8775,N_6537);
or U11006 (N_11006,N_6493,N_8495);
nand U11007 (N_11007,N_7732,N_7366);
nor U11008 (N_11008,N_8020,N_7299);
xnor U11009 (N_11009,N_8037,N_8138);
or U11010 (N_11010,N_7686,N_7847);
nand U11011 (N_11011,N_6188,N_8460);
nand U11012 (N_11012,N_8236,N_8536);
and U11013 (N_11013,N_6570,N_8206);
and U11014 (N_11014,N_6465,N_8206);
and U11015 (N_11015,N_6552,N_7990);
or U11016 (N_11016,N_6285,N_6119);
nand U11017 (N_11017,N_8970,N_7120);
or U11018 (N_11018,N_6493,N_8633);
or U11019 (N_11019,N_7124,N_6572);
and U11020 (N_11020,N_7972,N_7577);
nor U11021 (N_11021,N_7139,N_7749);
and U11022 (N_11022,N_8718,N_6586);
or U11023 (N_11023,N_7412,N_7448);
nand U11024 (N_11024,N_8731,N_7656);
or U11025 (N_11025,N_7357,N_7019);
and U11026 (N_11026,N_8716,N_8241);
or U11027 (N_11027,N_6691,N_8294);
nand U11028 (N_11028,N_8275,N_6687);
nand U11029 (N_11029,N_7373,N_7639);
nor U11030 (N_11030,N_8964,N_7486);
nand U11031 (N_11031,N_6406,N_8480);
nand U11032 (N_11032,N_6152,N_8147);
and U11033 (N_11033,N_8692,N_7393);
nor U11034 (N_11034,N_7341,N_8121);
nand U11035 (N_11035,N_7208,N_6707);
xor U11036 (N_11036,N_6829,N_8903);
xor U11037 (N_11037,N_6001,N_6546);
or U11038 (N_11038,N_6482,N_7616);
xnor U11039 (N_11039,N_7859,N_7148);
nand U11040 (N_11040,N_7299,N_7779);
and U11041 (N_11041,N_8298,N_7866);
nand U11042 (N_11042,N_7758,N_7708);
nand U11043 (N_11043,N_6091,N_7790);
nand U11044 (N_11044,N_8163,N_8345);
and U11045 (N_11045,N_6180,N_8585);
or U11046 (N_11046,N_7803,N_8983);
and U11047 (N_11047,N_6349,N_7446);
xor U11048 (N_11048,N_6929,N_6872);
nor U11049 (N_11049,N_7256,N_7837);
or U11050 (N_11050,N_6678,N_8788);
or U11051 (N_11051,N_8436,N_8525);
and U11052 (N_11052,N_8113,N_8638);
and U11053 (N_11053,N_8105,N_8335);
or U11054 (N_11054,N_8285,N_8480);
nor U11055 (N_11055,N_7629,N_7892);
or U11056 (N_11056,N_6841,N_7592);
nor U11057 (N_11057,N_7424,N_7574);
nand U11058 (N_11058,N_7439,N_7028);
nand U11059 (N_11059,N_8396,N_7628);
and U11060 (N_11060,N_8054,N_8747);
nor U11061 (N_11061,N_7114,N_6304);
xnor U11062 (N_11062,N_8094,N_6198);
or U11063 (N_11063,N_7429,N_6765);
nor U11064 (N_11064,N_7459,N_7737);
and U11065 (N_11065,N_7614,N_6613);
nor U11066 (N_11066,N_6122,N_6435);
or U11067 (N_11067,N_6504,N_8463);
nor U11068 (N_11068,N_7715,N_7574);
and U11069 (N_11069,N_6243,N_7930);
nand U11070 (N_11070,N_7552,N_7086);
and U11071 (N_11071,N_7014,N_8584);
nor U11072 (N_11072,N_6533,N_8515);
or U11073 (N_11073,N_6089,N_7433);
and U11074 (N_11074,N_7021,N_6632);
and U11075 (N_11075,N_8363,N_7636);
nor U11076 (N_11076,N_6209,N_8708);
or U11077 (N_11077,N_8707,N_6252);
nor U11078 (N_11078,N_6986,N_8576);
or U11079 (N_11079,N_7881,N_8798);
nand U11080 (N_11080,N_8380,N_7180);
nor U11081 (N_11081,N_6852,N_6742);
nand U11082 (N_11082,N_8375,N_6386);
and U11083 (N_11083,N_7646,N_8662);
nor U11084 (N_11084,N_7694,N_6132);
nor U11085 (N_11085,N_8912,N_8157);
or U11086 (N_11086,N_6556,N_8677);
or U11087 (N_11087,N_8701,N_6093);
nor U11088 (N_11088,N_7194,N_6891);
nor U11089 (N_11089,N_7736,N_8595);
nor U11090 (N_11090,N_6353,N_8601);
and U11091 (N_11091,N_8297,N_6383);
or U11092 (N_11092,N_6466,N_6952);
or U11093 (N_11093,N_8760,N_8099);
nor U11094 (N_11094,N_8307,N_8990);
nor U11095 (N_11095,N_7438,N_6771);
nor U11096 (N_11096,N_6877,N_7147);
nor U11097 (N_11097,N_8968,N_7288);
nand U11098 (N_11098,N_6604,N_6589);
nor U11099 (N_11099,N_6154,N_6861);
xor U11100 (N_11100,N_7775,N_7612);
and U11101 (N_11101,N_6101,N_6330);
nand U11102 (N_11102,N_6620,N_8477);
or U11103 (N_11103,N_8512,N_6038);
and U11104 (N_11104,N_6324,N_6833);
xor U11105 (N_11105,N_8887,N_6713);
nor U11106 (N_11106,N_7310,N_8004);
nor U11107 (N_11107,N_6716,N_7891);
nor U11108 (N_11108,N_8882,N_6251);
or U11109 (N_11109,N_8003,N_6267);
nand U11110 (N_11110,N_6054,N_7581);
nor U11111 (N_11111,N_8082,N_8769);
nor U11112 (N_11112,N_8087,N_7004);
and U11113 (N_11113,N_7698,N_8243);
or U11114 (N_11114,N_7390,N_8826);
nor U11115 (N_11115,N_7136,N_8695);
nor U11116 (N_11116,N_6719,N_6215);
nor U11117 (N_11117,N_6951,N_7019);
nand U11118 (N_11118,N_6909,N_8958);
xnor U11119 (N_11119,N_6071,N_6196);
xnor U11120 (N_11120,N_8264,N_6024);
and U11121 (N_11121,N_8279,N_6980);
nand U11122 (N_11122,N_6877,N_7135);
nand U11123 (N_11123,N_6717,N_7088);
xnor U11124 (N_11124,N_8977,N_8410);
nor U11125 (N_11125,N_8292,N_6071);
and U11126 (N_11126,N_7592,N_8978);
nand U11127 (N_11127,N_8046,N_6890);
nor U11128 (N_11128,N_7741,N_6314);
nand U11129 (N_11129,N_8568,N_8475);
and U11130 (N_11130,N_8804,N_8085);
or U11131 (N_11131,N_6057,N_6026);
nand U11132 (N_11132,N_6065,N_8525);
and U11133 (N_11133,N_7083,N_8968);
or U11134 (N_11134,N_8323,N_7169);
or U11135 (N_11135,N_6574,N_8567);
and U11136 (N_11136,N_8869,N_8457);
or U11137 (N_11137,N_7662,N_8036);
nand U11138 (N_11138,N_8276,N_6275);
nand U11139 (N_11139,N_6924,N_7956);
xnor U11140 (N_11140,N_6503,N_6641);
and U11141 (N_11141,N_8036,N_7450);
nand U11142 (N_11142,N_7639,N_8645);
and U11143 (N_11143,N_6922,N_7399);
nand U11144 (N_11144,N_6692,N_6976);
nor U11145 (N_11145,N_8751,N_6753);
nand U11146 (N_11146,N_8391,N_6999);
and U11147 (N_11147,N_6738,N_7744);
xor U11148 (N_11148,N_8409,N_7814);
nor U11149 (N_11149,N_8904,N_7373);
and U11150 (N_11150,N_8688,N_7882);
nand U11151 (N_11151,N_8664,N_6223);
nand U11152 (N_11152,N_6508,N_8410);
or U11153 (N_11153,N_6844,N_6535);
or U11154 (N_11154,N_8389,N_8423);
nand U11155 (N_11155,N_7922,N_8231);
nand U11156 (N_11156,N_7645,N_6138);
xnor U11157 (N_11157,N_6185,N_7302);
nand U11158 (N_11158,N_8841,N_8557);
nand U11159 (N_11159,N_8250,N_8866);
nor U11160 (N_11160,N_8321,N_8099);
or U11161 (N_11161,N_7684,N_6102);
nor U11162 (N_11162,N_6247,N_6533);
and U11163 (N_11163,N_7427,N_7994);
nand U11164 (N_11164,N_7290,N_6612);
and U11165 (N_11165,N_7761,N_6609);
and U11166 (N_11166,N_7407,N_7149);
and U11167 (N_11167,N_8473,N_6729);
xor U11168 (N_11168,N_8829,N_7208);
and U11169 (N_11169,N_8675,N_6376);
or U11170 (N_11170,N_6012,N_8709);
and U11171 (N_11171,N_8828,N_6354);
and U11172 (N_11172,N_7235,N_6493);
and U11173 (N_11173,N_7172,N_8200);
and U11174 (N_11174,N_6825,N_7606);
nand U11175 (N_11175,N_6755,N_8789);
and U11176 (N_11176,N_7976,N_7779);
or U11177 (N_11177,N_7713,N_8847);
and U11178 (N_11178,N_7984,N_6952);
and U11179 (N_11179,N_8331,N_6095);
or U11180 (N_11180,N_8440,N_7060);
or U11181 (N_11181,N_6561,N_8722);
nor U11182 (N_11182,N_8805,N_7451);
and U11183 (N_11183,N_8358,N_7885);
or U11184 (N_11184,N_6088,N_7351);
and U11185 (N_11185,N_6082,N_6667);
nor U11186 (N_11186,N_6532,N_6702);
nand U11187 (N_11187,N_8461,N_6165);
nor U11188 (N_11188,N_7343,N_8795);
or U11189 (N_11189,N_7675,N_8020);
nand U11190 (N_11190,N_8378,N_8456);
and U11191 (N_11191,N_6971,N_6173);
and U11192 (N_11192,N_7928,N_8659);
xor U11193 (N_11193,N_8803,N_8043);
and U11194 (N_11194,N_8992,N_8522);
and U11195 (N_11195,N_8637,N_6830);
and U11196 (N_11196,N_7144,N_6867);
or U11197 (N_11197,N_8338,N_6610);
or U11198 (N_11198,N_6459,N_8527);
or U11199 (N_11199,N_6478,N_7204);
nand U11200 (N_11200,N_6576,N_6611);
or U11201 (N_11201,N_7079,N_6009);
and U11202 (N_11202,N_6490,N_7399);
nor U11203 (N_11203,N_6932,N_7661);
nor U11204 (N_11204,N_6508,N_7343);
nor U11205 (N_11205,N_8684,N_6063);
xor U11206 (N_11206,N_7983,N_8796);
nor U11207 (N_11207,N_7507,N_8731);
nand U11208 (N_11208,N_6106,N_8161);
nor U11209 (N_11209,N_8584,N_8572);
nor U11210 (N_11210,N_7983,N_8418);
nand U11211 (N_11211,N_6921,N_6094);
nor U11212 (N_11212,N_7933,N_6792);
and U11213 (N_11213,N_6324,N_6506);
nor U11214 (N_11214,N_6536,N_7708);
or U11215 (N_11215,N_7801,N_6503);
or U11216 (N_11216,N_6658,N_8445);
xor U11217 (N_11217,N_8257,N_7561);
or U11218 (N_11218,N_7031,N_7165);
or U11219 (N_11219,N_8414,N_6427);
or U11220 (N_11220,N_7104,N_7718);
xor U11221 (N_11221,N_8502,N_7071);
nor U11222 (N_11222,N_7065,N_7059);
or U11223 (N_11223,N_6655,N_7721);
and U11224 (N_11224,N_6704,N_8080);
and U11225 (N_11225,N_6770,N_8889);
nand U11226 (N_11226,N_7721,N_7126);
nor U11227 (N_11227,N_8218,N_8993);
and U11228 (N_11228,N_8901,N_6770);
and U11229 (N_11229,N_8633,N_6081);
nor U11230 (N_11230,N_7441,N_7571);
and U11231 (N_11231,N_8607,N_7829);
nor U11232 (N_11232,N_6731,N_8769);
or U11233 (N_11233,N_8618,N_7989);
nor U11234 (N_11234,N_6367,N_7006);
and U11235 (N_11235,N_8961,N_7696);
nand U11236 (N_11236,N_6534,N_7302);
nand U11237 (N_11237,N_6306,N_6241);
nand U11238 (N_11238,N_7026,N_6742);
or U11239 (N_11239,N_6573,N_7192);
and U11240 (N_11240,N_8377,N_8865);
nor U11241 (N_11241,N_6949,N_8787);
nor U11242 (N_11242,N_6169,N_7292);
or U11243 (N_11243,N_8382,N_8627);
nand U11244 (N_11244,N_8072,N_6225);
and U11245 (N_11245,N_7306,N_6878);
nor U11246 (N_11246,N_6296,N_6038);
and U11247 (N_11247,N_6228,N_6635);
nor U11248 (N_11248,N_7272,N_6173);
and U11249 (N_11249,N_8534,N_6702);
or U11250 (N_11250,N_8881,N_8427);
nor U11251 (N_11251,N_8468,N_8712);
nand U11252 (N_11252,N_6878,N_7029);
and U11253 (N_11253,N_8791,N_8858);
nand U11254 (N_11254,N_6466,N_6830);
nand U11255 (N_11255,N_7401,N_6296);
nor U11256 (N_11256,N_6944,N_6046);
and U11257 (N_11257,N_7389,N_7417);
or U11258 (N_11258,N_7421,N_6404);
nand U11259 (N_11259,N_7066,N_7334);
or U11260 (N_11260,N_6125,N_7379);
and U11261 (N_11261,N_6861,N_8908);
xnor U11262 (N_11262,N_6764,N_8297);
or U11263 (N_11263,N_7977,N_7581);
and U11264 (N_11264,N_6920,N_6105);
nand U11265 (N_11265,N_6324,N_7637);
xnor U11266 (N_11266,N_8737,N_6771);
nand U11267 (N_11267,N_6362,N_6180);
xnor U11268 (N_11268,N_7676,N_7452);
nand U11269 (N_11269,N_7666,N_7109);
or U11270 (N_11270,N_8323,N_8020);
or U11271 (N_11271,N_7652,N_7568);
and U11272 (N_11272,N_6003,N_8896);
nor U11273 (N_11273,N_7666,N_7031);
and U11274 (N_11274,N_6418,N_6980);
or U11275 (N_11275,N_8885,N_7151);
nand U11276 (N_11276,N_7675,N_6083);
or U11277 (N_11277,N_8103,N_6878);
nand U11278 (N_11278,N_6706,N_8891);
and U11279 (N_11279,N_8710,N_7995);
or U11280 (N_11280,N_7257,N_8351);
and U11281 (N_11281,N_6756,N_7414);
and U11282 (N_11282,N_7688,N_8794);
nor U11283 (N_11283,N_6730,N_6346);
and U11284 (N_11284,N_8021,N_7888);
nor U11285 (N_11285,N_7359,N_7619);
nand U11286 (N_11286,N_6747,N_7514);
or U11287 (N_11287,N_7518,N_7629);
nand U11288 (N_11288,N_7747,N_7330);
and U11289 (N_11289,N_7597,N_7188);
and U11290 (N_11290,N_7278,N_7061);
and U11291 (N_11291,N_6438,N_6524);
nand U11292 (N_11292,N_7720,N_7520);
nor U11293 (N_11293,N_6506,N_8615);
nand U11294 (N_11294,N_7433,N_7168);
or U11295 (N_11295,N_6546,N_8291);
and U11296 (N_11296,N_8047,N_8728);
or U11297 (N_11297,N_8727,N_7149);
or U11298 (N_11298,N_6132,N_8786);
nor U11299 (N_11299,N_6738,N_7043);
nand U11300 (N_11300,N_6659,N_8966);
nand U11301 (N_11301,N_6441,N_8329);
xor U11302 (N_11302,N_8326,N_6787);
xnor U11303 (N_11303,N_7781,N_6258);
nor U11304 (N_11304,N_7022,N_6662);
and U11305 (N_11305,N_7996,N_6322);
nand U11306 (N_11306,N_7664,N_8836);
or U11307 (N_11307,N_6692,N_8370);
nand U11308 (N_11308,N_8356,N_7962);
nand U11309 (N_11309,N_7595,N_8619);
nand U11310 (N_11310,N_7217,N_7245);
nor U11311 (N_11311,N_8875,N_7535);
nor U11312 (N_11312,N_6951,N_7509);
and U11313 (N_11313,N_6532,N_8873);
nor U11314 (N_11314,N_7749,N_8691);
nand U11315 (N_11315,N_6341,N_7498);
nor U11316 (N_11316,N_6911,N_6595);
nor U11317 (N_11317,N_8014,N_7923);
or U11318 (N_11318,N_6902,N_6313);
xnor U11319 (N_11319,N_8928,N_6918);
and U11320 (N_11320,N_8725,N_7838);
nand U11321 (N_11321,N_7549,N_7124);
or U11322 (N_11322,N_6007,N_6054);
and U11323 (N_11323,N_7530,N_7806);
nand U11324 (N_11324,N_7988,N_6842);
or U11325 (N_11325,N_7964,N_8394);
nor U11326 (N_11326,N_8563,N_6494);
and U11327 (N_11327,N_7874,N_6134);
nor U11328 (N_11328,N_8173,N_6789);
nor U11329 (N_11329,N_6345,N_7524);
and U11330 (N_11330,N_6409,N_7229);
and U11331 (N_11331,N_8940,N_6841);
and U11332 (N_11332,N_7107,N_8992);
nand U11333 (N_11333,N_7661,N_8443);
and U11334 (N_11334,N_7757,N_6620);
or U11335 (N_11335,N_8459,N_7009);
nand U11336 (N_11336,N_8869,N_7858);
or U11337 (N_11337,N_6258,N_7110);
nor U11338 (N_11338,N_7522,N_7737);
and U11339 (N_11339,N_8593,N_8484);
nand U11340 (N_11340,N_8630,N_8490);
nor U11341 (N_11341,N_7078,N_6923);
nand U11342 (N_11342,N_8114,N_6076);
nand U11343 (N_11343,N_6742,N_8919);
nand U11344 (N_11344,N_6763,N_7312);
or U11345 (N_11345,N_8560,N_7263);
nor U11346 (N_11346,N_8336,N_8662);
or U11347 (N_11347,N_8209,N_7855);
or U11348 (N_11348,N_7117,N_8063);
or U11349 (N_11349,N_6311,N_6797);
nor U11350 (N_11350,N_7779,N_7184);
or U11351 (N_11351,N_6180,N_8907);
or U11352 (N_11352,N_6296,N_7873);
or U11353 (N_11353,N_7071,N_6195);
nand U11354 (N_11354,N_7089,N_7123);
nor U11355 (N_11355,N_7106,N_8907);
and U11356 (N_11356,N_6578,N_6424);
nor U11357 (N_11357,N_6546,N_7833);
or U11358 (N_11358,N_7081,N_7425);
and U11359 (N_11359,N_7929,N_8624);
nand U11360 (N_11360,N_8804,N_6017);
and U11361 (N_11361,N_8136,N_8977);
nand U11362 (N_11362,N_8599,N_7929);
or U11363 (N_11363,N_6126,N_6051);
nand U11364 (N_11364,N_6817,N_6326);
xnor U11365 (N_11365,N_6181,N_7002);
nor U11366 (N_11366,N_6601,N_8050);
nor U11367 (N_11367,N_8814,N_6319);
xnor U11368 (N_11368,N_8542,N_6240);
nor U11369 (N_11369,N_8341,N_7206);
nor U11370 (N_11370,N_6487,N_8801);
nor U11371 (N_11371,N_6873,N_6007);
nand U11372 (N_11372,N_6301,N_6281);
nand U11373 (N_11373,N_8415,N_7172);
nand U11374 (N_11374,N_7823,N_8054);
nand U11375 (N_11375,N_6956,N_6755);
xnor U11376 (N_11376,N_6192,N_8964);
xnor U11377 (N_11377,N_8479,N_7638);
nand U11378 (N_11378,N_6018,N_8861);
xor U11379 (N_11379,N_6335,N_8983);
or U11380 (N_11380,N_8754,N_6944);
and U11381 (N_11381,N_7458,N_8468);
nor U11382 (N_11382,N_6744,N_8797);
or U11383 (N_11383,N_6570,N_7275);
nor U11384 (N_11384,N_8010,N_7418);
xnor U11385 (N_11385,N_7525,N_8818);
or U11386 (N_11386,N_7084,N_6414);
and U11387 (N_11387,N_6601,N_6857);
or U11388 (N_11388,N_6911,N_8595);
nor U11389 (N_11389,N_7709,N_8567);
nand U11390 (N_11390,N_6892,N_7659);
and U11391 (N_11391,N_7152,N_8848);
and U11392 (N_11392,N_7220,N_7251);
xnor U11393 (N_11393,N_8936,N_6148);
or U11394 (N_11394,N_8055,N_8797);
nand U11395 (N_11395,N_8654,N_8793);
nand U11396 (N_11396,N_8896,N_6130);
xor U11397 (N_11397,N_6913,N_7147);
xnor U11398 (N_11398,N_6801,N_8983);
nor U11399 (N_11399,N_8716,N_8319);
or U11400 (N_11400,N_6825,N_6808);
xnor U11401 (N_11401,N_6519,N_6879);
and U11402 (N_11402,N_6460,N_8949);
nor U11403 (N_11403,N_7880,N_6629);
and U11404 (N_11404,N_6930,N_6872);
nand U11405 (N_11405,N_7702,N_6767);
nand U11406 (N_11406,N_7074,N_8999);
or U11407 (N_11407,N_7334,N_8555);
or U11408 (N_11408,N_8522,N_7014);
and U11409 (N_11409,N_7112,N_6024);
and U11410 (N_11410,N_8139,N_8692);
or U11411 (N_11411,N_7073,N_7063);
or U11412 (N_11412,N_6535,N_8016);
nand U11413 (N_11413,N_7055,N_6358);
or U11414 (N_11414,N_6499,N_8881);
nor U11415 (N_11415,N_6846,N_6008);
nor U11416 (N_11416,N_7106,N_6375);
or U11417 (N_11417,N_6141,N_8834);
nor U11418 (N_11418,N_7212,N_8137);
or U11419 (N_11419,N_8515,N_8195);
or U11420 (N_11420,N_6970,N_6728);
or U11421 (N_11421,N_7327,N_6379);
nor U11422 (N_11422,N_7127,N_6440);
nor U11423 (N_11423,N_7879,N_6435);
nand U11424 (N_11424,N_8687,N_7917);
nor U11425 (N_11425,N_7250,N_6923);
and U11426 (N_11426,N_7457,N_8305);
nor U11427 (N_11427,N_8883,N_6469);
or U11428 (N_11428,N_7293,N_7246);
nor U11429 (N_11429,N_6187,N_6130);
or U11430 (N_11430,N_7221,N_6434);
nor U11431 (N_11431,N_6574,N_7973);
and U11432 (N_11432,N_7425,N_7546);
and U11433 (N_11433,N_8301,N_6157);
xnor U11434 (N_11434,N_6624,N_7415);
or U11435 (N_11435,N_7400,N_8741);
xnor U11436 (N_11436,N_6096,N_6902);
xnor U11437 (N_11437,N_6146,N_7113);
nand U11438 (N_11438,N_8770,N_8531);
nor U11439 (N_11439,N_7606,N_7318);
xor U11440 (N_11440,N_7445,N_6857);
nor U11441 (N_11441,N_8329,N_8705);
and U11442 (N_11442,N_7061,N_8315);
nand U11443 (N_11443,N_7391,N_6674);
and U11444 (N_11444,N_6705,N_8738);
and U11445 (N_11445,N_6362,N_6812);
xnor U11446 (N_11446,N_7373,N_8210);
xor U11447 (N_11447,N_7668,N_6315);
nand U11448 (N_11448,N_6227,N_8499);
xor U11449 (N_11449,N_7456,N_6421);
nor U11450 (N_11450,N_8699,N_6088);
xnor U11451 (N_11451,N_8161,N_6985);
nor U11452 (N_11452,N_8724,N_7968);
xnor U11453 (N_11453,N_6767,N_8747);
or U11454 (N_11454,N_6343,N_8780);
nand U11455 (N_11455,N_6708,N_7497);
nor U11456 (N_11456,N_6281,N_8999);
xnor U11457 (N_11457,N_8063,N_8387);
xor U11458 (N_11458,N_7238,N_6597);
xor U11459 (N_11459,N_6951,N_7244);
nand U11460 (N_11460,N_7834,N_8968);
nor U11461 (N_11461,N_8945,N_8480);
nand U11462 (N_11462,N_6467,N_7896);
and U11463 (N_11463,N_6242,N_8226);
or U11464 (N_11464,N_7323,N_7388);
or U11465 (N_11465,N_7522,N_6716);
and U11466 (N_11466,N_6411,N_8469);
and U11467 (N_11467,N_8608,N_7159);
nor U11468 (N_11468,N_6432,N_7924);
and U11469 (N_11469,N_7921,N_6373);
nor U11470 (N_11470,N_6792,N_6022);
nor U11471 (N_11471,N_7303,N_7336);
nand U11472 (N_11472,N_7615,N_8043);
or U11473 (N_11473,N_8592,N_8348);
nand U11474 (N_11474,N_7008,N_6767);
and U11475 (N_11475,N_7824,N_8265);
or U11476 (N_11476,N_6643,N_7704);
and U11477 (N_11477,N_6211,N_6067);
or U11478 (N_11478,N_8613,N_6543);
nand U11479 (N_11479,N_7593,N_6485);
or U11480 (N_11480,N_8664,N_8033);
nor U11481 (N_11481,N_8179,N_7095);
xnor U11482 (N_11482,N_6685,N_8224);
nand U11483 (N_11483,N_8400,N_8876);
and U11484 (N_11484,N_8184,N_8305);
nand U11485 (N_11485,N_7217,N_8799);
and U11486 (N_11486,N_8373,N_7755);
nor U11487 (N_11487,N_6091,N_6670);
and U11488 (N_11488,N_6363,N_8963);
or U11489 (N_11489,N_8810,N_8397);
and U11490 (N_11490,N_7830,N_7825);
and U11491 (N_11491,N_6549,N_8183);
nand U11492 (N_11492,N_6963,N_6997);
or U11493 (N_11493,N_6213,N_8428);
nand U11494 (N_11494,N_6674,N_7065);
nor U11495 (N_11495,N_7030,N_7426);
xor U11496 (N_11496,N_6876,N_6497);
or U11497 (N_11497,N_7063,N_6083);
nand U11498 (N_11498,N_6019,N_8183);
and U11499 (N_11499,N_7408,N_6165);
nor U11500 (N_11500,N_7959,N_7881);
nor U11501 (N_11501,N_7436,N_8597);
or U11502 (N_11502,N_6048,N_6055);
and U11503 (N_11503,N_8258,N_6092);
or U11504 (N_11504,N_7161,N_7876);
and U11505 (N_11505,N_8023,N_6528);
and U11506 (N_11506,N_7709,N_7512);
or U11507 (N_11507,N_6092,N_8625);
xnor U11508 (N_11508,N_6348,N_8680);
xnor U11509 (N_11509,N_7792,N_6948);
and U11510 (N_11510,N_8928,N_8398);
and U11511 (N_11511,N_7318,N_6398);
nand U11512 (N_11512,N_6946,N_8465);
or U11513 (N_11513,N_7297,N_7740);
or U11514 (N_11514,N_8812,N_6429);
nor U11515 (N_11515,N_8496,N_7279);
and U11516 (N_11516,N_8639,N_6408);
and U11517 (N_11517,N_8728,N_8909);
or U11518 (N_11518,N_8325,N_6374);
or U11519 (N_11519,N_8427,N_8037);
or U11520 (N_11520,N_8403,N_6915);
nand U11521 (N_11521,N_7291,N_6182);
nand U11522 (N_11522,N_6261,N_8776);
or U11523 (N_11523,N_6837,N_8075);
and U11524 (N_11524,N_8093,N_7486);
or U11525 (N_11525,N_6911,N_7753);
and U11526 (N_11526,N_6255,N_7089);
nand U11527 (N_11527,N_7033,N_7695);
or U11528 (N_11528,N_6155,N_8233);
and U11529 (N_11529,N_7895,N_8830);
and U11530 (N_11530,N_6850,N_6810);
and U11531 (N_11531,N_8153,N_8852);
nand U11532 (N_11532,N_7720,N_8275);
nand U11533 (N_11533,N_8055,N_6025);
or U11534 (N_11534,N_7253,N_6447);
nor U11535 (N_11535,N_8934,N_6925);
and U11536 (N_11536,N_7563,N_7201);
or U11537 (N_11537,N_8810,N_6581);
nand U11538 (N_11538,N_7595,N_6119);
or U11539 (N_11539,N_7147,N_6924);
or U11540 (N_11540,N_8819,N_8148);
nand U11541 (N_11541,N_6393,N_8683);
xnor U11542 (N_11542,N_6389,N_7669);
or U11543 (N_11543,N_8404,N_6339);
nor U11544 (N_11544,N_6871,N_8989);
and U11545 (N_11545,N_8530,N_7198);
nand U11546 (N_11546,N_6658,N_6456);
or U11547 (N_11547,N_8535,N_8948);
or U11548 (N_11548,N_6695,N_8644);
nor U11549 (N_11549,N_7441,N_6141);
nor U11550 (N_11550,N_7897,N_6719);
nor U11551 (N_11551,N_8211,N_8899);
nor U11552 (N_11552,N_8143,N_7966);
nand U11553 (N_11553,N_8472,N_6583);
and U11554 (N_11554,N_8445,N_7061);
nand U11555 (N_11555,N_7484,N_6020);
or U11556 (N_11556,N_8942,N_7967);
and U11557 (N_11557,N_6610,N_6100);
and U11558 (N_11558,N_8576,N_7140);
and U11559 (N_11559,N_7815,N_8902);
nand U11560 (N_11560,N_8294,N_8033);
and U11561 (N_11561,N_6529,N_6499);
and U11562 (N_11562,N_6660,N_6675);
nand U11563 (N_11563,N_6193,N_8324);
nand U11564 (N_11564,N_8855,N_7508);
or U11565 (N_11565,N_8223,N_6392);
and U11566 (N_11566,N_7366,N_7058);
or U11567 (N_11567,N_7035,N_7001);
or U11568 (N_11568,N_8532,N_6062);
and U11569 (N_11569,N_8391,N_6223);
nor U11570 (N_11570,N_7976,N_8773);
nand U11571 (N_11571,N_6227,N_6202);
xor U11572 (N_11572,N_7960,N_7575);
xnor U11573 (N_11573,N_8281,N_8436);
xor U11574 (N_11574,N_6077,N_6360);
or U11575 (N_11575,N_6079,N_8691);
and U11576 (N_11576,N_8328,N_8674);
nand U11577 (N_11577,N_6718,N_6638);
nor U11578 (N_11578,N_6424,N_8965);
or U11579 (N_11579,N_7594,N_6197);
nand U11580 (N_11580,N_6464,N_6944);
and U11581 (N_11581,N_7457,N_6791);
or U11582 (N_11582,N_8111,N_7431);
or U11583 (N_11583,N_7650,N_6642);
nor U11584 (N_11584,N_7797,N_8304);
or U11585 (N_11585,N_6854,N_6713);
and U11586 (N_11586,N_8959,N_7094);
and U11587 (N_11587,N_8100,N_8261);
nand U11588 (N_11588,N_6271,N_8043);
or U11589 (N_11589,N_6213,N_7392);
and U11590 (N_11590,N_6028,N_7530);
nor U11591 (N_11591,N_8213,N_8512);
xnor U11592 (N_11592,N_6904,N_8941);
or U11593 (N_11593,N_8423,N_8792);
nand U11594 (N_11594,N_8929,N_7106);
or U11595 (N_11595,N_7545,N_6447);
nor U11596 (N_11596,N_8870,N_7828);
xnor U11597 (N_11597,N_7832,N_8683);
nand U11598 (N_11598,N_7181,N_7228);
or U11599 (N_11599,N_8222,N_8662);
nand U11600 (N_11600,N_7900,N_6300);
and U11601 (N_11601,N_8411,N_8337);
xor U11602 (N_11602,N_6796,N_6195);
xor U11603 (N_11603,N_8687,N_7229);
nand U11604 (N_11604,N_6458,N_8808);
or U11605 (N_11605,N_6275,N_6264);
nand U11606 (N_11606,N_6336,N_7706);
or U11607 (N_11607,N_8939,N_7711);
or U11608 (N_11608,N_7501,N_7324);
nand U11609 (N_11609,N_6803,N_8736);
and U11610 (N_11610,N_7858,N_8637);
nand U11611 (N_11611,N_6532,N_8178);
and U11612 (N_11612,N_7642,N_8403);
and U11613 (N_11613,N_8643,N_8230);
nor U11614 (N_11614,N_8184,N_6833);
nor U11615 (N_11615,N_8412,N_6089);
and U11616 (N_11616,N_7806,N_8385);
or U11617 (N_11617,N_7823,N_7524);
and U11618 (N_11618,N_6820,N_8636);
or U11619 (N_11619,N_8443,N_6087);
nor U11620 (N_11620,N_6623,N_6283);
xor U11621 (N_11621,N_6650,N_6620);
nand U11622 (N_11622,N_6158,N_8137);
xor U11623 (N_11623,N_8698,N_6039);
and U11624 (N_11624,N_7700,N_7304);
nand U11625 (N_11625,N_7762,N_6097);
or U11626 (N_11626,N_6521,N_8990);
nor U11627 (N_11627,N_8671,N_6705);
nor U11628 (N_11628,N_6095,N_8572);
nand U11629 (N_11629,N_6754,N_8247);
nor U11630 (N_11630,N_6978,N_7745);
nand U11631 (N_11631,N_6316,N_6246);
nand U11632 (N_11632,N_7182,N_8394);
nand U11633 (N_11633,N_8019,N_7122);
nand U11634 (N_11634,N_8013,N_8481);
or U11635 (N_11635,N_7829,N_6322);
nand U11636 (N_11636,N_7087,N_8634);
and U11637 (N_11637,N_8234,N_7147);
or U11638 (N_11638,N_7769,N_8900);
and U11639 (N_11639,N_6133,N_6379);
and U11640 (N_11640,N_7018,N_7817);
xor U11641 (N_11641,N_7550,N_6752);
or U11642 (N_11642,N_7149,N_8976);
nand U11643 (N_11643,N_7796,N_6719);
xnor U11644 (N_11644,N_7701,N_7607);
and U11645 (N_11645,N_8393,N_7362);
nand U11646 (N_11646,N_8918,N_7531);
or U11647 (N_11647,N_7502,N_6682);
or U11648 (N_11648,N_7791,N_6100);
and U11649 (N_11649,N_6420,N_6441);
xor U11650 (N_11650,N_7954,N_7434);
nand U11651 (N_11651,N_8421,N_7601);
and U11652 (N_11652,N_6336,N_8231);
nand U11653 (N_11653,N_8844,N_8023);
nor U11654 (N_11654,N_8334,N_6505);
nor U11655 (N_11655,N_8785,N_6111);
and U11656 (N_11656,N_7271,N_8705);
nand U11657 (N_11657,N_7190,N_8390);
nor U11658 (N_11658,N_7373,N_6867);
nand U11659 (N_11659,N_6897,N_6581);
nand U11660 (N_11660,N_6506,N_8602);
and U11661 (N_11661,N_6252,N_7854);
and U11662 (N_11662,N_6989,N_6459);
or U11663 (N_11663,N_8585,N_6045);
nand U11664 (N_11664,N_8572,N_6289);
nand U11665 (N_11665,N_7795,N_6504);
xnor U11666 (N_11666,N_6198,N_8305);
nand U11667 (N_11667,N_8156,N_8463);
nor U11668 (N_11668,N_8459,N_6247);
and U11669 (N_11669,N_8354,N_8294);
nor U11670 (N_11670,N_8738,N_6716);
nor U11671 (N_11671,N_7907,N_6266);
nand U11672 (N_11672,N_6909,N_6348);
and U11673 (N_11673,N_7705,N_6749);
or U11674 (N_11674,N_8589,N_7583);
nand U11675 (N_11675,N_7209,N_7064);
nor U11676 (N_11676,N_6641,N_6584);
nand U11677 (N_11677,N_8963,N_6453);
and U11678 (N_11678,N_7488,N_7896);
nand U11679 (N_11679,N_7954,N_7686);
or U11680 (N_11680,N_8744,N_6590);
nand U11681 (N_11681,N_7352,N_7760);
or U11682 (N_11682,N_8454,N_6344);
or U11683 (N_11683,N_8115,N_8347);
nor U11684 (N_11684,N_6975,N_7232);
or U11685 (N_11685,N_6446,N_8045);
and U11686 (N_11686,N_8717,N_6645);
and U11687 (N_11687,N_6920,N_6182);
nor U11688 (N_11688,N_8794,N_8007);
xor U11689 (N_11689,N_7928,N_6024);
or U11690 (N_11690,N_7370,N_8749);
nand U11691 (N_11691,N_7129,N_7669);
nand U11692 (N_11692,N_8144,N_6958);
nor U11693 (N_11693,N_8260,N_8209);
nand U11694 (N_11694,N_8696,N_7549);
and U11695 (N_11695,N_8108,N_7940);
and U11696 (N_11696,N_6842,N_8238);
or U11697 (N_11697,N_7490,N_6597);
nand U11698 (N_11698,N_8675,N_8220);
and U11699 (N_11699,N_8381,N_6963);
and U11700 (N_11700,N_7896,N_8001);
and U11701 (N_11701,N_7595,N_7481);
or U11702 (N_11702,N_6553,N_7111);
nor U11703 (N_11703,N_8513,N_6209);
or U11704 (N_11704,N_8038,N_8227);
nand U11705 (N_11705,N_7263,N_8096);
and U11706 (N_11706,N_8836,N_8477);
nor U11707 (N_11707,N_7041,N_8067);
and U11708 (N_11708,N_6328,N_7357);
or U11709 (N_11709,N_6732,N_7500);
and U11710 (N_11710,N_8922,N_6153);
nor U11711 (N_11711,N_7698,N_8400);
and U11712 (N_11712,N_8930,N_8352);
nor U11713 (N_11713,N_6288,N_8259);
nand U11714 (N_11714,N_6541,N_6945);
nor U11715 (N_11715,N_8574,N_8429);
nand U11716 (N_11716,N_7622,N_8246);
and U11717 (N_11717,N_8313,N_7509);
or U11718 (N_11718,N_6252,N_7687);
nor U11719 (N_11719,N_8759,N_8380);
nor U11720 (N_11720,N_8567,N_7950);
nor U11721 (N_11721,N_8662,N_6153);
or U11722 (N_11722,N_6479,N_8933);
xor U11723 (N_11723,N_7642,N_6280);
nor U11724 (N_11724,N_6430,N_6964);
nor U11725 (N_11725,N_8967,N_8903);
or U11726 (N_11726,N_6044,N_8679);
xor U11727 (N_11727,N_7094,N_8504);
or U11728 (N_11728,N_7636,N_7345);
nand U11729 (N_11729,N_6180,N_7901);
and U11730 (N_11730,N_6683,N_7385);
and U11731 (N_11731,N_6028,N_7520);
and U11732 (N_11732,N_8272,N_7672);
xnor U11733 (N_11733,N_8496,N_7472);
xnor U11734 (N_11734,N_7695,N_7503);
nand U11735 (N_11735,N_7926,N_8414);
and U11736 (N_11736,N_7625,N_8187);
nor U11737 (N_11737,N_8866,N_6282);
and U11738 (N_11738,N_8780,N_7375);
or U11739 (N_11739,N_6328,N_7386);
and U11740 (N_11740,N_6999,N_8612);
and U11741 (N_11741,N_6893,N_6794);
nand U11742 (N_11742,N_8091,N_6569);
and U11743 (N_11743,N_7664,N_8418);
nor U11744 (N_11744,N_6826,N_8563);
or U11745 (N_11745,N_6770,N_7860);
and U11746 (N_11746,N_7871,N_8505);
nor U11747 (N_11747,N_6287,N_8352);
or U11748 (N_11748,N_6038,N_6827);
nand U11749 (N_11749,N_8704,N_7091);
and U11750 (N_11750,N_8708,N_8965);
or U11751 (N_11751,N_8889,N_7582);
nand U11752 (N_11752,N_7269,N_7997);
nand U11753 (N_11753,N_6985,N_7906);
nand U11754 (N_11754,N_8215,N_7090);
and U11755 (N_11755,N_6071,N_7570);
or U11756 (N_11756,N_6150,N_6586);
nand U11757 (N_11757,N_7601,N_6376);
and U11758 (N_11758,N_6044,N_6834);
nand U11759 (N_11759,N_6110,N_7446);
and U11760 (N_11760,N_7371,N_8347);
xnor U11761 (N_11761,N_8496,N_8977);
and U11762 (N_11762,N_6019,N_8462);
nor U11763 (N_11763,N_7652,N_8879);
nor U11764 (N_11764,N_8202,N_8976);
nand U11765 (N_11765,N_6795,N_8068);
nand U11766 (N_11766,N_8080,N_8266);
nand U11767 (N_11767,N_7947,N_6072);
nor U11768 (N_11768,N_8052,N_6665);
or U11769 (N_11769,N_6424,N_6962);
and U11770 (N_11770,N_7305,N_8687);
nor U11771 (N_11771,N_8973,N_8399);
xnor U11772 (N_11772,N_7268,N_8681);
or U11773 (N_11773,N_8088,N_6296);
nand U11774 (N_11774,N_7531,N_7156);
and U11775 (N_11775,N_6232,N_8486);
and U11776 (N_11776,N_6672,N_8320);
nor U11777 (N_11777,N_6085,N_7462);
and U11778 (N_11778,N_6017,N_8861);
and U11779 (N_11779,N_6303,N_6748);
and U11780 (N_11780,N_8551,N_6173);
nand U11781 (N_11781,N_6841,N_7148);
nand U11782 (N_11782,N_6020,N_7861);
and U11783 (N_11783,N_6756,N_7198);
nor U11784 (N_11784,N_8990,N_7912);
nand U11785 (N_11785,N_7780,N_7319);
nand U11786 (N_11786,N_7845,N_7962);
or U11787 (N_11787,N_6720,N_8536);
nand U11788 (N_11788,N_8161,N_8094);
nand U11789 (N_11789,N_7629,N_8237);
nor U11790 (N_11790,N_6159,N_6161);
nand U11791 (N_11791,N_8596,N_6904);
nand U11792 (N_11792,N_7175,N_7801);
nand U11793 (N_11793,N_7632,N_6329);
and U11794 (N_11794,N_6527,N_6496);
xnor U11795 (N_11795,N_8309,N_8026);
or U11796 (N_11796,N_8296,N_6288);
nand U11797 (N_11797,N_8377,N_6516);
nand U11798 (N_11798,N_8917,N_8853);
nor U11799 (N_11799,N_6039,N_8776);
nand U11800 (N_11800,N_7348,N_7111);
xnor U11801 (N_11801,N_8077,N_7326);
or U11802 (N_11802,N_8589,N_7192);
nand U11803 (N_11803,N_7277,N_7677);
nand U11804 (N_11804,N_8830,N_6736);
nor U11805 (N_11805,N_8482,N_7158);
nand U11806 (N_11806,N_7336,N_6559);
or U11807 (N_11807,N_6327,N_8018);
nor U11808 (N_11808,N_6037,N_8770);
xor U11809 (N_11809,N_6105,N_8958);
and U11810 (N_11810,N_6815,N_6119);
or U11811 (N_11811,N_6931,N_6374);
and U11812 (N_11812,N_7579,N_7437);
nor U11813 (N_11813,N_8975,N_7494);
and U11814 (N_11814,N_7089,N_7498);
nor U11815 (N_11815,N_7994,N_6789);
or U11816 (N_11816,N_6126,N_6557);
or U11817 (N_11817,N_7769,N_6417);
or U11818 (N_11818,N_8265,N_7418);
nor U11819 (N_11819,N_8599,N_8880);
nand U11820 (N_11820,N_6586,N_8137);
and U11821 (N_11821,N_7490,N_6702);
nor U11822 (N_11822,N_6141,N_7049);
nor U11823 (N_11823,N_7258,N_7938);
xnor U11824 (N_11824,N_8218,N_6581);
nor U11825 (N_11825,N_8581,N_6176);
xnor U11826 (N_11826,N_6334,N_8928);
nor U11827 (N_11827,N_6712,N_8910);
nand U11828 (N_11828,N_7101,N_7638);
nor U11829 (N_11829,N_7903,N_6084);
and U11830 (N_11830,N_8650,N_7432);
nor U11831 (N_11831,N_6334,N_6135);
or U11832 (N_11832,N_6298,N_6032);
or U11833 (N_11833,N_8889,N_7091);
nor U11834 (N_11834,N_8933,N_7952);
or U11835 (N_11835,N_6768,N_6912);
nor U11836 (N_11836,N_8547,N_7769);
or U11837 (N_11837,N_6561,N_8758);
and U11838 (N_11838,N_8216,N_7980);
and U11839 (N_11839,N_7688,N_7346);
nand U11840 (N_11840,N_8900,N_6497);
nor U11841 (N_11841,N_6716,N_8542);
nor U11842 (N_11842,N_7366,N_8398);
or U11843 (N_11843,N_7151,N_7340);
and U11844 (N_11844,N_6431,N_7517);
or U11845 (N_11845,N_7950,N_6183);
nor U11846 (N_11846,N_7363,N_6839);
or U11847 (N_11847,N_7302,N_7100);
nor U11848 (N_11848,N_7869,N_7822);
nor U11849 (N_11849,N_8790,N_7813);
xor U11850 (N_11850,N_8473,N_7591);
nand U11851 (N_11851,N_8303,N_7945);
and U11852 (N_11852,N_7020,N_7168);
nand U11853 (N_11853,N_7346,N_7134);
and U11854 (N_11854,N_7374,N_8308);
nor U11855 (N_11855,N_8787,N_6572);
and U11856 (N_11856,N_6834,N_8354);
nand U11857 (N_11857,N_6896,N_6397);
xnor U11858 (N_11858,N_8048,N_7415);
nand U11859 (N_11859,N_8914,N_8417);
or U11860 (N_11860,N_7970,N_7449);
and U11861 (N_11861,N_7421,N_7107);
nand U11862 (N_11862,N_8604,N_7511);
nand U11863 (N_11863,N_7832,N_6919);
nor U11864 (N_11864,N_6552,N_7433);
nand U11865 (N_11865,N_7038,N_6068);
or U11866 (N_11866,N_6838,N_8466);
or U11867 (N_11867,N_7059,N_6457);
nor U11868 (N_11868,N_8997,N_6596);
nor U11869 (N_11869,N_7897,N_6638);
or U11870 (N_11870,N_8045,N_8321);
nor U11871 (N_11871,N_7007,N_8884);
nand U11872 (N_11872,N_6448,N_6854);
xnor U11873 (N_11873,N_6012,N_6411);
and U11874 (N_11874,N_8069,N_6789);
and U11875 (N_11875,N_7055,N_8751);
nand U11876 (N_11876,N_8230,N_7689);
and U11877 (N_11877,N_6069,N_8294);
nor U11878 (N_11878,N_8150,N_7919);
or U11879 (N_11879,N_6286,N_8268);
xnor U11880 (N_11880,N_8550,N_8184);
or U11881 (N_11881,N_6495,N_6301);
xnor U11882 (N_11882,N_6173,N_7004);
and U11883 (N_11883,N_6808,N_6033);
nand U11884 (N_11884,N_8007,N_6002);
nor U11885 (N_11885,N_6163,N_6017);
or U11886 (N_11886,N_6698,N_8953);
and U11887 (N_11887,N_8012,N_7486);
or U11888 (N_11888,N_6600,N_8029);
nor U11889 (N_11889,N_6117,N_6882);
xor U11890 (N_11890,N_7833,N_8860);
nand U11891 (N_11891,N_7257,N_6177);
and U11892 (N_11892,N_6427,N_6158);
nor U11893 (N_11893,N_7937,N_6807);
or U11894 (N_11894,N_8359,N_6133);
or U11895 (N_11895,N_7327,N_7020);
nand U11896 (N_11896,N_8300,N_7071);
nor U11897 (N_11897,N_7752,N_6150);
nand U11898 (N_11898,N_8870,N_6462);
and U11899 (N_11899,N_8972,N_8587);
nand U11900 (N_11900,N_8422,N_8346);
nor U11901 (N_11901,N_6631,N_6519);
xnor U11902 (N_11902,N_6486,N_8844);
or U11903 (N_11903,N_7551,N_7185);
and U11904 (N_11904,N_7954,N_8172);
nand U11905 (N_11905,N_8475,N_7211);
or U11906 (N_11906,N_7252,N_8499);
or U11907 (N_11907,N_8117,N_8508);
nor U11908 (N_11908,N_7915,N_7213);
or U11909 (N_11909,N_8911,N_8750);
xnor U11910 (N_11910,N_7374,N_6232);
nand U11911 (N_11911,N_6004,N_7865);
or U11912 (N_11912,N_6664,N_6343);
and U11913 (N_11913,N_6112,N_6055);
nand U11914 (N_11914,N_7207,N_6580);
and U11915 (N_11915,N_6744,N_7897);
nor U11916 (N_11916,N_7688,N_7786);
nand U11917 (N_11917,N_8284,N_7225);
nor U11918 (N_11918,N_8674,N_7668);
or U11919 (N_11919,N_6035,N_6923);
nor U11920 (N_11920,N_6966,N_6495);
nor U11921 (N_11921,N_8438,N_8639);
or U11922 (N_11922,N_7470,N_7052);
nor U11923 (N_11923,N_6948,N_8140);
or U11924 (N_11924,N_6480,N_6554);
or U11925 (N_11925,N_6436,N_8010);
nand U11926 (N_11926,N_6071,N_7991);
xnor U11927 (N_11927,N_7322,N_6115);
nand U11928 (N_11928,N_7416,N_7046);
and U11929 (N_11929,N_7016,N_7537);
nor U11930 (N_11930,N_6270,N_7288);
and U11931 (N_11931,N_8117,N_8045);
nand U11932 (N_11932,N_6424,N_8709);
xnor U11933 (N_11933,N_7375,N_8308);
or U11934 (N_11934,N_6017,N_7039);
nor U11935 (N_11935,N_7679,N_6333);
or U11936 (N_11936,N_7334,N_8035);
or U11937 (N_11937,N_7071,N_7229);
nand U11938 (N_11938,N_7398,N_8440);
nor U11939 (N_11939,N_7351,N_7740);
nand U11940 (N_11940,N_8204,N_7476);
or U11941 (N_11941,N_8827,N_8803);
nor U11942 (N_11942,N_8116,N_8935);
or U11943 (N_11943,N_8866,N_6526);
xor U11944 (N_11944,N_6685,N_7439);
and U11945 (N_11945,N_8794,N_8494);
nor U11946 (N_11946,N_7894,N_7930);
and U11947 (N_11947,N_7710,N_8994);
nor U11948 (N_11948,N_7620,N_7488);
nand U11949 (N_11949,N_8916,N_8908);
or U11950 (N_11950,N_6965,N_8321);
or U11951 (N_11951,N_6046,N_8993);
or U11952 (N_11952,N_8959,N_7341);
or U11953 (N_11953,N_6638,N_6506);
and U11954 (N_11954,N_8474,N_8731);
xor U11955 (N_11955,N_7553,N_7985);
and U11956 (N_11956,N_8245,N_7440);
nand U11957 (N_11957,N_8262,N_8291);
nand U11958 (N_11958,N_6236,N_6765);
nand U11959 (N_11959,N_6694,N_8826);
nand U11960 (N_11960,N_6124,N_8949);
nor U11961 (N_11961,N_8601,N_7806);
nand U11962 (N_11962,N_6706,N_7428);
nand U11963 (N_11963,N_6888,N_6277);
nor U11964 (N_11964,N_7524,N_8534);
xnor U11965 (N_11965,N_8251,N_8474);
nor U11966 (N_11966,N_6956,N_6560);
or U11967 (N_11967,N_7812,N_7427);
nor U11968 (N_11968,N_6214,N_6207);
or U11969 (N_11969,N_6103,N_6146);
xor U11970 (N_11970,N_6836,N_6527);
nand U11971 (N_11971,N_6835,N_7846);
or U11972 (N_11972,N_8463,N_6695);
or U11973 (N_11973,N_8756,N_6354);
and U11974 (N_11974,N_8282,N_6071);
xor U11975 (N_11975,N_7522,N_7673);
nand U11976 (N_11976,N_8635,N_6932);
xor U11977 (N_11977,N_8725,N_8230);
and U11978 (N_11978,N_6860,N_7816);
and U11979 (N_11979,N_7839,N_6880);
nand U11980 (N_11980,N_6568,N_8665);
or U11981 (N_11981,N_6119,N_8187);
and U11982 (N_11982,N_8413,N_8715);
or U11983 (N_11983,N_7559,N_7925);
nand U11984 (N_11984,N_8429,N_7676);
or U11985 (N_11985,N_7557,N_8744);
nor U11986 (N_11986,N_6265,N_7716);
and U11987 (N_11987,N_6561,N_8220);
and U11988 (N_11988,N_7201,N_6547);
xnor U11989 (N_11989,N_7139,N_6476);
nor U11990 (N_11990,N_7514,N_6351);
xor U11991 (N_11991,N_7793,N_6885);
or U11992 (N_11992,N_8207,N_6561);
or U11993 (N_11993,N_7505,N_7904);
nand U11994 (N_11994,N_6299,N_7583);
nand U11995 (N_11995,N_7759,N_7028);
nand U11996 (N_11996,N_6165,N_8957);
and U11997 (N_11997,N_7637,N_8417);
and U11998 (N_11998,N_7024,N_6516);
nor U11999 (N_11999,N_6042,N_6171);
or U12000 (N_12000,N_10747,N_9134);
and U12001 (N_12001,N_11827,N_9703);
nor U12002 (N_12002,N_10587,N_10285);
nor U12003 (N_12003,N_11400,N_10194);
and U12004 (N_12004,N_9082,N_10143);
and U12005 (N_12005,N_11088,N_11715);
nor U12006 (N_12006,N_9810,N_10419);
or U12007 (N_12007,N_11387,N_9272);
nor U12008 (N_12008,N_10907,N_11897);
or U12009 (N_12009,N_10482,N_10139);
or U12010 (N_12010,N_11368,N_9233);
or U12011 (N_12011,N_11029,N_11484);
nor U12012 (N_12012,N_11834,N_10961);
nand U12013 (N_12013,N_11024,N_10734);
nand U12014 (N_12014,N_9452,N_9959);
and U12015 (N_12015,N_9459,N_10763);
xor U12016 (N_12016,N_11016,N_10371);
nor U12017 (N_12017,N_10556,N_9508);
nand U12018 (N_12018,N_9294,N_10025);
and U12019 (N_12019,N_10436,N_11052);
or U12020 (N_12020,N_11039,N_11151);
and U12021 (N_12021,N_11091,N_10665);
nand U12022 (N_12022,N_10233,N_11251);
or U12023 (N_12023,N_11272,N_9185);
nor U12024 (N_12024,N_11855,N_11623);
or U12025 (N_12025,N_10700,N_10687);
or U12026 (N_12026,N_11448,N_11796);
and U12027 (N_12027,N_9364,N_9660);
nor U12028 (N_12028,N_9505,N_11301);
xnor U12029 (N_12029,N_10093,N_11226);
nor U12030 (N_12030,N_10924,N_10465);
nor U12031 (N_12031,N_11450,N_11722);
nand U12032 (N_12032,N_9168,N_10495);
or U12033 (N_12033,N_11338,N_11010);
and U12034 (N_12034,N_9483,N_10534);
or U12035 (N_12035,N_9126,N_11859);
or U12036 (N_12036,N_9656,N_11232);
and U12037 (N_12037,N_9326,N_10200);
xor U12038 (N_12038,N_9414,N_9993);
nor U12039 (N_12039,N_9994,N_11688);
and U12040 (N_12040,N_11723,N_10420);
nor U12041 (N_12041,N_10794,N_9178);
and U12042 (N_12042,N_11517,N_11981);
nand U12043 (N_12043,N_9276,N_10122);
or U12044 (N_12044,N_10856,N_11528);
nor U12045 (N_12045,N_10211,N_10305);
or U12046 (N_12046,N_11491,N_11324);
or U12047 (N_12047,N_9963,N_10859);
nor U12048 (N_12048,N_10248,N_11069);
nor U12049 (N_12049,N_10038,N_10485);
nor U12050 (N_12050,N_11611,N_9740);
nor U12051 (N_12051,N_11483,N_11989);
and U12052 (N_12052,N_9197,N_10456);
nand U12053 (N_12053,N_9847,N_10113);
nor U12054 (N_12054,N_9407,N_10952);
nor U12055 (N_12055,N_9028,N_9282);
or U12056 (N_12056,N_9211,N_10701);
nand U12057 (N_12057,N_11181,N_10380);
or U12058 (N_12058,N_11939,N_10271);
nand U12059 (N_12059,N_11873,N_10294);
nor U12060 (N_12060,N_9779,N_11988);
nor U12061 (N_12061,N_11093,N_10350);
or U12062 (N_12062,N_9650,N_11830);
xnor U12063 (N_12063,N_11804,N_9658);
and U12064 (N_12064,N_10065,N_9125);
and U12065 (N_12065,N_10150,N_11601);
nand U12066 (N_12066,N_11529,N_9796);
nand U12067 (N_12067,N_9066,N_11319);
xnor U12068 (N_12068,N_9752,N_9540);
or U12069 (N_12069,N_11706,N_10207);
nor U12070 (N_12070,N_11413,N_11256);
nand U12071 (N_12071,N_10489,N_11568);
or U12072 (N_12072,N_9306,N_10652);
nor U12073 (N_12073,N_9422,N_9413);
nor U12074 (N_12074,N_11695,N_10133);
nand U12075 (N_12075,N_9045,N_11747);
or U12076 (N_12076,N_11173,N_11027);
nor U12077 (N_12077,N_11655,N_11705);
nand U12078 (N_12078,N_10120,N_9893);
nor U12079 (N_12079,N_10850,N_10676);
and U12080 (N_12080,N_10240,N_9635);
nand U12081 (N_12081,N_9990,N_10932);
xor U12082 (N_12082,N_11519,N_10826);
or U12083 (N_12083,N_11671,N_11214);
or U12084 (N_12084,N_9627,N_10068);
nand U12085 (N_12085,N_10016,N_10135);
and U12086 (N_12086,N_11328,N_10315);
nand U12087 (N_12087,N_11584,N_10396);
or U12088 (N_12088,N_9983,N_9536);
nand U12089 (N_12089,N_11128,N_9002);
or U12090 (N_12090,N_9149,N_10881);
nor U12091 (N_12091,N_11750,N_11917);
nor U12092 (N_12092,N_9463,N_11878);
and U12093 (N_12093,N_11577,N_9914);
xnor U12094 (N_12094,N_11546,N_10384);
xnor U12095 (N_12095,N_11635,N_11185);
xor U12096 (N_12096,N_10158,N_11990);
and U12097 (N_12097,N_10639,N_11773);
nor U12098 (N_12098,N_11107,N_9746);
and U12099 (N_12099,N_11877,N_10114);
nand U12100 (N_12100,N_11221,N_10003);
nand U12101 (N_12101,N_10594,N_10748);
xnor U12102 (N_12102,N_10376,N_11753);
nor U12103 (N_12103,N_11087,N_10653);
nand U12104 (N_12104,N_11143,N_9894);
xnor U12105 (N_12105,N_11759,N_9203);
xnor U12106 (N_12106,N_9794,N_11157);
nor U12107 (N_12107,N_11680,N_9049);
xnor U12108 (N_12108,N_10429,N_9039);
and U12109 (N_12109,N_10921,N_9661);
and U12110 (N_12110,N_11691,N_10867);
nand U12111 (N_12111,N_9288,N_10678);
nor U12112 (N_12112,N_9095,N_10812);
nor U12113 (N_12113,N_10742,N_10781);
nand U12114 (N_12114,N_10631,N_11478);
or U12115 (N_12115,N_9121,N_11224);
nor U12116 (N_12116,N_10744,N_11971);
nor U12117 (N_12117,N_10985,N_10664);
or U12118 (N_12118,N_10833,N_10272);
or U12119 (N_12119,N_9051,N_9652);
xor U12120 (N_12120,N_10595,N_9972);
and U12121 (N_12121,N_11071,N_10868);
nor U12122 (N_12122,N_9360,N_9885);
xor U12123 (N_12123,N_10731,N_9113);
and U12124 (N_12124,N_11238,N_11512);
or U12125 (N_12125,N_10815,N_10872);
nor U12126 (N_12126,N_11514,N_9322);
nor U12127 (N_12127,N_9227,N_9410);
or U12128 (N_12128,N_9996,N_9030);
nor U12129 (N_12129,N_11973,N_9176);
nand U12130 (N_12130,N_10521,N_11240);
and U12131 (N_12131,N_9576,N_10142);
or U12132 (N_12132,N_11282,N_10131);
nand U12133 (N_12133,N_10788,N_10360);
or U12134 (N_12134,N_10566,N_10501);
or U12135 (N_12135,N_10963,N_10909);
nor U12136 (N_12136,N_10746,N_10453);
xnor U12137 (N_12137,N_9995,N_11381);
nand U12138 (N_12138,N_9783,N_9940);
or U12139 (N_12139,N_10450,N_9547);
xor U12140 (N_12140,N_10182,N_9036);
or U12141 (N_12141,N_10879,N_9135);
or U12142 (N_12142,N_9630,N_9755);
and U12143 (N_12143,N_11094,N_10259);
xnor U12144 (N_12144,N_9150,N_11443);
or U12145 (N_12145,N_11742,N_10757);
nand U12146 (N_12146,N_9938,N_10344);
and U12147 (N_12147,N_11525,N_9921);
nand U12148 (N_12148,N_10713,N_11649);
nand U12149 (N_12149,N_10972,N_9965);
or U12150 (N_12150,N_11497,N_9878);
and U12151 (N_12151,N_9849,N_11408);
nor U12152 (N_12152,N_10488,N_11234);
nand U12153 (N_12153,N_10497,N_10264);
nor U12154 (N_12154,N_11672,N_11465);
nand U12155 (N_12155,N_10729,N_11521);
and U12156 (N_12156,N_11875,N_9432);
nor U12157 (N_12157,N_11829,N_9757);
or U12158 (N_12158,N_11686,N_10255);
nor U12159 (N_12159,N_10662,N_9496);
nor U12160 (N_12160,N_10507,N_11122);
nand U12161 (N_12161,N_11175,N_11144);
or U12162 (N_12162,N_11086,N_10765);
nand U12163 (N_12163,N_10999,N_10537);
and U12164 (N_12164,N_10931,N_10399);
nor U12165 (N_12165,N_11476,N_10171);
nand U12166 (N_12166,N_9420,N_10836);
xnor U12167 (N_12167,N_9817,N_9260);
xor U12168 (N_12168,N_10401,N_10353);
or U12169 (N_12169,N_10818,N_10823);
and U12170 (N_12170,N_11007,N_10159);
nor U12171 (N_12171,N_10839,N_10252);
nand U12172 (N_12172,N_9874,N_10598);
and U12173 (N_12173,N_9477,N_9475);
nand U12174 (N_12174,N_9533,N_9926);
nor U12175 (N_12175,N_9469,N_11113);
nor U12176 (N_12176,N_10899,N_9927);
nand U12177 (N_12177,N_9281,N_11660);
or U12178 (N_12178,N_10659,N_9816);
and U12179 (N_12179,N_9307,N_11762);
and U12180 (N_12180,N_10636,N_11719);
or U12181 (N_12181,N_11161,N_10571);
or U12182 (N_12182,N_9587,N_10220);
nand U12183 (N_12183,N_10953,N_10364);
and U12184 (N_12184,N_10692,N_11460);
or U12185 (N_12185,N_10716,N_11906);
and U12186 (N_12186,N_10983,N_10679);
or U12187 (N_12187,N_9860,N_10616);
and U12188 (N_12188,N_11812,N_10984);
nor U12189 (N_12189,N_11409,N_9657);
and U12190 (N_12190,N_9270,N_10004);
nor U12191 (N_12191,N_10882,N_11970);
and U12192 (N_12192,N_10434,N_11624);
nand U12193 (N_12193,N_9200,N_11800);
and U12194 (N_12194,N_9356,N_9648);
nand U12195 (N_12195,N_10814,N_10052);
or U12196 (N_12196,N_11698,N_9062);
nand U12197 (N_12197,N_11178,N_11535);
and U12198 (N_12198,N_9730,N_11882);
nor U12199 (N_12199,N_10469,N_11211);
nor U12200 (N_12200,N_10613,N_10413);
or U12201 (N_12201,N_10722,N_11427);
nand U12202 (N_12202,N_11269,N_10261);
xnor U12203 (N_12203,N_11236,N_10253);
or U12204 (N_12204,N_10714,N_11560);
and U12205 (N_12205,N_11890,N_9212);
xnor U12206 (N_12206,N_9058,N_11502);
or U12207 (N_12207,N_11229,N_9727);
nand U12208 (N_12208,N_10050,N_10109);
nor U12209 (N_12209,N_9237,N_10042);
and U12210 (N_12210,N_9418,N_9397);
and U12211 (N_12211,N_9968,N_9786);
nor U12212 (N_12212,N_11543,N_11960);
nand U12213 (N_12213,N_10449,N_9844);
nand U12214 (N_12214,N_11189,N_11956);
or U12215 (N_12215,N_11083,N_9218);
and U12216 (N_12216,N_11752,N_9962);
and U12217 (N_12217,N_9341,N_10110);
or U12218 (N_12218,N_11850,N_10715);
nor U12219 (N_12219,N_9831,N_10494);
xor U12220 (N_12220,N_10165,N_11940);
and U12221 (N_12221,N_10599,N_10368);
nor U12222 (N_12222,N_10809,N_11851);
and U12223 (N_12223,N_10090,N_11239);
and U12224 (N_12224,N_11202,N_10876);
nor U12225 (N_12225,N_11455,N_10394);
nand U12226 (N_12226,N_11761,N_9585);
and U12227 (N_12227,N_9298,N_9381);
nor U12228 (N_12228,N_11740,N_9782);
and U12229 (N_12229,N_10550,N_10915);
nand U12230 (N_12230,N_9772,N_10979);
nand U12231 (N_12231,N_9229,N_9456);
or U12232 (N_12232,N_10130,N_9009);
nand U12233 (N_12233,N_11223,N_9239);
and U12234 (N_12234,N_9524,N_9527);
nor U12235 (N_12235,N_11072,N_10440);
or U12236 (N_12236,N_11000,N_10307);
and U12237 (N_12237,N_10655,N_10926);
or U12238 (N_12238,N_9194,N_11669);
or U12239 (N_12239,N_9479,N_9908);
nand U12240 (N_12240,N_9526,N_10414);
nand U12241 (N_12241,N_10783,N_9900);
nor U12242 (N_12242,N_9099,N_9287);
or U12243 (N_12243,N_9154,N_9956);
xor U12244 (N_12244,N_9924,N_10922);
nor U12245 (N_12245,N_9266,N_11291);
nand U12246 (N_12246,N_9631,N_11146);
nor U12247 (N_12247,N_10835,N_10381);
nor U12248 (N_12248,N_10056,N_11821);
or U12249 (N_12249,N_10483,N_11541);
or U12250 (N_12250,N_9224,N_11275);
nor U12251 (N_12251,N_11588,N_10905);
and U12252 (N_12252,N_10508,N_10768);
and U12253 (N_12253,N_10925,N_11627);
nand U12254 (N_12254,N_9106,N_11515);
or U12255 (N_12255,N_11365,N_11857);
xor U12256 (N_12256,N_11997,N_10441);
and U12257 (N_12257,N_10906,N_10303);
xor U12258 (N_12258,N_10333,N_9254);
or U12259 (N_12259,N_9726,N_9430);
or U12260 (N_12260,N_10164,N_9735);
and U12261 (N_12261,N_10709,N_11589);
nor U12262 (N_12262,N_10018,N_11808);
and U12263 (N_12263,N_9166,N_9445);
and U12264 (N_12264,N_10597,N_11955);
and U12265 (N_12265,N_9883,N_10178);
nand U12266 (N_12266,N_10893,N_9992);
or U12267 (N_12267,N_9472,N_9593);
nor U12268 (N_12268,N_10124,N_9554);
and U12269 (N_12269,N_9471,N_11192);
nor U12270 (N_12270,N_10204,N_10877);
nand U12271 (N_12271,N_9674,N_11929);
or U12272 (N_12272,N_11789,N_10047);
or U12273 (N_12273,N_11662,N_10367);
xor U12274 (N_12274,N_9513,N_9791);
and U12275 (N_12275,N_9283,N_9812);
nand U12276 (N_12276,N_9174,N_11676);
xor U12277 (N_12277,N_10035,N_9119);
nor U12278 (N_12278,N_9171,N_11074);
and U12279 (N_12279,N_10919,N_10094);
and U12280 (N_12280,N_10752,N_9615);
or U12281 (N_12281,N_11505,N_9493);
nor U12282 (N_12282,N_11458,N_11042);
and U12283 (N_12283,N_10184,N_11243);
nand U12284 (N_12284,N_11966,N_10431);
nor U12285 (N_12285,N_9638,N_10321);
nor U12286 (N_12286,N_10417,N_9415);
and U12287 (N_12287,N_11123,N_10189);
nand U12288 (N_12288,N_11165,N_10874);
or U12289 (N_12289,N_9611,N_9309);
or U12290 (N_12290,N_9987,N_9625);
nand U12291 (N_12291,N_9152,N_11060);
or U12292 (N_12292,N_10504,N_11526);
or U12293 (N_12293,N_9047,N_10002);
and U12294 (N_12294,N_9750,N_9440);
xor U12295 (N_12295,N_11618,N_9424);
nor U12296 (N_12296,N_10945,N_9167);
or U12297 (N_12297,N_9699,N_11656);
nand U12298 (N_12298,N_9512,N_11756);
or U12299 (N_12299,N_9428,N_9075);
and U12300 (N_12300,N_11090,N_9614);
or U12301 (N_12301,N_10470,N_10481);
xor U12302 (N_12302,N_10523,N_9000);
and U12303 (N_12303,N_10478,N_11566);
or U12304 (N_12304,N_11297,N_11119);
xor U12305 (N_12305,N_10551,N_11145);
or U12306 (N_12306,N_11023,N_10445);
and U12307 (N_12307,N_9115,N_9623);
and U12308 (N_12308,N_9856,N_9158);
xnor U12309 (N_12309,N_11089,N_9186);
nand U12310 (N_12310,N_11798,N_10549);
nand U12311 (N_12311,N_10741,N_11444);
nand U12312 (N_12312,N_11516,N_10954);
or U12313 (N_12313,N_11567,N_10548);
and U12314 (N_12314,N_9853,N_11166);
nand U12315 (N_12315,N_10432,N_10437);
and U12316 (N_12316,N_9142,N_9426);
and U12317 (N_12317,N_11564,N_10672);
nand U12318 (N_12318,N_10279,N_9988);
or U12319 (N_12319,N_9519,N_10357);
or U12320 (N_12320,N_9712,N_10438);
nand U12321 (N_12321,N_9235,N_11429);
nor U12322 (N_12322,N_9767,N_11210);
nor U12323 (N_12323,N_11580,N_11558);
nand U12324 (N_12324,N_10820,N_10095);
nor U12325 (N_12325,N_11975,N_9120);
nand U12326 (N_12326,N_10338,N_10822);
and U12327 (N_12327,N_9013,N_9668);
xnor U12328 (N_12328,N_11542,N_9435);
or U12329 (N_12329,N_10258,N_10174);
and U12330 (N_12330,N_10006,N_10973);
and U12331 (N_12331,N_11823,N_11280);
nor U12332 (N_12332,N_10318,N_11325);
nand U12333 (N_12333,N_11925,N_10694);
nor U12334 (N_12334,N_10009,N_11341);
or U12335 (N_12335,N_10282,N_10039);
nand U12336 (N_12336,N_10570,N_9653);
and U12337 (N_12337,N_9466,N_9534);
nor U12338 (N_12338,N_10074,N_10810);
or U12339 (N_12339,N_9012,N_11292);
or U12340 (N_12340,N_11401,N_11288);
nor U12341 (N_12341,N_11704,N_11776);
nor U12342 (N_12342,N_9811,N_9494);
and U12343 (N_12343,N_11106,N_9843);
nand U12344 (N_12344,N_9226,N_10971);
or U12345 (N_12345,N_9347,N_10317);
or U12346 (N_12346,N_10468,N_10390);
nor U12347 (N_12347,N_9634,N_10575);
xor U12348 (N_12348,N_11844,N_9562);
and U12349 (N_12349,N_9080,N_11035);
and U12350 (N_12350,N_11816,N_11435);
or U12351 (N_12351,N_11734,N_10198);
or U12352 (N_12352,N_10785,N_9497);
nand U12353 (N_12353,N_10319,N_11911);
and U12354 (N_12354,N_9495,N_11574);
and U12355 (N_12355,N_11331,N_11352);
and U12356 (N_12356,N_9128,N_11417);
nand U12357 (N_12357,N_9588,N_9838);
xnor U12358 (N_12358,N_10132,N_10447);
or U12359 (N_12359,N_9041,N_11944);
and U12360 (N_12360,N_11664,N_9136);
nor U12361 (N_12361,N_10354,N_11510);
and U12362 (N_12362,N_9510,N_9912);
or U12363 (N_12363,N_10270,N_11570);
nor U12364 (N_12364,N_11279,N_9403);
nand U12365 (N_12365,N_11498,N_11138);
nand U12366 (N_12366,N_10502,N_11538);
nor U12367 (N_12367,N_10772,N_10855);
xnor U12368 (N_12368,N_11885,N_9217);
nand U12369 (N_12369,N_10402,N_9243);
nand U12370 (N_12370,N_11907,N_11986);
and U12371 (N_12371,N_9258,N_11037);
or U12372 (N_12372,N_9780,N_10256);
or U12373 (N_12373,N_11233,N_10103);
nand U12374 (N_12374,N_9798,N_11696);
nor U12375 (N_12375,N_9457,N_10476);
and U12376 (N_12376,N_11025,N_10115);
and U12377 (N_12377,N_11692,N_10439);
or U12378 (N_12378,N_9346,N_11569);
and U12379 (N_12379,N_9803,N_11363);
or U12380 (N_12380,N_9261,N_10011);
or U12381 (N_12381,N_10176,N_11342);
or U12382 (N_12382,N_11622,N_10965);
nand U12383 (N_12383,N_11822,N_10335);
xnor U12384 (N_12384,N_9771,N_9970);
or U12385 (N_12385,N_11654,N_10552);
nand U12386 (N_12386,N_10300,N_9643);
and U12387 (N_12387,N_9967,N_9369);
nand U12388 (N_12388,N_11082,N_9131);
nor U12389 (N_12389,N_11732,N_10167);
nand U12390 (N_12390,N_11109,N_10591);
xor U12391 (N_12391,N_11390,N_10392);
xor U12392 (N_12392,N_11343,N_9586);
and U12393 (N_12393,N_9589,N_10276);
nand U12394 (N_12394,N_11679,N_11246);
nor U12395 (N_12395,N_11076,N_10627);
or U12396 (N_12396,N_9873,N_9455);
and U12397 (N_12397,N_10843,N_11041);
nand U12398 (N_12398,N_9303,N_10179);
xor U12399 (N_12399,N_10473,N_10228);
and U12400 (N_12400,N_10711,N_11969);
nand U12401 (N_12401,N_11818,N_11063);
and U12402 (N_12402,N_9324,N_11994);
nand U12403 (N_12403,N_10407,N_10980);
and U12404 (N_12404,N_9603,N_10683);
nand U12405 (N_12405,N_9690,N_9597);
nand U12406 (N_12406,N_11923,N_10491);
and U12407 (N_12407,N_11043,N_11315);
nor U12408 (N_12408,N_9180,N_11265);
nand U12409 (N_12409,N_11631,N_10190);
or U12410 (N_12410,N_10202,N_9758);
and U12411 (N_12411,N_10331,N_11394);
or U12412 (N_12412,N_11281,N_11849);
xor U12413 (N_12413,N_10986,N_9724);
and U12414 (N_12414,N_9248,N_11118);
or U12415 (N_12415,N_11922,N_10212);
nor U12416 (N_12416,N_9351,N_9087);
nand U12417 (N_12417,N_11194,N_11530);
or U12418 (N_12418,N_11702,N_11914);
or U12419 (N_12419,N_9419,N_10543);
nand U12420 (N_12420,N_9552,N_10448);
or U12421 (N_12421,N_10624,N_9948);
and U12422 (N_12422,N_11196,N_9467);
or U12423 (N_12423,N_10000,N_9899);
xor U12424 (N_12424,N_10728,N_9026);
nor U12425 (N_12425,N_9901,N_11021);
nor U12426 (N_12426,N_10119,N_11426);
nand U12427 (N_12427,N_9887,N_11926);
nand U12428 (N_12428,N_9319,N_9292);
nor U12429 (N_12429,N_10807,N_9209);
nand U12430 (N_12430,N_11299,N_9001);
nor U12431 (N_12431,N_11501,N_9144);
nand U12432 (N_12432,N_11121,N_10435);
or U12433 (N_12433,N_9183,N_9442);
and U12434 (N_12434,N_10037,N_9008);
xor U12435 (N_12435,N_9913,N_11078);
or U12436 (N_12436,N_10584,N_9362);
nand U12437 (N_12437,N_11665,N_10254);
and U12438 (N_12438,N_9368,N_9295);
or U12439 (N_12439,N_10528,N_9023);
xor U12440 (N_12440,N_9482,N_9837);
nor U12441 (N_12441,N_11054,N_9925);
nand U12442 (N_12442,N_9792,N_9569);
or U12443 (N_12443,N_11428,N_11746);
nand U12444 (N_12444,N_10960,N_10887);
and U12445 (N_12445,N_9101,N_11227);
or U12446 (N_12446,N_10216,N_11242);
nand U12447 (N_12447,N_11967,N_9964);
or U12448 (N_12448,N_10625,N_9808);
and U12449 (N_12449,N_11262,N_10296);
nor U12450 (N_12450,N_9622,N_10128);
nand U12451 (N_12451,N_10739,N_11527);
nand U12452 (N_12452,N_10871,N_11261);
and U12453 (N_12453,N_11137,N_10975);
and U12454 (N_12454,N_10218,N_11828);
xor U12455 (N_12455,N_10588,N_9877);
nand U12456 (N_12456,N_10430,N_11894);
nand U12457 (N_12457,N_9502,N_10069);
xnor U12458 (N_12458,N_9257,N_10341);
nor U12459 (N_12459,N_10295,N_9108);
nor U12460 (N_12460,N_11638,N_10949);
nor U12461 (N_12461,N_10287,N_9377);
and U12462 (N_12462,N_10474,N_11609);
or U12463 (N_12463,N_11729,N_9891);
xor U12464 (N_12464,N_10241,N_10541);
nor U12465 (N_12465,N_9195,N_9840);
nand U12466 (N_12466,N_9775,N_10870);
nor U12467 (N_12467,N_9416,N_11718);
nand U12468 (N_12468,N_10695,N_9788);
and U12469 (N_12469,N_9943,N_11965);
or U12470 (N_12470,N_9715,N_10289);
nor U12471 (N_12471,N_9476,N_9328);
or U12472 (N_12472,N_10503,N_9365);
and U12473 (N_12473,N_11479,N_9999);
nand U12474 (N_12474,N_11913,N_11213);
nor U12475 (N_12475,N_10361,N_11938);
and U12476 (N_12476,N_9400,N_11404);
and U12477 (N_12477,N_9694,N_9641);
or U12478 (N_12478,N_10796,N_9725);
and U12479 (N_12479,N_11422,N_10185);
and U12480 (N_12480,N_11884,N_11371);
or U12481 (N_12481,N_9280,N_11389);
nor U12482 (N_12482,N_11728,N_11646);
or U12483 (N_12483,N_10416,N_11613);
nor U12484 (N_12484,N_10145,N_9939);
nor U12485 (N_12485,N_11345,N_9692);
nand U12486 (N_12486,N_9388,N_9664);
and U12487 (N_12487,N_11561,N_11678);
and U12488 (N_12488,N_10590,N_10192);
nor U12489 (N_12489,N_9517,N_9998);
or U12490 (N_12490,N_10998,N_11650);
nor U12491 (N_12491,N_9454,N_11001);
and U12492 (N_12492,N_11625,N_9175);
and U12493 (N_12493,N_11399,N_9329);
and U12494 (N_12494,N_11209,N_10735);
nor U12495 (N_12495,N_10334,N_10832);
and U12496 (N_12496,N_10828,N_9773);
or U12497 (N_12497,N_11703,N_10337);
nand U12498 (N_12498,N_9404,N_10302);
nor U12499 (N_12499,N_10446,N_11603);
or U12500 (N_12500,N_11957,N_9114);
nand U12501 (N_12501,N_10217,N_10831);
or U12502 (N_12502,N_11861,N_10671);
nor U12503 (N_12503,N_9818,N_11477);
nor U12504 (N_12504,N_9210,N_9716);
nand U12505 (N_12505,N_10857,N_10654);
and U12506 (N_12506,N_11252,N_10043);
or U12507 (N_12507,N_11405,N_10203);
and U12508 (N_12508,N_9104,N_9070);
nor U12509 (N_12509,N_10247,N_10989);
or U12510 (N_12510,N_10499,N_10916);
xnor U12511 (N_12511,N_10576,N_10804);
nor U12512 (N_12512,N_10929,N_10129);
or U12513 (N_12513,N_11807,N_11865);
or U12514 (N_12514,N_11916,N_11153);
and U12515 (N_12515,N_9153,N_11848);
nand U12516 (N_12516,N_9405,N_9359);
nor U12517 (N_12517,N_10284,N_11306);
nor U12518 (N_12518,N_10071,N_11931);
or U12519 (N_12519,N_9551,N_11220);
nand U12520 (N_12520,N_11357,N_11395);
and U12521 (N_12521,N_9704,N_11295);
nand U12522 (N_12522,N_10278,N_10177);
nor U12523 (N_12523,N_10845,N_11760);
nor U12524 (N_12524,N_10637,N_11805);
nor U12525 (N_12525,N_9285,N_11053);
xnor U12526 (N_12526,N_11263,N_10391);
nand U12527 (N_12527,N_11996,N_11819);
nor U12528 (N_12528,N_11311,N_10422);
and U12529 (N_12529,N_9697,N_9563);
and U12530 (N_12530,N_11434,N_10323);
and U12531 (N_12531,N_9645,N_9875);
nand U12532 (N_12532,N_9685,N_11470);
or U12533 (N_12533,N_9279,N_9762);
or U12534 (N_12534,N_10606,N_9338);
xor U12535 (N_12535,N_10288,N_9204);
or U12536 (N_12536,N_10015,N_9275);
and U12537 (N_12537,N_9580,N_9003);
nor U12538 (N_12538,N_10789,N_10733);
and U12539 (N_12539,N_9357,N_11933);
and U12540 (N_12540,N_10567,N_11987);
nand U12541 (N_12541,N_11847,N_9866);
nand U12542 (N_12542,N_11757,N_11572);
or U12543 (N_12543,N_9785,N_10829);
nand U12544 (N_12544,N_9907,N_9054);
and U12545 (N_12545,N_11636,N_9545);
xor U12546 (N_12546,N_10615,N_10316);
xnor U12547 (N_12547,N_11051,N_9754);
or U12548 (N_12548,N_9876,N_9184);
nand U12549 (N_12549,N_9986,N_10108);
or U12550 (N_12550,N_9515,N_11059);
and U12551 (N_12551,N_9129,N_11675);
xnor U12552 (N_12552,N_9971,N_10644);
xor U12553 (N_12553,N_11710,N_9453);
and U12554 (N_12554,N_10869,N_10538);
and U12555 (N_12555,N_11207,N_9271);
nor U12556 (N_12556,N_10097,N_9805);
nor U12557 (N_12557,N_9680,N_9091);
xor U12558 (N_12558,N_9919,N_9332);
or U12559 (N_12559,N_11190,N_9343);
or U12560 (N_12560,N_11117,N_9065);
and U12561 (N_12561,N_9507,N_9441);
nand U12562 (N_12562,N_9067,N_10620);
or U12563 (N_12563,N_10726,N_9639);
nor U12564 (N_12564,N_11049,N_11754);
or U12565 (N_12565,N_9382,N_10269);
nand U12566 (N_12566,N_9981,N_9278);
nand U12567 (N_12567,N_11290,N_10937);
nor U12568 (N_12568,N_11098,N_10487);
and U12569 (N_12569,N_10642,N_9208);
xor U12570 (N_12570,N_11788,N_9707);
and U12571 (N_12571,N_10816,N_9709);
nand U12572 (N_12572,N_10612,N_9997);
nand U12573 (N_12573,N_10904,N_11416);
or U12574 (N_12574,N_10032,N_9646);
nor U12575 (N_12575,N_11817,N_9544);
nor U12576 (N_12576,N_11846,N_9916);
nand U12577 (N_12577,N_10239,N_10260);
xnor U12578 (N_12578,N_11592,N_11633);
or U12579 (N_12579,N_10950,N_11425);
nor U12580 (N_12580,N_10425,N_10967);
and U12581 (N_12581,N_9969,N_9738);
or U12582 (N_12582,N_9706,N_11260);
nand U12583 (N_12583,N_10460,N_9826);
xnor U12584 (N_12584,N_10680,N_11046);
xnor U12585 (N_12585,N_11854,N_11508);
xnor U12586 (N_12586,N_9745,N_10824);
nor U12587 (N_12587,N_10565,N_10806);
nor U12588 (N_12588,N_10805,N_10490);
nor U12589 (N_12589,N_9465,N_9610);
or U12590 (N_12590,N_11858,N_10049);
nand U12591 (N_12591,N_9446,N_9678);
nor U12592 (N_12592,N_10498,N_9179);
xnor U12593 (N_12593,N_9743,N_11026);
nand U12594 (N_12594,N_9093,N_9068);
xor U12595 (N_12595,N_9354,N_10324);
nand U12596 (N_12596,N_9116,N_11036);
xnor U12597 (N_12597,N_10863,N_9470);
nand U12598 (N_12598,N_11255,N_10996);
and U12599 (N_12599,N_9825,N_10520);
and U12600 (N_12600,N_10140,N_9005);
nand U12601 (N_12601,N_9695,N_9124);
or U12602 (N_12602,N_10340,N_9044);
nor U12603 (N_12603,N_11370,N_10691);
nand U12604 (N_12604,N_9189,N_11713);
and U12605 (N_12605,N_11276,N_9572);
or U12606 (N_12606,N_9094,N_10935);
and U12607 (N_12607,N_9213,N_11104);
nor U12608 (N_12608,N_9460,N_9263);
and U12609 (N_12609,N_11310,N_10799);
xor U12610 (N_12610,N_10134,N_10154);
and U12611 (N_12611,N_10941,N_10411);
nor U12612 (N_12612,N_11084,N_9799);
and U12613 (N_12613,N_10210,N_10593);
or U12614 (N_12614,N_9161,N_11790);
and U12615 (N_12615,N_9096,N_11193);
nand U12616 (N_12616,N_10808,N_9409);
and U12617 (N_12617,N_10088,N_10718);
xnor U12618 (N_12618,N_10496,N_11459);
and U12619 (N_12619,N_11201,N_11253);
nand U12620 (N_12620,N_9433,N_10512);
nor U12621 (N_12621,N_9553,N_11974);
nor U12622 (N_12622,N_10974,N_9011);
and U12623 (N_12623,N_10387,N_11547);
nor U12624 (N_12624,N_10860,N_10306);
xor U12625 (N_12625,N_9579,N_11329);
or U12626 (N_12626,N_10732,N_10086);
xnor U12627 (N_12627,N_9567,N_11895);
xor U12628 (N_12628,N_9015,N_11681);
or U12629 (N_12629,N_10675,N_10619);
or U12630 (N_12630,N_9267,N_11333);
and U12631 (N_12631,N_9954,N_9334);
nand U12632 (N_12632,N_10667,N_10638);
or U12633 (N_12633,N_11383,N_10792);
or U12634 (N_12634,N_11838,N_11581);
or U12635 (N_12635,N_11103,N_9321);
and U12636 (N_12636,N_9489,N_9596);
nor U12637 (N_12637,N_11163,N_11402);
nand U12638 (N_12638,N_9118,N_11392);
and U12639 (N_12639,N_10061,N_10320);
nand U12640 (N_12640,N_9708,N_9936);
or U12641 (N_12641,N_11991,N_11831);
nor U12642 (N_12642,N_10426,N_9835);
nor U12643 (N_12643,N_11068,N_10834);
nand U12644 (N_12644,N_10981,N_11347);
nor U12645 (N_12645,N_11340,N_11839);
or U12646 (N_12646,N_11344,N_9313);
xnor U12647 (N_12647,N_10075,N_10773);
nor U12648 (N_12648,N_11441,N_11195);
or U12649 (N_12649,N_9673,N_11158);
nor U12650 (N_12650,N_11724,N_10023);
nor U12651 (N_12651,N_9766,N_9804);
and U12652 (N_12652,N_11386,N_9350);
nor U12653 (N_12653,N_9765,N_9606);
and U12654 (N_12654,N_10707,N_11741);
nor U12655 (N_12655,N_11454,N_9345);
xnor U12656 (N_12656,N_9024,N_9083);
nor U12657 (N_12657,N_11978,N_11388);
nand U12658 (N_12658,N_9702,N_10682);
or U12659 (N_12659,N_11959,N_11585);
or U12660 (N_12660,N_10685,N_10524);
or U12661 (N_12661,N_11901,N_9806);
nand U12662 (N_12662,N_10647,N_11952);
and U12663 (N_12663,N_10634,N_10775);
nor U12664 (N_12664,N_9447,N_10947);
or U12665 (N_12665,N_9599,N_9392);
nand U12666 (N_12666,N_10569,N_11135);
or U12667 (N_12667,N_11259,N_11019);
nor U12668 (N_12668,N_11167,N_10301);
nor U12669 (N_12669,N_9148,N_11350);
nand U12670 (N_12670,N_9262,N_11414);
nand U12671 (N_12671,N_11110,N_9889);
nand U12672 (N_12672,N_9284,N_10546);
or U12673 (N_12673,N_11487,N_9079);
and U12674 (N_12674,N_9531,N_10632);
nor U12675 (N_12675,N_10891,N_11912);
and U12676 (N_12676,N_11397,N_9626);
xnor U12677 (N_12677,N_11205,N_9386);
nor U12678 (N_12678,N_11531,N_11919);
and U12679 (N_12679,N_9879,N_10155);
and U12680 (N_12680,N_10712,N_9221);
and U12681 (N_12681,N_10379,N_10890);
and U12682 (N_12682,N_10553,N_11204);
nor U12683 (N_12683,N_10423,N_10215);
nor U12684 (N_12684,N_10310,N_11946);
xnor U12685 (N_12685,N_10014,N_11898);
nor U12686 (N_12686,N_10365,N_10618);
nand U12687 (N_12687,N_9187,N_9427);
nand U12688 (N_12688,N_9071,N_10268);
or U12689 (N_12689,N_10208,N_10646);
or U12690 (N_12690,N_9541,N_9686);
nor U12691 (N_12691,N_11267,N_10313);
nor U12692 (N_12692,N_11908,N_11534);
and U12693 (N_12693,N_10355,N_10670);
xor U12694 (N_12694,N_11418,N_10730);
xnor U12695 (N_12695,N_10180,N_9797);
and U12696 (N_12696,N_9696,N_10045);
or U12697 (N_12697,N_11463,N_11257);
or U12698 (N_12698,N_10697,N_9801);
xor U12699 (N_12699,N_9361,N_10755);
or U12700 (N_12700,N_10183,N_11079);
nand U12701 (N_12701,N_9549,N_10163);
or U12702 (N_12702,N_11384,N_9205);
or U12703 (N_12703,N_11300,N_10896);
and U12704 (N_12704,N_11670,N_10738);
or U12705 (N_12705,N_11159,N_10751);
nor U12706 (N_12706,N_9311,N_9402);
nor U12707 (N_12707,N_10250,N_11360);
xnor U12708 (N_12708,N_11721,N_9050);
nor U12709 (N_12709,N_9421,N_9029);
nor U12710 (N_12710,N_11769,N_10166);
or U12711 (N_12711,N_11540,N_11867);
nand U12712 (N_12712,N_10601,N_10943);
or U12713 (N_12713,N_10886,N_9575);
nor U12714 (N_12714,N_11327,N_10542);
nor U12715 (N_12715,N_11141,N_11406);
nand U12716 (N_12716,N_10914,N_9761);
nand U12717 (N_12717,N_9888,N_11148);
and U12718 (N_12718,N_10795,N_10706);
nor U12719 (N_12719,N_10514,N_11266);
or U12720 (N_12720,N_9145,N_11888);
nor U12721 (N_12721,N_10105,N_10944);
nor U12722 (N_12722,N_9201,N_11149);
nand U12723 (N_12723,N_11199,N_11640);
or U12724 (N_12724,N_10977,N_11462);
and U12725 (N_12725,N_11833,N_9398);
or U12726 (N_12726,N_9862,N_10404);
nand U12727 (N_12727,N_10293,N_11140);
nor U12728 (N_12728,N_11766,N_9865);
nor U12729 (N_12729,N_9383,N_11755);
nor U12730 (N_12730,N_9501,N_10243);
and U12731 (N_12731,N_9640,N_11881);
nor U12732 (N_12732,N_9017,N_11608);
or U12733 (N_12733,N_10892,N_10770);
nor U12734 (N_12734,N_10583,N_10767);
and U12735 (N_12735,N_9247,N_11910);
nand U12736 (N_12736,N_9112,N_9958);
or U12737 (N_12737,N_10760,N_9719);
xor U12738 (N_12738,N_10743,N_9701);
nand U12739 (N_12739,N_10092,N_10136);
nand U12740 (N_12740,N_11733,N_11774);
nand U12741 (N_12741,N_10753,N_10862);
nor U12742 (N_12742,N_9558,N_11661);
nand U12743 (N_12743,N_11915,N_9688);
nand U12744 (N_12744,N_10082,N_9842);
and U12745 (N_12745,N_9090,N_10123);
or U12746 (N_12746,N_9355,N_9560);
nand U12747 (N_12747,N_10397,N_9930);
xor U12748 (N_12748,N_9850,N_11382);
or U12749 (N_12749,N_11006,N_11250);
nand U12750 (N_12750,N_10027,N_11614);
nor U12751 (N_12751,N_11028,N_9234);
and U12752 (N_12752,N_11899,N_10920);
or U12753 (N_12753,N_9548,N_9813);
and U12754 (N_12754,N_10312,N_10299);
or U12755 (N_12755,N_10621,N_10698);
nor U12756 (N_12756,N_9301,N_10573);
nand U12757 (N_12757,N_9374,N_11632);
and U12758 (N_12758,N_11056,N_9528);
nor U12759 (N_12759,N_9820,N_11587);
nand U12760 (N_12760,N_9957,N_9034);
or U12761 (N_12761,N_11556,N_11507);
nand U12762 (N_12762,N_11576,N_9451);
and U12763 (N_12763,N_10825,N_9437);
or U12764 (N_12764,N_11375,N_9157);
or U12765 (N_12765,N_10152,N_9349);
nand U12766 (N_12766,N_10982,N_11687);
xor U12767 (N_12767,N_11235,N_11369);
and U12768 (N_12768,N_11985,N_9649);
and U12769 (N_12769,N_10611,N_11644);
xnor U12770 (N_12770,N_11593,N_11442);
and U12771 (N_12771,N_9613,N_9616);
and U12772 (N_12772,N_10666,N_11903);
nand U12773 (N_12773,N_10020,N_11489);
nor U12774 (N_12774,N_9378,N_10342);
or U12775 (N_12775,N_9568,N_10895);
nand U12776 (N_12776,N_10554,N_9778);
or U12777 (N_12777,N_9975,N_10510);
or U12778 (N_12778,N_9802,N_10801);
nor U12779 (N_12779,N_9107,N_11735);
and U12780 (N_12780,N_11307,N_10081);
nor U12781 (N_12781,N_9103,N_11203);
nor U12782 (N_12782,N_10511,N_9385);
nor U12783 (N_12783,N_9488,N_11999);
and U12784 (N_12784,N_9252,N_11353);
xnor U12785 (N_12785,N_9251,N_10547);
and U12786 (N_12786,N_10585,N_11468);
nor U12787 (N_12787,N_9834,N_10172);
and U12788 (N_12788,N_9490,N_11452);
xor U12789 (N_12789,N_11599,N_9829);
nor U12790 (N_12790,N_10580,N_9905);
nor U12791 (N_12791,N_9947,N_9618);
nor U12792 (N_12792,N_11551,N_10536);
and U12793 (N_12793,N_9315,N_9736);
and U12794 (N_12794,N_9789,N_9583);
and U12795 (N_12795,N_11606,N_10790);
and U12796 (N_12796,N_11977,N_10900);
or U12797 (N_12797,N_10717,N_11598);
nor U12798 (N_12798,N_9010,N_9259);
or U12799 (N_12799,N_11586,N_11617);
nand U12800 (N_12800,N_11689,N_10242);
or U12801 (N_12801,N_9219,N_9728);
and U12802 (N_12802,N_10091,N_9933);
and U12803 (N_12803,N_9684,N_9191);
nand U12804 (N_12804,N_11403,N_11168);
nor U12805 (N_12805,N_9314,N_9604);
and U12806 (N_12806,N_9296,N_11182);
and U12807 (N_12807,N_11615,N_10918);
nand U12808 (N_12808,N_11962,N_9057);
and U12809 (N_12809,N_11017,N_11751);
nor U12810 (N_12810,N_10227,N_11781);
nand U12811 (N_12811,N_11963,N_11154);
and U12812 (N_12812,N_9130,N_10544);
or U12813 (N_12813,N_10614,N_10842);
nor U12814 (N_12814,N_10629,N_10084);
and U12815 (N_12815,N_11843,N_10298);
or U12816 (N_12816,N_11612,N_10137);
and U12817 (N_12817,N_11467,N_9892);
nand U12818 (N_12818,N_9854,N_9741);
or U12819 (N_12819,N_10385,N_10608);
or U12820 (N_12820,N_11764,N_10079);
xnor U12821 (N_12821,N_9529,N_9910);
nand U12822 (N_12822,N_10702,N_10191);
nor U12823 (N_12823,N_9516,N_9064);
nor U12824 (N_12824,N_9570,N_9774);
xnor U12825 (N_12825,N_11659,N_10325);
nor U12826 (N_12826,N_10181,N_9833);
or U12827 (N_12827,N_11423,N_9081);
and U12828 (N_12828,N_10539,N_11791);
xor U12829 (N_12829,N_10162,N_9481);
nand U12830 (N_12830,N_9713,N_11811);
or U12831 (N_12831,N_11809,N_11731);
xnor U12832 (N_12832,N_9565,N_11065);
nand U12833 (N_12833,N_11642,N_10096);
xnor U12834 (N_12834,N_9172,N_11924);
nor U12835 (N_12835,N_10033,N_11092);
and U12836 (N_12836,N_11302,N_9439);
nor U12837 (N_12837,N_10800,N_11814);
nor U12838 (N_12838,N_9867,N_10054);
nand U12839 (N_12839,N_9637,N_11180);
or U12840 (N_12840,N_10774,N_11142);
and U12841 (N_12841,N_10581,N_10651);
or U12842 (N_12842,N_10848,N_10723);
nor U12843 (N_12843,N_9890,N_10477);
and U12844 (N_12844,N_10388,N_10640);
and U12845 (N_12845,N_10838,N_10911);
xnor U12846 (N_12846,N_10745,N_9330);
or U12847 (N_12847,N_11616,N_9941);
and U12848 (N_12848,N_10291,N_11284);
and U12849 (N_12849,N_10966,N_10837);
and U12850 (N_12850,N_11583,N_11379);
and U12851 (N_12851,N_11495,N_11445);
nor U12852 (N_12852,N_10912,N_10756);
nand U12853 (N_12853,N_11685,N_9942);
nor U12854 (N_12854,N_11883,N_9518);
nand U12855 (N_12855,N_11075,N_9886);
nand U12856 (N_12856,N_10463,N_9207);
xor U12857 (N_12857,N_11336,N_10066);
and U12858 (N_12858,N_11779,N_10121);
and U12859 (N_12859,N_11287,N_10525);
nor U12860 (N_12860,N_10622,N_11298);
nor U12861 (N_12861,N_10661,N_9264);
and U12862 (N_12862,N_11247,N_11398);
nand U12863 (N_12863,N_11918,N_10067);
nor U12864 (N_12864,N_11554,N_11863);
nor U12865 (N_12865,N_9084,N_10451);
and U12866 (N_12866,N_9682,N_11820);
or U12867 (N_12867,N_9871,N_9061);
or U12868 (N_12868,N_9256,N_11490);
nor U12869 (N_12869,N_10861,N_9299);
or U12870 (N_12870,N_11739,N_11518);
nand U12871 (N_12871,N_10214,N_9052);
and U12872 (N_12872,N_9344,N_9487);
nor U12873 (N_12873,N_9600,N_9027);
nand U12874 (N_12874,N_10029,N_10457);
xnor U12875 (N_12875,N_9431,N_11935);
nor U12876 (N_12876,N_10221,N_9700);
or U12877 (N_12877,N_10500,N_9255);
and U12878 (N_12878,N_9390,N_11131);
or U12879 (N_12879,N_11552,N_11116);
or U12880 (N_12880,N_11602,N_11095);
nand U12881 (N_12881,N_9016,N_10948);
xor U12882 (N_12882,N_11003,N_10024);
or U12883 (N_12883,N_9007,N_9985);
nand U12884 (N_12884,N_11983,N_11902);
nor U12885 (N_12885,N_9423,N_11222);
nand U12886 (N_12886,N_9450,N_11183);
nand U12887 (N_12887,N_11571,N_11869);
or U12888 (N_12888,N_10993,N_9372);
nand U12889 (N_12889,N_11317,N_9852);
nor U12890 (N_12890,N_10046,N_10873);
and U12891 (N_12891,N_9286,N_10749);
nor U12892 (N_12892,N_10724,N_9784);
xnor U12893 (N_12893,N_9216,N_10188);
and U12894 (N_12894,N_11099,N_10428);
xor U12895 (N_12895,N_11031,N_9594);
and U12896 (N_12896,N_9164,N_9499);
nand U12897 (N_12897,N_11437,N_11446);
and U12898 (N_12898,N_9323,N_11013);
or U12899 (N_12899,N_9676,N_10994);
and U12900 (N_12900,N_10803,N_10297);
and U12901 (N_12901,N_11419,N_10237);
nand U12902 (N_12902,N_10351,N_10266);
or U12903 (N_12903,N_11845,N_11545);
nor U12904 (N_12904,N_11126,N_11198);
nand U12905 (N_12905,N_9644,N_11777);
xor U12906 (N_12906,N_11979,N_9399);
nand U12907 (N_12907,N_11597,N_11620);
nand U12908 (N_12908,N_11356,N_9737);
or U12909 (N_12909,N_9744,N_10062);
nand U12910 (N_12910,N_11451,N_11553);
nor U12911 (N_12911,N_9739,N_9800);
xnor U12912 (N_12912,N_11532,N_10910);
nor U12913 (N_12913,N_10308,N_11945);
nor U12914 (N_12914,N_11111,N_10853);
or U12915 (N_12915,N_11590,N_10527);
and U12916 (N_12916,N_10663,N_9828);
nor U12917 (N_12917,N_9681,N_11277);
and U12918 (N_12918,N_11475,N_9305);
nor U12919 (N_12919,N_11509,N_9830);
nand U12920 (N_12920,N_9859,N_10102);
nor U12921 (N_12921,N_9268,N_11930);
xor U12922 (N_12922,N_10778,N_9363);
xnor U12923 (N_12923,N_10251,N_9436);
nand U12924 (N_12924,N_11102,N_9734);
nand U12925 (N_12925,N_10889,N_11772);
nor U12926 (N_12926,N_9675,N_10349);
nand U12927 (N_12927,N_11015,N_11871);
and U12928 (N_12928,N_10988,N_10106);
nand U12929 (N_12929,N_9122,N_10147);
or U12930 (N_12930,N_9181,N_11115);
nor U12931 (N_12931,N_10405,N_9669);
nor U12932 (N_12932,N_10633,N_11758);
or U12933 (N_12933,N_10938,N_9814);
and U12934 (N_12934,N_11407,N_9504);
nor U12935 (N_12935,N_11862,N_9612);
nand U12936 (N_12936,N_9915,N_11998);
and U12937 (N_12937,N_11951,N_11810);
or U12938 (N_12938,N_11050,N_11870);
or U12939 (N_12939,N_9573,N_10959);
nand U12940 (N_12940,N_10249,N_11022);
and U12941 (N_12941,N_11480,N_10187);
nor U12942 (N_12942,N_9577,N_11802);
nand U12943 (N_12943,N_10710,N_11868);
nand U12944 (N_12944,N_11968,N_11964);
nor U12945 (N_12945,N_11637,N_11314);
xor U12946 (N_12946,N_9732,N_9729);
and U12947 (N_12947,N_10112,N_11594);
nor U12948 (N_12948,N_11825,N_10330);
or U12949 (N_12949,N_10382,N_10776);
and U12950 (N_12950,N_11245,N_11061);
and U12951 (N_12951,N_10257,N_10127);
or U12952 (N_12952,N_10345,N_11544);
xor U12953 (N_12953,N_10557,N_11948);
nand U12954 (N_12954,N_11674,N_10199);
nand U12955 (N_12955,N_10696,N_11274);
nand U12956 (N_12956,N_11663,N_10442);
and U12957 (N_12957,N_10238,N_9370);
or U12958 (N_12958,N_10708,N_10995);
xor U12959 (N_12959,N_9293,N_10846);
nand U12960 (N_12960,N_9123,N_10010);
and U12961 (N_12961,N_9751,N_9953);
nor U12962 (N_12962,N_10076,N_10472);
nor U12963 (N_12963,N_9542,N_11909);
nand U12964 (N_12964,N_11793,N_11038);
and U12965 (N_12965,N_10458,N_11690);
and U12966 (N_12966,N_9864,N_10997);
nand U12967 (N_12967,N_10309,N_9046);
and U12968 (N_12968,N_9602,N_11943);
or U12969 (N_12969,N_10486,N_11749);
nor U12970 (N_12970,N_11433,N_10762);
and U12971 (N_12971,N_10600,N_9063);
nor U12972 (N_12972,N_9698,N_11523);
and U12973 (N_12973,N_11947,N_11212);
and U12974 (N_12974,N_11188,N_11320);
or U12975 (N_12975,N_10720,N_10031);
or U12976 (N_12976,N_9434,N_10568);
and U12977 (N_12977,N_11485,N_11801);
nor U12978 (N_12978,N_10459,N_11785);
and U12979 (N_12979,N_10782,N_9621);
nand U12980 (N_12980,N_9367,N_10197);
or U12981 (N_12981,N_9376,N_10533);
and U12982 (N_12982,N_10418,N_11164);
and U12983 (N_12983,N_9097,N_11533);
or U12984 (N_12984,N_9206,N_9863);
and U12985 (N_12985,N_10329,N_9514);
nor U12986 (N_12986,N_10160,N_11420);
or U12987 (N_12987,N_11139,N_10262);
or U12988 (N_12988,N_10193,N_10101);
xor U12989 (N_12989,N_9317,N_9980);
or U12990 (N_12990,N_10311,N_9117);
xnor U12991 (N_12991,N_11727,N_10048);
and U12992 (N_12992,N_11579,N_10725);
nor U12993 (N_12993,N_9111,N_11803);
or U12994 (N_12994,N_11316,N_11582);
xnor U12995 (N_12995,N_10087,N_11206);
and U12996 (N_12996,N_10484,N_9348);
or U12997 (N_12997,N_11768,N_9845);
nand U12998 (N_12998,N_10894,N_9950);
or U12999 (N_12999,N_9448,N_9592);
or U13000 (N_13000,N_11647,N_11070);
or U13001 (N_13001,N_11449,N_9438);
and U13002 (N_13002,N_9723,N_11682);
nor U13003 (N_13003,N_9214,N_11002);
nand U13004 (N_13004,N_10630,N_10245);
and U13005 (N_13005,N_11009,N_10699);
nand U13006 (N_13006,N_10053,N_10116);
nand U13007 (N_13007,N_10908,N_10780);
and U13008 (N_13008,N_9846,N_11321);
nor U13009 (N_13009,N_11228,N_9632);
and U13010 (N_13010,N_10902,N_9537);
and U13011 (N_13011,N_11787,N_11972);
nor U13012 (N_13012,N_11412,N_11044);
xnor U13013 (N_13013,N_10244,N_10403);
nor U13014 (N_13014,N_10574,N_9133);
xor U13015 (N_13015,N_9391,N_10564);
xor U13016 (N_13016,N_10070,N_9146);
and U13017 (N_13017,N_11334,N_9960);
nand U13018 (N_13018,N_11376,N_9076);
or U13019 (N_13019,N_11557,N_9693);
nand U13020 (N_13020,N_9055,N_10777);
nor U13021 (N_13021,N_11905,N_10946);
or U13022 (N_13022,N_9591,N_9241);
nor U13023 (N_13023,N_11359,N_9633);
or U13024 (N_13024,N_11077,N_11129);
and U13025 (N_13025,N_9138,N_10786);
or U13026 (N_13026,N_11358,N_10467);
nor U13027 (N_13027,N_10138,N_10933);
nand U13028 (N_13028,N_11643,N_10677);
or U13029 (N_13029,N_9595,N_10206);
nand U13030 (N_13030,N_10347,N_10515);
and U13031 (N_13031,N_11629,N_11700);
or U13032 (N_13032,N_10875,N_11120);
or U13033 (N_13033,N_10607,N_10693);
or U13034 (N_13034,N_9320,N_9855);
nor U13035 (N_13035,N_11995,N_10479);
nand U13036 (N_13036,N_10374,N_9498);
xor U13037 (N_13037,N_9393,N_9228);
nand U13038 (N_13038,N_10605,N_9340);
and U13039 (N_13039,N_11693,N_9777);
nor U13040 (N_13040,N_11770,N_11782);
nor U13041 (N_13041,N_10230,N_10821);
and U13042 (N_13042,N_10668,N_9764);
nand U13043 (N_13043,N_9098,N_11440);
and U13044 (N_13044,N_9609,N_9961);
and U13045 (N_13045,N_9776,N_9747);
nand U13046 (N_13046,N_10531,N_10516);
nor U13047 (N_13047,N_11992,N_11005);
nor U13048 (N_13048,N_11934,N_10609);
and U13049 (N_13049,N_11892,N_11112);
nor U13050 (N_13050,N_11504,N_11364);
and U13051 (N_13051,N_11684,N_10148);
nand U13052 (N_13052,N_11506,N_9539);
nand U13053 (N_13053,N_9371,N_9793);
and U13054 (N_13054,N_10530,N_10518);
nor U13055 (N_13055,N_11836,N_9300);
xnor U13056 (N_13056,N_10383,N_10265);
and U13057 (N_13057,N_11474,N_10213);
or U13058 (N_13058,N_9086,N_9979);
nor U13059 (N_13059,N_9277,N_9977);
nand U13060 (N_13060,N_9903,N_9333);
nand U13061 (N_13061,N_11737,N_11874);
or U13062 (N_13062,N_9598,N_9077);
nor U13063 (N_13063,N_9358,N_11421);
or U13064 (N_13064,N_9302,N_9053);
nor U13065 (N_13065,N_11191,N_9795);
and U13066 (N_13066,N_9072,N_11034);
xor U13067 (N_13067,N_9532,N_9202);
or U13068 (N_13068,N_9937,N_9069);
nand U13069 (N_13069,N_10787,N_10055);
nand U13070 (N_13070,N_9043,N_11230);
xnor U13071 (N_13071,N_9401,N_10641);
or U13072 (N_13072,N_9815,N_9672);
or U13073 (N_13073,N_11954,N_9088);
xnor U13074 (N_13074,N_9379,N_9731);
nand U13075 (N_13075,N_11066,N_11332);
or U13076 (N_13076,N_9809,N_9220);
nand U13077 (N_13077,N_10461,N_9821);
nand U13078 (N_13078,N_10689,N_11936);
nand U13079 (N_13079,N_10505,N_10563);
nor U13080 (N_13080,N_11283,N_10793);
nand U13081 (N_13081,N_10034,N_9550);
or U13082 (N_13082,N_10346,N_9132);
nand U13083 (N_13083,N_11539,N_9882);
or U13084 (N_13084,N_9486,N_9500);
and U13085 (N_13085,N_9155,N_11305);
nor U13086 (N_13086,N_11488,N_9192);
nand U13087 (N_13087,N_11562,N_10840);
xnor U13088 (N_13088,N_11652,N_11355);
nor U13089 (N_13089,N_9156,N_10635);
and U13090 (N_13090,N_9177,N_11621);
and U13091 (N_13091,N_10471,N_11694);
and U13092 (N_13092,N_10226,N_11499);
or U13093 (N_13093,N_9928,N_9711);
or U13094 (N_13094,N_11826,N_9624);
nand U13095 (N_13095,N_9273,N_11666);
xnor U13096 (N_13096,N_11725,N_10326);
and U13097 (N_13097,N_10526,N_9236);
nor U13098 (N_13098,N_11150,N_10923);
and U13099 (N_13099,N_10409,N_9807);
nor U13100 (N_13100,N_9411,N_10149);
and U13101 (N_13101,N_10917,N_10784);
nand U13102 (N_13102,N_9753,N_10864);
and U13103 (N_13103,N_10492,N_11186);
or U13104 (N_13104,N_10545,N_11707);
nand U13105 (N_13105,N_11155,N_11004);
nor U13106 (N_13106,N_10851,N_11330);
and U13107 (N_13107,N_9654,N_9574);
and U13108 (N_13108,N_10754,N_9429);
or U13109 (N_13109,N_10769,N_9110);
nor U13110 (N_13110,N_11447,N_10901);
nor U13111 (N_13111,N_10532,N_10604);
nor U13112 (N_13112,N_10427,N_10144);
nor U13113 (N_13113,N_10290,N_11950);
or U13114 (N_13114,N_9170,N_10791);
xnor U13115 (N_13115,N_9444,N_9312);
and U13116 (N_13116,N_9714,N_10304);
nand U13117 (N_13117,N_10366,N_10958);
and U13118 (N_13118,N_9417,N_9025);
nand U13119 (N_13119,N_9909,N_9718);
and U13120 (N_13120,N_9952,N_9449);
nor U13121 (N_13121,N_10386,N_11842);
nor U13122 (N_13122,N_9395,N_10406);
or U13123 (N_13123,N_10610,N_11264);
and U13124 (N_13124,N_9667,N_9666);
nand U13125 (N_13125,N_10811,N_10369);
and U13126 (N_13126,N_10064,N_9352);
or U13127 (N_13127,N_9555,N_9683);
nand U13128 (N_13128,N_11697,N_11607);
nor U13129 (N_13129,N_10878,N_10830);
nand U13130 (N_13130,N_11852,N_10205);
nor U13131 (N_13131,N_9464,N_10030);
nand U13132 (N_13132,N_10146,N_9318);
and U13133 (N_13133,N_10466,N_11249);
and U13134 (N_13134,N_9511,N_9822);
and U13135 (N_13135,N_9509,N_11743);
and U13136 (N_13136,N_10849,N_11591);
or U13137 (N_13137,N_9710,N_10078);
nand U13138 (N_13138,N_11658,N_11730);
nor U13139 (N_13139,N_11372,N_10562);
nand U13140 (N_13140,N_11208,N_9492);
nand U13141 (N_13141,N_11471,N_10072);
nor U13142 (N_13142,N_10125,N_11876);
or U13143 (N_13143,N_10643,N_11639);
or U13144 (N_13144,N_9523,N_10400);
nor U13145 (N_13145,N_10222,N_11171);
or U13146 (N_13146,N_11466,N_9677);
or U13147 (N_13147,N_10578,N_10903);
xnor U13148 (N_13148,N_9389,N_9556);
and U13149 (N_13149,N_11271,N_10596);
or U13150 (N_13150,N_11351,N_10395);
nor U13151 (N_13151,N_10421,N_10168);
nand U13152 (N_13152,N_9160,N_10582);
nand U13153 (N_13153,N_10314,N_11464);
and U13154 (N_13154,N_10674,N_11339);
nor U13155 (N_13155,N_9923,N_11073);
or U13156 (N_13156,N_9443,N_9832);
nor U13157 (N_13157,N_9733,N_10464);
nand U13158 (N_13158,N_9037,N_11896);
or U13159 (N_13159,N_9564,N_10201);
and U13160 (N_13160,N_9872,N_11653);
nor U13161 (N_13161,N_10978,N_9485);
nor U13162 (N_13162,N_11736,N_9375);
or U13163 (N_13163,N_11160,N_10540);
nand U13164 (N_13164,N_10022,N_11701);
nor U13165 (N_13165,N_11237,N_10111);
nor U13166 (N_13166,N_11980,N_10927);
or U13167 (N_13167,N_11348,N_11303);
xnor U13168 (N_13168,N_11806,N_9749);
or U13169 (N_13169,N_11920,N_11278);
or U13170 (N_13170,N_10195,N_10017);
and U13171 (N_13171,N_11136,N_11548);
nand U13172 (N_13172,N_11080,N_10322);
xnor U13173 (N_13173,N_9503,N_11323);
nor U13174 (N_13174,N_9147,N_11513);
and U13175 (N_13175,N_11008,N_10658);
xor U13176 (N_13176,N_10519,N_9869);
xor U13177 (N_13177,N_11378,N_9139);
nand U13178 (N_13178,N_10173,N_10339);
nand U13179 (N_13179,N_11575,N_11500);
or U13180 (N_13180,N_11134,N_10005);
xor U13181 (N_13181,N_10854,N_9491);
nor U13182 (N_13182,N_11014,N_9223);
or U13183 (N_13183,N_10327,N_9032);
nor U13184 (N_13184,N_11604,N_11887);
nor U13185 (N_13185,N_11296,N_9408);
and U13186 (N_13186,N_11380,N_9480);
and U13187 (N_13187,N_10771,N_11254);
and U13188 (N_13188,N_9100,N_10883);
nor U13189 (N_13189,N_9973,N_11786);
nand U13190 (N_13190,N_9193,N_11699);
nor U13191 (N_13191,N_9035,N_9396);
nand U13192 (N_13192,N_11105,N_11219);
and U13193 (N_13193,N_9839,N_10219);
and U13194 (N_13194,N_10077,N_9590);
or U13195 (N_13195,N_9188,N_9335);
or U13196 (N_13196,N_11169,N_9253);
and U13197 (N_13197,N_9102,N_10719);
or U13198 (N_13198,N_10847,N_9868);
xor U13199 (N_13199,N_10412,N_10362);
or U13200 (N_13200,N_11373,N_11840);
nand U13201 (N_13201,N_10378,N_11322);
xor U13202 (N_13202,N_10844,N_10273);
nand U13203 (N_13203,N_9022,N_11217);
and U13204 (N_13204,N_10085,N_11744);
xnor U13205 (N_13205,N_11200,N_9141);
xnor U13206 (N_13206,N_10956,N_9085);
nor U13207 (N_13207,N_9406,N_10645);
or U13208 (N_13208,N_11778,N_9989);
nor U13209 (N_13209,N_9143,N_9898);
nand U13210 (N_13210,N_10955,N_10373);
or U13211 (N_13211,N_10083,N_9561);
nand U13212 (N_13212,N_11927,N_10280);
nor U13213 (N_13213,N_11853,N_10558);
nand U13214 (N_13214,N_9651,N_11893);
and U13215 (N_13215,N_11374,N_10650);
or U13216 (N_13216,N_11045,N_10928);
nor U13217 (N_13217,N_9265,N_11763);
or U13218 (N_13218,N_11472,N_10968);
nand U13219 (N_13219,N_9048,N_10234);
or U13220 (N_13220,N_11248,N_10681);
or U13221 (N_13221,N_10827,N_9019);
or U13222 (N_13222,N_9525,N_11595);
nand U13223 (N_13223,N_10758,N_10626);
nand U13224 (N_13224,N_10572,N_9127);
or U13225 (N_13225,N_11285,N_9074);
or U13226 (N_13226,N_10930,N_9040);
nor U13227 (N_13227,N_10740,N_10475);
and U13228 (N_13228,N_11346,N_11176);
or U13229 (N_13229,N_10617,N_11683);
or U13230 (N_13230,N_11124,N_11815);
or U13231 (N_13231,N_11048,N_11555);
and U13232 (N_13232,N_9159,N_11794);
nand U13233 (N_13233,N_10343,N_11668);
nand U13234 (N_13234,N_11377,N_9060);
or U13235 (N_13235,N_10603,N_9663);
nand U13236 (N_13236,N_9038,N_9269);
or U13237 (N_13237,N_9169,N_9906);
or U13238 (N_13238,N_11716,N_10443);
xor U13239 (N_13239,N_9244,N_9790);
or U13240 (N_13240,N_9342,N_9601);
nand U13241 (N_13241,N_11162,N_9824);
nor U13242 (N_13242,N_10286,N_9289);
xor U13243 (N_13243,N_10223,N_9920);
xor U13244 (N_13244,N_9137,N_9966);
nand U13245 (N_13245,N_9249,N_11030);
nand U13246 (N_13246,N_11921,N_11667);
nor U13247 (N_13247,N_9769,N_11573);
nand U13248 (N_13248,N_9557,N_11958);
nor U13249 (N_13249,N_9978,N_11366);
nand U13250 (N_13250,N_9857,N_11879);
nor U13251 (N_13251,N_9339,N_11775);
and U13252 (N_13252,N_9222,N_11293);
nor U13253 (N_13253,N_11436,N_11012);
or U13254 (N_13254,N_9671,N_9297);
nor U13255 (N_13255,N_11550,N_9722);
and U13256 (N_13256,N_9240,N_11438);
xnor U13257 (N_13257,N_9331,N_10156);
and U13258 (N_13258,N_11904,N_9904);
nand U13259 (N_13259,N_10962,N_9689);
and U13260 (N_13260,N_11496,N_9917);
nand U13261 (N_13261,N_10480,N_9291);
xor U13262 (N_13262,N_9705,N_9190);
nand U13263 (N_13263,N_11062,N_10592);
or U13264 (N_13264,N_11047,N_9918);
or U13265 (N_13265,N_10969,N_10224);
nand U13266 (N_13266,N_11641,N_10991);
or U13267 (N_13267,N_11765,N_10686);
and U13268 (N_13268,N_11795,N_10231);
and U13269 (N_13269,N_11174,N_11767);
and U13270 (N_13270,N_9578,N_10186);
nor U13271 (N_13271,N_11835,N_10936);
and U13272 (N_13272,N_9310,N_9629);
or U13273 (N_13273,N_11244,N_10766);
and U13274 (N_13274,N_10370,N_11481);
nand U13275 (N_13275,N_11648,N_9020);
nor U13276 (N_13276,N_10375,N_9092);
and U13277 (N_13277,N_9215,N_11101);
and U13278 (N_13278,N_11738,N_9182);
and U13279 (N_13279,N_10041,N_9151);
nand U13280 (N_13280,N_11411,N_11726);
and U13281 (N_13281,N_11928,N_9461);
xnor U13282 (N_13282,N_11096,N_9911);
nand U13283 (N_13283,N_9109,N_9014);
nand U13284 (N_13284,N_11866,N_9520);
and U13285 (N_13285,N_10992,N_11503);
or U13286 (N_13286,N_10688,N_11837);
xor U13287 (N_13287,N_11326,N_10410);
xor U13288 (N_13288,N_11537,N_9232);
nand U13289 (N_13289,N_10348,N_11832);
xor U13290 (N_13290,N_10865,N_11172);
nand U13291 (N_13291,N_9897,N_11953);
xor U13292 (N_13292,N_10063,N_11799);
and U13293 (N_13293,N_11032,N_10263);
nor U13294 (N_13294,N_9238,N_10209);
nand U13295 (N_13295,N_9530,N_11486);
nor U13296 (N_13296,N_11657,N_10036);
and U13297 (N_13297,N_11273,N_11367);
nand U13298 (N_13298,N_10555,N_11453);
or U13299 (N_13299,N_9665,N_11824);
nand U13300 (N_13300,N_9018,N_9327);
nand U13301 (N_13301,N_10852,N_9742);
xor U13302 (N_13302,N_9721,N_9246);
nor U13303 (N_13303,N_9473,N_10389);
and U13304 (N_13304,N_9605,N_11841);
or U13305 (N_13305,N_11289,N_9006);
nor U13306 (N_13306,N_11197,N_11294);
nand U13307 (N_13307,N_11520,N_9823);
nand U13308 (N_13308,N_9089,N_11385);
nor U13309 (N_13309,N_9870,N_11563);
and U13310 (N_13310,N_9717,N_9004);
nand U13311 (N_13311,N_11313,N_10433);
nand U13312 (N_13312,N_9691,N_10225);
or U13313 (N_13313,N_11304,N_10026);
or U13314 (N_13314,N_9198,N_11108);
nand U13315 (N_13315,N_9768,N_10802);
nor U13316 (N_13316,N_11020,N_11524);
and U13317 (N_13317,N_10157,N_10957);
and U13318 (N_13318,N_10454,N_11937);
and U13319 (N_13319,N_10100,N_10359);
nor U13320 (N_13320,N_10452,N_11147);
or U13321 (N_13321,N_10073,N_10858);
or U13322 (N_13322,N_11391,N_11482);
or U13323 (N_13323,N_11941,N_11745);
or U13324 (N_13324,N_11456,N_11976);
xor U13325 (N_13325,N_9881,N_10363);
or U13326 (N_13326,N_10493,N_9521);
nand U13327 (N_13327,N_9336,N_9162);
nor U13328 (N_13328,N_11610,N_10274);
and U13329 (N_13329,N_9506,N_11349);
or U13330 (N_13330,N_10602,N_10669);
nand U13331 (N_13331,N_9679,N_11100);
or U13332 (N_13332,N_9308,N_10561);
or U13333 (N_13333,N_10577,N_9607);
nor U13334 (N_13334,N_11057,N_11984);
or U13335 (N_13335,N_11677,N_11856);
nand U13336 (N_13336,N_10660,N_10232);
or U13337 (N_13337,N_10080,N_11130);
nand U13338 (N_13338,N_11748,N_9922);
nand U13339 (N_13339,N_10934,N_10153);
nand U13340 (N_13340,N_11431,N_9384);
xnor U13341 (N_13341,N_9078,N_9929);
xor U13342 (N_13342,N_10880,N_9425);
nor U13343 (N_13343,N_11549,N_11619);
xor U13344 (N_13344,N_11309,N_11932);
nor U13345 (N_13345,N_11097,N_9770);
and U13346 (N_13346,N_11215,N_11040);
or U13347 (N_13347,N_10657,N_11651);
and U13348 (N_13348,N_9290,N_9387);
and U13349 (N_13349,N_9140,N_11880);
nand U13350 (N_13350,N_10267,N_11792);
nand U13351 (N_13351,N_9242,N_10277);
and U13352 (N_13352,N_11511,N_11886);
nand U13353 (N_13353,N_9642,N_11156);
and U13354 (N_13354,N_9373,N_10008);
and U13355 (N_13355,N_11714,N_10151);
or U13356 (N_13356,N_10951,N_9522);
xnor U13357 (N_13357,N_9934,N_9478);
or U13358 (N_13358,N_9662,N_10703);
nand U13359 (N_13359,N_11058,N_10888);
nor U13360 (N_13360,N_11170,N_9546);
or U13361 (N_13361,N_11626,N_9559);
xor U13362 (N_13362,N_9932,N_10898);
or U13363 (N_13363,N_10057,N_9945);
or U13364 (N_13364,N_9836,N_9617);
xor U13365 (N_13365,N_11362,N_10336);
and U13366 (N_13366,N_9225,N_10586);
and U13367 (N_13367,N_9670,N_10684);
nand U13368 (N_13368,N_11286,N_10517);
xnor U13369 (N_13369,N_9647,N_10704);
and U13370 (N_13370,N_9105,N_10012);
nand U13371 (N_13371,N_10721,N_10819);
or U13372 (N_13372,N_10866,N_9819);
xnor U13373 (N_13373,N_10964,N_10058);
nor U13374 (N_13374,N_10736,N_11494);
nand U13375 (N_13375,N_9620,N_11630);
xor U13376 (N_13376,N_11337,N_10098);
nand U13377 (N_13377,N_9173,N_10976);
or U13378 (N_13378,N_9458,N_11064);
nor U13379 (N_13379,N_11127,N_11055);
xnor U13380 (N_13380,N_10275,N_9687);
nand U13381 (N_13381,N_11565,N_9042);
and U13382 (N_13382,N_9196,N_9861);
xnor U13383 (N_13383,N_10737,N_10021);
or U13384 (N_13384,N_11393,N_9380);
nand U13385 (N_13385,N_11942,N_10117);
nor U13386 (N_13386,N_11720,N_9412);
nor U13387 (N_13387,N_10509,N_11184);
xnor U13388 (N_13388,N_11461,N_10377);
nand U13389 (N_13389,N_11634,N_10332);
or U13390 (N_13390,N_10649,N_11011);
or U13391 (N_13391,N_10126,N_10089);
or U13392 (N_13392,N_11114,N_9628);
or U13393 (N_13393,N_10535,N_10455);
and U13394 (N_13394,N_10236,N_10246);
nor U13395 (N_13395,N_10690,N_11067);
xnor U13396 (N_13396,N_11889,N_11270);
or U13397 (N_13397,N_11457,N_10044);
nand U13398 (N_13398,N_11177,N_9851);
nor U13399 (N_13399,N_9394,N_11891);
and U13400 (N_13400,N_11860,N_9337);
nand U13401 (N_13401,N_11628,N_11018);
and U13402 (N_13402,N_11717,N_9245);
nand U13403 (N_13403,N_9250,N_9462);
nor U13404 (N_13404,N_10970,N_11469);
and U13405 (N_13405,N_9659,N_9944);
xor U13406 (N_13406,N_9566,N_9619);
xnor U13407 (N_13407,N_11396,N_11216);
nor U13408 (N_13408,N_9827,N_10797);
and U13409 (N_13409,N_11605,N_10007);
nand U13410 (N_13410,N_9316,N_10328);
xor U13411 (N_13411,N_9974,N_9608);
xor U13412 (N_13412,N_10628,N_9031);
or U13413 (N_13413,N_11152,N_11335);
nand U13414 (N_13414,N_9199,N_9468);
and U13415 (N_13415,N_10759,N_9841);
nor U13416 (N_13416,N_11864,N_11578);
nor U13417 (N_13417,N_9535,N_9484);
nand U13418 (N_13418,N_10656,N_10051);
or U13419 (N_13419,N_10559,N_10913);
and U13420 (N_13420,N_10408,N_9582);
nor U13421 (N_13421,N_10727,N_11218);
xor U13422 (N_13422,N_11780,N_11709);
or U13423 (N_13423,N_9073,N_10579);
xnor U13424 (N_13424,N_10175,N_11361);
xnor U13425 (N_13425,N_11993,N_10798);
or U13426 (N_13426,N_10118,N_11179);
nand U13427 (N_13427,N_11268,N_11258);
nand U13428 (N_13428,N_9902,N_11415);
nor U13429 (N_13429,N_11432,N_11318);
nor U13430 (N_13430,N_10885,N_11813);
nand U13431 (N_13431,N_11712,N_10060);
and U13432 (N_13432,N_9366,N_9304);
nor U13433 (N_13433,N_9584,N_11081);
and U13434 (N_13434,N_10623,N_10393);
nor U13435 (N_13435,N_9756,N_10059);
and U13436 (N_13436,N_10283,N_11982);
and U13437 (N_13437,N_10099,N_11085);
or U13438 (N_13438,N_9951,N_9325);
or U13439 (N_13439,N_9274,N_10462);
nand U13440 (N_13440,N_10161,N_10884);
nor U13441 (N_13441,N_11187,N_10415);
xor U13442 (N_13442,N_11125,N_9984);
nor U13443 (N_13443,N_11771,N_9976);
nor U13444 (N_13444,N_10779,N_10281);
nor U13445 (N_13445,N_9991,N_9880);
or U13446 (N_13446,N_9474,N_11559);
or U13447 (N_13447,N_11241,N_9787);
nor U13448 (N_13448,N_10372,N_11711);
and U13449 (N_13449,N_9858,N_11783);
nor U13450 (N_13450,N_9760,N_10104);
or U13451 (N_13451,N_10424,N_10040);
and U13452 (N_13452,N_10589,N_11225);
xor U13453 (N_13453,N_11784,N_9720);
nand U13454 (N_13454,N_9033,N_10141);
and U13455 (N_13455,N_9763,N_9163);
and U13456 (N_13456,N_10705,N_10001);
or U13457 (N_13457,N_9571,N_11536);
nand U13458 (N_13458,N_11492,N_10169);
nand U13459 (N_13459,N_10529,N_10107);
nand U13460 (N_13460,N_9949,N_10522);
or U13461 (N_13461,N_10444,N_10761);
and U13462 (N_13462,N_9353,N_10356);
or U13463 (N_13463,N_10648,N_11961);
or U13464 (N_13464,N_9896,N_9581);
xor U13465 (N_13465,N_9931,N_10170);
nand U13466 (N_13466,N_10897,N_11133);
or U13467 (N_13467,N_9230,N_11600);
nor U13468 (N_13468,N_11354,N_9781);
and U13469 (N_13469,N_10939,N_9165);
or U13470 (N_13470,N_9895,N_9935);
and U13471 (N_13471,N_9636,N_10942);
nand U13472 (N_13472,N_9955,N_11645);
or U13473 (N_13473,N_9759,N_10987);
xnor U13474 (N_13474,N_11231,N_10028);
xnor U13475 (N_13475,N_9538,N_11493);
or U13476 (N_13476,N_11410,N_11708);
nor U13477 (N_13477,N_11673,N_11424);
xnor U13478 (N_13478,N_10352,N_9231);
and U13479 (N_13479,N_10673,N_10358);
and U13480 (N_13480,N_9021,N_11900);
and U13481 (N_13481,N_11872,N_10292);
and U13482 (N_13482,N_11949,N_10817);
or U13483 (N_13483,N_11473,N_10513);
nor U13484 (N_13484,N_9543,N_10940);
xor U13485 (N_13485,N_9059,N_11596);
or U13486 (N_13486,N_9655,N_11439);
nand U13487 (N_13487,N_9848,N_9748);
xor U13488 (N_13488,N_11308,N_11033);
xor U13489 (N_13489,N_10750,N_9884);
nand U13490 (N_13490,N_10990,N_11312);
nand U13491 (N_13491,N_10560,N_9056);
nand U13492 (N_13492,N_10019,N_9946);
or U13493 (N_13493,N_10196,N_9982);
nand U13494 (N_13494,N_11430,N_11797);
or U13495 (N_13495,N_10841,N_11132);
or U13496 (N_13496,N_10813,N_10229);
nor U13497 (N_13497,N_10013,N_11522);
and U13498 (N_13498,N_10398,N_10235);
and U13499 (N_13499,N_10506,N_10764);
nand U13500 (N_13500,N_9249,N_9623);
nand U13501 (N_13501,N_11943,N_10587);
and U13502 (N_13502,N_11187,N_9500);
nand U13503 (N_13503,N_10378,N_9982);
or U13504 (N_13504,N_10650,N_11489);
nand U13505 (N_13505,N_10147,N_11449);
nand U13506 (N_13506,N_11137,N_11053);
or U13507 (N_13507,N_9617,N_9794);
nor U13508 (N_13508,N_10307,N_10052);
or U13509 (N_13509,N_10439,N_9794);
nor U13510 (N_13510,N_9513,N_10805);
nor U13511 (N_13511,N_10891,N_11225);
nand U13512 (N_13512,N_9960,N_10809);
or U13513 (N_13513,N_11995,N_11040);
nand U13514 (N_13514,N_9223,N_9530);
nand U13515 (N_13515,N_10863,N_9785);
nand U13516 (N_13516,N_9312,N_11516);
and U13517 (N_13517,N_9727,N_10299);
and U13518 (N_13518,N_9627,N_10568);
or U13519 (N_13519,N_10319,N_9133);
or U13520 (N_13520,N_9533,N_9037);
nand U13521 (N_13521,N_10127,N_10867);
nand U13522 (N_13522,N_9706,N_11823);
or U13523 (N_13523,N_10913,N_11374);
or U13524 (N_13524,N_11637,N_11653);
or U13525 (N_13525,N_9251,N_11920);
and U13526 (N_13526,N_10572,N_11606);
nand U13527 (N_13527,N_10187,N_11601);
or U13528 (N_13528,N_10077,N_9008);
xnor U13529 (N_13529,N_9076,N_9183);
or U13530 (N_13530,N_10906,N_10762);
xor U13531 (N_13531,N_9870,N_9335);
and U13532 (N_13532,N_11240,N_11114);
and U13533 (N_13533,N_11992,N_11793);
xnor U13534 (N_13534,N_10469,N_10346);
and U13535 (N_13535,N_11009,N_9596);
or U13536 (N_13536,N_10943,N_9544);
xnor U13537 (N_13537,N_10701,N_9283);
and U13538 (N_13538,N_11135,N_11029);
xnor U13539 (N_13539,N_11359,N_11713);
nand U13540 (N_13540,N_11027,N_9477);
or U13541 (N_13541,N_11991,N_11440);
nand U13542 (N_13542,N_9343,N_9623);
nand U13543 (N_13543,N_9397,N_10362);
nor U13544 (N_13544,N_10695,N_10952);
nand U13545 (N_13545,N_10225,N_10362);
nand U13546 (N_13546,N_10380,N_10798);
nand U13547 (N_13547,N_10839,N_11074);
nand U13548 (N_13548,N_9646,N_10014);
and U13549 (N_13549,N_9971,N_11203);
or U13550 (N_13550,N_9523,N_10424);
nand U13551 (N_13551,N_11883,N_10809);
nor U13552 (N_13552,N_9405,N_11421);
nor U13553 (N_13553,N_10791,N_10993);
and U13554 (N_13554,N_9260,N_10214);
nand U13555 (N_13555,N_10743,N_9231);
and U13556 (N_13556,N_10918,N_9512);
or U13557 (N_13557,N_10083,N_10708);
nor U13558 (N_13558,N_10681,N_10486);
or U13559 (N_13559,N_11963,N_10396);
xor U13560 (N_13560,N_9231,N_11376);
nand U13561 (N_13561,N_11189,N_9316);
nor U13562 (N_13562,N_9574,N_9629);
and U13563 (N_13563,N_11260,N_10884);
and U13564 (N_13564,N_11702,N_9618);
nor U13565 (N_13565,N_10355,N_11374);
nand U13566 (N_13566,N_11049,N_10925);
or U13567 (N_13567,N_10788,N_10686);
nor U13568 (N_13568,N_10852,N_9668);
or U13569 (N_13569,N_9456,N_9961);
and U13570 (N_13570,N_9904,N_10977);
and U13571 (N_13571,N_11651,N_11505);
nand U13572 (N_13572,N_9331,N_11471);
nor U13573 (N_13573,N_9408,N_9386);
and U13574 (N_13574,N_9184,N_9265);
and U13575 (N_13575,N_11329,N_11341);
nor U13576 (N_13576,N_11332,N_9087);
nor U13577 (N_13577,N_10097,N_11086);
nor U13578 (N_13578,N_9315,N_10037);
nor U13579 (N_13579,N_10354,N_10788);
xor U13580 (N_13580,N_11571,N_11767);
and U13581 (N_13581,N_9433,N_9195);
nor U13582 (N_13582,N_11612,N_9750);
xnor U13583 (N_13583,N_9697,N_10600);
xor U13584 (N_13584,N_9553,N_9853);
nor U13585 (N_13585,N_11005,N_11013);
or U13586 (N_13586,N_9164,N_10749);
nand U13587 (N_13587,N_9285,N_11357);
or U13588 (N_13588,N_9793,N_9751);
nand U13589 (N_13589,N_10085,N_11508);
nand U13590 (N_13590,N_9494,N_11275);
or U13591 (N_13591,N_11715,N_9254);
xnor U13592 (N_13592,N_9415,N_10143);
nand U13593 (N_13593,N_9955,N_11631);
or U13594 (N_13594,N_11175,N_11219);
or U13595 (N_13595,N_11082,N_9966);
nor U13596 (N_13596,N_10569,N_11172);
nand U13597 (N_13597,N_11044,N_11718);
xnor U13598 (N_13598,N_10260,N_10640);
nor U13599 (N_13599,N_10350,N_11828);
and U13600 (N_13600,N_10941,N_9191);
and U13601 (N_13601,N_9446,N_11015);
and U13602 (N_13602,N_11505,N_10964);
nand U13603 (N_13603,N_10502,N_9211);
nor U13604 (N_13604,N_11436,N_10006);
xnor U13605 (N_13605,N_11063,N_10303);
nor U13606 (N_13606,N_9809,N_11554);
nor U13607 (N_13607,N_10116,N_10461);
nor U13608 (N_13608,N_10170,N_10745);
xnor U13609 (N_13609,N_10984,N_9764);
or U13610 (N_13610,N_11423,N_11629);
or U13611 (N_13611,N_11458,N_11918);
nor U13612 (N_13612,N_11199,N_10071);
and U13613 (N_13613,N_11510,N_10031);
or U13614 (N_13614,N_9016,N_9098);
and U13615 (N_13615,N_9681,N_11889);
nor U13616 (N_13616,N_9188,N_10028);
nand U13617 (N_13617,N_11287,N_9846);
nor U13618 (N_13618,N_9915,N_11339);
nand U13619 (N_13619,N_9109,N_9444);
or U13620 (N_13620,N_9467,N_9392);
nand U13621 (N_13621,N_10140,N_10026);
and U13622 (N_13622,N_10621,N_11037);
nor U13623 (N_13623,N_11828,N_9408);
and U13624 (N_13624,N_10057,N_9483);
or U13625 (N_13625,N_11074,N_9179);
xor U13626 (N_13626,N_11261,N_10674);
and U13627 (N_13627,N_10756,N_9973);
and U13628 (N_13628,N_10946,N_11728);
nand U13629 (N_13629,N_9250,N_11296);
and U13630 (N_13630,N_9827,N_10150);
nor U13631 (N_13631,N_11773,N_11463);
nand U13632 (N_13632,N_9416,N_9744);
and U13633 (N_13633,N_9500,N_9619);
and U13634 (N_13634,N_9679,N_11890);
or U13635 (N_13635,N_9411,N_10513);
or U13636 (N_13636,N_9966,N_11371);
and U13637 (N_13637,N_11425,N_10737);
nor U13638 (N_13638,N_10117,N_9757);
xor U13639 (N_13639,N_10953,N_10946);
or U13640 (N_13640,N_10166,N_10448);
nor U13641 (N_13641,N_10466,N_11421);
nor U13642 (N_13642,N_11326,N_9361);
nor U13643 (N_13643,N_11956,N_11325);
or U13644 (N_13644,N_11472,N_11808);
nor U13645 (N_13645,N_9770,N_11945);
or U13646 (N_13646,N_11919,N_9006);
nand U13647 (N_13647,N_10757,N_10146);
xor U13648 (N_13648,N_10789,N_11130);
nand U13649 (N_13649,N_10967,N_9388);
nor U13650 (N_13650,N_9191,N_9284);
or U13651 (N_13651,N_9172,N_9097);
and U13652 (N_13652,N_11498,N_10577);
nor U13653 (N_13653,N_11545,N_11540);
or U13654 (N_13654,N_10235,N_11585);
or U13655 (N_13655,N_11206,N_9474);
nand U13656 (N_13656,N_11991,N_10528);
nand U13657 (N_13657,N_10465,N_11869);
nand U13658 (N_13658,N_9256,N_9982);
and U13659 (N_13659,N_11064,N_10103);
nor U13660 (N_13660,N_10525,N_11216);
nor U13661 (N_13661,N_10017,N_10514);
nand U13662 (N_13662,N_10102,N_9989);
or U13663 (N_13663,N_10111,N_9904);
or U13664 (N_13664,N_10264,N_9207);
nor U13665 (N_13665,N_11076,N_9166);
nand U13666 (N_13666,N_11229,N_10003);
or U13667 (N_13667,N_11852,N_9188);
and U13668 (N_13668,N_10467,N_9909);
and U13669 (N_13669,N_10016,N_10626);
and U13670 (N_13670,N_10926,N_11154);
nor U13671 (N_13671,N_10239,N_9463);
and U13672 (N_13672,N_11315,N_10608);
or U13673 (N_13673,N_10337,N_10364);
nor U13674 (N_13674,N_11624,N_10581);
nand U13675 (N_13675,N_11135,N_10372);
xor U13676 (N_13676,N_9252,N_10839);
nor U13677 (N_13677,N_9102,N_11899);
and U13678 (N_13678,N_9224,N_11656);
and U13679 (N_13679,N_9657,N_9499);
nor U13680 (N_13680,N_9333,N_9577);
nand U13681 (N_13681,N_10933,N_10771);
nor U13682 (N_13682,N_11077,N_10518);
nor U13683 (N_13683,N_10426,N_11236);
or U13684 (N_13684,N_9099,N_10186);
or U13685 (N_13685,N_11336,N_10613);
and U13686 (N_13686,N_10843,N_9492);
and U13687 (N_13687,N_10606,N_9638);
nor U13688 (N_13688,N_9812,N_11671);
or U13689 (N_13689,N_11591,N_11210);
nand U13690 (N_13690,N_9639,N_11387);
xor U13691 (N_13691,N_11623,N_10145);
and U13692 (N_13692,N_9110,N_10319);
nor U13693 (N_13693,N_9619,N_10321);
or U13694 (N_13694,N_11548,N_11709);
and U13695 (N_13695,N_10018,N_11706);
and U13696 (N_13696,N_10652,N_11551);
or U13697 (N_13697,N_11481,N_9888);
xnor U13698 (N_13698,N_9251,N_11544);
nand U13699 (N_13699,N_10397,N_9507);
nor U13700 (N_13700,N_11757,N_9594);
and U13701 (N_13701,N_11170,N_9873);
nor U13702 (N_13702,N_9037,N_9494);
nand U13703 (N_13703,N_10334,N_9560);
xnor U13704 (N_13704,N_10988,N_10368);
and U13705 (N_13705,N_10476,N_9029);
nor U13706 (N_13706,N_10949,N_11410);
nor U13707 (N_13707,N_10288,N_10015);
nand U13708 (N_13708,N_10346,N_10986);
xor U13709 (N_13709,N_11384,N_10857);
nor U13710 (N_13710,N_10689,N_11096);
or U13711 (N_13711,N_9282,N_9393);
nor U13712 (N_13712,N_9303,N_10986);
or U13713 (N_13713,N_9452,N_11641);
or U13714 (N_13714,N_11049,N_10189);
nand U13715 (N_13715,N_10837,N_11491);
nand U13716 (N_13716,N_11358,N_10307);
or U13717 (N_13717,N_9476,N_11321);
xor U13718 (N_13718,N_10393,N_11046);
xor U13719 (N_13719,N_11332,N_10619);
or U13720 (N_13720,N_11275,N_11575);
and U13721 (N_13721,N_9762,N_9505);
nor U13722 (N_13722,N_11103,N_9061);
or U13723 (N_13723,N_11403,N_10070);
or U13724 (N_13724,N_11522,N_10394);
and U13725 (N_13725,N_10912,N_11503);
and U13726 (N_13726,N_11339,N_10463);
nand U13727 (N_13727,N_10029,N_10532);
nor U13728 (N_13728,N_10838,N_11558);
or U13729 (N_13729,N_11743,N_11518);
and U13730 (N_13730,N_9140,N_9676);
and U13731 (N_13731,N_9886,N_11638);
and U13732 (N_13732,N_10230,N_11161);
xor U13733 (N_13733,N_11772,N_10228);
xnor U13734 (N_13734,N_9180,N_11054);
nand U13735 (N_13735,N_10115,N_11496);
and U13736 (N_13736,N_11676,N_10564);
or U13737 (N_13737,N_11977,N_11420);
or U13738 (N_13738,N_11519,N_9549);
xnor U13739 (N_13739,N_10412,N_10327);
nand U13740 (N_13740,N_10185,N_10235);
or U13741 (N_13741,N_11047,N_9520);
nor U13742 (N_13742,N_9346,N_10601);
or U13743 (N_13743,N_9281,N_9535);
xnor U13744 (N_13744,N_9086,N_10443);
or U13745 (N_13745,N_11047,N_10596);
nand U13746 (N_13746,N_9371,N_9813);
nand U13747 (N_13747,N_9477,N_9566);
and U13748 (N_13748,N_11176,N_11078);
and U13749 (N_13749,N_11482,N_11261);
or U13750 (N_13750,N_9226,N_11753);
and U13751 (N_13751,N_11956,N_11340);
xor U13752 (N_13752,N_9556,N_11883);
or U13753 (N_13753,N_11669,N_11054);
or U13754 (N_13754,N_11602,N_9363);
or U13755 (N_13755,N_9103,N_10802);
or U13756 (N_13756,N_9369,N_11698);
nor U13757 (N_13757,N_9299,N_10042);
and U13758 (N_13758,N_11362,N_10732);
nor U13759 (N_13759,N_10183,N_10466);
and U13760 (N_13760,N_11755,N_9308);
nor U13761 (N_13761,N_9521,N_11428);
xnor U13762 (N_13762,N_11960,N_11555);
and U13763 (N_13763,N_10348,N_11578);
or U13764 (N_13764,N_11533,N_10800);
nand U13765 (N_13765,N_9134,N_9641);
xnor U13766 (N_13766,N_9224,N_9768);
and U13767 (N_13767,N_9366,N_11140);
and U13768 (N_13768,N_9008,N_10233);
nand U13769 (N_13769,N_10992,N_9589);
nand U13770 (N_13770,N_9204,N_9361);
xor U13771 (N_13771,N_11210,N_9416);
nand U13772 (N_13772,N_11326,N_11504);
and U13773 (N_13773,N_9808,N_9803);
nor U13774 (N_13774,N_10887,N_11647);
xor U13775 (N_13775,N_10720,N_11904);
and U13776 (N_13776,N_11695,N_10608);
and U13777 (N_13777,N_10390,N_11777);
and U13778 (N_13778,N_11194,N_11355);
nand U13779 (N_13779,N_11910,N_11121);
xor U13780 (N_13780,N_11927,N_11170);
nor U13781 (N_13781,N_11622,N_11537);
or U13782 (N_13782,N_11250,N_10748);
and U13783 (N_13783,N_11389,N_9457);
nand U13784 (N_13784,N_9771,N_9910);
and U13785 (N_13785,N_9048,N_10477);
or U13786 (N_13786,N_11377,N_9984);
nor U13787 (N_13787,N_10003,N_10655);
nand U13788 (N_13788,N_10392,N_10193);
nor U13789 (N_13789,N_10848,N_11098);
xnor U13790 (N_13790,N_11568,N_11565);
nand U13791 (N_13791,N_10254,N_11920);
and U13792 (N_13792,N_10938,N_10656);
and U13793 (N_13793,N_9836,N_11201);
nor U13794 (N_13794,N_11051,N_10308);
nor U13795 (N_13795,N_9560,N_11312);
and U13796 (N_13796,N_10184,N_9960);
nand U13797 (N_13797,N_11140,N_10136);
nor U13798 (N_13798,N_10391,N_9353);
xor U13799 (N_13799,N_10019,N_9523);
nor U13800 (N_13800,N_11794,N_11442);
nor U13801 (N_13801,N_10144,N_11572);
and U13802 (N_13802,N_11964,N_11923);
nor U13803 (N_13803,N_10153,N_9380);
nand U13804 (N_13804,N_10488,N_11683);
nand U13805 (N_13805,N_9098,N_11243);
nor U13806 (N_13806,N_11764,N_10870);
nand U13807 (N_13807,N_11674,N_11379);
nand U13808 (N_13808,N_11722,N_9288);
and U13809 (N_13809,N_10681,N_10113);
nor U13810 (N_13810,N_11356,N_9995);
nand U13811 (N_13811,N_11754,N_9279);
xnor U13812 (N_13812,N_10032,N_11058);
or U13813 (N_13813,N_11248,N_10211);
nor U13814 (N_13814,N_10378,N_9286);
nor U13815 (N_13815,N_9796,N_9563);
nor U13816 (N_13816,N_10067,N_11169);
xnor U13817 (N_13817,N_11044,N_10257);
xnor U13818 (N_13818,N_11496,N_9155);
xnor U13819 (N_13819,N_9928,N_9296);
and U13820 (N_13820,N_11978,N_11968);
xnor U13821 (N_13821,N_9722,N_10375);
and U13822 (N_13822,N_9109,N_10527);
nand U13823 (N_13823,N_10650,N_11124);
xnor U13824 (N_13824,N_11056,N_10336);
nand U13825 (N_13825,N_9413,N_11658);
nor U13826 (N_13826,N_9912,N_11177);
and U13827 (N_13827,N_11792,N_11770);
or U13828 (N_13828,N_9351,N_9836);
and U13829 (N_13829,N_9422,N_9237);
and U13830 (N_13830,N_10733,N_10845);
nand U13831 (N_13831,N_10676,N_9826);
or U13832 (N_13832,N_10276,N_9165);
nand U13833 (N_13833,N_9135,N_11170);
xnor U13834 (N_13834,N_11047,N_9180);
or U13835 (N_13835,N_10741,N_11208);
or U13836 (N_13836,N_10068,N_9518);
and U13837 (N_13837,N_11492,N_11949);
nor U13838 (N_13838,N_9324,N_9589);
xor U13839 (N_13839,N_11296,N_11670);
or U13840 (N_13840,N_11534,N_11517);
or U13841 (N_13841,N_11461,N_11357);
xor U13842 (N_13842,N_10797,N_11582);
or U13843 (N_13843,N_10041,N_10790);
and U13844 (N_13844,N_10989,N_11319);
or U13845 (N_13845,N_9347,N_9906);
nand U13846 (N_13846,N_10386,N_11230);
or U13847 (N_13847,N_10832,N_11364);
nor U13848 (N_13848,N_11974,N_11450);
nand U13849 (N_13849,N_10996,N_11177);
nand U13850 (N_13850,N_9591,N_10505);
xnor U13851 (N_13851,N_11963,N_9776);
and U13852 (N_13852,N_11565,N_10972);
xnor U13853 (N_13853,N_11057,N_10841);
or U13854 (N_13854,N_11515,N_9587);
and U13855 (N_13855,N_10272,N_10265);
and U13856 (N_13856,N_10765,N_11123);
or U13857 (N_13857,N_9418,N_11983);
xor U13858 (N_13858,N_9395,N_9453);
and U13859 (N_13859,N_9771,N_9083);
nor U13860 (N_13860,N_10181,N_11502);
or U13861 (N_13861,N_10943,N_11064);
nor U13862 (N_13862,N_10407,N_10272);
nand U13863 (N_13863,N_9059,N_9585);
or U13864 (N_13864,N_9692,N_10346);
nor U13865 (N_13865,N_9160,N_9516);
and U13866 (N_13866,N_10315,N_9547);
xnor U13867 (N_13867,N_11872,N_11735);
xnor U13868 (N_13868,N_11340,N_9757);
and U13869 (N_13869,N_9066,N_11318);
nand U13870 (N_13870,N_10629,N_11412);
xnor U13871 (N_13871,N_11075,N_11770);
or U13872 (N_13872,N_10219,N_10469);
nor U13873 (N_13873,N_11408,N_11532);
xor U13874 (N_13874,N_11292,N_9773);
nand U13875 (N_13875,N_10554,N_9832);
nor U13876 (N_13876,N_11376,N_10215);
nand U13877 (N_13877,N_9069,N_11334);
nand U13878 (N_13878,N_9944,N_10522);
nor U13879 (N_13879,N_10888,N_10999);
nand U13880 (N_13880,N_10133,N_10348);
or U13881 (N_13881,N_10232,N_9211);
or U13882 (N_13882,N_11045,N_9656);
and U13883 (N_13883,N_10633,N_11043);
nor U13884 (N_13884,N_11239,N_9189);
nor U13885 (N_13885,N_11059,N_11378);
or U13886 (N_13886,N_10225,N_9509);
nor U13887 (N_13887,N_11284,N_9297);
xnor U13888 (N_13888,N_10868,N_11496);
and U13889 (N_13889,N_9632,N_11607);
nand U13890 (N_13890,N_11206,N_10494);
and U13891 (N_13891,N_10778,N_11198);
or U13892 (N_13892,N_9116,N_10372);
or U13893 (N_13893,N_11157,N_10946);
and U13894 (N_13894,N_10404,N_10189);
xor U13895 (N_13895,N_9821,N_9308);
nand U13896 (N_13896,N_10057,N_10483);
nand U13897 (N_13897,N_11684,N_11801);
nor U13898 (N_13898,N_9150,N_9575);
or U13899 (N_13899,N_11030,N_11450);
nand U13900 (N_13900,N_9393,N_11645);
xor U13901 (N_13901,N_9337,N_11768);
xnor U13902 (N_13902,N_11178,N_10902);
and U13903 (N_13903,N_10900,N_10498);
xnor U13904 (N_13904,N_9881,N_9774);
nor U13905 (N_13905,N_11021,N_11368);
or U13906 (N_13906,N_10600,N_11957);
or U13907 (N_13907,N_10817,N_9707);
or U13908 (N_13908,N_11425,N_10871);
xnor U13909 (N_13909,N_11530,N_9429);
or U13910 (N_13910,N_10386,N_10945);
nand U13911 (N_13911,N_9444,N_9946);
and U13912 (N_13912,N_10190,N_11305);
nand U13913 (N_13913,N_10292,N_10089);
nor U13914 (N_13914,N_10153,N_10310);
or U13915 (N_13915,N_11341,N_10830);
nor U13916 (N_13916,N_10777,N_9536);
nand U13917 (N_13917,N_10807,N_9242);
nand U13918 (N_13918,N_10368,N_10619);
nor U13919 (N_13919,N_9276,N_11991);
xnor U13920 (N_13920,N_10234,N_9127);
or U13921 (N_13921,N_9972,N_9743);
and U13922 (N_13922,N_10597,N_10034);
nor U13923 (N_13923,N_10298,N_9839);
xor U13924 (N_13924,N_11152,N_9726);
nand U13925 (N_13925,N_11204,N_10118);
and U13926 (N_13926,N_9256,N_9211);
or U13927 (N_13927,N_10096,N_11801);
or U13928 (N_13928,N_10347,N_10905);
or U13929 (N_13929,N_10670,N_10588);
nand U13930 (N_13930,N_11216,N_9601);
nor U13931 (N_13931,N_11874,N_11242);
nor U13932 (N_13932,N_10155,N_11038);
xnor U13933 (N_13933,N_10120,N_11233);
or U13934 (N_13934,N_9799,N_11450);
nand U13935 (N_13935,N_10410,N_11663);
nor U13936 (N_13936,N_10794,N_10923);
or U13937 (N_13937,N_9852,N_10175);
nor U13938 (N_13938,N_10999,N_9329);
or U13939 (N_13939,N_11333,N_11649);
or U13940 (N_13940,N_10222,N_9930);
nand U13941 (N_13941,N_10577,N_11199);
xor U13942 (N_13942,N_11573,N_11199);
nor U13943 (N_13943,N_10674,N_9143);
nor U13944 (N_13944,N_11766,N_9259);
nand U13945 (N_13945,N_10804,N_10240);
xor U13946 (N_13946,N_9258,N_9995);
nand U13947 (N_13947,N_11103,N_10945);
and U13948 (N_13948,N_11547,N_10855);
nor U13949 (N_13949,N_9897,N_11628);
xnor U13950 (N_13950,N_10416,N_11897);
nor U13951 (N_13951,N_9929,N_10092);
nand U13952 (N_13952,N_10644,N_11373);
and U13953 (N_13953,N_10072,N_10178);
nor U13954 (N_13954,N_9143,N_9700);
or U13955 (N_13955,N_11655,N_11226);
nand U13956 (N_13956,N_9053,N_10840);
nor U13957 (N_13957,N_9867,N_10196);
and U13958 (N_13958,N_10291,N_9245);
or U13959 (N_13959,N_11118,N_10849);
or U13960 (N_13960,N_11595,N_11705);
and U13961 (N_13961,N_11007,N_11323);
or U13962 (N_13962,N_9699,N_10671);
nand U13963 (N_13963,N_9182,N_11327);
and U13964 (N_13964,N_9894,N_11187);
nor U13965 (N_13965,N_11865,N_9610);
nor U13966 (N_13966,N_10219,N_10668);
nand U13967 (N_13967,N_10357,N_10604);
and U13968 (N_13968,N_9625,N_11083);
nor U13969 (N_13969,N_11474,N_10037);
nor U13970 (N_13970,N_9393,N_9969);
nor U13971 (N_13971,N_10999,N_11513);
or U13972 (N_13972,N_9717,N_10820);
or U13973 (N_13973,N_10399,N_11549);
nor U13974 (N_13974,N_9074,N_10986);
and U13975 (N_13975,N_11580,N_10782);
nand U13976 (N_13976,N_10795,N_11944);
nand U13977 (N_13977,N_9411,N_10787);
xnor U13978 (N_13978,N_10336,N_9725);
nand U13979 (N_13979,N_10793,N_10188);
and U13980 (N_13980,N_10277,N_9548);
nand U13981 (N_13981,N_9129,N_9560);
and U13982 (N_13982,N_10236,N_10497);
nor U13983 (N_13983,N_9491,N_9802);
nor U13984 (N_13984,N_9536,N_10673);
nand U13985 (N_13985,N_11574,N_10022);
or U13986 (N_13986,N_10361,N_9311);
and U13987 (N_13987,N_11203,N_11387);
nand U13988 (N_13988,N_11516,N_10753);
nand U13989 (N_13989,N_9810,N_11954);
nor U13990 (N_13990,N_11676,N_11974);
nor U13991 (N_13991,N_11068,N_10424);
or U13992 (N_13992,N_9897,N_10747);
nand U13993 (N_13993,N_9864,N_10692);
nor U13994 (N_13994,N_10622,N_10040);
xor U13995 (N_13995,N_9314,N_11441);
nand U13996 (N_13996,N_10301,N_9939);
nor U13997 (N_13997,N_9675,N_9084);
or U13998 (N_13998,N_10373,N_9369);
or U13999 (N_13999,N_10125,N_10123);
xor U14000 (N_14000,N_11287,N_10165);
nand U14001 (N_14001,N_11126,N_9193);
nor U14002 (N_14002,N_11863,N_11878);
or U14003 (N_14003,N_9659,N_10311);
nand U14004 (N_14004,N_10883,N_11560);
nand U14005 (N_14005,N_11983,N_10949);
xor U14006 (N_14006,N_10154,N_9428);
and U14007 (N_14007,N_11870,N_11522);
xor U14008 (N_14008,N_9704,N_11251);
xor U14009 (N_14009,N_9671,N_9169);
nor U14010 (N_14010,N_10284,N_11268);
nor U14011 (N_14011,N_9118,N_10219);
and U14012 (N_14012,N_10462,N_9543);
or U14013 (N_14013,N_11552,N_10598);
nor U14014 (N_14014,N_11769,N_11498);
and U14015 (N_14015,N_10334,N_10506);
nand U14016 (N_14016,N_10136,N_10279);
nand U14017 (N_14017,N_11159,N_11942);
xor U14018 (N_14018,N_10617,N_10772);
nor U14019 (N_14019,N_10213,N_9643);
nor U14020 (N_14020,N_11996,N_9888);
nand U14021 (N_14021,N_10714,N_11744);
and U14022 (N_14022,N_11152,N_9125);
or U14023 (N_14023,N_9381,N_9907);
and U14024 (N_14024,N_10025,N_9963);
nand U14025 (N_14025,N_11081,N_10261);
and U14026 (N_14026,N_10599,N_11503);
or U14027 (N_14027,N_11989,N_9469);
or U14028 (N_14028,N_9590,N_10638);
nand U14029 (N_14029,N_11261,N_11057);
nor U14030 (N_14030,N_9912,N_10326);
nor U14031 (N_14031,N_9303,N_9242);
nand U14032 (N_14032,N_10681,N_9691);
and U14033 (N_14033,N_11278,N_9545);
nand U14034 (N_14034,N_10533,N_9750);
nor U14035 (N_14035,N_11587,N_10833);
nand U14036 (N_14036,N_10930,N_10704);
nand U14037 (N_14037,N_11373,N_10865);
nand U14038 (N_14038,N_9220,N_11029);
and U14039 (N_14039,N_10116,N_9620);
nand U14040 (N_14040,N_10326,N_9529);
nand U14041 (N_14041,N_10900,N_10207);
nor U14042 (N_14042,N_11859,N_10244);
or U14043 (N_14043,N_9115,N_10563);
xor U14044 (N_14044,N_10068,N_11951);
xor U14045 (N_14045,N_10963,N_11630);
or U14046 (N_14046,N_11184,N_9798);
nor U14047 (N_14047,N_11865,N_11344);
nand U14048 (N_14048,N_9589,N_11798);
or U14049 (N_14049,N_11753,N_9318);
nor U14050 (N_14050,N_11846,N_9577);
or U14051 (N_14051,N_9741,N_9427);
or U14052 (N_14052,N_11199,N_10579);
and U14053 (N_14053,N_11380,N_11340);
nor U14054 (N_14054,N_11557,N_10845);
nor U14055 (N_14055,N_9236,N_11004);
nand U14056 (N_14056,N_11171,N_11631);
nand U14057 (N_14057,N_9593,N_9526);
nand U14058 (N_14058,N_10067,N_10533);
or U14059 (N_14059,N_9695,N_9360);
xor U14060 (N_14060,N_10760,N_11075);
xor U14061 (N_14061,N_11235,N_9484);
nand U14062 (N_14062,N_11954,N_9181);
xnor U14063 (N_14063,N_11439,N_9094);
or U14064 (N_14064,N_9573,N_11199);
xor U14065 (N_14065,N_9291,N_9692);
nand U14066 (N_14066,N_10912,N_10769);
nand U14067 (N_14067,N_9770,N_10614);
and U14068 (N_14068,N_10389,N_10682);
nand U14069 (N_14069,N_9214,N_11495);
or U14070 (N_14070,N_9115,N_9809);
nor U14071 (N_14071,N_10375,N_10707);
and U14072 (N_14072,N_10886,N_11244);
nand U14073 (N_14073,N_9717,N_10850);
nor U14074 (N_14074,N_9330,N_10746);
xor U14075 (N_14075,N_10426,N_11332);
or U14076 (N_14076,N_11395,N_11292);
xor U14077 (N_14077,N_10585,N_10647);
and U14078 (N_14078,N_10628,N_9912);
and U14079 (N_14079,N_11028,N_10497);
nand U14080 (N_14080,N_11542,N_10856);
xnor U14081 (N_14081,N_9920,N_9505);
nor U14082 (N_14082,N_9907,N_9875);
nor U14083 (N_14083,N_9603,N_9938);
nand U14084 (N_14084,N_11987,N_11532);
nor U14085 (N_14085,N_11875,N_10270);
and U14086 (N_14086,N_11420,N_10781);
nor U14087 (N_14087,N_9176,N_9063);
and U14088 (N_14088,N_9913,N_10755);
or U14089 (N_14089,N_9533,N_9513);
and U14090 (N_14090,N_10456,N_9878);
xnor U14091 (N_14091,N_11628,N_9441);
xor U14092 (N_14092,N_10152,N_11838);
nand U14093 (N_14093,N_11062,N_10120);
nand U14094 (N_14094,N_10816,N_10062);
xor U14095 (N_14095,N_9414,N_10696);
xor U14096 (N_14096,N_9469,N_10889);
xor U14097 (N_14097,N_10809,N_11968);
or U14098 (N_14098,N_11530,N_10319);
and U14099 (N_14099,N_9735,N_10229);
and U14100 (N_14100,N_10227,N_9638);
nand U14101 (N_14101,N_10305,N_10125);
or U14102 (N_14102,N_9639,N_9704);
xnor U14103 (N_14103,N_10818,N_10100);
or U14104 (N_14104,N_11887,N_9093);
xnor U14105 (N_14105,N_10068,N_10454);
or U14106 (N_14106,N_10566,N_10946);
xnor U14107 (N_14107,N_11545,N_11955);
and U14108 (N_14108,N_9165,N_11720);
nand U14109 (N_14109,N_10928,N_10242);
nand U14110 (N_14110,N_11750,N_9341);
nand U14111 (N_14111,N_11908,N_11182);
or U14112 (N_14112,N_10549,N_11547);
and U14113 (N_14113,N_11680,N_11145);
and U14114 (N_14114,N_11025,N_10104);
xor U14115 (N_14115,N_11940,N_10190);
or U14116 (N_14116,N_10823,N_10984);
nor U14117 (N_14117,N_9564,N_9226);
or U14118 (N_14118,N_10343,N_9210);
nor U14119 (N_14119,N_10973,N_9299);
or U14120 (N_14120,N_10512,N_11547);
or U14121 (N_14121,N_9180,N_11579);
nor U14122 (N_14122,N_9899,N_11090);
nor U14123 (N_14123,N_11223,N_9813);
and U14124 (N_14124,N_10951,N_11415);
or U14125 (N_14125,N_9605,N_11146);
nor U14126 (N_14126,N_9870,N_9317);
nand U14127 (N_14127,N_11683,N_11581);
nand U14128 (N_14128,N_9808,N_11802);
or U14129 (N_14129,N_9347,N_10600);
or U14130 (N_14130,N_11412,N_11735);
nand U14131 (N_14131,N_10840,N_10237);
nand U14132 (N_14132,N_10559,N_9030);
nand U14133 (N_14133,N_11961,N_11928);
nand U14134 (N_14134,N_9420,N_9180);
nor U14135 (N_14135,N_10132,N_11165);
nand U14136 (N_14136,N_10786,N_9836);
nand U14137 (N_14137,N_10321,N_10716);
or U14138 (N_14138,N_11185,N_9518);
nor U14139 (N_14139,N_11365,N_11801);
and U14140 (N_14140,N_9016,N_11883);
and U14141 (N_14141,N_11039,N_9420);
nand U14142 (N_14142,N_10783,N_9503);
nand U14143 (N_14143,N_11718,N_9382);
and U14144 (N_14144,N_10566,N_10320);
and U14145 (N_14145,N_11637,N_10165);
or U14146 (N_14146,N_11554,N_10966);
nand U14147 (N_14147,N_9117,N_11950);
xor U14148 (N_14148,N_10998,N_9148);
nor U14149 (N_14149,N_9113,N_10543);
nand U14150 (N_14150,N_11466,N_10069);
nor U14151 (N_14151,N_10663,N_11739);
or U14152 (N_14152,N_11296,N_11742);
and U14153 (N_14153,N_10480,N_11598);
or U14154 (N_14154,N_9615,N_10528);
nand U14155 (N_14155,N_9870,N_9408);
and U14156 (N_14156,N_10005,N_9879);
or U14157 (N_14157,N_11466,N_9786);
nand U14158 (N_14158,N_10631,N_10062);
nor U14159 (N_14159,N_11540,N_11103);
xor U14160 (N_14160,N_10599,N_10561);
nand U14161 (N_14161,N_11566,N_10789);
nor U14162 (N_14162,N_11181,N_9414);
or U14163 (N_14163,N_11584,N_9718);
and U14164 (N_14164,N_10813,N_9770);
xor U14165 (N_14165,N_9409,N_9746);
or U14166 (N_14166,N_9835,N_11181);
or U14167 (N_14167,N_9747,N_10258);
nand U14168 (N_14168,N_10090,N_9902);
xnor U14169 (N_14169,N_9058,N_10588);
nand U14170 (N_14170,N_11106,N_11208);
nand U14171 (N_14171,N_10747,N_10814);
nor U14172 (N_14172,N_9489,N_11151);
or U14173 (N_14173,N_11399,N_9665);
nand U14174 (N_14174,N_11492,N_10360);
nor U14175 (N_14175,N_10669,N_10152);
nor U14176 (N_14176,N_11900,N_10411);
nor U14177 (N_14177,N_11676,N_9500);
and U14178 (N_14178,N_10880,N_11017);
and U14179 (N_14179,N_11024,N_10450);
xnor U14180 (N_14180,N_11838,N_10055);
nand U14181 (N_14181,N_9980,N_9936);
nand U14182 (N_14182,N_9503,N_10167);
nor U14183 (N_14183,N_10527,N_10119);
nor U14184 (N_14184,N_11909,N_11448);
or U14185 (N_14185,N_10157,N_11842);
nor U14186 (N_14186,N_11384,N_11358);
and U14187 (N_14187,N_9618,N_11864);
and U14188 (N_14188,N_9195,N_10990);
or U14189 (N_14189,N_11027,N_11077);
and U14190 (N_14190,N_10070,N_10328);
nand U14191 (N_14191,N_10277,N_9387);
nand U14192 (N_14192,N_11941,N_9142);
xnor U14193 (N_14193,N_11089,N_10177);
nand U14194 (N_14194,N_10756,N_11320);
and U14195 (N_14195,N_10828,N_11353);
xor U14196 (N_14196,N_10619,N_11952);
nand U14197 (N_14197,N_11825,N_10013);
and U14198 (N_14198,N_10843,N_10445);
nor U14199 (N_14199,N_11959,N_9027);
or U14200 (N_14200,N_10325,N_9200);
xor U14201 (N_14201,N_11898,N_11307);
xor U14202 (N_14202,N_10156,N_11796);
nand U14203 (N_14203,N_10788,N_10603);
xor U14204 (N_14204,N_9351,N_9869);
and U14205 (N_14205,N_10081,N_11356);
or U14206 (N_14206,N_11428,N_11499);
or U14207 (N_14207,N_9131,N_11386);
nor U14208 (N_14208,N_10817,N_9727);
and U14209 (N_14209,N_11361,N_11128);
or U14210 (N_14210,N_10434,N_9730);
xor U14211 (N_14211,N_11585,N_11222);
nand U14212 (N_14212,N_11790,N_11956);
or U14213 (N_14213,N_10610,N_10665);
nand U14214 (N_14214,N_11683,N_11030);
or U14215 (N_14215,N_9923,N_11581);
xnor U14216 (N_14216,N_10817,N_11459);
or U14217 (N_14217,N_10416,N_10606);
or U14218 (N_14218,N_10167,N_9932);
or U14219 (N_14219,N_9526,N_11470);
nand U14220 (N_14220,N_9921,N_9740);
and U14221 (N_14221,N_10312,N_9897);
and U14222 (N_14222,N_9024,N_11171);
nand U14223 (N_14223,N_9466,N_11901);
and U14224 (N_14224,N_9550,N_11743);
nand U14225 (N_14225,N_9264,N_11583);
and U14226 (N_14226,N_9491,N_11596);
nand U14227 (N_14227,N_11738,N_11846);
xnor U14228 (N_14228,N_9741,N_9190);
or U14229 (N_14229,N_9787,N_11914);
nand U14230 (N_14230,N_9128,N_9301);
or U14231 (N_14231,N_9556,N_10003);
nand U14232 (N_14232,N_11635,N_10286);
and U14233 (N_14233,N_9925,N_9961);
nand U14234 (N_14234,N_9565,N_10486);
nand U14235 (N_14235,N_9875,N_10015);
nor U14236 (N_14236,N_11121,N_9452);
nor U14237 (N_14237,N_9230,N_9827);
or U14238 (N_14238,N_11517,N_11342);
xnor U14239 (N_14239,N_11348,N_10628);
or U14240 (N_14240,N_9707,N_9173);
and U14241 (N_14241,N_9408,N_10986);
xor U14242 (N_14242,N_9080,N_10132);
and U14243 (N_14243,N_9972,N_9756);
or U14244 (N_14244,N_9029,N_9415);
nor U14245 (N_14245,N_10645,N_9040);
or U14246 (N_14246,N_10244,N_11083);
nor U14247 (N_14247,N_11729,N_11259);
or U14248 (N_14248,N_11016,N_9403);
and U14249 (N_14249,N_11511,N_10770);
nand U14250 (N_14250,N_11312,N_9349);
or U14251 (N_14251,N_9280,N_9639);
nand U14252 (N_14252,N_9874,N_9259);
xnor U14253 (N_14253,N_9806,N_10635);
or U14254 (N_14254,N_9675,N_10621);
nor U14255 (N_14255,N_9215,N_11866);
nand U14256 (N_14256,N_10665,N_9952);
or U14257 (N_14257,N_11956,N_10335);
and U14258 (N_14258,N_10608,N_11956);
nor U14259 (N_14259,N_10128,N_10226);
and U14260 (N_14260,N_11267,N_10590);
and U14261 (N_14261,N_10846,N_11233);
and U14262 (N_14262,N_9304,N_10608);
nand U14263 (N_14263,N_10930,N_9471);
nor U14264 (N_14264,N_11309,N_11602);
nor U14265 (N_14265,N_9820,N_9183);
and U14266 (N_14266,N_11086,N_11931);
nor U14267 (N_14267,N_9064,N_10295);
nor U14268 (N_14268,N_11579,N_9768);
or U14269 (N_14269,N_11688,N_10920);
nor U14270 (N_14270,N_9688,N_11838);
nand U14271 (N_14271,N_10519,N_9455);
nor U14272 (N_14272,N_11340,N_10423);
nand U14273 (N_14273,N_10498,N_11670);
nor U14274 (N_14274,N_11620,N_11901);
or U14275 (N_14275,N_11767,N_9064);
nand U14276 (N_14276,N_9980,N_11614);
nor U14277 (N_14277,N_11807,N_9947);
nor U14278 (N_14278,N_9457,N_10250);
and U14279 (N_14279,N_9164,N_10375);
nand U14280 (N_14280,N_10419,N_10024);
nor U14281 (N_14281,N_11802,N_9654);
or U14282 (N_14282,N_9677,N_9263);
xnor U14283 (N_14283,N_11182,N_9071);
and U14284 (N_14284,N_9841,N_9101);
nand U14285 (N_14285,N_11881,N_11675);
and U14286 (N_14286,N_9244,N_10458);
nor U14287 (N_14287,N_11828,N_11027);
and U14288 (N_14288,N_9149,N_9240);
nand U14289 (N_14289,N_10585,N_9771);
nor U14290 (N_14290,N_9544,N_10328);
or U14291 (N_14291,N_10364,N_11897);
or U14292 (N_14292,N_11218,N_9309);
nor U14293 (N_14293,N_11696,N_10126);
and U14294 (N_14294,N_9682,N_11333);
nand U14295 (N_14295,N_9880,N_10954);
xnor U14296 (N_14296,N_9834,N_9713);
nor U14297 (N_14297,N_9625,N_11568);
nand U14298 (N_14298,N_11747,N_11824);
and U14299 (N_14299,N_9582,N_10072);
nor U14300 (N_14300,N_9480,N_11064);
nor U14301 (N_14301,N_9410,N_11967);
or U14302 (N_14302,N_11270,N_9549);
nor U14303 (N_14303,N_11118,N_11812);
or U14304 (N_14304,N_11912,N_11981);
nand U14305 (N_14305,N_9847,N_9883);
nand U14306 (N_14306,N_9439,N_9539);
and U14307 (N_14307,N_10667,N_11167);
and U14308 (N_14308,N_10700,N_9680);
nor U14309 (N_14309,N_9036,N_10298);
or U14310 (N_14310,N_11721,N_9808);
nor U14311 (N_14311,N_11803,N_9274);
or U14312 (N_14312,N_10896,N_11831);
xor U14313 (N_14313,N_9423,N_10963);
nor U14314 (N_14314,N_11688,N_11156);
xnor U14315 (N_14315,N_10619,N_11476);
xnor U14316 (N_14316,N_10803,N_10384);
or U14317 (N_14317,N_10082,N_10708);
nor U14318 (N_14318,N_9146,N_10861);
nor U14319 (N_14319,N_9860,N_9841);
nor U14320 (N_14320,N_11381,N_11564);
nand U14321 (N_14321,N_10982,N_11012);
xnor U14322 (N_14322,N_10459,N_11748);
or U14323 (N_14323,N_11751,N_11201);
and U14324 (N_14324,N_9126,N_10670);
nand U14325 (N_14325,N_10088,N_9446);
nand U14326 (N_14326,N_10959,N_11361);
and U14327 (N_14327,N_10032,N_9889);
nand U14328 (N_14328,N_9099,N_11977);
and U14329 (N_14329,N_9079,N_10686);
or U14330 (N_14330,N_9462,N_9553);
nor U14331 (N_14331,N_9724,N_11686);
or U14332 (N_14332,N_10398,N_11686);
nand U14333 (N_14333,N_10284,N_11415);
and U14334 (N_14334,N_11249,N_11184);
nor U14335 (N_14335,N_9901,N_10177);
nand U14336 (N_14336,N_9224,N_10883);
nor U14337 (N_14337,N_10628,N_10921);
nand U14338 (N_14338,N_9889,N_10157);
and U14339 (N_14339,N_9665,N_9888);
and U14340 (N_14340,N_10909,N_9684);
nand U14341 (N_14341,N_9365,N_11453);
and U14342 (N_14342,N_10401,N_9527);
and U14343 (N_14343,N_10868,N_9507);
and U14344 (N_14344,N_11216,N_9532);
nor U14345 (N_14345,N_9617,N_11389);
or U14346 (N_14346,N_10090,N_9666);
nor U14347 (N_14347,N_11565,N_11804);
and U14348 (N_14348,N_11400,N_11828);
nor U14349 (N_14349,N_10066,N_9119);
and U14350 (N_14350,N_9228,N_11164);
or U14351 (N_14351,N_9399,N_9186);
and U14352 (N_14352,N_9894,N_11589);
nor U14353 (N_14353,N_10077,N_9843);
nor U14354 (N_14354,N_9534,N_11286);
or U14355 (N_14355,N_9368,N_10938);
or U14356 (N_14356,N_11577,N_11755);
or U14357 (N_14357,N_10493,N_11255);
nand U14358 (N_14358,N_11284,N_11088);
or U14359 (N_14359,N_11041,N_11416);
nor U14360 (N_14360,N_11956,N_10892);
xnor U14361 (N_14361,N_10728,N_9551);
and U14362 (N_14362,N_11839,N_10768);
or U14363 (N_14363,N_11719,N_10924);
xnor U14364 (N_14364,N_11056,N_11222);
nand U14365 (N_14365,N_10228,N_11926);
nor U14366 (N_14366,N_9135,N_10938);
nor U14367 (N_14367,N_9817,N_10021);
and U14368 (N_14368,N_9837,N_10705);
and U14369 (N_14369,N_9741,N_9161);
xnor U14370 (N_14370,N_11145,N_11932);
and U14371 (N_14371,N_10336,N_9143);
and U14372 (N_14372,N_10646,N_9305);
nor U14373 (N_14373,N_10827,N_9751);
and U14374 (N_14374,N_9217,N_9964);
xnor U14375 (N_14375,N_10678,N_11715);
and U14376 (N_14376,N_9660,N_9818);
xor U14377 (N_14377,N_11811,N_9668);
nor U14378 (N_14378,N_10848,N_10491);
or U14379 (N_14379,N_10499,N_11026);
xor U14380 (N_14380,N_11879,N_11502);
or U14381 (N_14381,N_11354,N_11084);
nor U14382 (N_14382,N_11553,N_11745);
or U14383 (N_14383,N_10366,N_9063);
and U14384 (N_14384,N_9252,N_10040);
and U14385 (N_14385,N_10315,N_9954);
or U14386 (N_14386,N_11794,N_11650);
xor U14387 (N_14387,N_9562,N_11625);
nand U14388 (N_14388,N_11116,N_9010);
xnor U14389 (N_14389,N_10379,N_10969);
nor U14390 (N_14390,N_9035,N_10681);
nor U14391 (N_14391,N_9894,N_9483);
nor U14392 (N_14392,N_10784,N_9737);
nand U14393 (N_14393,N_9019,N_11831);
nor U14394 (N_14394,N_9452,N_9561);
nand U14395 (N_14395,N_11186,N_10632);
nor U14396 (N_14396,N_9523,N_11934);
and U14397 (N_14397,N_9791,N_11728);
nor U14398 (N_14398,N_10163,N_10205);
and U14399 (N_14399,N_11817,N_9181);
nor U14400 (N_14400,N_10885,N_11366);
nand U14401 (N_14401,N_10888,N_11184);
nand U14402 (N_14402,N_11701,N_11938);
nor U14403 (N_14403,N_10179,N_9977);
xnor U14404 (N_14404,N_11993,N_11591);
and U14405 (N_14405,N_11424,N_11546);
and U14406 (N_14406,N_11219,N_11052);
nor U14407 (N_14407,N_10298,N_10183);
nand U14408 (N_14408,N_10595,N_11218);
nand U14409 (N_14409,N_11052,N_10559);
nand U14410 (N_14410,N_9988,N_9514);
or U14411 (N_14411,N_10710,N_10016);
xnor U14412 (N_14412,N_10488,N_9984);
nor U14413 (N_14413,N_10521,N_10248);
nand U14414 (N_14414,N_11931,N_9618);
or U14415 (N_14415,N_9684,N_10033);
nand U14416 (N_14416,N_9250,N_11993);
xor U14417 (N_14417,N_11298,N_11453);
or U14418 (N_14418,N_11578,N_11667);
nand U14419 (N_14419,N_10338,N_10394);
and U14420 (N_14420,N_10591,N_9242);
nand U14421 (N_14421,N_10946,N_9471);
and U14422 (N_14422,N_11354,N_10635);
and U14423 (N_14423,N_11976,N_10131);
nor U14424 (N_14424,N_10129,N_11523);
nand U14425 (N_14425,N_11550,N_10310);
nor U14426 (N_14426,N_11520,N_10903);
nor U14427 (N_14427,N_10909,N_9300);
or U14428 (N_14428,N_10487,N_11207);
nand U14429 (N_14429,N_10525,N_11251);
and U14430 (N_14430,N_9623,N_9202);
xor U14431 (N_14431,N_11455,N_11493);
and U14432 (N_14432,N_9666,N_10636);
and U14433 (N_14433,N_9476,N_10640);
or U14434 (N_14434,N_10754,N_11933);
nand U14435 (N_14435,N_9405,N_9064);
or U14436 (N_14436,N_9216,N_10863);
nor U14437 (N_14437,N_11585,N_11217);
and U14438 (N_14438,N_10628,N_9550);
nand U14439 (N_14439,N_11671,N_10872);
nor U14440 (N_14440,N_11241,N_10870);
and U14441 (N_14441,N_10239,N_11583);
nand U14442 (N_14442,N_9185,N_11173);
or U14443 (N_14443,N_11344,N_11683);
and U14444 (N_14444,N_10145,N_9898);
nand U14445 (N_14445,N_10687,N_11191);
nor U14446 (N_14446,N_11178,N_11937);
and U14447 (N_14447,N_11282,N_11515);
nor U14448 (N_14448,N_9488,N_10540);
and U14449 (N_14449,N_11267,N_11061);
and U14450 (N_14450,N_10665,N_11197);
and U14451 (N_14451,N_10524,N_9182);
nor U14452 (N_14452,N_9791,N_11650);
nor U14453 (N_14453,N_9049,N_11384);
nand U14454 (N_14454,N_10884,N_11195);
nor U14455 (N_14455,N_11586,N_11304);
nand U14456 (N_14456,N_9801,N_10721);
nor U14457 (N_14457,N_9300,N_10839);
xnor U14458 (N_14458,N_10121,N_11219);
or U14459 (N_14459,N_11923,N_9226);
nor U14460 (N_14460,N_9983,N_9086);
and U14461 (N_14461,N_9322,N_11925);
or U14462 (N_14462,N_9920,N_11802);
or U14463 (N_14463,N_10717,N_10439);
nor U14464 (N_14464,N_10940,N_10657);
nand U14465 (N_14465,N_11589,N_9165);
nand U14466 (N_14466,N_10997,N_10841);
or U14467 (N_14467,N_11060,N_11865);
and U14468 (N_14468,N_9154,N_9858);
nor U14469 (N_14469,N_9277,N_10631);
and U14470 (N_14470,N_9380,N_9962);
and U14471 (N_14471,N_10742,N_11086);
or U14472 (N_14472,N_11653,N_9718);
or U14473 (N_14473,N_10444,N_9130);
or U14474 (N_14474,N_10632,N_10473);
and U14475 (N_14475,N_10288,N_10850);
nor U14476 (N_14476,N_11737,N_9384);
xnor U14477 (N_14477,N_11276,N_11185);
nand U14478 (N_14478,N_11932,N_9636);
xnor U14479 (N_14479,N_11526,N_10848);
nor U14480 (N_14480,N_10997,N_10503);
xnor U14481 (N_14481,N_9992,N_9335);
nand U14482 (N_14482,N_9214,N_10924);
and U14483 (N_14483,N_10603,N_10224);
and U14484 (N_14484,N_11704,N_10820);
nor U14485 (N_14485,N_11963,N_9917);
and U14486 (N_14486,N_9280,N_11083);
or U14487 (N_14487,N_9579,N_11199);
xor U14488 (N_14488,N_10096,N_10218);
nand U14489 (N_14489,N_11399,N_10420);
or U14490 (N_14490,N_9943,N_11846);
nand U14491 (N_14491,N_11466,N_9294);
or U14492 (N_14492,N_9266,N_10850);
and U14493 (N_14493,N_11960,N_11278);
nor U14494 (N_14494,N_11895,N_11257);
and U14495 (N_14495,N_10279,N_10099);
or U14496 (N_14496,N_9403,N_11266);
and U14497 (N_14497,N_9007,N_9336);
xnor U14498 (N_14498,N_10820,N_11846);
and U14499 (N_14499,N_11578,N_9851);
and U14500 (N_14500,N_10881,N_11525);
nand U14501 (N_14501,N_9293,N_10190);
or U14502 (N_14502,N_11568,N_11131);
and U14503 (N_14503,N_9008,N_9310);
nor U14504 (N_14504,N_9175,N_11579);
nor U14505 (N_14505,N_9204,N_11534);
or U14506 (N_14506,N_11864,N_10281);
and U14507 (N_14507,N_9503,N_11566);
nor U14508 (N_14508,N_10928,N_11348);
nand U14509 (N_14509,N_9368,N_9657);
nand U14510 (N_14510,N_9314,N_11225);
xnor U14511 (N_14511,N_9156,N_11767);
nor U14512 (N_14512,N_9187,N_9759);
and U14513 (N_14513,N_10436,N_11071);
nor U14514 (N_14514,N_10491,N_10306);
nand U14515 (N_14515,N_10686,N_11313);
or U14516 (N_14516,N_9948,N_9121);
nand U14517 (N_14517,N_10514,N_10250);
and U14518 (N_14518,N_9774,N_11705);
nor U14519 (N_14519,N_11936,N_9458);
nand U14520 (N_14520,N_11861,N_9855);
or U14521 (N_14521,N_9057,N_10513);
nand U14522 (N_14522,N_11412,N_9139);
nor U14523 (N_14523,N_11445,N_11648);
and U14524 (N_14524,N_10590,N_11819);
or U14525 (N_14525,N_9195,N_9923);
or U14526 (N_14526,N_11421,N_11251);
or U14527 (N_14527,N_11487,N_10705);
or U14528 (N_14528,N_11731,N_10633);
nand U14529 (N_14529,N_10045,N_11080);
and U14530 (N_14530,N_11480,N_9215);
or U14531 (N_14531,N_11776,N_11322);
and U14532 (N_14532,N_11883,N_10148);
or U14533 (N_14533,N_11580,N_10982);
nand U14534 (N_14534,N_11520,N_11402);
nor U14535 (N_14535,N_9990,N_10066);
or U14536 (N_14536,N_9858,N_9980);
and U14537 (N_14537,N_10132,N_11579);
or U14538 (N_14538,N_10197,N_11888);
or U14539 (N_14539,N_11662,N_10868);
nor U14540 (N_14540,N_11187,N_9504);
nand U14541 (N_14541,N_10271,N_9490);
or U14542 (N_14542,N_11336,N_9485);
nand U14543 (N_14543,N_9404,N_9422);
and U14544 (N_14544,N_11088,N_10612);
nand U14545 (N_14545,N_9550,N_11289);
nand U14546 (N_14546,N_11267,N_9036);
nor U14547 (N_14547,N_9902,N_11010);
nand U14548 (N_14548,N_11154,N_9495);
and U14549 (N_14549,N_9149,N_9231);
nand U14550 (N_14550,N_10033,N_9831);
or U14551 (N_14551,N_11219,N_11026);
or U14552 (N_14552,N_11346,N_10633);
or U14553 (N_14553,N_9059,N_9129);
nand U14554 (N_14554,N_9952,N_11443);
and U14555 (N_14555,N_10256,N_10671);
nand U14556 (N_14556,N_9078,N_9860);
and U14557 (N_14557,N_10684,N_11895);
or U14558 (N_14558,N_11802,N_10007);
nor U14559 (N_14559,N_10461,N_9792);
xor U14560 (N_14560,N_9205,N_11266);
nand U14561 (N_14561,N_9255,N_11427);
nand U14562 (N_14562,N_11240,N_10586);
nand U14563 (N_14563,N_10722,N_10488);
nand U14564 (N_14564,N_11470,N_9519);
nand U14565 (N_14565,N_11362,N_11503);
nor U14566 (N_14566,N_9416,N_10254);
and U14567 (N_14567,N_11275,N_11990);
and U14568 (N_14568,N_9207,N_11408);
nor U14569 (N_14569,N_10844,N_11044);
nor U14570 (N_14570,N_9217,N_11356);
and U14571 (N_14571,N_10298,N_9177);
nand U14572 (N_14572,N_9248,N_10811);
or U14573 (N_14573,N_9988,N_11127);
and U14574 (N_14574,N_11836,N_11870);
nor U14575 (N_14575,N_9529,N_9477);
or U14576 (N_14576,N_11442,N_9310);
nand U14577 (N_14577,N_10151,N_11074);
and U14578 (N_14578,N_11748,N_11293);
nor U14579 (N_14579,N_10432,N_11843);
and U14580 (N_14580,N_10648,N_9424);
or U14581 (N_14581,N_9280,N_11557);
nand U14582 (N_14582,N_10701,N_11120);
nor U14583 (N_14583,N_9999,N_11854);
nand U14584 (N_14584,N_9738,N_10155);
or U14585 (N_14585,N_11970,N_9688);
nor U14586 (N_14586,N_9841,N_9969);
xor U14587 (N_14587,N_11865,N_11799);
or U14588 (N_14588,N_9632,N_9991);
or U14589 (N_14589,N_10307,N_9788);
and U14590 (N_14590,N_9730,N_11474);
nor U14591 (N_14591,N_10246,N_10968);
xnor U14592 (N_14592,N_10990,N_11172);
nand U14593 (N_14593,N_10218,N_10877);
nor U14594 (N_14594,N_11697,N_11402);
nor U14595 (N_14595,N_10944,N_10600);
nor U14596 (N_14596,N_10376,N_11493);
and U14597 (N_14597,N_11357,N_10927);
and U14598 (N_14598,N_10031,N_9404);
nor U14599 (N_14599,N_11403,N_10189);
nand U14600 (N_14600,N_11310,N_11003);
or U14601 (N_14601,N_9710,N_11723);
xnor U14602 (N_14602,N_9254,N_11735);
xnor U14603 (N_14603,N_10095,N_9318);
nor U14604 (N_14604,N_9378,N_10197);
or U14605 (N_14605,N_10463,N_10906);
nand U14606 (N_14606,N_9656,N_11052);
nor U14607 (N_14607,N_9898,N_10609);
or U14608 (N_14608,N_9194,N_10967);
or U14609 (N_14609,N_10797,N_11871);
and U14610 (N_14610,N_9392,N_10099);
nand U14611 (N_14611,N_9102,N_11092);
nand U14612 (N_14612,N_9533,N_10222);
nand U14613 (N_14613,N_10029,N_9901);
and U14614 (N_14614,N_11282,N_10336);
nor U14615 (N_14615,N_11955,N_9989);
nand U14616 (N_14616,N_10586,N_10554);
or U14617 (N_14617,N_9969,N_10066);
or U14618 (N_14618,N_9308,N_9917);
and U14619 (N_14619,N_9216,N_9615);
nor U14620 (N_14620,N_10106,N_9612);
or U14621 (N_14621,N_11662,N_10651);
and U14622 (N_14622,N_9479,N_11827);
nor U14623 (N_14623,N_11190,N_10828);
and U14624 (N_14624,N_11908,N_9963);
xnor U14625 (N_14625,N_11382,N_11440);
nand U14626 (N_14626,N_11540,N_10079);
nor U14627 (N_14627,N_9495,N_10698);
and U14628 (N_14628,N_11280,N_11128);
xnor U14629 (N_14629,N_11186,N_9689);
or U14630 (N_14630,N_10789,N_11588);
nand U14631 (N_14631,N_10195,N_10953);
nand U14632 (N_14632,N_11266,N_11961);
nand U14633 (N_14633,N_11393,N_9538);
and U14634 (N_14634,N_9390,N_11047);
and U14635 (N_14635,N_11051,N_10190);
nand U14636 (N_14636,N_11787,N_10355);
xor U14637 (N_14637,N_9777,N_9667);
and U14638 (N_14638,N_10605,N_9934);
or U14639 (N_14639,N_9940,N_11030);
nor U14640 (N_14640,N_9767,N_11642);
nor U14641 (N_14641,N_10350,N_9415);
nor U14642 (N_14642,N_9380,N_9703);
nor U14643 (N_14643,N_10969,N_9762);
nand U14644 (N_14644,N_11537,N_11169);
xor U14645 (N_14645,N_10016,N_10443);
nand U14646 (N_14646,N_9750,N_9399);
nor U14647 (N_14647,N_10115,N_11026);
and U14648 (N_14648,N_10621,N_10037);
and U14649 (N_14649,N_9296,N_10300);
nor U14650 (N_14650,N_11343,N_9165);
nor U14651 (N_14651,N_10460,N_9020);
nor U14652 (N_14652,N_10759,N_10366);
or U14653 (N_14653,N_9143,N_9997);
or U14654 (N_14654,N_11762,N_10316);
nand U14655 (N_14655,N_10753,N_11313);
and U14656 (N_14656,N_11894,N_11900);
nand U14657 (N_14657,N_11092,N_9362);
or U14658 (N_14658,N_11129,N_9861);
nor U14659 (N_14659,N_10653,N_9645);
and U14660 (N_14660,N_10958,N_11816);
nand U14661 (N_14661,N_9426,N_9981);
nand U14662 (N_14662,N_11533,N_11280);
or U14663 (N_14663,N_10900,N_11012);
nor U14664 (N_14664,N_10028,N_11752);
xor U14665 (N_14665,N_9423,N_10795);
nand U14666 (N_14666,N_9262,N_10996);
nor U14667 (N_14667,N_10546,N_9139);
nor U14668 (N_14668,N_11881,N_11577);
or U14669 (N_14669,N_11503,N_9943);
xnor U14670 (N_14670,N_10852,N_11653);
nor U14671 (N_14671,N_11959,N_11372);
xor U14672 (N_14672,N_10032,N_9391);
nor U14673 (N_14673,N_11272,N_11166);
xnor U14674 (N_14674,N_10448,N_11983);
nor U14675 (N_14675,N_10389,N_11458);
xor U14676 (N_14676,N_10632,N_11788);
xnor U14677 (N_14677,N_11627,N_11030);
nor U14678 (N_14678,N_11784,N_10196);
or U14679 (N_14679,N_11182,N_10296);
nand U14680 (N_14680,N_10554,N_11702);
nand U14681 (N_14681,N_9401,N_11856);
nand U14682 (N_14682,N_10971,N_9663);
nand U14683 (N_14683,N_11444,N_10159);
and U14684 (N_14684,N_11974,N_11181);
xnor U14685 (N_14685,N_10763,N_9430);
or U14686 (N_14686,N_11668,N_9773);
nand U14687 (N_14687,N_9719,N_10686);
and U14688 (N_14688,N_9348,N_9134);
nand U14689 (N_14689,N_9980,N_11058);
or U14690 (N_14690,N_10156,N_9026);
nor U14691 (N_14691,N_11708,N_11121);
nor U14692 (N_14692,N_11161,N_9597);
or U14693 (N_14693,N_9344,N_10763);
and U14694 (N_14694,N_10768,N_10340);
nor U14695 (N_14695,N_9967,N_11991);
nand U14696 (N_14696,N_9775,N_10181);
nor U14697 (N_14697,N_11626,N_11289);
or U14698 (N_14698,N_11882,N_10784);
and U14699 (N_14699,N_11630,N_10581);
xor U14700 (N_14700,N_9947,N_9871);
and U14701 (N_14701,N_10854,N_10556);
and U14702 (N_14702,N_9890,N_9461);
or U14703 (N_14703,N_9665,N_9621);
nand U14704 (N_14704,N_10348,N_10555);
and U14705 (N_14705,N_11950,N_9945);
nand U14706 (N_14706,N_10755,N_10631);
nand U14707 (N_14707,N_10367,N_11812);
or U14708 (N_14708,N_10800,N_9411);
nor U14709 (N_14709,N_11174,N_9539);
or U14710 (N_14710,N_11447,N_9912);
xnor U14711 (N_14711,N_10892,N_11641);
nor U14712 (N_14712,N_11636,N_10526);
xor U14713 (N_14713,N_9580,N_10770);
or U14714 (N_14714,N_11455,N_11915);
or U14715 (N_14715,N_11524,N_9071);
nand U14716 (N_14716,N_10824,N_11955);
nand U14717 (N_14717,N_10675,N_11069);
nor U14718 (N_14718,N_10591,N_10605);
nor U14719 (N_14719,N_11964,N_11780);
nor U14720 (N_14720,N_9916,N_9966);
and U14721 (N_14721,N_9939,N_10416);
nor U14722 (N_14722,N_9591,N_9202);
or U14723 (N_14723,N_11809,N_11255);
nor U14724 (N_14724,N_10749,N_9198);
or U14725 (N_14725,N_11655,N_10231);
nand U14726 (N_14726,N_11721,N_9078);
xnor U14727 (N_14727,N_10033,N_11864);
nand U14728 (N_14728,N_11359,N_9621);
xnor U14729 (N_14729,N_10726,N_9978);
or U14730 (N_14730,N_9798,N_9742);
nand U14731 (N_14731,N_10370,N_10439);
xor U14732 (N_14732,N_9645,N_9161);
and U14733 (N_14733,N_10021,N_9408);
and U14734 (N_14734,N_11750,N_11825);
and U14735 (N_14735,N_10188,N_9420);
nand U14736 (N_14736,N_10220,N_11352);
xor U14737 (N_14737,N_9419,N_9599);
nand U14738 (N_14738,N_9474,N_11251);
nor U14739 (N_14739,N_11114,N_10944);
nand U14740 (N_14740,N_11725,N_11063);
and U14741 (N_14741,N_9204,N_9932);
nor U14742 (N_14742,N_9659,N_11932);
nor U14743 (N_14743,N_10039,N_10026);
nand U14744 (N_14744,N_10459,N_10438);
or U14745 (N_14745,N_10694,N_9804);
or U14746 (N_14746,N_11224,N_9563);
nand U14747 (N_14747,N_11289,N_10723);
nor U14748 (N_14748,N_10729,N_10786);
and U14749 (N_14749,N_9253,N_10169);
or U14750 (N_14750,N_9411,N_10893);
nor U14751 (N_14751,N_11458,N_9531);
and U14752 (N_14752,N_9423,N_11321);
nor U14753 (N_14753,N_11379,N_10581);
nand U14754 (N_14754,N_10935,N_10770);
nor U14755 (N_14755,N_10754,N_9557);
nor U14756 (N_14756,N_11306,N_11874);
nor U14757 (N_14757,N_10055,N_10739);
or U14758 (N_14758,N_10139,N_10926);
and U14759 (N_14759,N_11572,N_11045);
and U14760 (N_14760,N_11218,N_10069);
or U14761 (N_14761,N_11099,N_11852);
nand U14762 (N_14762,N_11208,N_9836);
and U14763 (N_14763,N_9236,N_9703);
nor U14764 (N_14764,N_11356,N_10106);
nand U14765 (N_14765,N_11412,N_10779);
or U14766 (N_14766,N_9886,N_9777);
nor U14767 (N_14767,N_9521,N_10864);
and U14768 (N_14768,N_10462,N_11817);
nor U14769 (N_14769,N_11179,N_10602);
and U14770 (N_14770,N_11187,N_9637);
xnor U14771 (N_14771,N_9457,N_10808);
or U14772 (N_14772,N_9619,N_9682);
nand U14773 (N_14773,N_10330,N_11137);
or U14774 (N_14774,N_10555,N_10207);
nor U14775 (N_14775,N_9712,N_11159);
nor U14776 (N_14776,N_11302,N_9180);
or U14777 (N_14777,N_11111,N_10118);
or U14778 (N_14778,N_9919,N_11389);
or U14779 (N_14779,N_9048,N_9199);
nand U14780 (N_14780,N_11604,N_9861);
xor U14781 (N_14781,N_10492,N_9532);
nand U14782 (N_14782,N_10658,N_11880);
nor U14783 (N_14783,N_10126,N_11966);
nand U14784 (N_14784,N_11559,N_9720);
or U14785 (N_14785,N_9826,N_11832);
xnor U14786 (N_14786,N_10137,N_9035);
and U14787 (N_14787,N_11688,N_10517);
nand U14788 (N_14788,N_10849,N_10498);
nor U14789 (N_14789,N_11628,N_9914);
or U14790 (N_14790,N_9276,N_9693);
nand U14791 (N_14791,N_11547,N_10524);
and U14792 (N_14792,N_9106,N_11141);
nor U14793 (N_14793,N_10852,N_10379);
and U14794 (N_14794,N_9654,N_10941);
or U14795 (N_14795,N_9235,N_11405);
xnor U14796 (N_14796,N_11051,N_10349);
and U14797 (N_14797,N_10622,N_10615);
nor U14798 (N_14798,N_11159,N_11262);
or U14799 (N_14799,N_10320,N_10909);
and U14800 (N_14800,N_9015,N_10753);
xor U14801 (N_14801,N_11035,N_10500);
nor U14802 (N_14802,N_11145,N_9746);
nor U14803 (N_14803,N_9545,N_10615);
xor U14804 (N_14804,N_11273,N_9125);
nor U14805 (N_14805,N_10012,N_10642);
and U14806 (N_14806,N_11292,N_9638);
xnor U14807 (N_14807,N_11653,N_11414);
and U14808 (N_14808,N_10943,N_11022);
xnor U14809 (N_14809,N_11817,N_11831);
nand U14810 (N_14810,N_11106,N_9808);
nor U14811 (N_14811,N_9893,N_10367);
nor U14812 (N_14812,N_9383,N_11554);
nor U14813 (N_14813,N_9802,N_11767);
nand U14814 (N_14814,N_9897,N_9278);
and U14815 (N_14815,N_11449,N_11537);
nor U14816 (N_14816,N_10811,N_9443);
nand U14817 (N_14817,N_9650,N_10807);
xor U14818 (N_14818,N_10486,N_11110);
nor U14819 (N_14819,N_9359,N_9416);
nor U14820 (N_14820,N_9266,N_10763);
and U14821 (N_14821,N_9197,N_10442);
or U14822 (N_14822,N_11114,N_9234);
or U14823 (N_14823,N_9970,N_9211);
nand U14824 (N_14824,N_10327,N_9211);
nand U14825 (N_14825,N_9799,N_9595);
nand U14826 (N_14826,N_11100,N_10575);
and U14827 (N_14827,N_10747,N_9282);
and U14828 (N_14828,N_11650,N_11131);
nand U14829 (N_14829,N_10851,N_11381);
xnor U14830 (N_14830,N_9811,N_9240);
nor U14831 (N_14831,N_10695,N_9164);
nor U14832 (N_14832,N_10803,N_11198);
or U14833 (N_14833,N_9276,N_11084);
xor U14834 (N_14834,N_10364,N_10512);
or U14835 (N_14835,N_10401,N_11407);
or U14836 (N_14836,N_9158,N_9395);
and U14837 (N_14837,N_10303,N_11549);
nand U14838 (N_14838,N_10439,N_9342);
or U14839 (N_14839,N_9353,N_9342);
nand U14840 (N_14840,N_10798,N_11336);
nand U14841 (N_14841,N_10325,N_10950);
and U14842 (N_14842,N_10052,N_10373);
and U14843 (N_14843,N_9990,N_9812);
or U14844 (N_14844,N_10094,N_9392);
or U14845 (N_14845,N_10224,N_11154);
and U14846 (N_14846,N_9251,N_10122);
and U14847 (N_14847,N_11614,N_11769);
xnor U14848 (N_14848,N_11249,N_10107);
and U14849 (N_14849,N_11002,N_11820);
nor U14850 (N_14850,N_10480,N_10434);
and U14851 (N_14851,N_10465,N_11468);
nand U14852 (N_14852,N_11100,N_10771);
nand U14853 (N_14853,N_11743,N_11240);
nor U14854 (N_14854,N_10557,N_10672);
and U14855 (N_14855,N_11100,N_10564);
nand U14856 (N_14856,N_11208,N_9172);
or U14857 (N_14857,N_9681,N_10034);
nor U14858 (N_14858,N_10394,N_11835);
or U14859 (N_14859,N_9650,N_10597);
nor U14860 (N_14860,N_10054,N_11370);
and U14861 (N_14861,N_9851,N_9791);
nor U14862 (N_14862,N_10361,N_11949);
and U14863 (N_14863,N_9545,N_10282);
nand U14864 (N_14864,N_11939,N_10507);
or U14865 (N_14865,N_9751,N_11522);
and U14866 (N_14866,N_11411,N_11049);
and U14867 (N_14867,N_9622,N_10656);
xor U14868 (N_14868,N_10751,N_11859);
or U14869 (N_14869,N_9777,N_11645);
xnor U14870 (N_14870,N_9982,N_11104);
or U14871 (N_14871,N_9311,N_10068);
or U14872 (N_14872,N_10538,N_11200);
nor U14873 (N_14873,N_9225,N_9073);
or U14874 (N_14874,N_9113,N_9795);
nand U14875 (N_14875,N_11898,N_11570);
or U14876 (N_14876,N_11397,N_10284);
nand U14877 (N_14877,N_10931,N_11661);
or U14878 (N_14878,N_10914,N_10817);
nand U14879 (N_14879,N_10588,N_9262);
and U14880 (N_14880,N_10227,N_11363);
nand U14881 (N_14881,N_11664,N_9854);
or U14882 (N_14882,N_9384,N_10744);
and U14883 (N_14883,N_11989,N_11621);
and U14884 (N_14884,N_9874,N_9595);
or U14885 (N_14885,N_10779,N_10296);
nand U14886 (N_14886,N_11022,N_10559);
and U14887 (N_14887,N_11321,N_11010);
xnor U14888 (N_14888,N_9116,N_11816);
and U14889 (N_14889,N_9788,N_11187);
and U14890 (N_14890,N_11187,N_9803);
or U14891 (N_14891,N_11688,N_10384);
nand U14892 (N_14892,N_11187,N_11085);
nand U14893 (N_14893,N_10221,N_10874);
or U14894 (N_14894,N_9545,N_9789);
nand U14895 (N_14895,N_9378,N_9094);
and U14896 (N_14896,N_11995,N_9329);
and U14897 (N_14897,N_10577,N_9548);
and U14898 (N_14898,N_10572,N_10437);
nand U14899 (N_14899,N_9675,N_9811);
nor U14900 (N_14900,N_9129,N_11343);
nand U14901 (N_14901,N_10419,N_11673);
and U14902 (N_14902,N_9031,N_11416);
nor U14903 (N_14903,N_9782,N_11647);
and U14904 (N_14904,N_11861,N_9994);
or U14905 (N_14905,N_11848,N_11369);
nand U14906 (N_14906,N_11476,N_11231);
nor U14907 (N_14907,N_10848,N_9249);
nor U14908 (N_14908,N_9981,N_11060);
and U14909 (N_14909,N_11844,N_10622);
xor U14910 (N_14910,N_11016,N_9024);
nor U14911 (N_14911,N_9659,N_10114);
or U14912 (N_14912,N_10409,N_9222);
or U14913 (N_14913,N_10239,N_9746);
and U14914 (N_14914,N_11783,N_9550);
nand U14915 (N_14915,N_10541,N_11362);
or U14916 (N_14916,N_9917,N_9103);
nand U14917 (N_14917,N_9273,N_10878);
and U14918 (N_14918,N_9549,N_10876);
nand U14919 (N_14919,N_10533,N_11467);
nand U14920 (N_14920,N_9310,N_11467);
and U14921 (N_14921,N_10771,N_11607);
nand U14922 (N_14922,N_9175,N_10102);
xnor U14923 (N_14923,N_11553,N_11601);
and U14924 (N_14924,N_10200,N_11836);
or U14925 (N_14925,N_11706,N_9326);
nor U14926 (N_14926,N_10160,N_9732);
nand U14927 (N_14927,N_10515,N_9379);
nor U14928 (N_14928,N_10769,N_10117);
nand U14929 (N_14929,N_11084,N_11937);
nand U14930 (N_14930,N_10768,N_9583);
and U14931 (N_14931,N_9490,N_11213);
nand U14932 (N_14932,N_9866,N_10242);
nand U14933 (N_14933,N_10513,N_10418);
nor U14934 (N_14934,N_11186,N_11675);
or U14935 (N_14935,N_11054,N_10284);
nor U14936 (N_14936,N_9406,N_11337);
nor U14937 (N_14937,N_10441,N_9820);
or U14938 (N_14938,N_10295,N_9444);
xnor U14939 (N_14939,N_9221,N_10928);
and U14940 (N_14940,N_9558,N_11407);
xor U14941 (N_14941,N_10770,N_10171);
nor U14942 (N_14942,N_9689,N_9508);
xnor U14943 (N_14943,N_11308,N_11697);
or U14944 (N_14944,N_10845,N_11273);
or U14945 (N_14945,N_10021,N_10384);
or U14946 (N_14946,N_10986,N_9893);
and U14947 (N_14947,N_9866,N_10750);
nor U14948 (N_14948,N_9062,N_10339);
nor U14949 (N_14949,N_9211,N_10826);
nand U14950 (N_14950,N_10315,N_9508);
nor U14951 (N_14951,N_9065,N_10457);
xor U14952 (N_14952,N_11173,N_11771);
and U14953 (N_14953,N_10646,N_10464);
xor U14954 (N_14954,N_11070,N_11663);
nor U14955 (N_14955,N_9303,N_9761);
and U14956 (N_14956,N_11652,N_10800);
nand U14957 (N_14957,N_11638,N_9184);
nor U14958 (N_14958,N_10813,N_10625);
or U14959 (N_14959,N_11071,N_11746);
xnor U14960 (N_14960,N_11154,N_9682);
or U14961 (N_14961,N_9558,N_10878);
and U14962 (N_14962,N_9740,N_9017);
or U14963 (N_14963,N_10359,N_11514);
and U14964 (N_14964,N_10684,N_9505);
and U14965 (N_14965,N_10610,N_10854);
nor U14966 (N_14966,N_11264,N_9908);
and U14967 (N_14967,N_11761,N_11183);
or U14968 (N_14968,N_10886,N_9784);
nand U14969 (N_14969,N_10972,N_9128);
nand U14970 (N_14970,N_9880,N_9163);
xor U14971 (N_14971,N_11121,N_10831);
and U14972 (N_14972,N_10294,N_9406);
or U14973 (N_14973,N_11258,N_10971);
and U14974 (N_14974,N_9613,N_11483);
and U14975 (N_14975,N_10860,N_11737);
or U14976 (N_14976,N_9910,N_11544);
and U14977 (N_14977,N_11665,N_11455);
nand U14978 (N_14978,N_10726,N_10698);
or U14979 (N_14979,N_11765,N_10291);
nor U14980 (N_14980,N_9862,N_11460);
nand U14981 (N_14981,N_11116,N_10235);
nand U14982 (N_14982,N_11302,N_10250);
nand U14983 (N_14983,N_11685,N_11502);
or U14984 (N_14984,N_10312,N_11513);
nor U14985 (N_14985,N_11902,N_11527);
and U14986 (N_14986,N_11766,N_9893);
nor U14987 (N_14987,N_9310,N_11095);
and U14988 (N_14988,N_11823,N_10413);
nor U14989 (N_14989,N_11446,N_11550);
nand U14990 (N_14990,N_10688,N_10985);
nor U14991 (N_14991,N_11093,N_10859);
or U14992 (N_14992,N_9377,N_10432);
or U14993 (N_14993,N_11305,N_11977);
nand U14994 (N_14994,N_9332,N_10236);
xor U14995 (N_14995,N_10772,N_10055);
xor U14996 (N_14996,N_9264,N_10489);
or U14997 (N_14997,N_9021,N_11754);
nor U14998 (N_14998,N_10061,N_9782);
nand U14999 (N_14999,N_10640,N_9457);
or UO_0 (O_0,N_12467,N_14743);
and UO_1 (O_1,N_14301,N_14079);
nand UO_2 (O_2,N_13911,N_12485);
nor UO_3 (O_3,N_14159,N_12086);
and UO_4 (O_4,N_13136,N_12650);
xnor UO_5 (O_5,N_14285,N_12255);
or UO_6 (O_6,N_13485,N_12788);
nor UO_7 (O_7,N_14997,N_13410);
xor UO_8 (O_8,N_14987,N_13089);
xnor UO_9 (O_9,N_12819,N_14684);
nand UO_10 (O_10,N_13026,N_12143);
or UO_11 (O_11,N_12980,N_12428);
nor UO_12 (O_12,N_12663,N_14668);
nand UO_13 (O_13,N_14686,N_12187);
nand UO_14 (O_14,N_13658,N_13888);
nand UO_15 (O_15,N_12034,N_13066);
nor UO_16 (O_16,N_12988,N_13320);
xor UO_17 (O_17,N_13542,N_12498);
and UO_18 (O_18,N_14227,N_12948);
or UO_19 (O_19,N_12276,N_14157);
xor UO_20 (O_20,N_14822,N_14208);
and UO_21 (O_21,N_13204,N_12212);
nor UO_22 (O_22,N_14274,N_12122);
and UO_23 (O_23,N_12533,N_13522);
or UO_24 (O_24,N_14190,N_12400);
nor UO_25 (O_25,N_14846,N_13424);
nor UO_26 (O_26,N_14031,N_12053);
and UO_27 (O_27,N_14189,N_13982);
or UO_28 (O_28,N_14792,N_13920);
nand UO_29 (O_29,N_14739,N_12188);
nand UO_30 (O_30,N_12447,N_13802);
nand UO_31 (O_31,N_12911,N_14331);
or UO_32 (O_32,N_13960,N_14417);
or UO_33 (O_33,N_14590,N_12454);
or UO_34 (O_34,N_12453,N_13489);
nand UO_35 (O_35,N_12012,N_13878);
and UO_36 (O_36,N_13285,N_13723);
and UO_37 (O_37,N_14669,N_12360);
xnor UO_38 (O_38,N_14772,N_12801);
nor UO_39 (O_39,N_13994,N_14513);
nand UO_40 (O_40,N_14477,N_13684);
or UO_41 (O_41,N_12140,N_12517);
nor UO_42 (O_42,N_13762,N_12662);
nand UO_43 (O_43,N_14631,N_13668);
xnor UO_44 (O_44,N_12219,N_12719);
or UO_45 (O_45,N_14712,N_14880);
nor UO_46 (O_46,N_13850,N_14185);
nand UO_47 (O_47,N_12218,N_12385);
xor UO_48 (O_48,N_13074,N_12446);
and UO_49 (O_49,N_13621,N_12025);
nor UO_50 (O_50,N_13192,N_12304);
nand UO_51 (O_51,N_12977,N_13397);
xor UO_52 (O_52,N_12828,N_14788);
xor UO_53 (O_53,N_13166,N_14089);
or UO_54 (O_54,N_13647,N_12114);
nor UO_55 (O_55,N_12322,N_12826);
or UO_56 (O_56,N_13387,N_12279);
and UO_57 (O_57,N_12550,N_14926);
nand UO_58 (O_58,N_13771,N_13624);
nor UO_59 (O_59,N_14213,N_13447);
nor UO_60 (O_60,N_13296,N_12127);
nor UO_61 (O_61,N_13707,N_12995);
xor UO_62 (O_62,N_14796,N_13495);
or UO_63 (O_63,N_13774,N_13239);
xor UO_64 (O_64,N_14807,N_12370);
and UO_65 (O_65,N_14884,N_12990);
and UO_66 (O_66,N_14637,N_13950);
and UO_67 (O_67,N_14550,N_13270);
nand UO_68 (O_68,N_13109,N_12777);
nand UO_69 (O_69,N_13217,N_14183);
nand UO_70 (O_70,N_13949,N_12561);
xor UO_71 (O_71,N_14278,N_12445);
nand UO_72 (O_72,N_13813,N_12104);
nand UO_73 (O_73,N_14528,N_14670);
or UO_74 (O_74,N_12917,N_12366);
xor UO_75 (O_75,N_13246,N_13745);
and UO_76 (O_76,N_13251,N_13797);
and UO_77 (O_77,N_14971,N_14257);
and UO_78 (O_78,N_14965,N_14072);
and UO_79 (O_79,N_13313,N_13206);
nor UO_80 (O_80,N_12426,N_14959);
and UO_81 (O_81,N_14800,N_14137);
and UO_82 (O_82,N_12307,N_12209);
or UO_83 (O_83,N_14962,N_14354);
nand UO_84 (O_84,N_14107,N_14479);
nor UO_85 (O_85,N_12331,N_13283);
nand UO_86 (O_86,N_14972,N_12480);
and UO_87 (O_87,N_12141,N_13778);
xnor UO_88 (O_88,N_14705,N_13901);
nand UO_89 (O_89,N_14587,N_13929);
or UO_90 (O_90,N_13677,N_13195);
and UO_91 (O_91,N_14936,N_13405);
xnor UO_92 (O_92,N_12644,N_14828);
or UO_93 (O_93,N_12891,N_14174);
and UO_94 (O_94,N_13683,N_13930);
nand UO_95 (O_95,N_14088,N_13606);
nand UO_96 (O_96,N_14261,N_12146);
xor UO_97 (O_97,N_13386,N_12548);
nor UO_98 (O_98,N_12349,N_13008);
nor UO_99 (O_99,N_14724,N_13655);
or UO_100 (O_100,N_14140,N_12878);
nor UO_101 (O_101,N_14533,N_13198);
nor UO_102 (O_102,N_14702,N_14620);
nor UO_103 (O_103,N_12392,N_14503);
and UO_104 (O_104,N_14225,N_12634);
and UO_105 (O_105,N_12551,N_13775);
or UO_106 (O_106,N_12513,N_12975);
nand UO_107 (O_107,N_12200,N_12386);
and UO_108 (O_108,N_12721,N_13098);
or UO_109 (O_109,N_13629,N_13880);
xnor UO_110 (O_110,N_12302,N_13600);
nor UO_111 (O_111,N_13943,N_13072);
nand UO_112 (O_112,N_13815,N_13203);
and UO_113 (O_113,N_13404,N_12181);
or UO_114 (O_114,N_13602,N_13838);
or UO_115 (O_115,N_14166,N_12001);
and UO_116 (O_116,N_13961,N_14595);
nor UO_117 (O_117,N_13037,N_13071);
and UO_118 (O_118,N_14740,N_14141);
or UO_119 (O_119,N_14838,N_14639);
nor UO_120 (O_120,N_14333,N_14520);
xnor UO_121 (O_121,N_13486,N_13261);
and UO_122 (O_122,N_12088,N_14224);
nand UO_123 (O_123,N_14614,N_13147);
xor UO_124 (O_124,N_13401,N_14570);
nor UO_125 (O_125,N_13443,N_13471);
or UO_126 (O_126,N_12961,N_12866);
xor UO_127 (O_127,N_13371,N_12616);
nand UO_128 (O_128,N_12482,N_14797);
nand UO_129 (O_129,N_13384,N_12109);
or UO_130 (O_130,N_13383,N_14835);
and UO_131 (O_131,N_12903,N_14019);
nor UO_132 (O_132,N_13228,N_14658);
and UO_133 (O_133,N_14554,N_14397);
and UO_134 (O_134,N_13230,N_12611);
nand UO_135 (O_135,N_13288,N_14337);
nand UO_136 (O_136,N_12741,N_14351);
nand UO_137 (O_137,N_14234,N_13141);
nor UO_138 (O_138,N_12997,N_13693);
nor UO_139 (O_139,N_13804,N_12003);
xor UO_140 (O_140,N_12887,N_13400);
and UO_141 (O_141,N_12798,N_14130);
nor UO_142 (O_142,N_13127,N_12247);
nor UO_143 (O_143,N_12009,N_12087);
xnor UO_144 (O_144,N_12309,N_14223);
nand UO_145 (O_145,N_13987,N_12368);
nor UO_146 (O_146,N_14707,N_14110);
nor UO_147 (O_147,N_13157,N_12857);
xnor UO_148 (O_148,N_12052,N_12672);
nand UO_149 (O_149,N_12422,N_14194);
nand UO_150 (O_150,N_12110,N_12591);
or UO_151 (O_151,N_14402,N_12364);
and UO_152 (O_152,N_14470,N_12335);
and UO_153 (O_153,N_13682,N_13910);
or UO_154 (O_154,N_13014,N_13879);
nand UO_155 (O_155,N_13069,N_13044);
nor UO_156 (O_156,N_12680,N_14552);
nand UO_157 (O_157,N_12705,N_13670);
nand UO_158 (O_158,N_14853,N_12198);
xnor UO_159 (O_159,N_14051,N_13211);
nand UO_160 (O_160,N_13795,N_14603);
nor UO_161 (O_161,N_14693,N_14217);
and UO_162 (O_162,N_14376,N_14336);
nand UO_163 (O_163,N_14370,N_12691);
or UO_164 (O_164,N_14934,N_12115);
nand UO_165 (O_165,N_13500,N_13526);
and UO_166 (O_166,N_13169,N_13000);
nand UO_167 (O_167,N_14499,N_12068);
and UO_168 (O_168,N_12885,N_14979);
or UO_169 (O_169,N_13926,N_12633);
or UO_170 (O_170,N_12005,N_13590);
or UO_171 (O_171,N_12210,N_14395);
or UO_172 (O_172,N_12154,N_13005);
and UO_173 (O_173,N_13364,N_14429);
xnor UO_174 (O_174,N_13913,N_14472);
xnor UO_175 (O_175,N_13969,N_14868);
nor UO_176 (O_176,N_12519,N_12372);
xor UO_177 (O_177,N_13488,N_13808);
nand UO_178 (O_178,N_13610,N_14725);
and UO_179 (O_179,N_13341,N_14640);
or UO_180 (O_180,N_12531,N_12888);
and UO_181 (O_181,N_13751,N_14540);
and UO_182 (O_182,N_12135,N_12176);
or UO_183 (O_183,N_13536,N_14327);
nand UO_184 (O_184,N_13126,N_12676);
nor UO_185 (O_185,N_14302,N_14632);
nand UO_186 (O_186,N_14268,N_13783);
nor UO_187 (O_187,N_13855,N_14296);
xnor UO_188 (O_188,N_12503,N_12293);
and UO_189 (O_189,N_12946,N_13422);
nand UO_190 (O_190,N_13511,N_13963);
nand UO_191 (O_191,N_12105,N_12500);
or UO_192 (O_192,N_13053,N_13001);
xor UO_193 (O_193,N_12424,N_14978);
or UO_194 (O_194,N_12021,N_14392);
and UO_195 (O_195,N_13437,N_13561);
nor UO_196 (O_196,N_14332,N_12452);
nand UO_197 (O_197,N_12677,N_13361);
and UO_198 (O_198,N_13247,N_12556);
nand UO_199 (O_199,N_13968,N_14451);
or UO_200 (O_200,N_13193,N_13108);
nor UO_201 (O_201,N_13667,N_13235);
nor UO_202 (O_202,N_12745,N_12472);
nor UO_203 (O_203,N_14678,N_13923);
or UO_204 (O_204,N_14087,N_12404);
nand UO_205 (O_205,N_13517,N_12681);
and UO_206 (O_206,N_12092,N_13036);
nand UO_207 (O_207,N_12489,N_14131);
nand UO_208 (O_208,N_13845,N_12495);
and UO_209 (O_209,N_12768,N_12215);
xor UO_210 (O_210,N_13398,N_14720);
and UO_211 (O_211,N_14653,N_13591);
nand UO_212 (O_212,N_13138,N_14326);
and UO_213 (O_213,N_14044,N_14246);
nand UO_214 (O_214,N_12241,N_12189);
nand UO_215 (O_215,N_14214,N_14318);
and UO_216 (O_216,N_14601,N_13290);
nor UO_217 (O_217,N_14985,N_14976);
nand UO_218 (O_218,N_14467,N_12994);
nor UO_219 (O_219,N_13777,N_12282);
or UO_220 (O_220,N_14761,N_12195);
nand UO_221 (O_221,N_12553,N_12317);
or UO_222 (O_222,N_14888,N_12585);
xor UO_223 (O_223,N_13515,N_12466);
and UO_224 (O_224,N_12343,N_13834);
nor UO_225 (O_225,N_14875,N_14991);
or UO_226 (O_226,N_12753,N_12532);
nor UO_227 (O_227,N_12406,N_13535);
or UO_228 (O_228,N_13043,N_14464);
and UO_229 (O_229,N_12675,N_14685);
or UO_230 (O_230,N_13651,N_13832);
nand UO_231 (O_231,N_14852,N_13440);
and UO_232 (O_232,N_13004,N_12514);
nand UO_233 (O_233,N_14945,N_12837);
nor UO_234 (O_234,N_14617,N_12265);
nand UO_235 (O_235,N_12256,N_12496);
nand UO_236 (O_236,N_13986,N_13512);
nor UO_237 (O_237,N_13611,N_14924);
and UO_238 (O_238,N_12225,N_12733);
nor UO_239 (O_239,N_12197,N_12940);
or UO_240 (O_240,N_13249,N_12038);
or UO_241 (O_241,N_12968,N_14633);
nand UO_242 (O_242,N_13978,N_14903);
or UO_243 (O_243,N_14308,N_14018);
nand UO_244 (O_244,N_13831,N_12341);
xnor UO_245 (O_245,N_12403,N_12702);
nor UO_246 (O_246,N_13612,N_13349);
nor UO_247 (O_247,N_12699,N_14917);
xnor UO_248 (O_248,N_13750,N_12574);
and UO_249 (O_249,N_14375,N_12145);
nor UO_250 (O_250,N_12336,N_12421);
nor UO_251 (O_251,N_13768,N_12600);
or UO_252 (O_252,N_12128,N_12919);
and UO_253 (O_253,N_14241,N_13367);
nor UO_254 (O_254,N_13639,N_13685);
nor UO_255 (O_255,N_14656,N_14863);
nand UO_256 (O_256,N_13408,N_13946);
and UO_257 (O_257,N_14950,N_12880);
nor UO_258 (O_258,N_12061,N_13273);
or UO_259 (O_259,N_12910,N_13353);
nor UO_260 (O_260,N_13550,N_12642);
or UO_261 (O_261,N_12897,N_14607);
nand UO_262 (O_262,N_14267,N_12410);
xnor UO_263 (O_263,N_13406,N_12180);
or UO_264 (O_264,N_14999,N_12593);
nor UO_265 (O_265,N_14476,N_14886);
or UO_266 (O_266,N_13415,N_13182);
and UO_267 (O_267,N_14430,N_14841);
and UO_268 (O_268,N_12230,N_12383);
or UO_269 (O_269,N_13102,N_13174);
or UO_270 (O_270,N_14180,N_13105);
nor UO_271 (O_271,N_14054,N_13974);
or UO_272 (O_272,N_13359,N_13029);
or UO_273 (O_273,N_12795,N_12484);
nor UO_274 (O_274,N_12831,N_14855);
nand UO_275 (O_275,N_12543,N_12814);
nor UO_276 (O_276,N_12070,N_12079);
or UO_277 (O_277,N_12545,N_13128);
and UO_278 (O_278,N_14168,N_14240);
xnor UO_279 (O_279,N_14303,N_12344);
nor UO_280 (O_280,N_13900,N_14592);
and UO_281 (O_281,N_12435,N_13445);
and UO_282 (O_282,N_13819,N_14857);
nor UO_283 (O_283,N_14004,N_12757);
nand UO_284 (O_284,N_13856,N_13134);
xnor UO_285 (O_285,N_13977,N_13653);
nor UO_286 (O_286,N_14751,N_13393);
xor UO_287 (O_287,N_14727,N_13649);
or UO_288 (O_288,N_12048,N_14277);
nand UO_289 (O_289,N_14813,N_13899);
nor UO_290 (O_290,N_13333,N_13483);
or UO_291 (O_291,N_12520,N_13593);
and UO_292 (O_292,N_14650,N_14039);
and UO_293 (O_293,N_14275,N_14981);
nand UO_294 (O_294,N_14239,N_14534);
nor UO_295 (O_295,N_13112,N_12799);
or UO_296 (O_296,N_12779,N_12217);
nor UO_297 (O_297,N_12129,N_13788);
xor UO_298 (O_298,N_12505,N_12248);
nand UO_299 (O_299,N_12440,N_13948);
xnor UO_300 (O_300,N_14272,N_14803);
and UO_301 (O_301,N_14372,N_14027);
and UO_302 (O_302,N_13881,N_14635);
or UO_303 (O_303,N_13708,N_14742);
or UO_304 (O_304,N_14488,N_12050);
nor UO_305 (O_305,N_13081,N_12017);
nand UO_306 (O_306,N_12729,N_12182);
nor UO_307 (O_307,N_13730,N_12027);
or UO_308 (O_308,N_13318,N_12029);
and UO_309 (O_309,N_14613,N_13478);
and UO_310 (O_310,N_13742,N_14427);
nand UO_311 (O_311,N_12504,N_12155);
nand UO_312 (O_312,N_14634,N_12627);
nand UO_313 (O_313,N_14485,N_14290);
nand UO_314 (O_314,N_14755,N_12340);
or UO_315 (O_315,N_13619,N_14484);
or UO_316 (O_316,N_13620,N_13958);
xnor UO_317 (O_317,N_12853,N_14573);
nor UO_318 (O_318,N_14134,N_13458);
nor UO_319 (O_319,N_14314,N_13291);
nor UO_320 (O_320,N_14776,N_12950);
nand UO_321 (O_321,N_14989,N_12413);
and UO_322 (O_322,N_12186,N_13385);
nand UO_323 (O_323,N_14942,N_14226);
nand UO_324 (O_324,N_13570,N_14017);
nand UO_325 (O_325,N_13565,N_14728);
nand UO_326 (O_326,N_12235,N_14567);
nor UO_327 (O_327,N_12151,N_14569);
nand UO_328 (O_328,N_12486,N_12414);
nand UO_329 (O_329,N_13010,N_14309);
and UO_330 (O_330,N_12572,N_13094);
nor UO_331 (O_331,N_14921,N_14457);
nand UO_332 (O_332,N_14220,N_14594);
nand UO_333 (O_333,N_12024,N_13068);
nand UO_334 (O_334,N_12196,N_13727);
or UO_335 (O_335,N_13197,N_13914);
and UO_336 (O_336,N_13607,N_13477);
and UO_337 (O_337,N_12631,N_12264);
nor UO_338 (O_338,N_13316,N_13173);
nor UO_339 (O_339,N_14008,N_14930);
nand UO_340 (O_340,N_14894,N_12571);
or UO_341 (O_341,N_13379,N_12771);
and UO_342 (O_342,N_14709,N_13549);
and UO_343 (O_343,N_14698,N_13547);
or UO_344 (O_344,N_12845,N_12071);
and UO_345 (O_345,N_13148,N_12957);
nor UO_346 (O_346,N_12947,N_13711);
and UO_347 (O_347,N_12666,N_12442);
and UO_348 (O_348,N_14568,N_13916);
xnor UO_349 (O_349,N_14064,N_13703);
and UO_350 (O_350,N_14492,N_14010);
xor UO_351 (O_351,N_12286,N_13733);
nand UO_352 (O_352,N_12359,N_14167);
and UO_353 (O_353,N_14150,N_14135);
nand UO_354 (O_354,N_14919,N_12530);
nand UO_355 (O_355,N_13131,N_12494);
nand UO_356 (O_356,N_12327,N_14915);
and UO_357 (O_357,N_13934,N_14906);
and UO_358 (O_358,N_12091,N_13671);
or UO_359 (O_359,N_12963,N_12417);
or UO_360 (O_360,N_12874,N_12546);
nor UO_361 (O_361,N_14366,N_12684);
nor UO_362 (O_362,N_12405,N_12624);
nor UO_363 (O_363,N_14374,N_13221);
nand UO_364 (O_364,N_13669,N_12773);
nand UO_365 (O_365,N_12010,N_13793);
or UO_366 (O_366,N_14348,N_13842);
nor UO_367 (O_367,N_14901,N_12808);
and UO_368 (O_368,N_12082,N_12904);
and UO_369 (O_369,N_13862,N_12746);
nor UO_370 (O_370,N_13487,N_13678);
or UO_371 (O_371,N_12185,N_12369);
and UO_372 (O_372,N_14158,N_12588);
nand UO_373 (O_373,N_14862,N_14378);
nand UO_374 (O_374,N_13013,N_13431);
nor UO_375 (O_375,N_14877,N_12085);
xnor UO_376 (O_376,N_13566,N_12156);
nand UO_377 (O_377,N_12411,N_12342);
nor UO_378 (O_378,N_13334,N_12796);
nand UO_379 (O_379,N_13971,N_12031);
xor UO_380 (O_380,N_12475,N_12610);
nand UO_381 (O_381,N_13615,N_14016);
and UO_382 (O_382,N_12685,N_14462);
or UO_383 (O_383,N_12626,N_12657);
or UO_384 (O_384,N_12924,N_13338);
xnor UO_385 (O_385,N_14491,N_14145);
nor UO_386 (O_386,N_12867,N_14029);
and UO_387 (O_387,N_14094,N_13799);
nor UO_388 (O_388,N_12351,N_12352);
nand UO_389 (O_389,N_13731,N_13265);
nand UO_390 (O_390,N_13079,N_14316);
nor UO_391 (O_391,N_13409,N_13854);
and UO_392 (O_392,N_12178,N_12620);
and UO_393 (O_393,N_12328,N_12438);
nand UO_394 (O_394,N_12075,N_12204);
nand UO_395 (O_395,N_12966,N_13597);
and UO_396 (O_396,N_14898,N_13114);
or UO_397 (O_397,N_14300,N_13552);
xnor UO_398 (O_398,N_13695,N_14970);
nand UO_399 (O_399,N_14990,N_12488);
or UO_400 (O_400,N_13618,N_12169);
or UO_401 (O_401,N_13705,N_13048);
nor UO_402 (O_402,N_14746,N_13609);
nor UO_403 (O_403,N_13534,N_13321);
xor UO_404 (O_404,N_14619,N_13787);
and UO_405 (O_405,N_14806,N_14923);
nor UO_406 (O_406,N_13186,N_12971);
nand UO_407 (O_407,N_14505,N_13663);
nor UO_408 (O_408,N_14986,N_12938);
or UO_409 (O_409,N_12784,N_13311);
nor UO_410 (O_410,N_14791,N_14249);
or UO_411 (O_411,N_13820,N_12066);
nor UO_412 (O_412,N_12497,N_12415);
nand UO_413 (O_413,N_13202,N_14691);
and UO_414 (O_414,N_14666,N_13399);
or UO_415 (O_415,N_14416,N_12764);
nand UO_416 (O_416,N_14322,N_13065);
nand UO_417 (O_417,N_14683,N_14897);
and UO_418 (O_418,N_14993,N_12858);
nor UO_419 (O_419,N_12555,N_12371);
xnor UO_420 (O_420,N_12308,N_14773);
or UO_421 (O_421,N_14817,N_12022);
and UO_422 (O_422,N_14022,N_14273);
nor UO_423 (O_423,N_13137,N_14182);
nor UO_424 (O_424,N_13622,N_14338);
or UO_425 (O_425,N_13501,N_13664);
xnor UO_426 (O_426,N_12639,N_12348);
xnor UO_427 (O_427,N_13248,N_13741);
and UO_428 (O_428,N_14958,N_12823);
xnor UO_429 (O_429,N_12043,N_14968);
xnor UO_430 (O_430,N_12292,N_12817);
or UO_431 (O_431,N_13067,N_12688);
and UO_432 (O_432,N_14695,N_13282);
or UO_433 (O_433,N_12515,N_12338);
nor UO_434 (O_434,N_14892,N_13699);
and UO_435 (O_435,N_13633,N_13275);
nor UO_436 (O_436,N_13375,N_12875);
or UO_437 (O_437,N_13421,N_12587);
nand UO_438 (O_438,N_12617,N_14536);
or UO_439 (O_439,N_12076,N_13363);
nor UO_440 (O_440,N_13608,N_12802);
nor UO_441 (O_441,N_13964,N_14280);
xor UO_442 (O_442,N_14541,N_12395);
nor UO_443 (O_443,N_12843,N_13631);
or UO_444 (O_444,N_13906,N_13464);
nor UO_445 (O_445,N_12989,N_12266);
nor UO_446 (O_446,N_14809,N_14516);
nor UO_447 (O_447,N_13821,N_12566);
nand UO_448 (O_448,N_14527,N_14202);
nand UO_449 (O_449,N_14344,N_12873);
or UO_450 (O_450,N_13738,N_13583);
nand UO_451 (O_451,N_13706,N_12646);
nor UO_452 (O_452,N_12298,N_14933);
and UO_453 (O_453,N_14198,N_12905);
or UO_454 (O_454,N_14252,N_12173);
nand UO_455 (O_455,N_12608,N_14657);
nor UO_456 (O_456,N_12237,N_13352);
nand UO_457 (O_457,N_13272,N_12936);
nand UO_458 (O_458,N_13687,N_13319);
nand UO_459 (O_459,N_13064,N_13234);
xnor UO_460 (O_460,N_12430,N_13133);
xnor UO_461 (O_461,N_14245,N_12992);
xnor UO_462 (O_462,N_12490,N_13945);
or UO_463 (O_463,N_14621,N_12429);
nand UO_464 (O_464,N_13915,N_13973);
nor UO_465 (O_465,N_12060,N_13567);
xnor UO_466 (O_466,N_14099,N_13446);
or UO_467 (O_467,N_14526,N_13190);
or UO_468 (O_468,N_12725,N_13376);
or UO_469 (O_469,N_13019,N_13849);
or UO_470 (O_470,N_14144,N_13308);
or UO_471 (O_471,N_14545,N_13274);
nor UO_472 (O_472,N_13902,N_13581);
and UO_473 (O_473,N_12310,N_13990);
and UO_474 (O_474,N_13419,N_12002);
xor UO_475 (O_475,N_13191,N_13231);
nand UO_476 (O_476,N_13207,N_14057);
nand UO_477 (O_477,N_13205,N_13729);
nand UO_478 (O_478,N_14823,N_13761);
and UO_479 (O_479,N_13944,N_14365);
and UO_480 (O_480,N_14098,N_14932);
nand UO_481 (O_481,N_14410,N_13144);
nand UO_482 (O_482,N_14049,N_14500);
and UO_483 (O_483,N_12559,N_14565);
nor UO_484 (O_484,N_13860,N_13080);
nor UO_485 (O_485,N_14982,N_12747);
nor UO_486 (O_486,N_12019,N_12791);
and UO_487 (O_487,N_12419,N_13891);
or UO_488 (O_488,N_13335,N_12996);
xnor UO_489 (O_489,N_14576,N_14518);
nand UO_490 (O_490,N_14538,N_13253);
xor UO_491 (O_491,N_14584,N_13942);
nand UO_492 (O_492,N_12014,N_12597);
and UO_493 (O_493,N_13996,N_13345);
or UO_494 (O_494,N_14081,N_13011);
or UO_495 (O_495,N_13689,N_14086);
nor UO_496 (O_496,N_13697,N_14007);
nand UO_497 (O_497,N_14649,N_13225);
xnor UO_498 (O_498,N_13473,N_13613);
or UO_499 (O_499,N_12922,N_13055);
nor UO_500 (O_500,N_14313,N_13666);
and UO_501 (O_501,N_12535,N_12923);
or UO_502 (O_502,N_12337,N_13800);
xnor UO_503 (O_503,N_12300,N_12149);
or UO_504 (O_504,N_12810,N_13056);
nand UO_505 (O_505,N_13165,N_12638);
nand UO_506 (O_506,N_13937,N_13301);
nor UO_507 (O_507,N_13213,N_13472);
nor UO_508 (O_508,N_12578,N_13524);
and UO_509 (O_509,N_13630,N_12201);
and UO_510 (O_510,N_14170,N_12899);
and UO_511 (O_511,N_14895,N_14943);
xnor UO_512 (O_512,N_14889,N_12640);
nor UO_513 (O_513,N_14222,N_14701);
nor UO_514 (O_514,N_12125,N_13113);
nor UO_515 (O_515,N_12269,N_14095);
and UO_516 (O_516,N_14381,N_14544);
xor UO_517 (O_517,N_12660,N_14449);
or UO_518 (O_518,N_13719,N_12973);
or UO_519 (O_519,N_13388,N_14865);
nor UO_520 (O_520,N_12516,N_14251);
or UO_521 (O_521,N_12781,N_12157);
nand UO_522 (O_522,N_13007,N_14328);
nand UO_523 (O_523,N_12894,N_13339);
and UO_524 (O_524,N_12208,N_13040);
nor UO_525 (O_525,N_12907,N_14553);
and UO_526 (O_526,N_14474,N_14164);
nand UO_527 (O_527,N_13784,N_14385);
nand UO_528 (O_528,N_12261,N_13662);
nor UO_529 (O_529,N_14784,N_12493);
xnor UO_530 (O_530,N_13219,N_14101);
and UO_531 (O_531,N_13972,N_13521);
nand UO_532 (O_532,N_14831,N_12199);
and UO_533 (O_533,N_12123,N_14711);
or UO_534 (O_534,N_13728,N_13051);
nor UO_535 (O_535,N_14952,N_12730);
nor UO_536 (O_536,N_13786,N_12929);
xnor UO_537 (O_537,N_14181,N_13470);
nand UO_538 (O_538,N_12776,N_14061);
nand UO_539 (O_539,N_13380,N_12981);
xor UO_540 (O_540,N_12399,N_12621);
or UO_541 (O_541,N_13822,N_12306);
nand UO_542 (O_542,N_12117,N_14789);
nand UO_543 (O_543,N_13830,N_13455);
xnor UO_544 (O_544,N_14660,N_13857);
nor UO_545 (O_545,N_12096,N_14264);
nand UO_546 (O_546,N_12761,N_12635);
nand UO_547 (O_547,N_13932,N_14045);
and UO_548 (O_548,N_12770,N_12321);
nor UO_549 (O_549,N_14187,N_14368);
or UO_550 (O_550,N_13256,N_13243);
and UO_551 (O_551,N_12815,N_14913);
and UO_552 (O_552,N_12964,N_14816);
or UO_553 (O_553,N_13870,N_13402);
xor UO_554 (O_554,N_14078,N_13764);
nand UO_555 (O_555,N_12315,N_14748);
xor UO_556 (O_556,N_13546,N_13450);
or UO_557 (O_557,N_12373,N_12704);
and UO_558 (O_558,N_14342,N_13954);
or UO_559 (O_559,N_14539,N_13598);
xor UO_560 (O_560,N_12103,N_12203);
and UO_561 (O_561,N_12107,N_12982);
or UO_562 (O_562,N_12737,N_12257);
nor UO_563 (O_563,N_13263,N_12769);
nand UO_564 (O_564,N_13720,N_13578);
nand UO_565 (O_565,N_14269,N_12731);
and UO_566 (O_566,N_12668,N_13589);
or UO_567 (O_567,N_14242,N_13149);
and UO_568 (O_568,N_13603,N_13344);
and UO_569 (O_569,N_13616,N_12877);
nor UO_570 (O_570,N_14311,N_12972);
xnor UO_571 (O_571,N_13289,N_12649);
nand UO_572 (O_572,N_13718,N_13518);
nor UO_573 (O_573,N_12120,N_13840);
or UO_574 (O_574,N_14357,N_13414);
nand UO_575 (O_575,N_12920,N_12080);
or UO_576 (O_576,N_12312,N_12775);
and UO_577 (O_577,N_13087,N_12742);
nand UO_578 (O_578,N_13110,N_13882);
or UO_579 (O_579,N_12686,N_14644);
or UO_580 (O_580,N_13434,N_12756);
or UO_581 (O_581,N_13041,N_14287);
nand UO_582 (O_582,N_12464,N_13356);
nor UO_583 (O_583,N_12865,N_14994);
nor UO_584 (O_584,N_14811,N_12382);
and UO_585 (O_585,N_12554,N_12067);
and UO_586 (O_586,N_12441,N_14973);
and UO_587 (O_587,N_12735,N_14036);
nor UO_588 (O_588,N_12388,N_13827);
or UO_589 (O_589,N_12126,N_12049);
and UO_590 (O_590,N_12171,N_13369);
xor UO_591 (O_591,N_13242,N_12701);
or UO_592 (O_592,N_14615,N_14404);
or UO_593 (O_593,N_12223,N_13257);
nor UO_594 (O_594,N_12868,N_14802);
nand UO_595 (O_595,N_14641,N_13156);
nor UO_596 (O_596,N_13161,N_13171);
nand UO_597 (O_597,N_13596,N_13277);
and UO_598 (O_598,N_13143,N_14148);
nand UO_599 (O_599,N_12708,N_12160);
nand UO_600 (O_600,N_12356,N_14622);
xnor UO_601 (O_601,N_12509,N_12527);
and UO_602 (O_602,N_12238,N_13227);
or UO_603 (O_603,N_12653,N_13045);
nand UO_604 (O_604,N_13563,N_12462);
nor UO_605 (O_605,N_13803,N_14747);
and UO_606 (O_606,N_14722,N_12111);
nand UO_607 (O_607,N_14799,N_13617);
xnor UO_608 (O_608,N_13656,N_12803);
nand UO_609 (O_609,N_14256,N_14840);
nand UO_610 (O_610,N_12792,N_12809);
xor UO_611 (O_611,N_14961,N_13645);
or UO_612 (O_612,N_12007,N_13264);
nor UO_613 (O_613,N_12134,N_12645);
xor UO_614 (O_614,N_12758,N_12084);
nor UO_615 (O_615,N_14352,N_12131);
xnor UO_616 (O_616,N_12692,N_14065);
nor UO_617 (O_617,N_12744,N_12280);
xor UO_618 (O_618,N_13883,N_12037);
or UO_619 (O_619,N_12268,N_13350);
nand UO_620 (O_620,N_14126,N_13347);
nor UO_621 (O_621,N_13919,N_14638);
or UO_622 (O_622,N_14787,N_12778);
or UO_623 (O_623,N_13099,N_13538);
nor UO_624 (O_624,N_14383,N_12570);
nand UO_625 (O_625,N_13429,N_12690);
or UO_626 (O_626,N_12324,N_13528);
or UO_627 (O_627,N_14454,N_14918);
nor UO_628 (O_628,N_14142,N_14362);
nand UO_629 (O_629,N_12658,N_14793);
and UO_630 (O_630,N_13180,N_14495);
nand UO_631 (O_631,N_13817,N_12636);
and UO_632 (O_632,N_12436,N_12013);
and UO_633 (O_633,N_13456,N_14785);
nand UO_634 (O_634,N_13871,N_12881);
nand UO_635 (O_635,N_13710,N_12471);
and UO_636 (O_636,N_14726,N_12833);
xnor UO_637 (O_637,N_12813,N_13370);
nor UO_638 (O_638,N_12786,N_14216);
nor UO_639 (O_639,N_14219,N_12113);
nor UO_640 (O_640,N_14953,N_13676);
nor UO_641 (O_641,N_12147,N_13130);
nor UO_642 (O_642,N_14764,N_14184);
nor UO_643 (O_643,N_14922,N_13049);
and UO_644 (O_644,N_13463,N_13543);
nor UO_645 (O_645,N_14891,N_14040);
or UO_646 (O_646,N_12346,N_14232);
xor UO_647 (O_647,N_13328,N_14253);
or UO_648 (O_648,N_14364,N_13562);
nand UO_649 (O_649,N_12501,N_14734);
nor UO_650 (O_650,N_12673,N_14422);
nor UO_651 (O_651,N_14403,N_12380);
nor UO_652 (O_652,N_13428,N_14703);
nor UO_653 (O_653,N_14262,N_13586);
xnor UO_654 (O_654,N_13152,N_14446);
nor UO_655 (O_655,N_12381,N_12528);
nand UO_656 (O_656,N_12409,N_14448);
nand UO_657 (O_657,N_13084,N_14859);
xnor UO_658 (O_658,N_13299,N_14468);
xnor UO_659 (O_659,N_12056,N_13579);
or UO_660 (O_660,N_13092,N_14829);
xor UO_661 (O_661,N_14902,N_14125);
and UO_662 (O_662,N_14320,N_12394);
nand UO_663 (O_663,N_12713,N_13760);
xnor UO_664 (O_664,N_12121,N_12062);
or UO_665 (O_665,N_14652,N_14914);
or UO_666 (O_666,N_14343,N_14904);
or UO_667 (O_667,N_13807,N_13674);
and UO_668 (O_668,N_14718,N_13995);
and UO_669 (O_669,N_13358,N_14597);
nor UO_670 (O_670,N_12391,N_13085);
nor UO_671 (O_671,N_13201,N_14882);
xor UO_672 (O_672,N_14780,N_14887);
nand UO_673 (O_673,N_13502,N_13984);
xor UO_674 (O_674,N_14419,N_12262);
nor UO_675 (O_675,N_13317,N_14100);
or UO_676 (O_676,N_14689,N_12194);
nand UO_677 (O_677,N_12958,N_12142);
and UO_678 (O_678,N_13490,N_12598);
nor UO_679 (O_679,N_13846,N_14405);
or UO_680 (O_680,N_14676,N_14655);
nor UO_681 (O_681,N_13449,N_14593);
xor UO_682 (O_682,N_14988,N_13713);
or UO_683 (O_683,N_14478,N_12760);
and UO_684 (O_684,N_14626,N_12296);
nor UO_685 (O_685,N_12579,N_14583);
nand UO_686 (O_686,N_13117,N_13163);
and UO_687 (O_687,N_13241,N_14390);
nor UO_688 (O_688,N_14206,N_12748);
nand UO_689 (O_689,N_12908,N_12431);
nand UO_690 (O_690,N_12124,N_14733);
nor UO_691 (O_691,N_13734,N_12046);
nand UO_692 (O_692,N_13872,N_12205);
or UO_693 (O_693,N_12601,N_12696);
nor UO_694 (O_694,N_14317,N_12541);
or UO_695 (O_695,N_12249,N_14512);
nand UO_696 (O_696,N_14156,N_13425);
and UO_697 (O_697,N_12000,N_13336);
xnor UO_698 (O_698,N_14043,N_12333);
and UO_699 (O_699,N_14123,N_14203);
or UO_700 (O_700,N_12362,N_14138);
or UO_701 (O_701,N_14437,N_14371);
nor UO_702 (O_702,N_14947,N_12211);
nor UO_703 (O_703,N_14878,N_14723);
or UO_704 (O_704,N_13232,N_12207);
nor UO_705 (O_705,N_14579,N_12683);
or UO_706 (O_706,N_14247,N_12363);
nor UO_707 (O_707,N_13047,N_14384);
and UO_708 (O_708,N_12921,N_13107);
and UO_709 (O_709,N_14814,N_14905);
or UO_710 (O_710,N_14304,N_12323);
nand UO_711 (O_711,N_14795,N_14292);
nand UO_712 (O_712,N_13588,N_12542);
nor UO_713 (O_713,N_14323,N_14177);
or UO_714 (O_714,N_12615,N_12726);
or UO_715 (O_715,N_12884,N_14805);
xor UO_716 (O_716,N_14821,N_14147);
nand UO_717 (O_717,N_14176,N_13781);
nand UO_718 (O_718,N_12407,N_12625);
or UO_719 (O_719,N_12239,N_12932);
and UO_720 (O_720,N_14794,N_14026);
and UO_721 (O_721,N_14555,N_12539);
or UO_722 (O_722,N_14489,N_14420);
and UO_723 (O_723,N_14760,N_12848);
nor UO_724 (O_724,N_12433,N_14608);
or UO_725 (O_725,N_14586,N_12750);
and UO_726 (O_726,N_12326,N_14704);
or UO_727 (O_727,N_12580,N_13999);
or UO_728 (O_728,N_12825,N_14186);
and UO_729 (O_729,N_12281,N_13255);
xnor UO_730 (O_730,N_12842,N_14346);
and UO_731 (O_731,N_14116,N_14842);
or UO_732 (O_732,N_13594,N_14609);
and UO_733 (O_733,N_12896,N_13506);
or UO_734 (O_734,N_14127,N_13912);
nand UO_735 (O_735,N_13438,N_12273);
xnor UO_736 (O_736,N_14046,N_13330);
or UO_737 (O_737,N_14737,N_12854);
and UO_738 (O_738,N_14845,N_14874);
or UO_739 (O_739,N_14377,N_12682);
nand UO_740 (O_740,N_12789,N_14254);
or UO_741 (O_741,N_14011,N_12192);
nand UO_742 (O_742,N_13514,N_14175);
nand UO_743 (O_743,N_13185,N_14271);
and UO_744 (O_744,N_12985,N_12836);
xnor UO_745 (O_745,N_12595,N_14319);
or UO_746 (O_746,N_12216,N_12220);
and UO_747 (O_747,N_14756,N_13031);
nand UO_748 (O_748,N_12785,N_12318);
and UO_749 (O_749,N_14386,N_12174);
or UO_750 (O_750,N_12073,N_14589);
xor UO_751 (O_751,N_14063,N_12191);
nand UO_752 (O_752,N_14128,N_14710);
and UO_753 (O_753,N_13214,N_13869);
xor UO_754 (O_754,N_12643,N_12805);
nand UO_755 (O_755,N_14109,N_13763);
nor UO_756 (O_756,N_13172,N_13892);
nor UO_757 (O_757,N_14667,N_14288);
and UO_758 (O_758,N_12518,N_14460);
and UO_759 (O_759,N_12507,N_13918);
or UO_760 (O_760,N_13189,N_14321);
and UO_761 (O_761,N_13545,N_12669);
or UO_762 (O_762,N_13372,N_14928);
and UO_763 (O_763,N_13091,N_12133);
nor UO_764 (O_764,N_12609,N_14104);
and UO_765 (O_765,N_13427,N_12707);
nand UO_766 (O_766,N_13058,N_13887);
or UO_767 (O_767,N_12892,N_13164);
or UO_768 (O_768,N_12102,N_12782);
nor UO_769 (O_769,N_12028,N_12727);
nand UO_770 (O_770,N_14165,N_12148);
or UO_771 (O_771,N_13139,N_12752);
nand UO_772 (O_772,N_13836,N_13841);
or UO_773 (O_773,N_12345,N_14060);
or UO_774 (O_774,N_13886,N_13480);
or UO_775 (O_775,N_12190,N_14334);
nor UO_776 (O_776,N_14530,N_14907);
and UO_777 (O_777,N_14591,N_13196);
or UO_778 (O_778,N_12330,N_13659);
and UO_779 (O_779,N_13050,N_12998);
and UO_780 (O_780,N_14529,N_14400);
or UO_781 (O_781,N_12720,N_14774);
and UO_782 (O_782,N_13648,N_13641);
or UO_783 (O_783,N_13508,N_13582);
and UO_784 (O_784,N_14169,N_13935);
or UO_785 (O_785,N_14757,N_14195);
nor UO_786 (O_786,N_13859,N_14037);
nand UO_787 (O_787,N_13479,N_14498);
nand UO_788 (O_788,N_12567,N_14542);
xor UO_789 (O_789,N_13922,N_14754);
or UO_790 (O_790,N_13772,N_12097);
nor UO_791 (O_791,N_14818,N_12614);
xnor UO_792 (O_792,N_12586,N_14315);
or UO_793 (O_793,N_14286,N_13411);
and UO_794 (O_794,N_13073,N_14744);
and UO_795 (O_795,N_12656,N_13046);
nand UO_796 (O_796,N_14665,N_14250);
nand UO_797 (O_797,N_14937,N_12396);
nand UO_798 (O_798,N_14112,N_13132);
nand UO_799 (O_799,N_12291,N_14409);
nand UO_800 (O_800,N_12648,N_13696);
nand UO_801 (O_801,N_13395,N_12557);
nor UO_802 (O_802,N_12450,N_14752);
nand UO_803 (O_803,N_12334,N_13158);
nor UO_804 (O_804,N_12299,N_14995);
nand UO_805 (O_805,N_12602,N_14014);
and UO_806 (O_806,N_13530,N_14523);
nand UO_807 (O_807,N_13461,N_12583);
or UO_808 (O_808,N_14340,N_12397);
or UO_809 (O_809,N_13898,N_14496);
and UO_810 (O_810,N_14967,N_12491);
nand UO_811 (O_811,N_12361,N_12011);
nor UO_812 (O_812,N_12448,N_14149);
nor UO_813 (O_813,N_13909,N_14957);
and UO_814 (O_814,N_12926,N_14585);
nand UO_815 (O_815,N_12271,N_12108);
nand UO_816 (O_816,N_12384,N_12969);
xnor UO_817 (O_817,N_14055,N_13222);
xor UO_818 (O_818,N_13833,N_13315);
and UO_819 (O_819,N_13155,N_13441);
nand UO_820 (O_820,N_14969,N_14801);
nand UO_821 (O_821,N_14876,N_14438);
xnor UO_822 (O_822,N_13660,N_13295);
xnor UO_823 (O_823,N_14136,N_14610);
or UO_824 (O_824,N_14771,N_13574);
nand UO_825 (O_825,N_12168,N_12763);
or UO_826 (O_826,N_13782,N_13753);
or UO_827 (O_827,N_14706,N_14486);
nor UO_828 (O_828,N_12365,N_12089);
or UO_829 (O_829,N_12674,N_14506);
and UO_830 (O_830,N_14834,N_13896);
nand UO_831 (O_831,N_13236,N_12165);
or UO_832 (O_832,N_12289,N_12655);
nand UO_833 (O_833,N_14096,N_14434);
and UO_834 (O_834,N_14456,N_14435);
nor UO_835 (O_835,N_13199,N_14578);
and UO_836 (O_836,N_14105,N_12427);
or UO_837 (O_837,N_14067,N_12311);
nand UO_838 (O_838,N_14908,N_12774);
and UO_839 (O_839,N_14525,N_12678);
and UO_840 (O_840,N_12081,N_13555);
and UO_841 (O_841,N_12956,N_14869);
nand UO_842 (O_842,N_14521,N_12458);
and UO_843 (O_843,N_13403,N_12589);
or UO_844 (O_844,N_14651,N_14848);
xnor UO_845 (O_845,N_14284,N_14535);
nand UO_846 (O_846,N_12818,N_12474);
nand UO_847 (O_847,N_12962,N_12694);
nor UO_848 (O_848,N_13374,N_13233);
nand UO_849 (O_849,N_14085,N_13129);
or UO_850 (O_850,N_12116,N_13724);
xor UO_851 (O_851,N_12558,N_13090);
nor UO_852 (O_852,N_13322,N_12272);
and UO_853 (O_853,N_14549,N_12955);
nand UO_854 (O_854,N_14114,N_12839);
nor UO_855 (O_855,N_13941,N_14487);
xnor UO_856 (O_856,N_12297,N_14407);
xor UO_857 (O_857,N_14092,N_12628);
or UO_858 (O_858,N_14015,N_14738);
nand UO_859 (O_859,N_13020,N_12521);
nand UO_860 (O_860,N_14730,N_13801);
xnor UO_861 (O_861,N_13297,N_14741);
and UO_862 (O_862,N_14480,N_12667);
or UO_863 (O_863,N_13540,N_12941);
and UO_864 (O_864,N_12613,N_12879);
nor UO_865 (O_865,N_12144,N_13519);
or UO_866 (O_866,N_14210,N_13754);
nor UO_867 (O_867,N_14870,N_12267);
nand UO_868 (O_868,N_13743,N_14281);
nor UO_869 (O_869,N_13736,N_13962);
nor UO_870 (O_870,N_13452,N_13262);
and UO_871 (O_871,N_12401,N_12150);
and UO_872 (O_872,N_12074,N_13209);
and UO_873 (O_873,N_14517,N_14077);
nor UO_874 (O_874,N_14697,N_13281);
nand UO_875 (O_875,N_12243,N_13343);
nand UO_876 (O_876,N_12925,N_13975);
and UO_877 (O_877,N_12576,N_12379);
nand UO_878 (O_878,N_14654,N_12986);
nor UO_879 (O_879,N_13698,N_12039);
nor UO_880 (O_880,N_13866,N_12914);
xor UO_881 (O_881,N_14779,N_13885);
xor UO_882 (O_882,N_13497,N_13673);
or UO_883 (O_883,N_12953,N_12112);
nor UO_884 (O_884,N_13686,N_14394);
and UO_885 (O_885,N_13573,N_12738);
nand UO_886 (O_886,N_12132,N_12523);
nand UO_887 (O_887,N_14279,N_13654);
or UO_888 (O_888,N_12736,N_12449);
nor UO_889 (O_889,N_14896,N_14447);
nand UO_890 (O_890,N_12483,N_13571);
and UO_891 (O_891,N_14604,N_12416);
and UO_892 (O_892,N_13167,N_13025);
xor UO_893 (O_893,N_12065,N_14690);
or UO_894 (O_894,N_13966,N_14172);
nand UO_895 (O_895,N_12698,N_14745);
or UO_896 (O_896,N_12045,N_14084);
or UO_897 (O_897,N_13454,N_12820);
nor UO_898 (O_898,N_12350,N_14510);
nor UO_899 (O_899,N_14179,N_14260);
nand UO_900 (O_900,N_13298,N_12711);
and UO_901 (O_901,N_13927,N_14310);
and UO_902 (O_902,N_14777,N_14646);
nand UO_903 (O_903,N_14481,N_14255);
xnor UO_904 (O_904,N_12900,N_14564);
and UO_905 (O_905,N_12314,N_12016);
xor UO_906 (O_906,N_12402,N_14035);
nor UO_907 (O_907,N_13766,N_12536);
or UO_908 (O_908,N_13188,N_13592);
or UO_909 (O_909,N_14558,N_12952);
nand UO_910 (O_910,N_13348,N_13806);
or UO_911 (O_911,N_14444,N_13814);
and UO_912 (O_912,N_14879,N_13444);
and UO_913 (O_913,N_12918,N_14443);
and UO_914 (O_914,N_14716,N_13539);
and UO_915 (O_915,N_13062,N_13442);
and UO_916 (O_916,N_12320,N_14694);
and UO_917 (O_917,N_14582,N_14052);
nand UO_918 (O_918,N_13378,N_14674);
nand UO_919 (O_919,N_14941,N_12455);
or UO_920 (O_920,N_13492,N_14066);
nor UO_921 (O_921,N_14283,N_12859);
nand UO_922 (O_922,N_13722,N_14355);
nor UO_923 (O_923,N_14243,N_14866);
or UO_924 (O_924,N_14411,N_13794);
and UO_925 (O_925,N_12136,N_12094);
nand UO_926 (O_926,N_14501,N_13985);
or UO_927 (O_927,N_13776,N_14964);
and UO_928 (O_928,N_13389,N_13024);
and UO_929 (O_929,N_12999,N_14032);
nor UO_930 (O_930,N_12544,N_13448);
xnor UO_931 (O_931,N_12260,N_13529);
xor UO_932 (O_932,N_12661,N_13146);
nand UO_933 (O_933,N_12153,N_12274);
nor UO_934 (O_934,N_14949,N_12723);
and UO_935 (O_935,N_12759,N_13309);
and UO_936 (O_936,N_14196,N_14580);
nor UO_937 (O_937,N_13979,N_14204);
or UO_938 (O_938,N_13145,N_14475);
xnor UO_939 (O_939,N_14494,N_13200);
nor UO_940 (O_940,N_14664,N_12934);
nor UO_941 (O_941,N_13120,N_14483);
nor UO_942 (O_942,N_13575,N_14836);
xnor UO_943 (O_943,N_14473,N_14053);
and UO_944 (O_944,N_12706,N_13509);
nor UO_945 (O_945,N_13679,N_14790);
nor UO_946 (O_946,N_13829,N_12937);
or UO_947 (O_947,N_13634,N_13306);
or UO_948 (O_948,N_13992,N_14111);
nor UO_949 (O_949,N_13054,N_13269);
nand UO_950 (O_950,N_13825,N_14406);
nand UO_951 (O_951,N_12959,N_14345);
nand UO_952 (O_952,N_12978,N_12390);
and UO_953 (O_953,N_12743,N_12221);
or UO_954 (O_954,N_13577,N_14611);
nand UO_955 (O_955,N_12883,N_12063);
nor UO_956 (O_956,N_12470,N_13407);
or UO_957 (O_957,N_12119,N_14192);
or UO_958 (O_958,N_14171,N_12231);
or UO_959 (O_959,N_13268,N_13811);
or UO_960 (O_960,N_14960,N_14629);
and UO_961 (O_961,N_13773,N_14191);
nor UO_962 (O_962,N_13183,N_12632);
and UO_963 (O_963,N_14293,N_12479);
and UO_964 (O_964,N_12512,N_14721);
and UO_965 (O_965,N_14559,N_13796);
nand UO_966 (O_966,N_13329,N_12287);
nor UO_967 (O_967,N_14103,N_14762);
and UO_968 (O_968,N_12534,N_13861);
or UO_969 (O_969,N_14153,N_14600);
nor UO_970 (O_970,N_12473,N_14675);
and UO_971 (O_971,N_13194,N_12492);
nand UO_972 (O_972,N_13433,N_13323);
nand UO_973 (O_973,N_12715,N_12794);
xnor UO_974 (O_974,N_14129,N_12054);
nor UO_975 (O_975,N_13680,N_14075);
nor UO_976 (O_976,N_13181,N_13637);
and UO_977 (O_977,N_14050,N_12930);
or UO_978 (O_978,N_13810,N_13792);
and UO_979 (O_979,N_13791,N_13420);
nor UO_980 (O_980,N_12939,N_13252);
nor UO_981 (O_981,N_14679,N_14827);
and UO_982 (O_982,N_12057,N_13482);
nor UO_983 (O_983,N_14659,N_13976);
nand UO_984 (O_984,N_14091,N_14871);
and UO_985 (O_985,N_14940,N_13533);
xnor UO_986 (O_986,N_13837,N_14229);
and UO_987 (O_987,N_12592,N_14021);
xnor UO_988 (O_988,N_13691,N_13101);
and UO_989 (O_989,N_14162,N_13844);
and UO_990 (O_990,N_12834,N_14758);
nand UO_991 (O_991,N_14024,N_12652);
nor UO_992 (O_992,N_14482,N_12765);
nand UO_993 (O_993,N_12991,N_14770);
xor UO_994 (O_994,N_12984,N_14003);
or UO_995 (O_995,N_12927,N_14606);
nor UO_996 (O_996,N_12942,N_13646);
and UO_997 (O_997,N_14006,N_12259);
and UO_998 (O_998,N_13601,N_12222);
or UO_999 (O_999,N_13135,N_14596);
nand UO_1000 (O_1000,N_12849,N_13572);
nand UO_1001 (O_1001,N_13876,N_12035);
and UO_1002 (O_1002,N_14672,N_14663);
or UO_1003 (O_1003,N_14956,N_12864);
or UO_1004 (O_1004,N_12313,N_14696);
nand UO_1005 (O_1005,N_14058,N_13498);
nor UO_1006 (O_1006,N_13756,N_13847);
xor UO_1007 (O_1007,N_13357,N_13953);
or UO_1008 (O_1008,N_13993,N_12228);
nor UO_1009 (O_1009,N_13643,N_13097);
and UO_1010 (O_1010,N_12847,N_14557);
or UO_1011 (O_1011,N_12829,N_13042);
or UO_1012 (O_1012,N_12332,N_13867);
nand UO_1013 (O_1013,N_12967,N_12564);
and UO_1014 (O_1014,N_14161,N_14977);
or UO_1015 (O_1015,N_13798,N_12890);
nor UO_1016 (O_1016,N_14786,N_12251);
nor UO_1017 (O_1017,N_14511,N_13326);
xor UO_1018 (O_1018,N_13780,N_14920);
xnor UO_1019 (O_1019,N_14466,N_13531);
or UO_1020 (O_1020,N_14298,N_14860);
and UO_1021 (O_1021,N_13752,N_14900);
nand UO_1022 (O_1022,N_13018,N_14391);
nor UO_1023 (O_1023,N_12665,N_13293);
nor UO_1024 (O_1024,N_13244,N_13391);
nor UO_1025 (O_1025,N_13623,N_12355);
nor UO_1026 (O_1026,N_12800,N_14433);
nand UO_1027 (O_1027,N_12629,N_12234);
nor UO_1028 (O_1028,N_12928,N_14625);
and UO_1029 (O_1029,N_13280,N_13532);
and UO_1030 (O_1030,N_14749,N_12931);
or UO_1031 (O_1031,N_12563,N_12166);
or UO_1032 (O_1032,N_12376,N_14418);
xor UO_1033 (O_1033,N_13302,N_12303);
and UO_1034 (O_1034,N_13153,N_14849);
or UO_1035 (O_1035,N_13997,N_13119);
and UO_1036 (O_1036,N_14408,N_12090);
nor UO_1037 (O_1037,N_12224,N_14005);
nor UO_1038 (O_1038,N_13626,N_14335);
nor UO_1039 (O_1039,N_12851,N_13824);
nor UO_1040 (O_1040,N_12547,N_14294);
nand UO_1041 (O_1041,N_13016,N_13560);
xor UO_1042 (O_1042,N_12869,N_12560);
nand UO_1043 (O_1043,N_12830,N_14458);
nand UO_1044 (O_1044,N_14946,N_13088);
and UO_1045 (O_1045,N_12098,N_12051);
nor UO_1046 (O_1046,N_13022,N_12993);
nor UO_1047 (O_1047,N_12787,N_12717);
nand UO_1048 (O_1048,N_14235,N_12526);
nor UO_1049 (O_1049,N_12783,N_14209);
or UO_1050 (O_1050,N_14561,N_14396);
or UO_1051 (O_1051,N_13423,N_14938);
and UO_1052 (O_1052,N_14380,N_14810);
nor UO_1053 (O_1053,N_14358,N_12912);
xnor UO_1054 (O_1054,N_12766,N_13828);
or UO_1055 (O_1055,N_14382,N_12647);
nand UO_1056 (O_1056,N_12821,N_13140);
nand UO_1057 (O_1057,N_14543,N_13991);
nand UO_1058 (O_1058,N_14824,N_13468);
nand UO_1059 (O_1059,N_13725,N_13033);
nand UO_1060 (O_1060,N_13537,N_12838);
nand UO_1061 (O_1061,N_12004,N_12290);
nor UO_1062 (O_1062,N_12604,N_13587);
nand UO_1063 (O_1063,N_12270,N_12213);
or UO_1064 (O_1064,N_14992,N_12184);
nand UO_1065 (O_1065,N_14341,N_14642);
xnor UO_1066 (O_1066,N_13154,N_13366);
nor UO_1067 (O_1067,N_14954,N_13853);
nand UO_1068 (O_1068,N_14677,N_14163);
xor UO_1069 (O_1069,N_12549,N_12790);
nand UO_1070 (O_1070,N_13988,N_13061);
nand UO_1071 (O_1071,N_14228,N_12058);
or UO_1072 (O_1072,N_14455,N_13739);
nor UO_1073 (O_1073,N_14312,N_14121);
nand UO_1074 (O_1074,N_14963,N_12055);
xor UO_1075 (O_1075,N_13907,N_13160);
and UO_1076 (O_1076,N_14471,N_12714);
nor UO_1077 (O_1077,N_14532,N_12023);
nand UO_1078 (O_1078,N_14093,N_12099);
nor UO_1079 (O_1079,N_12214,N_13661);
nand UO_1080 (O_1080,N_12398,N_14854);
nand UO_1081 (O_1081,N_13924,N_12870);
or UO_1082 (O_1082,N_12354,N_12951);
nand UO_1083 (O_1083,N_13908,N_13436);
nor UO_1084 (O_1084,N_13541,N_13355);
nor UO_1085 (O_1085,N_12316,N_13553);
xor UO_1086 (O_1086,N_14297,N_14441);
nand UO_1087 (O_1087,N_13324,N_13060);
and UO_1088 (O_1088,N_14266,N_13933);
nand UO_1089 (O_1089,N_12974,N_12443);
nor UO_1090 (O_1090,N_14571,N_12064);
xor UO_1091 (O_1091,N_13627,N_12319);
nand UO_1092 (O_1092,N_13312,N_14996);
xor UO_1093 (O_1093,N_13789,N_12006);
nand UO_1094 (O_1094,N_14537,N_14798);
or UO_1095 (O_1095,N_12712,N_14155);
or UO_1096 (O_1096,N_14350,N_12487);
and UO_1097 (O_1097,N_13714,N_13704);
and UO_1098 (O_1098,N_13938,N_13170);
nor UO_1099 (O_1099,N_14778,N_13816);
xor UO_1100 (O_1100,N_12245,N_12170);
or UO_1101 (O_1101,N_12258,N_13556);
nand UO_1102 (O_1102,N_14566,N_14680);
or UO_1103 (O_1103,N_14708,N_14980);
and UO_1104 (O_1104,N_12902,N_13749);
or UO_1105 (O_1105,N_13716,N_14120);
nor UO_1106 (O_1106,N_13874,N_13595);
nand UO_1107 (O_1107,N_13702,N_13121);
nand UO_1108 (O_1108,N_12444,N_13106);
nand UO_1109 (O_1109,N_13826,N_14912);
or UO_1110 (O_1110,N_13520,N_13717);
nor UO_1111 (O_1111,N_12502,N_13240);
or UO_1112 (O_1112,N_14160,N_12375);
and UO_1113 (O_1113,N_14825,N_14425);
nand UO_1114 (O_1114,N_12425,N_13177);
nand UO_1115 (O_1115,N_13481,N_12242);
xnor UO_1116 (O_1116,N_13215,N_12499);
and UO_1117 (O_1117,N_12069,N_14524);
nor UO_1118 (O_1118,N_13095,N_12233);
and UO_1119 (O_1119,N_14560,N_13747);
nand UO_1120 (O_1120,N_14599,N_14102);
or UO_1121 (O_1121,N_13503,N_14673);
nand UO_1122 (O_1122,N_13250,N_13709);
and UO_1123 (O_1123,N_13096,N_12456);
or UO_1124 (O_1124,N_14025,N_13715);
and UO_1125 (O_1125,N_14325,N_13224);
and UO_1126 (O_1126,N_14459,N_12606);
xor UO_1127 (O_1127,N_14839,N_14453);
nand UO_1128 (O_1128,N_12695,N_14826);
or UO_1129 (O_1129,N_13418,N_14736);
nor UO_1130 (O_1130,N_12954,N_14258);
nand UO_1131 (O_1131,N_12250,N_14339);
nand UO_1132 (O_1132,N_14910,N_13638);
xnor UO_1133 (O_1133,N_12040,N_14207);
or UO_1134 (O_1134,N_12960,N_14360);
and UO_1135 (O_1135,N_14899,N_12301);
nand UO_1136 (O_1136,N_14002,N_13340);
xnor UO_1137 (O_1137,N_12898,N_14431);
or UO_1138 (O_1138,N_13245,N_13394);
nand UO_1139 (O_1139,N_14387,N_14042);
nand UO_1140 (O_1140,N_14076,N_13544);
xor UO_1141 (O_1141,N_13672,N_12459);
nor UO_1142 (O_1142,N_12889,N_14630);
xnor UO_1143 (O_1143,N_13229,N_12718);
and UO_1144 (O_1144,N_12393,N_12762);
and UO_1145 (O_1145,N_12538,N_12596);
or UO_1146 (O_1146,N_12202,N_13017);
or UO_1147 (O_1147,N_13086,N_12909);
nand UO_1148 (O_1148,N_12226,N_14236);
nor UO_1149 (O_1149,N_14423,N_13851);
and UO_1150 (O_1150,N_12236,N_12886);
nand UO_1151 (O_1151,N_14041,N_14398);
or UO_1152 (O_1152,N_13554,N_14023);
and UO_1153 (O_1153,N_13125,N_13210);
and UO_1154 (O_1154,N_12284,N_13430);
xor UO_1155 (O_1155,N_13735,N_12945);
nor UO_1156 (O_1156,N_13510,N_14452);
or UO_1157 (O_1157,N_14519,N_14363);
and UO_1158 (O_1158,N_14671,N_14133);
and UO_1159 (O_1159,N_12751,N_14753);
or UO_1160 (O_1160,N_14643,N_14493);
nor UO_1161 (O_1161,N_14244,N_14815);
and UO_1162 (O_1162,N_12697,N_13965);
and UO_1163 (O_1163,N_14623,N_13417);
or UO_1164 (O_1164,N_12573,N_13310);
or UO_1165 (O_1165,N_14819,N_13267);
xnor UO_1166 (O_1166,N_13865,N_12476);
xor UO_1167 (O_1167,N_12387,N_13835);
or UO_1168 (O_1168,N_13925,N_12408);
nor UO_1169 (O_1169,N_14605,N_14305);
or UO_1170 (O_1170,N_14154,N_13078);
nor UO_1171 (O_1171,N_14955,N_12913);
nor UO_1172 (O_1172,N_14373,N_14068);
and UO_1173 (O_1173,N_14636,N_14812);
nor UO_1174 (O_1174,N_14193,N_13957);
or UO_1175 (O_1175,N_13331,N_13475);
or UO_1176 (O_1176,N_14551,N_13459);
or UO_1177 (O_1177,N_13548,N_13076);
nand UO_1178 (O_1178,N_14850,N_13124);
nor UO_1179 (O_1179,N_12036,N_12844);
nor UO_1180 (O_1180,N_12850,N_14804);
xnor UO_1181 (O_1181,N_13959,N_12347);
nand UO_1182 (O_1182,N_13260,N_13259);
or UO_1183 (O_1183,N_12722,N_14146);
nor UO_1184 (O_1184,N_13765,N_13012);
nand UO_1185 (O_1185,N_12525,N_14295);
nor UO_1186 (O_1186,N_13644,N_14233);
xnor UO_1187 (O_1187,N_14259,N_12575);
or UO_1188 (O_1188,N_12423,N_12139);
nor UO_1189 (O_1189,N_13884,N_13758);
and UO_1190 (O_1190,N_14379,N_13216);
or UO_1191 (O_1191,N_14263,N_12703);
nor UO_1192 (O_1192,N_13070,N_12358);
nor UO_1193 (O_1193,N_13726,N_12565);
nor UO_1194 (O_1194,N_12229,N_13362);
nor UO_1195 (O_1195,N_12095,N_12032);
and UO_1196 (O_1196,N_13516,N_12357);
nor UO_1197 (O_1197,N_13360,N_13218);
nor UO_1198 (O_1198,N_14047,N_13721);
nor UO_1199 (O_1199,N_12767,N_12524);
or UO_1200 (O_1200,N_13955,N_13757);
and UO_1201 (O_1201,N_13457,N_13740);
nor UO_1202 (O_1202,N_13006,N_12294);
and UO_1203 (O_1203,N_13009,N_14490);
or UO_1204 (O_1204,N_13585,N_13168);
nand UO_1205 (O_1205,N_13023,N_14000);
nor UO_1206 (O_1206,N_13632,N_12568);
nand UO_1207 (O_1207,N_13839,N_12679);
nand UO_1208 (O_1208,N_13111,N_12295);
and UO_1209 (O_1209,N_14151,N_14514);
nor UO_1210 (O_1210,N_12118,N_14766);
nor UO_1211 (O_1211,N_12477,N_12943);
xor UO_1212 (O_1212,N_12582,N_14389);
nor UO_1213 (O_1213,N_12824,N_13021);
xnor UO_1214 (O_1214,N_13779,N_12841);
xnor UO_1215 (O_1215,N_14911,N_13304);
nor UO_1216 (O_1216,N_12072,N_14265);
nor UO_1217 (O_1217,N_14356,N_14531);
or UO_1218 (O_1218,N_14117,N_13279);
nand UO_1219 (O_1219,N_14421,N_12158);
nor UO_1220 (O_1220,N_13212,N_13928);
or UO_1221 (O_1221,N_13694,N_13805);
nor UO_1222 (O_1222,N_14083,N_14890);
and UO_1223 (O_1223,N_13159,N_13650);
nor UO_1224 (O_1224,N_13665,N_14661);
nor UO_1225 (O_1225,N_13287,N_14867);
nor UO_1226 (O_1226,N_13337,N_14847);
or UO_1227 (O_1227,N_13767,N_12855);
or UO_1228 (O_1228,N_14012,N_14090);
nand UO_1229 (O_1229,N_14347,N_14616);
nand UO_1230 (O_1230,N_14844,N_14074);
nor UO_1231 (O_1231,N_12840,N_14211);
and UO_1232 (O_1232,N_13142,N_14463);
nor UO_1233 (O_1233,N_14864,N_14030);
nor UO_1234 (O_1234,N_14289,N_13104);
nor UO_1235 (O_1235,N_13462,N_12641);
and UO_1236 (O_1236,N_14881,N_13325);
and UO_1237 (O_1237,N_13276,N_12152);
xor UO_1238 (O_1238,N_13956,N_12434);
or UO_1239 (O_1239,N_14502,N_12511);
nand UO_1240 (O_1240,N_13642,N_14808);
or UO_1241 (O_1241,N_12510,N_14401);
and UO_1242 (O_1242,N_13354,N_14574);
nor UO_1243 (O_1243,N_13342,N_13314);
xor UO_1244 (O_1244,N_13179,N_12671);
nor UO_1245 (O_1245,N_12253,N_12420);
nand UO_1246 (O_1246,N_12590,N_14508);
or UO_1247 (O_1247,N_14687,N_12015);
nand UO_1248 (O_1248,N_12901,N_14173);
nand UO_1249 (O_1249,N_12378,N_12275);
nand UO_1250 (O_1250,N_12872,N_13904);
nand UO_1251 (O_1251,N_14034,N_13895);
nand UO_1252 (O_1252,N_13150,N_12412);
and UO_1253 (O_1253,N_13755,N_13093);
nand UO_1254 (O_1254,N_12130,N_13605);
or UO_1255 (O_1255,N_12044,N_13770);
and UO_1256 (O_1256,N_14237,N_14547);
nand UO_1257 (O_1257,N_13476,N_14218);
and UO_1258 (O_1258,N_12976,N_12876);
nand UO_1259 (O_1259,N_14119,N_12906);
and UO_1260 (O_1260,N_12732,N_12734);
nor UO_1261 (O_1261,N_13890,N_13681);
nor UO_1262 (O_1262,N_13675,N_13769);
and UO_1263 (O_1263,N_12893,N_14361);
xor UO_1264 (O_1264,N_14188,N_12552);
or UO_1265 (O_1265,N_12529,N_13493);
and UO_1266 (O_1266,N_12179,N_13584);
or UO_1267 (O_1267,N_13103,N_12970);
or UO_1268 (O_1268,N_13238,N_14048);
and UO_1269 (O_1269,N_12755,N_13952);
nor UO_1270 (O_1270,N_14699,N_13377);
or UO_1271 (O_1271,N_14948,N_13940);
nand UO_1272 (O_1272,N_13015,N_14546);
and UO_1273 (O_1273,N_14507,N_14883);
nand UO_1274 (O_1274,N_13118,N_13294);
nand UO_1275 (O_1275,N_13625,N_12607);
or UO_1276 (O_1276,N_13115,N_14450);
and UO_1277 (O_1277,N_12797,N_12915);
nand UO_1278 (O_1278,N_13873,N_14688);
and UO_1279 (O_1279,N_14143,N_14108);
nor UO_1280 (O_1280,N_12577,N_13426);
xor UO_1281 (O_1281,N_13258,N_13759);
nand UO_1282 (O_1282,N_12806,N_14359);
and UO_1283 (O_1283,N_14221,N_13484);
or UO_1284 (O_1284,N_13551,N_14509);
nand UO_1285 (O_1285,N_13223,N_13652);
nand UO_1286 (O_1286,N_14106,N_13569);
and UO_1287 (O_1287,N_13746,N_12175);
xor UO_1288 (O_1288,N_12522,N_13513);
and UO_1289 (O_1289,N_13640,N_12042);
nand UO_1290 (O_1290,N_13877,N_12389);
or UO_1291 (O_1291,N_13894,N_12846);
and UO_1292 (O_1292,N_12339,N_14832);
and UO_1293 (O_1293,N_12687,N_13868);
or UO_1294 (O_1294,N_14974,N_14782);
nor UO_1295 (O_1295,N_13576,N_12618);
nand UO_1296 (O_1296,N_12377,N_12305);
nor UO_1297 (O_1297,N_13897,N_13863);
nand UO_1298 (O_1298,N_14577,N_13451);
or UO_1299 (O_1299,N_13848,N_14445);
and UO_1300 (O_1300,N_14436,N_13507);
nor UO_1301 (O_1301,N_12812,N_13083);
xnor UO_1302 (O_1302,N_12856,N_12460);
and UO_1303 (O_1303,N_12018,N_12077);
nand UO_1304 (O_1304,N_13237,N_14612);
and UO_1305 (O_1305,N_13967,N_13028);
xnor UO_1306 (O_1306,N_14966,N_12935);
and UO_1307 (O_1307,N_12654,N_12965);
nor UO_1308 (O_1308,N_12278,N_14951);
and UO_1309 (O_1309,N_13082,N_12700);
and UO_1310 (O_1310,N_14588,N_14522);
nand UO_1311 (O_1311,N_14729,N_13505);
nor UO_1312 (O_1312,N_13286,N_12933);
xnor UO_1313 (O_1313,N_14925,N_14856);
or UO_1314 (O_1314,N_14692,N_14178);
nor UO_1315 (O_1315,N_12163,N_14282);
and UO_1316 (O_1316,N_13635,N_13390);
nand UO_1317 (O_1317,N_13151,N_12603);
nand UO_1318 (O_1318,N_12811,N_14851);
or UO_1319 (O_1319,N_14215,N_13453);
nor UO_1320 (O_1320,N_13983,N_12451);
and UO_1321 (O_1321,N_12709,N_13628);
or UO_1322 (O_1322,N_12716,N_12983);
or UO_1323 (O_1323,N_14681,N_14080);
nor UO_1324 (O_1324,N_12353,N_13327);
and UO_1325 (O_1325,N_12916,N_12252);
nand UO_1326 (O_1326,N_13059,N_14662);
nand UO_1327 (O_1327,N_13504,N_14944);
and UO_1328 (O_1328,N_13614,N_12693);
nand UO_1329 (O_1329,N_13491,N_13300);
or UO_1330 (O_1330,N_13700,N_12463);
nand UO_1331 (O_1331,N_13466,N_14001);
nand UO_1332 (O_1332,N_14765,N_13527);
and UO_1333 (O_1333,N_14927,N_12083);
nor UO_1334 (O_1334,N_12871,N_12754);
nor UO_1335 (O_1335,N_12183,N_12374);
or UO_1336 (O_1336,N_13465,N_12106);
nor UO_1337 (O_1337,N_14939,N_12540);
or UO_1338 (O_1338,N_13381,N_14122);
and UO_1339 (O_1339,N_12594,N_14872);
nor UO_1340 (O_1340,N_14562,N_12670);
nor UO_1341 (O_1341,N_14324,N_12807);
nor UO_1342 (O_1342,N_14497,N_14399);
or UO_1343 (O_1343,N_14556,N_12244);
and UO_1344 (O_1344,N_12461,N_12138);
nand UO_1345 (O_1345,N_14013,N_14763);
or UO_1346 (O_1346,N_12159,N_14201);
nand UO_1347 (O_1347,N_13032,N_13208);
nand UO_1348 (O_1348,N_13474,N_12569);
xnor UO_1349 (O_1349,N_14975,N_12895);
nor UO_1350 (O_1350,N_14873,N_13812);
nand UO_1351 (O_1351,N_14627,N_14929);
or UO_1352 (O_1352,N_13100,N_13303);
nand UO_1353 (O_1353,N_13178,N_14069);
and UO_1354 (O_1354,N_12728,N_12437);
and UO_1355 (O_1355,N_14199,N_14717);
nand UO_1356 (O_1356,N_13496,N_13864);
nor UO_1357 (O_1357,N_14575,N_13809);
nand UO_1358 (O_1358,N_14775,N_14307);
xor UO_1359 (O_1359,N_14998,N_12465);
nand UO_1360 (O_1360,N_14369,N_14893);
and UO_1361 (O_1361,N_12739,N_12651);
nor UO_1362 (O_1362,N_14073,N_14414);
or UO_1363 (O_1363,N_14598,N_13875);
nand UO_1364 (O_1364,N_12835,N_12457);
nor UO_1365 (O_1365,N_14837,N_12740);
and UO_1366 (O_1366,N_13692,N_12852);
nand UO_1367 (O_1367,N_14843,N_12288);
and UO_1368 (O_1368,N_12283,N_12100);
nand UO_1369 (O_1369,N_12232,N_12710);
nor UO_1370 (O_1370,N_13038,N_13175);
xor UO_1371 (O_1371,N_13284,N_12078);
xnor UO_1372 (O_1372,N_13003,N_14759);
xor UO_1373 (O_1373,N_12623,N_12008);
xnor UO_1374 (O_1374,N_13460,N_12944);
nor UO_1375 (O_1375,N_14428,N_13939);
xnor UO_1376 (O_1376,N_14440,N_14291);
and UO_1377 (O_1377,N_12137,N_12367);
nor UO_1378 (O_1378,N_14750,N_12093);
and UO_1379 (O_1379,N_14735,N_14118);
nand UO_1380 (O_1380,N_13499,N_12030);
and UO_1381 (O_1381,N_13732,N_14935);
nor UO_1382 (O_1382,N_14861,N_13432);
nand UO_1383 (O_1383,N_13494,N_13396);
or UO_1384 (O_1384,N_12059,N_14349);
and UO_1385 (O_1385,N_13271,N_12637);
or UO_1386 (O_1386,N_12630,N_14885);
and UO_1387 (O_1387,N_14768,N_14070);
nand UO_1388 (O_1388,N_14719,N_14469);
or UO_1389 (O_1389,N_13057,N_14071);
and UO_1390 (O_1390,N_13123,N_12033);
or UO_1391 (O_1391,N_12659,N_12882);
nor UO_1392 (O_1392,N_14624,N_13525);
nor UO_1393 (O_1393,N_14028,N_14330);
nand UO_1394 (O_1394,N_12804,N_12949);
nand UO_1395 (O_1395,N_12822,N_14238);
and UO_1396 (O_1396,N_14715,N_12987);
xor UO_1397 (O_1397,N_14714,N_14648);
or UO_1398 (O_1398,N_13852,N_13981);
nand UO_1399 (O_1399,N_14432,N_12101);
nand UO_1400 (O_1400,N_12749,N_14858);
xnor UO_1401 (O_1401,N_12164,N_13568);
nand UO_1402 (O_1402,N_14329,N_12047);
or UO_1403 (O_1403,N_13690,N_12026);
nor UO_1404 (O_1404,N_13416,N_14082);
nand UO_1405 (O_1405,N_13382,N_13002);
and UO_1406 (O_1406,N_13523,N_12020);
nand UO_1407 (O_1407,N_14412,N_14152);
or UO_1408 (O_1408,N_13905,N_14388);
and UO_1409 (O_1409,N_13469,N_14113);
nand UO_1410 (O_1410,N_13559,N_13351);
nor UO_1411 (O_1411,N_12581,N_14248);
nand UO_1412 (O_1412,N_14270,N_13368);
nand UO_1413 (O_1413,N_13599,N_12418);
or UO_1414 (O_1414,N_12860,N_14461);
nor UO_1415 (O_1415,N_13947,N_13657);
and UO_1416 (O_1416,N_14230,N_14393);
or UO_1417 (O_1417,N_14132,N_12439);
nor UO_1418 (O_1418,N_13346,N_12325);
nor UO_1419 (O_1419,N_13122,N_14769);
nand UO_1420 (O_1420,N_13557,N_12664);
and UO_1421 (O_1421,N_12193,N_14931);
and UO_1422 (O_1422,N_12622,N_12041);
or UO_1423 (O_1423,N_14212,N_13823);
or UO_1424 (O_1424,N_14647,N_12246);
nand UO_1425 (O_1425,N_13748,N_13936);
nor UO_1426 (O_1426,N_12162,N_14200);
nor UO_1427 (O_1427,N_14628,N_14645);
nand UO_1428 (O_1428,N_13332,N_14833);
or UO_1429 (O_1429,N_14731,N_12861);
nand UO_1430 (O_1430,N_14442,N_14139);
nand UO_1431 (O_1431,N_13254,N_14306);
nand UO_1432 (O_1432,N_12177,N_13413);
nand UO_1433 (O_1433,N_14038,N_13970);
nor UO_1434 (O_1434,N_13921,N_14009);
and UO_1435 (O_1435,N_14984,N_13039);
or UO_1436 (O_1436,N_14781,N_12254);
nor UO_1437 (O_1437,N_13030,N_13558);
nand UO_1438 (O_1438,N_12862,N_12172);
and UO_1439 (O_1439,N_13162,N_14515);
nor UO_1440 (O_1440,N_13187,N_14056);
nand UO_1441 (O_1441,N_13220,N_14682);
nor UO_1442 (O_1442,N_14732,N_14563);
and UO_1443 (O_1443,N_14062,N_14909);
and UO_1444 (O_1444,N_14276,N_12612);
nand UO_1445 (O_1445,N_12793,N_12285);
nor UO_1446 (O_1446,N_12206,N_13903);
nor UO_1447 (O_1447,N_12979,N_13435);
nor UO_1448 (O_1448,N_12605,N_14231);
nand UO_1449 (O_1449,N_13412,N_12329);
and UO_1450 (O_1450,N_12277,N_13688);
nand UO_1451 (O_1451,N_12832,N_13790);
or UO_1452 (O_1452,N_14413,N_14504);
nand UO_1453 (O_1453,N_14033,N_13063);
xnor UO_1454 (O_1454,N_13604,N_12432);
nand UO_1455 (O_1455,N_12167,N_13712);
or UO_1456 (O_1456,N_12772,N_13392);
and UO_1457 (O_1457,N_12584,N_13266);
nand UO_1458 (O_1458,N_14367,N_14097);
xor UO_1459 (O_1459,N_13636,N_13889);
and UO_1460 (O_1460,N_13052,N_13034);
and UO_1461 (O_1461,N_12724,N_12468);
nand UO_1462 (O_1462,N_14115,N_12227);
nor UO_1463 (O_1463,N_13989,N_14983);
nand UO_1464 (O_1464,N_13564,N_13893);
nor UO_1465 (O_1465,N_12619,N_12599);
nand UO_1466 (O_1466,N_13439,N_14548);
xor UO_1467 (O_1467,N_14439,N_14581);
nand UO_1468 (O_1468,N_13818,N_14426);
and UO_1469 (O_1469,N_13951,N_13365);
or UO_1470 (O_1470,N_13858,N_13307);
nand UO_1471 (O_1471,N_13035,N_12863);
nand UO_1472 (O_1472,N_14767,N_13226);
nand UO_1473 (O_1473,N_14353,N_12780);
nor UO_1474 (O_1474,N_14783,N_14205);
or UO_1475 (O_1475,N_12263,N_12827);
nand UO_1476 (O_1476,N_12240,N_12469);
and UO_1477 (O_1477,N_13980,N_13467);
or UO_1478 (O_1478,N_14299,N_13744);
nor UO_1479 (O_1479,N_14197,N_13917);
xor UO_1480 (O_1480,N_14713,N_13077);
and UO_1481 (O_1481,N_13027,N_13116);
and UO_1482 (O_1482,N_14618,N_12562);
nor UO_1483 (O_1483,N_14830,N_13843);
or UO_1484 (O_1484,N_14415,N_14916);
and UO_1485 (O_1485,N_13278,N_12537);
nand UO_1486 (O_1486,N_14700,N_12508);
or UO_1487 (O_1487,N_13373,N_13785);
nor UO_1488 (O_1488,N_12816,N_14572);
nor UO_1489 (O_1489,N_13998,N_12481);
nand UO_1490 (O_1490,N_14820,N_13737);
xnor UO_1491 (O_1491,N_13580,N_14059);
xnor UO_1492 (O_1492,N_14465,N_13305);
and UO_1493 (O_1493,N_13931,N_14602);
nor UO_1494 (O_1494,N_12689,N_14020);
and UO_1495 (O_1495,N_14424,N_13184);
nand UO_1496 (O_1496,N_12161,N_12478);
nand UO_1497 (O_1497,N_13075,N_13292);
nor UO_1498 (O_1498,N_12506,N_13176);
nor UO_1499 (O_1499,N_13701,N_14124);
nor UO_1500 (O_1500,N_14055,N_14660);
nand UO_1501 (O_1501,N_12511,N_12825);
xnor UO_1502 (O_1502,N_13737,N_14134);
or UO_1503 (O_1503,N_12252,N_13987);
nand UO_1504 (O_1504,N_12548,N_14026);
or UO_1505 (O_1505,N_14498,N_12499);
and UO_1506 (O_1506,N_14695,N_13861);
nor UO_1507 (O_1507,N_13168,N_14949);
nand UO_1508 (O_1508,N_12103,N_13712);
or UO_1509 (O_1509,N_13905,N_14493);
nand UO_1510 (O_1510,N_13055,N_13496);
or UO_1511 (O_1511,N_12762,N_12967);
or UO_1512 (O_1512,N_13743,N_12483);
or UO_1513 (O_1513,N_14690,N_12357);
nor UO_1514 (O_1514,N_14247,N_13906);
or UO_1515 (O_1515,N_14113,N_12221);
nor UO_1516 (O_1516,N_13170,N_14416);
nand UO_1517 (O_1517,N_13939,N_12690);
and UO_1518 (O_1518,N_14514,N_12470);
nor UO_1519 (O_1519,N_14750,N_13445);
or UO_1520 (O_1520,N_13749,N_12233);
xnor UO_1521 (O_1521,N_13717,N_12843);
and UO_1522 (O_1522,N_12039,N_13229);
nor UO_1523 (O_1523,N_14281,N_14562);
nand UO_1524 (O_1524,N_12063,N_13469);
and UO_1525 (O_1525,N_12130,N_13342);
nor UO_1526 (O_1526,N_13334,N_12153);
nor UO_1527 (O_1527,N_12789,N_14121);
nor UO_1528 (O_1528,N_13221,N_14873);
nand UO_1529 (O_1529,N_14170,N_14527);
and UO_1530 (O_1530,N_14412,N_13257);
nand UO_1531 (O_1531,N_13282,N_13280);
nand UO_1532 (O_1532,N_12378,N_12428);
or UO_1533 (O_1533,N_14567,N_13501);
nor UO_1534 (O_1534,N_12637,N_12746);
nor UO_1535 (O_1535,N_12348,N_14495);
nor UO_1536 (O_1536,N_13441,N_14116);
and UO_1537 (O_1537,N_14231,N_12701);
nor UO_1538 (O_1538,N_14414,N_13714);
xor UO_1539 (O_1539,N_14559,N_12810);
nor UO_1540 (O_1540,N_13033,N_12276);
nand UO_1541 (O_1541,N_12567,N_12712);
or UO_1542 (O_1542,N_12180,N_13223);
or UO_1543 (O_1543,N_12156,N_14933);
or UO_1544 (O_1544,N_13131,N_13948);
nand UO_1545 (O_1545,N_14742,N_14260);
and UO_1546 (O_1546,N_14270,N_13265);
and UO_1547 (O_1547,N_13457,N_14983);
nor UO_1548 (O_1548,N_12897,N_14234);
nor UO_1549 (O_1549,N_14634,N_14148);
or UO_1550 (O_1550,N_14815,N_12147);
and UO_1551 (O_1551,N_12423,N_13524);
xnor UO_1552 (O_1552,N_14363,N_14639);
nor UO_1553 (O_1553,N_12317,N_12567);
nor UO_1554 (O_1554,N_13908,N_12268);
and UO_1555 (O_1555,N_14863,N_14313);
or UO_1556 (O_1556,N_12758,N_14044);
or UO_1557 (O_1557,N_14809,N_13119);
or UO_1558 (O_1558,N_13692,N_13953);
nand UO_1559 (O_1559,N_12201,N_12698);
nand UO_1560 (O_1560,N_12891,N_12397);
xor UO_1561 (O_1561,N_13384,N_14062);
nor UO_1562 (O_1562,N_13629,N_14807);
nor UO_1563 (O_1563,N_12020,N_13220);
or UO_1564 (O_1564,N_12579,N_12686);
nand UO_1565 (O_1565,N_12566,N_13005);
and UO_1566 (O_1566,N_13940,N_12153);
or UO_1567 (O_1567,N_12445,N_13180);
or UO_1568 (O_1568,N_14347,N_12744);
and UO_1569 (O_1569,N_12001,N_13590);
or UO_1570 (O_1570,N_13436,N_14422);
nand UO_1571 (O_1571,N_13950,N_13086);
xor UO_1572 (O_1572,N_12911,N_14015);
or UO_1573 (O_1573,N_13271,N_13470);
nor UO_1574 (O_1574,N_14542,N_14379);
and UO_1575 (O_1575,N_12574,N_14797);
nor UO_1576 (O_1576,N_13916,N_13914);
or UO_1577 (O_1577,N_14624,N_12983);
and UO_1578 (O_1578,N_12817,N_13585);
nand UO_1579 (O_1579,N_12559,N_13122);
xor UO_1580 (O_1580,N_14139,N_14285);
or UO_1581 (O_1581,N_12732,N_12943);
nor UO_1582 (O_1582,N_12520,N_12936);
and UO_1583 (O_1583,N_14257,N_13896);
nor UO_1584 (O_1584,N_13153,N_13117);
and UO_1585 (O_1585,N_12888,N_14499);
or UO_1586 (O_1586,N_12995,N_14894);
and UO_1587 (O_1587,N_13432,N_13815);
nand UO_1588 (O_1588,N_14210,N_13331);
nand UO_1589 (O_1589,N_12226,N_13998);
or UO_1590 (O_1590,N_13682,N_14992);
or UO_1591 (O_1591,N_13476,N_12203);
and UO_1592 (O_1592,N_12790,N_13672);
xor UO_1593 (O_1593,N_12255,N_13721);
and UO_1594 (O_1594,N_13245,N_13660);
nand UO_1595 (O_1595,N_12222,N_13605);
and UO_1596 (O_1596,N_14635,N_14504);
xnor UO_1597 (O_1597,N_12669,N_13273);
and UO_1598 (O_1598,N_14332,N_12458);
or UO_1599 (O_1599,N_13899,N_12691);
or UO_1600 (O_1600,N_12326,N_12280);
or UO_1601 (O_1601,N_14811,N_14946);
or UO_1602 (O_1602,N_14160,N_14275);
and UO_1603 (O_1603,N_12278,N_13102);
or UO_1604 (O_1604,N_14425,N_13506);
and UO_1605 (O_1605,N_13483,N_14075);
and UO_1606 (O_1606,N_14788,N_12792);
nand UO_1607 (O_1607,N_12765,N_12342);
nor UO_1608 (O_1608,N_12164,N_13133);
nand UO_1609 (O_1609,N_13190,N_12476);
nor UO_1610 (O_1610,N_14095,N_13761);
nor UO_1611 (O_1611,N_13682,N_12705);
nand UO_1612 (O_1612,N_12365,N_13811);
nor UO_1613 (O_1613,N_12140,N_13633);
or UO_1614 (O_1614,N_14146,N_13769);
or UO_1615 (O_1615,N_12833,N_14107);
nor UO_1616 (O_1616,N_14053,N_12851);
nor UO_1617 (O_1617,N_13572,N_13192);
nand UO_1618 (O_1618,N_14835,N_14943);
or UO_1619 (O_1619,N_12528,N_12162);
and UO_1620 (O_1620,N_12776,N_14918);
or UO_1621 (O_1621,N_12362,N_14697);
and UO_1622 (O_1622,N_12917,N_14499);
or UO_1623 (O_1623,N_12541,N_13935);
nand UO_1624 (O_1624,N_13320,N_12706);
and UO_1625 (O_1625,N_14414,N_14103);
nand UO_1626 (O_1626,N_12944,N_14836);
nor UO_1627 (O_1627,N_14871,N_13490);
and UO_1628 (O_1628,N_14159,N_13978);
nor UO_1629 (O_1629,N_14371,N_12078);
nor UO_1630 (O_1630,N_13148,N_13039);
or UO_1631 (O_1631,N_13608,N_12449);
nor UO_1632 (O_1632,N_14382,N_14585);
or UO_1633 (O_1633,N_14180,N_14596);
nand UO_1634 (O_1634,N_13775,N_13234);
or UO_1635 (O_1635,N_12124,N_14164);
nor UO_1636 (O_1636,N_14238,N_12779);
nor UO_1637 (O_1637,N_13434,N_13071);
and UO_1638 (O_1638,N_13523,N_13476);
xnor UO_1639 (O_1639,N_14039,N_14229);
xor UO_1640 (O_1640,N_14879,N_12185);
nand UO_1641 (O_1641,N_14467,N_13371);
nand UO_1642 (O_1642,N_13393,N_12916);
or UO_1643 (O_1643,N_12317,N_13565);
or UO_1644 (O_1644,N_13392,N_12196);
and UO_1645 (O_1645,N_12495,N_13395);
and UO_1646 (O_1646,N_13772,N_12289);
nand UO_1647 (O_1647,N_13171,N_14585);
nand UO_1648 (O_1648,N_12934,N_12366);
or UO_1649 (O_1649,N_14648,N_14764);
and UO_1650 (O_1650,N_12843,N_12051);
and UO_1651 (O_1651,N_13484,N_14251);
nand UO_1652 (O_1652,N_13404,N_12426);
nor UO_1653 (O_1653,N_13036,N_14641);
nand UO_1654 (O_1654,N_12690,N_13209);
and UO_1655 (O_1655,N_14846,N_12362);
or UO_1656 (O_1656,N_13258,N_12217);
xor UO_1657 (O_1657,N_14215,N_14737);
nand UO_1658 (O_1658,N_12791,N_14356);
nor UO_1659 (O_1659,N_13426,N_14550);
nor UO_1660 (O_1660,N_12183,N_14563);
and UO_1661 (O_1661,N_12439,N_12912);
and UO_1662 (O_1662,N_14131,N_12689);
nor UO_1663 (O_1663,N_14735,N_13952);
or UO_1664 (O_1664,N_14991,N_12100);
and UO_1665 (O_1665,N_14201,N_12124);
nand UO_1666 (O_1666,N_13195,N_13584);
or UO_1667 (O_1667,N_13624,N_14540);
or UO_1668 (O_1668,N_12630,N_13248);
and UO_1669 (O_1669,N_14839,N_14358);
xor UO_1670 (O_1670,N_12774,N_14311);
or UO_1671 (O_1671,N_13773,N_13838);
nand UO_1672 (O_1672,N_13320,N_12306);
xnor UO_1673 (O_1673,N_13381,N_13653);
and UO_1674 (O_1674,N_14955,N_13915);
xnor UO_1675 (O_1675,N_13183,N_13607);
nor UO_1676 (O_1676,N_12236,N_14486);
nor UO_1677 (O_1677,N_14637,N_14333);
and UO_1678 (O_1678,N_12329,N_13596);
nor UO_1679 (O_1679,N_12087,N_14103);
nor UO_1680 (O_1680,N_13923,N_14163);
or UO_1681 (O_1681,N_13202,N_14066);
or UO_1682 (O_1682,N_14011,N_13030);
nor UO_1683 (O_1683,N_12794,N_13623);
xor UO_1684 (O_1684,N_14060,N_14204);
xnor UO_1685 (O_1685,N_14637,N_13855);
or UO_1686 (O_1686,N_14689,N_12795);
or UO_1687 (O_1687,N_12509,N_13606);
and UO_1688 (O_1688,N_12288,N_14877);
nor UO_1689 (O_1689,N_13622,N_13821);
nor UO_1690 (O_1690,N_12850,N_13048);
and UO_1691 (O_1691,N_14121,N_12454);
or UO_1692 (O_1692,N_12762,N_14830);
xor UO_1693 (O_1693,N_14203,N_13090);
xor UO_1694 (O_1694,N_13724,N_12262);
nor UO_1695 (O_1695,N_14057,N_13510);
or UO_1696 (O_1696,N_14077,N_12519);
or UO_1697 (O_1697,N_12338,N_13805);
and UO_1698 (O_1698,N_12695,N_12665);
or UO_1699 (O_1699,N_13363,N_12795);
nor UO_1700 (O_1700,N_13142,N_12273);
nand UO_1701 (O_1701,N_14800,N_13654);
xor UO_1702 (O_1702,N_12759,N_12565);
nand UO_1703 (O_1703,N_14232,N_13844);
nor UO_1704 (O_1704,N_12337,N_13037);
and UO_1705 (O_1705,N_12151,N_12636);
or UO_1706 (O_1706,N_12678,N_12169);
and UO_1707 (O_1707,N_14078,N_14257);
and UO_1708 (O_1708,N_13797,N_14826);
and UO_1709 (O_1709,N_13024,N_13605);
nor UO_1710 (O_1710,N_13030,N_13541);
or UO_1711 (O_1711,N_12261,N_13768);
or UO_1712 (O_1712,N_13137,N_12131);
or UO_1713 (O_1713,N_12044,N_14403);
nand UO_1714 (O_1714,N_12441,N_13497);
nand UO_1715 (O_1715,N_12624,N_13931);
nor UO_1716 (O_1716,N_14633,N_12836);
and UO_1717 (O_1717,N_13898,N_13389);
and UO_1718 (O_1718,N_14875,N_14261);
nor UO_1719 (O_1719,N_12698,N_12593);
nor UO_1720 (O_1720,N_14439,N_13253);
or UO_1721 (O_1721,N_14678,N_13722);
nand UO_1722 (O_1722,N_14394,N_13682);
or UO_1723 (O_1723,N_12058,N_13364);
nand UO_1724 (O_1724,N_13289,N_13255);
or UO_1725 (O_1725,N_13778,N_13395);
and UO_1726 (O_1726,N_14382,N_14512);
or UO_1727 (O_1727,N_13405,N_12976);
xor UO_1728 (O_1728,N_14542,N_13187);
or UO_1729 (O_1729,N_12969,N_13127);
and UO_1730 (O_1730,N_14635,N_13364);
nand UO_1731 (O_1731,N_13456,N_12792);
nand UO_1732 (O_1732,N_13199,N_13239);
xnor UO_1733 (O_1733,N_13441,N_12156);
or UO_1734 (O_1734,N_13418,N_13432);
or UO_1735 (O_1735,N_14029,N_12539);
nand UO_1736 (O_1736,N_13771,N_13582);
or UO_1737 (O_1737,N_14891,N_14802);
nand UO_1738 (O_1738,N_13533,N_14614);
nand UO_1739 (O_1739,N_12036,N_12208);
nor UO_1740 (O_1740,N_12598,N_12018);
or UO_1741 (O_1741,N_14973,N_14210);
nor UO_1742 (O_1742,N_13189,N_12855);
nor UO_1743 (O_1743,N_13150,N_14803);
nor UO_1744 (O_1744,N_12442,N_12249);
nand UO_1745 (O_1745,N_12761,N_13875);
and UO_1746 (O_1746,N_13577,N_14037);
or UO_1747 (O_1747,N_14749,N_13135);
nor UO_1748 (O_1748,N_12344,N_12766);
and UO_1749 (O_1749,N_12136,N_14703);
or UO_1750 (O_1750,N_14393,N_14263);
nor UO_1751 (O_1751,N_14248,N_12695);
or UO_1752 (O_1752,N_12610,N_13606);
and UO_1753 (O_1753,N_12748,N_12944);
and UO_1754 (O_1754,N_13231,N_14297);
nand UO_1755 (O_1755,N_13373,N_13824);
xor UO_1756 (O_1756,N_14418,N_14883);
and UO_1757 (O_1757,N_13411,N_14605);
nand UO_1758 (O_1758,N_13624,N_12057);
or UO_1759 (O_1759,N_14085,N_13995);
or UO_1760 (O_1760,N_14265,N_12624);
xor UO_1761 (O_1761,N_12145,N_12619);
or UO_1762 (O_1762,N_12234,N_14139);
nor UO_1763 (O_1763,N_14591,N_12871);
nand UO_1764 (O_1764,N_13068,N_13103);
and UO_1765 (O_1765,N_13296,N_13739);
and UO_1766 (O_1766,N_12781,N_14528);
nor UO_1767 (O_1767,N_14687,N_13339);
nor UO_1768 (O_1768,N_14565,N_12751);
nand UO_1769 (O_1769,N_13724,N_12363);
or UO_1770 (O_1770,N_14769,N_12805);
xnor UO_1771 (O_1771,N_14592,N_12942);
nand UO_1772 (O_1772,N_12530,N_13430);
and UO_1773 (O_1773,N_13599,N_13846);
and UO_1774 (O_1774,N_13951,N_14492);
xor UO_1775 (O_1775,N_14819,N_14503);
and UO_1776 (O_1776,N_14892,N_14475);
nand UO_1777 (O_1777,N_14059,N_14624);
nor UO_1778 (O_1778,N_12007,N_12479);
nor UO_1779 (O_1779,N_13689,N_12676);
and UO_1780 (O_1780,N_12875,N_14897);
nor UO_1781 (O_1781,N_12881,N_14685);
and UO_1782 (O_1782,N_12808,N_12468);
or UO_1783 (O_1783,N_13498,N_12721);
nor UO_1784 (O_1784,N_12281,N_13929);
nor UO_1785 (O_1785,N_12175,N_14017);
and UO_1786 (O_1786,N_14617,N_12871);
nand UO_1787 (O_1787,N_13717,N_13695);
and UO_1788 (O_1788,N_14746,N_13793);
nor UO_1789 (O_1789,N_13341,N_12763);
and UO_1790 (O_1790,N_13547,N_13332);
xnor UO_1791 (O_1791,N_13151,N_14739);
or UO_1792 (O_1792,N_12381,N_12969);
or UO_1793 (O_1793,N_13043,N_12447);
xor UO_1794 (O_1794,N_13304,N_12970);
nand UO_1795 (O_1795,N_13589,N_12890);
nor UO_1796 (O_1796,N_12122,N_13804);
and UO_1797 (O_1797,N_12336,N_14252);
and UO_1798 (O_1798,N_12359,N_12772);
and UO_1799 (O_1799,N_13773,N_13644);
and UO_1800 (O_1800,N_13392,N_13784);
nand UO_1801 (O_1801,N_12634,N_12423);
nand UO_1802 (O_1802,N_13389,N_14914);
or UO_1803 (O_1803,N_14385,N_13736);
nor UO_1804 (O_1804,N_14639,N_13494);
nor UO_1805 (O_1805,N_12113,N_12650);
or UO_1806 (O_1806,N_12601,N_13288);
nand UO_1807 (O_1807,N_12010,N_14103);
nand UO_1808 (O_1808,N_13134,N_13513);
and UO_1809 (O_1809,N_13705,N_13262);
or UO_1810 (O_1810,N_12148,N_13790);
or UO_1811 (O_1811,N_14713,N_14926);
and UO_1812 (O_1812,N_12153,N_13861);
xnor UO_1813 (O_1813,N_13510,N_13672);
nor UO_1814 (O_1814,N_12099,N_14119);
and UO_1815 (O_1815,N_13548,N_14750);
nor UO_1816 (O_1816,N_14177,N_13393);
or UO_1817 (O_1817,N_14317,N_12095);
xnor UO_1818 (O_1818,N_12835,N_13987);
nor UO_1819 (O_1819,N_13173,N_13563);
nand UO_1820 (O_1820,N_14244,N_12207);
and UO_1821 (O_1821,N_14804,N_12055);
nor UO_1822 (O_1822,N_14266,N_14312);
or UO_1823 (O_1823,N_14687,N_12321);
nand UO_1824 (O_1824,N_13865,N_14264);
nand UO_1825 (O_1825,N_13318,N_13470);
and UO_1826 (O_1826,N_13001,N_12852);
and UO_1827 (O_1827,N_14356,N_12461);
or UO_1828 (O_1828,N_14715,N_14258);
nand UO_1829 (O_1829,N_12076,N_13570);
or UO_1830 (O_1830,N_14393,N_14016);
nand UO_1831 (O_1831,N_12328,N_14316);
nand UO_1832 (O_1832,N_14327,N_12645);
or UO_1833 (O_1833,N_13843,N_12955);
or UO_1834 (O_1834,N_14936,N_13864);
xnor UO_1835 (O_1835,N_13388,N_14470);
or UO_1836 (O_1836,N_14215,N_14528);
or UO_1837 (O_1837,N_13244,N_14071);
and UO_1838 (O_1838,N_14270,N_13171);
nand UO_1839 (O_1839,N_14866,N_12274);
or UO_1840 (O_1840,N_14745,N_13513);
nand UO_1841 (O_1841,N_14353,N_14923);
xnor UO_1842 (O_1842,N_14440,N_12970);
nor UO_1843 (O_1843,N_14757,N_12437);
and UO_1844 (O_1844,N_14156,N_12167);
nand UO_1845 (O_1845,N_14486,N_14178);
nor UO_1846 (O_1846,N_13676,N_13297);
nor UO_1847 (O_1847,N_14570,N_13087);
and UO_1848 (O_1848,N_12985,N_14382);
or UO_1849 (O_1849,N_12195,N_12518);
nand UO_1850 (O_1850,N_14582,N_14980);
nor UO_1851 (O_1851,N_12763,N_14012);
and UO_1852 (O_1852,N_13591,N_14581);
xnor UO_1853 (O_1853,N_12327,N_12983);
xor UO_1854 (O_1854,N_14240,N_13954);
nand UO_1855 (O_1855,N_13230,N_14479);
and UO_1856 (O_1856,N_14339,N_14523);
nand UO_1857 (O_1857,N_14367,N_13858);
nand UO_1858 (O_1858,N_13661,N_12251);
or UO_1859 (O_1859,N_12278,N_14237);
and UO_1860 (O_1860,N_14867,N_12681);
nand UO_1861 (O_1861,N_13841,N_14574);
or UO_1862 (O_1862,N_12338,N_13935);
or UO_1863 (O_1863,N_14661,N_14653);
or UO_1864 (O_1864,N_14071,N_12394);
or UO_1865 (O_1865,N_14742,N_13763);
or UO_1866 (O_1866,N_13112,N_13630);
or UO_1867 (O_1867,N_14550,N_12838);
xnor UO_1868 (O_1868,N_12476,N_12318);
nand UO_1869 (O_1869,N_12325,N_13740);
and UO_1870 (O_1870,N_12908,N_14345);
nor UO_1871 (O_1871,N_14664,N_14345);
nor UO_1872 (O_1872,N_12309,N_14428);
nand UO_1873 (O_1873,N_14982,N_12363);
nor UO_1874 (O_1874,N_12040,N_14949);
nor UO_1875 (O_1875,N_14911,N_12991);
nor UO_1876 (O_1876,N_12629,N_12871);
nor UO_1877 (O_1877,N_12807,N_14127);
xor UO_1878 (O_1878,N_12982,N_14586);
nor UO_1879 (O_1879,N_13871,N_12672);
and UO_1880 (O_1880,N_13494,N_13794);
nand UO_1881 (O_1881,N_14528,N_14492);
nand UO_1882 (O_1882,N_12406,N_12683);
nand UO_1883 (O_1883,N_14823,N_14290);
nor UO_1884 (O_1884,N_14402,N_13218);
or UO_1885 (O_1885,N_14052,N_12220);
or UO_1886 (O_1886,N_12190,N_14839);
nand UO_1887 (O_1887,N_13314,N_14762);
or UO_1888 (O_1888,N_12393,N_13701);
nand UO_1889 (O_1889,N_13252,N_12291);
nor UO_1890 (O_1890,N_12839,N_14363);
and UO_1891 (O_1891,N_13851,N_14763);
and UO_1892 (O_1892,N_14428,N_13220);
and UO_1893 (O_1893,N_12269,N_13976);
xor UO_1894 (O_1894,N_13440,N_12727);
nor UO_1895 (O_1895,N_12436,N_13595);
nand UO_1896 (O_1896,N_13418,N_12720);
nor UO_1897 (O_1897,N_14596,N_12456);
nor UO_1898 (O_1898,N_14844,N_12738);
nor UO_1899 (O_1899,N_13429,N_13931);
or UO_1900 (O_1900,N_14132,N_13032);
nor UO_1901 (O_1901,N_12428,N_13152);
or UO_1902 (O_1902,N_13487,N_12923);
nor UO_1903 (O_1903,N_13647,N_12755);
nand UO_1904 (O_1904,N_12945,N_13647);
nand UO_1905 (O_1905,N_12932,N_14941);
nand UO_1906 (O_1906,N_13995,N_12399);
and UO_1907 (O_1907,N_12624,N_12128);
nand UO_1908 (O_1908,N_12819,N_12543);
xnor UO_1909 (O_1909,N_14482,N_14109);
or UO_1910 (O_1910,N_14122,N_14052);
and UO_1911 (O_1911,N_13936,N_12884);
xnor UO_1912 (O_1912,N_13193,N_14953);
and UO_1913 (O_1913,N_12851,N_13395);
or UO_1914 (O_1914,N_12696,N_13402);
or UO_1915 (O_1915,N_14705,N_13129);
and UO_1916 (O_1916,N_13882,N_13714);
xnor UO_1917 (O_1917,N_14013,N_12327);
nor UO_1918 (O_1918,N_12452,N_13875);
nand UO_1919 (O_1919,N_12268,N_14722);
or UO_1920 (O_1920,N_14149,N_14446);
nand UO_1921 (O_1921,N_14202,N_14147);
nor UO_1922 (O_1922,N_13954,N_12041);
nor UO_1923 (O_1923,N_14546,N_13311);
nor UO_1924 (O_1924,N_12351,N_14708);
nand UO_1925 (O_1925,N_12065,N_14017);
nand UO_1926 (O_1926,N_14938,N_14152);
and UO_1927 (O_1927,N_12791,N_14992);
nand UO_1928 (O_1928,N_12190,N_14055);
or UO_1929 (O_1929,N_12297,N_12340);
nand UO_1930 (O_1930,N_13344,N_14971);
nand UO_1931 (O_1931,N_13830,N_13792);
nand UO_1932 (O_1932,N_13367,N_14939);
nand UO_1933 (O_1933,N_13938,N_12628);
or UO_1934 (O_1934,N_14205,N_13429);
nand UO_1935 (O_1935,N_13099,N_12874);
xor UO_1936 (O_1936,N_12507,N_13434);
or UO_1937 (O_1937,N_12029,N_13351);
and UO_1938 (O_1938,N_14192,N_13744);
xnor UO_1939 (O_1939,N_14680,N_14041);
nand UO_1940 (O_1940,N_14157,N_12218);
or UO_1941 (O_1941,N_14864,N_12961);
nor UO_1942 (O_1942,N_14311,N_14598);
or UO_1943 (O_1943,N_14622,N_13362);
nand UO_1944 (O_1944,N_14602,N_13414);
or UO_1945 (O_1945,N_14071,N_14488);
xnor UO_1946 (O_1946,N_14566,N_12727);
and UO_1947 (O_1947,N_13776,N_14941);
nand UO_1948 (O_1948,N_12403,N_13560);
and UO_1949 (O_1949,N_12402,N_13645);
or UO_1950 (O_1950,N_14342,N_12357);
or UO_1951 (O_1951,N_13594,N_14712);
or UO_1952 (O_1952,N_13437,N_13172);
nor UO_1953 (O_1953,N_13456,N_12467);
or UO_1954 (O_1954,N_13820,N_13547);
and UO_1955 (O_1955,N_14666,N_12904);
nand UO_1956 (O_1956,N_12962,N_13757);
nor UO_1957 (O_1957,N_12026,N_14020);
nand UO_1958 (O_1958,N_13482,N_12158);
nand UO_1959 (O_1959,N_12928,N_13154);
nand UO_1960 (O_1960,N_12359,N_14534);
or UO_1961 (O_1961,N_13612,N_14643);
and UO_1962 (O_1962,N_12613,N_13372);
nor UO_1963 (O_1963,N_12457,N_14954);
nand UO_1964 (O_1964,N_13270,N_14829);
or UO_1965 (O_1965,N_12844,N_13346);
or UO_1966 (O_1966,N_13587,N_14713);
xor UO_1967 (O_1967,N_14966,N_14781);
nand UO_1968 (O_1968,N_13615,N_13534);
or UO_1969 (O_1969,N_12339,N_14554);
and UO_1970 (O_1970,N_14191,N_14114);
xor UO_1971 (O_1971,N_14183,N_13398);
or UO_1972 (O_1972,N_12802,N_13349);
nor UO_1973 (O_1973,N_13718,N_12264);
and UO_1974 (O_1974,N_14988,N_14173);
xnor UO_1975 (O_1975,N_13468,N_12309);
nand UO_1976 (O_1976,N_12282,N_12175);
or UO_1977 (O_1977,N_14407,N_13934);
nor UO_1978 (O_1978,N_14294,N_14144);
and UO_1979 (O_1979,N_14166,N_12103);
nand UO_1980 (O_1980,N_12634,N_13532);
and UO_1981 (O_1981,N_14398,N_12581);
nor UO_1982 (O_1982,N_13501,N_14618);
nand UO_1983 (O_1983,N_14956,N_12184);
nor UO_1984 (O_1984,N_14763,N_12975);
and UO_1985 (O_1985,N_13213,N_12347);
nor UO_1986 (O_1986,N_13152,N_14783);
nand UO_1987 (O_1987,N_13366,N_12611);
and UO_1988 (O_1988,N_12120,N_12385);
or UO_1989 (O_1989,N_12741,N_13250);
or UO_1990 (O_1990,N_14488,N_14337);
nor UO_1991 (O_1991,N_13612,N_12500);
nand UO_1992 (O_1992,N_14011,N_14045);
nand UO_1993 (O_1993,N_14004,N_14244);
or UO_1994 (O_1994,N_12229,N_13720);
xor UO_1995 (O_1995,N_12190,N_12991);
or UO_1996 (O_1996,N_14963,N_12539);
and UO_1997 (O_1997,N_13684,N_12484);
nor UO_1998 (O_1998,N_13263,N_13926);
nand UO_1999 (O_1999,N_13225,N_13549);
endmodule