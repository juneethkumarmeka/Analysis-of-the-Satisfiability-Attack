module basic_1000_10000_1500_20_levels_10xor_7(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999;
nor U0 (N_0,In_387,In_118);
nand U1 (N_1,In_677,In_306);
and U2 (N_2,In_325,In_432);
or U3 (N_3,In_887,In_304);
xnor U4 (N_4,In_319,In_159);
nor U5 (N_5,In_23,In_795);
or U6 (N_6,In_721,In_616);
and U7 (N_7,In_285,In_389);
nor U8 (N_8,In_402,In_386);
or U9 (N_9,In_859,In_660);
nor U10 (N_10,In_261,In_152);
nor U11 (N_11,In_61,In_326);
nand U12 (N_12,In_580,In_236);
nor U13 (N_13,In_6,In_674);
and U14 (N_14,In_364,In_665);
xnor U15 (N_15,In_802,In_273);
nand U16 (N_16,In_33,In_164);
nand U17 (N_17,In_936,In_866);
nand U18 (N_18,In_209,In_301);
and U19 (N_19,In_498,In_652);
xor U20 (N_20,In_403,In_920);
or U21 (N_21,In_262,In_300);
nand U22 (N_22,In_67,In_756);
xor U23 (N_23,In_27,In_14);
nand U24 (N_24,In_452,In_267);
and U25 (N_25,In_295,In_987);
nor U26 (N_26,In_438,In_450);
nand U27 (N_27,In_58,In_957);
nand U28 (N_28,In_686,In_345);
and U29 (N_29,In_829,In_318);
xnor U30 (N_30,In_979,In_373);
nand U31 (N_31,In_34,In_971);
nand U32 (N_32,In_896,In_603);
xnor U33 (N_33,In_716,In_828);
or U34 (N_34,In_395,In_631);
xnor U35 (N_35,In_800,In_535);
xnor U36 (N_36,In_976,In_230);
and U37 (N_37,In_843,In_197);
nand U38 (N_38,In_410,In_915);
nand U39 (N_39,In_64,In_258);
and U40 (N_40,In_767,In_298);
and U41 (N_41,In_992,In_259);
or U42 (N_42,In_11,In_500);
xnor U43 (N_43,In_534,In_529);
or U44 (N_44,In_695,In_292);
nor U45 (N_45,In_321,In_142);
and U46 (N_46,In_1,In_646);
and U47 (N_47,In_173,In_494);
xor U48 (N_48,In_248,In_71);
and U49 (N_49,In_693,In_350);
nand U50 (N_50,In_485,In_542);
or U51 (N_51,In_384,In_45);
and U52 (N_52,In_80,In_909);
xnor U53 (N_53,In_531,In_539);
nand U54 (N_54,In_931,In_997);
or U55 (N_55,In_825,In_816);
or U56 (N_56,In_963,In_483);
nor U57 (N_57,In_264,In_73);
xor U58 (N_58,In_35,In_769);
nor U59 (N_59,In_691,In_25);
and U60 (N_60,In_464,In_840);
xor U61 (N_61,In_311,In_481);
nor U62 (N_62,In_833,In_585);
nor U63 (N_63,In_359,In_251);
and U64 (N_64,In_933,In_240);
nor U65 (N_65,In_889,In_290);
and U66 (N_66,In_553,In_85);
and U67 (N_67,In_948,In_794);
or U68 (N_68,In_676,In_569);
nand U69 (N_69,In_469,In_703);
and U70 (N_70,In_516,In_145);
nand U71 (N_71,In_898,In_893);
xnor U72 (N_72,In_678,In_351);
or U73 (N_73,In_120,In_89);
nand U74 (N_74,In_999,In_761);
nand U75 (N_75,In_133,In_658);
and U76 (N_76,In_48,In_86);
xor U77 (N_77,In_265,In_177);
nor U78 (N_78,In_137,In_227);
nor U79 (N_79,In_499,In_930);
and U80 (N_80,In_755,In_174);
xnor U81 (N_81,In_30,In_907);
or U82 (N_82,In_683,In_482);
nand U83 (N_83,In_396,In_592);
and U84 (N_84,In_18,In_617);
xor U85 (N_85,In_923,In_200);
and U86 (N_86,In_50,In_108);
xnor U87 (N_87,In_718,In_596);
xor U88 (N_88,In_562,In_773);
xor U89 (N_89,In_892,In_332);
xnor U90 (N_90,In_161,In_671);
or U91 (N_91,In_966,In_226);
nor U92 (N_92,In_731,In_586);
and U93 (N_93,In_620,In_330);
nand U94 (N_94,In_183,In_782);
xnor U95 (N_95,In_908,In_737);
or U96 (N_96,In_975,In_745);
xnor U97 (N_97,In_256,In_629);
nor U98 (N_98,In_286,In_94);
and U99 (N_99,In_198,In_688);
nor U100 (N_100,In_932,In_626);
xnor U101 (N_101,In_119,In_187);
nand U102 (N_102,In_572,In_751);
or U103 (N_103,In_947,In_143);
xor U104 (N_104,In_278,In_93);
nor U105 (N_105,In_995,In_730);
and U106 (N_106,In_827,In_867);
or U107 (N_107,In_453,In_110);
nor U108 (N_108,In_554,In_451);
and U109 (N_109,In_700,In_138);
and U110 (N_110,In_771,In_69);
and U111 (N_111,In_759,In_548);
and U112 (N_112,In_766,In_103);
or U113 (N_113,In_416,In_502);
xnor U114 (N_114,In_447,In_566);
xor U115 (N_115,In_232,In_507);
nand U116 (N_116,In_266,In_503);
and U117 (N_117,In_281,In_939);
nor U118 (N_118,In_40,In_28);
nor U119 (N_119,In_153,In_725);
xor U120 (N_120,In_715,In_692);
and U121 (N_121,In_314,In_925);
or U122 (N_122,In_400,In_466);
or U123 (N_123,In_984,In_68);
or U124 (N_124,In_91,In_943);
and U125 (N_125,In_564,In_231);
nand U126 (N_126,In_515,In_918);
nor U127 (N_127,In_55,In_269);
nand U128 (N_128,In_765,In_853);
or U129 (N_129,In_916,In_207);
nand U130 (N_130,In_220,In_659);
nand U131 (N_131,In_633,In_215);
or U132 (N_132,In_533,In_129);
xor U133 (N_133,In_747,In_121);
nand U134 (N_134,In_537,In_905);
and U135 (N_135,In_437,In_238);
nand U136 (N_136,In_62,In_393);
nor U137 (N_137,In_710,In_574);
or U138 (N_138,In_17,In_399);
and U139 (N_139,In_599,In_112);
nand U140 (N_140,In_824,In_848);
and U141 (N_141,In_397,In_666);
or U142 (N_142,In_970,In_670);
nand U143 (N_143,In_127,In_317);
or U144 (N_144,In_783,In_216);
nor U145 (N_145,In_409,In_699);
nand U146 (N_146,In_77,In_435);
and U147 (N_147,In_561,In_817);
xnor U148 (N_148,In_974,In_170);
nor U149 (N_149,In_37,In_263);
nand U150 (N_150,In_775,In_168);
or U151 (N_151,In_799,In_444);
nand U152 (N_152,In_850,In_21);
nand U153 (N_153,In_883,In_346);
and U154 (N_154,In_282,In_547);
nor U155 (N_155,In_97,In_358);
or U156 (N_156,In_792,In_29);
xnor U157 (N_157,In_377,In_211);
nand U158 (N_158,In_880,In_615);
nor U159 (N_159,In_74,In_307);
nor U160 (N_160,In_863,In_5);
xnor U161 (N_161,In_627,In_556);
nor U162 (N_162,In_856,In_910);
xor U163 (N_163,In_308,In_582);
or U164 (N_164,In_54,In_272);
and U165 (N_165,In_808,In_162);
or U166 (N_166,In_870,In_949);
and U167 (N_167,In_839,In_696);
nand U168 (N_168,In_640,In_495);
nand U169 (N_169,In_944,In_496);
xor U170 (N_170,In_965,In_937);
or U171 (N_171,In_293,In_519);
nor U172 (N_172,In_4,In_151);
xor U173 (N_173,In_900,In_147);
or U174 (N_174,In_988,In_229);
or U175 (N_175,In_770,In_237);
nor U176 (N_176,In_568,In_789);
xor U177 (N_177,In_541,In_487);
xor U178 (N_178,In_919,In_175);
xor U179 (N_179,In_128,In_316);
and U180 (N_180,In_679,In_525);
nand U181 (N_181,In_320,In_842);
nand U182 (N_182,In_876,In_977);
and U183 (N_183,In_489,In_875);
or U184 (N_184,In_218,In_102);
xnor U185 (N_185,In_834,In_36);
and U186 (N_186,In_166,In_189);
nand U187 (N_187,In_945,In_478);
nand U188 (N_188,In_419,In_90);
and U189 (N_189,In_604,In_854);
or U190 (N_190,In_449,In_296);
xor U191 (N_191,In_47,In_309);
nand U192 (N_192,In_878,In_811);
or U193 (N_193,In_92,In_407);
or U194 (N_194,In_99,In_15);
nor U195 (N_195,In_331,In_849);
nor U196 (N_196,In_764,In_980);
nand U197 (N_197,In_714,In_224);
xor U198 (N_198,In_376,In_440);
or U199 (N_199,In_148,In_532);
nor U200 (N_200,In_899,In_906);
or U201 (N_201,In_903,In_322);
nand U202 (N_202,In_549,In_504);
or U203 (N_203,In_433,In_46);
xor U204 (N_204,In_647,In_342);
xor U205 (N_205,In_347,In_101);
or U206 (N_206,In_378,In_134);
xor U207 (N_207,In_881,In_621);
and U208 (N_208,In_669,In_821);
xor U209 (N_209,In_902,In_914);
or U210 (N_210,In_459,In_978);
or U211 (N_211,In_202,In_705);
or U212 (N_212,In_690,In_78);
nand U213 (N_213,In_911,In_401);
and U214 (N_214,In_753,In_605);
and U215 (N_215,In_135,In_571);
or U216 (N_216,In_368,In_420);
nand U217 (N_217,In_897,In_831);
and U218 (N_218,In_774,In_38);
xnor U219 (N_219,In_847,In_823);
and U220 (N_220,In_157,In_122);
xnor U221 (N_221,In_105,In_559);
or U222 (N_222,In_412,In_868);
nor U223 (N_223,In_830,In_423);
nor U224 (N_224,In_536,In_501);
and U225 (N_225,In_221,In_565);
nand U226 (N_226,In_512,In_841);
xor U227 (N_227,In_191,In_860);
nor U228 (N_228,In_362,In_171);
nand U229 (N_229,In_461,In_467);
or U230 (N_230,In_19,In_934);
xnor U231 (N_231,In_245,In_20);
or U232 (N_232,In_154,In_382);
and U233 (N_233,In_355,In_472);
nand U234 (N_234,In_740,In_645);
and U235 (N_235,In_927,In_380);
or U236 (N_236,In_363,In_846);
nand U237 (N_237,In_476,In_510);
and U238 (N_238,In_668,In_323);
and U239 (N_239,In_832,In_370);
and U240 (N_240,In_257,In_426);
nor U241 (N_241,In_521,In_194);
and U242 (N_242,In_624,In_720);
and U243 (N_243,In_124,In_252);
or U244 (N_244,In_722,In_131);
or U245 (N_245,In_356,In_780);
or U246 (N_246,In_294,In_610);
and U247 (N_247,In_815,In_219);
nor U248 (N_248,In_594,In_760);
nand U249 (N_249,In_391,In_369);
and U250 (N_250,In_637,In_96);
xor U251 (N_251,In_702,In_804);
and U252 (N_252,In_809,In_732);
xnor U253 (N_253,In_283,In_754);
nor U254 (N_254,In_82,In_155);
xor U255 (N_255,In_819,In_711);
or U256 (N_256,In_374,In_540);
nor U257 (N_257,In_492,In_648);
xnor U258 (N_258,In_2,In_338);
and U259 (N_259,In_528,In_836);
or U260 (N_260,In_588,In_682);
and U261 (N_261,In_468,In_383);
or U262 (N_262,In_743,In_595);
and U263 (N_263,In_26,In_408);
and U264 (N_264,In_3,In_104);
and U265 (N_265,In_404,In_201);
nor U266 (N_266,In_681,In_336);
and U267 (N_267,In_655,In_417);
nand U268 (N_268,In_244,In_150);
xnor U269 (N_269,In_584,In_81);
nor U270 (N_270,In_247,In_334);
and U271 (N_271,In_884,In_511);
or U272 (N_272,In_434,In_805);
and U273 (N_273,In_341,In_852);
and U274 (N_274,In_276,In_284);
xor U275 (N_275,In_79,In_776);
nor U276 (N_276,In_886,In_538);
xor U277 (N_277,In_190,In_635);
and U278 (N_278,In_814,In_845);
or U279 (N_279,In_872,In_136);
nor U280 (N_280,In_694,In_287);
and U281 (N_281,In_664,In_208);
nor U282 (N_282,In_513,In_777);
nor U283 (N_283,In_518,In_195);
and U284 (N_284,In_750,In_680);
nand U285 (N_285,In_508,In_176);
nand U286 (N_286,In_583,In_357);
nor U287 (N_287,In_630,In_701);
or U288 (N_288,In_60,In_455);
or U289 (N_289,In_969,In_545);
or U290 (N_290,In_9,In_994);
nor U291 (N_291,In_313,In_738);
and U292 (N_292,In_563,In_844);
nand U293 (N_293,In_593,In_768);
or U294 (N_294,In_921,In_784);
and U295 (N_295,In_798,In_490);
or U296 (N_296,In_479,In_797);
and U297 (N_297,In_673,In_953);
or U298 (N_298,In_552,In_591);
nand U299 (N_299,In_462,In_100);
or U300 (N_300,In_608,In_203);
nor U301 (N_301,In_858,In_749);
nor U302 (N_302,In_644,In_310);
nand U303 (N_303,In_813,In_418);
nor U304 (N_304,In_430,In_70);
nor U305 (N_305,In_53,In_113);
nand U306 (N_306,In_172,In_7);
or U307 (N_307,In_274,In_49);
nor U308 (N_308,In_106,In_952);
xnor U309 (N_309,In_182,In_998);
or U310 (N_310,In_422,In_303);
nor U311 (N_311,In_810,In_851);
nand U312 (N_312,In_111,In_885);
or U313 (N_313,In_289,In_439);
nand U314 (N_314,In_958,In_243);
xor U315 (N_315,In_178,In_360);
or U316 (N_316,In_390,In_935);
xor U317 (N_317,In_835,In_299);
or U318 (N_318,In_411,In_653);
xor U319 (N_319,In_184,In_879);
nand U320 (N_320,In_117,In_985);
or U321 (N_321,In_506,In_526);
nor U322 (N_322,In_838,In_546);
or U323 (N_323,In_758,In_260);
or U324 (N_324,In_139,In_857);
nor U325 (N_325,In_855,In_375);
or U326 (N_326,In_114,In_398);
and U327 (N_327,In_56,In_372);
nand U328 (N_328,In_406,In_597);
xor U329 (N_329,In_144,In_75);
and U330 (N_330,In_405,In_0);
and U331 (N_331,In_891,In_385);
or U332 (N_332,In_589,In_991);
nor U333 (N_333,In_522,In_448);
nand U334 (N_334,In_733,In_329);
xor U335 (N_335,In_149,In_280);
and U336 (N_336,In_180,In_895);
nor U337 (N_337,In_165,In_348);
nor U338 (N_338,In_712,In_199);
nor U339 (N_339,In_457,In_491);
and U340 (N_340,In_651,In_454);
nand U341 (N_341,In_217,In_661);
and U342 (N_342,In_475,In_188);
nor U343 (N_343,In_442,In_109);
nand U344 (N_344,In_126,In_689);
and U345 (N_345,In_581,In_865);
and U346 (N_346,In_946,In_788);
nand U347 (N_347,In_44,In_793);
or U348 (N_348,In_163,In_598);
or U349 (N_349,In_729,In_115);
nand U350 (N_350,In_928,In_734);
or U351 (N_351,In_606,In_486);
and U352 (N_352,In_622,In_312);
xor U353 (N_353,In_972,In_781);
nor U354 (N_354,In_901,In_523);
or U355 (N_355,In_728,In_654);
xor U356 (N_356,In_578,In_253);
xnor U357 (N_357,In_477,In_748);
nand U358 (N_358,In_570,In_636);
xnor U359 (N_359,In_638,In_223);
or U360 (N_360,In_107,In_337);
xnor U361 (N_361,In_288,In_590);
and U362 (N_362,In_663,In_632);
and U363 (N_363,In_576,In_463);
xnor U364 (N_364,In_826,In_233);
xor U365 (N_365,In_912,In_31);
nor U366 (N_366,In_505,In_353);
xnor U367 (N_367,In_98,In_667);
nor U368 (N_368,In_277,In_926);
xnor U369 (N_369,In_707,In_941);
xnor U370 (N_370,In_41,In_882);
xnor U371 (N_371,In_675,In_305);
nor U372 (N_372,In_140,In_302);
and U373 (N_373,In_735,In_874);
nand U374 (N_374,In_602,In_268);
and U375 (N_375,In_429,In_837);
xnor U376 (N_376,In_394,In_324);
and U377 (N_377,In_801,In_973);
nand U378 (N_378,In_116,In_613);
or U379 (N_379,In_196,In_822);
nor U380 (N_380,In_787,In_806);
xnor U381 (N_381,In_460,In_315);
nor U382 (N_382,In_960,In_614);
xnor U383 (N_383,In_123,In_672);
nand U384 (N_384,In_255,In_132);
and U385 (N_385,In_388,In_600);
nand U386 (N_386,In_577,In_657);
nand U387 (N_387,In_704,In_752);
or U388 (N_388,In_993,In_210);
and U389 (N_389,In_924,In_959);
or U390 (N_390,In_685,In_786);
nand U391 (N_391,In_65,In_275);
nor U392 (N_392,In_950,In_697);
nor U393 (N_393,In_982,In_968);
and U394 (N_394,In_962,In_634);
xnor U395 (N_395,In_543,In_989);
and U396 (N_396,In_76,In_803);
nand U397 (N_397,In_352,In_146);
nor U398 (N_398,In_524,In_328);
xor U399 (N_399,In_192,In_441);
or U400 (N_400,In_241,In_361);
and U401 (N_401,In_642,In_130);
xnor U402 (N_402,In_996,In_392);
nand U403 (N_403,In_807,In_790);
nor U404 (N_404,In_8,In_990);
xor U405 (N_405,In_443,In_739);
nand U406 (N_406,In_343,In_558);
nor U407 (N_407,In_986,In_557);
and U408 (N_408,In_493,In_954);
nor U409 (N_409,In_726,In_160);
nor U410 (N_410,In_234,In_88);
nand U411 (N_411,In_961,In_32);
and U412 (N_412,In_480,In_51);
xor U413 (N_413,In_530,In_249);
and U414 (N_414,In_888,In_141);
nor U415 (N_415,In_421,In_193);
and U416 (N_416,In_861,In_723);
xnor U417 (N_417,In_942,In_650);
or U418 (N_418,In_785,In_550);
nand U419 (N_419,In_213,In_242);
xnor U420 (N_420,In_239,In_57);
nand U421 (N_421,In_222,In_517);
and U422 (N_422,In_59,In_291);
nand U423 (N_423,In_611,In_938);
xor U424 (N_424,In_763,In_24);
nor U425 (N_425,In_618,In_354);
or U426 (N_426,In_560,In_717);
nor U427 (N_427,In_297,In_371);
nand U428 (N_428,In_713,In_779);
xor U429 (N_429,In_649,In_156);
xor U430 (N_430,In_465,In_13);
nor U431 (N_431,In_250,In_656);
and U432 (N_432,In_379,In_956);
nand U433 (N_433,In_708,In_16);
nor U434 (N_434,In_709,In_497);
and U435 (N_435,In_981,In_922);
and U436 (N_436,In_340,In_551);
nand U437 (N_437,In_367,In_473);
or U438 (N_438,In_625,In_349);
nor U439 (N_439,In_818,In_509);
nand U440 (N_440,In_279,In_520);
nand U441 (N_441,In_169,In_87);
nand U442 (N_442,In_333,In_52);
nor U443 (N_443,In_95,In_84);
nor U444 (N_444,In_365,In_873);
or U445 (N_445,In_158,In_414);
or U446 (N_446,In_964,In_864);
or U447 (N_447,In_544,In_43);
xor U448 (N_448,In_488,In_167);
xnor U449 (N_449,In_66,In_951);
nand U450 (N_450,In_254,In_869);
nor U451 (N_451,In_967,In_125);
xnor U452 (N_452,In_890,In_778);
or U453 (N_453,In_474,In_185);
nand U454 (N_454,In_601,In_179);
nand U455 (N_455,In_270,In_762);
xor U456 (N_456,In_514,In_772);
and U457 (N_457,In_344,In_271);
xnor U458 (N_458,In_820,In_427);
xor U459 (N_459,In_746,In_366);
and U460 (N_460,In_225,In_204);
or U461 (N_461,In_698,In_63);
and U462 (N_462,In_22,In_228);
nor U463 (N_463,In_757,In_662);
nand U464 (N_464,In_612,In_12);
nand U465 (N_465,In_10,In_706);
nor U466 (N_466,In_471,In_415);
or U467 (N_467,In_424,In_796);
and U468 (N_468,In_235,In_246);
xor U469 (N_469,In_862,In_575);
xor U470 (N_470,In_684,In_623);
xnor U471 (N_471,In_428,In_527);
nand U472 (N_472,In_791,In_470);
or U473 (N_473,In_327,In_381);
and U474 (N_474,In_955,In_335);
or U475 (N_475,In_212,In_214);
nand U476 (N_476,In_719,In_425);
nand U477 (N_477,In_436,In_940);
and U478 (N_478,In_643,In_579);
nand U479 (N_479,In_812,In_181);
nor U480 (N_480,In_628,In_871);
nor U481 (N_481,In_456,In_929);
nand U482 (N_482,In_983,In_339);
xor U483 (N_483,In_72,In_913);
and U484 (N_484,In_917,In_186);
and U485 (N_485,In_413,In_587);
nor U486 (N_486,In_555,In_42);
xnor U487 (N_487,In_724,In_736);
and U488 (N_488,In_904,In_877);
or U489 (N_489,In_446,In_894);
xnor U490 (N_490,In_458,In_445);
or U491 (N_491,In_619,In_609);
and U492 (N_492,In_205,In_641);
nand U493 (N_493,In_567,In_431);
or U494 (N_494,In_607,In_744);
nand U495 (N_495,In_639,In_206);
nor U496 (N_496,In_687,In_39);
nor U497 (N_497,In_742,In_727);
and U498 (N_498,In_83,In_741);
nor U499 (N_499,In_484,In_573);
nand U500 (N_500,N_493,N_307);
xnor U501 (N_501,N_211,N_375);
and U502 (N_502,N_97,N_248);
or U503 (N_503,N_132,N_356);
xor U504 (N_504,N_325,N_62);
and U505 (N_505,N_368,N_155);
or U506 (N_506,N_227,N_498);
xor U507 (N_507,N_321,N_203);
or U508 (N_508,N_401,N_138);
xor U509 (N_509,N_428,N_96);
xor U510 (N_510,N_295,N_141);
nor U511 (N_511,N_3,N_188);
nor U512 (N_512,N_404,N_56);
xor U513 (N_513,N_250,N_270);
xnor U514 (N_514,N_350,N_335);
nand U515 (N_515,N_158,N_165);
and U516 (N_516,N_216,N_242);
and U517 (N_517,N_137,N_492);
or U518 (N_518,N_148,N_84);
nor U519 (N_519,N_59,N_2);
and U520 (N_520,N_71,N_127);
xor U521 (N_521,N_433,N_16);
and U522 (N_522,N_277,N_414);
nor U523 (N_523,N_247,N_479);
and U524 (N_524,N_345,N_457);
or U525 (N_525,N_6,N_175);
or U526 (N_526,N_394,N_234);
nand U527 (N_527,N_108,N_347);
or U528 (N_528,N_205,N_218);
nor U529 (N_529,N_66,N_301);
xnor U530 (N_530,N_320,N_448);
nor U531 (N_531,N_495,N_147);
and U532 (N_532,N_109,N_252);
xnor U533 (N_533,N_161,N_40);
nor U534 (N_534,N_432,N_5);
nand U535 (N_535,N_213,N_27);
or U536 (N_536,N_11,N_463);
nor U537 (N_537,N_131,N_288);
nand U538 (N_538,N_456,N_14);
xnor U539 (N_539,N_53,N_225);
nor U540 (N_540,N_219,N_346);
and U541 (N_541,N_51,N_263);
nand U542 (N_542,N_387,N_173);
nand U543 (N_543,N_180,N_371);
xnor U544 (N_544,N_296,N_358);
xor U545 (N_545,N_76,N_224);
or U546 (N_546,N_251,N_168);
xor U547 (N_547,N_69,N_65);
and U548 (N_548,N_171,N_133);
nor U549 (N_549,N_145,N_440);
and U550 (N_550,N_260,N_489);
nand U551 (N_551,N_476,N_82);
nand U552 (N_552,N_328,N_123);
and U553 (N_553,N_67,N_149);
and U554 (N_554,N_402,N_395);
nand U555 (N_555,N_327,N_336);
nor U556 (N_556,N_119,N_7);
and U557 (N_557,N_416,N_300);
xor U558 (N_558,N_88,N_241);
xnor U559 (N_559,N_160,N_409);
nor U560 (N_560,N_343,N_391);
and U561 (N_561,N_272,N_298);
and U562 (N_562,N_421,N_264);
nand U563 (N_563,N_112,N_129);
xor U564 (N_564,N_130,N_118);
and U565 (N_565,N_172,N_232);
nand U566 (N_566,N_1,N_243);
or U567 (N_567,N_196,N_284);
xor U568 (N_568,N_355,N_61);
nand U569 (N_569,N_128,N_318);
and U570 (N_570,N_192,N_342);
nand U571 (N_571,N_309,N_326);
xor U572 (N_572,N_93,N_255);
nand U573 (N_573,N_156,N_41);
nor U574 (N_574,N_177,N_72);
and U575 (N_575,N_50,N_310);
or U576 (N_576,N_73,N_437);
xnor U577 (N_577,N_446,N_338);
xnor U578 (N_578,N_89,N_245);
and U579 (N_579,N_68,N_386);
or U580 (N_580,N_208,N_229);
nor U581 (N_581,N_206,N_434);
and U582 (N_582,N_254,N_302);
nand U583 (N_583,N_114,N_262);
xnor U584 (N_584,N_366,N_42);
or U585 (N_585,N_266,N_392);
xor U586 (N_586,N_98,N_238);
nand U587 (N_587,N_222,N_329);
nand U588 (N_588,N_190,N_441);
xor U589 (N_589,N_44,N_341);
nor U590 (N_590,N_289,N_267);
or U591 (N_591,N_33,N_210);
nor U592 (N_592,N_367,N_55);
xnor U593 (N_593,N_236,N_166);
xnor U594 (N_594,N_484,N_85);
and U595 (N_595,N_36,N_458);
and U596 (N_596,N_87,N_223);
and U597 (N_597,N_363,N_430);
nand U598 (N_598,N_348,N_101);
nor U599 (N_599,N_439,N_269);
and U600 (N_600,N_58,N_120);
xor U601 (N_601,N_461,N_151);
nor U602 (N_602,N_417,N_377);
xor U603 (N_603,N_285,N_103);
and U604 (N_604,N_80,N_246);
or U605 (N_605,N_94,N_212);
xor U606 (N_606,N_146,N_256);
and U607 (N_607,N_418,N_316);
or U608 (N_608,N_372,N_46);
and U609 (N_609,N_468,N_60);
nor U610 (N_610,N_423,N_75);
or U611 (N_611,N_322,N_469);
or U612 (N_612,N_273,N_426);
and U613 (N_613,N_201,N_104);
nand U614 (N_614,N_150,N_275);
xnor U615 (N_615,N_233,N_249);
or U616 (N_616,N_305,N_344);
or U617 (N_617,N_81,N_390);
nor U618 (N_618,N_78,N_47);
nand U619 (N_619,N_235,N_91);
and U620 (N_620,N_189,N_239);
and U621 (N_621,N_497,N_220);
nor U622 (N_622,N_185,N_195);
or U623 (N_623,N_162,N_429);
and U624 (N_624,N_373,N_444);
nor U625 (N_625,N_12,N_125);
and U626 (N_626,N_200,N_420);
nand U627 (N_627,N_351,N_228);
nor U628 (N_628,N_369,N_370);
and U629 (N_629,N_317,N_281);
nor U630 (N_630,N_257,N_470);
and U631 (N_631,N_28,N_465);
and U632 (N_632,N_349,N_265);
xor U633 (N_633,N_202,N_452);
or U634 (N_634,N_293,N_276);
nor U635 (N_635,N_453,N_475);
xor U636 (N_636,N_261,N_140);
nor U637 (N_637,N_31,N_306);
nand U638 (N_638,N_226,N_477);
nor U639 (N_639,N_63,N_334);
xnor U640 (N_640,N_279,N_411);
nor U641 (N_641,N_32,N_384);
nand U642 (N_642,N_435,N_126);
and U643 (N_643,N_396,N_198);
xor U644 (N_644,N_193,N_186);
xnor U645 (N_645,N_111,N_214);
xor U646 (N_646,N_354,N_385);
xor U647 (N_647,N_70,N_100);
nor U648 (N_648,N_481,N_17);
or U649 (N_649,N_122,N_333);
nand U650 (N_650,N_121,N_464);
nor U651 (N_651,N_74,N_454);
xnor U652 (N_652,N_378,N_451);
xnor U653 (N_653,N_25,N_178);
and U654 (N_654,N_144,N_142);
nor U655 (N_655,N_4,N_379);
nor U656 (N_656,N_187,N_174);
or U657 (N_657,N_331,N_244);
nor U658 (N_658,N_412,N_135);
or U659 (N_659,N_34,N_37);
or U660 (N_660,N_134,N_380);
and U661 (N_661,N_291,N_92);
xnor U662 (N_662,N_191,N_442);
nand U663 (N_663,N_436,N_106);
and U664 (N_664,N_313,N_480);
and U665 (N_665,N_443,N_39);
nor U666 (N_666,N_8,N_447);
and U667 (N_667,N_381,N_398);
nand U668 (N_668,N_183,N_54);
nor U669 (N_669,N_374,N_20);
nor U670 (N_670,N_410,N_405);
xor U671 (N_671,N_207,N_107);
nand U672 (N_672,N_319,N_115);
and U673 (N_673,N_268,N_10);
or U674 (N_674,N_176,N_152);
or U675 (N_675,N_153,N_15);
nand U676 (N_676,N_491,N_460);
or U677 (N_677,N_340,N_167);
and U678 (N_678,N_376,N_332);
nand U679 (N_679,N_286,N_0);
nor U680 (N_680,N_474,N_312);
and U681 (N_681,N_455,N_294);
nor U682 (N_682,N_314,N_399);
xor U683 (N_683,N_365,N_159);
and U684 (N_684,N_330,N_154);
or U685 (N_685,N_360,N_353);
and U686 (N_686,N_95,N_215);
and U687 (N_687,N_164,N_482);
nand U688 (N_688,N_424,N_18);
and U689 (N_689,N_311,N_494);
and U690 (N_690,N_304,N_19);
xnor U691 (N_691,N_445,N_184);
nor U692 (N_692,N_240,N_466);
nand U693 (N_693,N_48,N_413);
or U694 (N_694,N_357,N_221);
and U695 (N_695,N_170,N_79);
or U696 (N_696,N_86,N_315);
and U697 (N_697,N_449,N_419);
nand U698 (N_698,N_179,N_139);
nand U699 (N_699,N_487,N_471);
xnor U700 (N_700,N_283,N_397);
nand U701 (N_701,N_499,N_393);
nand U702 (N_702,N_431,N_303);
xnor U703 (N_703,N_105,N_230);
or U704 (N_704,N_462,N_362);
nor U705 (N_705,N_259,N_64);
or U706 (N_706,N_278,N_486);
xnor U707 (N_707,N_485,N_258);
and U708 (N_708,N_299,N_90);
nor U709 (N_709,N_467,N_157);
nor U710 (N_710,N_117,N_483);
or U711 (N_711,N_21,N_297);
or U712 (N_712,N_361,N_77);
xnor U713 (N_713,N_49,N_422);
xnor U714 (N_714,N_24,N_163);
and U715 (N_715,N_490,N_181);
nor U716 (N_716,N_339,N_406);
nor U717 (N_717,N_83,N_408);
or U718 (N_718,N_450,N_427);
or U719 (N_719,N_237,N_13);
nor U720 (N_720,N_102,N_364);
nor U721 (N_721,N_274,N_308);
nor U722 (N_722,N_52,N_271);
xor U723 (N_723,N_382,N_359);
nand U724 (N_724,N_472,N_38);
and U725 (N_725,N_57,N_438);
and U726 (N_726,N_110,N_99);
nor U727 (N_727,N_388,N_352);
and U728 (N_728,N_199,N_113);
or U729 (N_729,N_407,N_478);
or U730 (N_730,N_323,N_136);
and U731 (N_731,N_425,N_290);
nand U732 (N_732,N_9,N_292);
and U733 (N_733,N_337,N_473);
or U734 (N_734,N_204,N_282);
nor U735 (N_735,N_287,N_488);
xor U736 (N_736,N_280,N_209);
and U737 (N_737,N_415,N_29);
and U738 (N_738,N_45,N_324);
nand U739 (N_739,N_231,N_26);
and U740 (N_740,N_496,N_197);
nor U741 (N_741,N_253,N_217);
or U742 (N_742,N_169,N_124);
nand U743 (N_743,N_30,N_23);
or U744 (N_744,N_389,N_383);
nand U745 (N_745,N_22,N_182);
nor U746 (N_746,N_194,N_459);
xnor U747 (N_747,N_403,N_400);
xor U748 (N_748,N_43,N_143);
nand U749 (N_749,N_35,N_116);
or U750 (N_750,N_169,N_254);
or U751 (N_751,N_455,N_356);
nor U752 (N_752,N_310,N_499);
xor U753 (N_753,N_135,N_320);
and U754 (N_754,N_435,N_312);
or U755 (N_755,N_334,N_389);
nand U756 (N_756,N_289,N_177);
or U757 (N_757,N_248,N_165);
xor U758 (N_758,N_377,N_401);
and U759 (N_759,N_282,N_471);
xor U760 (N_760,N_29,N_378);
and U761 (N_761,N_461,N_317);
and U762 (N_762,N_247,N_310);
xor U763 (N_763,N_111,N_98);
and U764 (N_764,N_325,N_162);
nor U765 (N_765,N_308,N_87);
nor U766 (N_766,N_437,N_286);
and U767 (N_767,N_111,N_367);
nor U768 (N_768,N_253,N_52);
and U769 (N_769,N_137,N_71);
or U770 (N_770,N_257,N_171);
xor U771 (N_771,N_343,N_462);
or U772 (N_772,N_476,N_273);
nand U773 (N_773,N_394,N_414);
or U774 (N_774,N_394,N_121);
nand U775 (N_775,N_322,N_328);
xnor U776 (N_776,N_97,N_30);
nor U777 (N_777,N_484,N_447);
and U778 (N_778,N_407,N_219);
xor U779 (N_779,N_85,N_32);
and U780 (N_780,N_38,N_42);
nor U781 (N_781,N_49,N_443);
xnor U782 (N_782,N_446,N_250);
xor U783 (N_783,N_181,N_57);
nor U784 (N_784,N_464,N_336);
nor U785 (N_785,N_396,N_131);
nand U786 (N_786,N_72,N_282);
or U787 (N_787,N_242,N_413);
nor U788 (N_788,N_99,N_47);
nor U789 (N_789,N_93,N_281);
xnor U790 (N_790,N_349,N_386);
xor U791 (N_791,N_472,N_231);
or U792 (N_792,N_52,N_296);
and U793 (N_793,N_212,N_336);
xor U794 (N_794,N_259,N_30);
nand U795 (N_795,N_433,N_184);
and U796 (N_796,N_133,N_124);
nand U797 (N_797,N_321,N_424);
nor U798 (N_798,N_135,N_236);
nand U799 (N_799,N_470,N_405);
nor U800 (N_800,N_418,N_173);
nor U801 (N_801,N_460,N_160);
or U802 (N_802,N_487,N_459);
xnor U803 (N_803,N_114,N_215);
or U804 (N_804,N_257,N_212);
or U805 (N_805,N_497,N_223);
and U806 (N_806,N_262,N_186);
xor U807 (N_807,N_20,N_493);
xor U808 (N_808,N_106,N_364);
nand U809 (N_809,N_317,N_495);
nor U810 (N_810,N_122,N_94);
nand U811 (N_811,N_302,N_44);
nand U812 (N_812,N_229,N_255);
xnor U813 (N_813,N_196,N_378);
nand U814 (N_814,N_39,N_419);
xnor U815 (N_815,N_267,N_131);
nor U816 (N_816,N_235,N_399);
xor U817 (N_817,N_209,N_400);
or U818 (N_818,N_489,N_127);
and U819 (N_819,N_201,N_297);
nand U820 (N_820,N_224,N_101);
and U821 (N_821,N_6,N_49);
and U822 (N_822,N_55,N_58);
nand U823 (N_823,N_9,N_10);
or U824 (N_824,N_195,N_484);
nand U825 (N_825,N_301,N_2);
xor U826 (N_826,N_122,N_104);
nand U827 (N_827,N_65,N_77);
nand U828 (N_828,N_284,N_329);
xnor U829 (N_829,N_250,N_301);
or U830 (N_830,N_469,N_181);
or U831 (N_831,N_192,N_22);
xor U832 (N_832,N_310,N_441);
nor U833 (N_833,N_325,N_418);
xor U834 (N_834,N_183,N_239);
xor U835 (N_835,N_122,N_131);
nor U836 (N_836,N_417,N_27);
xnor U837 (N_837,N_467,N_297);
xor U838 (N_838,N_194,N_406);
or U839 (N_839,N_32,N_229);
and U840 (N_840,N_412,N_60);
nor U841 (N_841,N_39,N_452);
and U842 (N_842,N_50,N_187);
and U843 (N_843,N_371,N_189);
or U844 (N_844,N_33,N_231);
nand U845 (N_845,N_371,N_340);
nand U846 (N_846,N_391,N_44);
and U847 (N_847,N_62,N_348);
and U848 (N_848,N_278,N_12);
or U849 (N_849,N_109,N_184);
and U850 (N_850,N_370,N_408);
nand U851 (N_851,N_88,N_198);
xnor U852 (N_852,N_328,N_432);
xor U853 (N_853,N_267,N_446);
or U854 (N_854,N_353,N_359);
nand U855 (N_855,N_45,N_461);
or U856 (N_856,N_220,N_328);
and U857 (N_857,N_434,N_184);
and U858 (N_858,N_11,N_44);
nor U859 (N_859,N_392,N_11);
nor U860 (N_860,N_121,N_150);
and U861 (N_861,N_174,N_7);
xnor U862 (N_862,N_319,N_281);
or U863 (N_863,N_266,N_386);
nor U864 (N_864,N_258,N_51);
nand U865 (N_865,N_388,N_151);
xnor U866 (N_866,N_414,N_153);
nor U867 (N_867,N_69,N_319);
nor U868 (N_868,N_302,N_222);
nor U869 (N_869,N_459,N_156);
or U870 (N_870,N_130,N_473);
and U871 (N_871,N_106,N_420);
xnor U872 (N_872,N_337,N_153);
nor U873 (N_873,N_48,N_155);
and U874 (N_874,N_251,N_177);
or U875 (N_875,N_352,N_5);
nand U876 (N_876,N_8,N_488);
xor U877 (N_877,N_490,N_443);
xor U878 (N_878,N_262,N_51);
or U879 (N_879,N_463,N_235);
and U880 (N_880,N_402,N_455);
or U881 (N_881,N_374,N_346);
nand U882 (N_882,N_326,N_266);
nand U883 (N_883,N_455,N_82);
nor U884 (N_884,N_200,N_444);
or U885 (N_885,N_244,N_426);
or U886 (N_886,N_103,N_378);
xor U887 (N_887,N_356,N_464);
nand U888 (N_888,N_102,N_280);
and U889 (N_889,N_259,N_49);
xnor U890 (N_890,N_428,N_202);
nand U891 (N_891,N_238,N_247);
and U892 (N_892,N_301,N_241);
and U893 (N_893,N_286,N_220);
and U894 (N_894,N_161,N_333);
and U895 (N_895,N_144,N_367);
and U896 (N_896,N_91,N_426);
nor U897 (N_897,N_126,N_107);
xnor U898 (N_898,N_133,N_409);
nand U899 (N_899,N_141,N_349);
xnor U900 (N_900,N_425,N_343);
and U901 (N_901,N_407,N_154);
nor U902 (N_902,N_302,N_292);
xnor U903 (N_903,N_156,N_449);
nor U904 (N_904,N_229,N_422);
xnor U905 (N_905,N_151,N_477);
and U906 (N_906,N_178,N_405);
or U907 (N_907,N_458,N_369);
xor U908 (N_908,N_380,N_492);
xnor U909 (N_909,N_9,N_495);
nand U910 (N_910,N_141,N_335);
xor U911 (N_911,N_277,N_475);
xor U912 (N_912,N_241,N_15);
and U913 (N_913,N_141,N_172);
xor U914 (N_914,N_1,N_102);
xor U915 (N_915,N_374,N_211);
xor U916 (N_916,N_498,N_418);
nand U917 (N_917,N_274,N_446);
and U918 (N_918,N_484,N_252);
nand U919 (N_919,N_463,N_403);
nand U920 (N_920,N_430,N_110);
or U921 (N_921,N_36,N_32);
nor U922 (N_922,N_453,N_193);
nand U923 (N_923,N_189,N_451);
xnor U924 (N_924,N_147,N_227);
nor U925 (N_925,N_209,N_258);
and U926 (N_926,N_116,N_342);
nand U927 (N_927,N_414,N_110);
and U928 (N_928,N_359,N_196);
or U929 (N_929,N_17,N_117);
or U930 (N_930,N_182,N_352);
xor U931 (N_931,N_142,N_90);
or U932 (N_932,N_472,N_428);
xnor U933 (N_933,N_154,N_364);
nor U934 (N_934,N_468,N_59);
and U935 (N_935,N_479,N_265);
and U936 (N_936,N_272,N_231);
and U937 (N_937,N_154,N_303);
xnor U938 (N_938,N_238,N_6);
or U939 (N_939,N_72,N_494);
xor U940 (N_940,N_155,N_264);
nand U941 (N_941,N_456,N_419);
nand U942 (N_942,N_488,N_123);
and U943 (N_943,N_105,N_468);
or U944 (N_944,N_246,N_202);
or U945 (N_945,N_217,N_254);
nor U946 (N_946,N_450,N_419);
or U947 (N_947,N_265,N_460);
nor U948 (N_948,N_20,N_368);
and U949 (N_949,N_209,N_351);
nand U950 (N_950,N_91,N_206);
nor U951 (N_951,N_163,N_246);
nor U952 (N_952,N_72,N_447);
xnor U953 (N_953,N_103,N_430);
nor U954 (N_954,N_380,N_475);
xor U955 (N_955,N_465,N_208);
or U956 (N_956,N_310,N_38);
or U957 (N_957,N_300,N_275);
xnor U958 (N_958,N_301,N_363);
xnor U959 (N_959,N_406,N_232);
nor U960 (N_960,N_177,N_252);
and U961 (N_961,N_37,N_172);
or U962 (N_962,N_143,N_181);
nand U963 (N_963,N_149,N_433);
and U964 (N_964,N_199,N_398);
nand U965 (N_965,N_368,N_35);
or U966 (N_966,N_92,N_30);
nor U967 (N_967,N_270,N_129);
and U968 (N_968,N_207,N_454);
nor U969 (N_969,N_184,N_145);
and U970 (N_970,N_215,N_393);
nand U971 (N_971,N_159,N_63);
nand U972 (N_972,N_427,N_127);
and U973 (N_973,N_146,N_391);
and U974 (N_974,N_381,N_168);
and U975 (N_975,N_119,N_424);
nand U976 (N_976,N_419,N_72);
nor U977 (N_977,N_98,N_446);
nor U978 (N_978,N_188,N_283);
and U979 (N_979,N_168,N_135);
nand U980 (N_980,N_289,N_355);
nor U981 (N_981,N_360,N_433);
xnor U982 (N_982,N_447,N_286);
nand U983 (N_983,N_73,N_384);
nand U984 (N_984,N_199,N_344);
or U985 (N_985,N_45,N_427);
xor U986 (N_986,N_410,N_109);
or U987 (N_987,N_244,N_369);
or U988 (N_988,N_7,N_493);
xnor U989 (N_989,N_93,N_360);
and U990 (N_990,N_149,N_178);
nand U991 (N_991,N_304,N_233);
nand U992 (N_992,N_35,N_416);
nand U993 (N_993,N_273,N_450);
xnor U994 (N_994,N_307,N_406);
and U995 (N_995,N_26,N_259);
nand U996 (N_996,N_218,N_276);
nor U997 (N_997,N_291,N_473);
or U998 (N_998,N_160,N_284);
nor U999 (N_999,N_8,N_97);
or U1000 (N_1000,N_774,N_627);
or U1001 (N_1001,N_554,N_725);
nor U1002 (N_1002,N_777,N_762);
and U1003 (N_1003,N_682,N_704);
nor U1004 (N_1004,N_826,N_874);
xnor U1005 (N_1005,N_688,N_800);
or U1006 (N_1006,N_972,N_693);
nor U1007 (N_1007,N_565,N_661);
nand U1008 (N_1008,N_644,N_843);
or U1009 (N_1009,N_651,N_946);
and U1010 (N_1010,N_775,N_541);
xnor U1011 (N_1011,N_809,N_765);
and U1012 (N_1012,N_860,N_539);
and U1013 (N_1013,N_957,N_700);
nand U1014 (N_1014,N_681,N_965);
and U1015 (N_1015,N_636,N_863);
and U1016 (N_1016,N_701,N_764);
xor U1017 (N_1017,N_572,N_746);
and U1018 (N_1018,N_550,N_755);
nor U1019 (N_1019,N_721,N_510);
xnor U1020 (N_1020,N_973,N_886);
nand U1021 (N_1021,N_632,N_538);
xnor U1022 (N_1022,N_571,N_989);
and U1023 (N_1023,N_808,N_859);
nor U1024 (N_1024,N_606,N_514);
nand U1025 (N_1025,N_730,N_828);
nor U1026 (N_1026,N_602,N_930);
or U1027 (N_1027,N_570,N_870);
nor U1028 (N_1028,N_903,N_729);
nor U1029 (N_1029,N_789,N_779);
nand U1030 (N_1030,N_821,N_824);
nand U1031 (N_1031,N_884,N_614);
or U1032 (N_1032,N_537,N_825);
nor U1033 (N_1033,N_502,N_898);
nor U1034 (N_1034,N_739,N_831);
and U1035 (N_1035,N_840,N_987);
nand U1036 (N_1036,N_761,N_677);
xnor U1037 (N_1037,N_519,N_995);
and U1038 (N_1038,N_668,N_861);
xnor U1039 (N_1039,N_592,N_735);
nor U1040 (N_1040,N_933,N_871);
or U1041 (N_1041,N_913,N_698);
nand U1042 (N_1042,N_782,N_689);
nand U1043 (N_1043,N_918,N_691);
nand U1044 (N_1044,N_937,N_696);
nor U1045 (N_1045,N_917,N_947);
or U1046 (N_1046,N_692,N_620);
and U1047 (N_1047,N_717,N_535);
or U1048 (N_1048,N_934,N_685);
or U1049 (N_1049,N_561,N_567);
or U1050 (N_1050,N_806,N_991);
and U1051 (N_1051,N_936,N_619);
nor U1052 (N_1052,N_798,N_635);
xor U1053 (N_1053,N_653,N_551);
nor U1054 (N_1054,N_659,N_842);
or U1055 (N_1055,N_815,N_885);
nor U1056 (N_1056,N_950,N_888);
or U1057 (N_1057,N_813,N_740);
xnor U1058 (N_1058,N_756,N_594);
nor U1059 (N_1059,N_734,N_747);
nor U1060 (N_1060,N_801,N_894);
xnor U1061 (N_1061,N_807,N_949);
and U1062 (N_1062,N_967,N_818);
or U1063 (N_1063,N_549,N_852);
and U1064 (N_1064,N_922,N_584);
nand U1065 (N_1065,N_948,N_679);
or U1066 (N_1066,N_683,N_736);
and U1067 (N_1067,N_643,N_770);
nand U1068 (N_1068,N_941,N_883);
nand U1069 (N_1069,N_568,N_797);
nor U1070 (N_1070,N_791,N_667);
nor U1071 (N_1071,N_992,N_545);
xor U1072 (N_1072,N_796,N_654);
nand U1073 (N_1073,N_556,N_881);
and U1074 (N_1074,N_981,N_626);
and U1075 (N_1075,N_858,N_846);
nor U1076 (N_1076,N_823,N_686);
xor U1077 (N_1077,N_799,N_687);
xnor U1078 (N_1078,N_942,N_641);
nor U1079 (N_1079,N_513,N_925);
nand U1080 (N_1080,N_910,N_999);
and U1081 (N_1081,N_562,N_805);
and U1082 (N_1082,N_601,N_959);
nand U1083 (N_1083,N_624,N_904);
nor U1084 (N_1084,N_962,N_715);
or U1085 (N_1085,N_508,N_994);
nor U1086 (N_1086,N_975,N_705);
xnor U1087 (N_1087,N_583,N_766);
and U1088 (N_1088,N_652,N_604);
xnor U1089 (N_1089,N_540,N_822);
nand U1090 (N_1090,N_605,N_776);
and U1091 (N_1091,N_684,N_882);
or U1092 (N_1092,N_971,N_889);
xnor U1093 (N_1093,N_811,N_866);
xnor U1094 (N_1094,N_678,N_986);
nor U1095 (N_1095,N_720,N_982);
nor U1096 (N_1096,N_945,N_623);
or U1097 (N_1097,N_517,N_956);
and U1098 (N_1098,N_980,N_613);
xor U1099 (N_1099,N_522,N_656);
nor U1100 (N_1100,N_996,N_841);
or U1101 (N_1101,N_763,N_964);
xor U1102 (N_1102,N_512,N_712);
nor U1103 (N_1103,N_820,N_585);
nor U1104 (N_1104,N_507,N_608);
nor U1105 (N_1105,N_836,N_768);
or U1106 (N_1106,N_771,N_915);
xnor U1107 (N_1107,N_690,N_914);
xor U1108 (N_1108,N_542,N_504);
or U1109 (N_1109,N_543,N_548);
and U1110 (N_1110,N_500,N_979);
or U1111 (N_1111,N_590,N_579);
xor U1112 (N_1112,N_607,N_629);
xnor U1113 (N_1113,N_530,N_639);
xnor U1114 (N_1114,N_680,N_521);
nand U1115 (N_1115,N_990,N_575);
or U1116 (N_1116,N_544,N_891);
xnor U1117 (N_1117,N_598,N_617);
nand U1118 (N_1118,N_829,N_560);
and U1119 (N_1119,N_976,N_812);
nand U1120 (N_1120,N_657,N_977);
nand U1121 (N_1121,N_878,N_753);
xor U1122 (N_1122,N_634,N_529);
and U1123 (N_1123,N_531,N_932);
xor U1124 (N_1124,N_612,N_788);
xor U1125 (N_1125,N_911,N_819);
xnor U1126 (N_1126,N_804,N_610);
nand U1127 (N_1127,N_928,N_781);
and U1128 (N_1128,N_912,N_961);
xor U1129 (N_1129,N_552,N_867);
nand U1130 (N_1130,N_640,N_926);
and U1131 (N_1131,N_752,N_618);
or U1132 (N_1132,N_837,N_616);
or U1133 (N_1133,N_719,N_877);
nand U1134 (N_1134,N_897,N_699);
nor U1135 (N_1135,N_650,N_713);
xor U1136 (N_1136,N_759,N_511);
or U1137 (N_1137,N_716,N_767);
nor U1138 (N_1138,N_649,N_662);
and U1139 (N_1139,N_576,N_953);
or U1140 (N_1140,N_710,N_940);
nand U1141 (N_1141,N_533,N_875);
and U1142 (N_1142,N_534,N_707);
or U1143 (N_1143,N_869,N_893);
and U1144 (N_1144,N_865,N_983);
nand U1145 (N_1145,N_527,N_833);
and U1146 (N_1146,N_666,N_553);
or U1147 (N_1147,N_974,N_939);
and U1148 (N_1148,N_603,N_827);
nand U1149 (N_1149,N_757,N_750);
nor U1150 (N_1150,N_726,N_851);
xnor U1151 (N_1151,N_890,N_853);
nand U1152 (N_1152,N_645,N_923);
and U1153 (N_1153,N_520,N_574);
xnor U1154 (N_1154,N_787,N_802);
or U1155 (N_1155,N_785,N_954);
nand U1156 (N_1156,N_773,N_960);
xnor U1157 (N_1157,N_742,N_839);
xnor U1158 (N_1158,N_563,N_966);
nor U1159 (N_1159,N_694,N_835);
nor U1160 (N_1160,N_745,N_929);
or U1161 (N_1161,N_803,N_525);
xnor U1162 (N_1162,N_648,N_708);
or U1163 (N_1163,N_862,N_834);
and U1164 (N_1164,N_738,N_921);
xor U1165 (N_1165,N_501,N_793);
nand U1166 (N_1166,N_783,N_864);
nand U1167 (N_1167,N_557,N_628);
nor U1168 (N_1168,N_581,N_615);
and U1169 (N_1169,N_792,N_887);
or U1170 (N_1170,N_951,N_952);
nor U1171 (N_1171,N_873,N_595);
or U1172 (N_1172,N_577,N_564);
and U1173 (N_1173,N_795,N_670);
nand U1174 (N_1174,N_969,N_532);
xnor U1175 (N_1175,N_943,N_896);
nor U1176 (N_1176,N_599,N_609);
nor U1177 (N_1177,N_855,N_856);
xor U1178 (N_1178,N_600,N_892);
and U1179 (N_1179,N_997,N_732);
xor U1180 (N_1180,N_630,N_676);
or U1181 (N_1181,N_963,N_523);
nor U1182 (N_1182,N_998,N_518);
nand U1183 (N_1183,N_727,N_978);
xnor U1184 (N_1184,N_728,N_944);
xor U1185 (N_1185,N_907,N_868);
and U1186 (N_1186,N_611,N_968);
xnor U1187 (N_1187,N_731,N_810);
or U1188 (N_1188,N_879,N_832);
nor U1189 (N_1189,N_637,N_931);
nor U1190 (N_1190,N_588,N_880);
and U1191 (N_1191,N_744,N_794);
and U1192 (N_1192,N_633,N_587);
nor U1193 (N_1193,N_596,N_503);
nor U1194 (N_1194,N_769,N_737);
and U1195 (N_1195,N_622,N_638);
xnor U1196 (N_1196,N_760,N_524);
nand U1197 (N_1197,N_516,N_786);
nand U1198 (N_1198,N_895,N_569);
xor U1199 (N_1199,N_669,N_749);
nand U1200 (N_1200,N_900,N_586);
xnor U1201 (N_1201,N_665,N_847);
xnor U1202 (N_1202,N_849,N_672);
or U1203 (N_1203,N_555,N_816);
xnor U1204 (N_1204,N_566,N_850);
nor U1205 (N_1205,N_758,N_642);
nor U1206 (N_1206,N_984,N_814);
nor U1207 (N_1207,N_702,N_660);
nand U1208 (N_1208,N_848,N_723);
or U1209 (N_1209,N_955,N_724);
and U1210 (N_1210,N_558,N_709);
nor U1211 (N_1211,N_547,N_784);
or U1212 (N_1212,N_695,N_817);
xor U1213 (N_1213,N_748,N_647);
xnor U1214 (N_1214,N_905,N_845);
and U1215 (N_1215,N_582,N_625);
or U1216 (N_1216,N_790,N_573);
or U1217 (N_1217,N_938,N_854);
xor U1218 (N_1218,N_909,N_658);
nand U1219 (N_1219,N_772,N_578);
nor U1220 (N_1220,N_580,N_902);
and U1221 (N_1221,N_993,N_671);
nand U1222 (N_1222,N_631,N_857);
or U1223 (N_1223,N_778,N_985);
nand U1224 (N_1224,N_935,N_697);
xnor U1225 (N_1225,N_664,N_714);
nand U1226 (N_1226,N_920,N_655);
xnor U1227 (N_1227,N_916,N_703);
xor U1228 (N_1228,N_528,N_733);
xor U1229 (N_1229,N_718,N_838);
nor U1230 (N_1230,N_597,N_663);
and U1231 (N_1231,N_743,N_722);
and U1232 (N_1232,N_536,N_546);
xnor U1233 (N_1233,N_970,N_646);
xnor U1234 (N_1234,N_901,N_675);
and U1235 (N_1235,N_830,N_526);
nor U1236 (N_1236,N_559,N_780);
nor U1237 (N_1237,N_876,N_673);
or U1238 (N_1238,N_509,N_593);
xnor U1239 (N_1239,N_674,N_741);
nand U1240 (N_1240,N_919,N_506);
and U1241 (N_1241,N_872,N_505);
or U1242 (N_1242,N_754,N_515);
or U1243 (N_1243,N_899,N_751);
nand U1244 (N_1244,N_988,N_589);
nand U1245 (N_1245,N_711,N_591);
nand U1246 (N_1246,N_706,N_958);
and U1247 (N_1247,N_927,N_908);
and U1248 (N_1248,N_621,N_906);
and U1249 (N_1249,N_844,N_924);
or U1250 (N_1250,N_964,N_999);
and U1251 (N_1251,N_698,N_703);
nor U1252 (N_1252,N_762,N_685);
nand U1253 (N_1253,N_769,N_575);
or U1254 (N_1254,N_886,N_580);
nor U1255 (N_1255,N_554,N_695);
nor U1256 (N_1256,N_774,N_709);
and U1257 (N_1257,N_988,N_856);
or U1258 (N_1258,N_945,N_653);
and U1259 (N_1259,N_653,N_929);
and U1260 (N_1260,N_833,N_614);
xnor U1261 (N_1261,N_806,N_871);
nand U1262 (N_1262,N_801,N_710);
xor U1263 (N_1263,N_514,N_560);
nand U1264 (N_1264,N_957,N_702);
or U1265 (N_1265,N_631,N_861);
and U1266 (N_1266,N_822,N_775);
or U1267 (N_1267,N_674,N_953);
and U1268 (N_1268,N_907,N_616);
nand U1269 (N_1269,N_765,N_655);
nand U1270 (N_1270,N_547,N_601);
nor U1271 (N_1271,N_890,N_906);
xor U1272 (N_1272,N_991,N_794);
nand U1273 (N_1273,N_615,N_791);
or U1274 (N_1274,N_678,N_548);
nand U1275 (N_1275,N_825,N_758);
and U1276 (N_1276,N_629,N_780);
and U1277 (N_1277,N_679,N_710);
and U1278 (N_1278,N_638,N_962);
or U1279 (N_1279,N_907,N_644);
xor U1280 (N_1280,N_807,N_880);
nand U1281 (N_1281,N_524,N_649);
nand U1282 (N_1282,N_736,N_905);
xnor U1283 (N_1283,N_634,N_816);
nor U1284 (N_1284,N_667,N_987);
nor U1285 (N_1285,N_784,N_690);
nand U1286 (N_1286,N_786,N_728);
and U1287 (N_1287,N_559,N_829);
nand U1288 (N_1288,N_516,N_743);
or U1289 (N_1289,N_576,N_787);
or U1290 (N_1290,N_675,N_580);
xnor U1291 (N_1291,N_621,N_767);
or U1292 (N_1292,N_991,N_700);
and U1293 (N_1293,N_899,N_971);
and U1294 (N_1294,N_801,N_993);
nand U1295 (N_1295,N_709,N_501);
nor U1296 (N_1296,N_798,N_842);
and U1297 (N_1297,N_770,N_974);
or U1298 (N_1298,N_828,N_778);
and U1299 (N_1299,N_701,N_708);
nand U1300 (N_1300,N_795,N_974);
nand U1301 (N_1301,N_917,N_987);
and U1302 (N_1302,N_668,N_827);
nand U1303 (N_1303,N_667,N_836);
or U1304 (N_1304,N_559,N_963);
nand U1305 (N_1305,N_818,N_792);
xor U1306 (N_1306,N_640,N_636);
nand U1307 (N_1307,N_576,N_720);
nand U1308 (N_1308,N_819,N_871);
and U1309 (N_1309,N_903,N_704);
nand U1310 (N_1310,N_967,N_968);
or U1311 (N_1311,N_787,N_571);
nor U1312 (N_1312,N_685,N_785);
xor U1313 (N_1313,N_555,N_982);
nand U1314 (N_1314,N_769,N_586);
nand U1315 (N_1315,N_646,N_776);
xor U1316 (N_1316,N_595,N_644);
xor U1317 (N_1317,N_875,N_511);
nand U1318 (N_1318,N_511,N_967);
or U1319 (N_1319,N_958,N_880);
or U1320 (N_1320,N_925,N_863);
nor U1321 (N_1321,N_786,N_671);
or U1322 (N_1322,N_577,N_810);
nor U1323 (N_1323,N_514,N_571);
or U1324 (N_1324,N_881,N_829);
nor U1325 (N_1325,N_993,N_618);
nand U1326 (N_1326,N_857,N_625);
and U1327 (N_1327,N_738,N_659);
and U1328 (N_1328,N_512,N_597);
and U1329 (N_1329,N_717,N_877);
nand U1330 (N_1330,N_915,N_828);
xnor U1331 (N_1331,N_975,N_750);
and U1332 (N_1332,N_952,N_507);
or U1333 (N_1333,N_702,N_788);
xnor U1334 (N_1334,N_727,N_935);
nand U1335 (N_1335,N_841,N_760);
xor U1336 (N_1336,N_850,N_842);
xnor U1337 (N_1337,N_553,N_967);
and U1338 (N_1338,N_793,N_580);
and U1339 (N_1339,N_699,N_691);
xor U1340 (N_1340,N_876,N_816);
or U1341 (N_1341,N_687,N_745);
or U1342 (N_1342,N_867,N_890);
and U1343 (N_1343,N_893,N_525);
and U1344 (N_1344,N_635,N_540);
xor U1345 (N_1345,N_948,N_607);
nand U1346 (N_1346,N_896,N_909);
nand U1347 (N_1347,N_805,N_531);
nand U1348 (N_1348,N_791,N_650);
nor U1349 (N_1349,N_648,N_701);
nor U1350 (N_1350,N_589,N_844);
nand U1351 (N_1351,N_918,N_738);
nand U1352 (N_1352,N_950,N_799);
nand U1353 (N_1353,N_547,N_855);
or U1354 (N_1354,N_891,N_671);
nor U1355 (N_1355,N_586,N_710);
or U1356 (N_1356,N_995,N_761);
nor U1357 (N_1357,N_862,N_676);
and U1358 (N_1358,N_559,N_816);
or U1359 (N_1359,N_923,N_747);
or U1360 (N_1360,N_658,N_601);
nor U1361 (N_1361,N_600,N_972);
nand U1362 (N_1362,N_714,N_644);
nand U1363 (N_1363,N_558,N_957);
or U1364 (N_1364,N_584,N_668);
nand U1365 (N_1365,N_637,N_942);
xnor U1366 (N_1366,N_641,N_606);
or U1367 (N_1367,N_577,N_966);
and U1368 (N_1368,N_764,N_645);
nand U1369 (N_1369,N_987,N_629);
nand U1370 (N_1370,N_641,N_996);
or U1371 (N_1371,N_672,N_556);
nor U1372 (N_1372,N_588,N_502);
or U1373 (N_1373,N_763,N_915);
nor U1374 (N_1374,N_939,N_517);
xnor U1375 (N_1375,N_773,N_873);
or U1376 (N_1376,N_704,N_816);
and U1377 (N_1377,N_831,N_560);
or U1378 (N_1378,N_799,N_526);
nand U1379 (N_1379,N_578,N_905);
nor U1380 (N_1380,N_515,N_659);
and U1381 (N_1381,N_840,N_543);
xnor U1382 (N_1382,N_809,N_572);
xor U1383 (N_1383,N_706,N_933);
nand U1384 (N_1384,N_940,N_917);
or U1385 (N_1385,N_845,N_520);
nor U1386 (N_1386,N_904,N_524);
and U1387 (N_1387,N_708,N_889);
xnor U1388 (N_1388,N_724,N_538);
xor U1389 (N_1389,N_640,N_709);
and U1390 (N_1390,N_966,N_700);
and U1391 (N_1391,N_718,N_927);
nand U1392 (N_1392,N_782,N_586);
xor U1393 (N_1393,N_987,N_827);
nand U1394 (N_1394,N_624,N_721);
or U1395 (N_1395,N_529,N_703);
xnor U1396 (N_1396,N_728,N_986);
nand U1397 (N_1397,N_948,N_767);
nor U1398 (N_1398,N_525,N_995);
nor U1399 (N_1399,N_646,N_973);
and U1400 (N_1400,N_552,N_993);
or U1401 (N_1401,N_858,N_658);
nand U1402 (N_1402,N_833,N_851);
and U1403 (N_1403,N_521,N_918);
or U1404 (N_1404,N_627,N_892);
xnor U1405 (N_1405,N_906,N_816);
xnor U1406 (N_1406,N_501,N_748);
xnor U1407 (N_1407,N_529,N_501);
nand U1408 (N_1408,N_775,N_620);
xor U1409 (N_1409,N_672,N_948);
or U1410 (N_1410,N_777,N_614);
nor U1411 (N_1411,N_806,N_980);
nand U1412 (N_1412,N_972,N_662);
nand U1413 (N_1413,N_500,N_952);
xor U1414 (N_1414,N_991,N_529);
nand U1415 (N_1415,N_918,N_901);
or U1416 (N_1416,N_699,N_957);
or U1417 (N_1417,N_749,N_621);
nand U1418 (N_1418,N_792,N_730);
or U1419 (N_1419,N_688,N_667);
or U1420 (N_1420,N_731,N_817);
or U1421 (N_1421,N_918,N_538);
xor U1422 (N_1422,N_853,N_745);
xnor U1423 (N_1423,N_641,N_504);
nand U1424 (N_1424,N_883,N_837);
or U1425 (N_1425,N_936,N_514);
xor U1426 (N_1426,N_942,N_872);
and U1427 (N_1427,N_865,N_578);
or U1428 (N_1428,N_714,N_619);
nor U1429 (N_1429,N_675,N_862);
and U1430 (N_1430,N_625,N_649);
nand U1431 (N_1431,N_734,N_849);
or U1432 (N_1432,N_990,N_777);
and U1433 (N_1433,N_531,N_543);
nand U1434 (N_1434,N_719,N_793);
and U1435 (N_1435,N_873,N_916);
or U1436 (N_1436,N_767,N_551);
and U1437 (N_1437,N_561,N_982);
or U1438 (N_1438,N_777,N_516);
or U1439 (N_1439,N_505,N_735);
xor U1440 (N_1440,N_543,N_665);
nor U1441 (N_1441,N_903,N_658);
or U1442 (N_1442,N_698,N_932);
or U1443 (N_1443,N_922,N_711);
or U1444 (N_1444,N_608,N_943);
xor U1445 (N_1445,N_956,N_686);
nand U1446 (N_1446,N_796,N_993);
nand U1447 (N_1447,N_568,N_614);
nand U1448 (N_1448,N_550,N_687);
or U1449 (N_1449,N_916,N_721);
or U1450 (N_1450,N_791,N_613);
or U1451 (N_1451,N_759,N_886);
or U1452 (N_1452,N_594,N_617);
xnor U1453 (N_1453,N_554,N_576);
or U1454 (N_1454,N_768,N_561);
nand U1455 (N_1455,N_551,N_953);
or U1456 (N_1456,N_637,N_587);
nor U1457 (N_1457,N_976,N_520);
or U1458 (N_1458,N_852,N_935);
nand U1459 (N_1459,N_769,N_563);
or U1460 (N_1460,N_804,N_670);
nor U1461 (N_1461,N_603,N_898);
or U1462 (N_1462,N_777,N_570);
nand U1463 (N_1463,N_994,N_734);
nand U1464 (N_1464,N_967,N_775);
or U1465 (N_1465,N_762,N_892);
nor U1466 (N_1466,N_586,N_628);
or U1467 (N_1467,N_525,N_991);
nor U1468 (N_1468,N_992,N_555);
nand U1469 (N_1469,N_720,N_757);
nor U1470 (N_1470,N_608,N_877);
or U1471 (N_1471,N_609,N_882);
and U1472 (N_1472,N_894,N_827);
nand U1473 (N_1473,N_712,N_709);
and U1474 (N_1474,N_840,N_652);
nand U1475 (N_1475,N_509,N_654);
xnor U1476 (N_1476,N_543,N_973);
or U1477 (N_1477,N_880,N_684);
nor U1478 (N_1478,N_688,N_781);
nor U1479 (N_1479,N_554,N_705);
and U1480 (N_1480,N_646,N_816);
xnor U1481 (N_1481,N_629,N_658);
nand U1482 (N_1482,N_699,N_570);
and U1483 (N_1483,N_691,N_776);
nor U1484 (N_1484,N_762,N_933);
and U1485 (N_1485,N_925,N_761);
nor U1486 (N_1486,N_729,N_662);
and U1487 (N_1487,N_858,N_635);
or U1488 (N_1488,N_570,N_979);
nor U1489 (N_1489,N_907,N_525);
nor U1490 (N_1490,N_922,N_916);
nand U1491 (N_1491,N_911,N_608);
xor U1492 (N_1492,N_800,N_702);
or U1493 (N_1493,N_881,N_717);
xor U1494 (N_1494,N_741,N_582);
nor U1495 (N_1495,N_678,N_881);
and U1496 (N_1496,N_946,N_580);
nor U1497 (N_1497,N_752,N_909);
nor U1498 (N_1498,N_933,N_797);
and U1499 (N_1499,N_809,N_942);
xnor U1500 (N_1500,N_1138,N_1301);
or U1501 (N_1501,N_1213,N_1099);
or U1502 (N_1502,N_1416,N_1445);
and U1503 (N_1503,N_1177,N_1371);
nor U1504 (N_1504,N_1407,N_1386);
xnor U1505 (N_1505,N_1450,N_1186);
and U1506 (N_1506,N_1264,N_1352);
xor U1507 (N_1507,N_1114,N_1305);
and U1508 (N_1508,N_1346,N_1269);
and U1509 (N_1509,N_1265,N_1102);
nand U1510 (N_1510,N_1408,N_1061);
nand U1511 (N_1511,N_1317,N_1419);
nor U1512 (N_1512,N_1032,N_1350);
or U1513 (N_1513,N_1146,N_1312);
nand U1514 (N_1514,N_1329,N_1081);
and U1515 (N_1515,N_1476,N_1261);
or U1516 (N_1516,N_1428,N_1420);
or U1517 (N_1517,N_1007,N_1343);
and U1518 (N_1518,N_1166,N_1117);
and U1519 (N_1519,N_1396,N_1197);
nand U1520 (N_1520,N_1479,N_1040);
or U1521 (N_1521,N_1018,N_1489);
and U1522 (N_1522,N_1154,N_1108);
nand U1523 (N_1523,N_1015,N_1124);
or U1524 (N_1524,N_1313,N_1341);
or U1525 (N_1525,N_1185,N_1452);
or U1526 (N_1526,N_1252,N_1315);
and U1527 (N_1527,N_1057,N_1482);
or U1528 (N_1528,N_1337,N_1283);
xor U1529 (N_1529,N_1339,N_1063);
and U1530 (N_1530,N_1226,N_1424);
or U1531 (N_1531,N_1498,N_1430);
and U1532 (N_1532,N_1228,N_1409);
or U1533 (N_1533,N_1161,N_1029);
or U1534 (N_1534,N_1323,N_1326);
xnor U1535 (N_1535,N_1413,N_1249);
nand U1536 (N_1536,N_1179,N_1297);
nand U1537 (N_1537,N_1493,N_1441);
nand U1538 (N_1538,N_1333,N_1172);
nor U1539 (N_1539,N_1463,N_1244);
or U1540 (N_1540,N_1336,N_1480);
xor U1541 (N_1541,N_1483,N_1318);
and U1542 (N_1542,N_1028,N_1242);
and U1543 (N_1543,N_1142,N_1306);
xor U1544 (N_1544,N_1435,N_1487);
nor U1545 (N_1545,N_1077,N_1250);
nor U1546 (N_1546,N_1291,N_1023);
nand U1547 (N_1547,N_1144,N_1072);
nand U1548 (N_1548,N_1403,N_1240);
nand U1549 (N_1549,N_1017,N_1270);
and U1550 (N_1550,N_1314,N_1257);
or U1551 (N_1551,N_1207,N_1140);
or U1552 (N_1552,N_1034,N_1293);
xnor U1553 (N_1553,N_1405,N_1376);
and U1554 (N_1554,N_1472,N_1495);
xor U1555 (N_1555,N_1021,N_1120);
nor U1556 (N_1556,N_1211,N_1043);
or U1557 (N_1557,N_1436,N_1049);
xor U1558 (N_1558,N_1074,N_1204);
nor U1559 (N_1559,N_1488,N_1135);
xnor U1560 (N_1560,N_1158,N_1360);
nor U1561 (N_1561,N_1279,N_1263);
or U1562 (N_1562,N_1009,N_1221);
or U1563 (N_1563,N_1434,N_1176);
and U1564 (N_1564,N_1110,N_1109);
and U1565 (N_1565,N_1200,N_1453);
xnor U1566 (N_1566,N_1107,N_1098);
nor U1567 (N_1567,N_1397,N_1066);
nand U1568 (N_1568,N_1225,N_1069);
or U1569 (N_1569,N_1369,N_1275);
xor U1570 (N_1570,N_1481,N_1392);
nor U1571 (N_1571,N_1295,N_1382);
nand U1572 (N_1572,N_1347,N_1444);
xnor U1573 (N_1573,N_1359,N_1274);
nand U1574 (N_1574,N_1000,N_1169);
nand U1575 (N_1575,N_1327,N_1237);
xnor U1576 (N_1576,N_1067,N_1082);
or U1577 (N_1577,N_1367,N_1319);
nor U1578 (N_1578,N_1272,N_1459);
xor U1579 (N_1579,N_1147,N_1006);
and U1580 (N_1580,N_1073,N_1348);
xor U1581 (N_1581,N_1189,N_1393);
xor U1582 (N_1582,N_1182,N_1448);
nor U1583 (N_1583,N_1202,N_1457);
and U1584 (N_1584,N_1255,N_1206);
nor U1585 (N_1585,N_1302,N_1433);
and U1586 (N_1586,N_1203,N_1119);
nor U1587 (N_1587,N_1080,N_1148);
nand U1588 (N_1588,N_1273,N_1451);
or U1589 (N_1589,N_1022,N_1462);
nor U1590 (N_1590,N_1159,N_1229);
and U1591 (N_1591,N_1310,N_1331);
nor U1592 (N_1592,N_1192,N_1175);
nand U1593 (N_1593,N_1247,N_1042);
or U1594 (N_1594,N_1011,N_1193);
xnor U1595 (N_1595,N_1231,N_1103);
nand U1596 (N_1596,N_1027,N_1150);
xor U1597 (N_1597,N_1054,N_1385);
xnor U1598 (N_1598,N_1092,N_1288);
and U1599 (N_1599,N_1012,N_1342);
xor U1600 (N_1600,N_1025,N_1289);
nor U1601 (N_1601,N_1366,N_1473);
or U1602 (N_1602,N_1093,N_1438);
and U1603 (N_1603,N_1139,N_1155);
or U1604 (N_1604,N_1128,N_1113);
nand U1605 (N_1605,N_1276,N_1222);
nand U1606 (N_1606,N_1432,N_1187);
and U1607 (N_1607,N_1490,N_1129);
xnor U1608 (N_1608,N_1469,N_1351);
and U1609 (N_1609,N_1078,N_1245);
xnor U1610 (N_1610,N_1446,N_1227);
nand U1611 (N_1611,N_1091,N_1149);
or U1612 (N_1612,N_1036,N_1431);
and U1613 (N_1613,N_1165,N_1060);
and U1614 (N_1614,N_1168,N_1131);
nor U1615 (N_1615,N_1344,N_1132);
nor U1616 (N_1616,N_1358,N_1191);
or U1617 (N_1617,N_1353,N_1497);
nand U1618 (N_1618,N_1217,N_1425);
and U1619 (N_1619,N_1335,N_1118);
and U1620 (N_1620,N_1001,N_1477);
or U1621 (N_1621,N_1111,N_1033);
and U1622 (N_1622,N_1308,N_1485);
xor U1623 (N_1623,N_1259,N_1447);
or U1624 (N_1624,N_1404,N_1039);
nand U1625 (N_1625,N_1389,N_1475);
nand U1626 (N_1626,N_1285,N_1127);
and U1627 (N_1627,N_1031,N_1373);
nor U1628 (N_1628,N_1121,N_1160);
nor U1629 (N_1629,N_1090,N_1105);
nor U1630 (N_1630,N_1375,N_1426);
or U1631 (N_1631,N_1461,N_1126);
and U1632 (N_1632,N_1325,N_1048);
xnor U1633 (N_1633,N_1079,N_1084);
xor U1634 (N_1634,N_1095,N_1300);
and U1635 (N_1635,N_1356,N_1152);
nand U1636 (N_1636,N_1307,N_1429);
xor U1637 (N_1637,N_1051,N_1232);
xor U1638 (N_1638,N_1384,N_1330);
and U1639 (N_1639,N_1097,N_1387);
or U1640 (N_1640,N_1471,N_1423);
nand U1641 (N_1641,N_1381,N_1468);
xor U1642 (N_1642,N_1088,N_1047);
or U1643 (N_1643,N_1454,N_1209);
xor U1644 (N_1644,N_1220,N_1440);
nand U1645 (N_1645,N_1253,N_1374);
nand U1646 (N_1646,N_1096,N_1201);
or U1647 (N_1647,N_1418,N_1156);
nand U1648 (N_1648,N_1294,N_1398);
xnor U1649 (N_1649,N_1071,N_1205);
and U1650 (N_1650,N_1492,N_1068);
nor U1651 (N_1651,N_1284,N_1062);
or U1652 (N_1652,N_1467,N_1458);
xnor U1653 (N_1653,N_1134,N_1016);
xor U1654 (N_1654,N_1199,N_1290);
nand U1655 (N_1655,N_1410,N_1280);
or U1656 (N_1656,N_1194,N_1399);
nor U1657 (N_1657,N_1085,N_1266);
or U1658 (N_1658,N_1198,N_1024);
nand U1659 (N_1659,N_1173,N_1181);
or U1660 (N_1660,N_1286,N_1046);
nand U1661 (N_1661,N_1122,N_1484);
nand U1662 (N_1662,N_1070,N_1125);
and U1663 (N_1663,N_1422,N_1298);
and U1664 (N_1664,N_1013,N_1143);
xor U1665 (N_1665,N_1215,N_1162);
xnor U1666 (N_1666,N_1170,N_1234);
and U1667 (N_1667,N_1157,N_1010);
or U1668 (N_1668,N_1238,N_1402);
nand U1669 (N_1669,N_1180,N_1401);
and U1670 (N_1670,N_1052,N_1491);
and U1671 (N_1671,N_1241,N_1395);
nand U1672 (N_1672,N_1421,N_1328);
xor U1673 (N_1673,N_1045,N_1026);
or U1674 (N_1674,N_1439,N_1456);
xnor U1675 (N_1675,N_1390,N_1377);
xor U1676 (N_1676,N_1355,N_1038);
nor U1677 (N_1677,N_1246,N_1044);
nor U1678 (N_1678,N_1388,N_1478);
nand U1679 (N_1679,N_1267,N_1400);
nor U1680 (N_1680,N_1208,N_1239);
nand U1681 (N_1681,N_1230,N_1311);
xnor U1682 (N_1682,N_1171,N_1271);
nand U1683 (N_1683,N_1104,N_1055);
nand U1684 (N_1684,N_1100,N_1304);
or U1685 (N_1685,N_1368,N_1087);
nor U1686 (N_1686,N_1299,N_1281);
nor U1687 (N_1687,N_1136,N_1406);
and U1688 (N_1688,N_1106,N_1212);
nor U1689 (N_1689,N_1035,N_1145);
or U1690 (N_1690,N_1365,N_1195);
or U1691 (N_1691,N_1362,N_1449);
and U1692 (N_1692,N_1364,N_1260);
nand U1693 (N_1693,N_1464,N_1417);
or U1694 (N_1694,N_1496,N_1332);
nor U1695 (N_1695,N_1460,N_1218);
or U1696 (N_1696,N_1075,N_1470);
nor U1697 (N_1697,N_1334,N_1494);
nand U1698 (N_1698,N_1278,N_1003);
nand U1699 (N_1699,N_1383,N_1123);
and U1700 (N_1700,N_1465,N_1014);
nor U1701 (N_1701,N_1214,N_1316);
nor U1702 (N_1702,N_1020,N_1303);
nor U1703 (N_1703,N_1361,N_1277);
and U1704 (N_1704,N_1268,N_1041);
nor U1705 (N_1705,N_1223,N_1196);
xnor U1706 (N_1706,N_1059,N_1499);
xnor U1707 (N_1707,N_1378,N_1065);
or U1708 (N_1708,N_1235,N_1379);
xor U1709 (N_1709,N_1455,N_1474);
nor U1710 (N_1710,N_1151,N_1320);
nand U1711 (N_1711,N_1322,N_1258);
or U1712 (N_1712,N_1053,N_1050);
xor U1713 (N_1713,N_1058,N_1019);
nor U1714 (N_1714,N_1101,N_1427);
or U1715 (N_1715,N_1183,N_1345);
or U1716 (N_1716,N_1370,N_1137);
xnor U1717 (N_1717,N_1357,N_1094);
nand U1718 (N_1718,N_1236,N_1251);
or U1719 (N_1719,N_1321,N_1248);
nor U1720 (N_1720,N_1210,N_1153);
and U1721 (N_1721,N_1442,N_1292);
and U1722 (N_1722,N_1415,N_1443);
or U1723 (N_1723,N_1338,N_1008);
nand U1724 (N_1724,N_1064,N_1394);
nand U1725 (N_1725,N_1086,N_1219);
nor U1726 (N_1726,N_1167,N_1133);
nand U1727 (N_1727,N_1340,N_1349);
and U1728 (N_1728,N_1412,N_1004);
or U1729 (N_1729,N_1324,N_1233);
nor U1730 (N_1730,N_1116,N_1002);
and U1731 (N_1731,N_1282,N_1163);
and U1732 (N_1732,N_1112,N_1190);
nor U1733 (N_1733,N_1287,N_1262);
xnor U1734 (N_1734,N_1466,N_1254);
and U1735 (N_1735,N_1411,N_1380);
xnor U1736 (N_1736,N_1141,N_1486);
or U1737 (N_1737,N_1089,N_1224);
or U1738 (N_1738,N_1164,N_1243);
nand U1739 (N_1739,N_1309,N_1391);
nor U1740 (N_1740,N_1184,N_1363);
nor U1741 (N_1741,N_1174,N_1056);
or U1742 (N_1742,N_1256,N_1372);
xor U1743 (N_1743,N_1037,N_1296);
xor U1744 (N_1744,N_1076,N_1216);
nand U1745 (N_1745,N_1437,N_1354);
and U1746 (N_1746,N_1115,N_1178);
xnor U1747 (N_1747,N_1188,N_1414);
nand U1748 (N_1748,N_1030,N_1005);
or U1749 (N_1749,N_1130,N_1083);
xnor U1750 (N_1750,N_1012,N_1392);
nor U1751 (N_1751,N_1011,N_1182);
and U1752 (N_1752,N_1097,N_1244);
and U1753 (N_1753,N_1150,N_1113);
or U1754 (N_1754,N_1288,N_1165);
or U1755 (N_1755,N_1334,N_1397);
xor U1756 (N_1756,N_1320,N_1093);
and U1757 (N_1757,N_1066,N_1454);
xor U1758 (N_1758,N_1123,N_1069);
and U1759 (N_1759,N_1301,N_1353);
xor U1760 (N_1760,N_1242,N_1284);
nor U1761 (N_1761,N_1026,N_1194);
or U1762 (N_1762,N_1300,N_1441);
nand U1763 (N_1763,N_1084,N_1243);
xnor U1764 (N_1764,N_1014,N_1123);
and U1765 (N_1765,N_1257,N_1224);
or U1766 (N_1766,N_1426,N_1005);
and U1767 (N_1767,N_1439,N_1301);
xnor U1768 (N_1768,N_1032,N_1436);
nor U1769 (N_1769,N_1233,N_1114);
nand U1770 (N_1770,N_1405,N_1114);
xnor U1771 (N_1771,N_1278,N_1292);
or U1772 (N_1772,N_1359,N_1388);
or U1773 (N_1773,N_1214,N_1213);
xnor U1774 (N_1774,N_1245,N_1289);
xor U1775 (N_1775,N_1113,N_1337);
nor U1776 (N_1776,N_1263,N_1478);
xnor U1777 (N_1777,N_1330,N_1446);
and U1778 (N_1778,N_1227,N_1374);
or U1779 (N_1779,N_1022,N_1426);
xnor U1780 (N_1780,N_1113,N_1222);
nor U1781 (N_1781,N_1460,N_1356);
and U1782 (N_1782,N_1233,N_1190);
nand U1783 (N_1783,N_1305,N_1470);
and U1784 (N_1784,N_1007,N_1287);
xor U1785 (N_1785,N_1355,N_1397);
nor U1786 (N_1786,N_1120,N_1171);
nor U1787 (N_1787,N_1157,N_1041);
nand U1788 (N_1788,N_1452,N_1489);
nand U1789 (N_1789,N_1365,N_1381);
nand U1790 (N_1790,N_1357,N_1365);
or U1791 (N_1791,N_1090,N_1311);
nand U1792 (N_1792,N_1128,N_1323);
and U1793 (N_1793,N_1090,N_1205);
nor U1794 (N_1794,N_1350,N_1270);
xnor U1795 (N_1795,N_1094,N_1216);
nand U1796 (N_1796,N_1408,N_1343);
nand U1797 (N_1797,N_1002,N_1033);
xor U1798 (N_1798,N_1437,N_1372);
nor U1799 (N_1799,N_1050,N_1237);
and U1800 (N_1800,N_1187,N_1264);
and U1801 (N_1801,N_1302,N_1371);
xor U1802 (N_1802,N_1379,N_1483);
xor U1803 (N_1803,N_1355,N_1069);
or U1804 (N_1804,N_1455,N_1108);
or U1805 (N_1805,N_1212,N_1222);
xor U1806 (N_1806,N_1436,N_1304);
and U1807 (N_1807,N_1054,N_1464);
nand U1808 (N_1808,N_1053,N_1373);
xor U1809 (N_1809,N_1316,N_1075);
nand U1810 (N_1810,N_1080,N_1179);
nor U1811 (N_1811,N_1451,N_1218);
or U1812 (N_1812,N_1375,N_1205);
nand U1813 (N_1813,N_1068,N_1224);
and U1814 (N_1814,N_1101,N_1144);
xor U1815 (N_1815,N_1018,N_1325);
and U1816 (N_1816,N_1495,N_1277);
or U1817 (N_1817,N_1215,N_1430);
xnor U1818 (N_1818,N_1146,N_1007);
xor U1819 (N_1819,N_1249,N_1340);
and U1820 (N_1820,N_1291,N_1295);
or U1821 (N_1821,N_1017,N_1055);
xor U1822 (N_1822,N_1119,N_1340);
and U1823 (N_1823,N_1405,N_1340);
and U1824 (N_1824,N_1079,N_1377);
and U1825 (N_1825,N_1290,N_1166);
and U1826 (N_1826,N_1464,N_1072);
xor U1827 (N_1827,N_1461,N_1351);
nand U1828 (N_1828,N_1154,N_1063);
or U1829 (N_1829,N_1131,N_1099);
nor U1830 (N_1830,N_1210,N_1368);
nand U1831 (N_1831,N_1487,N_1348);
xnor U1832 (N_1832,N_1253,N_1142);
or U1833 (N_1833,N_1298,N_1473);
xnor U1834 (N_1834,N_1068,N_1375);
nand U1835 (N_1835,N_1319,N_1088);
nor U1836 (N_1836,N_1045,N_1070);
nor U1837 (N_1837,N_1259,N_1218);
xnor U1838 (N_1838,N_1497,N_1039);
xnor U1839 (N_1839,N_1490,N_1213);
nor U1840 (N_1840,N_1010,N_1340);
nor U1841 (N_1841,N_1023,N_1087);
and U1842 (N_1842,N_1135,N_1221);
nor U1843 (N_1843,N_1082,N_1487);
or U1844 (N_1844,N_1396,N_1109);
or U1845 (N_1845,N_1477,N_1016);
xnor U1846 (N_1846,N_1103,N_1497);
or U1847 (N_1847,N_1178,N_1097);
or U1848 (N_1848,N_1464,N_1237);
nand U1849 (N_1849,N_1439,N_1223);
xor U1850 (N_1850,N_1387,N_1015);
nor U1851 (N_1851,N_1424,N_1143);
nand U1852 (N_1852,N_1198,N_1014);
nand U1853 (N_1853,N_1304,N_1427);
nand U1854 (N_1854,N_1099,N_1408);
xor U1855 (N_1855,N_1000,N_1200);
or U1856 (N_1856,N_1282,N_1240);
xor U1857 (N_1857,N_1410,N_1055);
or U1858 (N_1858,N_1375,N_1266);
or U1859 (N_1859,N_1055,N_1352);
nor U1860 (N_1860,N_1293,N_1006);
or U1861 (N_1861,N_1097,N_1237);
and U1862 (N_1862,N_1353,N_1378);
nand U1863 (N_1863,N_1451,N_1133);
xor U1864 (N_1864,N_1252,N_1001);
and U1865 (N_1865,N_1046,N_1077);
nand U1866 (N_1866,N_1171,N_1110);
and U1867 (N_1867,N_1155,N_1142);
or U1868 (N_1868,N_1005,N_1327);
xor U1869 (N_1869,N_1038,N_1013);
and U1870 (N_1870,N_1433,N_1266);
nor U1871 (N_1871,N_1136,N_1218);
nor U1872 (N_1872,N_1458,N_1378);
or U1873 (N_1873,N_1129,N_1244);
xnor U1874 (N_1874,N_1319,N_1447);
or U1875 (N_1875,N_1377,N_1225);
or U1876 (N_1876,N_1225,N_1419);
nand U1877 (N_1877,N_1321,N_1314);
and U1878 (N_1878,N_1092,N_1027);
and U1879 (N_1879,N_1154,N_1109);
nand U1880 (N_1880,N_1193,N_1134);
and U1881 (N_1881,N_1247,N_1305);
nand U1882 (N_1882,N_1445,N_1325);
nand U1883 (N_1883,N_1189,N_1458);
nand U1884 (N_1884,N_1482,N_1176);
xnor U1885 (N_1885,N_1308,N_1459);
or U1886 (N_1886,N_1127,N_1278);
and U1887 (N_1887,N_1269,N_1257);
or U1888 (N_1888,N_1370,N_1028);
nand U1889 (N_1889,N_1040,N_1376);
and U1890 (N_1890,N_1464,N_1225);
and U1891 (N_1891,N_1355,N_1099);
or U1892 (N_1892,N_1163,N_1460);
or U1893 (N_1893,N_1246,N_1450);
nand U1894 (N_1894,N_1466,N_1337);
nand U1895 (N_1895,N_1092,N_1023);
nand U1896 (N_1896,N_1494,N_1387);
or U1897 (N_1897,N_1035,N_1302);
nand U1898 (N_1898,N_1299,N_1108);
or U1899 (N_1899,N_1009,N_1334);
nor U1900 (N_1900,N_1064,N_1043);
and U1901 (N_1901,N_1241,N_1100);
or U1902 (N_1902,N_1256,N_1007);
xnor U1903 (N_1903,N_1168,N_1488);
or U1904 (N_1904,N_1343,N_1477);
xor U1905 (N_1905,N_1070,N_1242);
or U1906 (N_1906,N_1346,N_1226);
nand U1907 (N_1907,N_1176,N_1083);
or U1908 (N_1908,N_1213,N_1323);
nand U1909 (N_1909,N_1041,N_1171);
nor U1910 (N_1910,N_1404,N_1436);
nand U1911 (N_1911,N_1372,N_1106);
and U1912 (N_1912,N_1183,N_1313);
nand U1913 (N_1913,N_1310,N_1081);
xor U1914 (N_1914,N_1464,N_1211);
and U1915 (N_1915,N_1033,N_1109);
and U1916 (N_1916,N_1451,N_1232);
nand U1917 (N_1917,N_1256,N_1021);
xnor U1918 (N_1918,N_1068,N_1437);
nor U1919 (N_1919,N_1055,N_1487);
xnor U1920 (N_1920,N_1316,N_1228);
nand U1921 (N_1921,N_1497,N_1318);
or U1922 (N_1922,N_1316,N_1162);
nor U1923 (N_1923,N_1465,N_1044);
xor U1924 (N_1924,N_1260,N_1473);
nand U1925 (N_1925,N_1457,N_1174);
or U1926 (N_1926,N_1321,N_1443);
xnor U1927 (N_1927,N_1118,N_1331);
xnor U1928 (N_1928,N_1382,N_1445);
or U1929 (N_1929,N_1386,N_1398);
or U1930 (N_1930,N_1286,N_1433);
nand U1931 (N_1931,N_1313,N_1196);
nor U1932 (N_1932,N_1125,N_1045);
or U1933 (N_1933,N_1133,N_1339);
or U1934 (N_1934,N_1226,N_1460);
nor U1935 (N_1935,N_1079,N_1276);
and U1936 (N_1936,N_1307,N_1041);
nand U1937 (N_1937,N_1468,N_1356);
nor U1938 (N_1938,N_1083,N_1235);
nor U1939 (N_1939,N_1084,N_1071);
xor U1940 (N_1940,N_1279,N_1446);
or U1941 (N_1941,N_1142,N_1230);
xor U1942 (N_1942,N_1166,N_1064);
nand U1943 (N_1943,N_1140,N_1360);
nor U1944 (N_1944,N_1385,N_1392);
and U1945 (N_1945,N_1026,N_1095);
nor U1946 (N_1946,N_1027,N_1091);
xnor U1947 (N_1947,N_1053,N_1041);
nor U1948 (N_1948,N_1469,N_1140);
or U1949 (N_1949,N_1425,N_1249);
or U1950 (N_1950,N_1451,N_1382);
xnor U1951 (N_1951,N_1388,N_1401);
and U1952 (N_1952,N_1370,N_1349);
and U1953 (N_1953,N_1185,N_1379);
and U1954 (N_1954,N_1222,N_1330);
nand U1955 (N_1955,N_1163,N_1311);
or U1956 (N_1956,N_1332,N_1066);
nand U1957 (N_1957,N_1209,N_1183);
or U1958 (N_1958,N_1259,N_1434);
nor U1959 (N_1959,N_1196,N_1127);
nor U1960 (N_1960,N_1038,N_1160);
and U1961 (N_1961,N_1393,N_1492);
nand U1962 (N_1962,N_1427,N_1136);
and U1963 (N_1963,N_1143,N_1132);
or U1964 (N_1964,N_1129,N_1059);
or U1965 (N_1965,N_1106,N_1062);
xor U1966 (N_1966,N_1404,N_1291);
nor U1967 (N_1967,N_1114,N_1109);
or U1968 (N_1968,N_1323,N_1398);
nor U1969 (N_1969,N_1157,N_1020);
xor U1970 (N_1970,N_1083,N_1257);
and U1971 (N_1971,N_1003,N_1253);
xor U1972 (N_1972,N_1368,N_1342);
nor U1973 (N_1973,N_1116,N_1195);
or U1974 (N_1974,N_1430,N_1128);
xor U1975 (N_1975,N_1048,N_1410);
nand U1976 (N_1976,N_1164,N_1387);
nand U1977 (N_1977,N_1261,N_1160);
or U1978 (N_1978,N_1495,N_1453);
nand U1979 (N_1979,N_1135,N_1243);
xnor U1980 (N_1980,N_1352,N_1026);
or U1981 (N_1981,N_1064,N_1267);
or U1982 (N_1982,N_1100,N_1077);
nand U1983 (N_1983,N_1448,N_1037);
xnor U1984 (N_1984,N_1426,N_1208);
or U1985 (N_1985,N_1334,N_1237);
nor U1986 (N_1986,N_1303,N_1354);
or U1987 (N_1987,N_1463,N_1253);
or U1988 (N_1988,N_1495,N_1172);
or U1989 (N_1989,N_1059,N_1494);
xnor U1990 (N_1990,N_1128,N_1172);
or U1991 (N_1991,N_1174,N_1182);
and U1992 (N_1992,N_1341,N_1249);
nor U1993 (N_1993,N_1163,N_1382);
nand U1994 (N_1994,N_1174,N_1102);
nor U1995 (N_1995,N_1452,N_1232);
xnor U1996 (N_1996,N_1244,N_1008);
nand U1997 (N_1997,N_1351,N_1263);
or U1998 (N_1998,N_1436,N_1132);
or U1999 (N_1999,N_1443,N_1241);
xor U2000 (N_2000,N_1699,N_1993);
and U2001 (N_2001,N_1503,N_1578);
nor U2002 (N_2002,N_1537,N_1531);
nor U2003 (N_2003,N_1764,N_1944);
or U2004 (N_2004,N_1637,N_1974);
nand U2005 (N_2005,N_1703,N_1852);
xor U2006 (N_2006,N_1639,N_1806);
nor U2007 (N_2007,N_1573,N_1522);
and U2008 (N_2008,N_1584,N_1773);
xor U2009 (N_2009,N_1548,N_1770);
nand U2010 (N_2010,N_1929,N_1595);
or U2011 (N_2011,N_1952,N_1611);
xnor U2012 (N_2012,N_1765,N_1543);
or U2013 (N_2013,N_1758,N_1742);
nand U2014 (N_2014,N_1879,N_1804);
nand U2015 (N_2015,N_1908,N_1851);
or U2016 (N_2016,N_1702,N_1886);
nand U2017 (N_2017,N_1977,N_1811);
or U2018 (N_2018,N_1867,N_1866);
nor U2019 (N_2019,N_1570,N_1817);
and U2020 (N_2020,N_1823,N_1677);
nor U2021 (N_2021,N_1981,N_1831);
nor U2022 (N_2022,N_1756,N_1655);
or U2023 (N_2023,N_1845,N_1784);
nor U2024 (N_2024,N_1885,N_1854);
xnor U2025 (N_2025,N_1840,N_1897);
and U2026 (N_2026,N_1988,N_1751);
and U2027 (N_2027,N_1515,N_1945);
xor U2028 (N_2028,N_1839,N_1906);
nor U2029 (N_2029,N_1964,N_1871);
nand U2030 (N_2030,N_1524,N_1794);
nand U2031 (N_2031,N_1819,N_1646);
xnor U2032 (N_2032,N_1684,N_1902);
and U2033 (N_2033,N_1690,N_1842);
nor U2034 (N_2034,N_1701,N_1553);
xor U2035 (N_2035,N_1685,N_1846);
nand U2036 (N_2036,N_1506,N_1568);
xnor U2037 (N_2037,N_1510,N_1545);
xnor U2038 (N_2038,N_1526,N_1715);
xor U2039 (N_2039,N_1735,N_1528);
or U2040 (N_2040,N_1750,N_1962);
and U2041 (N_2041,N_1922,N_1853);
nand U2042 (N_2042,N_1591,N_1574);
nor U2043 (N_2043,N_1694,N_1599);
xor U2044 (N_2044,N_1587,N_1513);
and U2045 (N_2045,N_1920,N_1518);
or U2046 (N_2046,N_1713,N_1552);
nor U2047 (N_2047,N_1716,N_1753);
nand U2048 (N_2048,N_1905,N_1579);
nor U2049 (N_2049,N_1719,N_1641);
or U2050 (N_2050,N_1627,N_1673);
nor U2051 (N_2051,N_1900,N_1856);
and U2052 (N_2052,N_1927,N_1803);
nor U2053 (N_2053,N_1665,N_1911);
and U2054 (N_2054,N_1728,N_1752);
nand U2055 (N_2055,N_1951,N_1547);
nand U2056 (N_2056,N_1829,N_1877);
or U2057 (N_2057,N_1890,N_1561);
and U2058 (N_2058,N_1912,N_1650);
xnor U2059 (N_2059,N_1682,N_1805);
xnor U2060 (N_2060,N_1663,N_1833);
or U2061 (N_2061,N_1527,N_1914);
xnor U2062 (N_2062,N_1585,N_1630);
and U2063 (N_2063,N_1670,N_1828);
or U2064 (N_2064,N_1843,N_1538);
nand U2065 (N_2065,N_1982,N_1849);
nor U2066 (N_2066,N_1994,N_1799);
and U2067 (N_2067,N_1542,N_1653);
nor U2068 (N_2068,N_1950,N_1558);
and U2069 (N_2069,N_1657,N_1672);
nand U2070 (N_2070,N_1645,N_1940);
xor U2071 (N_2071,N_1941,N_1631);
and U2072 (N_2072,N_1855,N_1969);
nand U2073 (N_2073,N_1638,N_1978);
or U2074 (N_2074,N_1590,N_1678);
xor U2075 (N_2075,N_1668,N_1942);
nand U2076 (N_2076,N_1550,N_1620);
or U2077 (N_2077,N_1777,N_1825);
and U2078 (N_2078,N_1581,N_1733);
xnor U2079 (N_2079,N_1661,N_1909);
xor U2080 (N_2080,N_1863,N_1971);
and U2081 (N_2081,N_1603,N_1776);
or U2082 (N_2082,N_1894,N_1624);
nand U2083 (N_2083,N_1659,N_1870);
nand U2084 (N_2084,N_1747,N_1946);
and U2085 (N_2085,N_1830,N_1516);
or U2086 (N_2086,N_1575,N_1676);
nand U2087 (N_2087,N_1774,N_1647);
or U2088 (N_2088,N_1996,N_1614);
and U2089 (N_2089,N_1544,N_1896);
and U2090 (N_2090,N_1718,N_1723);
or U2091 (N_2091,N_1862,N_1727);
xor U2092 (N_2092,N_1623,N_1529);
xor U2093 (N_2093,N_1610,N_1714);
nor U2094 (N_2094,N_1635,N_1976);
or U2095 (N_2095,N_1539,N_1874);
and U2096 (N_2096,N_1725,N_1907);
and U2097 (N_2097,N_1688,N_1802);
xor U2098 (N_2098,N_1743,N_1613);
and U2099 (N_2099,N_1608,N_1824);
or U2100 (N_2100,N_1671,N_1762);
nor U2101 (N_2101,N_1546,N_1625);
xnor U2102 (N_2102,N_1788,N_1893);
or U2103 (N_2103,N_1636,N_1642);
or U2104 (N_2104,N_1633,N_1954);
xor U2105 (N_2105,N_1586,N_1744);
or U2106 (N_2106,N_1734,N_1536);
and U2107 (N_2107,N_1760,N_1606);
xnor U2108 (N_2108,N_1720,N_1991);
xnor U2109 (N_2109,N_1998,N_1564);
xor U2110 (N_2110,N_1571,N_1999);
or U2111 (N_2111,N_1939,N_1592);
and U2112 (N_2112,N_1605,N_1966);
xor U2113 (N_2113,N_1895,N_1957);
xnor U2114 (N_2114,N_1980,N_1680);
xnor U2115 (N_2115,N_1860,N_1557);
xor U2116 (N_2116,N_1616,N_1933);
or U2117 (N_2117,N_1541,N_1949);
and U2118 (N_2118,N_1704,N_1847);
nor U2119 (N_2119,N_1683,N_1782);
nor U2120 (N_2120,N_1757,N_1888);
nor U2121 (N_2121,N_1577,N_1918);
or U2122 (N_2122,N_1961,N_1617);
nor U2123 (N_2123,N_1901,N_1724);
and U2124 (N_2124,N_1698,N_1511);
xor U2125 (N_2125,N_1746,N_1508);
nand U2126 (N_2126,N_1903,N_1565);
nand U2127 (N_2127,N_1640,N_1809);
or U2128 (N_2128,N_1540,N_1593);
xnor U2129 (N_2129,N_1594,N_1622);
nor U2130 (N_2130,N_1726,N_1669);
and U2131 (N_2131,N_1973,N_1768);
and U2132 (N_2132,N_1869,N_1555);
xnor U2133 (N_2133,N_1987,N_1705);
or U2134 (N_2134,N_1958,N_1972);
nor U2135 (N_2135,N_1995,N_1722);
nor U2136 (N_2136,N_1928,N_1779);
nor U2137 (N_2137,N_1797,N_1648);
and U2138 (N_2138,N_1523,N_1968);
or U2139 (N_2139,N_1754,N_1604);
xor U2140 (N_2140,N_1868,N_1618);
nor U2141 (N_2141,N_1514,N_1721);
xor U2142 (N_2142,N_1749,N_1923);
and U2143 (N_2143,N_1857,N_1807);
nor U2144 (N_2144,N_1795,N_1674);
and U2145 (N_2145,N_1960,N_1876);
or U2146 (N_2146,N_1687,N_1935);
nand U2147 (N_2147,N_1836,N_1916);
xor U2148 (N_2148,N_1984,N_1850);
and U2149 (N_2149,N_1566,N_1559);
xor U2150 (N_2150,N_1965,N_1602);
nor U2151 (N_2151,N_1891,N_1931);
xnor U2152 (N_2152,N_1500,N_1848);
nor U2153 (N_2153,N_1649,N_1934);
or U2154 (N_2154,N_1562,N_1667);
nor U2155 (N_2155,N_1643,N_1769);
xnor U2156 (N_2156,N_1959,N_1838);
and U2157 (N_2157,N_1864,N_1505);
nand U2158 (N_2158,N_1801,N_1808);
or U2159 (N_2159,N_1986,N_1821);
or U2160 (N_2160,N_1948,N_1915);
and U2161 (N_2161,N_1582,N_1793);
nand U2162 (N_2162,N_1740,N_1861);
nand U2163 (N_2163,N_1576,N_1686);
and U2164 (N_2164,N_1589,N_1696);
nor U2165 (N_2165,N_1588,N_1706);
xor U2166 (N_2166,N_1859,N_1992);
nand U2167 (N_2167,N_1525,N_1601);
xnor U2168 (N_2168,N_1832,N_1741);
nor U2169 (N_2169,N_1772,N_1621);
or U2170 (N_2170,N_1810,N_1745);
or U2171 (N_2171,N_1873,N_1551);
nor U2172 (N_2172,N_1975,N_1781);
xnor U2173 (N_2173,N_1953,N_1512);
or U2174 (N_2174,N_1947,N_1679);
nand U2175 (N_2175,N_1712,N_1883);
or U2176 (N_2176,N_1549,N_1597);
or U2177 (N_2177,N_1681,N_1609);
and U2178 (N_2178,N_1739,N_1619);
nand U2179 (N_2179,N_1729,N_1732);
and U2180 (N_2180,N_1985,N_1798);
nor U2181 (N_2181,N_1600,N_1736);
nand U2182 (N_2182,N_1664,N_1535);
and U2183 (N_2183,N_1533,N_1880);
and U2184 (N_2184,N_1790,N_1932);
and U2185 (N_2185,N_1708,N_1737);
xnor U2186 (N_2186,N_1813,N_1759);
nand U2187 (N_2187,N_1697,N_1583);
or U2188 (N_2188,N_1783,N_1707);
nor U2189 (N_2189,N_1632,N_1658);
and U2190 (N_2190,N_1930,N_1904);
nand U2191 (N_2191,N_1615,N_1693);
and U2192 (N_2192,N_1937,N_1709);
or U2193 (N_2193,N_1654,N_1956);
and U2194 (N_2194,N_1748,N_1926);
nor U2195 (N_2195,N_1634,N_1569);
or U2196 (N_2196,N_1792,N_1924);
nand U2197 (N_2197,N_1519,N_1983);
and U2198 (N_2198,N_1717,N_1865);
nor U2199 (N_2199,N_1785,N_1607);
xor U2200 (N_2200,N_1730,N_1501);
and U2201 (N_2201,N_1738,N_1919);
and U2202 (N_2202,N_1651,N_1507);
nor U2203 (N_2203,N_1675,N_1652);
xnor U2204 (N_2204,N_1656,N_1755);
and U2205 (N_2205,N_1556,N_1521);
nor U2206 (N_2206,N_1816,N_1789);
xnor U2207 (N_2207,N_1612,N_1884);
nor U2208 (N_2208,N_1820,N_1892);
nor U2209 (N_2209,N_1509,N_1970);
and U2210 (N_2210,N_1689,N_1628);
nor U2211 (N_2211,N_1881,N_1530);
xnor U2212 (N_2212,N_1967,N_1989);
nand U2213 (N_2213,N_1812,N_1761);
nor U2214 (N_2214,N_1938,N_1629);
xnor U2215 (N_2215,N_1800,N_1660);
or U2216 (N_2216,N_1872,N_1796);
and U2217 (N_2217,N_1560,N_1692);
or U2218 (N_2218,N_1841,N_1711);
xnor U2219 (N_2219,N_1834,N_1925);
xnor U2220 (N_2220,N_1791,N_1858);
xnor U2221 (N_2221,N_1520,N_1936);
nor U2222 (N_2222,N_1786,N_1943);
nor U2223 (N_2223,N_1818,N_1778);
xor U2224 (N_2224,N_1898,N_1534);
xor U2225 (N_2225,N_1580,N_1567);
nor U2226 (N_2226,N_1710,N_1763);
or U2227 (N_2227,N_1691,N_1814);
nor U2228 (N_2228,N_1666,N_1775);
xor U2229 (N_2229,N_1921,N_1844);
nor U2230 (N_2230,N_1517,N_1822);
nor U2231 (N_2231,N_1979,N_1554);
nor U2232 (N_2232,N_1596,N_1780);
xnor U2233 (N_2233,N_1990,N_1787);
and U2234 (N_2234,N_1835,N_1910);
nor U2235 (N_2235,N_1887,N_1731);
nor U2236 (N_2236,N_1913,N_1532);
nand U2237 (N_2237,N_1695,N_1917);
and U2238 (N_2238,N_1899,N_1955);
nand U2239 (N_2239,N_1882,N_1815);
or U2240 (N_2240,N_1598,N_1767);
xor U2241 (N_2241,N_1837,N_1572);
xnor U2242 (N_2242,N_1626,N_1644);
xor U2243 (N_2243,N_1700,N_1504);
nor U2244 (N_2244,N_1878,N_1889);
nor U2245 (N_2245,N_1766,N_1502);
nand U2246 (N_2246,N_1771,N_1827);
nand U2247 (N_2247,N_1963,N_1662);
and U2248 (N_2248,N_1563,N_1875);
nor U2249 (N_2249,N_1826,N_1997);
nand U2250 (N_2250,N_1662,N_1836);
nor U2251 (N_2251,N_1917,N_1818);
and U2252 (N_2252,N_1630,N_1668);
nand U2253 (N_2253,N_1758,N_1673);
xnor U2254 (N_2254,N_1781,N_1865);
or U2255 (N_2255,N_1583,N_1853);
or U2256 (N_2256,N_1728,N_1789);
or U2257 (N_2257,N_1808,N_1760);
xnor U2258 (N_2258,N_1817,N_1642);
nor U2259 (N_2259,N_1614,N_1910);
xor U2260 (N_2260,N_1769,N_1553);
and U2261 (N_2261,N_1803,N_1511);
nor U2262 (N_2262,N_1886,N_1797);
or U2263 (N_2263,N_1663,N_1563);
nor U2264 (N_2264,N_1974,N_1829);
xor U2265 (N_2265,N_1881,N_1722);
nor U2266 (N_2266,N_1617,N_1952);
and U2267 (N_2267,N_1797,N_1740);
xnor U2268 (N_2268,N_1909,N_1770);
or U2269 (N_2269,N_1674,N_1818);
or U2270 (N_2270,N_1743,N_1919);
and U2271 (N_2271,N_1973,N_1988);
or U2272 (N_2272,N_1649,N_1984);
xnor U2273 (N_2273,N_1598,N_1797);
xor U2274 (N_2274,N_1786,N_1592);
or U2275 (N_2275,N_1911,N_1746);
xnor U2276 (N_2276,N_1620,N_1822);
or U2277 (N_2277,N_1620,N_1836);
or U2278 (N_2278,N_1699,N_1942);
xor U2279 (N_2279,N_1833,N_1741);
or U2280 (N_2280,N_1845,N_1795);
nand U2281 (N_2281,N_1633,N_1729);
nor U2282 (N_2282,N_1949,N_1512);
nand U2283 (N_2283,N_1875,N_1547);
nor U2284 (N_2284,N_1949,N_1872);
xnor U2285 (N_2285,N_1683,N_1708);
and U2286 (N_2286,N_1557,N_1797);
nor U2287 (N_2287,N_1925,N_1572);
nor U2288 (N_2288,N_1819,N_1866);
and U2289 (N_2289,N_1713,N_1866);
nand U2290 (N_2290,N_1505,N_1567);
or U2291 (N_2291,N_1907,N_1983);
and U2292 (N_2292,N_1789,N_1742);
or U2293 (N_2293,N_1837,N_1582);
nor U2294 (N_2294,N_1723,N_1837);
nor U2295 (N_2295,N_1922,N_1918);
nand U2296 (N_2296,N_1564,N_1699);
nor U2297 (N_2297,N_1755,N_1738);
and U2298 (N_2298,N_1576,N_1589);
xnor U2299 (N_2299,N_1845,N_1861);
nor U2300 (N_2300,N_1599,N_1828);
and U2301 (N_2301,N_1592,N_1713);
or U2302 (N_2302,N_1890,N_1855);
nand U2303 (N_2303,N_1725,N_1729);
or U2304 (N_2304,N_1779,N_1876);
nor U2305 (N_2305,N_1728,N_1621);
and U2306 (N_2306,N_1726,N_1865);
nand U2307 (N_2307,N_1653,N_1710);
and U2308 (N_2308,N_1797,N_1614);
nand U2309 (N_2309,N_1656,N_1597);
nor U2310 (N_2310,N_1698,N_1563);
nand U2311 (N_2311,N_1758,N_1613);
xor U2312 (N_2312,N_1561,N_1526);
nand U2313 (N_2313,N_1930,N_1876);
and U2314 (N_2314,N_1615,N_1746);
and U2315 (N_2315,N_1929,N_1598);
and U2316 (N_2316,N_1512,N_1708);
nand U2317 (N_2317,N_1740,N_1529);
xnor U2318 (N_2318,N_1636,N_1530);
nand U2319 (N_2319,N_1781,N_1771);
nor U2320 (N_2320,N_1906,N_1691);
xor U2321 (N_2321,N_1917,N_1789);
and U2322 (N_2322,N_1589,N_1954);
nor U2323 (N_2323,N_1700,N_1841);
nor U2324 (N_2324,N_1879,N_1725);
xor U2325 (N_2325,N_1675,N_1969);
xor U2326 (N_2326,N_1909,N_1538);
xor U2327 (N_2327,N_1821,N_1505);
or U2328 (N_2328,N_1583,N_1762);
nor U2329 (N_2329,N_1679,N_1886);
xnor U2330 (N_2330,N_1829,N_1840);
or U2331 (N_2331,N_1787,N_1605);
and U2332 (N_2332,N_1501,N_1719);
and U2333 (N_2333,N_1663,N_1789);
xor U2334 (N_2334,N_1635,N_1574);
nor U2335 (N_2335,N_1790,N_1937);
and U2336 (N_2336,N_1542,N_1639);
and U2337 (N_2337,N_1922,N_1714);
xnor U2338 (N_2338,N_1617,N_1766);
and U2339 (N_2339,N_1540,N_1756);
nand U2340 (N_2340,N_1589,N_1586);
nand U2341 (N_2341,N_1631,N_1750);
and U2342 (N_2342,N_1742,N_1869);
nor U2343 (N_2343,N_1847,N_1936);
xor U2344 (N_2344,N_1849,N_1665);
xnor U2345 (N_2345,N_1943,N_1847);
nand U2346 (N_2346,N_1596,N_1727);
xor U2347 (N_2347,N_1927,N_1889);
or U2348 (N_2348,N_1631,N_1768);
nor U2349 (N_2349,N_1863,N_1921);
xnor U2350 (N_2350,N_1501,N_1902);
nor U2351 (N_2351,N_1705,N_1962);
xnor U2352 (N_2352,N_1985,N_1972);
or U2353 (N_2353,N_1940,N_1619);
xor U2354 (N_2354,N_1734,N_1945);
xor U2355 (N_2355,N_1913,N_1820);
or U2356 (N_2356,N_1779,N_1570);
nand U2357 (N_2357,N_1751,N_1605);
and U2358 (N_2358,N_1849,N_1835);
nor U2359 (N_2359,N_1918,N_1640);
nand U2360 (N_2360,N_1637,N_1653);
nand U2361 (N_2361,N_1858,N_1589);
or U2362 (N_2362,N_1985,N_1714);
nand U2363 (N_2363,N_1777,N_1519);
nor U2364 (N_2364,N_1902,N_1799);
or U2365 (N_2365,N_1516,N_1955);
or U2366 (N_2366,N_1938,N_1892);
nand U2367 (N_2367,N_1516,N_1566);
nand U2368 (N_2368,N_1937,N_1537);
or U2369 (N_2369,N_1872,N_1820);
nand U2370 (N_2370,N_1783,N_1595);
xnor U2371 (N_2371,N_1614,N_1724);
nor U2372 (N_2372,N_1528,N_1515);
nor U2373 (N_2373,N_1650,N_1936);
nor U2374 (N_2374,N_1878,N_1722);
and U2375 (N_2375,N_1897,N_1575);
nor U2376 (N_2376,N_1883,N_1901);
nand U2377 (N_2377,N_1799,N_1990);
or U2378 (N_2378,N_1888,N_1927);
nand U2379 (N_2379,N_1923,N_1977);
nor U2380 (N_2380,N_1938,N_1901);
nor U2381 (N_2381,N_1638,N_1656);
or U2382 (N_2382,N_1695,N_1723);
nor U2383 (N_2383,N_1639,N_1938);
nor U2384 (N_2384,N_1873,N_1819);
or U2385 (N_2385,N_1792,N_1747);
or U2386 (N_2386,N_1645,N_1582);
or U2387 (N_2387,N_1774,N_1851);
xor U2388 (N_2388,N_1940,N_1923);
or U2389 (N_2389,N_1556,N_1908);
xnor U2390 (N_2390,N_1847,N_1855);
xor U2391 (N_2391,N_1619,N_1978);
xnor U2392 (N_2392,N_1962,N_1979);
xor U2393 (N_2393,N_1505,N_1694);
nor U2394 (N_2394,N_1515,N_1893);
nand U2395 (N_2395,N_1596,N_1511);
nor U2396 (N_2396,N_1931,N_1999);
and U2397 (N_2397,N_1930,N_1619);
or U2398 (N_2398,N_1514,N_1867);
nor U2399 (N_2399,N_1860,N_1984);
or U2400 (N_2400,N_1651,N_1737);
nand U2401 (N_2401,N_1836,N_1554);
nor U2402 (N_2402,N_1567,N_1629);
or U2403 (N_2403,N_1526,N_1860);
or U2404 (N_2404,N_1861,N_1783);
and U2405 (N_2405,N_1876,N_1991);
nor U2406 (N_2406,N_1631,N_1704);
and U2407 (N_2407,N_1585,N_1639);
xnor U2408 (N_2408,N_1585,N_1565);
and U2409 (N_2409,N_1964,N_1788);
and U2410 (N_2410,N_1556,N_1876);
or U2411 (N_2411,N_1799,N_1813);
xor U2412 (N_2412,N_1732,N_1994);
xnor U2413 (N_2413,N_1949,N_1615);
nand U2414 (N_2414,N_1884,N_1667);
and U2415 (N_2415,N_1835,N_1866);
or U2416 (N_2416,N_1879,N_1614);
xnor U2417 (N_2417,N_1559,N_1509);
and U2418 (N_2418,N_1904,N_1817);
xor U2419 (N_2419,N_1538,N_1903);
and U2420 (N_2420,N_1829,N_1632);
or U2421 (N_2421,N_1773,N_1985);
xnor U2422 (N_2422,N_1537,N_1944);
or U2423 (N_2423,N_1957,N_1548);
xnor U2424 (N_2424,N_1809,N_1660);
nand U2425 (N_2425,N_1710,N_1652);
nand U2426 (N_2426,N_1781,N_1648);
nor U2427 (N_2427,N_1551,N_1776);
and U2428 (N_2428,N_1997,N_1708);
and U2429 (N_2429,N_1747,N_1808);
nor U2430 (N_2430,N_1824,N_1725);
nand U2431 (N_2431,N_1968,N_1956);
nand U2432 (N_2432,N_1948,N_1523);
nand U2433 (N_2433,N_1850,N_1512);
and U2434 (N_2434,N_1563,N_1966);
xor U2435 (N_2435,N_1679,N_1690);
nor U2436 (N_2436,N_1676,N_1712);
and U2437 (N_2437,N_1754,N_1528);
xnor U2438 (N_2438,N_1505,N_1665);
xor U2439 (N_2439,N_1909,N_1958);
xnor U2440 (N_2440,N_1967,N_1992);
or U2441 (N_2441,N_1500,N_1964);
or U2442 (N_2442,N_1940,N_1795);
nor U2443 (N_2443,N_1967,N_1862);
xor U2444 (N_2444,N_1808,N_1886);
and U2445 (N_2445,N_1543,N_1517);
or U2446 (N_2446,N_1920,N_1979);
or U2447 (N_2447,N_1615,N_1983);
xnor U2448 (N_2448,N_1823,N_1655);
nor U2449 (N_2449,N_1536,N_1560);
and U2450 (N_2450,N_1610,N_1750);
nand U2451 (N_2451,N_1713,N_1842);
or U2452 (N_2452,N_1765,N_1989);
and U2453 (N_2453,N_1847,N_1724);
and U2454 (N_2454,N_1646,N_1884);
and U2455 (N_2455,N_1815,N_1538);
xnor U2456 (N_2456,N_1695,N_1594);
and U2457 (N_2457,N_1520,N_1711);
nand U2458 (N_2458,N_1819,N_1592);
nand U2459 (N_2459,N_1545,N_1913);
nor U2460 (N_2460,N_1949,N_1622);
or U2461 (N_2461,N_1737,N_1822);
and U2462 (N_2462,N_1514,N_1752);
xor U2463 (N_2463,N_1761,N_1935);
or U2464 (N_2464,N_1886,N_1569);
and U2465 (N_2465,N_1843,N_1638);
nand U2466 (N_2466,N_1838,N_1816);
xor U2467 (N_2467,N_1808,N_1695);
xor U2468 (N_2468,N_1621,N_1813);
xnor U2469 (N_2469,N_1753,N_1964);
or U2470 (N_2470,N_1507,N_1652);
xor U2471 (N_2471,N_1942,N_1863);
nor U2472 (N_2472,N_1984,N_1847);
or U2473 (N_2473,N_1899,N_1803);
nand U2474 (N_2474,N_1984,N_1921);
or U2475 (N_2475,N_1578,N_1781);
nor U2476 (N_2476,N_1529,N_1531);
nand U2477 (N_2477,N_1891,N_1582);
nand U2478 (N_2478,N_1724,N_1838);
nand U2479 (N_2479,N_1953,N_1616);
nand U2480 (N_2480,N_1658,N_1531);
and U2481 (N_2481,N_1910,N_1552);
and U2482 (N_2482,N_1776,N_1977);
and U2483 (N_2483,N_1760,N_1731);
or U2484 (N_2484,N_1650,N_1506);
nor U2485 (N_2485,N_1785,N_1923);
nand U2486 (N_2486,N_1541,N_1549);
and U2487 (N_2487,N_1899,N_1585);
and U2488 (N_2488,N_1691,N_1677);
nand U2489 (N_2489,N_1930,N_1725);
nand U2490 (N_2490,N_1713,N_1655);
xnor U2491 (N_2491,N_1628,N_1661);
nand U2492 (N_2492,N_1980,N_1727);
nand U2493 (N_2493,N_1831,N_1961);
nor U2494 (N_2494,N_1734,N_1717);
xor U2495 (N_2495,N_1763,N_1944);
or U2496 (N_2496,N_1949,N_1906);
nand U2497 (N_2497,N_1574,N_1844);
or U2498 (N_2498,N_1725,N_1886);
or U2499 (N_2499,N_1873,N_1989);
xnor U2500 (N_2500,N_2196,N_2223);
and U2501 (N_2501,N_2391,N_2475);
nor U2502 (N_2502,N_2377,N_2346);
or U2503 (N_2503,N_2247,N_2118);
nor U2504 (N_2504,N_2380,N_2256);
nand U2505 (N_2505,N_2032,N_2108);
nor U2506 (N_2506,N_2075,N_2498);
xor U2507 (N_2507,N_2365,N_2202);
and U2508 (N_2508,N_2422,N_2402);
or U2509 (N_2509,N_2191,N_2338);
nand U2510 (N_2510,N_2178,N_2213);
or U2511 (N_2511,N_2471,N_2084);
nand U2512 (N_2512,N_2340,N_2214);
nor U2513 (N_2513,N_2451,N_2427);
xnor U2514 (N_2514,N_2296,N_2418);
xnor U2515 (N_2515,N_2160,N_2155);
xor U2516 (N_2516,N_2269,N_2231);
or U2517 (N_2517,N_2126,N_2114);
nand U2518 (N_2518,N_2326,N_2490);
or U2519 (N_2519,N_2112,N_2021);
xnor U2520 (N_2520,N_2235,N_2428);
xor U2521 (N_2521,N_2203,N_2210);
xor U2522 (N_2522,N_2394,N_2024);
and U2523 (N_2523,N_2388,N_2455);
nand U2524 (N_2524,N_2005,N_2392);
nand U2525 (N_2525,N_2122,N_2264);
xor U2526 (N_2526,N_2142,N_2423);
nand U2527 (N_2527,N_2218,N_2016);
nor U2528 (N_2528,N_2248,N_2329);
nor U2529 (N_2529,N_2305,N_2297);
nand U2530 (N_2530,N_2258,N_2336);
nand U2531 (N_2531,N_2023,N_2315);
or U2532 (N_2532,N_2077,N_2290);
or U2533 (N_2533,N_2435,N_2378);
nand U2534 (N_2534,N_2182,N_2458);
nor U2535 (N_2535,N_2390,N_2104);
nand U2536 (N_2536,N_2241,N_2197);
or U2537 (N_2537,N_2148,N_2113);
or U2538 (N_2538,N_2071,N_2496);
nand U2539 (N_2539,N_2445,N_2224);
nand U2540 (N_2540,N_2366,N_2416);
nor U2541 (N_2541,N_2288,N_2403);
xnor U2542 (N_2542,N_2470,N_2359);
nor U2543 (N_2543,N_2041,N_2204);
xor U2544 (N_2544,N_2215,N_2281);
or U2545 (N_2545,N_2385,N_2234);
nor U2546 (N_2546,N_2065,N_2335);
xor U2547 (N_2547,N_2370,N_2246);
nor U2548 (N_2548,N_2238,N_2389);
xnor U2549 (N_2549,N_2372,N_2439);
nand U2550 (N_2550,N_2141,N_2476);
nor U2551 (N_2551,N_2276,N_2482);
nor U2552 (N_2552,N_2310,N_2229);
xor U2553 (N_2553,N_2300,N_2056);
xor U2554 (N_2554,N_2183,N_2250);
nand U2555 (N_2555,N_2257,N_2134);
and U2556 (N_2556,N_2230,N_2199);
xor U2557 (N_2557,N_2173,N_2293);
and U2558 (N_2558,N_2187,N_2322);
or U2559 (N_2559,N_2103,N_2325);
xor U2560 (N_2560,N_2059,N_2170);
xor U2561 (N_2561,N_2344,N_2318);
and U2562 (N_2562,N_2384,N_2282);
nor U2563 (N_2563,N_2363,N_2468);
xnor U2564 (N_2564,N_2124,N_2164);
and U2565 (N_2565,N_2254,N_2031);
nor U2566 (N_2566,N_2180,N_2186);
nor U2567 (N_2567,N_2376,N_2312);
and U2568 (N_2568,N_2437,N_2003);
or U2569 (N_2569,N_2062,N_2166);
and U2570 (N_2570,N_2261,N_2401);
nand U2571 (N_2571,N_2111,N_2280);
nor U2572 (N_2572,N_2324,N_2371);
nand U2573 (N_2573,N_2440,N_2308);
and U2574 (N_2574,N_2125,N_2117);
or U2575 (N_2575,N_2342,N_2047);
or U2576 (N_2576,N_2158,N_2253);
and U2577 (N_2577,N_2063,N_2429);
nand U2578 (N_2578,N_2162,N_2013);
nand U2579 (N_2579,N_2441,N_2033);
or U2580 (N_2580,N_2074,N_2138);
xor U2581 (N_2581,N_2036,N_2414);
nor U2582 (N_2582,N_2201,N_2494);
and U2583 (N_2583,N_2327,N_2045);
nand U2584 (N_2584,N_2069,N_2129);
nand U2585 (N_2585,N_2337,N_2452);
nand U2586 (N_2586,N_2053,N_2292);
or U2587 (N_2587,N_2497,N_2265);
nand U2588 (N_2588,N_2219,N_2167);
and U2589 (N_2589,N_2017,N_2382);
nand U2590 (N_2590,N_2145,N_2472);
nand U2591 (N_2591,N_2492,N_2369);
or U2592 (N_2592,N_2454,N_2188);
nand U2593 (N_2593,N_2298,N_2448);
nand U2594 (N_2594,N_2411,N_2493);
and U2595 (N_2595,N_2295,N_2050);
xnor U2596 (N_2596,N_2347,N_2198);
nor U2597 (N_2597,N_2499,N_2128);
or U2598 (N_2598,N_2172,N_2110);
and U2599 (N_2599,N_2192,N_2177);
or U2600 (N_2600,N_2115,N_2473);
nor U2601 (N_2601,N_2152,N_2027);
nor U2602 (N_2602,N_2406,N_2139);
or U2603 (N_2603,N_2156,N_2130);
nand U2604 (N_2604,N_2207,N_2102);
and U2605 (N_2605,N_2465,N_2267);
nor U2606 (N_2606,N_2277,N_2467);
and U2607 (N_2607,N_2011,N_2009);
xnor U2608 (N_2608,N_2474,N_2284);
and U2609 (N_2609,N_2132,N_2313);
or U2610 (N_2610,N_2463,N_2189);
nand U2611 (N_2611,N_2133,N_2299);
nand U2612 (N_2612,N_2405,N_2044);
and U2613 (N_2613,N_2309,N_2285);
xor U2614 (N_2614,N_2030,N_2483);
nand U2615 (N_2615,N_2099,N_2195);
nor U2616 (N_2616,N_2491,N_2485);
or U2617 (N_2617,N_2364,N_2002);
or U2618 (N_2618,N_2398,N_2438);
xnor U2619 (N_2619,N_2457,N_2413);
xnor U2620 (N_2620,N_2123,N_2239);
or U2621 (N_2621,N_2143,N_2205);
nor U2622 (N_2622,N_2450,N_2120);
or U2623 (N_2623,N_2449,N_2456);
xor U2624 (N_2624,N_2286,N_2028);
or U2625 (N_2625,N_2150,N_2354);
and U2626 (N_2626,N_2080,N_2109);
xor U2627 (N_2627,N_2147,N_2291);
nor U2628 (N_2628,N_2159,N_2270);
nor U2629 (N_2629,N_2131,N_2168);
nor U2630 (N_2630,N_2090,N_2049);
xnor U2631 (N_2631,N_2311,N_2228);
xor U2632 (N_2632,N_2443,N_2176);
nand U2633 (N_2633,N_2432,N_2034);
nor U2634 (N_2634,N_2301,N_2420);
and U2635 (N_2635,N_2067,N_2426);
xnor U2636 (N_2636,N_2073,N_2092);
and U2637 (N_2637,N_2208,N_2442);
nor U2638 (N_2638,N_2042,N_2165);
or U2639 (N_2639,N_2360,N_2163);
and U2640 (N_2640,N_2070,N_2051);
or U2641 (N_2641,N_2477,N_2430);
xnor U2642 (N_2642,N_2237,N_2425);
and U2643 (N_2643,N_2357,N_2466);
or U2644 (N_2644,N_2105,N_2040);
nor U2645 (N_2645,N_2140,N_2400);
nand U2646 (N_2646,N_2495,N_2415);
xnor U2647 (N_2647,N_2333,N_2314);
nand U2648 (N_2648,N_2351,N_2343);
or U2649 (N_2649,N_2144,N_2091);
or U2650 (N_2650,N_2339,N_2487);
nor U2651 (N_2651,N_2025,N_2259);
nor U2652 (N_2652,N_2368,N_2096);
nor U2653 (N_2653,N_2236,N_2227);
or U2654 (N_2654,N_2066,N_2043);
nand U2655 (N_2655,N_2396,N_2233);
nand U2656 (N_2656,N_2181,N_2184);
xor U2657 (N_2657,N_2484,N_2319);
nor U2658 (N_2658,N_2085,N_2054);
nand U2659 (N_2659,N_2387,N_2263);
and U2660 (N_2660,N_2345,N_2375);
xnor U2661 (N_2661,N_2060,N_2022);
or U2662 (N_2662,N_2464,N_2217);
nand U2663 (N_2663,N_2107,N_2433);
xnor U2664 (N_2664,N_2179,N_2412);
xnor U2665 (N_2665,N_2057,N_2149);
nand U2666 (N_2666,N_2193,N_2459);
nand U2667 (N_2667,N_2006,N_2037);
xor U2668 (N_2668,N_2220,N_2079);
or U2669 (N_2669,N_2488,N_2287);
nand U2670 (N_2670,N_2331,N_2424);
and U2671 (N_2671,N_2018,N_2101);
nand U2672 (N_2672,N_2489,N_2175);
nor U2673 (N_2673,N_2244,N_2279);
or U2674 (N_2674,N_2039,N_2012);
nor U2675 (N_2675,N_2094,N_2408);
xor U2676 (N_2676,N_2431,N_2206);
and U2677 (N_2677,N_2446,N_2081);
or U2678 (N_2678,N_2478,N_2019);
nor U2679 (N_2679,N_2086,N_2061);
xor U2680 (N_2680,N_2272,N_2460);
and U2681 (N_2681,N_2127,N_2255);
xnor U2682 (N_2682,N_2260,N_2444);
nand U2683 (N_2683,N_2352,N_2209);
nor U2684 (N_2684,N_2146,N_2232);
nand U2685 (N_2685,N_2038,N_2046);
xor U2686 (N_2686,N_2216,N_2356);
xnor U2687 (N_2687,N_2243,N_2151);
and U2688 (N_2688,N_2303,N_2082);
and U2689 (N_2689,N_2273,N_2486);
and U2690 (N_2690,N_2137,N_2447);
xor U2691 (N_2691,N_2421,N_2302);
xor U2692 (N_2692,N_2271,N_2020);
xor U2693 (N_2693,N_2349,N_2383);
or U2694 (N_2694,N_2350,N_2095);
nand U2695 (N_2695,N_2434,N_2266);
xnor U2696 (N_2696,N_2479,N_2397);
nand U2697 (N_2697,N_2328,N_2221);
xnor U2698 (N_2698,N_2058,N_2323);
xor U2699 (N_2699,N_2007,N_2334);
and U2700 (N_2700,N_2268,N_2171);
and U2701 (N_2701,N_2409,N_2222);
nor U2702 (N_2702,N_2367,N_2100);
xor U2703 (N_2703,N_2010,N_2064);
nand U2704 (N_2704,N_2052,N_2190);
xor U2705 (N_2705,N_2275,N_2317);
nand U2706 (N_2706,N_2461,N_2076);
nand U2707 (N_2707,N_2395,N_2078);
nor U2708 (N_2708,N_2035,N_2481);
nor U2709 (N_2709,N_2161,N_2157);
and U2710 (N_2710,N_2136,N_2278);
nor U2711 (N_2711,N_2393,N_2245);
or U2712 (N_2712,N_2304,N_2174);
and U2713 (N_2713,N_2361,N_2307);
and U2714 (N_2714,N_2226,N_2469);
nand U2715 (N_2715,N_2055,N_2306);
nor U2716 (N_2716,N_2154,N_2194);
nor U2717 (N_2717,N_2320,N_2480);
nand U2718 (N_2718,N_2294,N_2249);
and U2719 (N_2719,N_2410,N_2088);
nor U2720 (N_2720,N_2212,N_2097);
nor U2721 (N_2721,N_2316,N_2262);
nand U2722 (N_2722,N_2211,N_2106);
and U2723 (N_2723,N_2083,N_2341);
xor U2724 (N_2724,N_2386,N_2283);
xor U2725 (N_2725,N_2252,N_2251);
nand U2726 (N_2726,N_2321,N_2072);
xor U2727 (N_2727,N_2355,N_2381);
nand U2728 (N_2728,N_2332,N_2116);
nand U2729 (N_2729,N_2169,N_2004);
nand U2730 (N_2730,N_2225,N_2358);
nor U2731 (N_2731,N_2153,N_2015);
xnor U2732 (N_2732,N_2121,N_2119);
xnor U2733 (N_2733,N_2379,N_2242);
nor U2734 (N_2734,N_2419,N_2200);
or U2735 (N_2735,N_2399,N_2014);
xnor U2736 (N_2736,N_2048,N_2362);
and U2737 (N_2737,N_2404,N_2135);
nand U2738 (N_2738,N_2353,N_2436);
or U2739 (N_2739,N_2000,N_2407);
or U2740 (N_2740,N_2289,N_2029);
nor U2741 (N_2741,N_2417,N_2008);
xnor U2742 (N_2742,N_2453,N_2274);
nor U2743 (N_2743,N_2462,N_2374);
xnor U2744 (N_2744,N_2330,N_2098);
xor U2745 (N_2745,N_2026,N_2240);
nand U2746 (N_2746,N_2087,N_2089);
and U2747 (N_2747,N_2185,N_2068);
nor U2748 (N_2748,N_2093,N_2348);
and U2749 (N_2749,N_2001,N_2373);
nand U2750 (N_2750,N_2337,N_2450);
xnor U2751 (N_2751,N_2481,N_2255);
nor U2752 (N_2752,N_2069,N_2157);
nor U2753 (N_2753,N_2148,N_2075);
nand U2754 (N_2754,N_2072,N_2120);
nand U2755 (N_2755,N_2090,N_2323);
or U2756 (N_2756,N_2259,N_2188);
nand U2757 (N_2757,N_2305,N_2194);
xnor U2758 (N_2758,N_2029,N_2154);
xor U2759 (N_2759,N_2125,N_2357);
or U2760 (N_2760,N_2128,N_2049);
or U2761 (N_2761,N_2014,N_2235);
or U2762 (N_2762,N_2217,N_2432);
and U2763 (N_2763,N_2135,N_2209);
nor U2764 (N_2764,N_2109,N_2280);
or U2765 (N_2765,N_2214,N_2236);
or U2766 (N_2766,N_2371,N_2157);
nand U2767 (N_2767,N_2164,N_2408);
or U2768 (N_2768,N_2313,N_2396);
nand U2769 (N_2769,N_2002,N_2394);
and U2770 (N_2770,N_2331,N_2219);
or U2771 (N_2771,N_2499,N_2026);
and U2772 (N_2772,N_2314,N_2328);
or U2773 (N_2773,N_2415,N_2403);
or U2774 (N_2774,N_2307,N_2006);
nand U2775 (N_2775,N_2236,N_2354);
xor U2776 (N_2776,N_2112,N_2469);
nor U2777 (N_2777,N_2189,N_2432);
nand U2778 (N_2778,N_2238,N_2164);
nand U2779 (N_2779,N_2231,N_2079);
nor U2780 (N_2780,N_2109,N_2375);
and U2781 (N_2781,N_2395,N_2157);
nor U2782 (N_2782,N_2151,N_2407);
or U2783 (N_2783,N_2420,N_2094);
and U2784 (N_2784,N_2360,N_2331);
xor U2785 (N_2785,N_2294,N_2291);
xor U2786 (N_2786,N_2017,N_2059);
or U2787 (N_2787,N_2214,N_2439);
xnor U2788 (N_2788,N_2147,N_2053);
nand U2789 (N_2789,N_2480,N_2248);
xor U2790 (N_2790,N_2274,N_2268);
and U2791 (N_2791,N_2194,N_2204);
nand U2792 (N_2792,N_2242,N_2358);
nand U2793 (N_2793,N_2262,N_2139);
or U2794 (N_2794,N_2105,N_2252);
nor U2795 (N_2795,N_2065,N_2030);
nand U2796 (N_2796,N_2062,N_2206);
xor U2797 (N_2797,N_2110,N_2077);
and U2798 (N_2798,N_2356,N_2104);
nand U2799 (N_2799,N_2013,N_2405);
xor U2800 (N_2800,N_2192,N_2327);
nor U2801 (N_2801,N_2430,N_2253);
xnor U2802 (N_2802,N_2200,N_2085);
nor U2803 (N_2803,N_2203,N_2401);
nand U2804 (N_2804,N_2289,N_2317);
nand U2805 (N_2805,N_2475,N_2000);
and U2806 (N_2806,N_2070,N_2258);
nand U2807 (N_2807,N_2291,N_2323);
xnor U2808 (N_2808,N_2048,N_2328);
nand U2809 (N_2809,N_2359,N_2316);
or U2810 (N_2810,N_2357,N_2283);
and U2811 (N_2811,N_2419,N_2151);
nor U2812 (N_2812,N_2495,N_2227);
nand U2813 (N_2813,N_2470,N_2125);
or U2814 (N_2814,N_2064,N_2185);
xor U2815 (N_2815,N_2444,N_2051);
and U2816 (N_2816,N_2487,N_2216);
or U2817 (N_2817,N_2475,N_2371);
and U2818 (N_2818,N_2459,N_2427);
xor U2819 (N_2819,N_2253,N_2217);
nor U2820 (N_2820,N_2383,N_2396);
or U2821 (N_2821,N_2197,N_2075);
and U2822 (N_2822,N_2258,N_2166);
nor U2823 (N_2823,N_2116,N_2416);
xnor U2824 (N_2824,N_2227,N_2205);
and U2825 (N_2825,N_2245,N_2388);
and U2826 (N_2826,N_2257,N_2456);
nor U2827 (N_2827,N_2004,N_2493);
or U2828 (N_2828,N_2323,N_2077);
nor U2829 (N_2829,N_2075,N_2115);
nand U2830 (N_2830,N_2250,N_2335);
xnor U2831 (N_2831,N_2212,N_2294);
nand U2832 (N_2832,N_2237,N_2130);
and U2833 (N_2833,N_2445,N_2481);
and U2834 (N_2834,N_2392,N_2366);
xnor U2835 (N_2835,N_2382,N_2240);
xnor U2836 (N_2836,N_2351,N_2494);
nor U2837 (N_2837,N_2022,N_2339);
xor U2838 (N_2838,N_2313,N_2035);
xnor U2839 (N_2839,N_2038,N_2239);
xor U2840 (N_2840,N_2042,N_2262);
and U2841 (N_2841,N_2435,N_2280);
and U2842 (N_2842,N_2202,N_2214);
nand U2843 (N_2843,N_2109,N_2068);
nor U2844 (N_2844,N_2473,N_2325);
and U2845 (N_2845,N_2259,N_2320);
xor U2846 (N_2846,N_2434,N_2485);
nand U2847 (N_2847,N_2369,N_2102);
nand U2848 (N_2848,N_2419,N_2244);
and U2849 (N_2849,N_2194,N_2321);
or U2850 (N_2850,N_2386,N_2463);
nand U2851 (N_2851,N_2230,N_2485);
or U2852 (N_2852,N_2452,N_2314);
or U2853 (N_2853,N_2125,N_2426);
nand U2854 (N_2854,N_2136,N_2496);
xnor U2855 (N_2855,N_2173,N_2444);
xor U2856 (N_2856,N_2467,N_2203);
nand U2857 (N_2857,N_2342,N_2108);
and U2858 (N_2858,N_2151,N_2147);
or U2859 (N_2859,N_2070,N_2313);
nand U2860 (N_2860,N_2073,N_2046);
and U2861 (N_2861,N_2041,N_2487);
or U2862 (N_2862,N_2146,N_2041);
xnor U2863 (N_2863,N_2079,N_2058);
or U2864 (N_2864,N_2270,N_2156);
nor U2865 (N_2865,N_2496,N_2450);
nand U2866 (N_2866,N_2347,N_2062);
nor U2867 (N_2867,N_2382,N_2373);
nor U2868 (N_2868,N_2004,N_2402);
nor U2869 (N_2869,N_2210,N_2099);
or U2870 (N_2870,N_2107,N_2434);
xnor U2871 (N_2871,N_2197,N_2322);
nor U2872 (N_2872,N_2150,N_2102);
and U2873 (N_2873,N_2492,N_2257);
nor U2874 (N_2874,N_2215,N_2213);
or U2875 (N_2875,N_2041,N_2109);
nand U2876 (N_2876,N_2372,N_2480);
nor U2877 (N_2877,N_2355,N_2426);
and U2878 (N_2878,N_2027,N_2351);
or U2879 (N_2879,N_2220,N_2030);
and U2880 (N_2880,N_2311,N_2221);
xor U2881 (N_2881,N_2483,N_2097);
and U2882 (N_2882,N_2177,N_2319);
nor U2883 (N_2883,N_2003,N_2140);
xnor U2884 (N_2884,N_2140,N_2224);
nand U2885 (N_2885,N_2222,N_2485);
nor U2886 (N_2886,N_2403,N_2359);
xnor U2887 (N_2887,N_2391,N_2261);
nand U2888 (N_2888,N_2251,N_2141);
and U2889 (N_2889,N_2306,N_2101);
and U2890 (N_2890,N_2340,N_2396);
xor U2891 (N_2891,N_2333,N_2227);
nor U2892 (N_2892,N_2048,N_2112);
nand U2893 (N_2893,N_2455,N_2287);
nor U2894 (N_2894,N_2348,N_2062);
nor U2895 (N_2895,N_2170,N_2164);
nand U2896 (N_2896,N_2444,N_2023);
xnor U2897 (N_2897,N_2169,N_2150);
nand U2898 (N_2898,N_2322,N_2078);
and U2899 (N_2899,N_2353,N_2413);
and U2900 (N_2900,N_2087,N_2387);
or U2901 (N_2901,N_2414,N_2331);
and U2902 (N_2902,N_2209,N_2138);
xor U2903 (N_2903,N_2192,N_2157);
nand U2904 (N_2904,N_2232,N_2005);
or U2905 (N_2905,N_2280,N_2496);
xnor U2906 (N_2906,N_2143,N_2064);
nor U2907 (N_2907,N_2427,N_2298);
and U2908 (N_2908,N_2109,N_2197);
or U2909 (N_2909,N_2320,N_2292);
nand U2910 (N_2910,N_2204,N_2491);
nor U2911 (N_2911,N_2210,N_2161);
xor U2912 (N_2912,N_2416,N_2341);
xnor U2913 (N_2913,N_2286,N_2031);
nor U2914 (N_2914,N_2433,N_2285);
nor U2915 (N_2915,N_2406,N_2005);
nand U2916 (N_2916,N_2154,N_2018);
nand U2917 (N_2917,N_2346,N_2016);
xor U2918 (N_2918,N_2375,N_2024);
xnor U2919 (N_2919,N_2358,N_2032);
nor U2920 (N_2920,N_2489,N_2462);
nor U2921 (N_2921,N_2372,N_2155);
nor U2922 (N_2922,N_2004,N_2497);
nor U2923 (N_2923,N_2192,N_2075);
nand U2924 (N_2924,N_2176,N_2066);
or U2925 (N_2925,N_2333,N_2356);
and U2926 (N_2926,N_2186,N_2290);
or U2927 (N_2927,N_2009,N_2216);
or U2928 (N_2928,N_2154,N_2198);
xor U2929 (N_2929,N_2390,N_2043);
nand U2930 (N_2930,N_2009,N_2064);
or U2931 (N_2931,N_2045,N_2194);
nand U2932 (N_2932,N_2137,N_2302);
nor U2933 (N_2933,N_2335,N_2130);
xnor U2934 (N_2934,N_2438,N_2217);
nand U2935 (N_2935,N_2161,N_2066);
xor U2936 (N_2936,N_2182,N_2394);
nand U2937 (N_2937,N_2065,N_2474);
xnor U2938 (N_2938,N_2087,N_2070);
or U2939 (N_2939,N_2350,N_2188);
and U2940 (N_2940,N_2410,N_2161);
and U2941 (N_2941,N_2180,N_2060);
or U2942 (N_2942,N_2383,N_2152);
or U2943 (N_2943,N_2167,N_2435);
or U2944 (N_2944,N_2087,N_2450);
and U2945 (N_2945,N_2364,N_2036);
xor U2946 (N_2946,N_2159,N_2306);
nand U2947 (N_2947,N_2340,N_2115);
xor U2948 (N_2948,N_2430,N_2378);
nand U2949 (N_2949,N_2485,N_2196);
and U2950 (N_2950,N_2342,N_2307);
nor U2951 (N_2951,N_2495,N_2278);
nand U2952 (N_2952,N_2125,N_2018);
nor U2953 (N_2953,N_2070,N_2323);
and U2954 (N_2954,N_2328,N_2077);
or U2955 (N_2955,N_2368,N_2020);
and U2956 (N_2956,N_2336,N_2288);
nand U2957 (N_2957,N_2100,N_2396);
and U2958 (N_2958,N_2189,N_2176);
nand U2959 (N_2959,N_2034,N_2301);
or U2960 (N_2960,N_2454,N_2397);
nand U2961 (N_2961,N_2184,N_2164);
or U2962 (N_2962,N_2134,N_2043);
or U2963 (N_2963,N_2447,N_2338);
and U2964 (N_2964,N_2490,N_2183);
and U2965 (N_2965,N_2058,N_2121);
or U2966 (N_2966,N_2255,N_2296);
nor U2967 (N_2967,N_2336,N_2444);
and U2968 (N_2968,N_2121,N_2179);
and U2969 (N_2969,N_2055,N_2002);
nand U2970 (N_2970,N_2298,N_2291);
nor U2971 (N_2971,N_2023,N_2012);
and U2972 (N_2972,N_2245,N_2477);
or U2973 (N_2973,N_2276,N_2165);
or U2974 (N_2974,N_2475,N_2256);
nand U2975 (N_2975,N_2137,N_2083);
nor U2976 (N_2976,N_2176,N_2124);
nand U2977 (N_2977,N_2141,N_2309);
nand U2978 (N_2978,N_2473,N_2351);
nand U2979 (N_2979,N_2447,N_2441);
xnor U2980 (N_2980,N_2348,N_2043);
and U2981 (N_2981,N_2447,N_2284);
nor U2982 (N_2982,N_2209,N_2341);
nor U2983 (N_2983,N_2342,N_2111);
and U2984 (N_2984,N_2187,N_2412);
and U2985 (N_2985,N_2234,N_2240);
nand U2986 (N_2986,N_2378,N_2233);
and U2987 (N_2987,N_2039,N_2463);
xor U2988 (N_2988,N_2169,N_2259);
nand U2989 (N_2989,N_2496,N_2160);
or U2990 (N_2990,N_2418,N_2426);
nand U2991 (N_2991,N_2405,N_2123);
or U2992 (N_2992,N_2023,N_2302);
and U2993 (N_2993,N_2087,N_2152);
nand U2994 (N_2994,N_2324,N_2079);
nor U2995 (N_2995,N_2199,N_2114);
nor U2996 (N_2996,N_2376,N_2226);
or U2997 (N_2997,N_2091,N_2138);
and U2998 (N_2998,N_2278,N_2276);
or U2999 (N_2999,N_2433,N_2331);
and U3000 (N_3000,N_2850,N_2794);
nor U3001 (N_3001,N_2975,N_2685);
and U3002 (N_3002,N_2510,N_2872);
xor U3003 (N_3003,N_2670,N_2675);
xor U3004 (N_3004,N_2797,N_2764);
nor U3005 (N_3005,N_2545,N_2526);
nand U3006 (N_3006,N_2821,N_2658);
and U3007 (N_3007,N_2557,N_2827);
or U3008 (N_3008,N_2819,N_2576);
or U3009 (N_3009,N_2965,N_2911);
nand U3010 (N_3010,N_2815,N_2762);
or U3011 (N_3011,N_2739,N_2852);
nand U3012 (N_3012,N_2532,N_2808);
or U3013 (N_3013,N_2640,N_2707);
xnor U3014 (N_3014,N_2743,N_2980);
xor U3015 (N_3015,N_2527,N_2951);
and U3016 (N_3016,N_2867,N_2514);
nand U3017 (N_3017,N_2522,N_2773);
nor U3018 (N_3018,N_2676,N_2654);
nand U3019 (N_3019,N_2881,N_2958);
and U3020 (N_3020,N_2521,N_2584);
nand U3021 (N_3021,N_2548,N_2864);
nand U3022 (N_3022,N_2542,N_2740);
nand U3023 (N_3023,N_2775,N_2801);
and U3024 (N_3024,N_2563,N_2895);
nor U3025 (N_3025,N_2826,N_2729);
and U3026 (N_3026,N_2841,N_2623);
nand U3027 (N_3027,N_2929,N_2506);
xnor U3028 (N_3028,N_2962,N_2880);
or U3029 (N_3029,N_2870,N_2838);
xnor U3030 (N_3030,N_2596,N_2734);
xnor U3031 (N_3031,N_2984,N_2909);
or U3032 (N_3032,N_2677,N_2611);
or U3033 (N_3033,N_2949,N_2721);
xnor U3034 (N_3034,N_2788,N_2802);
nand U3035 (N_3035,N_2551,N_2568);
nor U3036 (N_3036,N_2846,N_2871);
nand U3037 (N_3037,N_2747,N_2698);
nor U3038 (N_3038,N_2622,N_2795);
or U3039 (N_3039,N_2615,N_2502);
nand U3040 (N_3040,N_2777,N_2631);
xnor U3041 (N_3041,N_2998,N_2919);
and U3042 (N_3042,N_2566,N_2689);
and U3043 (N_3043,N_2784,N_2937);
or U3044 (N_3044,N_2726,N_2778);
and U3045 (N_3045,N_2679,N_2771);
or U3046 (N_3046,N_2508,N_2793);
and U3047 (N_3047,N_2578,N_2530);
and U3048 (N_3048,N_2600,N_2609);
nand U3049 (N_3049,N_2843,N_2603);
nand U3050 (N_3050,N_2905,N_2671);
and U3051 (N_3051,N_2672,N_2684);
xor U3052 (N_3052,N_2883,N_2626);
or U3053 (N_3053,N_2877,N_2644);
nor U3054 (N_3054,N_2906,N_2716);
and U3055 (N_3055,N_2621,N_2928);
or U3056 (N_3056,N_2858,N_2931);
or U3057 (N_3057,N_2760,N_2653);
and U3058 (N_3058,N_2845,N_2755);
xnor U3059 (N_3059,N_2890,N_2648);
nand U3060 (N_3060,N_2925,N_2810);
xnor U3061 (N_3061,N_2770,N_2637);
or U3062 (N_3062,N_2681,N_2702);
xor U3063 (N_3063,N_2878,N_2577);
or U3064 (N_3064,N_2767,N_2590);
or U3065 (N_3065,N_2800,N_2805);
nor U3066 (N_3066,N_2848,N_2900);
xnor U3067 (N_3067,N_2924,N_2692);
xor U3068 (N_3068,N_2572,N_2970);
and U3069 (N_3069,N_2564,N_2741);
nand U3070 (N_3070,N_2941,N_2501);
nor U3071 (N_3071,N_2923,N_2896);
nor U3072 (N_3072,N_2892,N_2792);
xnor U3073 (N_3073,N_2628,N_2632);
or U3074 (N_3074,N_2519,N_2574);
nor U3075 (N_3075,N_2573,N_2515);
xnor U3076 (N_3076,N_2851,N_2948);
and U3077 (N_3077,N_2686,N_2759);
nand U3078 (N_3078,N_2700,N_2668);
and U3079 (N_3079,N_2605,N_2525);
nand U3080 (N_3080,N_2952,N_2853);
and U3081 (N_3081,N_2995,N_2938);
nand U3082 (N_3082,N_2981,N_2765);
xnor U3083 (N_3083,N_2583,N_2649);
nand U3084 (N_3084,N_2823,N_2907);
or U3085 (N_3085,N_2718,N_2855);
xor U3086 (N_3086,N_2917,N_2804);
nor U3087 (N_3087,N_2944,N_2866);
nand U3088 (N_3088,N_2731,N_2604);
xnor U3089 (N_3089,N_2835,N_2816);
xor U3090 (N_3090,N_2575,N_2736);
or U3091 (N_3091,N_2597,N_2818);
nor U3092 (N_3092,N_2921,N_2663);
or U3093 (N_3093,N_2733,N_2599);
nor U3094 (N_3094,N_2592,N_2885);
and U3095 (N_3095,N_2837,N_2939);
or U3096 (N_3096,N_2969,N_2886);
or U3097 (N_3097,N_2918,N_2633);
or U3098 (N_3098,N_2735,N_2666);
and U3099 (N_3099,N_2593,N_2546);
and U3100 (N_3100,N_2636,N_2897);
and U3101 (N_3101,N_2674,N_2505);
nor U3102 (N_3102,N_2558,N_2585);
xnor U3103 (N_3103,N_2610,N_2687);
or U3104 (N_3104,N_2796,N_2562);
nor U3105 (N_3105,N_2624,N_2516);
and U3106 (N_3106,N_2964,N_2961);
nor U3107 (N_3107,N_2591,N_2646);
or U3108 (N_3108,N_2954,N_2507);
nor U3109 (N_3109,N_2865,N_2857);
nor U3110 (N_3110,N_2667,N_2701);
xor U3111 (N_3111,N_2703,N_2744);
xnor U3112 (N_3112,N_2955,N_2738);
or U3113 (N_3113,N_2774,N_2748);
or U3114 (N_3114,N_2717,N_2882);
nand U3115 (N_3115,N_2614,N_2887);
xor U3116 (N_3116,N_2859,N_2641);
and U3117 (N_3117,N_2559,N_2678);
nand U3118 (N_3118,N_2647,N_2732);
or U3119 (N_3119,N_2868,N_2607);
nand U3120 (N_3120,N_2776,N_2634);
xnor U3121 (N_3121,N_2673,N_2799);
or U3122 (N_3122,N_2842,N_2688);
and U3123 (N_3123,N_2638,N_2655);
nor U3124 (N_3124,N_2543,N_2779);
nor U3125 (N_3125,N_2803,N_2511);
or U3126 (N_3126,N_2983,N_2856);
nor U3127 (N_3127,N_2751,N_2512);
and U3128 (N_3128,N_2758,N_2960);
nand U3129 (N_3129,N_2791,N_2669);
xnor U3130 (N_3130,N_2694,N_2992);
nand U3131 (N_3131,N_2839,N_2645);
or U3132 (N_3132,N_2728,N_2709);
xnor U3133 (N_3133,N_2533,N_2783);
or U3134 (N_3134,N_2891,N_2953);
nand U3135 (N_3135,N_2724,N_2898);
nand U3136 (N_3136,N_2997,N_2696);
and U3137 (N_3137,N_2782,N_2769);
nand U3138 (N_3138,N_2549,N_2832);
nand U3139 (N_3139,N_2824,N_2531);
xor U3140 (N_3140,N_2587,N_2651);
or U3141 (N_3141,N_2695,N_2817);
or U3142 (N_3142,N_2869,N_2986);
nand U3143 (N_3143,N_2982,N_2812);
nor U3144 (N_3144,N_2503,N_2656);
xor U3145 (N_3145,N_2565,N_2567);
and U3146 (N_3146,N_2772,N_2761);
and U3147 (N_3147,N_2840,N_2556);
xor U3148 (N_3148,N_2520,N_2926);
and U3149 (N_3149,N_2571,N_2753);
nor U3150 (N_3150,N_2547,N_2664);
or U3151 (N_3151,N_2754,N_2993);
nor U3152 (N_3152,N_2612,N_2936);
xnor U3153 (N_3153,N_2705,N_2560);
xor U3154 (N_3154,N_2594,N_2586);
xnor U3155 (N_3155,N_2580,N_2756);
nor U3156 (N_3156,N_2589,N_2787);
xnor U3157 (N_3157,N_2830,N_2537);
or U3158 (N_3158,N_2706,N_2643);
or U3159 (N_3159,N_2908,N_2935);
nand U3160 (N_3160,N_2608,N_2978);
or U3161 (N_3161,N_2509,N_2639);
and U3162 (N_3162,N_2598,N_2544);
or U3163 (N_3163,N_2524,N_2627);
nand U3164 (N_3164,N_2683,N_2972);
nand U3165 (N_3165,N_2836,N_2915);
xnor U3166 (N_3166,N_2806,N_2699);
and U3167 (N_3167,N_2539,N_2541);
xnor U3168 (N_3168,N_2723,N_2844);
nor U3169 (N_3169,N_2697,N_2650);
and U3170 (N_3170,N_2809,N_2899);
or U3171 (N_3171,N_2875,N_2595);
nand U3172 (N_3172,N_2873,N_2956);
nor U3173 (N_3173,N_2554,N_2693);
nand U3174 (N_3174,N_2635,N_2889);
or U3175 (N_3175,N_2999,N_2825);
xnor U3176 (N_3176,N_2963,N_2976);
nand U3177 (N_3177,N_2813,N_2932);
and U3178 (N_3178,N_2712,N_2704);
and U3179 (N_3179,N_2629,N_2660);
and U3180 (N_3180,N_2725,N_2719);
or U3181 (N_3181,N_2985,N_2973);
nor U3182 (N_3182,N_2988,N_2902);
nand U3183 (N_3183,N_2553,N_2933);
nor U3184 (N_3184,N_2523,N_2934);
nand U3185 (N_3185,N_2517,N_2613);
nand U3186 (N_3186,N_2752,N_2529);
and U3187 (N_3187,N_2862,N_2990);
and U3188 (N_3188,N_2968,N_2942);
nor U3189 (N_3189,N_2714,N_2713);
nor U3190 (N_3190,N_2737,N_2996);
and U3191 (N_3191,N_2659,N_2922);
nand U3192 (N_3192,N_2722,N_2884);
and U3193 (N_3193,N_2581,N_2947);
and U3194 (N_3194,N_2500,N_2642);
or U3195 (N_3195,N_2989,N_2849);
nor U3196 (N_3196,N_2617,N_2711);
and U3197 (N_3197,N_2967,N_2528);
nor U3198 (N_3198,N_2763,N_2619);
or U3199 (N_3199,N_2863,N_2987);
and U3200 (N_3200,N_2786,N_2834);
nand U3201 (N_3201,N_2876,N_2757);
nor U3202 (N_3202,N_2822,N_2831);
or U3203 (N_3203,N_2727,N_2829);
nand U3204 (N_3204,N_2820,N_2540);
nand U3205 (N_3205,N_2513,N_2582);
nor U3206 (N_3206,N_2789,N_2974);
or U3207 (N_3207,N_2994,N_2879);
xnor U3208 (N_3208,N_2618,N_2912);
nand U3209 (N_3209,N_2749,N_2781);
nand U3210 (N_3210,N_2661,N_2957);
nand U3211 (N_3211,N_2977,N_2888);
or U3212 (N_3212,N_2940,N_2588);
xnor U3213 (N_3213,N_2916,N_2602);
nor U3214 (N_3214,N_2847,N_2798);
or U3215 (N_3215,N_2691,N_2959);
and U3216 (N_3216,N_2534,N_2746);
xor U3217 (N_3217,N_2715,N_2950);
or U3218 (N_3218,N_2971,N_2903);
and U3219 (N_3219,N_2652,N_2550);
and U3220 (N_3220,N_2930,N_2720);
and U3221 (N_3221,N_2552,N_2504);
xor U3222 (N_3222,N_2807,N_2570);
or U3223 (N_3223,N_2742,N_2657);
xnor U3224 (N_3224,N_2893,N_2745);
xor U3225 (N_3225,N_2601,N_2680);
and U3226 (N_3226,N_2665,N_2914);
xnor U3227 (N_3227,N_2828,N_2569);
xnor U3228 (N_3228,N_2894,N_2536);
nor U3229 (N_3229,N_2625,N_2979);
nand U3230 (N_3230,N_2690,N_2966);
nor U3231 (N_3231,N_2710,N_2785);
or U3232 (N_3232,N_2913,N_2616);
and U3233 (N_3233,N_2538,N_2630);
and U3234 (N_3234,N_2943,N_2768);
and U3235 (N_3235,N_2920,N_2561);
and U3236 (N_3236,N_2874,N_2579);
nand U3237 (N_3237,N_2790,N_2750);
and U3238 (N_3238,N_2766,N_2606);
xnor U3239 (N_3239,N_2708,N_2854);
xor U3240 (N_3240,N_2991,N_2682);
nand U3241 (N_3241,N_2780,N_2861);
xor U3242 (N_3242,N_2620,N_2904);
and U3243 (N_3243,N_2833,N_2860);
nor U3244 (N_3244,N_2535,N_2946);
or U3245 (N_3245,N_2814,N_2662);
xnor U3246 (N_3246,N_2945,N_2518);
xor U3247 (N_3247,N_2730,N_2901);
nor U3248 (N_3248,N_2811,N_2910);
nand U3249 (N_3249,N_2555,N_2927);
nor U3250 (N_3250,N_2871,N_2679);
xor U3251 (N_3251,N_2827,N_2934);
nor U3252 (N_3252,N_2538,N_2615);
or U3253 (N_3253,N_2783,N_2992);
and U3254 (N_3254,N_2806,N_2554);
and U3255 (N_3255,N_2733,N_2641);
and U3256 (N_3256,N_2568,N_2648);
or U3257 (N_3257,N_2848,N_2884);
nor U3258 (N_3258,N_2511,N_2590);
nor U3259 (N_3259,N_2642,N_2847);
nand U3260 (N_3260,N_2732,N_2661);
xnor U3261 (N_3261,N_2595,N_2685);
nand U3262 (N_3262,N_2711,N_2873);
nand U3263 (N_3263,N_2820,N_2970);
xor U3264 (N_3264,N_2879,N_2633);
and U3265 (N_3265,N_2756,N_2616);
xnor U3266 (N_3266,N_2697,N_2657);
xor U3267 (N_3267,N_2851,N_2926);
nand U3268 (N_3268,N_2962,N_2528);
xnor U3269 (N_3269,N_2521,N_2678);
xnor U3270 (N_3270,N_2875,N_2659);
or U3271 (N_3271,N_2838,N_2697);
nand U3272 (N_3272,N_2552,N_2717);
nor U3273 (N_3273,N_2867,N_2675);
nor U3274 (N_3274,N_2713,N_2536);
xor U3275 (N_3275,N_2667,N_2914);
or U3276 (N_3276,N_2908,N_2730);
nor U3277 (N_3277,N_2957,N_2950);
nand U3278 (N_3278,N_2525,N_2750);
or U3279 (N_3279,N_2626,N_2950);
and U3280 (N_3280,N_2975,N_2724);
xnor U3281 (N_3281,N_2888,N_2970);
or U3282 (N_3282,N_2584,N_2759);
and U3283 (N_3283,N_2884,N_2606);
nor U3284 (N_3284,N_2922,N_2889);
nor U3285 (N_3285,N_2751,N_2839);
nor U3286 (N_3286,N_2808,N_2587);
nor U3287 (N_3287,N_2541,N_2892);
and U3288 (N_3288,N_2632,N_2790);
nor U3289 (N_3289,N_2729,N_2633);
or U3290 (N_3290,N_2833,N_2645);
or U3291 (N_3291,N_2966,N_2581);
and U3292 (N_3292,N_2559,N_2725);
xor U3293 (N_3293,N_2626,N_2819);
or U3294 (N_3294,N_2814,N_2661);
and U3295 (N_3295,N_2708,N_2552);
or U3296 (N_3296,N_2903,N_2734);
or U3297 (N_3297,N_2869,N_2711);
or U3298 (N_3298,N_2895,N_2643);
nand U3299 (N_3299,N_2633,N_2663);
nand U3300 (N_3300,N_2874,N_2633);
nor U3301 (N_3301,N_2711,N_2915);
or U3302 (N_3302,N_2634,N_2717);
and U3303 (N_3303,N_2887,N_2575);
or U3304 (N_3304,N_2649,N_2910);
or U3305 (N_3305,N_2902,N_2592);
xnor U3306 (N_3306,N_2881,N_2909);
nand U3307 (N_3307,N_2617,N_2972);
or U3308 (N_3308,N_2569,N_2837);
or U3309 (N_3309,N_2736,N_2690);
xor U3310 (N_3310,N_2589,N_2754);
xor U3311 (N_3311,N_2590,N_2916);
xor U3312 (N_3312,N_2525,N_2813);
xor U3313 (N_3313,N_2903,N_2755);
xor U3314 (N_3314,N_2700,N_2896);
nand U3315 (N_3315,N_2624,N_2904);
xnor U3316 (N_3316,N_2650,N_2796);
xnor U3317 (N_3317,N_2791,N_2604);
nand U3318 (N_3318,N_2773,N_2895);
nand U3319 (N_3319,N_2754,N_2842);
and U3320 (N_3320,N_2971,N_2564);
nand U3321 (N_3321,N_2517,N_2806);
nand U3322 (N_3322,N_2629,N_2814);
or U3323 (N_3323,N_2572,N_2697);
and U3324 (N_3324,N_2742,N_2551);
nor U3325 (N_3325,N_2757,N_2966);
nand U3326 (N_3326,N_2623,N_2804);
or U3327 (N_3327,N_2682,N_2578);
nand U3328 (N_3328,N_2999,N_2788);
and U3329 (N_3329,N_2679,N_2501);
and U3330 (N_3330,N_2919,N_2584);
and U3331 (N_3331,N_2652,N_2647);
xor U3332 (N_3332,N_2947,N_2807);
nor U3333 (N_3333,N_2582,N_2520);
nand U3334 (N_3334,N_2899,N_2612);
xnor U3335 (N_3335,N_2654,N_2739);
or U3336 (N_3336,N_2915,N_2569);
or U3337 (N_3337,N_2960,N_2855);
nand U3338 (N_3338,N_2819,N_2827);
nand U3339 (N_3339,N_2885,N_2636);
or U3340 (N_3340,N_2996,N_2766);
or U3341 (N_3341,N_2910,N_2834);
or U3342 (N_3342,N_2550,N_2692);
or U3343 (N_3343,N_2920,N_2725);
nand U3344 (N_3344,N_2539,N_2929);
and U3345 (N_3345,N_2966,N_2875);
xnor U3346 (N_3346,N_2683,N_2768);
or U3347 (N_3347,N_2701,N_2688);
and U3348 (N_3348,N_2873,N_2742);
nand U3349 (N_3349,N_2914,N_2759);
nand U3350 (N_3350,N_2971,N_2511);
xnor U3351 (N_3351,N_2526,N_2673);
or U3352 (N_3352,N_2929,N_2841);
or U3353 (N_3353,N_2900,N_2980);
and U3354 (N_3354,N_2550,N_2852);
and U3355 (N_3355,N_2843,N_2933);
or U3356 (N_3356,N_2898,N_2989);
or U3357 (N_3357,N_2983,N_2512);
and U3358 (N_3358,N_2672,N_2517);
nor U3359 (N_3359,N_2696,N_2740);
nand U3360 (N_3360,N_2543,N_2724);
and U3361 (N_3361,N_2653,N_2578);
xor U3362 (N_3362,N_2785,N_2563);
or U3363 (N_3363,N_2574,N_2628);
xor U3364 (N_3364,N_2616,N_2579);
nand U3365 (N_3365,N_2596,N_2917);
or U3366 (N_3366,N_2725,N_2894);
and U3367 (N_3367,N_2757,N_2735);
and U3368 (N_3368,N_2825,N_2703);
nor U3369 (N_3369,N_2891,N_2669);
and U3370 (N_3370,N_2899,N_2594);
nor U3371 (N_3371,N_2970,N_2532);
xnor U3372 (N_3372,N_2804,N_2863);
xnor U3373 (N_3373,N_2564,N_2809);
or U3374 (N_3374,N_2755,N_2632);
and U3375 (N_3375,N_2917,N_2800);
and U3376 (N_3376,N_2972,N_2616);
nand U3377 (N_3377,N_2753,N_2576);
nor U3378 (N_3378,N_2662,N_2987);
xor U3379 (N_3379,N_2939,N_2524);
xnor U3380 (N_3380,N_2670,N_2806);
xnor U3381 (N_3381,N_2982,N_2770);
nand U3382 (N_3382,N_2564,N_2577);
nand U3383 (N_3383,N_2637,N_2896);
and U3384 (N_3384,N_2829,N_2956);
nand U3385 (N_3385,N_2505,N_2812);
and U3386 (N_3386,N_2536,N_2580);
xor U3387 (N_3387,N_2691,N_2562);
or U3388 (N_3388,N_2528,N_2561);
nor U3389 (N_3389,N_2552,N_2596);
nor U3390 (N_3390,N_2986,N_2826);
xor U3391 (N_3391,N_2961,N_2552);
or U3392 (N_3392,N_2571,N_2952);
nor U3393 (N_3393,N_2992,N_2881);
nor U3394 (N_3394,N_2904,N_2830);
nand U3395 (N_3395,N_2536,N_2729);
nand U3396 (N_3396,N_2703,N_2913);
xnor U3397 (N_3397,N_2609,N_2922);
xnor U3398 (N_3398,N_2760,N_2660);
xnor U3399 (N_3399,N_2708,N_2802);
xor U3400 (N_3400,N_2838,N_2964);
or U3401 (N_3401,N_2651,N_2552);
and U3402 (N_3402,N_2626,N_2549);
nor U3403 (N_3403,N_2820,N_2685);
or U3404 (N_3404,N_2925,N_2886);
nor U3405 (N_3405,N_2544,N_2532);
or U3406 (N_3406,N_2906,N_2915);
or U3407 (N_3407,N_2504,N_2654);
xnor U3408 (N_3408,N_2972,N_2819);
xor U3409 (N_3409,N_2685,N_2580);
or U3410 (N_3410,N_2757,N_2514);
nor U3411 (N_3411,N_2630,N_2595);
xnor U3412 (N_3412,N_2929,N_2815);
and U3413 (N_3413,N_2966,N_2958);
nand U3414 (N_3414,N_2675,N_2896);
or U3415 (N_3415,N_2835,N_2737);
nand U3416 (N_3416,N_2538,N_2812);
xnor U3417 (N_3417,N_2677,N_2913);
or U3418 (N_3418,N_2504,N_2749);
xnor U3419 (N_3419,N_2501,N_2662);
nand U3420 (N_3420,N_2757,N_2516);
and U3421 (N_3421,N_2822,N_2626);
xnor U3422 (N_3422,N_2847,N_2933);
nand U3423 (N_3423,N_2872,N_2544);
or U3424 (N_3424,N_2651,N_2515);
or U3425 (N_3425,N_2666,N_2971);
and U3426 (N_3426,N_2575,N_2951);
nand U3427 (N_3427,N_2744,N_2931);
nand U3428 (N_3428,N_2638,N_2692);
nand U3429 (N_3429,N_2777,N_2971);
nand U3430 (N_3430,N_2516,N_2771);
and U3431 (N_3431,N_2613,N_2967);
nor U3432 (N_3432,N_2601,N_2878);
xnor U3433 (N_3433,N_2608,N_2700);
or U3434 (N_3434,N_2744,N_2692);
or U3435 (N_3435,N_2617,N_2672);
nand U3436 (N_3436,N_2967,N_2649);
nor U3437 (N_3437,N_2778,N_2886);
or U3438 (N_3438,N_2569,N_2939);
and U3439 (N_3439,N_2609,N_2711);
and U3440 (N_3440,N_2975,N_2515);
nor U3441 (N_3441,N_2995,N_2894);
nand U3442 (N_3442,N_2538,N_2566);
or U3443 (N_3443,N_2917,N_2953);
nand U3444 (N_3444,N_2580,N_2732);
nand U3445 (N_3445,N_2853,N_2504);
or U3446 (N_3446,N_2995,N_2627);
and U3447 (N_3447,N_2959,N_2542);
nand U3448 (N_3448,N_2590,N_2996);
or U3449 (N_3449,N_2912,N_2595);
or U3450 (N_3450,N_2712,N_2763);
and U3451 (N_3451,N_2848,N_2946);
nor U3452 (N_3452,N_2610,N_2606);
xor U3453 (N_3453,N_2575,N_2612);
nand U3454 (N_3454,N_2749,N_2983);
or U3455 (N_3455,N_2894,N_2643);
and U3456 (N_3456,N_2512,N_2793);
nor U3457 (N_3457,N_2525,N_2665);
nor U3458 (N_3458,N_2511,N_2535);
nor U3459 (N_3459,N_2954,N_2696);
xor U3460 (N_3460,N_2614,N_2556);
xor U3461 (N_3461,N_2532,N_2573);
nand U3462 (N_3462,N_2889,N_2582);
nor U3463 (N_3463,N_2532,N_2502);
nor U3464 (N_3464,N_2589,N_2894);
xor U3465 (N_3465,N_2717,N_2807);
xnor U3466 (N_3466,N_2824,N_2562);
nand U3467 (N_3467,N_2969,N_2830);
and U3468 (N_3468,N_2686,N_2666);
and U3469 (N_3469,N_2584,N_2666);
xnor U3470 (N_3470,N_2517,N_2906);
nor U3471 (N_3471,N_2852,N_2672);
or U3472 (N_3472,N_2783,N_2718);
or U3473 (N_3473,N_2647,N_2963);
or U3474 (N_3474,N_2631,N_2911);
nand U3475 (N_3475,N_2964,N_2560);
xor U3476 (N_3476,N_2946,N_2669);
or U3477 (N_3477,N_2578,N_2620);
nor U3478 (N_3478,N_2805,N_2932);
xnor U3479 (N_3479,N_2933,N_2613);
nor U3480 (N_3480,N_2973,N_2796);
or U3481 (N_3481,N_2845,N_2964);
or U3482 (N_3482,N_2895,N_2738);
xor U3483 (N_3483,N_2531,N_2584);
or U3484 (N_3484,N_2654,N_2991);
xnor U3485 (N_3485,N_2691,N_2988);
nand U3486 (N_3486,N_2930,N_2683);
or U3487 (N_3487,N_2850,N_2662);
or U3488 (N_3488,N_2580,N_2968);
nand U3489 (N_3489,N_2997,N_2857);
nand U3490 (N_3490,N_2815,N_2961);
xor U3491 (N_3491,N_2782,N_2791);
or U3492 (N_3492,N_2913,N_2570);
nand U3493 (N_3493,N_2954,N_2866);
xnor U3494 (N_3494,N_2863,N_2962);
nand U3495 (N_3495,N_2776,N_2961);
nor U3496 (N_3496,N_2880,N_2726);
nor U3497 (N_3497,N_2721,N_2870);
or U3498 (N_3498,N_2774,N_2961);
or U3499 (N_3499,N_2720,N_2689);
or U3500 (N_3500,N_3477,N_3443);
nand U3501 (N_3501,N_3160,N_3356);
or U3502 (N_3502,N_3372,N_3458);
nand U3503 (N_3503,N_3236,N_3272);
nor U3504 (N_3504,N_3471,N_3310);
or U3505 (N_3505,N_3419,N_3393);
or U3506 (N_3506,N_3429,N_3385);
xor U3507 (N_3507,N_3162,N_3407);
and U3508 (N_3508,N_3350,N_3432);
and U3509 (N_3509,N_3357,N_3193);
xor U3510 (N_3510,N_3247,N_3460);
nand U3511 (N_3511,N_3260,N_3007);
and U3512 (N_3512,N_3353,N_3103);
nand U3513 (N_3513,N_3342,N_3220);
nand U3514 (N_3514,N_3448,N_3205);
and U3515 (N_3515,N_3416,N_3055);
nor U3516 (N_3516,N_3031,N_3254);
nor U3517 (N_3517,N_3309,N_3163);
nor U3518 (N_3518,N_3312,N_3324);
xor U3519 (N_3519,N_3266,N_3206);
nand U3520 (N_3520,N_3200,N_3225);
xor U3521 (N_3521,N_3013,N_3437);
xor U3522 (N_3522,N_3280,N_3070);
nor U3523 (N_3523,N_3188,N_3177);
xnor U3524 (N_3524,N_3131,N_3089);
and U3525 (N_3525,N_3119,N_3445);
xor U3526 (N_3526,N_3190,N_3010);
nor U3527 (N_3527,N_3008,N_3347);
and U3528 (N_3528,N_3164,N_3112);
and U3529 (N_3529,N_3168,N_3198);
nand U3530 (N_3530,N_3343,N_3078);
nor U3531 (N_3531,N_3191,N_3136);
nor U3532 (N_3532,N_3498,N_3242);
xnor U3533 (N_3533,N_3151,N_3394);
nor U3534 (N_3534,N_3386,N_3492);
nor U3535 (N_3535,N_3082,N_3387);
xnor U3536 (N_3536,N_3406,N_3428);
nand U3537 (N_3537,N_3380,N_3287);
xor U3538 (N_3538,N_3130,N_3487);
nand U3539 (N_3539,N_3115,N_3041);
nand U3540 (N_3540,N_3421,N_3039);
nor U3541 (N_3541,N_3321,N_3173);
nor U3542 (N_3542,N_3392,N_3391);
and U3543 (N_3543,N_3100,N_3431);
or U3544 (N_3544,N_3472,N_3358);
nor U3545 (N_3545,N_3124,N_3488);
xor U3546 (N_3546,N_3439,N_3384);
xor U3547 (N_3547,N_3122,N_3085);
or U3548 (N_3548,N_3355,N_3269);
nor U3549 (N_3549,N_3117,N_3049);
and U3550 (N_3550,N_3113,N_3067);
or U3551 (N_3551,N_3019,N_3025);
and U3552 (N_3552,N_3189,N_3241);
and U3553 (N_3553,N_3228,N_3064);
or U3554 (N_3554,N_3376,N_3468);
or U3555 (N_3555,N_3106,N_3073);
nor U3556 (N_3556,N_3230,N_3395);
nor U3557 (N_3557,N_3268,N_3054);
nand U3558 (N_3558,N_3011,N_3056);
xnor U3559 (N_3559,N_3261,N_3462);
and U3560 (N_3560,N_3370,N_3301);
and U3561 (N_3561,N_3479,N_3227);
or U3562 (N_3562,N_3390,N_3375);
or U3563 (N_3563,N_3118,N_3022);
nor U3564 (N_3564,N_3265,N_3399);
xor U3565 (N_3565,N_3036,N_3090);
xor U3566 (N_3566,N_3340,N_3322);
nand U3567 (N_3567,N_3108,N_3238);
nand U3568 (N_3568,N_3410,N_3181);
or U3569 (N_3569,N_3137,N_3121);
nor U3570 (N_3570,N_3361,N_3180);
nor U3571 (N_3571,N_3330,N_3065);
or U3572 (N_3572,N_3497,N_3296);
nand U3573 (N_3573,N_3223,N_3434);
xor U3574 (N_3574,N_3305,N_3478);
nand U3575 (N_3575,N_3414,N_3125);
and U3576 (N_3576,N_3377,N_3438);
xnor U3577 (N_3577,N_3367,N_3217);
nand U3578 (N_3578,N_3048,N_3229);
nor U3579 (N_3579,N_3159,N_3405);
nand U3580 (N_3580,N_3222,N_3398);
xnor U3581 (N_3581,N_3291,N_3294);
nand U3582 (N_3582,N_3126,N_3298);
and U3583 (N_3583,N_3249,N_3026);
and U3584 (N_3584,N_3476,N_3303);
or U3585 (N_3585,N_3133,N_3311);
or U3586 (N_3586,N_3493,N_3182);
and U3587 (N_3587,N_3021,N_3156);
nand U3588 (N_3588,N_3032,N_3359);
nand U3589 (N_3589,N_3446,N_3210);
or U3590 (N_3590,N_3145,N_3084);
and U3591 (N_3591,N_3491,N_3232);
xnor U3592 (N_3592,N_3346,N_3231);
or U3593 (N_3593,N_3326,N_3494);
or U3594 (N_3594,N_3283,N_3299);
or U3595 (N_3595,N_3216,N_3235);
or U3596 (N_3596,N_3348,N_3344);
xnor U3597 (N_3597,N_3104,N_3331);
xnor U3598 (N_3598,N_3307,N_3098);
nand U3599 (N_3599,N_3071,N_3009);
xor U3600 (N_3600,N_3282,N_3378);
nand U3601 (N_3601,N_3316,N_3127);
and U3602 (N_3602,N_3092,N_3207);
nand U3603 (N_3603,N_3051,N_3132);
nor U3604 (N_3604,N_3218,N_3139);
nor U3605 (N_3605,N_3044,N_3338);
and U3606 (N_3606,N_3456,N_3172);
nor U3607 (N_3607,N_3194,N_3475);
xnor U3608 (N_3608,N_3000,N_3457);
nand U3609 (N_3609,N_3363,N_3034);
xor U3610 (N_3610,N_3074,N_3178);
xnor U3611 (N_3611,N_3058,N_3485);
and U3612 (N_3612,N_3063,N_3224);
and U3613 (N_3613,N_3110,N_3273);
or U3614 (N_3614,N_3369,N_3441);
or U3615 (N_3615,N_3470,N_3183);
xnor U3616 (N_3616,N_3023,N_3080);
or U3617 (N_3617,N_3114,N_3455);
nand U3618 (N_3618,N_3374,N_3215);
xor U3619 (N_3619,N_3461,N_3449);
nor U3620 (N_3620,N_3246,N_3204);
nor U3621 (N_3621,N_3454,N_3081);
nand U3622 (N_3622,N_3364,N_3105);
or U3623 (N_3623,N_3295,N_3373);
nand U3624 (N_3624,N_3499,N_3417);
nand U3625 (N_3625,N_3027,N_3033);
nand U3626 (N_3626,N_3086,N_3288);
nand U3627 (N_3627,N_3195,N_3286);
nand U3628 (N_3628,N_3404,N_3111);
nand U3629 (N_3629,N_3016,N_3142);
xnor U3630 (N_3630,N_3425,N_3256);
nand U3631 (N_3631,N_3057,N_3275);
xor U3632 (N_3632,N_3144,N_3362);
xor U3633 (N_3633,N_3382,N_3379);
and U3634 (N_3634,N_3094,N_3096);
or U3635 (N_3635,N_3042,N_3465);
and U3636 (N_3636,N_3097,N_3134);
nor U3637 (N_3637,N_3109,N_3459);
or U3638 (N_3638,N_3069,N_3251);
nor U3639 (N_3639,N_3239,N_3244);
nor U3640 (N_3640,N_3495,N_3199);
and U3641 (N_3641,N_3452,N_3253);
or U3642 (N_3642,N_3252,N_3187);
xnor U3643 (N_3643,N_3146,N_3066);
nand U3644 (N_3644,N_3444,N_3167);
or U3645 (N_3645,N_3175,N_3046);
or U3646 (N_3646,N_3334,N_3150);
or U3647 (N_3647,N_3208,N_3371);
and U3648 (N_3648,N_3061,N_3018);
or U3649 (N_3649,N_3352,N_3262);
or U3650 (N_3650,N_3473,N_3427);
or U3651 (N_3651,N_3388,N_3169);
xor U3652 (N_3652,N_3052,N_3480);
or U3653 (N_3653,N_3165,N_3481);
nand U3654 (N_3654,N_3004,N_3209);
or U3655 (N_3655,N_3001,N_3091);
nand U3656 (N_3656,N_3258,N_3102);
nor U3657 (N_3657,N_3381,N_3426);
or U3658 (N_3658,N_3333,N_3463);
and U3659 (N_3659,N_3420,N_3143);
nor U3660 (N_3660,N_3368,N_3400);
or U3661 (N_3661,N_3196,N_3323);
nor U3662 (N_3662,N_3289,N_3171);
nand U3663 (N_3663,N_3327,N_3176);
xor U3664 (N_3664,N_3453,N_3469);
and U3665 (N_3665,N_3413,N_3147);
xor U3666 (N_3666,N_3430,N_3270);
nand U3667 (N_3667,N_3271,N_3237);
nand U3668 (N_3668,N_3318,N_3332);
nor U3669 (N_3669,N_3401,N_3138);
and U3670 (N_3670,N_3213,N_3128);
and U3671 (N_3671,N_3093,N_3116);
nor U3672 (N_3672,N_3255,N_3366);
nor U3673 (N_3673,N_3408,N_3202);
nand U3674 (N_3674,N_3319,N_3192);
xor U3675 (N_3675,N_3135,N_3038);
and U3676 (N_3676,N_3012,N_3313);
and U3677 (N_3677,N_3467,N_3141);
xnor U3678 (N_3678,N_3450,N_3047);
xor U3679 (N_3679,N_3075,N_3412);
and U3680 (N_3680,N_3101,N_3014);
and U3681 (N_3681,N_3197,N_3440);
and U3682 (N_3682,N_3297,N_3274);
and U3683 (N_3683,N_3257,N_3120);
or U3684 (N_3684,N_3099,N_3259);
and U3685 (N_3685,N_3422,N_3017);
xnor U3686 (N_3686,N_3403,N_3402);
xnor U3687 (N_3687,N_3474,N_3464);
nor U3688 (N_3688,N_3015,N_3030);
xor U3689 (N_3689,N_3140,N_3335);
xnor U3690 (N_3690,N_3293,N_3050);
nor U3691 (N_3691,N_3281,N_3077);
nand U3692 (N_3692,N_3020,N_3170);
nor U3693 (N_3693,N_3029,N_3002);
xnor U3694 (N_3694,N_3317,N_3129);
and U3695 (N_3695,N_3415,N_3447);
and U3696 (N_3696,N_3214,N_3221);
nor U3697 (N_3697,N_3186,N_3088);
nor U3698 (N_3698,N_3157,N_3442);
or U3699 (N_3699,N_3148,N_3300);
nor U3700 (N_3700,N_3423,N_3240);
xnor U3701 (N_3701,N_3284,N_3212);
or U3702 (N_3702,N_3005,N_3158);
nand U3703 (N_3703,N_3277,N_3152);
or U3704 (N_3704,N_3234,N_3336);
or U3705 (N_3705,N_3435,N_3349);
xor U3706 (N_3706,N_3339,N_3486);
and U3707 (N_3707,N_3045,N_3483);
nand U3708 (N_3708,N_3087,N_3325);
and U3709 (N_3709,N_3360,N_3490);
or U3710 (N_3710,N_3006,N_3062);
and U3711 (N_3711,N_3482,N_3060);
nand U3712 (N_3712,N_3059,N_3418);
or U3713 (N_3713,N_3351,N_3396);
and U3714 (N_3714,N_3226,N_3466);
nor U3715 (N_3715,N_3365,N_3329);
nor U3716 (N_3716,N_3345,N_3174);
and U3717 (N_3717,N_3245,N_3267);
xor U3718 (N_3718,N_3161,N_3233);
nor U3719 (N_3719,N_3451,N_3328);
xor U3720 (N_3720,N_3436,N_3276);
xor U3721 (N_3721,N_3278,N_3028);
and U3722 (N_3722,N_3389,N_3264);
or U3723 (N_3723,N_3083,N_3149);
or U3724 (N_3724,N_3076,N_3079);
or U3725 (N_3725,N_3219,N_3304);
nor U3726 (N_3726,N_3107,N_3496);
nor U3727 (N_3727,N_3433,N_3040);
or U3728 (N_3728,N_3341,N_3153);
xor U3729 (N_3729,N_3397,N_3354);
xnor U3730 (N_3730,N_3279,N_3285);
nand U3731 (N_3731,N_3292,N_3489);
xor U3732 (N_3732,N_3184,N_3053);
nor U3733 (N_3733,N_3072,N_3383);
nor U3734 (N_3734,N_3263,N_3320);
nand U3735 (N_3735,N_3248,N_3250);
and U3736 (N_3736,N_3179,N_3155);
and U3737 (N_3737,N_3003,N_3203);
or U3738 (N_3738,N_3095,N_3035);
and U3739 (N_3739,N_3243,N_3201);
nand U3740 (N_3740,N_3306,N_3308);
and U3741 (N_3741,N_3154,N_3409);
and U3742 (N_3742,N_3211,N_3424);
nand U3743 (N_3743,N_3037,N_3411);
nand U3744 (N_3744,N_3290,N_3185);
xor U3745 (N_3745,N_3315,N_3024);
xor U3746 (N_3746,N_3068,N_3166);
or U3747 (N_3747,N_3123,N_3484);
or U3748 (N_3748,N_3314,N_3043);
or U3749 (N_3749,N_3337,N_3302);
or U3750 (N_3750,N_3105,N_3246);
or U3751 (N_3751,N_3011,N_3127);
xor U3752 (N_3752,N_3000,N_3409);
nor U3753 (N_3753,N_3451,N_3274);
nor U3754 (N_3754,N_3473,N_3178);
and U3755 (N_3755,N_3014,N_3369);
nand U3756 (N_3756,N_3102,N_3171);
xor U3757 (N_3757,N_3393,N_3355);
nor U3758 (N_3758,N_3327,N_3031);
xnor U3759 (N_3759,N_3260,N_3028);
or U3760 (N_3760,N_3436,N_3298);
xor U3761 (N_3761,N_3213,N_3071);
and U3762 (N_3762,N_3014,N_3226);
and U3763 (N_3763,N_3209,N_3128);
nor U3764 (N_3764,N_3157,N_3056);
xnor U3765 (N_3765,N_3255,N_3437);
nand U3766 (N_3766,N_3378,N_3206);
or U3767 (N_3767,N_3076,N_3350);
and U3768 (N_3768,N_3077,N_3037);
or U3769 (N_3769,N_3424,N_3047);
and U3770 (N_3770,N_3477,N_3029);
nand U3771 (N_3771,N_3009,N_3088);
xnor U3772 (N_3772,N_3303,N_3178);
xor U3773 (N_3773,N_3259,N_3429);
nand U3774 (N_3774,N_3094,N_3035);
nor U3775 (N_3775,N_3408,N_3231);
nand U3776 (N_3776,N_3158,N_3227);
and U3777 (N_3777,N_3125,N_3020);
xnor U3778 (N_3778,N_3298,N_3369);
xnor U3779 (N_3779,N_3094,N_3496);
or U3780 (N_3780,N_3495,N_3179);
xnor U3781 (N_3781,N_3460,N_3363);
nor U3782 (N_3782,N_3020,N_3244);
xnor U3783 (N_3783,N_3497,N_3272);
and U3784 (N_3784,N_3414,N_3458);
xnor U3785 (N_3785,N_3058,N_3332);
and U3786 (N_3786,N_3183,N_3494);
nor U3787 (N_3787,N_3234,N_3128);
xor U3788 (N_3788,N_3296,N_3247);
or U3789 (N_3789,N_3306,N_3469);
nor U3790 (N_3790,N_3465,N_3252);
xnor U3791 (N_3791,N_3041,N_3292);
xor U3792 (N_3792,N_3482,N_3492);
or U3793 (N_3793,N_3265,N_3299);
and U3794 (N_3794,N_3262,N_3253);
nand U3795 (N_3795,N_3092,N_3168);
xnor U3796 (N_3796,N_3088,N_3052);
nor U3797 (N_3797,N_3009,N_3029);
nand U3798 (N_3798,N_3165,N_3352);
nor U3799 (N_3799,N_3217,N_3417);
xor U3800 (N_3800,N_3305,N_3254);
xor U3801 (N_3801,N_3294,N_3238);
or U3802 (N_3802,N_3439,N_3378);
or U3803 (N_3803,N_3332,N_3352);
or U3804 (N_3804,N_3225,N_3282);
nor U3805 (N_3805,N_3432,N_3335);
xor U3806 (N_3806,N_3479,N_3313);
and U3807 (N_3807,N_3370,N_3351);
and U3808 (N_3808,N_3184,N_3050);
nand U3809 (N_3809,N_3455,N_3088);
or U3810 (N_3810,N_3000,N_3125);
and U3811 (N_3811,N_3045,N_3323);
and U3812 (N_3812,N_3066,N_3455);
nor U3813 (N_3813,N_3185,N_3227);
or U3814 (N_3814,N_3261,N_3440);
nor U3815 (N_3815,N_3040,N_3188);
or U3816 (N_3816,N_3124,N_3308);
nand U3817 (N_3817,N_3365,N_3243);
xor U3818 (N_3818,N_3223,N_3440);
xor U3819 (N_3819,N_3246,N_3134);
and U3820 (N_3820,N_3433,N_3110);
and U3821 (N_3821,N_3117,N_3400);
and U3822 (N_3822,N_3315,N_3475);
and U3823 (N_3823,N_3007,N_3449);
and U3824 (N_3824,N_3002,N_3430);
xor U3825 (N_3825,N_3276,N_3069);
or U3826 (N_3826,N_3169,N_3156);
nor U3827 (N_3827,N_3301,N_3132);
xnor U3828 (N_3828,N_3179,N_3234);
and U3829 (N_3829,N_3238,N_3385);
and U3830 (N_3830,N_3475,N_3135);
nor U3831 (N_3831,N_3036,N_3278);
or U3832 (N_3832,N_3115,N_3409);
and U3833 (N_3833,N_3283,N_3215);
nand U3834 (N_3834,N_3249,N_3138);
nand U3835 (N_3835,N_3440,N_3462);
nand U3836 (N_3836,N_3320,N_3005);
xnor U3837 (N_3837,N_3359,N_3175);
and U3838 (N_3838,N_3391,N_3323);
nor U3839 (N_3839,N_3204,N_3095);
and U3840 (N_3840,N_3477,N_3333);
xnor U3841 (N_3841,N_3195,N_3173);
nand U3842 (N_3842,N_3413,N_3044);
nand U3843 (N_3843,N_3288,N_3108);
or U3844 (N_3844,N_3347,N_3057);
nor U3845 (N_3845,N_3146,N_3194);
or U3846 (N_3846,N_3054,N_3480);
xor U3847 (N_3847,N_3399,N_3154);
or U3848 (N_3848,N_3366,N_3351);
or U3849 (N_3849,N_3003,N_3009);
xnor U3850 (N_3850,N_3299,N_3244);
nand U3851 (N_3851,N_3084,N_3094);
or U3852 (N_3852,N_3436,N_3193);
xnor U3853 (N_3853,N_3423,N_3402);
nand U3854 (N_3854,N_3143,N_3433);
or U3855 (N_3855,N_3432,N_3158);
xor U3856 (N_3856,N_3207,N_3366);
xnor U3857 (N_3857,N_3148,N_3449);
or U3858 (N_3858,N_3277,N_3385);
and U3859 (N_3859,N_3340,N_3047);
nand U3860 (N_3860,N_3098,N_3488);
xnor U3861 (N_3861,N_3146,N_3328);
and U3862 (N_3862,N_3448,N_3423);
or U3863 (N_3863,N_3320,N_3211);
and U3864 (N_3864,N_3243,N_3040);
nor U3865 (N_3865,N_3041,N_3395);
nor U3866 (N_3866,N_3031,N_3378);
nor U3867 (N_3867,N_3006,N_3242);
nand U3868 (N_3868,N_3276,N_3349);
nand U3869 (N_3869,N_3440,N_3148);
and U3870 (N_3870,N_3247,N_3031);
nor U3871 (N_3871,N_3181,N_3309);
and U3872 (N_3872,N_3114,N_3382);
nor U3873 (N_3873,N_3065,N_3419);
nor U3874 (N_3874,N_3066,N_3268);
and U3875 (N_3875,N_3241,N_3494);
nand U3876 (N_3876,N_3025,N_3345);
nor U3877 (N_3877,N_3392,N_3266);
or U3878 (N_3878,N_3204,N_3403);
nor U3879 (N_3879,N_3134,N_3092);
nand U3880 (N_3880,N_3139,N_3266);
nand U3881 (N_3881,N_3080,N_3481);
or U3882 (N_3882,N_3067,N_3348);
nand U3883 (N_3883,N_3096,N_3437);
and U3884 (N_3884,N_3102,N_3337);
xor U3885 (N_3885,N_3183,N_3449);
nor U3886 (N_3886,N_3035,N_3184);
nor U3887 (N_3887,N_3169,N_3180);
or U3888 (N_3888,N_3355,N_3061);
nor U3889 (N_3889,N_3111,N_3105);
or U3890 (N_3890,N_3453,N_3042);
xnor U3891 (N_3891,N_3170,N_3246);
nand U3892 (N_3892,N_3490,N_3233);
xor U3893 (N_3893,N_3063,N_3412);
nor U3894 (N_3894,N_3057,N_3272);
and U3895 (N_3895,N_3200,N_3094);
nor U3896 (N_3896,N_3018,N_3177);
xnor U3897 (N_3897,N_3041,N_3003);
nor U3898 (N_3898,N_3492,N_3120);
nand U3899 (N_3899,N_3348,N_3414);
or U3900 (N_3900,N_3429,N_3267);
or U3901 (N_3901,N_3251,N_3303);
and U3902 (N_3902,N_3222,N_3063);
and U3903 (N_3903,N_3330,N_3293);
xnor U3904 (N_3904,N_3133,N_3204);
or U3905 (N_3905,N_3379,N_3024);
nor U3906 (N_3906,N_3139,N_3147);
and U3907 (N_3907,N_3365,N_3103);
xor U3908 (N_3908,N_3077,N_3421);
nor U3909 (N_3909,N_3202,N_3104);
nand U3910 (N_3910,N_3109,N_3198);
or U3911 (N_3911,N_3145,N_3263);
xnor U3912 (N_3912,N_3183,N_3369);
xnor U3913 (N_3913,N_3442,N_3028);
nor U3914 (N_3914,N_3357,N_3095);
and U3915 (N_3915,N_3212,N_3151);
and U3916 (N_3916,N_3161,N_3121);
nor U3917 (N_3917,N_3063,N_3348);
or U3918 (N_3918,N_3084,N_3107);
nor U3919 (N_3919,N_3273,N_3162);
and U3920 (N_3920,N_3213,N_3039);
xnor U3921 (N_3921,N_3366,N_3313);
or U3922 (N_3922,N_3460,N_3457);
nor U3923 (N_3923,N_3306,N_3017);
nor U3924 (N_3924,N_3167,N_3165);
and U3925 (N_3925,N_3399,N_3139);
xor U3926 (N_3926,N_3029,N_3210);
or U3927 (N_3927,N_3142,N_3191);
or U3928 (N_3928,N_3311,N_3205);
xnor U3929 (N_3929,N_3027,N_3030);
or U3930 (N_3930,N_3334,N_3081);
nor U3931 (N_3931,N_3168,N_3262);
and U3932 (N_3932,N_3099,N_3050);
nand U3933 (N_3933,N_3291,N_3099);
or U3934 (N_3934,N_3193,N_3126);
and U3935 (N_3935,N_3022,N_3366);
xnor U3936 (N_3936,N_3218,N_3214);
nand U3937 (N_3937,N_3301,N_3116);
nor U3938 (N_3938,N_3449,N_3127);
xnor U3939 (N_3939,N_3127,N_3312);
nor U3940 (N_3940,N_3191,N_3449);
nand U3941 (N_3941,N_3267,N_3368);
xor U3942 (N_3942,N_3329,N_3491);
nand U3943 (N_3943,N_3341,N_3217);
nand U3944 (N_3944,N_3107,N_3070);
xnor U3945 (N_3945,N_3027,N_3108);
nor U3946 (N_3946,N_3435,N_3485);
nor U3947 (N_3947,N_3411,N_3336);
or U3948 (N_3948,N_3280,N_3176);
and U3949 (N_3949,N_3112,N_3318);
nor U3950 (N_3950,N_3153,N_3095);
nor U3951 (N_3951,N_3296,N_3116);
and U3952 (N_3952,N_3453,N_3217);
nor U3953 (N_3953,N_3263,N_3201);
xnor U3954 (N_3954,N_3232,N_3008);
and U3955 (N_3955,N_3108,N_3325);
or U3956 (N_3956,N_3112,N_3172);
nand U3957 (N_3957,N_3007,N_3495);
nor U3958 (N_3958,N_3089,N_3177);
or U3959 (N_3959,N_3090,N_3344);
xnor U3960 (N_3960,N_3160,N_3016);
xor U3961 (N_3961,N_3248,N_3187);
and U3962 (N_3962,N_3437,N_3228);
and U3963 (N_3963,N_3202,N_3231);
nand U3964 (N_3964,N_3133,N_3182);
and U3965 (N_3965,N_3419,N_3245);
or U3966 (N_3966,N_3000,N_3313);
nand U3967 (N_3967,N_3006,N_3199);
xor U3968 (N_3968,N_3321,N_3107);
nand U3969 (N_3969,N_3162,N_3365);
and U3970 (N_3970,N_3390,N_3387);
nor U3971 (N_3971,N_3106,N_3322);
nand U3972 (N_3972,N_3405,N_3146);
and U3973 (N_3973,N_3258,N_3349);
or U3974 (N_3974,N_3098,N_3391);
or U3975 (N_3975,N_3221,N_3377);
nand U3976 (N_3976,N_3189,N_3365);
or U3977 (N_3977,N_3000,N_3252);
nor U3978 (N_3978,N_3221,N_3082);
nand U3979 (N_3979,N_3205,N_3172);
or U3980 (N_3980,N_3384,N_3392);
and U3981 (N_3981,N_3487,N_3221);
or U3982 (N_3982,N_3287,N_3254);
or U3983 (N_3983,N_3378,N_3476);
nand U3984 (N_3984,N_3446,N_3441);
nand U3985 (N_3985,N_3007,N_3069);
nor U3986 (N_3986,N_3078,N_3297);
nand U3987 (N_3987,N_3272,N_3392);
nand U3988 (N_3988,N_3437,N_3163);
and U3989 (N_3989,N_3397,N_3197);
or U3990 (N_3990,N_3458,N_3111);
and U3991 (N_3991,N_3473,N_3330);
nor U3992 (N_3992,N_3308,N_3073);
xor U3993 (N_3993,N_3178,N_3433);
xor U3994 (N_3994,N_3262,N_3370);
nand U3995 (N_3995,N_3437,N_3133);
nand U3996 (N_3996,N_3054,N_3047);
or U3997 (N_3997,N_3061,N_3360);
and U3998 (N_3998,N_3135,N_3011);
nor U3999 (N_3999,N_3309,N_3480);
or U4000 (N_4000,N_3555,N_3680);
and U4001 (N_4001,N_3939,N_3959);
nor U4002 (N_4002,N_3576,N_3588);
xnor U4003 (N_4003,N_3670,N_3945);
nor U4004 (N_4004,N_3971,N_3821);
and U4005 (N_4005,N_3630,N_3844);
nand U4006 (N_4006,N_3778,N_3819);
or U4007 (N_4007,N_3523,N_3758);
and U4008 (N_4008,N_3503,N_3747);
or U4009 (N_4009,N_3866,N_3584);
xor U4010 (N_4010,N_3922,N_3927);
nand U4011 (N_4011,N_3962,N_3804);
or U4012 (N_4012,N_3956,N_3817);
nand U4013 (N_4013,N_3687,N_3721);
or U4014 (N_4014,N_3530,N_3910);
and U4015 (N_4015,N_3659,N_3952);
and U4016 (N_4016,N_3571,N_3566);
and U4017 (N_4017,N_3665,N_3560);
xor U4018 (N_4018,N_3568,N_3859);
nand U4019 (N_4019,N_3547,N_3996);
and U4020 (N_4020,N_3890,N_3975);
or U4021 (N_4021,N_3789,N_3963);
and U4022 (N_4022,N_3760,N_3838);
nor U4023 (N_4023,N_3668,N_3694);
xor U4024 (N_4024,N_3896,N_3660);
or U4025 (N_4025,N_3920,N_3671);
nor U4026 (N_4026,N_3990,N_3647);
nor U4027 (N_4027,N_3869,N_3782);
nand U4028 (N_4028,N_3763,N_3925);
xnor U4029 (N_4029,N_3621,N_3973);
nor U4030 (N_4030,N_3750,N_3867);
xor U4031 (N_4031,N_3985,N_3638);
nor U4032 (N_4032,N_3807,N_3998);
or U4033 (N_4033,N_3801,N_3813);
nand U4034 (N_4034,N_3913,N_3752);
or U4035 (N_4035,N_3533,N_3504);
nor U4036 (N_4036,N_3928,N_3527);
nor U4037 (N_4037,N_3650,N_3643);
nand U4038 (N_4038,N_3662,N_3957);
nand U4039 (N_4039,N_3641,N_3683);
nand U4040 (N_4040,N_3886,N_3761);
xor U4041 (N_4041,N_3961,N_3577);
or U4042 (N_4042,N_3772,N_3969);
and U4043 (N_4043,N_3567,N_3934);
nand U4044 (N_4044,N_3861,N_3532);
xnor U4045 (N_4045,N_3907,N_3651);
and U4046 (N_4046,N_3581,N_3582);
or U4047 (N_4047,N_3551,N_3738);
nor U4048 (N_4048,N_3874,N_3977);
xor U4049 (N_4049,N_3798,N_3953);
and U4050 (N_4050,N_3775,N_3833);
nor U4051 (N_4051,N_3639,N_3848);
nand U4052 (N_4052,N_3766,N_3993);
and U4053 (N_4053,N_3751,N_3597);
nor U4054 (N_4054,N_3725,N_3876);
nor U4055 (N_4055,N_3964,N_3793);
nand U4056 (N_4056,N_3737,N_3525);
nand U4057 (N_4057,N_3629,N_3535);
nand U4058 (N_4058,N_3575,N_3949);
xor U4059 (N_4059,N_3723,N_3553);
xnor U4060 (N_4060,N_3968,N_3712);
nand U4061 (N_4061,N_3831,N_3693);
nand U4062 (N_4062,N_3989,N_3537);
nor U4063 (N_4063,N_3787,N_3678);
nor U4064 (N_4064,N_3814,N_3921);
and U4065 (N_4065,N_3633,N_3919);
xnor U4066 (N_4066,N_3826,N_3636);
nor U4067 (N_4067,N_3578,N_3600);
nand U4068 (N_4068,N_3524,N_3997);
or U4069 (N_4069,N_3682,N_3649);
xor U4070 (N_4070,N_3673,N_3938);
nor U4071 (N_4071,N_3843,N_3809);
nor U4072 (N_4072,N_3640,N_3792);
nor U4073 (N_4073,N_3900,N_3840);
or U4074 (N_4074,N_3544,N_3739);
xor U4075 (N_4075,N_3736,N_3733);
xnor U4076 (N_4076,N_3740,N_3856);
nand U4077 (N_4077,N_3880,N_3828);
or U4078 (N_4078,N_3602,N_3623);
nand U4079 (N_4079,N_3923,N_3515);
nand U4080 (N_4080,N_3987,N_3594);
nor U4081 (N_4081,N_3773,N_3879);
nand U4082 (N_4082,N_3864,N_3868);
or U4083 (N_4083,N_3716,N_3951);
or U4084 (N_4084,N_3958,N_3654);
and U4085 (N_4085,N_3730,N_3516);
nand U4086 (N_4086,N_3619,N_3847);
nand U4087 (N_4087,N_3824,N_3912);
nor U4088 (N_4088,N_3734,N_3679);
xor U4089 (N_4089,N_3877,N_3944);
nor U4090 (N_4090,N_3726,N_3875);
nand U4091 (N_4091,N_3507,N_3574);
and U4092 (N_4092,N_3634,N_3852);
or U4093 (N_4093,N_3719,N_3690);
or U4094 (N_4094,N_3748,N_3918);
nand U4095 (N_4095,N_3691,N_3837);
nor U4096 (N_4096,N_3911,N_3892);
xnor U4097 (N_4097,N_3697,N_3510);
and U4098 (N_4098,N_3930,N_3779);
or U4099 (N_4099,N_3933,N_3846);
xor U4100 (N_4100,N_3935,N_3502);
nor U4101 (N_4101,N_3889,N_3699);
xnor U4102 (N_4102,N_3981,N_3882);
or U4103 (N_4103,N_3573,N_3811);
xor U4104 (N_4104,N_3931,N_3937);
and U4105 (N_4105,N_3803,N_3810);
xnor U4106 (N_4106,N_3857,N_3686);
nor U4107 (N_4107,N_3509,N_3714);
and U4108 (N_4108,N_3520,N_3790);
nor U4109 (N_4109,N_3598,N_3521);
xor U4110 (N_4110,N_3842,N_3771);
and U4111 (N_4111,N_3563,N_3617);
nor U4112 (N_4112,N_3983,N_3822);
or U4113 (N_4113,N_3505,N_3802);
nor U4114 (N_4114,N_3756,N_3603);
nand U4115 (N_4115,N_3548,N_3565);
nor U4116 (N_4116,N_3820,N_3514);
xnor U4117 (N_4117,N_3542,N_3606);
nand U4118 (N_4118,N_3749,N_3622);
and U4119 (N_4119,N_3709,N_3854);
nand U4120 (N_4120,N_3589,N_3897);
and U4121 (N_4121,N_3627,N_3902);
or U4122 (N_4122,N_3967,N_3599);
nor U4123 (N_4123,N_3684,N_3765);
or U4124 (N_4124,N_3746,N_3988);
xnor U4125 (N_4125,N_3950,N_3620);
nand U4126 (N_4126,N_3796,N_3508);
nand U4127 (N_4127,N_3755,N_3853);
xnor U4128 (N_4128,N_3592,N_3863);
xor U4129 (N_4129,N_3917,N_3805);
xnor U4130 (N_4130,N_3591,N_3865);
xor U4131 (N_4131,N_3899,N_3669);
and U4132 (N_4132,N_3695,N_3731);
and U4133 (N_4133,N_3871,N_3710);
and U4134 (N_4134,N_3586,N_3529);
xor U4135 (N_4135,N_3705,N_3898);
xor U4136 (N_4136,N_3966,N_3556);
nor U4137 (N_4137,N_3830,N_3637);
nor U4138 (N_4138,N_3557,N_3727);
nor U4139 (N_4139,N_3906,N_3717);
xnor U4140 (N_4140,N_3829,N_3745);
nand U4141 (N_4141,N_3901,N_3653);
or U4142 (N_4142,N_3614,N_3645);
and U4143 (N_4143,N_3500,N_3720);
nor U4144 (N_4144,N_3827,N_3593);
xnor U4145 (N_4145,N_3994,N_3908);
nand U4146 (N_4146,N_3743,N_3940);
or U4147 (N_4147,N_3929,N_3943);
or U4148 (N_4148,N_3692,N_3744);
xnor U4149 (N_4149,N_3800,N_3561);
nand U4150 (N_4150,N_3832,N_3681);
nor U4151 (N_4151,N_3873,N_3770);
xnor U4152 (N_4152,N_3794,N_3795);
or U4153 (N_4153,N_3613,N_3870);
or U4154 (N_4154,N_3825,N_3808);
or U4155 (N_4155,N_3979,N_3932);
or U4156 (N_4156,N_3788,N_3522);
and U4157 (N_4157,N_3815,N_3596);
xnor U4158 (N_4158,N_3905,N_3531);
xnor U4159 (N_4159,N_3546,N_3728);
nor U4160 (N_4160,N_3835,N_3724);
xnor U4161 (N_4161,N_3888,N_3858);
and U4162 (N_4162,N_3608,N_3528);
or U4163 (N_4163,N_3626,N_3845);
or U4164 (N_4164,N_3657,N_3628);
nand U4165 (N_4165,N_3947,N_3777);
and U4166 (N_4166,N_3955,N_3982);
nor U4167 (N_4167,N_3526,N_3978);
nand U4168 (N_4168,N_3569,N_3767);
and U4169 (N_4169,N_3718,N_3534);
xnor U4170 (N_4170,N_3554,N_3583);
xnor U4171 (N_4171,N_3652,N_3540);
or U4172 (N_4172,N_3774,N_3580);
and U4173 (N_4173,N_3924,N_3541);
or U4174 (N_4174,N_3536,N_3538);
xor U4175 (N_4175,N_3834,N_3585);
nand U4176 (N_4176,N_3762,N_3936);
and U4177 (N_4177,N_3618,N_3658);
and U4178 (N_4178,N_3909,N_3980);
and U4179 (N_4179,N_3549,N_3999);
or U4180 (N_4180,N_3759,N_3839);
xor U4181 (N_4181,N_3860,N_3974);
xnor U4182 (N_4182,N_3707,N_3688);
or U4183 (N_4183,N_3648,N_3706);
nand U4184 (N_4184,N_3885,N_3612);
or U4185 (N_4185,N_3704,N_3768);
and U4186 (N_4186,N_3519,N_3685);
and U4187 (N_4187,N_3722,N_3946);
nor U4188 (N_4188,N_3545,N_3550);
xor U4189 (N_4189,N_3797,N_3661);
nor U4190 (N_4190,N_3501,N_3587);
xnor U4191 (N_4191,N_3732,N_3517);
nor U4192 (N_4192,N_3632,N_3689);
xor U4193 (N_4193,N_3970,N_3784);
or U4194 (N_4194,N_3635,N_3667);
nand U4195 (N_4195,N_3506,N_3903);
nand U4196 (N_4196,N_3672,N_3711);
nand U4197 (N_4197,N_3995,N_3812);
or U4198 (N_4198,N_3823,N_3893);
nand U4199 (N_4199,N_3703,N_3862);
nand U4200 (N_4200,N_3625,N_3700);
xor U4201 (N_4201,N_3590,N_3604);
nand U4202 (N_4202,N_3579,N_3610);
or U4203 (N_4203,N_3713,N_3791);
nor U4204 (N_4204,N_3511,N_3729);
and U4205 (N_4205,N_3753,N_3564);
and U4206 (N_4206,N_3769,N_3702);
nor U4207 (N_4207,N_3984,N_3754);
nand U4208 (N_4208,N_3701,N_3609);
or U4209 (N_4209,N_3675,N_3572);
and U4210 (N_4210,N_3757,N_3543);
nor U4211 (N_4211,N_3783,N_3676);
nand U4212 (N_4212,N_3786,N_3849);
nor U4213 (N_4213,N_3872,N_3816);
nand U4214 (N_4214,N_3677,N_3850);
xor U4215 (N_4215,N_3941,N_3735);
or U4216 (N_4216,N_3664,N_3926);
nand U4217 (N_4217,N_3764,N_3878);
nand U4218 (N_4218,N_3891,N_3570);
nand U4219 (N_4219,N_3887,N_3601);
and U4220 (N_4220,N_3855,N_3642);
nor U4221 (N_4221,N_3991,N_3799);
and U4222 (N_4222,N_3965,N_3972);
nand U4223 (N_4223,N_3960,N_3986);
nand U4224 (N_4224,N_3611,N_3605);
nand U4225 (N_4225,N_3818,N_3644);
xnor U4226 (N_4226,N_3836,N_3948);
or U4227 (N_4227,N_3780,N_3741);
nor U4228 (N_4228,N_3806,N_3904);
xor U4229 (N_4229,N_3884,N_3698);
nor U4230 (N_4230,N_3562,N_3595);
and U4231 (N_4231,N_3615,N_3646);
xnor U4232 (N_4232,N_3624,N_3607);
or U4233 (N_4233,N_3841,N_3663);
xor U4234 (N_4234,N_3559,N_3512);
or U4235 (N_4235,N_3976,N_3781);
or U4236 (N_4236,N_3992,N_3942);
xnor U4237 (N_4237,N_3552,N_3851);
xnor U4238 (N_4238,N_3915,N_3539);
xnor U4239 (N_4239,N_3914,N_3558);
nand U4240 (N_4240,N_3916,N_3883);
xor U4241 (N_4241,N_3655,N_3715);
and U4242 (N_4242,N_3513,N_3895);
or U4243 (N_4243,N_3666,N_3708);
or U4244 (N_4244,N_3616,N_3881);
or U4245 (N_4245,N_3656,N_3954);
or U4246 (N_4246,N_3776,N_3696);
xor U4247 (N_4247,N_3631,N_3674);
or U4248 (N_4248,N_3894,N_3742);
nor U4249 (N_4249,N_3518,N_3785);
nand U4250 (N_4250,N_3513,N_3736);
nand U4251 (N_4251,N_3560,N_3702);
xnor U4252 (N_4252,N_3573,N_3893);
xor U4253 (N_4253,N_3515,N_3952);
xnor U4254 (N_4254,N_3953,N_3639);
nor U4255 (N_4255,N_3633,N_3685);
nor U4256 (N_4256,N_3623,N_3563);
and U4257 (N_4257,N_3678,N_3790);
xnor U4258 (N_4258,N_3868,N_3567);
or U4259 (N_4259,N_3670,N_3704);
and U4260 (N_4260,N_3918,N_3866);
and U4261 (N_4261,N_3882,N_3749);
nor U4262 (N_4262,N_3973,N_3612);
nand U4263 (N_4263,N_3862,N_3650);
or U4264 (N_4264,N_3957,N_3592);
or U4265 (N_4265,N_3688,N_3990);
and U4266 (N_4266,N_3952,N_3682);
or U4267 (N_4267,N_3630,N_3524);
nand U4268 (N_4268,N_3545,N_3827);
nand U4269 (N_4269,N_3690,N_3888);
nand U4270 (N_4270,N_3820,N_3985);
or U4271 (N_4271,N_3728,N_3881);
or U4272 (N_4272,N_3894,N_3720);
nand U4273 (N_4273,N_3584,N_3996);
or U4274 (N_4274,N_3693,N_3851);
nand U4275 (N_4275,N_3763,N_3596);
nand U4276 (N_4276,N_3718,N_3635);
and U4277 (N_4277,N_3958,N_3503);
and U4278 (N_4278,N_3530,N_3638);
xor U4279 (N_4279,N_3668,N_3796);
xnor U4280 (N_4280,N_3641,N_3679);
or U4281 (N_4281,N_3917,N_3752);
xor U4282 (N_4282,N_3824,N_3931);
xnor U4283 (N_4283,N_3522,N_3520);
xnor U4284 (N_4284,N_3933,N_3978);
or U4285 (N_4285,N_3598,N_3881);
nor U4286 (N_4286,N_3809,N_3771);
nor U4287 (N_4287,N_3922,N_3847);
or U4288 (N_4288,N_3722,N_3615);
or U4289 (N_4289,N_3875,N_3576);
and U4290 (N_4290,N_3558,N_3502);
or U4291 (N_4291,N_3939,N_3877);
nor U4292 (N_4292,N_3715,N_3927);
or U4293 (N_4293,N_3634,N_3888);
xor U4294 (N_4294,N_3995,N_3676);
or U4295 (N_4295,N_3622,N_3588);
or U4296 (N_4296,N_3843,N_3627);
and U4297 (N_4297,N_3767,N_3700);
and U4298 (N_4298,N_3715,N_3874);
and U4299 (N_4299,N_3570,N_3971);
or U4300 (N_4300,N_3879,N_3999);
xnor U4301 (N_4301,N_3598,N_3563);
nor U4302 (N_4302,N_3661,N_3875);
xor U4303 (N_4303,N_3620,N_3793);
or U4304 (N_4304,N_3712,N_3601);
nand U4305 (N_4305,N_3893,N_3816);
or U4306 (N_4306,N_3729,N_3642);
or U4307 (N_4307,N_3872,N_3674);
xor U4308 (N_4308,N_3919,N_3930);
and U4309 (N_4309,N_3590,N_3819);
or U4310 (N_4310,N_3606,N_3971);
and U4311 (N_4311,N_3592,N_3994);
and U4312 (N_4312,N_3723,N_3733);
nand U4313 (N_4313,N_3972,N_3712);
and U4314 (N_4314,N_3973,N_3800);
nor U4315 (N_4315,N_3779,N_3927);
nor U4316 (N_4316,N_3810,N_3679);
or U4317 (N_4317,N_3584,N_3719);
or U4318 (N_4318,N_3599,N_3525);
and U4319 (N_4319,N_3572,N_3546);
nor U4320 (N_4320,N_3528,N_3810);
nand U4321 (N_4321,N_3692,N_3790);
nor U4322 (N_4322,N_3676,N_3692);
and U4323 (N_4323,N_3884,N_3544);
and U4324 (N_4324,N_3665,N_3789);
xnor U4325 (N_4325,N_3783,N_3674);
nand U4326 (N_4326,N_3973,N_3765);
nor U4327 (N_4327,N_3921,N_3649);
and U4328 (N_4328,N_3928,N_3889);
or U4329 (N_4329,N_3889,N_3515);
xor U4330 (N_4330,N_3792,N_3852);
nand U4331 (N_4331,N_3644,N_3552);
and U4332 (N_4332,N_3802,N_3615);
nand U4333 (N_4333,N_3992,N_3530);
nor U4334 (N_4334,N_3985,N_3993);
or U4335 (N_4335,N_3591,N_3993);
xnor U4336 (N_4336,N_3959,N_3958);
nor U4337 (N_4337,N_3536,N_3943);
xor U4338 (N_4338,N_3872,N_3682);
or U4339 (N_4339,N_3773,N_3625);
nor U4340 (N_4340,N_3655,N_3706);
nor U4341 (N_4341,N_3557,N_3806);
and U4342 (N_4342,N_3742,N_3654);
nand U4343 (N_4343,N_3927,N_3714);
xnor U4344 (N_4344,N_3929,N_3732);
nor U4345 (N_4345,N_3628,N_3744);
nand U4346 (N_4346,N_3506,N_3694);
nand U4347 (N_4347,N_3968,N_3946);
and U4348 (N_4348,N_3706,N_3928);
xnor U4349 (N_4349,N_3842,N_3719);
nand U4350 (N_4350,N_3573,N_3664);
or U4351 (N_4351,N_3814,N_3681);
and U4352 (N_4352,N_3625,N_3917);
nand U4353 (N_4353,N_3983,N_3842);
xnor U4354 (N_4354,N_3986,N_3513);
nand U4355 (N_4355,N_3854,N_3562);
xnor U4356 (N_4356,N_3927,N_3503);
or U4357 (N_4357,N_3727,N_3675);
nor U4358 (N_4358,N_3658,N_3811);
xor U4359 (N_4359,N_3530,N_3582);
nand U4360 (N_4360,N_3525,N_3843);
xor U4361 (N_4361,N_3753,N_3727);
nor U4362 (N_4362,N_3776,N_3653);
nand U4363 (N_4363,N_3585,N_3550);
nand U4364 (N_4364,N_3628,N_3849);
and U4365 (N_4365,N_3860,N_3827);
xnor U4366 (N_4366,N_3764,N_3973);
nor U4367 (N_4367,N_3883,N_3610);
xor U4368 (N_4368,N_3602,N_3715);
nand U4369 (N_4369,N_3521,N_3718);
and U4370 (N_4370,N_3804,N_3602);
nor U4371 (N_4371,N_3688,N_3861);
nor U4372 (N_4372,N_3609,N_3503);
nor U4373 (N_4373,N_3793,N_3833);
or U4374 (N_4374,N_3882,N_3958);
and U4375 (N_4375,N_3734,N_3974);
nor U4376 (N_4376,N_3627,N_3801);
and U4377 (N_4377,N_3958,N_3708);
or U4378 (N_4378,N_3977,N_3592);
nor U4379 (N_4379,N_3631,N_3810);
and U4380 (N_4380,N_3922,N_3565);
or U4381 (N_4381,N_3855,N_3718);
nor U4382 (N_4382,N_3870,N_3559);
and U4383 (N_4383,N_3613,N_3553);
and U4384 (N_4384,N_3796,N_3772);
nor U4385 (N_4385,N_3707,N_3974);
or U4386 (N_4386,N_3549,N_3694);
nand U4387 (N_4387,N_3679,N_3698);
xor U4388 (N_4388,N_3590,N_3577);
and U4389 (N_4389,N_3824,N_3598);
nand U4390 (N_4390,N_3756,N_3983);
nand U4391 (N_4391,N_3957,N_3535);
nor U4392 (N_4392,N_3579,N_3685);
and U4393 (N_4393,N_3791,N_3953);
nor U4394 (N_4394,N_3784,N_3627);
and U4395 (N_4395,N_3517,N_3766);
nand U4396 (N_4396,N_3907,N_3653);
nand U4397 (N_4397,N_3858,N_3862);
nor U4398 (N_4398,N_3747,N_3845);
nor U4399 (N_4399,N_3756,N_3755);
nand U4400 (N_4400,N_3543,N_3742);
xnor U4401 (N_4401,N_3506,N_3762);
nand U4402 (N_4402,N_3725,N_3750);
nand U4403 (N_4403,N_3831,N_3879);
xor U4404 (N_4404,N_3664,N_3823);
and U4405 (N_4405,N_3695,N_3957);
nor U4406 (N_4406,N_3932,N_3680);
and U4407 (N_4407,N_3610,N_3627);
xor U4408 (N_4408,N_3919,N_3547);
and U4409 (N_4409,N_3658,N_3972);
or U4410 (N_4410,N_3851,N_3612);
nor U4411 (N_4411,N_3588,N_3865);
and U4412 (N_4412,N_3757,N_3802);
nor U4413 (N_4413,N_3543,N_3579);
nand U4414 (N_4414,N_3815,N_3681);
nor U4415 (N_4415,N_3969,N_3845);
nor U4416 (N_4416,N_3980,N_3620);
nor U4417 (N_4417,N_3507,N_3586);
xnor U4418 (N_4418,N_3920,N_3692);
or U4419 (N_4419,N_3908,N_3881);
or U4420 (N_4420,N_3777,N_3855);
or U4421 (N_4421,N_3804,N_3689);
or U4422 (N_4422,N_3977,N_3932);
and U4423 (N_4423,N_3691,N_3790);
nand U4424 (N_4424,N_3684,N_3719);
nor U4425 (N_4425,N_3914,N_3861);
xor U4426 (N_4426,N_3741,N_3666);
nand U4427 (N_4427,N_3796,N_3551);
nand U4428 (N_4428,N_3669,N_3863);
and U4429 (N_4429,N_3929,N_3738);
or U4430 (N_4430,N_3599,N_3764);
nand U4431 (N_4431,N_3785,N_3595);
xnor U4432 (N_4432,N_3891,N_3542);
and U4433 (N_4433,N_3786,N_3652);
and U4434 (N_4434,N_3705,N_3909);
nand U4435 (N_4435,N_3956,N_3954);
and U4436 (N_4436,N_3969,N_3826);
xnor U4437 (N_4437,N_3861,N_3564);
nor U4438 (N_4438,N_3664,N_3647);
xor U4439 (N_4439,N_3559,N_3955);
nor U4440 (N_4440,N_3522,N_3915);
nand U4441 (N_4441,N_3545,N_3861);
nor U4442 (N_4442,N_3996,N_3883);
xnor U4443 (N_4443,N_3573,N_3624);
or U4444 (N_4444,N_3651,N_3756);
or U4445 (N_4445,N_3852,N_3637);
nor U4446 (N_4446,N_3550,N_3655);
nor U4447 (N_4447,N_3899,N_3898);
and U4448 (N_4448,N_3808,N_3612);
and U4449 (N_4449,N_3843,N_3690);
xor U4450 (N_4450,N_3885,N_3884);
and U4451 (N_4451,N_3876,N_3614);
and U4452 (N_4452,N_3653,N_3749);
nor U4453 (N_4453,N_3744,N_3924);
nor U4454 (N_4454,N_3576,N_3906);
and U4455 (N_4455,N_3822,N_3808);
xnor U4456 (N_4456,N_3713,N_3706);
xor U4457 (N_4457,N_3952,N_3994);
nand U4458 (N_4458,N_3925,N_3915);
nand U4459 (N_4459,N_3846,N_3874);
or U4460 (N_4460,N_3881,N_3942);
nor U4461 (N_4461,N_3912,N_3793);
xnor U4462 (N_4462,N_3844,N_3797);
xnor U4463 (N_4463,N_3689,N_3680);
xnor U4464 (N_4464,N_3935,N_3548);
nor U4465 (N_4465,N_3596,N_3836);
xor U4466 (N_4466,N_3654,N_3965);
and U4467 (N_4467,N_3852,N_3642);
nand U4468 (N_4468,N_3591,N_3544);
or U4469 (N_4469,N_3782,N_3794);
and U4470 (N_4470,N_3533,N_3576);
xor U4471 (N_4471,N_3933,N_3610);
and U4472 (N_4472,N_3842,N_3761);
nor U4473 (N_4473,N_3909,N_3968);
nand U4474 (N_4474,N_3743,N_3830);
nor U4475 (N_4475,N_3538,N_3574);
nand U4476 (N_4476,N_3714,N_3968);
nand U4477 (N_4477,N_3780,N_3538);
and U4478 (N_4478,N_3576,N_3629);
nor U4479 (N_4479,N_3838,N_3826);
nand U4480 (N_4480,N_3887,N_3683);
nor U4481 (N_4481,N_3502,N_3520);
xnor U4482 (N_4482,N_3809,N_3517);
nand U4483 (N_4483,N_3930,N_3662);
and U4484 (N_4484,N_3825,N_3559);
and U4485 (N_4485,N_3838,N_3598);
and U4486 (N_4486,N_3682,N_3502);
xnor U4487 (N_4487,N_3821,N_3546);
and U4488 (N_4488,N_3786,N_3598);
or U4489 (N_4489,N_3873,N_3857);
and U4490 (N_4490,N_3773,N_3546);
nor U4491 (N_4491,N_3846,N_3810);
nand U4492 (N_4492,N_3772,N_3907);
or U4493 (N_4493,N_3867,N_3592);
xor U4494 (N_4494,N_3746,N_3835);
or U4495 (N_4495,N_3657,N_3678);
nand U4496 (N_4496,N_3850,N_3750);
or U4497 (N_4497,N_3954,N_3796);
and U4498 (N_4498,N_3826,N_3727);
nor U4499 (N_4499,N_3913,N_3690);
nor U4500 (N_4500,N_4267,N_4195);
xnor U4501 (N_4501,N_4248,N_4445);
or U4502 (N_4502,N_4370,N_4108);
and U4503 (N_4503,N_4156,N_4043);
nand U4504 (N_4504,N_4202,N_4342);
nand U4505 (N_4505,N_4443,N_4192);
xor U4506 (N_4506,N_4327,N_4268);
or U4507 (N_4507,N_4377,N_4137);
nand U4508 (N_4508,N_4476,N_4091);
xor U4509 (N_4509,N_4279,N_4232);
nor U4510 (N_4510,N_4219,N_4012);
or U4511 (N_4511,N_4483,N_4425);
nor U4512 (N_4512,N_4170,N_4098);
nand U4513 (N_4513,N_4235,N_4274);
xor U4514 (N_4514,N_4255,N_4431);
xnor U4515 (N_4515,N_4101,N_4074);
nand U4516 (N_4516,N_4461,N_4228);
and U4517 (N_4517,N_4452,N_4462);
or U4518 (N_4518,N_4079,N_4496);
or U4519 (N_4519,N_4331,N_4336);
nor U4520 (N_4520,N_4239,N_4242);
nor U4521 (N_4521,N_4308,N_4045);
nand U4522 (N_4522,N_4402,N_4293);
nand U4523 (N_4523,N_4198,N_4215);
nand U4524 (N_4524,N_4493,N_4314);
or U4525 (N_4525,N_4066,N_4063);
xor U4526 (N_4526,N_4148,N_4460);
and U4527 (N_4527,N_4280,N_4480);
nor U4528 (N_4528,N_4001,N_4399);
xnor U4529 (N_4529,N_4379,N_4028);
and U4530 (N_4530,N_4019,N_4374);
nor U4531 (N_4531,N_4058,N_4311);
and U4532 (N_4532,N_4492,N_4354);
nand U4533 (N_4533,N_4253,N_4162);
nand U4534 (N_4534,N_4060,N_4053);
nand U4535 (N_4535,N_4265,N_4024);
or U4536 (N_4536,N_4498,N_4105);
xor U4537 (N_4537,N_4154,N_4263);
and U4538 (N_4538,N_4360,N_4134);
and U4539 (N_4539,N_4054,N_4018);
nand U4540 (N_4540,N_4025,N_4306);
nor U4541 (N_4541,N_4307,N_4348);
nor U4542 (N_4542,N_4276,N_4014);
or U4543 (N_4543,N_4488,N_4023);
and U4544 (N_4544,N_4015,N_4486);
or U4545 (N_4545,N_4102,N_4287);
nor U4546 (N_4546,N_4187,N_4266);
or U4547 (N_4547,N_4473,N_4005);
nor U4548 (N_4548,N_4117,N_4426);
nand U4549 (N_4549,N_4386,N_4298);
nor U4550 (N_4550,N_4448,N_4305);
nor U4551 (N_4551,N_4437,N_4254);
nor U4552 (N_4552,N_4381,N_4435);
nor U4553 (N_4553,N_4471,N_4050);
xnor U4554 (N_4554,N_4391,N_4164);
nand U4555 (N_4555,N_4051,N_4479);
nand U4556 (N_4556,N_4344,N_4127);
nor U4557 (N_4557,N_4070,N_4133);
or U4558 (N_4558,N_4189,N_4206);
and U4559 (N_4559,N_4466,N_4169);
nand U4560 (N_4560,N_4447,N_4086);
nor U4561 (N_4561,N_4459,N_4118);
or U4562 (N_4562,N_4286,N_4487);
or U4563 (N_4563,N_4294,N_4396);
xor U4564 (N_4564,N_4039,N_4126);
and U4565 (N_4565,N_4037,N_4046);
xnor U4566 (N_4566,N_4361,N_4324);
or U4567 (N_4567,N_4457,N_4099);
or U4568 (N_4568,N_4289,N_4095);
or U4569 (N_4569,N_4233,N_4246);
and U4570 (N_4570,N_4155,N_4347);
and U4571 (N_4571,N_4092,N_4303);
and U4572 (N_4572,N_4330,N_4428);
nor U4573 (N_4573,N_4107,N_4190);
nand U4574 (N_4574,N_4325,N_4113);
nor U4575 (N_4575,N_4358,N_4338);
or U4576 (N_4576,N_4318,N_4357);
or U4577 (N_4577,N_4109,N_4158);
and U4578 (N_4578,N_4068,N_4458);
nor U4579 (N_4579,N_4090,N_4069);
xor U4580 (N_4580,N_4131,N_4475);
xnor U4581 (N_4581,N_4184,N_4321);
and U4582 (N_4582,N_4281,N_4097);
or U4583 (N_4583,N_4301,N_4337);
nor U4584 (N_4584,N_4009,N_4359);
nor U4585 (N_4585,N_4427,N_4363);
xor U4586 (N_4586,N_4423,N_4432);
nand U4587 (N_4587,N_4010,N_4499);
xnor U4588 (N_4588,N_4094,N_4186);
nand U4589 (N_4589,N_4188,N_4193);
nor U4590 (N_4590,N_4081,N_4339);
nor U4591 (N_4591,N_4047,N_4110);
xor U4592 (N_4592,N_4218,N_4002);
and U4593 (N_4593,N_4430,N_4332);
xor U4594 (N_4594,N_4234,N_4389);
nor U4595 (N_4595,N_4210,N_4290);
nor U4596 (N_4596,N_4404,N_4482);
xnor U4597 (N_4597,N_4468,N_4035);
xnor U4598 (N_4598,N_4317,N_4007);
nand U4599 (N_4599,N_4229,N_4222);
nor U4600 (N_4600,N_4204,N_4153);
xnor U4601 (N_4601,N_4146,N_4375);
or U4602 (N_4602,N_4088,N_4185);
xor U4603 (N_4603,N_4196,N_4161);
xor U4604 (N_4604,N_4143,N_4477);
nand U4605 (N_4605,N_4030,N_4173);
and U4606 (N_4606,N_4271,N_4387);
and U4607 (N_4607,N_4104,N_4304);
or U4608 (N_4608,N_4072,N_4182);
or U4609 (N_4609,N_4084,N_4212);
nand U4610 (N_4610,N_4419,N_4481);
or U4611 (N_4611,N_4369,N_4328);
and U4612 (N_4612,N_4403,N_4390);
xnor U4613 (N_4613,N_4484,N_4297);
or U4614 (N_4614,N_4440,N_4128);
nand U4615 (N_4615,N_4411,N_4175);
and U4616 (N_4616,N_4291,N_4217);
nand U4617 (N_4617,N_4315,N_4371);
nand U4618 (N_4618,N_4197,N_4407);
nand U4619 (N_4619,N_4089,N_4406);
or U4620 (N_4620,N_4221,N_4145);
nand U4621 (N_4621,N_4416,N_4405);
or U4622 (N_4622,N_4418,N_4214);
or U4623 (N_4623,N_4183,N_4252);
and U4624 (N_4624,N_4455,N_4353);
and U4625 (N_4625,N_4119,N_4272);
nor U4626 (N_4626,N_4004,N_4200);
xnor U4627 (N_4627,N_4135,N_4124);
nor U4628 (N_4628,N_4115,N_4278);
and U4629 (N_4629,N_4413,N_4450);
nor U4630 (N_4630,N_4008,N_4073);
or U4631 (N_4631,N_4167,N_4453);
and U4632 (N_4632,N_4159,N_4456);
and U4633 (N_4633,N_4245,N_4415);
nand U4634 (N_4634,N_4142,N_4016);
xor U4635 (N_4635,N_4284,N_4042);
nor U4636 (N_4636,N_4241,N_4121);
or U4637 (N_4637,N_4351,N_4000);
xor U4638 (N_4638,N_4168,N_4201);
nand U4639 (N_4639,N_4463,N_4464);
or U4640 (N_4640,N_4224,N_4116);
and U4641 (N_4641,N_4078,N_4065);
or U4642 (N_4642,N_4299,N_4223);
nor U4643 (N_4643,N_4454,N_4313);
nand U4644 (N_4644,N_4130,N_4244);
and U4645 (N_4645,N_4259,N_4439);
and U4646 (N_4646,N_4112,N_4341);
and U4647 (N_4647,N_4021,N_4231);
or U4648 (N_4648,N_4038,N_4376);
nand U4649 (N_4649,N_4157,N_4478);
and U4650 (N_4650,N_4366,N_4467);
and U4651 (N_4651,N_4378,N_4160);
and U4652 (N_4652,N_4216,N_4257);
and U4653 (N_4653,N_4367,N_4075);
nand U4654 (N_4654,N_4199,N_4041);
or U4655 (N_4655,N_4136,N_4057);
xor U4656 (N_4656,N_4180,N_4236);
and U4657 (N_4657,N_4444,N_4260);
and U4658 (N_4658,N_4087,N_4433);
or U4659 (N_4659,N_4174,N_4151);
and U4660 (N_4660,N_4048,N_4326);
and U4661 (N_4661,N_4372,N_4397);
and U4662 (N_4662,N_4044,N_4264);
xor U4663 (N_4663,N_4398,N_4408);
xnor U4664 (N_4664,N_4491,N_4420);
and U4665 (N_4665,N_4288,N_4395);
xnor U4666 (N_4666,N_4003,N_4017);
xnor U4667 (N_4667,N_4149,N_4334);
or U4668 (N_4668,N_4040,N_4364);
nor U4669 (N_4669,N_4085,N_4230);
nor U4670 (N_4670,N_4400,N_4368);
xnor U4671 (N_4671,N_4208,N_4247);
or U4672 (N_4672,N_4132,N_4049);
nand U4673 (N_4673,N_4238,N_4320);
or U4674 (N_4674,N_4220,N_4495);
nand U4675 (N_4675,N_4129,N_4093);
xnor U4676 (N_4676,N_4122,N_4138);
or U4677 (N_4677,N_4421,N_4032);
nand U4678 (N_4678,N_4275,N_4106);
nand U4679 (N_4679,N_4385,N_4329);
nand U4680 (N_4680,N_4269,N_4365);
nor U4681 (N_4681,N_4026,N_4139);
nand U4682 (N_4682,N_4277,N_4424);
nor U4683 (N_4683,N_4258,N_4392);
or U4684 (N_4684,N_4029,N_4422);
xor U4685 (N_4685,N_4414,N_4147);
or U4686 (N_4686,N_4322,N_4470);
xnor U4687 (N_4687,N_4125,N_4191);
xnor U4688 (N_4688,N_4373,N_4438);
or U4689 (N_4689,N_4059,N_4176);
and U4690 (N_4690,N_4056,N_4465);
nand U4691 (N_4691,N_4349,N_4485);
and U4692 (N_4692,N_4261,N_4096);
xnor U4693 (N_4693,N_4243,N_4302);
nor U4694 (N_4694,N_4114,N_4451);
nor U4695 (N_4695,N_4285,N_4262);
xnor U4696 (N_4696,N_4022,N_4394);
nand U4697 (N_4697,N_4172,N_4150);
or U4698 (N_4698,N_4227,N_4031);
or U4699 (N_4699,N_4077,N_4449);
nor U4700 (N_4700,N_4380,N_4209);
nand U4701 (N_4701,N_4382,N_4383);
xnor U4702 (N_4702,N_4335,N_4080);
and U4703 (N_4703,N_4052,N_4434);
nand U4704 (N_4704,N_4494,N_4384);
and U4705 (N_4705,N_4071,N_4120);
xnor U4706 (N_4706,N_4062,N_4429);
xor U4707 (N_4707,N_4061,N_4282);
or U4708 (N_4708,N_4177,N_4034);
nor U4709 (N_4709,N_4006,N_4103);
and U4710 (N_4710,N_4442,N_4350);
xor U4711 (N_4711,N_4140,N_4144);
and U4712 (N_4712,N_4203,N_4251);
or U4713 (N_4713,N_4310,N_4163);
xor U4714 (N_4714,N_4207,N_4489);
nor U4715 (N_4715,N_4205,N_4273);
and U4716 (N_4716,N_4295,N_4166);
or U4717 (N_4717,N_4256,N_4469);
nor U4718 (N_4718,N_4076,N_4346);
nor U4719 (N_4719,N_4213,N_4011);
nor U4720 (N_4720,N_4123,N_4141);
nand U4721 (N_4721,N_4020,N_4165);
xor U4722 (N_4722,N_4319,N_4152);
or U4723 (N_4723,N_4417,N_4340);
nand U4724 (N_4724,N_4333,N_4446);
or U4725 (N_4725,N_4027,N_4309);
or U4726 (N_4726,N_4067,N_4225);
xnor U4727 (N_4727,N_4179,N_4055);
xor U4728 (N_4728,N_4409,N_4393);
or U4729 (N_4729,N_4490,N_4036);
xor U4730 (N_4730,N_4323,N_4250);
or U4731 (N_4731,N_4033,N_4474);
and U4732 (N_4732,N_4111,N_4441);
nor U4733 (N_4733,N_4345,N_4083);
or U4734 (N_4734,N_4300,N_4412);
or U4735 (N_4735,N_4362,N_4181);
or U4736 (N_4736,N_4352,N_4316);
and U4737 (N_4737,N_4064,N_4171);
or U4738 (N_4738,N_4249,N_4292);
and U4739 (N_4739,N_4178,N_4356);
nand U4740 (N_4740,N_4343,N_4240);
nand U4741 (N_4741,N_4226,N_4283);
xor U4742 (N_4742,N_4237,N_4436);
xor U4743 (N_4743,N_4296,N_4082);
or U4744 (N_4744,N_4401,N_4497);
nor U4745 (N_4745,N_4355,N_4472);
nor U4746 (N_4746,N_4312,N_4388);
nand U4747 (N_4747,N_4013,N_4270);
xnor U4748 (N_4748,N_4194,N_4211);
nor U4749 (N_4749,N_4100,N_4410);
xor U4750 (N_4750,N_4380,N_4037);
or U4751 (N_4751,N_4202,N_4002);
and U4752 (N_4752,N_4318,N_4289);
xnor U4753 (N_4753,N_4338,N_4484);
nor U4754 (N_4754,N_4464,N_4235);
xor U4755 (N_4755,N_4106,N_4322);
or U4756 (N_4756,N_4485,N_4420);
nor U4757 (N_4757,N_4109,N_4297);
or U4758 (N_4758,N_4350,N_4179);
nand U4759 (N_4759,N_4443,N_4360);
nor U4760 (N_4760,N_4129,N_4400);
nor U4761 (N_4761,N_4494,N_4050);
or U4762 (N_4762,N_4387,N_4043);
nand U4763 (N_4763,N_4491,N_4182);
xnor U4764 (N_4764,N_4329,N_4181);
xor U4765 (N_4765,N_4338,N_4427);
and U4766 (N_4766,N_4160,N_4435);
nor U4767 (N_4767,N_4194,N_4461);
or U4768 (N_4768,N_4247,N_4482);
nand U4769 (N_4769,N_4059,N_4048);
nor U4770 (N_4770,N_4228,N_4174);
and U4771 (N_4771,N_4012,N_4065);
xor U4772 (N_4772,N_4020,N_4496);
xnor U4773 (N_4773,N_4008,N_4281);
xnor U4774 (N_4774,N_4208,N_4345);
xnor U4775 (N_4775,N_4153,N_4483);
or U4776 (N_4776,N_4371,N_4424);
xor U4777 (N_4777,N_4192,N_4029);
and U4778 (N_4778,N_4119,N_4437);
or U4779 (N_4779,N_4310,N_4440);
nand U4780 (N_4780,N_4045,N_4265);
xor U4781 (N_4781,N_4335,N_4433);
or U4782 (N_4782,N_4361,N_4344);
nand U4783 (N_4783,N_4093,N_4199);
and U4784 (N_4784,N_4441,N_4219);
nand U4785 (N_4785,N_4382,N_4172);
xnor U4786 (N_4786,N_4347,N_4194);
or U4787 (N_4787,N_4354,N_4005);
and U4788 (N_4788,N_4378,N_4086);
nand U4789 (N_4789,N_4399,N_4470);
xor U4790 (N_4790,N_4372,N_4378);
or U4791 (N_4791,N_4222,N_4323);
xor U4792 (N_4792,N_4226,N_4313);
or U4793 (N_4793,N_4221,N_4275);
or U4794 (N_4794,N_4209,N_4405);
xor U4795 (N_4795,N_4323,N_4157);
or U4796 (N_4796,N_4157,N_4071);
nand U4797 (N_4797,N_4115,N_4135);
and U4798 (N_4798,N_4418,N_4392);
xor U4799 (N_4799,N_4299,N_4175);
and U4800 (N_4800,N_4353,N_4436);
xnor U4801 (N_4801,N_4049,N_4088);
or U4802 (N_4802,N_4034,N_4123);
nor U4803 (N_4803,N_4420,N_4199);
nand U4804 (N_4804,N_4138,N_4406);
and U4805 (N_4805,N_4464,N_4332);
nor U4806 (N_4806,N_4368,N_4200);
nand U4807 (N_4807,N_4133,N_4111);
or U4808 (N_4808,N_4453,N_4373);
or U4809 (N_4809,N_4472,N_4460);
and U4810 (N_4810,N_4161,N_4428);
or U4811 (N_4811,N_4283,N_4359);
xor U4812 (N_4812,N_4242,N_4452);
nor U4813 (N_4813,N_4166,N_4084);
or U4814 (N_4814,N_4265,N_4137);
xnor U4815 (N_4815,N_4267,N_4150);
nand U4816 (N_4816,N_4375,N_4289);
or U4817 (N_4817,N_4069,N_4162);
or U4818 (N_4818,N_4441,N_4144);
nand U4819 (N_4819,N_4252,N_4276);
xor U4820 (N_4820,N_4256,N_4232);
xnor U4821 (N_4821,N_4354,N_4358);
xor U4822 (N_4822,N_4134,N_4329);
or U4823 (N_4823,N_4364,N_4170);
or U4824 (N_4824,N_4446,N_4238);
or U4825 (N_4825,N_4015,N_4125);
and U4826 (N_4826,N_4131,N_4334);
xor U4827 (N_4827,N_4077,N_4179);
nand U4828 (N_4828,N_4151,N_4067);
and U4829 (N_4829,N_4046,N_4053);
or U4830 (N_4830,N_4298,N_4161);
nand U4831 (N_4831,N_4468,N_4291);
xor U4832 (N_4832,N_4277,N_4299);
xor U4833 (N_4833,N_4364,N_4055);
and U4834 (N_4834,N_4147,N_4380);
nor U4835 (N_4835,N_4379,N_4424);
nand U4836 (N_4836,N_4477,N_4187);
xnor U4837 (N_4837,N_4096,N_4357);
nand U4838 (N_4838,N_4080,N_4233);
nor U4839 (N_4839,N_4244,N_4320);
xnor U4840 (N_4840,N_4234,N_4280);
nor U4841 (N_4841,N_4277,N_4045);
xnor U4842 (N_4842,N_4468,N_4080);
xnor U4843 (N_4843,N_4045,N_4286);
nor U4844 (N_4844,N_4278,N_4209);
and U4845 (N_4845,N_4340,N_4262);
or U4846 (N_4846,N_4179,N_4059);
or U4847 (N_4847,N_4383,N_4297);
xor U4848 (N_4848,N_4421,N_4126);
xnor U4849 (N_4849,N_4412,N_4022);
nand U4850 (N_4850,N_4039,N_4205);
and U4851 (N_4851,N_4247,N_4497);
xor U4852 (N_4852,N_4346,N_4466);
nor U4853 (N_4853,N_4108,N_4358);
or U4854 (N_4854,N_4389,N_4347);
or U4855 (N_4855,N_4347,N_4248);
or U4856 (N_4856,N_4303,N_4164);
and U4857 (N_4857,N_4282,N_4357);
and U4858 (N_4858,N_4298,N_4240);
nand U4859 (N_4859,N_4191,N_4480);
or U4860 (N_4860,N_4355,N_4291);
and U4861 (N_4861,N_4250,N_4191);
nor U4862 (N_4862,N_4250,N_4279);
or U4863 (N_4863,N_4245,N_4326);
xor U4864 (N_4864,N_4121,N_4239);
and U4865 (N_4865,N_4393,N_4478);
nand U4866 (N_4866,N_4369,N_4263);
and U4867 (N_4867,N_4007,N_4099);
nor U4868 (N_4868,N_4385,N_4315);
nand U4869 (N_4869,N_4126,N_4120);
nand U4870 (N_4870,N_4023,N_4168);
or U4871 (N_4871,N_4459,N_4403);
or U4872 (N_4872,N_4045,N_4238);
and U4873 (N_4873,N_4143,N_4436);
and U4874 (N_4874,N_4177,N_4019);
nor U4875 (N_4875,N_4474,N_4127);
xor U4876 (N_4876,N_4310,N_4271);
and U4877 (N_4877,N_4160,N_4044);
xor U4878 (N_4878,N_4002,N_4148);
nand U4879 (N_4879,N_4107,N_4070);
or U4880 (N_4880,N_4433,N_4279);
nand U4881 (N_4881,N_4224,N_4409);
nor U4882 (N_4882,N_4468,N_4340);
or U4883 (N_4883,N_4346,N_4000);
or U4884 (N_4884,N_4114,N_4032);
and U4885 (N_4885,N_4039,N_4299);
xnor U4886 (N_4886,N_4400,N_4225);
nor U4887 (N_4887,N_4058,N_4233);
nand U4888 (N_4888,N_4100,N_4317);
or U4889 (N_4889,N_4003,N_4361);
or U4890 (N_4890,N_4110,N_4414);
nand U4891 (N_4891,N_4466,N_4326);
and U4892 (N_4892,N_4287,N_4058);
and U4893 (N_4893,N_4476,N_4147);
and U4894 (N_4894,N_4099,N_4422);
nor U4895 (N_4895,N_4167,N_4477);
nor U4896 (N_4896,N_4077,N_4038);
and U4897 (N_4897,N_4239,N_4495);
and U4898 (N_4898,N_4113,N_4105);
and U4899 (N_4899,N_4232,N_4025);
nor U4900 (N_4900,N_4284,N_4034);
nor U4901 (N_4901,N_4120,N_4483);
and U4902 (N_4902,N_4068,N_4442);
nand U4903 (N_4903,N_4004,N_4195);
nor U4904 (N_4904,N_4219,N_4157);
nand U4905 (N_4905,N_4345,N_4048);
nand U4906 (N_4906,N_4219,N_4482);
and U4907 (N_4907,N_4470,N_4491);
nand U4908 (N_4908,N_4292,N_4304);
nor U4909 (N_4909,N_4368,N_4086);
nor U4910 (N_4910,N_4035,N_4158);
nand U4911 (N_4911,N_4282,N_4314);
and U4912 (N_4912,N_4112,N_4493);
and U4913 (N_4913,N_4094,N_4161);
and U4914 (N_4914,N_4215,N_4325);
or U4915 (N_4915,N_4406,N_4422);
nand U4916 (N_4916,N_4258,N_4395);
and U4917 (N_4917,N_4159,N_4185);
nand U4918 (N_4918,N_4375,N_4207);
xor U4919 (N_4919,N_4384,N_4185);
or U4920 (N_4920,N_4078,N_4487);
or U4921 (N_4921,N_4051,N_4212);
or U4922 (N_4922,N_4183,N_4173);
nand U4923 (N_4923,N_4484,N_4224);
and U4924 (N_4924,N_4225,N_4243);
or U4925 (N_4925,N_4471,N_4254);
or U4926 (N_4926,N_4367,N_4183);
xor U4927 (N_4927,N_4049,N_4389);
or U4928 (N_4928,N_4056,N_4103);
nand U4929 (N_4929,N_4151,N_4128);
nor U4930 (N_4930,N_4059,N_4321);
nand U4931 (N_4931,N_4219,N_4285);
and U4932 (N_4932,N_4020,N_4395);
nor U4933 (N_4933,N_4492,N_4143);
nand U4934 (N_4934,N_4116,N_4304);
nand U4935 (N_4935,N_4478,N_4354);
nand U4936 (N_4936,N_4089,N_4429);
nand U4937 (N_4937,N_4076,N_4247);
nor U4938 (N_4938,N_4159,N_4297);
nand U4939 (N_4939,N_4332,N_4419);
and U4940 (N_4940,N_4100,N_4245);
or U4941 (N_4941,N_4217,N_4400);
nor U4942 (N_4942,N_4299,N_4004);
nand U4943 (N_4943,N_4119,N_4212);
xnor U4944 (N_4944,N_4368,N_4337);
and U4945 (N_4945,N_4262,N_4474);
nor U4946 (N_4946,N_4336,N_4458);
nand U4947 (N_4947,N_4442,N_4008);
and U4948 (N_4948,N_4059,N_4282);
xor U4949 (N_4949,N_4281,N_4495);
nor U4950 (N_4950,N_4286,N_4449);
nor U4951 (N_4951,N_4019,N_4208);
xnor U4952 (N_4952,N_4245,N_4421);
or U4953 (N_4953,N_4242,N_4009);
xnor U4954 (N_4954,N_4134,N_4260);
and U4955 (N_4955,N_4061,N_4269);
and U4956 (N_4956,N_4171,N_4239);
nor U4957 (N_4957,N_4020,N_4322);
xnor U4958 (N_4958,N_4327,N_4297);
nor U4959 (N_4959,N_4227,N_4123);
and U4960 (N_4960,N_4465,N_4345);
xor U4961 (N_4961,N_4105,N_4077);
xnor U4962 (N_4962,N_4179,N_4184);
nand U4963 (N_4963,N_4371,N_4458);
and U4964 (N_4964,N_4426,N_4442);
xor U4965 (N_4965,N_4395,N_4287);
nor U4966 (N_4966,N_4137,N_4250);
and U4967 (N_4967,N_4386,N_4464);
or U4968 (N_4968,N_4152,N_4031);
nor U4969 (N_4969,N_4333,N_4279);
and U4970 (N_4970,N_4378,N_4294);
xnor U4971 (N_4971,N_4193,N_4422);
nor U4972 (N_4972,N_4412,N_4237);
nor U4973 (N_4973,N_4382,N_4444);
xor U4974 (N_4974,N_4482,N_4080);
nor U4975 (N_4975,N_4457,N_4417);
nor U4976 (N_4976,N_4329,N_4248);
xor U4977 (N_4977,N_4133,N_4329);
xnor U4978 (N_4978,N_4475,N_4296);
and U4979 (N_4979,N_4447,N_4298);
xnor U4980 (N_4980,N_4424,N_4410);
xnor U4981 (N_4981,N_4364,N_4355);
xnor U4982 (N_4982,N_4427,N_4253);
or U4983 (N_4983,N_4333,N_4219);
nand U4984 (N_4984,N_4261,N_4395);
xor U4985 (N_4985,N_4302,N_4135);
nand U4986 (N_4986,N_4299,N_4358);
nor U4987 (N_4987,N_4421,N_4165);
and U4988 (N_4988,N_4354,N_4488);
nand U4989 (N_4989,N_4093,N_4186);
nor U4990 (N_4990,N_4334,N_4232);
nand U4991 (N_4991,N_4364,N_4331);
and U4992 (N_4992,N_4075,N_4065);
nand U4993 (N_4993,N_4462,N_4227);
nor U4994 (N_4994,N_4120,N_4429);
and U4995 (N_4995,N_4239,N_4327);
or U4996 (N_4996,N_4330,N_4433);
nand U4997 (N_4997,N_4251,N_4069);
and U4998 (N_4998,N_4241,N_4457);
nand U4999 (N_4999,N_4121,N_4305);
or U5000 (N_5000,N_4911,N_4720);
nand U5001 (N_5001,N_4953,N_4864);
or U5002 (N_5002,N_4549,N_4683);
or U5003 (N_5003,N_4939,N_4988);
xnor U5004 (N_5004,N_4680,N_4728);
nor U5005 (N_5005,N_4517,N_4718);
nor U5006 (N_5006,N_4971,N_4968);
nor U5007 (N_5007,N_4936,N_4938);
xnor U5008 (N_5008,N_4651,N_4861);
xor U5009 (N_5009,N_4559,N_4814);
and U5010 (N_5010,N_4986,N_4975);
nor U5011 (N_5011,N_4949,N_4838);
nand U5012 (N_5012,N_4627,N_4620);
and U5013 (N_5013,N_4818,N_4622);
xor U5014 (N_5014,N_4855,N_4591);
nand U5015 (N_5015,N_4777,N_4990);
nor U5016 (N_5016,N_4852,N_4802);
or U5017 (N_5017,N_4639,N_4950);
nor U5018 (N_5018,N_4666,N_4661);
and U5019 (N_5019,N_4600,N_4800);
or U5020 (N_5020,N_4616,N_4682);
nor U5021 (N_5021,N_4824,N_4645);
xor U5022 (N_5022,N_4757,N_4635);
nand U5023 (N_5023,N_4779,N_4510);
or U5024 (N_5024,N_4671,N_4691);
xnor U5025 (N_5025,N_4959,N_4750);
nand U5026 (N_5026,N_4804,N_4656);
and U5027 (N_5027,N_4684,N_4603);
xor U5028 (N_5028,N_4652,N_4500);
nand U5029 (N_5029,N_4801,N_4688);
nand U5030 (N_5030,N_4992,N_4741);
nand U5031 (N_5031,N_4980,N_4659);
and U5032 (N_5032,N_4563,N_4927);
nand U5033 (N_5033,N_4715,N_4809);
nor U5034 (N_5034,N_4704,N_4839);
nand U5035 (N_5035,N_4538,N_4686);
or U5036 (N_5036,N_4907,N_4769);
nor U5037 (N_5037,N_4925,N_4908);
and U5038 (N_5038,N_4605,N_4888);
or U5039 (N_5039,N_4565,N_4951);
nor U5040 (N_5040,N_4884,N_4572);
xor U5041 (N_5041,N_4943,N_4826);
xor U5042 (N_5042,N_4606,N_4940);
nand U5043 (N_5043,N_4817,N_4999);
nor U5044 (N_5044,N_4646,N_4760);
nor U5045 (N_5045,N_4593,N_4756);
nand U5046 (N_5046,N_4995,N_4825);
nand U5047 (N_5047,N_4531,N_4762);
nor U5048 (N_5048,N_4729,N_4746);
nor U5049 (N_5049,N_4921,N_4931);
or U5050 (N_5050,N_4708,N_4709);
nor U5051 (N_5051,N_4535,N_4707);
nand U5052 (N_5052,N_4764,N_4573);
and U5053 (N_5053,N_4689,N_4650);
and U5054 (N_5054,N_4732,N_4542);
nand U5055 (N_5055,N_4952,N_4854);
nand U5056 (N_5056,N_4737,N_4929);
nand U5057 (N_5057,N_4964,N_4883);
or U5058 (N_5058,N_4768,N_4853);
nor U5059 (N_5059,N_4906,N_4880);
or U5060 (N_5060,N_4663,N_4594);
xnor U5061 (N_5061,N_4653,N_4629);
or U5062 (N_5062,N_4521,N_4934);
xor U5063 (N_5063,N_4615,N_4654);
nand U5064 (N_5064,N_4905,N_4920);
nand U5065 (N_5065,N_4841,N_4974);
nor U5066 (N_5066,N_4845,N_4643);
xnor U5067 (N_5067,N_4621,N_4548);
xnor U5068 (N_5068,N_4785,N_4783);
or U5069 (N_5069,N_4896,N_4870);
or U5070 (N_5070,N_4808,N_4843);
or U5071 (N_5071,N_4690,N_4900);
and U5072 (N_5072,N_4797,N_4942);
and U5073 (N_5073,N_4978,N_4789);
xor U5074 (N_5074,N_4984,N_4744);
nand U5075 (N_5075,N_4566,N_4892);
xnor U5076 (N_5076,N_4631,N_4543);
xnor U5077 (N_5077,N_4915,N_4946);
nand U5078 (N_5078,N_4893,N_4641);
or U5079 (N_5079,N_4881,N_4633);
xor U5080 (N_5080,N_4669,N_4956);
nor U5081 (N_5081,N_4523,N_4842);
or U5082 (N_5082,N_4514,N_4873);
nor U5083 (N_5083,N_4714,N_4862);
nand U5084 (N_5084,N_4840,N_4618);
or U5085 (N_5085,N_4596,N_4773);
or U5086 (N_5086,N_4963,N_4597);
or U5087 (N_5087,N_4960,N_4501);
nor U5088 (N_5088,N_4899,N_4657);
xor U5089 (N_5089,N_4534,N_4851);
or U5090 (N_5090,N_4677,N_4726);
xor U5091 (N_5091,N_4681,N_4532);
or U5092 (N_5092,N_4793,N_4664);
xor U5093 (N_5093,N_4810,N_4580);
nor U5094 (N_5094,N_4617,N_4721);
nand U5095 (N_5095,N_4765,N_4869);
nor U5096 (N_5096,N_4519,N_4694);
nor U5097 (N_5097,N_4571,N_4527);
and U5098 (N_5098,N_4700,N_4736);
nand U5099 (N_5099,N_4567,N_4898);
or U5100 (N_5100,N_4752,N_4926);
xor U5101 (N_5101,N_4576,N_4528);
and U5102 (N_5102,N_4835,N_4857);
nor U5103 (N_5103,N_4649,N_4917);
or U5104 (N_5104,N_4928,N_4705);
nand U5105 (N_5105,N_4577,N_4679);
and U5106 (N_5106,N_4676,N_4608);
nor U5107 (N_5107,N_4697,N_4987);
or U5108 (N_5108,N_4828,N_4623);
xnor U5109 (N_5109,N_4582,N_4526);
xor U5110 (N_5110,N_4546,N_4515);
and U5111 (N_5111,N_4813,N_4660);
and U5112 (N_5112,N_4642,N_4636);
xor U5113 (N_5113,N_4973,N_4876);
nor U5114 (N_5114,N_4844,N_4539);
xnor U5115 (N_5115,N_4701,N_4699);
nand U5116 (N_5116,N_4748,N_4829);
nor U5117 (N_5117,N_4935,N_4958);
nand U5118 (N_5118,N_4590,N_4551);
nand U5119 (N_5119,N_4722,N_4787);
nand U5120 (N_5120,N_4733,N_4866);
and U5121 (N_5121,N_4912,N_4834);
nor U5122 (N_5122,N_4882,N_4710);
nor U5123 (N_5123,N_4919,N_4578);
nand U5124 (N_5124,N_4613,N_4875);
or U5125 (N_5125,N_4833,N_4922);
nand U5126 (N_5126,N_4821,N_4822);
nand U5127 (N_5127,N_4560,N_4584);
nand U5128 (N_5128,N_4879,N_4871);
and U5129 (N_5129,N_4923,N_4674);
or U5130 (N_5130,N_4745,N_4819);
and U5131 (N_5131,N_4966,N_4668);
and U5132 (N_5132,N_4947,N_4753);
xor U5133 (N_5133,N_4957,N_4511);
and U5134 (N_5134,N_4781,N_4589);
nand U5135 (N_5135,N_4742,N_4670);
xnor U5136 (N_5136,N_4823,N_4901);
xnor U5137 (N_5137,N_4820,N_4743);
xor U5138 (N_5138,N_4692,N_4524);
xor U5139 (N_5139,N_4948,N_4730);
nand U5140 (N_5140,N_4860,N_4913);
nand U5141 (N_5141,N_4738,N_4562);
xnor U5142 (N_5142,N_4513,N_4739);
xor U5143 (N_5143,N_4581,N_4522);
nor U5144 (N_5144,N_4767,N_4972);
and U5145 (N_5145,N_4993,N_4607);
nor U5146 (N_5146,N_4867,N_4696);
xnor U5147 (N_5147,N_4976,N_4868);
nand U5148 (N_5148,N_4885,N_4556);
nand U5149 (N_5149,N_4561,N_4609);
nand U5150 (N_5150,N_4574,N_4507);
and U5151 (N_5151,N_4547,N_4614);
and U5152 (N_5152,N_4827,N_4658);
nor U5153 (N_5153,N_4585,N_4610);
xnor U5154 (N_5154,N_4792,N_4897);
nor U5155 (N_5155,N_4890,N_4508);
nand U5156 (N_5156,N_4759,N_4655);
nor U5157 (N_5157,N_4595,N_4602);
nor U5158 (N_5158,N_4932,N_4889);
nor U5159 (N_5159,N_4982,N_4717);
nor U5160 (N_5160,N_4695,N_4916);
and U5161 (N_5161,N_4969,N_4918);
xnor U5162 (N_5162,N_4552,N_4761);
nand U5163 (N_5163,N_4994,N_4540);
or U5164 (N_5164,N_4503,N_4647);
and U5165 (N_5165,N_4944,N_4774);
xnor U5166 (N_5166,N_4985,N_4583);
xnor U5167 (N_5167,N_4640,N_4568);
or U5168 (N_5168,N_4557,N_4619);
nand U5169 (N_5169,N_4863,N_4533);
nand U5170 (N_5170,N_4634,N_4795);
and U5171 (N_5171,N_4933,N_4848);
nand U5172 (N_5172,N_4983,N_4702);
and U5173 (N_5173,N_4586,N_4806);
nor U5174 (N_5174,N_4846,N_4588);
xnor U5175 (N_5175,N_4665,N_4570);
nor U5176 (N_5176,N_4758,N_4638);
nand U5177 (N_5177,N_4989,N_4790);
nor U5178 (N_5178,N_4754,N_4678);
xnor U5179 (N_5179,N_4604,N_4811);
or U5180 (N_5180,N_4910,N_4598);
nor U5181 (N_5181,N_4772,N_4740);
xnor U5182 (N_5182,N_4816,N_4991);
xnor U5183 (N_5183,N_4856,N_4837);
nor U5184 (N_5184,N_4662,N_4849);
nor U5185 (N_5185,N_4713,N_4812);
nor U5186 (N_5186,N_4903,N_4706);
or U5187 (N_5187,N_4979,N_4504);
xnor U5188 (N_5188,N_4667,N_4770);
or U5189 (N_5189,N_4798,N_4796);
nand U5190 (N_5190,N_4763,N_4723);
or U5191 (N_5191,N_4865,N_4902);
or U5192 (N_5192,N_4687,N_4569);
nand U5193 (N_5193,N_4536,N_4611);
or U5194 (N_5194,N_4815,N_4516);
nor U5195 (N_5195,N_4505,N_4564);
and U5196 (N_5196,N_4799,N_4545);
or U5197 (N_5197,N_4945,N_4878);
xor U5198 (N_5198,N_4977,N_4555);
nor U5199 (N_5199,N_4719,N_4778);
or U5200 (N_5200,N_4771,N_4924);
nand U5201 (N_5201,N_4967,N_4727);
xor U5202 (N_5202,N_4766,N_4587);
or U5203 (N_5203,N_4731,N_4998);
and U5204 (N_5204,N_4937,N_4632);
nand U5205 (N_5205,N_4877,N_4859);
or U5206 (N_5206,N_4558,N_4612);
xor U5207 (N_5207,N_4685,N_4698);
and U5208 (N_5208,N_4914,N_4575);
and U5209 (N_5209,N_4831,N_4648);
xnor U5210 (N_5210,N_4506,N_4541);
nand U5211 (N_5211,N_4579,N_4693);
xor U5212 (N_5212,N_4904,N_4626);
nand U5213 (N_5213,N_4637,N_4537);
and U5214 (N_5214,N_4512,N_4847);
nand U5215 (N_5215,N_4599,N_4941);
and U5216 (N_5216,N_4711,N_4909);
nor U5217 (N_5217,N_4930,N_4601);
nor U5218 (N_5218,N_4544,N_4962);
nor U5219 (N_5219,N_4712,N_4734);
nor U5220 (N_5220,N_4775,N_4749);
nor U5221 (N_5221,N_4794,N_4755);
nand U5222 (N_5222,N_4887,N_4735);
nand U5223 (N_5223,N_4782,N_4724);
nor U5224 (N_5224,N_4529,N_4891);
and U5225 (N_5225,N_4803,N_4850);
and U5226 (N_5226,N_4895,N_4858);
and U5227 (N_5227,N_4630,N_4725);
nor U5228 (N_5228,N_4747,N_4550);
nand U5229 (N_5229,N_4751,N_4624);
and U5230 (N_5230,N_4780,N_4675);
nand U5231 (N_5231,N_4673,N_4961);
nor U5232 (N_5232,N_4786,N_4886);
xnor U5233 (N_5233,N_4554,N_4955);
xor U5234 (N_5234,N_4874,N_4502);
and U5235 (N_5235,N_4628,N_4996);
nand U5236 (N_5236,N_4791,N_4894);
or U5237 (N_5237,N_4518,N_4625);
xor U5238 (N_5238,N_4644,N_4836);
nand U5239 (N_5239,N_4965,N_4784);
and U5240 (N_5240,N_4520,N_4716);
nor U5241 (N_5241,N_4509,N_4776);
and U5242 (N_5242,N_4872,N_4981);
nand U5243 (N_5243,N_4954,N_4830);
nand U5244 (N_5244,N_4592,N_4703);
xnor U5245 (N_5245,N_4807,N_4553);
nor U5246 (N_5246,N_4530,N_4672);
and U5247 (N_5247,N_4970,N_4805);
nor U5248 (N_5248,N_4525,N_4997);
xor U5249 (N_5249,N_4788,N_4832);
nor U5250 (N_5250,N_4609,N_4724);
nor U5251 (N_5251,N_4966,N_4580);
nor U5252 (N_5252,N_4944,N_4530);
or U5253 (N_5253,N_4950,N_4626);
and U5254 (N_5254,N_4937,N_4959);
or U5255 (N_5255,N_4812,N_4762);
or U5256 (N_5256,N_4937,N_4935);
nand U5257 (N_5257,N_4638,N_4839);
or U5258 (N_5258,N_4913,N_4720);
xor U5259 (N_5259,N_4951,N_4814);
nand U5260 (N_5260,N_4856,N_4639);
nand U5261 (N_5261,N_4884,N_4880);
nand U5262 (N_5262,N_4756,N_4702);
and U5263 (N_5263,N_4985,N_4737);
and U5264 (N_5264,N_4731,N_4842);
nand U5265 (N_5265,N_4646,N_4691);
or U5266 (N_5266,N_4923,N_4567);
nor U5267 (N_5267,N_4742,N_4615);
or U5268 (N_5268,N_4678,N_4728);
or U5269 (N_5269,N_4505,N_4645);
and U5270 (N_5270,N_4916,N_4605);
and U5271 (N_5271,N_4627,N_4702);
nor U5272 (N_5272,N_4780,N_4913);
or U5273 (N_5273,N_4552,N_4514);
and U5274 (N_5274,N_4711,N_4992);
or U5275 (N_5275,N_4950,N_4516);
and U5276 (N_5276,N_4730,N_4607);
nand U5277 (N_5277,N_4509,N_4811);
nor U5278 (N_5278,N_4503,N_4995);
nand U5279 (N_5279,N_4623,N_4924);
or U5280 (N_5280,N_4634,N_4749);
and U5281 (N_5281,N_4515,N_4896);
xor U5282 (N_5282,N_4706,N_4664);
xor U5283 (N_5283,N_4998,N_4854);
nor U5284 (N_5284,N_4778,N_4814);
and U5285 (N_5285,N_4936,N_4869);
nand U5286 (N_5286,N_4979,N_4545);
xnor U5287 (N_5287,N_4858,N_4834);
or U5288 (N_5288,N_4912,N_4883);
nand U5289 (N_5289,N_4562,N_4531);
nand U5290 (N_5290,N_4858,N_4855);
and U5291 (N_5291,N_4882,N_4921);
nand U5292 (N_5292,N_4851,N_4842);
and U5293 (N_5293,N_4583,N_4655);
nor U5294 (N_5294,N_4598,N_4596);
or U5295 (N_5295,N_4839,N_4821);
xnor U5296 (N_5296,N_4892,N_4710);
xor U5297 (N_5297,N_4988,N_4997);
nand U5298 (N_5298,N_4946,N_4971);
nand U5299 (N_5299,N_4564,N_4562);
or U5300 (N_5300,N_4943,N_4768);
xor U5301 (N_5301,N_4551,N_4839);
or U5302 (N_5302,N_4593,N_4909);
and U5303 (N_5303,N_4823,N_4667);
xnor U5304 (N_5304,N_4965,N_4954);
xnor U5305 (N_5305,N_4929,N_4579);
and U5306 (N_5306,N_4699,N_4723);
or U5307 (N_5307,N_4535,N_4655);
nand U5308 (N_5308,N_4679,N_4871);
xnor U5309 (N_5309,N_4902,N_4776);
or U5310 (N_5310,N_4684,N_4775);
xor U5311 (N_5311,N_4859,N_4862);
nand U5312 (N_5312,N_4782,N_4727);
nor U5313 (N_5313,N_4679,N_4944);
nor U5314 (N_5314,N_4647,N_4757);
nand U5315 (N_5315,N_4586,N_4801);
and U5316 (N_5316,N_4910,N_4955);
nand U5317 (N_5317,N_4664,N_4959);
nand U5318 (N_5318,N_4709,N_4982);
and U5319 (N_5319,N_4706,N_4955);
or U5320 (N_5320,N_4904,N_4600);
xor U5321 (N_5321,N_4592,N_4721);
xnor U5322 (N_5322,N_4508,N_4506);
or U5323 (N_5323,N_4900,N_4644);
nand U5324 (N_5324,N_4948,N_4621);
nand U5325 (N_5325,N_4776,N_4556);
and U5326 (N_5326,N_4982,N_4800);
xor U5327 (N_5327,N_4787,N_4620);
and U5328 (N_5328,N_4930,N_4810);
xnor U5329 (N_5329,N_4994,N_4742);
nor U5330 (N_5330,N_4971,N_4621);
and U5331 (N_5331,N_4924,N_4728);
xor U5332 (N_5332,N_4607,N_4745);
and U5333 (N_5333,N_4600,N_4780);
nand U5334 (N_5334,N_4939,N_4693);
or U5335 (N_5335,N_4832,N_4782);
and U5336 (N_5336,N_4647,N_4733);
and U5337 (N_5337,N_4838,N_4993);
xnor U5338 (N_5338,N_4542,N_4640);
or U5339 (N_5339,N_4953,N_4751);
and U5340 (N_5340,N_4953,N_4525);
or U5341 (N_5341,N_4856,N_4934);
nand U5342 (N_5342,N_4703,N_4779);
xor U5343 (N_5343,N_4659,N_4845);
xnor U5344 (N_5344,N_4971,N_4641);
nand U5345 (N_5345,N_4529,N_4957);
and U5346 (N_5346,N_4559,N_4805);
xnor U5347 (N_5347,N_4803,N_4749);
or U5348 (N_5348,N_4870,N_4892);
xnor U5349 (N_5349,N_4574,N_4789);
or U5350 (N_5350,N_4648,N_4822);
and U5351 (N_5351,N_4576,N_4773);
and U5352 (N_5352,N_4611,N_4713);
nor U5353 (N_5353,N_4843,N_4875);
nor U5354 (N_5354,N_4770,N_4951);
xnor U5355 (N_5355,N_4513,N_4521);
or U5356 (N_5356,N_4833,N_4834);
and U5357 (N_5357,N_4563,N_4843);
nand U5358 (N_5358,N_4528,N_4944);
nand U5359 (N_5359,N_4597,N_4869);
nor U5360 (N_5360,N_4520,N_4696);
or U5361 (N_5361,N_4632,N_4649);
xor U5362 (N_5362,N_4986,N_4793);
nand U5363 (N_5363,N_4514,N_4632);
nand U5364 (N_5364,N_4716,N_4930);
nand U5365 (N_5365,N_4825,N_4932);
nor U5366 (N_5366,N_4974,N_4917);
nor U5367 (N_5367,N_4621,N_4655);
xor U5368 (N_5368,N_4805,N_4926);
xnor U5369 (N_5369,N_4908,N_4725);
nor U5370 (N_5370,N_4598,N_4667);
xnor U5371 (N_5371,N_4911,N_4585);
and U5372 (N_5372,N_4890,N_4656);
xnor U5373 (N_5373,N_4732,N_4977);
and U5374 (N_5374,N_4782,N_4656);
or U5375 (N_5375,N_4560,N_4523);
or U5376 (N_5376,N_4665,N_4609);
xor U5377 (N_5377,N_4787,N_4891);
nand U5378 (N_5378,N_4687,N_4873);
xnor U5379 (N_5379,N_4850,N_4567);
nor U5380 (N_5380,N_4927,N_4875);
or U5381 (N_5381,N_4834,N_4896);
nand U5382 (N_5382,N_4624,N_4925);
nand U5383 (N_5383,N_4790,N_4755);
xnor U5384 (N_5384,N_4509,N_4580);
or U5385 (N_5385,N_4703,N_4607);
or U5386 (N_5386,N_4875,N_4996);
nand U5387 (N_5387,N_4985,N_4922);
xnor U5388 (N_5388,N_4901,N_4657);
xnor U5389 (N_5389,N_4686,N_4635);
nor U5390 (N_5390,N_4683,N_4818);
xor U5391 (N_5391,N_4677,N_4632);
or U5392 (N_5392,N_4989,N_4729);
nor U5393 (N_5393,N_4897,N_4891);
xor U5394 (N_5394,N_4954,N_4983);
nand U5395 (N_5395,N_4858,N_4933);
or U5396 (N_5396,N_4963,N_4611);
nand U5397 (N_5397,N_4585,N_4822);
xnor U5398 (N_5398,N_4820,N_4585);
nand U5399 (N_5399,N_4553,N_4853);
and U5400 (N_5400,N_4716,N_4713);
and U5401 (N_5401,N_4804,N_4845);
nor U5402 (N_5402,N_4853,N_4938);
and U5403 (N_5403,N_4827,N_4805);
nand U5404 (N_5404,N_4807,N_4605);
xnor U5405 (N_5405,N_4850,N_4889);
xnor U5406 (N_5406,N_4710,N_4979);
nor U5407 (N_5407,N_4747,N_4634);
nand U5408 (N_5408,N_4661,N_4625);
nand U5409 (N_5409,N_4910,N_4633);
and U5410 (N_5410,N_4655,N_4593);
xor U5411 (N_5411,N_4733,N_4873);
or U5412 (N_5412,N_4632,N_4959);
xor U5413 (N_5413,N_4956,N_4500);
xnor U5414 (N_5414,N_4936,N_4632);
and U5415 (N_5415,N_4613,N_4843);
nor U5416 (N_5416,N_4903,N_4995);
or U5417 (N_5417,N_4697,N_4888);
and U5418 (N_5418,N_4672,N_4632);
or U5419 (N_5419,N_4690,N_4662);
xnor U5420 (N_5420,N_4516,N_4643);
nor U5421 (N_5421,N_4690,N_4897);
nor U5422 (N_5422,N_4746,N_4752);
xnor U5423 (N_5423,N_4978,N_4592);
or U5424 (N_5424,N_4548,N_4721);
xor U5425 (N_5425,N_4699,N_4742);
and U5426 (N_5426,N_4866,N_4601);
xor U5427 (N_5427,N_4601,N_4819);
or U5428 (N_5428,N_4992,N_4613);
xnor U5429 (N_5429,N_4914,N_4639);
nor U5430 (N_5430,N_4629,N_4667);
and U5431 (N_5431,N_4921,N_4736);
and U5432 (N_5432,N_4627,N_4791);
xor U5433 (N_5433,N_4893,N_4935);
xnor U5434 (N_5434,N_4682,N_4887);
nand U5435 (N_5435,N_4714,N_4741);
nor U5436 (N_5436,N_4562,N_4988);
xor U5437 (N_5437,N_4825,N_4604);
nand U5438 (N_5438,N_4861,N_4979);
xor U5439 (N_5439,N_4751,N_4927);
nor U5440 (N_5440,N_4936,N_4971);
nand U5441 (N_5441,N_4891,N_4820);
xor U5442 (N_5442,N_4767,N_4917);
nand U5443 (N_5443,N_4839,N_4679);
and U5444 (N_5444,N_4645,N_4882);
and U5445 (N_5445,N_4826,N_4903);
nor U5446 (N_5446,N_4631,N_4761);
xor U5447 (N_5447,N_4973,N_4700);
and U5448 (N_5448,N_4897,N_4869);
nand U5449 (N_5449,N_4540,N_4788);
nor U5450 (N_5450,N_4552,N_4554);
xor U5451 (N_5451,N_4818,N_4680);
nand U5452 (N_5452,N_4942,N_4609);
nand U5453 (N_5453,N_4749,N_4960);
or U5454 (N_5454,N_4559,N_4859);
and U5455 (N_5455,N_4906,N_4652);
nand U5456 (N_5456,N_4585,N_4693);
or U5457 (N_5457,N_4784,N_4833);
or U5458 (N_5458,N_4537,N_4914);
and U5459 (N_5459,N_4977,N_4685);
xnor U5460 (N_5460,N_4800,N_4572);
and U5461 (N_5461,N_4845,N_4970);
nor U5462 (N_5462,N_4781,N_4857);
nor U5463 (N_5463,N_4829,N_4678);
nand U5464 (N_5464,N_4775,N_4951);
nand U5465 (N_5465,N_4963,N_4886);
nor U5466 (N_5466,N_4732,N_4994);
nand U5467 (N_5467,N_4514,N_4659);
and U5468 (N_5468,N_4520,N_4622);
or U5469 (N_5469,N_4887,N_4729);
or U5470 (N_5470,N_4527,N_4629);
xnor U5471 (N_5471,N_4635,N_4539);
nand U5472 (N_5472,N_4898,N_4928);
and U5473 (N_5473,N_4689,N_4546);
and U5474 (N_5474,N_4781,N_4920);
and U5475 (N_5475,N_4880,N_4620);
or U5476 (N_5476,N_4779,N_4832);
and U5477 (N_5477,N_4690,N_4848);
xor U5478 (N_5478,N_4671,N_4881);
nor U5479 (N_5479,N_4712,N_4869);
nor U5480 (N_5480,N_4747,N_4892);
or U5481 (N_5481,N_4815,N_4954);
nor U5482 (N_5482,N_4739,N_4810);
or U5483 (N_5483,N_4522,N_4706);
or U5484 (N_5484,N_4868,N_4531);
nor U5485 (N_5485,N_4833,N_4607);
or U5486 (N_5486,N_4638,N_4504);
nor U5487 (N_5487,N_4982,N_4755);
nor U5488 (N_5488,N_4615,N_4853);
nand U5489 (N_5489,N_4502,N_4567);
xor U5490 (N_5490,N_4898,N_4710);
nand U5491 (N_5491,N_4886,N_4864);
or U5492 (N_5492,N_4806,N_4568);
xor U5493 (N_5493,N_4547,N_4698);
nor U5494 (N_5494,N_4991,N_4826);
or U5495 (N_5495,N_4727,N_4735);
nand U5496 (N_5496,N_4737,N_4612);
and U5497 (N_5497,N_4683,N_4848);
or U5498 (N_5498,N_4542,N_4661);
and U5499 (N_5499,N_4697,N_4717);
nor U5500 (N_5500,N_5473,N_5117);
nor U5501 (N_5501,N_5136,N_5306);
or U5502 (N_5502,N_5172,N_5255);
and U5503 (N_5503,N_5234,N_5256);
xor U5504 (N_5504,N_5343,N_5402);
or U5505 (N_5505,N_5395,N_5303);
nand U5506 (N_5506,N_5493,N_5074);
nand U5507 (N_5507,N_5382,N_5289);
nand U5508 (N_5508,N_5203,N_5463);
or U5509 (N_5509,N_5328,N_5272);
and U5510 (N_5510,N_5434,N_5362);
nor U5511 (N_5511,N_5167,N_5044);
xnor U5512 (N_5512,N_5386,N_5041);
or U5513 (N_5513,N_5424,N_5403);
nor U5514 (N_5514,N_5099,N_5495);
nor U5515 (N_5515,N_5292,N_5469);
xor U5516 (N_5516,N_5235,N_5072);
or U5517 (N_5517,N_5219,N_5441);
xnor U5518 (N_5518,N_5216,N_5060);
nand U5519 (N_5519,N_5271,N_5051);
nand U5520 (N_5520,N_5438,N_5000);
or U5521 (N_5521,N_5221,N_5465);
nor U5522 (N_5522,N_5092,N_5375);
nand U5523 (N_5523,N_5146,N_5214);
nand U5524 (N_5524,N_5419,N_5036);
nand U5525 (N_5525,N_5442,N_5475);
or U5526 (N_5526,N_5459,N_5162);
nand U5527 (N_5527,N_5327,N_5261);
or U5528 (N_5528,N_5211,N_5253);
nand U5529 (N_5529,N_5405,N_5288);
or U5530 (N_5530,N_5321,N_5389);
xor U5531 (N_5531,N_5308,N_5010);
xnor U5532 (N_5532,N_5397,N_5038);
and U5533 (N_5533,N_5200,N_5244);
nand U5534 (N_5534,N_5055,N_5012);
nor U5535 (N_5535,N_5432,N_5298);
nand U5536 (N_5536,N_5366,N_5447);
nor U5537 (N_5537,N_5263,N_5224);
xor U5538 (N_5538,N_5333,N_5478);
nor U5539 (N_5539,N_5490,N_5317);
nand U5540 (N_5540,N_5118,N_5090);
or U5541 (N_5541,N_5141,N_5322);
and U5542 (N_5542,N_5370,N_5340);
and U5543 (N_5543,N_5407,N_5057);
or U5544 (N_5544,N_5396,N_5264);
xnor U5545 (N_5545,N_5138,N_5229);
xor U5546 (N_5546,N_5128,N_5131);
nor U5547 (N_5547,N_5132,N_5309);
nor U5548 (N_5548,N_5470,N_5154);
and U5549 (N_5549,N_5350,N_5011);
xor U5550 (N_5550,N_5440,N_5159);
xor U5551 (N_5551,N_5013,N_5369);
nand U5552 (N_5552,N_5349,N_5363);
or U5553 (N_5553,N_5076,N_5058);
xor U5554 (N_5554,N_5399,N_5019);
nor U5555 (N_5555,N_5455,N_5086);
or U5556 (N_5556,N_5247,N_5102);
nor U5557 (N_5557,N_5173,N_5122);
nor U5558 (N_5558,N_5284,N_5079);
or U5559 (N_5559,N_5491,N_5178);
and U5560 (N_5560,N_5240,N_5135);
xor U5561 (N_5561,N_5291,N_5281);
or U5562 (N_5562,N_5191,N_5056);
xor U5563 (N_5563,N_5184,N_5144);
and U5564 (N_5564,N_5107,N_5300);
or U5565 (N_5565,N_5496,N_5006);
or U5566 (N_5566,N_5094,N_5116);
nor U5567 (N_5567,N_5242,N_5112);
xor U5568 (N_5568,N_5198,N_5104);
and U5569 (N_5569,N_5045,N_5276);
xnor U5570 (N_5570,N_5452,N_5464);
nor U5571 (N_5571,N_5279,N_5325);
and U5572 (N_5572,N_5319,N_5114);
xnor U5573 (N_5573,N_5422,N_5367);
nor U5574 (N_5574,N_5471,N_5228);
xor U5575 (N_5575,N_5212,N_5391);
and U5576 (N_5576,N_5275,N_5258);
nand U5577 (N_5577,N_5472,N_5476);
nand U5578 (N_5578,N_5220,N_5456);
nand U5579 (N_5579,N_5311,N_5278);
xnor U5580 (N_5580,N_5050,N_5341);
nand U5581 (N_5581,N_5048,N_5108);
or U5582 (N_5582,N_5194,N_5208);
nand U5583 (N_5583,N_5005,N_5286);
nand U5584 (N_5584,N_5204,N_5448);
xnor U5585 (N_5585,N_5449,N_5192);
or U5586 (N_5586,N_5037,N_5304);
and U5587 (N_5587,N_5357,N_5254);
nand U5588 (N_5588,N_5101,N_5302);
nand U5589 (N_5589,N_5123,N_5323);
nand U5590 (N_5590,N_5032,N_5031);
nor U5591 (N_5591,N_5338,N_5400);
or U5592 (N_5592,N_5065,N_5436);
xor U5593 (N_5593,N_5481,N_5001);
nor U5594 (N_5594,N_5140,N_5385);
or U5595 (N_5595,N_5195,N_5067);
xor U5596 (N_5596,N_5164,N_5046);
or U5597 (N_5597,N_5315,N_5273);
nand U5598 (N_5598,N_5175,N_5153);
nor U5599 (N_5599,N_5249,N_5433);
or U5600 (N_5600,N_5009,N_5166);
and U5601 (N_5601,N_5354,N_5207);
nand U5602 (N_5602,N_5411,N_5426);
nor U5603 (N_5603,N_5121,N_5115);
nand U5604 (N_5604,N_5125,N_5073);
and U5605 (N_5605,N_5316,N_5028);
xnor U5606 (N_5606,N_5295,N_5080);
nor U5607 (N_5607,N_5457,N_5398);
nand U5608 (N_5608,N_5324,N_5483);
xor U5609 (N_5609,N_5485,N_5494);
xnor U5610 (N_5610,N_5142,N_5205);
xor U5611 (N_5611,N_5071,N_5230);
or U5612 (N_5612,N_5078,N_5039);
or U5613 (N_5613,N_5344,N_5372);
or U5614 (N_5614,N_5181,N_5130);
nor U5615 (N_5615,N_5210,N_5042);
or U5616 (N_5616,N_5270,N_5280);
or U5617 (N_5617,N_5332,N_5008);
nor U5618 (N_5618,N_5353,N_5299);
nor U5619 (N_5619,N_5100,N_5085);
or U5620 (N_5620,N_5155,N_5186);
nor U5621 (N_5621,N_5081,N_5467);
or U5622 (N_5622,N_5149,N_5110);
nor U5623 (N_5623,N_5082,N_5285);
and U5624 (N_5624,N_5217,N_5177);
xnor U5625 (N_5625,N_5222,N_5035);
or U5626 (N_5626,N_5437,N_5474);
nand U5627 (N_5627,N_5176,N_5381);
nor U5628 (N_5628,N_5183,N_5106);
nor U5629 (N_5629,N_5413,N_5352);
xor U5630 (N_5630,N_5326,N_5346);
or U5631 (N_5631,N_5069,N_5018);
nor U5632 (N_5632,N_5064,N_5231);
nand U5633 (N_5633,N_5373,N_5160);
nor U5634 (N_5634,N_5297,N_5320);
or U5635 (N_5635,N_5282,N_5301);
nor U5636 (N_5636,N_5148,N_5283);
nor U5637 (N_5637,N_5068,N_5185);
nand U5638 (N_5638,N_5355,N_5239);
nor U5639 (N_5639,N_5499,N_5416);
nand U5640 (N_5640,N_5252,N_5040);
or U5641 (N_5641,N_5388,N_5245);
or U5642 (N_5642,N_5310,N_5417);
xor U5643 (N_5643,N_5250,N_5215);
nand U5644 (N_5644,N_5171,N_5133);
nand U5645 (N_5645,N_5268,N_5070);
xor U5646 (N_5646,N_5498,N_5336);
nor U5647 (N_5647,N_5151,N_5335);
and U5648 (N_5648,N_5443,N_5098);
xnor U5649 (N_5649,N_5294,N_5227);
nor U5650 (N_5650,N_5479,N_5023);
or U5651 (N_5651,N_5137,N_5423);
xor U5652 (N_5652,N_5487,N_5339);
or U5653 (N_5653,N_5356,N_5147);
and U5654 (N_5654,N_5265,N_5233);
xnor U5655 (N_5655,N_5034,N_5109);
nand U5656 (N_5656,N_5277,N_5414);
or U5657 (N_5657,N_5206,N_5190);
nor U5658 (N_5658,N_5097,N_5004);
and U5659 (N_5659,N_5016,N_5262);
and U5660 (N_5660,N_5152,N_5030);
or U5661 (N_5661,N_5358,N_5453);
nor U5662 (N_5662,N_5103,N_5484);
nand U5663 (N_5663,N_5095,N_5477);
xor U5664 (N_5664,N_5025,N_5248);
nor U5665 (N_5665,N_5084,N_5334);
nand U5666 (N_5666,N_5052,N_5488);
nand U5667 (N_5667,N_5458,N_5165);
nor U5668 (N_5668,N_5404,N_5492);
nor U5669 (N_5669,N_5421,N_5342);
and U5670 (N_5670,N_5017,N_5232);
xnor U5671 (N_5671,N_5296,N_5163);
nor U5672 (N_5672,N_5318,N_5157);
xnor U5673 (N_5673,N_5062,N_5409);
and U5674 (N_5674,N_5435,N_5466);
xor U5675 (N_5675,N_5460,N_5439);
or U5676 (N_5676,N_5111,N_5053);
or U5677 (N_5677,N_5075,N_5096);
and U5678 (N_5678,N_5364,N_5156);
nor U5679 (N_5679,N_5088,N_5168);
nor U5680 (N_5680,N_5089,N_5188);
or U5681 (N_5681,N_5120,N_5379);
and U5682 (N_5682,N_5047,N_5026);
nor U5683 (N_5683,N_5380,N_5347);
nand U5684 (N_5684,N_5179,N_5266);
nor U5685 (N_5685,N_5145,N_5237);
xor U5686 (N_5686,N_5374,N_5480);
nor U5687 (N_5687,N_5267,N_5161);
nor U5688 (N_5688,N_5083,N_5392);
and U5689 (N_5689,N_5331,N_5429);
nand U5690 (N_5690,N_5246,N_5377);
or U5691 (N_5691,N_5312,N_5223);
nand U5692 (N_5692,N_5015,N_5021);
or U5693 (N_5693,N_5345,N_5033);
or U5694 (N_5694,N_5189,N_5348);
or U5695 (N_5695,N_5127,N_5259);
or U5696 (N_5696,N_5390,N_5119);
nand U5697 (N_5697,N_5401,N_5077);
nor U5698 (N_5698,N_5209,N_5196);
nand U5699 (N_5699,N_5293,N_5158);
nand U5700 (N_5700,N_5287,N_5461);
xnor U5701 (N_5701,N_5043,N_5193);
nand U5702 (N_5702,N_5022,N_5225);
nor U5703 (N_5703,N_5170,N_5305);
or U5704 (N_5704,N_5425,N_5337);
nand U5705 (N_5705,N_5431,N_5139);
xnor U5706 (N_5706,N_5105,N_5361);
nand U5707 (N_5707,N_5126,N_5124);
xnor U5708 (N_5708,N_5383,N_5024);
xnor U5709 (N_5709,N_5027,N_5007);
or U5710 (N_5710,N_5243,N_5330);
nand U5711 (N_5711,N_5359,N_5054);
xnor U5712 (N_5712,N_5201,N_5420);
or U5713 (N_5713,N_5180,N_5451);
nand U5714 (N_5714,N_5087,N_5129);
or U5715 (N_5715,N_5260,N_5410);
nand U5716 (N_5716,N_5444,N_5412);
or U5717 (N_5717,N_5462,N_5049);
or U5718 (N_5718,N_5269,N_5384);
nor U5719 (N_5719,N_5427,N_5113);
nand U5720 (N_5720,N_5020,N_5482);
and U5721 (N_5721,N_5307,N_5226);
xnor U5722 (N_5722,N_5029,N_5059);
nor U5723 (N_5723,N_5134,N_5274);
nand U5724 (N_5724,N_5445,N_5387);
or U5725 (N_5725,N_5290,N_5489);
nor U5726 (N_5726,N_5091,N_5197);
xor U5727 (N_5727,N_5415,N_5454);
and U5728 (N_5728,N_5430,N_5468);
nor U5729 (N_5729,N_5313,N_5497);
nand U5730 (N_5730,N_5093,N_5428);
xnor U5731 (N_5731,N_5368,N_5393);
xnor U5732 (N_5732,N_5218,N_5061);
and U5733 (N_5733,N_5143,N_5150);
nand U5734 (N_5734,N_5351,N_5202);
nor U5735 (N_5735,N_5486,N_5251);
nor U5736 (N_5736,N_5003,N_5406);
or U5737 (N_5737,N_5371,N_5014);
nor U5738 (N_5738,N_5446,N_5241);
xor U5739 (N_5739,N_5187,N_5365);
nand U5740 (N_5740,N_5213,N_5450);
or U5741 (N_5741,N_5408,N_5314);
and U5742 (N_5742,N_5182,N_5329);
xnor U5743 (N_5743,N_5418,N_5360);
xor U5744 (N_5744,N_5169,N_5394);
and U5745 (N_5745,N_5199,N_5063);
nor U5746 (N_5746,N_5376,N_5238);
or U5747 (N_5747,N_5236,N_5257);
nand U5748 (N_5748,N_5002,N_5174);
or U5749 (N_5749,N_5066,N_5378);
and U5750 (N_5750,N_5428,N_5256);
nand U5751 (N_5751,N_5127,N_5153);
xnor U5752 (N_5752,N_5157,N_5028);
nor U5753 (N_5753,N_5412,N_5030);
nor U5754 (N_5754,N_5157,N_5378);
xnor U5755 (N_5755,N_5078,N_5436);
and U5756 (N_5756,N_5108,N_5123);
xnor U5757 (N_5757,N_5075,N_5236);
nor U5758 (N_5758,N_5313,N_5240);
and U5759 (N_5759,N_5132,N_5285);
nand U5760 (N_5760,N_5449,N_5013);
xnor U5761 (N_5761,N_5421,N_5000);
nand U5762 (N_5762,N_5103,N_5244);
and U5763 (N_5763,N_5247,N_5152);
xnor U5764 (N_5764,N_5255,N_5367);
nor U5765 (N_5765,N_5275,N_5007);
nand U5766 (N_5766,N_5220,N_5108);
xor U5767 (N_5767,N_5277,N_5418);
or U5768 (N_5768,N_5065,N_5176);
xnor U5769 (N_5769,N_5437,N_5371);
xnor U5770 (N_5770,N_5406,N_5467);
and U5771 (N_5771,N_5443,N_5184);
nand U5772 (N_5772,N_5004,N_5167);
or U5773 (N_5773,N_5449,N_5242);
and U5774 (N_5774,N_5291,N_5267);
xnor U5775 (N_5775,N_5215,N_5411);
and U5776 (N_5776,N_5382,N_5098);
xor U5777 (N_5777,N_5255,N_5265);
and U5778 (N_5778,N_5468,N_5229);
and U5779 (N_5779,N_5203,N_5417);
and U5780 (N_5780,N_5011,N_5204);
and U5781 (N_5781,N_5204,N_5214);
and U5782 (N_5782,N_5278,N_5445);
xor U5783 (N_5783,N_5172,N_5321);
nor U5784 (N_5784,N_5496,N_5120);
and U5785 (N_5785,N_5176,N_5037);
nor U5786 (N_5786,N_5125,N_5194);
nand U5787 (N_5787,N_5450,N_5137);
xor U5788 (N_5788,N_5152,N_5464);
nand U5789 (N_5789,N_5041,N_5442);
or U5790 (N_5790,N_5103,N_5315);
or U5791 (N_5791,N_5119,N_5294);
xnor U5792 (N_5792,N_5370,N_5320);
or U5793 (N_5793,N_5117,N_5339);
nor U5794 (N_5794,N_5319,N_5190);
nand U5795 (N_5795,N_5092,N_5186);
nand U5796 (N_5796,N_5268,N_5458);
or U5797 (N_5797,N_5141,N_5245);
and U5798 (N_5798,N_5086,N_5335);
or U5799 (N_5799,N_5485,N_5197);
xnor U5800 (N_5800,N_5474,N_5032);
or U5801 (N_5801,N_5419,N_5148);
and U5802 (N_5802,N_5002,N_5205);
and U5803 (N_5803,N_5289,N_5266);
xor U5804 (N_5804,N_5399,N_5495);
and U5805 (N_5805,N_5162,N_5223);
nor U5806 (N_5806,N_5401,N_5383);
xnor U5807 (N_5807,N_5370,N_5138);
xnor U5808 (N_5808,N_5381,N_5445);
nand U5809 (N_5809,N_5420,N_5385);
nand U5810 (N_5810,N_5220,N_5205);
xnor U5811 (N_5811,N_5000,N_5133);
or U5812 (N_5812,N_5398,N_5327);
or U5813 (N_5813,N_5024,N_5298);
xnor U5814 (N_5814,N_5015,N_5301);
nor U5815 (N_5815,N_5252,N_5362);
nand U5816 (N_5816,N_5192,N_5024);
and U5817 (N_5817,N_5268,N_5043);
xnor U5818 (N_5818,N_5370,N_5488);
and U5819 (N_5819,N_5281,N_5207);
nor U5820 (N_5820,N_5385,N_5405);
xnor U5821 (N_5821,N_5150,N_5065);
nor U5822 (N_5822,N_5063,N_5252);
nand U5823 (N_5823,N_5326,N_5242);
nor U5824 (N_5824,N_5381,N_5100);
nor U5825 (N_5825,N_5468,N_5098);
or U5826 (N_5826,N_5452,N_5053);
nor U5827 (N_5827,N_5332,N_5367);
nor U5828 (N_5828,N_5233,N_5335);
xor U5829 (N_5829,N_5074,N_5351);
or U5830 (N_5830,N_5487,N_5387);
and U5831 (N_5831,N_5428,N_5386);
and U5832 (N_5832,N_5441,N_5009);
xor U5833 (N_5833,N_5083,N_5081);
nor U5834 (N_5834,N_5076,N_5006);
xor U5835 (N_5835,N_5126,N_5339);
nor U5836 (N_5836,N_5015,N_5173);
xor U5837 (N_5837,N_5462,N_5484);
or U5838 (N_5838,N_5149,N_5165);
or U5839 (N_5839,N_5493,N_5311);
xor U5840 (N_5840,N_5414,N_5029);
or U5841 (N_5841,N_5287,N_5164);
nor U5842 (N_5842,N_5078,N_5034);
or U5843 (N_5843,N_5215,N_5259);
and U5844 (N_5844,N_5141,N_5454);
nor U5845 (N_5845,N_5489,N_5040);
nand U5846 (N_5846,N_5014,N_5325);
nor U5847 (N_5847,N_5499,N_5223);
nor U5848 (N_5848,N_5089,N_5439);
and U5849 (N_5849,N_5470,N_5285);
nand U5850 (N_5850,N_5236,N_5222);
and U5851 (N_5851,N_5308,N_5267);
or U5852 (N_5852,N_5013,N_5398);
nor U5853 (N_5853,N_5385,N_5096);
or U5854 (N_5854,N_5008,N_5243);
nor U5855 (N_5855,N_5070,N_5206);
and U5856 (N_5856,N_5251,N_5408);
nand U5857 (N_5857,N_5149,N_5354);
nand U5858 (N_5858,N_5431,N_5078);
and U5859 (N_5859,N_5127,N_5118);
nand U5860 (N_5860,N_5345,N_5188);
nor U5861 (N_5861,N_5399,N_5267);
and U5862 (N_5862,N_5301,N_5391);
nand U5863 (N_5863,N_5130,N_5223);
or U5864 (N_5864,N_5402,N_5220);
xor U5865 (N_5865,N_5225,N_5344);
or U5866 (N_5866,N_5247,N_5444);
and U5867 (N_5867,N_5195,N_5084);
and U5868 (N_5868,N_5052,N_5334);
xor U5869 (N_5869,N_5005,N_5395);
and U5870 (N_5870,N_5016,N_5476);
or U5871 (N_5871,N_5234,N_5239);
xor U5872 (N_5872,N_5175,N_5480);
nor U5873 (N_5873,N_5180,N_5170);
xor U5874 (N_5874,N_5191,N_5219);
nand U5875 (N_5875,N_5068,N_5348);
nand U5876 (N_5876,N_5271,N_5424);
nand U5877 (N_5877,N_5067,N_5373);
nand U5878 (N_5878,N_5225,N_5338);
or U5879 (N_5879,N_5080,N_5261);
nand U5880 (N_5880,N_5266,N_5151);
xnor U5881 (N_5881,N_5185,N_5241);
nor U5882 (N_5882,N_5188,N_5235);
xnor U5883 (N_5883,N_5463,N_5395);
nor U5884 (N_5884,N_5044,N_5397);
nand U5885 (N_5885,N_5238,N_5145);
nand U5886 (N_5886,N_5047,N_5405);
nor U5887 (N_5887,N_5026,N_5167);
nand U5888 (N_5888,N_5023,N_5021);
or U5889 (N_5889,N_5184,N_5444);
xor U5890 (N_5890,N_5399,N_5037);
xor U5891 (N_5891,N_5378,N_5029);
or U5892 (N_5892,N_5493,N_5259);
nor U5893 (N_5893,N_5148,N_5401);
nand U5894 (N_5894,N_5003,N_5384);
nor U5895 (N_5895,N_5347,N_5238);
nand U5896 (N_5896,N_5165,N_5218);
nand U5897 (N_5897,N_5130,N_5173);
nand U5898 (N_5898,N_5170,N_5274);
nor U5899 (N_5899,N_5492,N_5288);
or U5900 (N_5900,N_5242,N_5441);
nor U5901 (N_5901,N_5361,N_5204);
nand U5902 (N_5902,N_5314,N_5268);
and U5903 (N_5903,N_5483,N_5383);
nand U5904 (N_5904,N_5221,N_5430);
nor U5905 (N_5905,N_5393,N_5238);
and U5906 (N_5906,N_5458,N_5351);
and U5907 (N_5907,N_5000,N_5233);
nand U5908 (N_5908,N_5110,N_5398);
xor U5909 (N_5909,N_5461,N_5064);
xor U5910 (N_5910,N_5469,N_5154);
and U5911 (N_5911,N_5405,N_5298);
or U5912 (N_5912,N_5461,N_5030);
nor U5913 (N_5913,N_5176,N_5079);
nand U5914 (N_5914,N_5110,N_5380);
or U5915 (N_5915,N_5051,N_5314);
or U5916 (N_5916,N_5259,N_5001);
nor U5917 (N_5917,N_5216,N_5040);
or U5918 (N_5918,N_5036,N_5430);
nor U5919 (N_5919,N_5441,N_5244);
xnor U5920 (N_5920,N_5122,N_5060);
and U5921 (N_5921,N_5208,N_5054);
nand U5922 (N_5922,N_5104,N_5157);
and U5923 (N_5923,N_5035,N_5412);
nand U5924 (N_5924,N_5174,N_5183);
nor U5925 (N_5925,N_5437,N_5443);
xor U5926 (N_5926,N_5391,N_5060);
xnor U5927 (N_5927,N_5252,N_5438);
nor U5928 (N_5928,N_5496,N_5207);
and U5929 (N_5929,N_5254,N_5081);
and U5930 (N_5930,N_5106,N_5442);
nor U5931 (N_5931,N_5313,N_5070);
or U5932 (N_5932,N_5187,N_5251);
and U5933 (N_5933,N_5080,N_5039);
nor U5934 (N_5934,N_5471,N_5455);
nor U5935 (N_5935,N_5202,N_5448);
or U5936 (N_5936,N_5337,N_5381);
or U5937 (N_5937,N_5444,N_5123);
nor U5938 (N_5938,N_5411,N_5389);
xor U5939 (N_5939,N_5192,N_5165);
or U5940 (N_5940,N_5330,N_5206);
xnor U5941 (N_5941,N_5473,N_5059);
xor U5942 (N_5942,N_5219,N_5190);
nor U5943 (N_5943,N_5374,N_5034);
xor U5944 (N_5944,N_5137,N_5119);
nor U5945 (N_5945,N_5036,N_5165);
nand U5946 (N_5946,N_5348,N_5387);
nor U5947 (N_5947,N_5257,N_5229);
xnor U5948 (N_5948,N_5408,N_5029);
xnor U5949 (N_5949,N_5400,N_5193);
or U5950 (N_5950,N_5101,N_5356);
nand U5951 (N_5951,N_5298,N_5229);
and U5952 (N_5952,N_5334,N_5420);
nand U5953 (N_5953,N_5120,N_5308);
nand U5954 (N_5954,N_5111,N_5007);
nor U5955 (N_5955,N_5000,N_5079);
and U5956 (N_5956,N_5395,N_5119);
or U5957 (N_5957,N_5113,N_5451);
nor U5958 (N_5958,N_5130,N_5127);
xnor U5959 (N_5959,N_5486,N_5235);
or U5960 (N_5960,N_5454,N_5353);
xor U5961 (N_5961,N_5000,N_5089);
xor U5962 (N_5962,N_5380,N_5004);
nor U5963 (N_5963,N_5388,N_5316);
nor U5964 (N_5964,N_5358,N_5221);
nor U5965 (N_5965,N_5154,N_5122);
xnor U5966 (N_5966,N_5287,N_5194);
xor U5967 (N_5967,N_5331,N_5214);
nand U5968 (N_5968,N_5437,N_5098);
nand U5969 (N_5969,N_5121,N_5421);
and U5970 (N_5970,N_5192,N_5238);
and U5971 (N_5971,N_5145,N_5242);
nand U5972 (N_5972,N_5341,N_5307);
xor U5973 (N_5973,N_5452,N_5319);
and U5974 (N_5974,N_5158,N_5127);
xnor U5975 (N_5975,N_5189,N_5416);
or U5976 (N_5976,N_5110,N_5237);
nand U5977 (N_5977,N_5004,N_5137);
or U5978 (N_5978,N_5257,N_5158);
and U5979 (N_5979,N_5417,N_5070);
nand U5980 (N_5980,N_5342,N_5066);
nand U5981 (N_5981,N_5222,N_5457);
xnor U5982 (N_5982,N_5172,N_5167);
nand U5983 (N_5983,N_5355,N_5035);
nor U5984 (N_5984,N_5042,N_5245);
nand U5985 (N_5985,N_5227,N_5419);
nand U5986 (N_5986,N_5037,N_5078);
nand U5987 (N_5987,N_5310,N_5035);
nor U5988 (N_5988,N_5447,N_5251);
nand U5989 (N_5989,N_5382,N_5049);
nor U5990 (N_5990,N_5446,N_5045);
xor U5991 (N_5991,N_5128,N_5283);
and U5992 (N_5992,N_5189,N_5197);
xnor U5993 (N_5993,N_5225,N_5387);
xnor U5994 (N_5994,N_5373,N_5034);
xnor U5995 (N_5995,N_5183,N_5303);
xor U5996 (N_5996,N_5037,N_5181);
nand U5997 (N_5997,N_5401,N_5229);
and U5998 (N_5998,N_5244,N_5204);
xnor U5999 (N_5999,N_5485,N_5151);
and U6000 (N_6000,N_5817,N_5671);
xnor U6001 (N_6001,N_5723,N_5583);
nand U6002 (N_6002,N_5856,N_5822);
nand U6003 (N_6003,N_5612,N_5806);
and U6004 (N_6004,N_5592,N_5926);
nor U6005 (N_6005,N_5695,N_5974);
and U6006 (N_6006,N_5524,N_5575);
xnor U6007 (N_6007,N_5688,N_5648);
nor U6008 (N_6008,N_5643,N_5746);
and U6009 (N_6009,N_5938,N_5812);
and U6010 (N_6010,N_5752,N_5523);
nor U6011 (N_6011,N_5934,N_5999);
and U6012 (N_6012,N_5841,N_5654);
and U6013 (N_6013,N_5700,N_5620);
xnor U6014 (N_6014,N_5596,N_5534);
nor U6015 (N_6015,N_5814,N_5845);
or U6016 (N_6016,N_5830,N_5565);
xor U6017 (N_6017,N_5674,N_5715);
and U6018 (N_6018,N_5947,N_5662);
and U6019 (N_6019,N_5835,N_5663);
or U6020 (N_6020,N_5811,N_5667);
and U6021 (N_6021,N_5568,N_5740);
and U6022 (N_6022,N_5753,N_5771);
nand U6023 (N_6023,N_5866,N_5658);
nand U6024 (N_6024,N_5800,N_5833);
xnor U6025 (N_6025,N_5943,N_5961);
xor U6026 (N_6026,N_5895,N_5540);
nor U6027 (N_6027,N_5975,N_5980);
or U6028 (N_6028,N_5919,N_5883);
or U6029 (N_6029,N_5921,N_5680);
or U6030 (N_6030,N_5707,N_5692);
nand U6031 (N_6031,N_5726,N_5672);
nor U6032 (N_6032,N_5710,N_5923);
and U6033 (N_6033,N_5815,N_5908);
nor U6034 (N_6034,N_5652,N_5993);
xor U6035 (N_6035,N_5506,N_5511);
nor U6036 (N_6036,N_5874,N_5952);
and U6037 (N_6037,N_5824,N_5623);
xnor U6038 (N_6038,N_5530,N_5887);
and U6039 (N_6039,N_5910,N_5573);
xor U6040 (N_6040,N_5533,N_5584);
nand U6041 (N_6041,N_5765,N_5966);
or U6042 (N_6042,N_5786,N_5608);
xor U6043 (N_6043,N_5985,N_5621);
and U6044 (N_6044,N_5816,N_5642);
nor U6045 (N_6045,N_5760,N_5970);
xnor U6046 (N_6046,N_5732,N_5650);
nand U6047 (N_6047,N_5610,N_5837);
and U6048 (N_6048,N_5702,N_5802);
nand U6049 (N_6049,N_5748,N_5542);
nand U6050 (N_6050,N_5730,N_5510);
or U6051 (N_6051,N_5703,N_5528);
and U6052 (N_6052,N_5950,N_5867);
nand U6053 (N_6053,N_5944,N_5589);
and U6054 (N_6054,N_5544,N_5823);
nor U6055 (N_6055,N_5744,N_5987);
nand U6056 (N_6056,N_5770,N_5706);
and U6057 (N_6057,N_5977,N_5756);
and U6058 (N_6058,N_5601,N_5909);
nand U6059 (N_6059,N_5545,N_5945);
xnor U6060 (N_6060,N_5774,N_5792);
nor U6061 (N_6061,N_5547,N_5881);
nand U6062 (N_6062,N_5701,N_5920);
or U6063 (N_6063,N_5618,N_5720);
nor U6064 (N_6064,N_5858,N_5679);
nor U6065 (N_6065,N_5903,N_5925);
nor U6066 (N_6066,N_5754,N_5588);
and U6067 (N_6067,N_5735,N_5591);
nand U6068 (N_6068,N_5781,N_5935);
xnor U6069 (N_6069,N_5572,N_5724);
nand U6070 (N_6070,N_5803,N_5698);
xnor U6071 (N_6071,N_5846,N_5646);
or U6072 (N_6072,N_5779,N_5940);
or U6073 (N_6073,N_5790,N_5832);
nand U6074 (N_6074,N_5635,N_5791);
and U6075 (N_6075,N_5741,N_5912);
nor U6076 (N_6076,N_5670,N_5870);
nor U6077 (N_6077,N_5683,N_5891);
xnor U6078 (N_6078,N_5687,N_5512);
nand U6079 (N_6079,N_5651,N_5714);
xnor U6080 (N_6080,N_5598,N_5949);
nor U6081 (N_6081,N_5594,N_5902);
nand U6082 (N_6082,N_5820,N_5579);
and U6083 (N_6083,N_5625,N_5882);
and U6084 (N_6084,N_5638,N_5868);
nand U6085 (N_6085,N_5567,N_5622);
xor U6086 (N_6086,N_5969,N_5991);
or U6087 (N_6087,N_5529,N_5930);
nand U6088 (N_6088,N_5556,N_5637);
nor U6089 (N_6089,N_5965,N_5764);
xnor U6090 (N_6090,N_5990,N_5798);
xor U6091 (N_6091,N_5986,N_5879);
nand U6092 (N_6092,N_5761,N_5619);
nand U6093 (N_6093,N_5851,N_5501);
nand U6094 (N_6094,N_5932,N_5963);
or U6095 (N_6095,N_5995,N_5957);
nand U6096 (N_6096,N_5656,N_5745);
and U6097 (N_6097,N_5733,N_5614);
nor U6098 (N_6098,N_5772,N_5927);
or U6099 (N_6099,N_5872,N_5731);
nor U6100 (N_6100,N_5749,N_5853);
nor U6101 (N_6101,N_5628,N_5978);
xor U6102 (N_6102,N_5520,N_5759);
xnor U6103 (N_6103,N_5875,N_5500);
and U6104 (N_6104,N_5829,N_5827);
nand U6105 (N_6105,N_5766,N_5543);
and U6106 (N_6106,N_5526,N_5936);
nand U6107 (N_6107,N_5677,N_5795);
nand U6108 (N_6108,N_5629,N_5782);
xnor U6109 (N_6109,N_5942,N_5600);
nor U6110 (N_6110,N_5560,N_5937);
nand U6111 (N_6111,N_5834,N_5857);
nor U6112 (N_6112,N_5763,N_5862);
nor U6113 (N_6113,N_5804,N_5593);
xor U6114 (N_6114,N_5843,N_5994);
xnor U6115 (N_6115,N_5633,N_5665);
and U6116 (N_6116,N_5787,N_5647);
and U6117 (N_6117,N_5821,N_5988);
or U6118 (N_6118,N_5659,N_5640);
xor U6119 (N_6119,N_5539,N_5813);
and U6120 (N_6120,N_5886,N_5615);
and U6121 (N_6121,N_5900,N_5553);
xnor U6122 (N_6122,N_5634,N_5516);
or U6123 (N_6123,N_5668,N_5924);
or U6124 (N_6124,N_5563,N_5604);
or U6125 (N_6125,N_5639,N_5554);
nor U6126 (N_6126,N_5657,N_5951);
nor U6127 (N_6127,N_5535,N_5768);
nor U6128 (N_6128,N_5527,N_5721);
and U6129 (N_6129,N_5842,N_5848);
nor U6130 (N_6130,N_5799,N_5890);
and U6131 (N_6131,N_5597,N_5916);
and U6132 (N_6132,N_5789,N_5697);
nor U6133 (N_6133,N_5897,N_5775);
or U6134 (N_6134,N_5576,N_5655);
and U6135 (N_6135,N_5718,N_5611);
or U6136 (N_6136,N_5502,N_5836);
nand U6137 (N_6137,N_5508,N_5855);
nor U6138 (N_6138,N_5784,N_5840);
xor U6139 (N_6139,N_5825,N_5645);
nand U6140 (N_6140,N_5631,N_5982);
nor U6141 (N_6141,N_5541,N_5682);
and U6142 (N_6142,N_5580,N_5607);
or U6143 (N_6143,N_5705,N_5546);
and U6144 (N_6144,N_5854,N_5989);
nor U6145 (N_6145,N_5555,N_5630);
xnor U6146 (N_6146,N_5960,N_5661);
nand U6147 (N_6147,N_5953,N_5641);
nand U6148 (N_6148,N_5807,N_5581);
or U6149 (N_6149,N_5616,N_5971);
xnor U6150 (N_6150,N_5939,N_5574);
nand U6151 (N_6151,N_5998,N_5736);
and U6152 (N_6152,N_5847,N_5973);
or U6153 (N_6153,N_5899,N_5976);
and U6154 (N_6154,N_5653,N_5595);
nor U6155 (N_6155,N_5632,N_5801);
and U6156 (N_6156,N_5549,N_5742);
and U6157 (N_6157,N_5561,N_5582);
nor U6158 (N_6158,N_5757,N_5696);
or U6159 (N_6159,N_5933,N_5778);
xnor U6160 (N_6160,N_5562,N_5624);
nand U6161 (N_6161,N_5552,N_5863);
and U6162 (N_6162,N_5959,N_5962);
nor U6163 (N_6163,N_5831,N_5690);
and U6164 (N_6164,N_5922,N_5885);
nor U6165 (N_6165,N_5587,N_5603);
and U6166 (N_6166,N_5805,N_5888);
nor U6167 (N_6167,N_5751,N_5808);
or U6168 (N_6168,N_5901,N_5914);
or U6169 (N_6169,N_5709,N_5536);
and U6170 (N_6170,N_5602,N_5907);
nor U6171 (N_6171,N_5711,N_5954);
xor U6172 (N_6172,N_5776,N_5522);
and U6173 (N_6173,N_5649,N_5956);
xor U6174 (N_6174,N_5505,N_5955);
and U6175 (N_6175,N_5617,N_5996);
and U6176 (N_6176,N_5894,N_5948);
xor U6177 (N_6177,N_5570,N_5983);
nand U6178 (N_6178,N_5518,N_5810);
and U6179 (N_6179,N_5958,N_5551);
nor U6180 (N_6180,N_5917,N_5515);
or U6181 (N_6181,N_5737,N_5712);
nand U6182 (N_6182,N_5839,N_5678);
nand U6183 (N_6183,N_5780,N_5689);
nor U6184 (N_6184,N_5504,N_5613);
xor U6185 (N_6185,N_5738,N_5722);
or U6186 (N_6186,N_5675,N_5627);
xnor U6187 (N_6187,N_5777,N_5968);
or U6188 (N_6188,N_5794,N_5685);
nor U6189 (N_6189,N_5931,N_5519);
xnor U6190 (N_6190,N_5521,N_5704);
and U6191 (N_6191,N_5713,N_5928);
nand U6192 (N_6192,N_5538,N_5739);
xor U6193 (N_6193,N_5869,N_5981);
and U6194 (N_6194,N_5743,N_5758);
xor U6195 (N_6195,N_5513,N_5569);
or U6196 (N_6196,N_5606,N_5979);
and U6197 (N_6197,N_5531,N_5964);
and U6198 (N_6198,N_5509,N_5585);
or U6199 (N_6199,N_5525,N_5826);
and U6200 (N_6200,N_5838,N_5577);
xor U6201 (N_6201,N_5578,N_5664);
or U6202 (N_6202,N_5636,N_5693);
nand U6203 (N_6203,N_5725,N_5913);
or U6204 (N_6204,N_5929,N_5785);
nor U6205 (N_6205,N_5861,N_5666);
nand U6206 (N_6206,N_5676,N_5967);
nor U6207 (N_6207,N_5997,N_5717);
xor U6208 (N_6208,N_5880,N_5892);
and U6209 (N_6209,N_5558,N_5532);
nand U6210 (N_6210,N_5673,N_5972);
nor U6211 (N_6211,N_5694,N_5796);
nand U6212 (N_6212,N_5769,N_5905);
xnor U6213 (N_6213,N_5699,N_5877);
or U6214 (N_6214,N_5889,N_5849);
xnor U6215 (N_6215,N_5818,N_5797);
and U6216 (N_6216,N_5507,N_5884);
or U6217 (N_6217,N_5728,N_5734);
or U6218 (N_6218,N_5762,N_5915);
nor U6219 (N_6219,N_5809,N_5729);
nor U6220 (N_6220,N_5859,N_5871);
or U6221 (N_6221,N_5873,N_5864);
or U6222 (N_6222,N_5590,N_5898);
xor U6223 (N_6223,N_5644,N_5893);
xor U6224 (N_6224,N_5681,N_5605);
nand U6225 (N_6225,N_5686,N_5984);
and U6226 (N_6226,N_5918,N_5550);
xor U6227 (N_6227,N_5852,N_5946);
xor U6228 (N_6228,N_5828,N_5773);
xnor U6229 (N_6229,N_5684,N_5503);
and U6230 (N_6230,N_5911,N_5906);
xor U6231 (N_6231,N_5626,N_5517);
or U6232 (N_6232,N_5719,N_5564);
or U6233 (N_6233,N_5755,N_5819);
nand U6234 (N_6234,N_5865,N_5708);
nor U6235 (N_6235,N_5844,N_5747);
and U6236 (N_6236,N_5548,N_5691);
xnor U6237 (N_6237,N_5941,N_5559);
xor U6238 (N_6238,N_5571,N_5896);
nand U6239 (N_6239,N_5669,N_5850);
or U6240 (N_6240,N_5904,N_5878);
or U6241 (N_6241,N_5727,N_5660);
nor U6242 (N_6242,N_5716,N_5566);
or U6243 (N_6243,N_5876,N_5860);
and U6244 (N_6244,N_5599,N_5750);
xor U6245 (N_6245,N_5537,N_5609);
or U6246 (N_6246,N_5793,N_5783);
and U6247 (N_6247,N_5992,N_5514);
nor U6248 (N_6248,N_5788,N_5767);
nor U6249 (N_6249,N_5586,N_5557);
xnor U6250 (N_6250,N_5823,N_5906);
xor U6251 (N_6251,N_5756,N_5694);
or U6252 (N_6252,N_5738,N_5778);
nand U6253 (N_6253,N_5804,N_5739);
nand U6254 (N_6254,N_5857,N_5604);
or U6255 (N_6255,N_5556,N_5995);
nor U6256 (N_6256,N_5630,N_5664);
nand U6257 (N_6257,N_5611,N_5548);
xnor U6258 (N_6258,N_5793,N_5874);
or U6259 (N_6259,N_5870,N_5619);
nor U6260 (N_6260,N_5873,N_5754);
or U6261 (N_6261,N_5523,N_5806);
or U6262 (N_6262,N_5819,N_5954);
nor U6263 (N_6263,N_5779,N_5735);
xnor U6264 (N_6264,N_5566,N_5723);
xor U6265 (N_6265,N_5640,N_5914);
xnor U6266 (N_6266,N_5578,N_5688);
or U6267 (N_6267,N_5821,N_5958);
nor U6268 (N_6268,N_5536,N_5948);
xor U6269 (N_6269,N_5683,N_5599);
nor U6270 (N_6270,N_5684,N_5699);
nor U6271 (N_6271,N_5598,N_5725);
and U6272 (N_6272,N_5908,N_5698);
or U6273 (N_6273,N_5502,N_5776);
or U6274 (N_6274,N_5525,N_5724);
and U6275 (N_6275,N_5716,N_5626);
and U6276 (N_6276,N_5789,N_5563);
nor U6277 (N_6277,N_5603,N_5685);
nor U6278 (N_6278,N_5767,N_5743);
and U6279 (N_6279,N_5721,N_5596);
or U6280 (N_6280,N_5597,N_5831);
or U6281 (N_6281,N_5635,N_5874);
or U6282 (N_6282,N_5778,N_5524);
nor U6283 (N_6283,N_5620,N_5799);
xnor U6284 (N_6284,N_5965,N_5786);
nand U6285 (N_6285,N_5936,N_5830);
or U6286 (N_6286,N_5928,N_5914);
or U6287 (N_6287,N_5688,N_5526);
xnor U6288 (N_6288,N_5643,N_5977);
or U6289 (N_6289,N_5636,N_5960);
and U6290 (N_6290,N_5504,N_5966);
nor U6291 (N_6291,N_5641,N_5881);
and U6292 (N_6292,N_5631,N_5753);
and U6293 (N_6293,N_5533,N_5961);
xor U6294 (N_6294,N_5817,N_5525);
xnor U6295 (N_6295,N_5757,N_5556);
or U6296 (N_6296,N_5824,N_5662);
nand U6297 (N_6297,N_5688,N_5510);
and U6298 (N_6298,N_5849,N_5960);
or U6299 (N_6299,N_5617,N_5509);
nor U6300 (N_6300,N_5973,N_5758);
nor U6301 (N_6301,N_5726,N_5730);
nand U6302 (N_6302,N_5774,N_5542);
xnor U6303 (N_6303,N_5930,N_5603);
nand U6304 (N_6304,N_5592,N_5933);
or U6305 (N_6305,N_5944,N_5581);
or U6306 (N_6306,N_5708,N_5630);
nand U6307 (N_6307,N_5680,N_5774);
and U6308 (N_6308,N_5887,N_5745);
or U6309 (N_6309,N_5739,N_5728);
and U6310 (N_6310,N_5709,N_5522);
xor U6311 (N_6311,N_5901,N_5636);
nor U6312 (N_6312,N_5673,N_5702);
and U6313 (N_6313,N_5841,N_5692);
nand U6314 (N_6314,N_5796,N_5935);
nor U6315 (N_6315,N_5799,N_5693);
or U6316 (N_6316,N_5742,N_5744);
nand U6317 (N_6317,N_5626,N_5555);
nand U6318 (N_6318,N_5531,N_5579);
xnor U6319 (N_6319,N_5694,N_5907);
nor U6320 (N_6320,N_5551,N_5540);
xnor U6321 (N_6321,N_5910,N_5735);
or U6322 (N_6322,N_5519,N_5602);
nand U6323 (N_6323,N_5547,N_5828);
nand U6324 (N_6324,N_5949,N_5890);
nor U6325 (N_6325,N_5760,N_5642);
or U6326 (N_6326,N_5916,N_5930);
and U6327 (N_6327,N_5896,N_5582);
and U6328 (N_6328,N_5521,N_5979);
xor U6329 (N_6329,N_5529,N_5987);
and U6330 (N_6330,N_5728,N_5664);
nor U6331 (N_6331,N_5516,N_5602);
and U6332 (N_6332,N_5733,N_5937);
nand U6333 (N_6333,N_5805,N_5733);
or U6334 (N_6334,N_5703,N_5537);
or U6335 (N_6335,N_5819,N_5626);
or U6336 (N_6336,N_5671,N_5762);
nand U6337 (N_6337,N_5646,N_5648);
or U6338 (N_6338,N_5716,N_5829);
xnor U6339 (N_6339,N_5801,N_5951);
and U6340 (N_6340,N_5760,N_5814);
or U6341 (N_6341,N_5523,N_5567);
or U6342 (N_6342,N_5684,N_5566);
and U6343 (N_6343,N_5944,N_5675);
nor U6344 (N_6344,N_5984,N_5979);
nor U6345 (N_6345,N_5539,N_5905);
and U6346 (N_6346,N_5573,N_5560);
nor U6347 (N_6347,N_5555,N_5700);
and U6348 (N_6348,N_5573,N_5838);
nor U6349 (N_6349,N_5976,N_5595);
xnor U6350 (N_6350,N_5548,N_5502);
nand U6351 (N_6351,N_5540,N_5822);
and U6352 (N_6352,N_5510,N_5930);
nor U6353 (N_6353,N_5804,N_5709);
nand U6354 (N_6354,N_5872,N_5973);
nor U6355 (N_6355,N_5901,N_5945);
or U6356 (N_6356,N_5552,N_5880);
nand U6357 (N_6357,N_5641,N_5949);
and U6358 (N_6358,N_5920,N_5667);
nor U6359 (N_6359,N_5628,N_5653);
xor U6360 (N_6360,N_5694,N_5636);
or U6361 (N_6361,N_5973,N_5884);
xnor U6362 (N_6362,N_5883,N_5655);
nor U6363 (N_6363,N_5662,N_5635);
xor U6364 (N_6364,N_5516,N_5984);
nor U6365 (N_6365,N_5758,N_5789);
nand U6366 (N_6366,N_5646,N_5739);
and U6367 (N_6367,N_5549,N_5655);
nand U6368 (N_6368,N_5770,N_5831);
nand U6369 (N_6369,N_5536,N_5570);
nand U6370 (N_6370,N_5639,N_5918);
nor U6371 (N_6371,N_5758,N_5672);
and U6372 (N_6372,N_5948,N_5607);
nor U6373 (N_6373,N_5501,N_5520);
and U6374 (N_6374,N_5651,N_5947);
and U6375 (N_6375,N_5941,N_5874);
nor U6376 (N_6376,N_5681,N_5851);
and U6377 (N_6377,N_5884,N_5584);
xnor U6378 (N_6378,N_5773,N_5734);
xor U6379 (N_6379,N_5522,N_5824);
nand U6380 (N_6380,N_5797,N_5743);
nand U6381 (N_6381,N_5904,N_5560);
nand U6382 (N_6382,N_5895,N_5920);
nor U6383 (N_6383,N_5956,N_5569);
nor U6384 (N_6384,N_5759,N_5911);
nand U6385 (N_6385,N_5853,N_5866);
nor U6386 (N_6386,N_5833,N_5958);
xnor U6387 (N_6387,N_5937,N_5643);
nand U6388 (N_6388,N_5553,N_5954);
nor U6389 (N_6389,N_5956,N_5708);
or U6390 (N_6390,N_5874,N_5542);
nand U6391 (N_6391,N_5559,N_5567);
nor U6392 (N_6392,N_5604,N_5635);
or U6393 (N_6393,N_5834,N_5508);
xnor U6394 (N_6394,N_5664,N_5994);
nor U6395 (N_6395,N_5942,N_5667);
or U6396 (N_6396,N_5595,N_5820);
nor U6397 (N_6397,N_5592,N_5988);
nand U6398 (N_6398,N_5590,N_5800);
nand U6399 (N_6399,N_5893,N_5972);
and U6400 (N_6400,N_5951,N_5552);
and U6401 (N_6401,N_5796,N_5756);
xnor U6402 (N_6402,N_5672,N_5633);
nand U6403 (N_6403,N_5686,N_5820);
nand U6404 (N_6404,N_5552,N_5881);
or U6405 (N_6405,N_5991,N_5977);
and U6406 (N_6406,N_5922,N_5704);
or U6407 (N_6407,N_5545,N_5674);
and U6408 (N_6408,N_5926,N_5766);
and U6409 (N_6409,N_5912,N_5933);
or U6410 (N_6410,N_5913,N_5558);
nand U6411 (N_6411,N_5872,N_5816);
or U6412 (N_6412,N_5545,N_5629);
or U6413 (N_6413,N_5594,N_5654);
xnor U6414 (N_6414,N_5888,N_5997);
and U6415 (N_6415,N_5898,N_5654);
xnor U6416 (N_6416,N_5677,N_5534);
nand U6417 (N_6417,N_5801,N_5982);
nor U6418 (N_6418,N_5850,N_5769);
and U6419 (N_6419,N_5726,N_5892);
and U6420 (N_6420,N_5650,N_5932);
xnor U6421 (N_6421,N_5864,N_5559);
nand U6422 (N_6422,N_5732,N_5793);
nand U6423 (N_6423,N_5759,N_5819);
xor U6424 (N_6424,N_5590,N_5882);
and U6425 (N_6425,N_5550,N_5815);
nand U6426 (N_6426,N_5665,N_5628);
xnor U6427 (N_6427,N_5819,N_5851);
nor U6428 (N_6428,N_5986,N_5691);
nor U6429 (N_6429,N_5721,N_5600);
and U6430 (N_6430,N_5556,N_5833);
or U6431 (N_6431,N_5516,N_5734);
and U6432 (N_6432,N_5907,N_5932);
nor U6433 (N_6433,N_5699,N_5840);
and U6434 (N_6434,N_5654,N_5552);
and U6435 (N_6435,N_5617,N_5854);
and U6436 (N_6436,N_5802,N_5805);
or U6437 (N_6437,N_5930,N_5751);
or U6438 (N_6438,N_5966,N_5977);
nand U6439 (N_6439,N_5986,N_5642);
or U6440 (N_6440,N_5656,N_5520);
or U6441 (N_6441,N_5619,N_5503);
and U6442 (N_6442,N_5719,N_5918);
nor U6443 (N_6443,N_5719,N_5601);
nor U6444 (N_6444,N_5500,N_5879);
or U6445 (N_6445,N_5947,N_5904);
nand U6446 (N_6446,N_5902,N_5892);
xor U6447 (N_6447,N_5502,N_5503);
xnor U6448 (N_6448,N_5727,N_5797);
nand U6449 (N_6449,N_5723,N_5643);
or U6450 (N_6450,N_5630,N_5789);
nor U6451 (N_6451,N_5791,N_5510);
xnor U6452 (N_6452,N_5707,N_5718);
nand U6453 (N_6453,N_5617,N_5755);
nor U6454 (N_6454,N_5901,N_5622);
xnor U6455 (N_6455,N_5939,N_5777);
nand U6456 (N_6456,N_5989,N_5686);
xor U6457 (N_6457,N_5878,N_5892);
nor U6458 (N_6458,N_5623,N_5759);
and U6459 (N_6459,N_5569,N_5880);
nand U6460 (N_6460,N_5565,N_5940);
or U6461 (N_6461,N_5506,N_5515);
xor U6462 (N_6462,N_5959,N_5723);
or U6463 (N_6463,N_5989,N_5555);
nor U6464 (N_6464,N_5952,N_5766);
or U6465 (N_6465,N_5915,N_5927);
nand U6466 (N_6466,N_5886,N_5566);
xor U6467 (N_6467,N_5665,N_5923);
or U6468 (N_6468,N_5930,N_5600);
or U6469 (N_6469,N_5710,N_5692);
xor U6470 (N_6470,N_5783,N_5554);
and U6471 (N_6471,N_5966,N_5641);
nor U6472 (N_6472,N_5720,N_5896);
nand U6473 (N_6473,N_5763,N_5904);
and U6474 (N_6474,N_5785,N_5790);
or U6475 (N_6475,N_5968,N_5536);
xnor U6476 (N_6476,N_5563,N_5943);
or U6477 (N_6477,N_5620,N_5704);
or U6478 (N_6478,N_5546,N_5518);
nor U6479 (N_6479,N_5676,N_5810);
xor U6480 (N_6480,N_5695,N_5977);
nor U6481 (N_6481,N_5615,N_5747);
nor U6482 (N_6482,N_5552,N_5539);
and U6483 (N_6483,N_5886,N_5646);
or U6484 (N_6484,N_5585,N_5925);
and U6485 (N_6485,N_5512,N_5752);
nand U6486 (N_6486,N_5770,N_5581);
xor U6487 (N_6487,N_5864,N_5694);
nand U6488 (N_6488,N_5610,N_5761);
or U6489 (N_6489,N_5557,N_5966);
nand U6490 (N_6490,N_5863,N_5930);
and U6491 (N_6491,N_5797,N_5772);
or U6492 (N_6492,N_5601,N_5875);
nor U6493 (N_6493,N_5838,N_5724);
xnor U6494 (N_6494,N_5905,N_5847);
xnor U6495 (N_6495,N_5952,N_5771);
or U6496 (N_6496,N_5671,N_5981);
or U6497 (N_6497,N_5834,N_5574);
and U6498 (N_6498,N_5759,N_5996);
xnor U6499 (N_6499,N_5807,N_5555);
nor U6500 (N_6500,N_6299,N_6077);
or U6501 (N_6501,N_6270,N_6252);
and U6502 (N_6502,N_6263,N_6044);
or U6503 (N_6503,N_6100,N_6303);
xnor U6504 (N_6504,N_6045,N_6080);
and U6505 (N_6505,N_6250,N_6215);
and U6506 (N_6506,N_6223,N_6282);
or U6507 (N_6507,N_6142,N_6338);
or U6508 (N_6508,N_6022,N_6095);
nor U6509 (N_6509,N_6257,N_6278);
xnor U6510 (N_6510,N_6403,N_6144);
nor U6511 (N_6511,N_6297,N_6108);
xor U6512 (N_6512,N_6378,N_6047);
xor U6513 (N_6513,N_6099,N_6068);
and U6514 (N_6514,N_6391,N_6242);
or U6515 (N_6515,N_6477,N_6206);
and U6516 (N_6516,N_6186,N_6380);
and U6517 (N_6517,N_6332,N_6353);
and U6518 (N_6518,N_6266,N_6154);
and U6519 (N_6519,N_6057,N_6133);
nand U6520 (N_6520,N_6482,N_6447);
nor U6521 (N_6521,N_6193,N_6180);
xnor U6522 (N_6522,N_6205,N_6480);
and U6523 (N_6523,N_6341,N_6114);
nand U6524 (N_6524,N_6283,N_6470);
nand U6525 (N_6525,N_6286,N_6440);
nand U6526 (N_6526,N_6487,N_6295);
xnor U6527 (N_6527,N_6468,N_6217);
or U6528 (N_6528,N_6127,N_6402);
or U6529 (N_6529,N_6106,N_6085);
and U6530 (N_6530,N_6056,N_6113);
nand U6531 (N_6531,N_6156,N_6420);
and U6532 (N_6532,N_6126,N_6195);
or U6533 (N_6533,N_6018,N_6107);
nor U6534 (N_6534,N_6445,N_6102);
and U6535 (N_6535,N_6296,N_6393);
nand U6536 (N_6536,N_6368,N_6419);
or U6537 (N_6537,N_6494,N_6039);
nor U6538 (N_6538,N_6356,N_6199);
nand U6539 (N_6539,N_6227,N_6359);
and U6540 (N_6540,N_6115,N_6162);
nand U6541 (N_6541,N_6231,N_6149);
and U6542 (N_6542,N_6153,N_6130);
xnor U6543 (N_6543,N_6422,N_6082);
nor U6544 (N_6544,N_6170,N_6169);
nor U6545 (N_6545,N_6331,N_6435);
or U6546 (N_6546,N_6458,N_6481);
or U6547 (N_6547,N_6302,N_6221);
and U6548 (N_6548,N_6112,N_6473);
nor U6549 (N_6549,N_6009,N_6198);
xor U6550 (N_6550,N_6386,N_6049);
xnor U6551 (N_6551,N_6012,N_6456);
xor U6552 (N_6552,N_6497,N_6328);
or U6553 (N_6553,N_6385,N_6088);
nor U6554 (N_6554,N_6475,N_6004);
and U6555 (N_6555,N_6405,N_6204);
or U6556 (N_6556,N_6086,N_6267);
or U6557 (N_6557,N_6429,N_6061);
xnor U6558 (N_6558,N_6213,N_6432);
nand U6559 (N_6559,N_6312,N_6421);
and U6560 (N_6560,N_6373,N_6364);
nand U6561 (N_6561,N_6463,N_6390);
or U6562 (N_6562,N_6157,N_6003);
and U6563 (N_6563,N_6005,N_6471);
and U6564 (N_6564,N_6054,N_6074);
xnor U6565 (N_6565,N_6076,N_6277);
nand U6566 (N_6566,N_6182,N_6036);
and U6567 (N_6567,N_6374,N_6308);
nor U6568 (N_6568,N_6145,N_6179);
and U6569 (N_6569,N_6090,N_6249);
nand U6570 (N_6570,N_6272,N_6339);
or U6571 (N_6571,N_6098,N_6330);
nand U6572 (N_6572,N_6094,N_6219);
nor U6573 (N_6573,N_6132,N_6027);
xnor U6574 (N_6574,N_6316,N_6306);
or U6575 (N_6575,N_6140,N_6174);
and U6576 (N_6576,N_6387,N_6459);
and U6577 (N_6577,N_6218,N_6412);
and U6578 (N_6578,N_6448,N_6041);
or U6579 (N_6579,N_6097,N_6253);
and U6580 (N_6580,N_6371,N_6237);
nand U6581 (N_6581,N_6315,N_6268);
and U6582 (N_6582,N_6243,N_6318);
nand U6583 (N_6583,N_6409,N_6222);
nand U6584 (N_6584,N_6093,N_6210);
nand U6585 (N_6585,N_6189,N_6415);
and U6586 (N_6586,N_6065,N_6240);
xnor U6587 (N_6587,N_6388,N_6216);
nand U6588 (N_6588,N_6187,N_6247);
and U6589 (N_6589,N_6214,N_6367);
nand U6590 (N_6590,N_6234,N_6369);
xor U6591 (N_6591,N_6400,N_6064);
xor U6592 (N_6592,N_6490,N_6260);
nand U6593 (N_6593,N_6319,N_6478);
nor U6594 (N_6594,N_6434,N_6079);
and U6595 (N_6595,N_6376,N_6089);
nor U6596 (N_6596,N_6399,N_6357);
or U6597 (N_6597,N_6418,N_6483);
or U6598 (N_6598,N_6406,N_6466);
and U6599 (N_6599,N_6229,N_6361);
and U6600 (N_6600,N_6123,N_6486);
nand U6601 (N_6601,N_6016,N_6492);
or U6602 (N_6602,N_6336,N_6460);
xor U6603 (N_6603,N_6439,N_6105);
nor U6604 (N_6604,N_6209,N_6427);
nand U6605 (N_6605,N_6067,N_6398);
nor U6606 (N_6606,N_6158,N_6462);
and U6607 (N_6607,N_6350,N_6124);
nand U6608 (N_6608,N_6042,N_6334);
xor U6609 (N_6609,N_6053,N_6287);
xor U6610 (N_6610,N_6347,N_6352);
or U6611 (N_6611,N_6200,N_6069);
nand U6612 (N_6612,N_6175,N_6191);
nand U6613 (N_6613,N_6037,N_6355);
or U6614 (N_6614,N_6379,N_6034);
xnor U6615 (N_6615,N_6254,N_6464);
nor U6616 (N_6616,N_6327,N_6280);
and U6617 (N_6617,N_6203,N_6220);
and U6618 (N_6618,N_6394,N_6437);
nor U6619 (N_6619,N_6117,N_6116);
and U6620 (N_6620,N_6208,N_6461);
or U6621 (N_6621,N_6194,N_6196);
or U6622 (N_6622,N_6011,N_6424);
xor U6623 (N_6623,N_6058,N_6015);
nand U6624 (N_6624,N_6111,N_6317);
nand U6625 (N_6625,N_6185,N_6021);
or U6626 (N_6626,N_6395,N_6178);
xor U6627 (N_6627,N_6438,N_6101);
nand U6628 (N_6628,N_6363,N_6091);
nor U6629 (N_6629,N_6281,N_6006);
nand U6630 (N_6630,N_6232,N_6171);
xnor U6631 (N_6631,N_6365,N_6488);
nand U6632 (N_6632,N_6344,N_6024);
nor U6633 (N_6633,N_6320,N_6071);
xnor U6634 (N_6634,N_6259,N_6323);
nor U6635 (N_6635,N_6279,N_6288);
nor U6636 (N_6636,N_6310,N_6078);
nand U6637 (N_6637,N_6120,N_6301);
nor U6638 (N_6638,N_6150,N_6161);
nor U6639 (N_6639,N_6321,N_6104);
or U6640 (N_6640,N_6062,N_6165);
xor U6641 (N_6641,N_6014,N_6444);
and U6642 (N_6642,N_6177,N_6164);
and U6643 (N_6643,N_6329,N_6264);
and U6644 (N_6644,N_6383,N_6059);
or U6645 (N_6645,N_6426,N_6228);
or U6646 (N_6646,N_6457,N_6366);
nor U6647 (N_6647,N_6465,N_6026);
nand U6648 (N_6648,N_6294,N_6305);
and U6649 (N_6649,N_6256,N_6343);
or U6650 (N_6650,N_6147,N_6455);
nand U6651 (N_6651,N_6430,N_6322);
or U6652 (N_6652,N_6119,N_6493);
nor U6653 (N_6653,N_6392,N_6087);
and U6654 (N_6654,N_6413,N_6075);
and U6655 (N_6655,N_6030,N_6007);
nor U6656 (N_6656,N_6275,N_6351);
xnor U6657 (N_6657,N_6137,N_6212);
nor U6658 (N_6658,N_6246,N_6129);
nand U6659 (N_6659,N_6372,N_6146);
xnor U6660 (N_6660,N_6349,N_6184);
and U6661 (N_6661,N_6000,N_6375);
nand U6662 (N_6662,N_6188,N_6143);
nor U6663 (N_6663,N_6135,N_6055);
or U6664 (N_6664,N_6125,N_6051);
nand U6665 (N_6665,N_6013,N_6410);
xor U6666 (N_6666,N_6168,N_6211);
xor U6667 (N_6667,N_6407,N_6019);
nor U6668 (N_6668,N_6397,N_6038);
xnor U6669 (N_6669,N_6314,N_6224);
or U6670 (N_6670,N_6225,N_6273);
nor U6671 (N_6671,N_6148,N_6167);
nor U6672 (N_6672,N_6443,N_6333);
nand U6673 (N_6673,N_6284,N_6384);
nand U6674 (N_6674,N_6241,N_6300);
nand U6675 (N_6675,N_6202,N_6335);
nor U6676 (N_6676,N_6324,N_6382);
nand U6677 (N_6677,N_6173,N_6110);
nand U6678 (N_6678,N_6425,N_6431);
nor U6679 (N_6679,N_6311,N_6121);
and U6680 (N_6680,N_6269,N_6244);
and U6681 (N_6681,N_6498,N_6166);
nor U6682 (N_6682,N_6118,N_6495);
nand U6683 (N_6683,N_6416,N_6411);
xnor U6684 (N_6684,N_6485,N_6313);
nor U6685 (N_6685,N_6274,N_6201);
nand U6686 (N_6686,N_6136,N_6131);
xor U6687 (N_6687,N_6002,N_6096);
nand U6688 (N_6688,N_6360,N_6060);
and U6689 (N_6689,N_6446,N_6103);
nor U6690 (N_6690,N_6290,N_6479);
or U6691 (N_6691,N_6370,N_6176);
nand U6692 (N_6692,N_6307,N_6235);
xnor U6693 (N_6693,N_6381,N_6428);
nor U6694 (N_6694,N_6404,N_6417);
nor U6695 (N_6695,N_6238,N_6046);
nand U6696 (N_6696,N_6160,N_6337);
xnor U6697 (N_6697,N_6489,N_6325);
or U6698 (N_6698,N_6134,N_6377);
nand U6699 (N_6699,N_6197,N_6010);
nand U6700 (N_6700,N_6304,N_6251);
nor U6701 (N_6701,N_6261,N_6052);
or U6702 (N_6702,N_6081,N_6255);
nor U6703 (N_6703,N_6025,N_6396);
nand U6704 (N_6704,N_6138,N_6192);
nor U6705 (N_6705,N_6023,N_6122);
nand U6706 (N_6706,N_6362,N_6342);
nor U6707 (N_6707,N_6233,N_6032);
and U6708 (N_6708,N_6230,N_6291);
nor U6709 (N_6709,N_6072,N_6159);
and U6710 (N_6710,N_6063,N_6345);
nor U6711 (N_6711,N_6070,N_6474);
nand U6712 (N_6712,N_6151,N_6066);
nand U6713 (N_6713,N_6020,N_6028);
xnor U6714 (N_6714,N_6358,N_6083);
or U6715 (N_6715,N_6484,N_6155);
and U6716 (N_6716,N_6190,N_6472);
or U6717 (N_6717,N_6245,N_6401);
nand U6718 (N_6718,N_6207,N_6181);
xor U6719 (N_6719,N_6348,N_6340);
or U6720 (N_6720,N_6248,N_6262);
or U6721 (N_6721,N_6423,N_6452);
and U6722 (N_6722,N_6499,N_6084);
and U6723 (N_6723,N_6109,N_6271);
xnor U6724 (N_6724,N_6141,N_6265);
or U6725 (N_6725,N_6226,N_6408);
nand U6726 (N_6726,N_6496,N_6029);
and U6727 (N_6727,N_6276,N_6043);
and U6728 (N_6728,N_6442,N_6449);
or U6729 (N_6729,N_6048,N_6389);
nand U6730 (N_6730,N_6128,N_6469);
or U6731 (N_6731,N_6326,N_6258);
xnor U6732 (N_6732,N_6451,N_6040);
and U6733 (N_6733,N_6454,N_6354);
or U6734 (N_6734,N_6172,N_6017);
or U6735 (N_6735,N_6285,N_6163);
or U6736 (N_6736,N_6033,N_6139);
and U6737 (N_6737,N_6298,N_6073);
nor U6738 (N_6738,N_6491,N_6236);
nor U6739 (N_6739,N_6441,N_6183);
nand U6740 (N_6740,N_6239,N_6309);
or U6741 (N_6741,N_6008,N_6001);
and U6742 (N_6742,N_6453,N_6433);
and U6743 (N_6743,N_6436,N_6450);
xor U6744 (N_6744,N_6031,N_6467);
nand U6745 (N_6745,N_6035,N_6293);
nand U6746 (N_6746,N_6092,N_6292);
or U6747 (N_6747,N_6476,N_6050);
nand U6748 (N_6748,N_6414,N_6289);
nand U6749 (N_6749,N_6346,N_6152);
xor U6750 (N_6750,N_6358,N_6316);
xnor U6751 (N_6751,N_6261,N_6282);
and U6752 (N_6752,N_6039,N_6004);
nand U6753 (N_6753,N_6272,N_6449);
and U6754 (N_6754,N_6313,N_6486);
nand U6755 (N_6755,N_6479,N_6052);
nand U6756 (N_6756,N_6498,N_6007);
xor U6757 (N_6757,N_6379,N_6112);
xnor U6758 (N_6758,N_6034,N_6410);
xnor U6759 (N_6759,N_6067,N_6369);
or U6760 (N_6760,N_6130,N_6134);
and U6761 (N_6761,N_6348,N_6213);
nor U6762 (N_6762,N_6220,N_6484);
or U6763 (N_6763,N_6469,N_6345);
and U6764 (N_6764,N_6386,N_6200);
nor U6765 (N_6765,N_6304,N_6100);
nor U6766 (N_6766,N_6193,N_6086);
xnor U6767 (N_6767,N_6025,N_6265);
nand U6768 (N_6768,N_6030,N_6101);
nor U6769 (N_6769,N_6172,N_6115);
xnor U6770 (N_6770,N_6194,N_6065);
nor U6771 (N_6771,N_6324,N_6449);
or U6772 (N_6772,N_6433,N_6028);
nand U6773 (N_6773,N_6438,N_6057);
xor U6774 (N_6774,N_6101,N_6183);
or U6775 (N_6775,N_6199,N_6409);
or U6776 (N_6776,N_6456,N_6465);
and U6777 (N_6777,N_6197,N_6438);
and U6778 (N_6778,N_6104,N_6050);
and U6779 (N_6779,N_6294,N_6303);
xor U6780 (N_6780,N_6033,N_6268);
nand U6781 (N_6781,N_6384,N_6430);
xnor U6782 (N_6782,N_6077,N_6006);
nor U6783 (N_6783,N_6280,N_6144);
xnor U6784 (N_6784,N_6016,N_6143);
nor U6785 (N_6785,N_6171,N_6389);
nand U6786 (N_6786,N_6130,N_6254);
nor U6787 (N_6787,N_6121,N_6119);
nand U6788 (N_6788,N_6395,N_6237);
or U6789 (N_6789,N_6496,N_6380);
and U6790 (N_6790,N_6494,N_6291);
and U6791 (N_6791,N_6132,N_6203);
xnor U6792 (N_6792,N_6232,N_6158);
and U6793 (N_6793,N_6034,N_6299);
or U6794 (N_6794,N_6147,N_6038);
and U6795 (N_6795,N_6402,N_6079);
nor U6796 (N_6796,N_6033,N_6280);
and U6797 (N_6797,N_6078,N_6393);
and U6798 (N_6798,N_6005,N_6219);
nor U6799 (N_6799,N_6010,N_6049);
xor U6800 (N_6800,N_6224,N_6494);
or U6801 (N_6801,N_6226,N_6152);
nand U6802 (N_6802,N_6055,N_6326);
nor U6803 (N_6803,N_6336,N_6251);
nand U6804 (N_6804,N_6330,N_6039);
and U6805 (N_6805,N_6132,N_6106);
nand U6806 (N_6806,N_6267,N_6266);
nand U6807 (N_6807,N_6487,N_6371);
nand U6808 (N_6808,N_6177,N_6356);
nor U6809 (N_6809,N_6216,N_6162);
nand U6810 (N_6810,N_6410,N_6012);
xor U6811 (N_6811,N_6498,N_6297);
or U6812 (N_6812,N_6093,N_6056);
xor U6813 (N_6813,N_6374,N_6124);
nor U6814 (N_6814,N_6351,N_6044);
nand U6815 (N_6815,N_6323,N_6320);
and U6816 (N_6816,N_6441,N_6292);
or U6817 (N_6817,N_6419,N_6420);
nor U6818 (N_6818,N_6142,N_6375);
xor U6819 (N_6819,N_6298,N_6280);
nand U6820 (N_6820,N_6048,N_6384);
xor U6821 (N_6821,N_6227,N_6264);
xor U6822 (N_6822,N_6404,N_6393);
nor U6823 (N_6823,N_6272,N_6214);
and U6824 (N_6824,N_6135,N_6480);
and U6825 (N_6825,N_6383,N_6031);
xor U6826 (N_6826,N_6155,N_6397);
xnor U6827 (N_6827,N_6252,N_6033);
nor U6828 (N_6828,N_6473,N_6302);
or U6829 (N_6829,N_6399,N_6460);
and U6830 (N_6830,N_6426,N_6282);
and U6831 (N_6831,N_6108,N_6229);
nand U6832 (N_6832,N_6072,N_6280);
xor U6833 (N_6833,N_6174,N_6405);
nand U6834 (N_6834,N_6048,N_6237);
nor U6835 (N_6835,N_6156,N_6208);
nand U6836 (N_6836,N_6156,N_6151);
and U6837 (N_6837,N_6276,N_6460);
nor U6838 (N_6838,N_6066,N_6180);
nor U6839 (N_6839,N_6206,N_6486);
nor U6840 (N_6840,N_6070,N_6259);
nand U6841 (N_6841,N_6162,N_6339);
nand U6842 (N_6842,N_6069,N_6407);
or U6843 (N_6843,N_6009,N_6374);
xnor U6844 (N_6844,N_6086,N_6324);
or U6845 (N_6845,N_6346,N_6052);
nor U6846 (N_6846,N_6115,N_6306);
or U6847 (N_6847,N_6269,N_6290);
nor U6848 (N_6848,N_6021,N_6365);
and U6849 (N_6849,N_6491,N_6419);
nor U6850 (N_6850,N_6293,N_6019);
nor U6851 (N_6851,N_6290,N_6179);
xnor U6852 (N_6852,N_6189,N_6482);
nand U6853 (N_6853,N_6119,N_6220);
and U6854 (N_6854,N_6395,N_6390);
or U6855 (N_6855,N_6420,N_6198);
nor U6856 (N_6856,N_6276,N_6289);
nor U6857 (N_6857,N_6435,N_6482);
nor U6858 (N_6858,N_6095,N_6341);
and U6859 (N_6859,N_6336,N_6467);
nand U6860 (N_6860,N_6427,N_6491);
and U6861 (N_6861,N_6166,N_6234);
or U6862 (N_6862,N_6310,N_6245);
and U6863 (N_6863,N_6037,N_6142);
and U6864 (N_6864,N_6022,N_6092);
or U6865 (N_6865,N_6443,N_6257);
and U6866 (N_6866,N_6069,N_6218);
nor U6867 (N_6867,N_6067,N_6294);
nor U6868 (N_6868,N_6096,N_6391);
xor U6869 (N_6869,N_6013,N_6469);
nor U6870 (N_6870,N_6448,N_6129);
xnor U6871 (N_6871,N_6036,N_6210);
nand U6872 (N_6872,N_6047,N_6366);
and U6873 (N_6873,N_6468,N_6321);
nor U6874 (N_6874,N_6229,N_6104);
nand U6875 (N_6875,N_6014,N_6004);
nor U6876 (N_6876,N_6055,N_6295);
nand U6877 (N_6877,N_6287,N_6126);
and U6878 (N_6878,N_6357,N_6106);
and U6879 (N_6879,N_6017,N_6054);
nand U6880 (N_6880,N_6090,N_6328);
nor U6881 (N_6881,N_6022,N_6260);
or U6882 (N_6882,N_6322,N_6226);
nand U6883 (N_6883,N_6433,N_6422);
and U6884 (N_6884,N_6495,N_6012);
nand U6885 (N_6885,N_6408,N_6420);
nor U6886 (N_6886,N_6163,N_6080);
nor U6887 (N_6887,N_6252,N_6290);
nand U6888 (N_6888,N_6313,N_6095);
or U6889 (N_6889,N_6364,N_6187);
or U6890 (N_6890,N_6201,N_6289);
nor U6891 (N_6891,N_6342,N_6340);
nor U6892 (N_6892,N_6016,N_6352);
xnor U6893 (N_6893,N_6119,N_6171);
nor U6894 (N_6894,N_6435,N_6277);
xor U6895 (N_6895,N_6322,N_6158);
or U6896 (N_6896,N_6221,N_6035);
nor U6897 (N_6897,N_6129,N_6284);
and U6898 (N_6898,N_6050,N_6063);
nor U6899 (N_6899,N_6327,N_6054);
nand U6900 (N_6900,N_6497,N_6041);
or U6901 (N_6901,N_6091,N_6008);
or U6902 (N_6902,N_6061,N_6425);
xor U6903 (N_6903,N_6122,N_6141);
nor U6904 (N_6904,N_6409,N_6251);
nor U6905 (N_6905,N_6057,N_6169);
nand U6906 (N_6906,N_6193,N_6035);
nor U6907 (N_6907,N_6285,N_6202);
nand U6908 (N_6908,N_6287,N_6276);
nor U6909 (N_6909,N_6418,N_6134);
nand U6910 (N_6910,N_6449,N_6068);
or U6911 (N_6911,N_6198,N_6048);
nand U6912 (N_6912,N_6029,N_6451);
or U6913 (N_6913,N_6263,N_6231);
or U6914 (N_6914,N_6087,N_6083);
nand U6915 (N_6915,N_6054,N_6407);
nor U6916 (N_6916,N_6162,N_6080);
nor U6917 (N_6917,N_6333,N_6497);
nor U6918 (N_6918,N_6124,N_6178);
nand U6919 (N_6919,N_6148,N_6233);
or U6920 (N_6920,N_6456,N_6441);
nor U6921 (N_6921,N_6324,N_6107);
nor U6922 (N_6922,N_6428,N_6072);
or U6923 (N_6923,N_6147,N_6317);
xnor U6924 (N_6924,N_6108,N_6285);
nand U6925 (N_6925,N_6285,N_6169);
or U6926 (N_6926,N_6141,N_6419);
nand U6927 (N_6927,N_6231,N_6492);
and U6928 (N_6928,N_6393,N_6450);
nand U6929 (N_6929,N_6232,N_6019);
or U6930 (N_6930,N_6223,N_6398);
xnor U6931 (N_6931,N_6373,N_6415);
xor U6932 (N_6932,N_6221,N_6099);
and U6933 (N_6933,N_6479,N_6387);
xnor U6934 (N_6934,N_6302,N_6016);
nand U6935 (N_6935,N_6114,N_6382);
xor U6936 (N_6936,N_6176,N_6337);
nor U6937 (N_6937,N_6057,N_6232);
and U6938 (N_6938,N_6156,N_6458);
xor U6939 (N_6939,N_6478,N_6450);
nor U6940 (N_6940,N_6208,N_6333);
or U6941 (N_6941,N_6242,N_6299);
nand U6942 (N_6942,N_6246,N_6397);
nand U6943 (N_6943,N_6400,N_6355);
nor U6944 (N_6944,N_6018,N_6192);
and U6945 (N_6945,N_6016,N_6408);
or U6946 (N_6946,N_6116,N_6363);
or U6947 (N_6947,N_6433,N_6326);
and U6948 (N_6948,N_6259,N_6247);
nand U6949 (N_6949,N_6410,N_6141);
nand U6950 (N_6950,N_6103,N_6012);
xor U6951 (N_6951,N_6262,N_6446);
and U6952 (N_6952,N_6091,N_6493);
and U6953 (N_6953,N_6446,N_6265);
xnor U6954 (N_6954,N_6199,N_6446);
nor U6955 (N_6955,N_6087,N_6160);
nand U6956 (N_6956,N_6279,N_6491);
nand U6957 (N_6957,N_6299,N_6068);
nand U6958 (N_6958,N_6354,N_6384);
xnor U6959 (N_6959,N_6260,N_6337);
nand U6960 (N_6960,N_6172,N_6352);
or U6961 (N_6961,N_6180,N_6258);
nand U6962 (N_6962,N_6342,N_6241);
nor U6963 (N_6963,N_6450,N_6120);
and U6964 (N_6964,N_6035,N_6033);
xor U6965 (N_6965,N_6107,N_6029);
nand U6966 (N_6966,N_6171,N_6184);
or U6967 (N_6967,N_6362,N_6140);
and U6968 (N_6968,N_6181,N_6103);
and U6969 (N_6969,N_6370,N_6310);
nand U6970 (N_6970,N_6269,N_6395);
nand U6971 (N_6971,N_6035,N_6486);
and U6972 (N_6972,N_6173,N_6396);
and U6973 (N_6973,N_6071,N_6374);
nor U6974 (N_6974,N_6234,N_6312);
or U6975 (N_6975,N_6410,N_6362);
xnor U6976 (N_6976,N_6042,N_6342);
and U6977 (N_6977,N_6035,N_6263);
nand U6978 (N_6978,N_6210,N_6491);
nand U6979 (N_6979,N_6114,N_6359);
nand U6980 (N_6980,N_6447,N_6204);
nor U6981 (N_6981,N_6333,N_6416);
nand U6982 (N_6982,N_6445,N_6311);
nand U6983 (N_6983,N_6434,N_6188);
nand U6984 (N_6984,N_6223,N_6131);
nor U6985 (N_6985,N_6091,N_6486);
nor U6986 (N_6986,N_6420,N_6133);
nor U6987 (N_6987,N_6380,N_6356);
nor U6988 (N_6988,N_6376,N_6208);
xnor U6989 (N_6989,N_6335,N_6184);
and U6990 (N_6990,N_6230,N_6095);
nand U6991 (N_6991,N_6218,N_6247);
and U6992 (N_6992,N_6261,N_6480);
nand U6993 (N_6993,N_6140,N_6029);
nand U6994 (N_6994,N_6292,N_6146);
and U6995 (N_6995,N_6161,N_6400);
nor U6996 (N_6996,N_6319,N_6197);
xor U6997 (N_6997,N_6143,N_6388);
and U6998 (N_6998,N_6015,N_6023);
and U6999 (N_6999,N_6435,N_6460);
or U7000 (N_7000,N_6902,N_6586);
nor U7001 (N_7001,N_6804,N_6650);
nor U7002 (N_7002,N_6634,N_6709);
or U7003 (N_7003,N_6674,N_6906);
and U7004 (N_7004,N_6899,N_6578);
or U7005 (N_7005,N_6675,N_6544);
and U7006 (N_7006,N_6811,N_6830);
xor U7007 (N_7007,N_6620,N_6720);
or U7008 (N_7008,N_6657,N_6583);
or U7009 (N_7009,N_6907,N_6738);
and U7010 (N_7010,N_6856,N_6809);
and U7011 (N_7011,N_6575,N_6501);
nor U7012 (N_7012,N_6557,N_6695);
xnor U7013 (N_7013,N_6786,N_6669);
nor U7014 (N_7014,N_6952,N_6623);
and U7015 (N_7015,N_6996,N_6938);
nand U7016 (N_7016,N_6834,N_6849);
nand U7017 (N_7017,N_6537,N_6805);
nor U7018 (N_7018,N_6829,N_6933);
xor U7019 (N_7019,N_6713,N_6677);
xor U7020 (N_7020,N_6788,N_6982);
nor U7021 (N_7021,N_6812,N_6820);
nor U7022 (N_7022,N_6892,N_6552);
xor U7023 (N_7023,N_6573,N_6912);
nand U7024 (N_7024,N_6900,N_6966);
nand U7025 (N_7025,N_6896,N_6965);
and U7026 (N_7026,N_6886,N_6676);
nor U7027 (N_7027,N_6706,N_6962);
xnor U7028 (N_7028,N_6800,N_6869);
and U7029 (N_7029,N_6777,N_6646);
and U7030 (N_7030,N_6762,N_6701);
or U7031 (N_7031,N_6511,N_6993);
nor U7032 (N_7032,N_6672,N_6600);
nor U7033 (N_7033,N_6603,N_6958);
nor U7034 (N_7034,N_6795,N_6678);
nand U7035 (N_7035,N_6908,N_6719);
or U7036 (N_7036,N_6942,N_6684);
xnor U7037 (N_7037,N_6960,N_6585);
or U7038 (N_7038,N_6589,N_6517);
xor U7039 (N_7039,N_6584,N_6877);
nor U7040 (N_7040,N_6564,N_6512);
xor U7041 (N_7041,N_6858,N_6518);
nand U7042 (N_7042,N_6970,N_6825);
nand U7043 (N_7043,N_6602,N_6734);
and U7044 (N_7044,N_6770,N_6617);
and U7045 (N_7045,N_6502,N_6992);
or U7046 (N_7046,N_6898,N_6928);
nand U7047 (N_7047,N_6598,N_6526);
and U7048 (N_7048,N_6859,N_6727);
or U7049 (N_7049,N_6643,N_6755);
nand U7050 (N_7050,N_6757,N_6500);
nand U7051 (N_7051,N_6865,N_6660);
nand U7052 (N_7052,N_6976,N_6988);
nand U7053 (N_7053,N_6813,N_6721);
nor U7054 (N_7054,N_6924,N_6563);
nand U7055 (N_7055,N_6789,N_6611);
or U7056 (N_7056,N_6717,N_6522);
and U7057 (N_7057,N_6513,N_6772);
or U7058 (N_7058,N_6778,N_6887);
and U7059 (N_7059,N_6978,N_6625);
nor U7060 (N_7060,N_6685,N_6696);
and U7061 (N_7061,N_6860,N_6974);
nor U7062 (N_7062,N_6521,N_6776);
nor U7063 (N_7063,N_6889,N_6519);
xnor U7064 (N_7064,N_6547,N_6707);
or U7065 (N_7065,N_6711,N_6852);
xnor U7066 (N_7066,N_6704,N_6740);
or U7067 (N_7067,N_6588,N_6750);
nand U7068 (N_7068,N_6806,N_6991);
or U7069 (N_7069,N_6922,N_6828);
xor U7070 (N_7070,N_6909,N_6903);
xnor U7071 (N_7071,N_6664,N_6923);
nor U7072 (N_7072,N_6523,N_6937);
xor U7073 (N_7073,N_6831,N_6539);
xor U7074 (N_7074,N_6702,N_6724);
nor U7075 (N_7075,N_6668,N_6606);
nor U7076 (N_7076,N_6735,N_6961);
xnor U7077 (N_7077,N_6601,N_6599);
nor U7078 (N_7078,N_6569,N_6870);
xnor U7079 (N_7079,N_6723,N_6648);
nor U7080 (N_7080,N_6614,N_6821);
nor U7081 (N_7081,N_6885,N_6577);
xor U7082 (N_7082,N_6979,N_6998);
or U7083 (N_7083,N_6572,N_6725);
and U7084 (N_7084,N_6510,N_6580);
or U7085 (N_7085,N_6835,N_6642);
nor U7086 (N_7086,N_6932,N_6627);
or U7087 (N_7087,N_6609,N_6618);
nand U7088 (N_7088,N_6596,N_6853);
and U7089 (N_7089,N_6981,N_6558);
xnor U7090 (N_7090,N_6631,N_6566);
or U7091 (N_7091,N_6836,N_6504);
and U7092 (N_7092,N_6972,N_6917);
and U7093 (N_7093,N_6803,N_6774);
and U7094 (N_7094,N_6639,N_6659);
or U7095 (N_7095,N_6655,N_6651);
nand U7096 (N_7096,N_6934,N_6638);
and U7097 (N_7097,N_6525,N_6781);
nand U7098 (N_7098,N_6833,N_6763);
xor U7099 (N_7099,N_6871,N_6946);
or U7100 (N_7100,N_6953,N_6703);
or U7101 (N_7101,N_6878,N_6729);
and U7102 (N_7102,N_6808,N_6760);
and U7103 (N_7103,N_6691,N_6653);
and U7104 (N_7104,N_6839,N_6536);
nand U7105 (N_7105,N_6964,N_6787);
xnor U7106 (N_7106,N_6766,N_6841);
nor U7107 (N_7107,N_6528,N_6890);
and U7108 (N_7108,N_6570,N_6694);
nand U7109 (N_7109,N_6911,N_6541);
or U7110 (N_7110,N_6957,N_6973);
xnor U7111 (N_7111,N_6799,N_6635);
or U7112 (N_7112,N_6556,N_6716);
or U7113 (N_7113,N_6861,N_6571);
nand U7114 (N_7114,N_6748,N_6505);
or U7115 (N_7115,N_6881,N_6925);
nand U7116 (N_7116,N_6615,N_6851);
or U7117 (N_7117,N_6689,N_6904);
or U7118 (N_7118,N_6619,N_6782);
or U7119 (N_7119,N_6594,N_6710);
and U7120 (N_7120,N_6817,N_6910);
and U7121 (N_7121,N_6567,N_6951);
xor U7122 (N_7122,N_6607,N_6545);
nor U7123 (N_7123,N_6759,N_6944);
or U7124 (N_7124,N_6665,N_6661);
nand U7125 (N_7125,N_6773,N_6508);
nor U7126 (N_7126,N_6714,N_6793);
xor U7127 (N_7127,N_6816,N_6534);
or U7128 (N_7128,N_6936,N_6656);
or U7129 (N_7129,N_6832,N_6593);
xnor U7130 (N_7130,N_6527,N_6948);
and U7131 (N_7131,N_6801,N_6652);
and U7132 (N_7132,N_6524,N_6949);
nand U7133 (N_7133,N_6555,N_6985);
or U7134 (N_7134,N_6548,N_6968);
nor U7135 (N_7135,N_6531,N_6514);
nand U7136 (N_7136,N_6784,N_6785);
nand U7137 (N_7137,N_6969,N_6746);
nand U7138 (N_7138,N_6700,N_6814);
nor U7139 (N_7139,N_6956,N_6579);
and U7140 (N_7140,N_6509,N_6921);
nor U7141 (N_7141,N_6848,N_6561);
or U7142 (N_7142,N_6764,N_6679);
nor U7143 (N_7143,N_6919,N_6940);
nor U7144 (N_7144,N_6636,N_6975);
xnor U7145 (N_7145,N_6977,N_6914);
nor U7146 (N_7146,N_6765,N_6913);
xor U7147 (N_7147,N_6775,N_6824);
or U7148 (N_7148,N_6538,N_6810);
and U7149 (N_7149,N_6733,N_6743);
nand U7150 (N_7150,N_6927,N_6994);
xnor U7151 (N_7151,N_6761,N_6855);
nor U7152 (N_7152,N_6945,N_6649);
nand U7153 (N_7153,N_6752,N_6779);
nand U7154 (N_7154,N_6520,N_6613);
and U7155 (N_7155,N_6891,N_6726);
nand U7156 (N_7156,N_6741,N_6790);
and U7157 (N_7157,N_6591,N_6622);
nand U7158 (N_7158,N_6749,N_6582);
nand U7159 (N_7159,N_6901,N_6780);
nand U7160 (N_7160,N_6843,N_6670);
nand U7161 (N_7161,N_6529,N_6967);
xor U7162 (N_7162,N_6535,N_6797);
xor U7163 (N_7163,N_6872,N_6687);
and U7164 (N_7164,N_6632,N_6983);
nand U7165 (N_7165,N_6783,N_6666);
nor U7166 (N_7166,N_6918,N_6895);
or U7167 (N_7167,N_6604,N_6697);
xnor U7168 (N_7168,N_6915,N_6984);
nand U7169 (N_7169,N_6673,N_6882);
xor U7170 (N_7170,N_6875,N_6963);
nand U7171 (N_7171,N_6827,N_6647);
nor U7172 (N_7172,N_6612,N_6692);
nand U7173 (N_7173,N_6863,N_6715);
nand U7174 (N_7174,N_6605,N_6667);
and U7175 (N_7175,N_6862,N_6722);
nor U7176 (N_7176,N_6626,N_6837);
nor U7177 (N_7177,N_6767,N_6971);
nor U7178 (N_7178,N_6542,N_6530);
or U7179 (N_7179,N_6515,N_6641);
nand U7180 (N_7180,N_6616,N_6690);
or U7181 (N_7181,N_6873,N_6897);
nand U7182 (N_7182,N_6798,N_6840);
xnor U7183 (N_7183,N_6663,N_6728);
or U7184 (N_7184,N_6645,N_6562);
xor U7185 (N_7185,N_6796,N_6818);
xnor U7186 (N_7186,N_6565,N_6553);
nand U7187 (N_7187,N_6794,N_6929);
and U7188 (N_7188,N_6621,N_6559);
xnor U7189 (N_7189,N_6950,N_6920);
or U7190 (N_7190,N_6980,N_6543);
or U7191 (N_7191,N_6756,N_6595);
nor U7192 (N_7192,N_6597,N_6712);
and U7193 (N_7193,N_6718,N_6662);
nor U7194 (N_7194,N_6546,N_6705);
xor U7195 (N_7195,N_6751,N_6864);
nor U7196 (N_7196,N_6905,N_6815);
nor U7197 (N_7197,N_6995,N_6850);
and U7198 (N_7198,N_6532,N_6930);
and U7199 (N_7199,N_6628,N_6989);
nor U7200 (N_7200,N_6742,N_6879);
and U7201 (N_7201,N_6516,N_6866);
nor U7202 (N_7202,N_6999,N_6681);
or U7203 (N_7203,N_6874,N_6540);
or U7204 (N_7204,N_6854,N_6732);
nor U7205 (N_7205,N_6654,N_6758);
nand U7206 (N_7206,N_6629,N_6574);
nand U7207 (N_7207,N_6916,N_6633);
xor U7208 (N_7208,N_6826,N_6838);
and U7209 (N_7209,N_6847,N_6637);
and U7210 (N_7210,N_6744,N_6592);
or U7211 (N_7211,N_6739,N_6926);
and U7212 (N_7212,N_6644,N_6737);
and U7213 (N_7213,N_6802,N_6560);
nor U7214 (N_7214,N_6686,N_6943);
xor U7215 (N_7215,N_6883,N_6658);
nor U7216 (N_7216,N_6939,N_6941);
xnor U7217 (N_7217,N_6807,N_6819);
xnor U7218 (N_7218,N_6893,N_6507);
nand U7219 (N_7219,N_6754,N_6791);
nor U7220 (N_7220,N_6624,N_6792);
xnor U7221 (N_7221,N_6503,N_6888);
or U7222 (N_7222,N_6954,N_6506);
xor U7223 (N_7223,N_6680,N_6959);
nor U7224 (N_7224,N_6745,N_6688);
and U7225 (N_7225,N_6708,N_6880);
or U7226 (N_7226,N_6844,N_6576);
nor U7227 (N_7227,N_6568,N_6867);
and U7228 (N_7228,N_6587,N_6987);
xnor U7229 (N_7229,N_6581,N_6730);
xnor U7230 (N_7230,N_6894,N_6551);
nor U7231 (N_7231,N_6533,N_6671);
and U7232 (N_7232,N_6549,N_6822);
nor U7233 (N_7233,N_6736,N_6845);
xor U7234 (N_7234,N_6990,N_6590);
and U7235 (N_7235,N_6997,N_6693);
nand U7236 (N_7236,N_6935,N_6699);
xor U7237 (N_7237,N_6876,N_6683);
or U7238 (N_7238,N_6771,N_6550);
nor U7239 (N_7239,N_6931,N_6731);
and U7240 (N_7240,N_6640,N_6630);
xnor U7241 (N_7241,N_6842,N_6768);
or U7242 (N_7242,N_6823,N_6610);
and U7243 (N_7243,N_6884,N_6747);
and U7244 (N_7244,N_6955,N_6608);
and U7245 (N_7245,N_6868,N_6986);
and U7246 (N_7246,N_6682,N_6769);
or U7247 (N_7247,N_6698,N_6947);
and U7248 (N_7248,N_6857,N_6846);
and U7249 (N_7249,N_6753,N_6554);
xor U7250 (N_7250,N_6690,N_6853);
nor U7251 (N_7251,N_6541,N_6920);
or U7252 (N_7252,N_6571,N_6693);
nand U7253 (N_7253,N_6962,N_6894);
or U7254 (N_7254,N_6738,N_6742);
nor U7255 (N_7255,N_6855,N_6507);
nor U7256 (N_7256,N_6886,N_6724);
or U7257 (N_7257,N_6950,N_6687);
nor U7258 (N_7258,N_6974,N_6511);
nor U7259 (N_7259,N_6922,N_6717);
and U7260 (N_7260,N_6635,N_6786);
nor U7261 (N_7261,N_6758,N_6593);
and U7262 (N_7262,N_6737,N_6761);
nor U7263 (N_7263,N_6598,N_6906);
and U7264 (N_7264,N_6767,N_6889);
nor U7265 (N_7265,N_6790,N_6533);
xor U7266 (N_7266,N_6647,N_6793);
nand U7267 (N_7267,N_6988,N_6882);
or U7268 (N_7268,N_6684,N_6786);
or U7269 (N_7269,N_6814,N_6710);
xor U7270 (N_7270,N_6543,N_6875);
xnor U7271 (N_7271,N_6509,N_6731);
nor U7272 (N_7272,N_6768,N_6935);
nor U7273 (N_7273,N_6970,N_6648);
nand U7274 (N_7274,N_6843,N_6883);
and U7275 (N_7275,N_6765,N_6500);
and U7276 (N_7276,N_6664,N_6864);
nand U7277 (N_7277,N_6856,N_6889);
xor U7278 (N_7278,N_6947,N_6628);
nand U7279 (N_7279,N_6627,N_6935);
nand U7280 (N_7280,N_6892,N_6577);
and U7281 (N_7281,N_6904,N_6618);
xor U7282 (N_7282,N_6824,N_6791);
nor U7283 (N_7283,N_6950,N_6570);
nor U7284 (N_7284,N_6822,N_6815);
xnor U7285 (N_7285,N_6836,N_6521);
or U7286 (N_7286,N_6686,N_6992);
and U7287 (N_7287,N_6501,N_6981);
nand U7288 (N_7288,N_6565,N_6857);
and U7289 (N_7289,N_6689,N_6659);
nor U7290 (N_7290,N_6856,N_6556);
or U7291 (N_7291,N_6586,N_6623);
nand U7292 (N_7292,N_6733,N_6581);
nand U7293 (N_7293,N_6516,N_6978);
nor U7294 (N_7294,N_6926,N_6931);
xor U7295 (N_7295,N_6550,N_6670);
xor U7296 (N_7296,N_6770,N_6828);
or U7297 (N_7297,N_6811,N_6504);
and U7298 (N_7298,N_6633,N_6676);
nor U7299 (N_7299,N_6971,N_6511);
nand U7300 (N_7300,N_6583,N_6823);
xnor U7301 (N_7301,N_6891,N_6950);
or U7302 (N_7302,N_6646,N_6820);
nand U7303 (N_7303,N_6880,N_6926);
xnor U7304 (N_7304,N_6665,N_6657);
nand U7305 (N_7305,N_6611,N_6541);
nor U7306 (N_7306,N_6813,N_6599);
nand U7307 (N_7307,N_6902,N_6989);
or U7308 (N_7308,N_6885,N_6741);
nor U7309 (N_7309,N_6626,N_6631);
xnor U7310 (N_7310,N_6643,N_6895);
nor U7311 (N_7311,N_6752,N_6789);
nand U7312 (N_7312,N_6687,N_6990);
xor U7313 (N_7313,N_6982,N_6535);
nor U7314 (N_7314,N_6939,N_6713);
nand U7315 (N_7315,N_6747,N_6577);
xor U7316 (N_7316,N_6736,N_6722);
nand U7317 (N_7317,N_6675,N_6800);
or U7318 (N_7318,N_6810,N_6971);
nand U7319 (N_7319,N_6696,N_6512);
or U7320 (N_7320,N_6751,N_6722);
and U7321 (N_7321,N_6979,N_6917);
nand U7322 (N_7322,N_6802,N_6960);
nand U7323 (N_7323,N_6602,N_6913);
nor U7324 (N_7324,N_6830,N_6667);
nor U7325 (N_7325,N_6500,N_6691);
or U7326 (N_7326,N_6535,N_6849);
or U7327 (N_7327,N_6555,N_6894);
nor U7328 (N_7328,N_6524,N_6832);
nand U7329 (N_7329,N_6752,N_6807);
and U7330 (N_7330,N_6773,N_6655);
nand U7331 (N_7331,N_6920,N_6914);
nand U7332 (N_7332,N_6650,N_6793);
xnor U7333 (N_7333,N_6552,N_6614);
xnor U7334 (N_7334,N_6522,N_6819);
or U7335 (N_7335,N_6548,N_6972);
xnor U7336 (N_7336,N_6502,N_6785);
xor U7337 (N_7337,N_6576,N_6602);
or U7338 (N_7338,N_6894,N_6632);
or U7339 (N_7339,N_6832,N_6861);
nor U7340 (N_7340,N_6793,N_6732);
xor U7341 (N_7341,N_6639,N_6954);
or U7342 (N_7342,N_6927,N_6829);
nand U7343 (N_7343,N_6964,N_6916);
nor U7344 (N_7344,N_6763,N_6734);
nand U7345 (N_7345,N_6584,N_6897);
nor U7346 (N_7346,N_6576,N_6951);
nor U7347 (N_7347,N_6657,N_6774);
and U7348 (N_7348,N_6535,N_6859);
xor U7349 (N_7349,N_6811,N_6539);
nand U7350 (N_7350,N_6612,N_6870);
xnor U7351 (N_7351,N_6877,N_6742);
or U7352 (N_7352,N_6943,N_6980);
xnor U7353 (N_7353,N_6574,N_6929);
nor U7354 (N_7354,N_6986,N_6663);
nand U7355 (N_7355,N_6762,N_6995);
and U7356 (N_7356,N_6752,N_6915);
nand U7357 (N_7357,N_6835,N_6543);
and U7358 (N_7358,N_6625,N_6899);
and U7359 (N_7359,N_6758,N_6591);
nor U7360 (N_7360,N_6734,N_6977);
nand U7361 (N_7361,N_6852,N_6786);
xor U7362 (N_7362,N_6551,N_6568);
nand U7363 (N_7363,N_6566,N_6685);
nand U7364 (N_7364,N_6501,N_6730);
or U7365 (N_7365,N_6659,N_6622);
or U7366 (N_7366,N_6839,N_6521);
xor U7367 (N_7367,N_6927,N_6843);
xor U7368 (N_7368,N_6947,N_6864);
nand U7369 (N_7369,N_6769,N_6714);
and U7370 (N_7370,N_6563,N_6897);
and U7371 (N_7371,N_6815,N_6875);
and U7372 (N_7372,N_6933,N_6793);
and U7373 (N_7373,N_6758,N_6753);
nor U7374 (N_7374,N_6901,N_6726);
nor U7375 (N_7375,N_6884,N_6989);
and U7376 (N_7376,N_6833,N_6713);
xor U7377 (N_7377,N_6705,N_6579);
and U7378 (N_7378,N_6621,N_6757);
and U7379 (N_7379,N_6999,N_6694);
or U7380 (N_7380,N_6968,N_6674);
nand U7381 (N_7381,N_6771,N_6807);
xnor U7382 (N_7382,N_6550,N_6838);
nand U7383 (N_7383,N_6812,N_6985);
nor U7384 (N_7384,N_6840,N_6780);
and U7385 (N_7385,N_6977,N_6566);
and U7386 (N_7386,N_6766,N_6562);
nor U7387 (N_7387,N_6934,N_6747);
nor U7388 (N_7388,N_6616,N_6845);
or U7389 (N_7389,N_6551,N_6745);
xor U7390 (N_7390,N_6557,N_6906);
nor U7391 (N_7391,N_6651,N_6908);
xnor U7392 (N_7392,N_6966,N_6889);
nor U7393 (N_7393,N_6509,N_6551);
nor U7394 (N_7394,N_6933,N_6778);
nor U7395 (N_7395,N_6652,N_6708);
or U7396 (N_7396,N_6608,N_6778);
or U7397 (N_7397,N_6923,N_6525);
and U7398 (N_7398,N_6832,N_6858);
nand U7399 (N_7399,N_6611,N_6931);
and U7400 (N_7400,N_6939,N_6639);
nand U7401 (N_7401,N_6740,N_6803);
and U7402 (N_7402,N_6885,N_6679);
nand U7403 (N_7403,N_6913,N_6641);
xnor U7404 (N_7404,N_6589,N_6857);
or U7405 (N_7405,N_6959,N_6575);
nand U7406 (N_7406,N_6783,N_6615);
xor U7407 (N_7407,N_6971,N_6616);
and U7408 (N_7408,N_6513,N_6917);
and U7409 (N_7409,N_6990,N_6506);
nand U7410 (N_7410,N_6669,N_6749);
and U7411 (N_7411,N_6722,N_6901);
or U7412 (N_7412,N_6584,N_6662);
nor U7413 (N_7413,N_6502,N_6868);
xnor U7414 (N_7414,N_6639,N_6904);
nand U7415 (N_7415,N_6895,N_6530);
or U7416 (N_7416,N_6949,N_6708);
nor U7417 (N_7417,N_6833,N_6657);
or U7418 (N_7418,N_6930,N_6997);
and U7419 (N_7419,N_6982,N_6950);
or U7420 (N_7420,N_6716,N_6758);
xor U7421 (N_7421,N_6538,N_6694);
nand U7422 (N_7422,N_6889,N_6814);
xor U7423 (N_7423,N_6875,N_6563);
nand U7424 (N_7424,N_6734,N_6928);
nor U7425 (N_7425,N_6650,N_6660);
nor U7426 (N_7426,N_6881,N_6559);
nor U7427 (N_7427,N_6517,N_6800);
nand U7428 (N_7428,N_6892,N_6541);
xnor U7429 (N_7429,N_6910,N_6516);
nor U7430 (N_7430,N_6691,N_6574);
or U7431 (N_7431,N_6723,N_6669);
nand U7432 (N_7432,N_6502,N_6512);
and U7433 (N_7433,N_6951,N_6885);
xor U7434 (N_7434,N_6971,N_6823);
nor U7435 (N_7435,N_6915,N_6694);
nand U7436 (N_7436,N_6701,N_6932);
nor U7437 (N_7437,N_6909,N_6874);
xor U7438 (N_7438,N_6973,N_6868);
or U7439 (N_7439,N_6565,N_6908);
nand U7440 (N_7440,N_6661,N_6595);
or U7441 (N_7441,N_6688,N_6935);
and U7442 (N_7442,N_6574,N_6536);
nand U7443 (N_7443,N_6906,N_6646);
nor U7444 (N_7444,N_6918,N_6796);
nor U7445 (N_7445,N_6501,N_6615);
or U7446 (N_7446,N_6571,N_6836);
nor U7447 (N_7447,N_6526,N_6511);
or U7448 (N_7448,N_6857,N_6800);
xnor U7449 (N_7449,N_6889,N_6655);
nand U7450 (N_7450,N_6553,N_6566);
and U7451 (N_7451,N_6813,N_6676);
and U7452 (N_7452,N_6956,N_6939);
and U7453 (N_7453,N_6587,N_6554);
or U7454 (N_7454,N_6856,N_6796);
nand U7455 (N_7455,N_6591,N_6693);
and U7456 (N_7456,N_6729,N_6821);
or U7457 (N_7457,N_6611,N_6686);
xnor U7458 (N_7458,N_6853,N_6777);
and U7459 (N_7459,N_6626,N_6597);
xnor U7460 (N_7460,N_6943,N_6652);
nor U7461 (N_7461,N_6934,N_6795);
nand U7462 (N_7462,N_6980,N_6632);
nor U7463 (N_7463,N_6642,N_6659);
or U7464 (N_7464,N_6628,N_6575);
and U7465 (N_7465,N_6665,N_6762);
and U7466 (N_7466,N_6805,N_6754);
or U7467 (N_7467,N_6853,N_6869);
nor U7468 (N_7468,N_6798,N_6637);
and U7469 (N_7469,N_6646,N_6910);
nand U7470 (N_7470,N_6614,N_6694);
or U7471 (N_7471,N_6511,N_6643);
nor U7472 (N_7472,N_6903,N_6825);
nand U7473 (N_7473,N_6570,N_6835);
and U7474 (N_7474,N_6952,N_6773);
nor U7475 (N_7475,N_6616,N_6974);
nor U7476 (N_7476,N_6615,N_6766);
nor U7477 (N_7477,N_6975,N_6991);
and U7478 (N_7478,N_6961,N_6746);
nand U7479 (N_7479,N_6862,N_6819);
nor U7480 (N_7480,N_6751,N_6677);
nand U7481 (N_7481,N_6927,N_6686);
or U7482 (N_7482,N_6500,N_6956);
and U7483 (N_7483,N_6847,N_6870);
xnor U7484 (N_7484,N_6953,N_6716);
nor U7485 (N_7485,N_6991,N_6965);
or U7486 (N_7486,N_6985,N_6683);
nand U7487 (N_7487,N_6827,N_6945);
nand U7488 (N_7488,N_6837,N_6976);
nor U7489 (N_7489,N_6822,N_6925);
and U7490 (N_7490,N_6968,N_6854);
xor U7491 (N_7491,N_6940,N_6861);
nor U7492 (N_7492,N_6656,N_6800);
nor U7493 (N_7493,N_6906,N_6914);
and U7494 (N_7494,N_6910,N_6638);
and U7495 (N_7495,N_6953,N_6675);
or U7496 (N_7496,N_6799,N_6985);
nand U7497 (N_7497,N_6673,N_6618);
xor U7498 (N_7498,N_6938,N_6914);
or U7499 (N_7499,N_6660,N_6951);
nand U7500 (N_7500,N_7206,N_7469);
nand U7501 (N_7501,N_7311,N_7151);
or U7502 (N_7502,N_7461,N_7121);
nor U7503 (N_7503,N_7064,N_7336);
and U7504 (N_7504,N_7439,N_7371);
or U7505 (N_7505,N_7181,N_7490);
xor U7506 (N_7506,N_7250,N_7315);
nor U7507 (N_7507,N_7210,N_7015);
nand U7508 (N_7508,N_7377,N_7073);
or U7509 (N_7509,N_7182,N_7270);
nand U7510 (N_7510,N_7170,N_7186);
and U7511 (N_7511,N_7496,N_7264);
or U7512 (N_7512,N_7423,N_7018);
xor U7513 (N_7513,N_7128,N_7484);
nand U7514 (N_7514,N_7465,N_7014);
and U7515 (N_7515,N_7157,N_7414);
nand U7516 (N_7516,N_7456,N_7455);
xnor U7517 (N_7517,N_7180,N_7040);
nor U7518 (N_7518,N_7175,N_7196);
nor U7519 (N_7519,N_7050,N_7364);
xnor U7520 (N_7520,N_7269,N_7255);
xor U7521 (N_7521,N_7246,N_7229);
nand U7522 (N_7522,N_7072,N_7495);
nor U7523 (N_7523,N_7214,N_7091);
nand U7524 (N_7524,N_7174,N_7438);
nor U7525 (N_7525,N_7298,N_7322);
xnor U7526 (N_7526,N_7143,N_7079);
nand U7527 (N_7527,N_7382,N_7267);
nand U7528 (N_7528,N_7065,N_7286);
nand U7529 (N_7529,N_7357,N_7388);
nor U7530 (N_7530,N_7002,N_7419);
and U7531 (N_7531,N_7462,N_7070);
nand U7532 (N_7532,N_7329,N_7037);
and U7533 (N_7533,N_7265,N_7193);
xor U7534 (N_7534,N_7172,N_7370);
and U7535 (N_7535,N_7467,N_7476);
nand U7536 (N_7536,N_7062,N_7154);
xor U7537 (N_7537,N_7296,N_7260);
nor U7538 (N_7538,N_7138,N_7191);
xor U7539 (N_7539,N_7036,N_7375);
and U7540 (N_7540,N_7346,N_7249);
nor U7541 (N_7541,N_7284,N_7078);
xor U7542 (N_7542,N_7099,N_7188);
nor U7543 (N_7543,N_7258,N_7007);
xor U7544 (N_7544,N_7137,N_7245);
xnor U7545 (N_7545,N_7444,N_7297);
nand U7546 (N_7546,N_7351,N_7426);
or U7547 (N_7547,N_7092,N_7033);
nand U7548 (N_7548,N_7126,N_7123);
xor U7549 (N_7549,N_7204,N_7344);
and U7550 (N_7550,N_7392,N_7135);
nor U7551 (N_7551,N_7294,N_7082);
nand U7552 (N_7552,N_7118,N_7119);
and U7553 (N_7553,N_7316,N_7431);
nor U7554 (N_7554,N_7140,N_7363);
nor U7555 (N_7555,N_7242,N_7220);
or U7556 (N_7556,N_7049,N_7303);
nor U7557 (N_7557,N_7306,N_7468);
nor U7558 (N_7558,N_7323,N_7302);
and U7559 (N_7559,N_7086,N_7202);
and U7560 (N_7560,N_7068,N_7480);
or U7561 (N_7561,N_7057,N_7141);
and U7562 (N_7562,N_7254,N_7142);
nand U7563 (N_7563,N_7256,N_7261);
nand U7564 (N_7564,N_7027,N_7477);
nand U7565 (N_7565,N_7457,N_7360);
or U7566 (N_7566,N_7034,N_7418);
xnor U7567 (N_7567,N_7453,N_7084);
or U7568 (N_7568,N_7130,N_7083);
nor U7569 (N_7569,N_7032,N_7074);
nand U7570 (N_7570,N_7482,N_7061);
and U7571 (N_7571,N_7281,N_7402);
and U7572 (N_7572,N_7237,N_7103);
xor U7573 (N_7573,N_7272,N_7069);
or U7574 (N_7574,N_7285,N_7197);
or U7575 (N_7575,N_7077,N_7224);
or U7576 (N_7576,N_7328,N_7485);
nor U7577 (N_7577,N_7136,N_7163);
xor U7578 (N_7578,N_7190,N_7021);
or U7579 (N_7579,N_7177,N_7327);
nand U7580 (N_7580,N_7241,N_7248);
and U7581 (N_7581,N_7435,N_7359);
nand U7582 (N_7582,N_7029,N_7275);
or U7583 (N_7583,N_7318,N_7499);
and U7584 (N_7584,N_7454,N_7397);
nor U7585 (N_7585,N_7319,N_7189);
nor U7586 (N_7586,N_7301,N_7276);
nor U7587 (N_7587,N_7263,N_7024);
and U7588 (N_7588,N_7449,N_7113);
and U7589 (N_7589,N_7430,N_7347);
nor U7590 (N_7590,N_7404,N_7139);
or U7591 (N_7591,N_7479,N_7169);
or U7592 (N_7592,N_7432,N_7396);
nor U7593 (N_7593,N_7150,N_7109);
xnor U7594 (N_7594,N_7314,N_7259);
nor U7595 (N_7595,N_7108,N_7152);
nand U7596 (N_7596,N_7277,N_7350);
nand U7597 (N_7597,N_7039,N_7192);
and U7598 (N_7598,N_7195,N_7147);
nor U7599 (N_7599,N_7106,N_7464);
and U7600 (N_7600,N_7085,N_7112);
nand U7601 (N_7601,N_7216,N_7001);
or U7602 (N_7602,N_7425,N_7101);
xnor U7603 (N_7603,N_7310,N_7349);
xnor U7604 (N_7604,N_7299,N_7230);
or U7605 (N_7605,N_7361,N_7421);
nor U7606 (N_7606,N_7409,N_7131);
and U7607 (N_7607,N_7110,N_7107);
or U7608 (N_7608,N_7279,N_7096);
and U7609 (N_7609,N_7274,N_7307);
nand U7610 (N_7610,N_7129,N_7338);
xnor U7611 (N_7611,N_7355,N_7017);
nor U7612 (N_7612,N_7104,N_7341);
or U7613 (N_7613,N_7288,N_7162);
nor U7614 (N_7614,N_7395,N_7489);
nand U7615 (N_7615,N_7117,N_7333);
nand U7616 (N_7616,N_7293,N_7471);
nor U7617 (N_7617,N_7217,N_7058);
nand U7618 (N_7618,N_7443,N_7025);
nand U7619 (N_7619,N_7401,N_7013);
nand U7620 (N_7620,N_7168,N_7045);
nand U7621 (N_7621,N_7184,N_7451);
xnor U7622 (N_7622,N_7075,N_7097);
and U7623 (N_7623,N_7330,N_7226);
xor U7624 (N_7624,N_7011,N_7428);
or U7625 (N_7625,N_7046,N_7478);
xnor U7626 (N_7626,N_7098,N_7022);
or U7627 (N_7627,N_7199,N_7209);
or U7628 (N_7628,N_7362,N_7212);
and U7629 (N_7629,N_7283,N_7223);
nand U7630 (N_7630,N_7243,N_7134);
nand U7631 (N_7631,N_7146,N_7483);
xnor U7632 (N_7632,N_7056,N_7102);
nor U7633 (N_7633,N_7047,N_7312);
nand U7634 (N_7634,N_7387,N_7198);
and U7635 (N_7635,N_7358,N_7090);
xnor U7636 (N_7636,N_7400,N_7171);
or U7637 (N_7637,N_7187,N_7252);
nand U7638 (N_7638,N_7342,N_7234);
xor U7639 (N_7639,N_7394,N_7266);
xor U7640 (N_7640,N_7340,N_7020);
xnor U7641 (N_7641,N_7326,N_7491);
nand U7642 (N_7642,N_7348,N_7185);
nor U7643 (N_7643,N_7335,N_7459);
xor U7644 (N_7644,N_7390,N_7399);
xnor U7645 (N_7645,N_7164,N_7225);
xnor U7646 (N_7646,N_7417,N_7228);
nor U7647 (N_7647,N_7309,N_7376);
or U7648 (N_7648,N_7200,N_7010);
and U7649 (N_7649,N_7238,N_7379);
nor U7650 (N_7650,N_7089,N_7067);
xor U7651 (N_7651,N_7374,N_7161);
xnor U7652 (N_7652,N_7433,N_7145);
xnor U7653 (N_7653,N_7044,N_7203);
and U7654 (N_7654,N_7367,N_7095);
or U7655 (N_7655,N_7240,N_7247);
or U7656 (N_7656,N_7133,N_7236);
nand U7657 (N_7657,N_7369,N_7378);
xor U7658 (N_7658,N_7304,N_7295);
nor U7659 (N_7659,N_7475,N_7381);
nand U7660 (N_7660,N_7231,N_7012);
and U7661 (N_7661,N_7041,N_7268);
xnor U7662 (N_7662,N_7125,N_7087);
and U7663 (N_7663,N_7373,N_7043);
or U7664 (N_7664,N_7410,N_7415);
nand U7665 (N_7665,N_7324,N_7321);
or U7666 (N_7666,N_7159,N_7132);
and U7667 (N_7667,N_7149,N_7386);
and U7668 (N_7668,N_7116,N_7111);
nand U7669 (N_7669,N_7028,N_7160);
and U7670 (N_7670,N_7215,N_7127);
xor U7671 (N_7671,N_7420,N_7273);
or U7672 (N_7672,N_7218,N_7179);
nor U7673 (N_7673,N_7300,N_7019);
and U7674 (N_7674,N_7416,N_7144);
nor U7675 (N_7675,N_7004,N_7412);
and U7676 (N_7676,N_7262,N_7257);
or U7677 (N_7677,N_7317,N_7366);
and U7678 (N_7678,N_7406,N_7278);
or U7679 (N_7679,N_7447,N_7060);
nand U7680 (N_7680,N_7308,N_7365);
nand U7681 (N_7681,N_7398,N_7063);
or U7682 (N_7682,N_7282,N_7173);
or U7683 (N_7683,N_7081,N_7290);
and U7684 (N_7684,N_7385,N_7023);
and U7685 (N_7685,N_7411,N_7292);
and U7686 (N_7686,N_7492,N_7009);
nand U7687 (N_7687,N_7219,N_7059);
xor U7688 (N_7688,N_7393,N_7088);
nor U7689 (N_7689,N_7052,N_7035);
xor U7690 (N_7690,N_7337,N_7227);
nand U7691 (N_7691,N_7353,N_7251);
nor U7692 (N_7692,N_7194,N_7165);
nand U7693 (N_7693,N_7498,N_7093);
and U7694 (N_7694,N_7458,N_7466);
or U7695 (N_7695,N_7071,N_7222);
xor U7696 (N_7696,N_7384,N_7178);
xor U7697 (N_7697,N_7332,N_7114);
xnor U7698 (N_7698,N_7003,N_7481);
or U7699 (N_7699,N_7183,N_7094);
nor U7700 (N_7700,N_7497,N_7053);
nand U7701 (N_7701,N_7124,N_7354);
xor U7702 (N_7702,N_7372,N_7460);
or U7703 (N_7703,N_7474,N_7148);
nor U7704 (N_7704,N_7389,N_7166);
xor U7705 (N_7705,N_7427,N_7448);
nor U7706 (N_7706,N_7213,N_7105);
or U7707 (N_7707,N_7352,N_7100);
and U7708 (N_7708,N_7280,N_7331);
and U7709 (N_7709,N_7176,N_7445);
or U7710 (N_7710,N_7424,N_7383);
nand U7711 (N_7711,N_7452,N_7343);
xor U7712 (N_7712,N_7436,N_7473);
nor U7713 (N_7713,N_7155,N_7030);
nor U7714 (N_7714,N_7076,N_7472);
or U7715 (N_7715,N_7038,N_7334);
and U7716 (N_7716,N_7488,N_7016);
xnor U7717 (N_7717,N_7407,N_7391);
nand U7718 (N_7718,N_7313,N_7494);
nor U7719 (N_7719,N_7291,N_7211);
xor U7720 (N_7720,N_7325,N_7031);
or U7721 (N_7721,N_7320,N_7287);
xnor U7722 (N_7722,N_7120,N_7115);
and U7723 (N_7723,N_7403,N_7463);
nor U7724 (N_7724,N_7006,N_7493);
xnor U7725 (N_7725,N_7167,N_7413);
or U7726 (N_7726,N_7380,N_7158);
xnor U7727 (N_7727,N_7446,N_7305);
or U7728 (N_7728,N_7000,N_7405);
nand U7729 (N_7729,N_7048,N_7066);
nand U7730 (N_7730,N_7450,N_7440);
or U7731 (N_7731,N_7055,N_7487);
nand U7732 (N_7732,N_7345,N_7339);
xor U7733 (N_7733,N_7051,N_7235);
and U7734 (N_7734,N_7026,N_7122);
nand U7735 (N_7735,N_7244,N_7233);
and U7736 (N_7736,N_7208,N_7080);
nand U7737 (N_7737,N_7042,N_7205);
or U7738 (N_7738,N_7005,N_7008);
or U7739 (N_7739,N_7271,N_7221);
xnor U7740 (N_7740,N_7207,N_7442);
nor U7741 (N_7741,N_7408,N_7253);
nor U7742 (N_7742,N_7437,N_7441);
or U7743 (N_7743,N_7422,N_7232);
and U7744 (N_7744,N_7289,N_7156);
or U7745 (N_7745,N_7054,N_7434);
and U7746 (N_7746,N_7429,N_7153);
or U7747 (N_7747,N_7470,N_7368);
and U7748 (N_7748,N_7239,N_7201);
and U7749 (N_7749,N_7486,N_7356);
nor U7750 (N_7750,N_7008,N_7486);
and U7751 (N_7751,N_7225,N_7318);
and U7752 (N_7752,N_7221,N_7283);
xor U7753 (N_7753,N_7296,N_7417);
nand U7754 (N_7754,N_7033,N_7080);
or U7755 (N_7755,N_7447,N_7458);
nor U7756 (N_7756,N_7161,N_7326);
nor U7757 (N_7757,N_7404,N_7381);
and U7758 (N_7758,N_7242,N_7115);
and U7759 (N_7759,N_7165,N_7275);
or U7760 (N_7760,N_7437,N_7040);
nand U7761 (N_7761,N_7135,N_7314);
nand U7762 (N_7762,N_7481,N_7387);
nor U7763 (N_7763,N_7403,N_7416);
and U7764 (N_7764,N_7185,N_7124);
nand U7765 (N_7765,N_7168,N_7377);
nand U7766 (N_7766,N_7401,N_7156);
xnor U7767 (N_7767,N_7390,N_7311);
and U7768 (N_7768,N_7079,N_7477);
xor U7769 (N_7769,N_7212,N_7213);
nor U7770 (N_7770,N_7003,N_7256);
or U7771 (N_7771,N_7418,N_7226);
and U7772 (N_7772,N_7167,N_7221);
xor U7773 (N_7773,N_7218,N_7158);
and U7774 (N_7774,N_7344,N_7252);
nand U7775 (N_7775,N_7453,N_7197);
xnor U7776 (N_7776,N_7193,N_7121);
nand U7777 (N_7777,N_7495,N_7472);
xor U7778 (N_7778,N_7272,N_7153);
nand U7779 (N_7779,N_7106,N_7063);
and U7780 (N_7780,N_7476,N_7038);
and U7781 (N_7781,N_7134,N_7415);
and U7782 (N_7782,N_7403,N_7281);
xnor U7783 (N_7783,N_7308,N_7179);
nand U7784 (N_7784,N_7465,N_7017);
and U7785 (N_7785,N_7047,N_7415);
xnor U7786 (N_7786,N_7254,N_7198);
and U7787 (N_7787,N_7131,N_7473);
xnor U7788 (N_7788,N_7010,N_7313);
xor U7789 (N_7789,N_7082,N_7278);
nand U7790 (N_7790,N_7236,N_7270);
and U7791 (N_7791,N_7289,N_7316);
and U7792 (N_7792,N_7227,N_7242);
and U7793 (N_7793,N_7095,N_7008);
nor U7794 (N_7794,N_7108,N_7424);
nand U7795 (N_7795,N_7301,N_7416);
xor U7796 (N_7796,N_7049,N_7179);
nand U7797 (N_7797,N_7010,N_7304);
nand U7798 (N_7798,N_7113,N_7439);
nor U7799 (N_7799,N_7182,N_7324);
nand U7800 (N_7800,N_7369,N_7411);
and U7801 (N_7801,N_7442,N_7349);
xor U7802 (N_7802,N_7419,N_7400);
nand U7803 (N_7803,N_7356,N_7399);
nor U7804 (N_7804,N_7177,N_7385);
nor U7805 (N_7805,N_7038,N_7403);
and U7806 (N_7806,N_7095,N_7472);
or U7807 (N_7807,N_7352,N_7153);
and U7808 (N_7808,N_7080,N_7180);
and U7809 (N_7809,N_7203,N_7286);
and U7810 (N_7810,N_7266,N_7183);
nand U7811 (N_7811,N_7472,N_7068);
nand U7812 (N_7812,N_7058,N_7259);
nand U7813 (N_7813,N_7070,N_7104);
nand U7814 (N_7814,N_7235,N_7386);
nor U7815 (N_7815,N_7054,N_7310);
xor U7816 (N_7816,N_7291,N_7445);
nor U7817 (N_7817,N_7151,N_7107);
and U7818 (N_7818,N_7082,N_7293);
and U7819 (N_7819,N_7229,N_7294);
or U7820 (N_7820,N_7210,N_7125);
or U7821 (N_7821,N_7369,N_7124);
and U7822 (N_7822,N_7458,N_7090);
and U7823 (N_7823,N_7037,N_7356);
nor U7824 (N_7824,N_7407,N_7269);
xnor U7825 (N_7825,N_7323,N_7408);
nor U7826 (N_7826,N_7417,N_7268);
nor U7827 (N_7827,N_7423,N_7452);
xor U7828 (N_7828,N_7093,N_7130);
nand U7829 (N_7829,N_7393,N_7193);
and U7830 (N_7830,N_7304,N_7398);
xnor U7831 (N_7831,N_7186,N_7299);
or U7832 (N_7832,N_7219,N_7215);
or U7833 (N_7833,N_7469,N_7422);
and U7834 (N_7834,N_7301,N_7224);
nand U7835 (N_7835,N_7157,N_7172);
nand U7836 (N_7836,N_7141,N_7035);
nand U7837 (N_7837,N_7257,N_7161);
xor U7838 (N_7838,N_7172,N_7108);
nor U7839 (N_7839,N_7414,N_7235);
nand U7840 (N_7840,N_7418,N_7405);
or U7841 (N_7841,N_7178,N_7370);
or U7842 (N_7842,N_7339,N_7400);
and U7843 (N_7843,N_7030,N_7216);
nand U7844 (N_7844,N_7249,N_7405);
xnor U7845 (N_7845,N_7272,N_7454);
or U7846 (N_7846,N_7132,N_7253);
nand U7847 (N_7847,N_7030,N_7257);
and U7848 (N_7848,N_7497,N_7029);
xnor U7849 (N_7849,N_7426,N_7327);
nor U7850 (N_7850,N_7288,N_7035);
xnor U7851 (N_7851,N_7135,N_7231);
or U7852 (N_7852,N_7129,N_7402);
nand U7853 (N_7853,N_7323,N_7141);
nand U7854 (N_7854,N_7148,N_7368);
or U7855 (N_7855,N_7162,N_7457);
nand U7856 (N_7856,N_7072,N_7336);
or U7857 (N_7857,N_7270,N_7360);
and U7858 (N_7858,N_7352,N_7206);
nand U7859 (N_7859,N_7445,N_7013);
nor U7860 (N_7860,N_7066,N_7036);
and U7861 (N_7861,N_7303,N_7140);
xor U7862 (N_7862,N_7309,N_7485);
xor U7863 (N_7863,N_7022,N_7277);
or U7864 (N_7864,N_7265,N_7132);
xnor U7865 (N_7865,N_7275,N_7194);
xor U7866 (N_7866,N_7163,N_7042);
nand U7867 (N_7867,N_7348,N_7229);
xor U7868 (N_7868,N_7259,N_7286);
and U7869 (N_7869,N_7454,N_7100);
nand U7870 (N_7870,N_7046,N_7101);
or U7871 (N_7871,N_7259,N_7224);
and U7872 (N_7872,N_7002,N_7245);
nand U7873 (N_7873,N_7326,N_7413);
nor U7874 (N_7874,N_7258,N_7161);
and U7875 (N_7875,N_7381,N_7305);
or U7876 (N_7876,N_7010,N_7324);
xor U7877 (N_7877,N_7493,N_7255);
nand U7878 (N_7878,N_7417,N_7017);
and U7879 (N_7879,N_7481,N_7477);
xor U7880 (N_7880,N_7423,N_7132);
nor U7881 (N_7881,N_7004,N_7020);
nor U7882 (N_7882,N_7070,N_7409);
nor U7883 (N_7883,N_7247,N_7069);
nand U7884 (N_7884,N_7379,N_7486);
nor U7885 (N_7885,N_7184,N_7032);
and U7886 (N_7886,N_7252,N_7094);
nor U7887 (N_7887,N_7279,N_7134);
nor U7888 (N_7888,N_7243,N_7376);
xor U7889 (N_7889,N_7045,N_7359);
xor U7890 (N_7890,N_7200,N_7363);
xnor U7891 (N_7891,N_7444,N_7464);
and U7892 (N_7892,N_7146,N_7157);
xor U7893 (N_7893,N_7434,N_7319);
nand U7894 (N_7894,N_7440,N_7024);
and U7895 (N_7895,N_7071,N_7180);
nand U7896 (N_7896,N_7452,N_7199);
and U7897 (N_7897,N_7251,N_7315);
and U7898 (N_7898,N_7278,N_7159);
and U7899 (N_7899,N_7111,N_7335);
xor U7900 (N_7900,N_7133,N_7457);
or U7901 (N_7901,N_7164,N_7115);
or U7902 (N_7902,N_7472,N_7491);
and U7903 (N_7903,N_7484,N_7042);
xnor U7904 (N_7904,N_7252,N_7312);
or U7905 (N_7905,N_7224,N_7011);
nand U7906 (N_7906,N_7285,N_7345);
and U7907 (N_7907,N_7079,N_7499);
nor U7908 (N_7908,N_7145,N_7048);
and U7909 (N_7909,N_7228,N_7014);
and U7910 (N_7910,N_7218,N_7165);
or U7911 (N_7911,N_7190,N_7484);
and U7912 (N_7912,N_7179,N_7098);
nand U7913 (N_7913,N_7047,N_7340);
xor U7914 (N_7914,N_7225,N_7424);
or U7915 (N_7915,N_7176,N_7358);
nor U7916 (N_7916,N_7233,N_7258);
or U7917 (N_7917,N_7439,N_7184);
and U7918 (N_7918,N_7306,N_7028);
and U7919 (N_7919,N_7093,N_7020);
or U7920 (N_7920,N_7286,N_7173);
xor U7921 (N_7921,N_7449,N_7265);
xor U7922 (N_7922,N_7040,N_7350);
or U7923 (N_7923,N_7122,N_7324);
nor U7924 (N_7924,N_7004,N_7302);
nand U7925 (N_7925,N_7381,N_7353);
nor U7926 (N_7926,N_7016,N_7198);
and U7927 (N_7927,N_7057,N_7405);
and U7928 (N_7928,N_7268,N_7003);
nor U7929 (N_7929,N_7272,N_7335);
nand U7930 (N_7930,N_7020,N_7242);
xor U7931 (N_7931,N_7167,N_7275);
nand U7932 (N_7932,N_7094,N_7022);
nand U7933 (N_7933,N_7199,N_7192);
xnor U7934 (N_7934,N_7152,N_7285);
nand U7935 (N_7935,N_7409,N_7273);
and U7936 (N_7936,N_7240,N_7144);
and U7937 (N_7937,N_7237,N_7455);
nor U7938 (N_7938,N_7145,N_7211);
or U7939 (N_7939,N_7252,N_7318);
nand U7940 (N_7940,N_7230,N_7006);
nor U7941 (N_7941,N_7185,N_7026);
or U7942 (N_7942,N_7429,N_7234);
xnor U7943 (N_7943,N_7457,N_7487);
nand U7944 (N_7944,N_7371,N_7381);
and U7945 (N_7945,N_7483,N_7438);
nor U7946 (N_7946,N_7150,N_7395);
xnor U7947 (N_7947,N_7050,N_7360);
nor U7948 (N_7948,N_7033,N_7263);
xnor U7949 (N_7949,N_7312,N_7168);
nor U7950 (N_7950,N_7353,N_7462);
xnor U7951 (N_7951,N_7150,N_7104);
xnor U7952 (N_7952,N_7122,N_7051);
nand U7953 (N_7953,N_7188,N_7217);
or U7954 (N_7954,N_7196,N_7000);
nand U7955 (N_7955,N_7198,N_7181);
or U7956 (N_7956,N_7335,N_7465);
nand U7957 (N_7957,N_7286,N_7007);
nor U7958 (N_7958,N_7463,N_7172);
and U7959 (N_7959,N_7128,N_7152);
xor U7960 (N_7960,N_7091,N_7378);
nor U7961 (N_7961,N_7019,N_7124);
xnor U7962 (N_7962,N_7451,N_7291);
nand U7963 (N_7963,N_7345,N_7411);
nand U7964 (N_7964,N_7414,N_7434);
xnor U7965 (N_7965,N_7180,N_7447);
nand U7966 (N_7966,N_7165,N_7226);
nand U7967 (N_7967,N_7220,N_7126);
nor U7968 (N_7968,N_7286,N_7229);
nand U7969 (N_7969,N_7241,N_7325);
nor U7970 (N_7970,N_7390,N_7403);
and U7971 (N_7971,N_7006,N_7026);
xnor U7972 (N_7972,N_7160,N_7091);
nor U7973 (N_7973,N_7445,N_7224);
and U7974 (N_7974,N_7171,N_7104);
xor U7975 (N_7975,N_7421,N_7286);
or U7976 (N_7976,N_7073,N_7038);
nor U7977 (N_7977,N_7248,N_7370);
and U7978 (N_7978,N_7247,N_7342);
nor U7979 (N_7979,N_7448,N_7446);
xor U7980 (N_7980,N_7055,N_7054);
and U7981 (N_7981,N_7123,N_7124);
nand U7982 (N_7982,N_7264,N_7382);
or U7983 (N_7983,N_7097,N_7034);
and U7984 (N_7984,N_7119,N_7147);
nor U7985 (N_7985,N_7034,N_7135);
nor U7986 (N_7986,N_7256,N_7313);
and U7987 (N_7987,N_7498,N_7437);
nor U7988 (N_7988,N_7378,N_7135);
nand U7989 (N_7989,N_7120,N_7495);
xor U7990 (N_7990,N_7418,N_7179);
xnor U7991 (N_7991,N_7409,N_7249);
or U7992 (N_7992,N_7292,N_7438);
and U7993 (N_7993,N_7125,N_7325);
xnor U7994 (N_7994,N_7190,N_7295);
xnor U7995 (N_7995,N_7293,N_7001);
or U7996 (N_7996,N_7081,N_7135);
nor U7997 (N_7997,N_7241,N_7024);
nor U7998 (N_7998,N_7491,N_7258);
or U7999 (N_7999,N_7140,N_7243);
nor U8000 (N_8000,N_7801,N_7703);
xnor U8001 (N_8001,N_7831,N_7535);
nor U8002 (N_8002,N_7905,N_7805);
xnor U8003 (N_8003,N_7884,N_7862);
or U8004 (N_8004,N_7556,N_7625);
and U8005 (N_8005,N_7798,N_7820);
nor U8006 (N_8006,N_7968,N_7612);
xnor U8007 (N_8007,N_7903,N_7650);
nand U8008 (N_8008,N_7683,N_7666);
and U8009 (N_8009,N_7828,N_7700);
nor U8010 (N_8010,N_7967,N_7607);
or U8011 (N_8011,N_7997,N_7583);
nor U8012 (N_8012,N_7502,N_7649);
xor U8013 (N_8013,N_7540,N_7635);
and U8014 (N_8014,N_7648,N_7986);
or U8015 (N_8015,N_7678,N_7817);
nand U8016 (N_8016,N_7506,N_7926);
and U8017 (N_8017,N_7745,N_7925);
nor U8018 (N_8018,N_7713,N_7933);
xnor U8019 (N_8019,N_7936,N_7748);
xnor U8020 (N_8020,N_7503,N_7841);
and U8021 (N_8021,N_7768,N_7751);
nand U8022 (N_8022,N_7918,N_7771);
nor U8023 (N_8023,N_7657,N_7860);
nor U8024 (N_8024,N_7668,N_7786);
and U8025 (N_8025,N_7576,N_7562);
or U8026 (N_8026,N_7622,N_7646);
nor U8027 (N_8027,N_7911,N_7661);
and U8028 (N_8028,N_7791,N_7842);
or U8029 (N_8029,N_7707,N_7832);
and U8030 (N_8030,N_7715,N_7974);
xor U8031 (N_8031,N_7616,N_7824);
and U8032 (N_8032,N_7906,N_7833);
and U8033 (N_8033,N_7674,N_7916);
or U8034 (N_8034,N_7954,N_7520);
xor U8035 (N_8035,N_7890,N_7898);
nor U8036 (N_8036,N_7597,N_7510);
nor U8037 (N_8037,N_7919,N_7522);
or U8038 (N_8038,N_7682,N_7552);
and U8039 (N_8039,N_7896,N_7807);
and U8040 (N_8040,N_7859,N_7566);
nand U8041 (N_8041,N_7991,N_7928);
nand U8042 (N_8042,N_7721,N_7932);
or U8043 (N_8043,N_7655,N_7543);
xor U8044 (N_8044,N_7636,N_7675);
and U8045 (N_8045,N_7573,N_7923);
nor U8046 (N_8046,N_7688,N_7677);
xor U8047 (N_8047,N_7927,N_7642);
xor U8048 (N_8048,N_7691,N_7763);
and U8049 (N_8049,N_7821,N_7536);
nand U8050 (N_8050,N_7604,N_7901);
xor U8051 (N_8051,N_7571,N_7767);
or U8052 (N_8052,N_7962,N_7652);
and U8053 (N_8053,N_7594,N_7826);
and U8054 (N_8054,N_7812,N_7980);
nor U8055 (N_8055,N_7528,N_7656);
nor U8056 (N_8056,N_7871,N_7957);
and U8057 (N_8057,N_7984,N_7874);
nor U8058 (N_8058,N_7970,N_7982);
nor U8059 (N_8059,N_7727,N_7746);
and U8060 (N_8060,N_7773,N_7972);
xor U8061 (N_8061,N_7961,N_7784);
and U8062 (N_8062,N_7803,N_7846);
or U8063 (N_8063,N_7710,N_7588);
or U8064 (N_8064,N_7837,N_7796);
nor U8065 (N_8065,N_7719,N_7762);
or U8066 (N_8066,N_7910,N_7716);
and U8067 (N_8067,N_7709,N_7789);
xor U8068 (N_8068,N_7659,N_7759);
and U8069 (N_8069,N_7722,N_7813);
or U8070 (N_8070,N_7603,N_7626);
or U8071 (N_8071,N_7868,N_7613);
or U8072 (N_8072,N_7921,N_7814);
and U8073 (N_8073,N_7998,N_7845);
and U8074 (N_8074,N_7836,N_7952);
nor U8075 (N_8075,N_7887,N_7676);
or U8076 (N_8076,N_7627,N_7518);
nor U8077 (N_8077,N_7934,N_7720);
or U8078 (N_8078,N_7823,N_7654);
and U8079 (N_8079,N_7939,N_7985);
nand U8080 (N_8080,N_7662,N_7912);
nor U8081 (N_8081,N_7694,N_7899);
nor U8082 (N_8082,N_7645,N_7660);
and U8083 (N_8083,N_7511,N_7857);
nor U8084 (N_8084,N_7551,N_7882);
or U8085 (N_8085,N_7595,N_7712);
nor U8086 (N_8086,N_7608,N_7940);
or U8087 (N_8087,N_7752,N_7834);
or U8088 (N_8088,N_7711,N_7797);
nand U8089 (N_8089,N_7996,N_7983);
xnor U8090 (N_8090,N_7806,N_7598);
nand U8091 (N_8091,N_7570,N_7815);
or U8092 (N_8092,N_7731,N_7651);
nor U8093 (N_8093,N_7593,N_7760);
xor U8094 (N_8094,N_7769,N_7856);
nand U8095 (N_8095,N_7500,N_7877);
nand U8096 (N_8096,N_7808,N_7705);
nor U8097 (N_8097,N_7900,N_7726);
or U8098 (N_8098,N_7523,N_7718);
and U8099 (N_8099,N_7744,N_7764);
or U8100 (N_8100,N_7809,N_7739);
nand U8101 (N_8101,N_7852,N_7558);
and U8102 (N_8102,N_7581,N_7600);
xor U8103 (N_8103,N_7754,N_7605);
or U8104 (N_8104,N_7867,N_7738);
and U8105 (N_8105,N_7848,N_7737);
xor U8106 (N_8106,N_7541,N_7665);
nor U8107 (N_8107,N_7553,N_7742);
or U8108 (N_8108,N_7819,N_7730);
or U8109 (N_8109,N_7546,N_7561);
nand U8110 (N_8110,N_7617,N_7804);
xnor U8111 (N_8111,N_7942,N_7592);
xnor U8112 (N_8112,N_7792,N_7610);
nor U8113 (N_8113,N_7690,N_7672);
nor U8114 (N_8114,N_7565,N_7865);
nand U8115 (N_8115,N_7881,N_7514);
xnor U8116 (N_8116,N_7517,N_7995);
and U8117 (N_8117,N_7632,N_7790);
nor U8118 (N_8118,N_7647,N_7644);
or U8119 (N_8119,N_7578,N_7620);
nor U8120 (N_8120,N_7555,N_7534);
or U8121 (N_8121,N_7761,N_7658);
nand U8122 (N_8122,N_7964,N_7781);
and U8123 (N_8123,N_7669,N_7689);
nor U8124 (N_8124,N_7878,N_7537);
or U8125 (N_8125,N_7501,N_7866);
and U8126 (N_8126,N_7641,N_7516);
nor U8127 (N_8127,N_7897,N_7929);
or U8128 (N_8128,N_7981,N_7521);
xnor U8129 (N_8129,N_7508,N_7618);
nand U8130 (N_8130,N_7564,N_7750);
and U8131 (N_8131,N_7525,N_7956);
nand U8132 (N_8132,N_7589,N_7944);
nand U8133 (N_8133,N_7855,N_7875);
and U8134 (N_8134,N_7547,N_7863);
nand U8135 (N_8135,N_7671,N_7639);
xnor U8136 (N_8136,N_7992,N_7664);
nor U8137 (N_8137,N_7830,N_7989);
and U8138 (N_8138,N_7596,N_7849);
or U8139 (N_8139,N_7988,N_7854);
nand U8140 (N_8140,N_7844,N_7920);
xor U8141 (N_8141,N_7969,N_7851);
nand U8142 (N_8142,N_7704,N_7930);
nor U8143 (N_8143,N_7788,N_7601);
xnor U8144 (N_8144,N_7714,N_7567);
or U8145 (N_8145,N_7701,N_7542);
nand U8146 (N_8146,N_7765,N_7976);
nand U8147 (N_8147,N_7895,N_7515);
xnor U8148 (N_8148,N_7958,N_7870);
nand U8149 (N_8149,N_7602,N_7614);
nor U8150 (N_8150,N_7953,N_7586);
nor U8151 (N_8151,N_7913,N_7966);
nand U8152 (N_8152,N_7734,N_7825);
and U8153 (N_8153,N_7590,N_7949);
nor U8154 (N_8154,N_7959,N_7822);
nand U8155 (N_8155,N_7987,N_7680);
or U8156 (N_8156,N_7548,N_7785);
or U8157 (N_8157,N_7779,N_7615);
nand U8158 (N_8158,N_7793,N_7640);
or U8159 (N_8159,N_7638,N_7810);
or U8160 (N_8160,N_7915,N_7973);
nor U8161 (N_8161,N_7717,N_7941);
and U8162 (N_8162,N_7579,N_7584);
or U8163 (N_8163,N_7698,N_7559);
nand U8164 (N_8164,N_7893,N_7663);
or U8165 (N_8165,N_7917,N_7971);
or U8166 (N_8166,N_7741,N_7530);
and U8167 (N_8167,N_7529,N_7747);
and U8168 (N_8168,N_7743,N_7609);
or U8169 (N_8169,N_7544,N_7606);
and U8170 (N_8170,N_7943,N_7643);
xnor U8171 (N_8171,N_7740,N_7840);
nand U8172 (N_8172,N_7977,N_7766);
nand U8173 (N_8173,N_7587,N_7550);
and U8174 (N_8174,N_7706,N_7776);
or U8175 (N_8175,N_7724,N_7795);
or U8176 (N_8176,N_7729,N_7945);
and U8177 (N_8177,N_7507,N_7619);
or U8178 (N_8178,N_7653,N_7774);
nor U8179 (N_8179,N_7802,N_7847);
and U8180 (N_8180,N_7637,N_7876);
and U8181 (N_8181,N_7880,N_7693);
or U8182 (N_8182,N_7582,N_7549);
and U8183 (N_8183,N_7756,N_7532);
nor U8184 (N_8184,N_7979,N_7699);
and U8185 (N_8185,N_7839,N_7799);
xnor U8186 (N_8186,N_7753,N_7891);
and U8187 (N_8187,N_7557,N_7554);
or U8188 (N_8188,N_7736,N_7946);
or U8189 (N_8189,N_7563,N_7835);
and U8190 (N_8190,N_7950,N_7770);
and U8191 (N_8191,N_7960,N_7686);
and U8192 (N_8192,N_7585,N_7697);
or U8193 (N_8193,N_7872,N_7978);
or U8194 (N_8194,N_7560,N_7907);
or U8195 (N_8195,N_7629,N_7512);
nor U8196 (N_8196,N_7955,N_7667);
xnor U8197 (N_8197,N_7965,N_7990);
and U8198 (N_8198,N_7963,N_7908);
and U8199 (N_8199,N_7818,N_7599);
and U8200 (N_8200,N_7937,N_7999);
nand U8201 (N_8201,N_7947,N_7513);
nand U8202 (N_8202,N_7850,N_7811);
nor U8203 (N_8203,N_7994,N_7504);
xnor U8204 (N_8204,N_7621,N_7904);
nand U8205 (N_8205,N_7948,N_7755);
or U8206 (N_8206,N_7684,N_7695);
nand U8207 (N_8207,N_7538,N_7782);
xnor U8208 (N_8208,N_7922,N_7681);
xnor U8209 (N_8209,N_7531,N_7780);
nand U8210 (N_8210,N_7894,N_7758);
nand U8211 (N_8211,N_7509,N_7838);
nor U8212 (N_8212,N_7843,N_7539);
xor U8213 (N_8213,N_7591,N_7794);
nand U8214 (N_8214,N_7885,N_7864);
xor U8215 (N_8215,N_7829,N_7827);
and U8216 (N_8216,N_7909,N_7735);
and U8217 (N_8217,N_7902,N_7519);
or U8218 (N_8218,N_7670,N_7630);
nand U8219 (N_8219,N_7889,N_7631);
and U8220 (N_8220,N_7853,N_7732);
xor U8221 (N_8221,N_7924,N_7931);
nor U8222 (N_8222,N_7938,N_7858);
and U8223 (N_8223,N_7611,N_7775);
xnor U8224 (N_8224,N_7783,N_7708);
and U8225 (N_8225,N_7505,N_7728);
nor U8226 (N_8226,N_7935,N_7568);
nor U8227 (N_8227,N_7533,N_7778);
and U8228 (N_8228,N_7526,N_7577);
and U8229 (N_8229,N_7725,N_7527);
and U8230 (N_8230,N_7574,N_7623);
or U8231 (N_8231,N_7861,N_7624);
and U8232 (N_8232,N_7886,N_7673);
nor U8233 (N_8233,N_7575,N_7580);
or U8234 (N_8234,N_7892,N_7749);
xor U8235 (N_8235,N_7951,N_7545);
nor U8236 (N_8236,N_7634,N_7883);
nand U8237 (N_8237,N_7816,N_7873);
nor U8238 (N_8238,N_7975,N_7777);
xnor U8239 (N_8239,N_7800,N_7914);
nand U8240 (N_8240,N_7685,N_7687);
nor U8241 (N_8241,N_7993,N_7879);
nor U8242 (N_8242,N_7733,N_7633);
nor U8243 (N_8243,N_7628,N_7679);
and U8244 (N_8244,N_7692,N_7888);
or U8245 (N_8245,N_7869,N_7572);
xor U8246 (N_8246,N_7524,N_7787);
and U8247 (N_8247,N_7757,N_7696);
nand U8248 (N_8248,N_7569,N_7772);
or U8249 (N_8249,N_7702,N_7723);
nor U8250 (N_8250,N_7799,N_7929);
and U8251 (N_8251,N_7740,N_7506);
or U8252 (N_8252,N_7566,N_7941);
nand U8253 (N_8253,N_7746,N_7643);
and U8254 (N_8254,N_7583,N_7797);
nand U8255 (N_8255,N_7565,N_7800);
and U8256 (N_8256,N_7733,N_7903);
and U8257 (N_8257,N_7789,N_7539);
xnor U8258 (N_8258,N_7537,N_7598);
nand U8259 (N_8259,N_7744,N_7837);
nor U8260 (N_8260,N_7664,N_7548);
nand U8261 (N_8261,N_7554,N_7556);
nor U8262 (N_8262,N_7524,N_7988);
nor U8263 (N_8263,N_7986,N_7772);
or U8264 (N_8264,N_7713,N_7717);
nand U8265 (N_8265,N_7643,N_7917);
nand U8266 (N_8266,N_7849,N_7813);
xnor U8267 (N_8267,N_7739,N_7547);
nand U8268 (N_8268,N_7501,N_7946);
xnor U8269 (N_8269,N_7584,N_7733);
nor U8270 (N_8270,N_7746,N_7785);
nor U8271 (N_8271,N_7574,N_7591);
nor U8272 (N_8272,N_7663,N_7825);
or U8273 (N_8273,N_7570,N_7906);
nand U8274 (N_8274,N_7991,N_7673);
nand U8275 (N_8275,N_7763,N_7942);
nor U8276 (N_8276,N_7591,N_7957);
and U8277 (N_8277,N_7647,N_7988);
and U8278 (N_8278,N_7788,N_7920);
xnor U8279 (N_8279,N_7648,N_7923);
and U8280 (N_8280,N_7916,N_7812);
nor U8281 (N_8281,N_7751,N_7992);
or U8282 (N_8282,N_7824,N_7746);
nand U8283 (N_8283,N_7706,N_7504);
and U8284 (N_8284,N_7847,N_7727);
or U8285 (N_8285,N_7679,N_7735);
or U8286 (N_8286,N_7654,N_7728);
xnor U8287 (N_8287,N_7516,N_7832);
nor U8288 (N_8288,N_7713,N_7639);
nor U8289 (N_8289,N_7541,N_7965);
nand U8290 (N_8290,N_7666,N_7900);
nor U8291 (N_8291,N_7773,N_7775);
nor U8292 (N_8292,N_7864,N_7945);
and U8293 (N_8293,N_7970,N_7564);
and U8294 (N_8294,N_7689,N_7711);
and U8295 (N_8295,N_7671,N_7777);
nor U8296 (N_8296,N_7925,N_7744);
nand U8297 (N_8297,N_7582,N_7609);
or U8298 (N_8298,N_7919,N_7570);
nor U8299 (N_8299,N_7889,N_7797);
nand U8300 (N_8300,N_7775,N_7692);
nand U8301 (N_8301,N_7754,N_7786);
or U8302 (N_8302,N_7921,N_7556);
nand U8303 (N_8303,N_7565,N_7651);
nand U8304 (N_8304,N_7598,N_7906);
or U8305 (N_8305,N_7584,N_7766);
nand U8306 (N_8306,N_7867,N_7663);
nor U8307 (N_8307,N_7839,N_7627);
nand U8308 (N_8308,N_7906,N_7591);
and U8309 (N_8309,N_7969,N_7556);
nand U8310 (N_8310,N_7968,N_7534);
and U8311 (N_8311,N_7772,N_7816);
or U8312 (N_8312,N_7925,N_7678);
nand U8313 (N_8313,N_7927,N_7607);
nand U8314 (N_8314,N_7586,N_7788);
or U8315 (N_8315,N_7581,N_7977);
nand U8316 (N_8316,N_7911,N_7561);
or U8317 (N_8317,N_7574,N_7981);
nor U8318 (N_8318,N_7698,N_7617);
or U8319 (N_8319,N_7565,N_7840);
nor U8320 (N_8320,N_7506,N_7573);
xor U8321 (N_8321,N_7594,N_7971);
xor U8322 (N_8322,N_7906,N_7658);
nor U8323 (N_8323,N_7627,N_7656);
nand U8324 (N_8324,N_7614,N_7818);
xnor U8325 (N_8325,N_7869,N_7699);
or U8326 (N_8326,N_7568,N_7607);
xnor U8327 (N_8327,N_7916,N_7576);
nor U8328 (N_8328,N_7711,N_7775);
and U8329 (N_8329,N_7589,N_7886);
nand U8330 (N_8330,N_7869,N_7717);
xor U8331 (N_8331,N_7995,N_7927);
xnor U8332 (N_8332,N_7648,N_7586);
xnor U8333 (N_8333,N_7589,N_7709);
or U8334 (N_8334,N_7827,N_7997);
xnor U8335 (N_8335,N_7731,N_7947);
or U8336 (N_8336,N_7563,N_7999);
xor U8337 (N_8337,N_7689,N_7875);
xnor U8338 (N_8338,N_7617,N_7991);
xor U8339 (N_8339,N_7524,N_7535);
and U8340 (N_8340,N_7748,N_7597);
nor U8341 (N_8341,N_7543,N_7632);
nand U8342 (N_8342,N_7794,N_7684);
or U8343 (N_8343,N_7610,N_7839);
nand U8344 (N_8344,N_7866,N_7875);
xnor U8345 (N_8345,N_7679,N_7844);
xnor U8346 (N_8346,N_7960,N_7684);
nor U8347 (N_8347,N_7710,N_7855);
nand U8348 (N_8348,N_7604,N_7556);
xor U8349 (N_8349,N_7876,N_7532);
nand U8350 (N_8350,N_7901,N_7790);
or U8351 (N_8351,N_7700,N_7566);
nand U8352 (N_8352,N_7638,N_7721);
nor U8353 (N_8353,N_7790,N_7832);
nor U8354 (N_8354,N_7558,N_7901);
nor U8355 (N_8355,N_7870,N_7561);
and U8356 (N_8356,N_7793,N_7570);
nand U8357 (N_8357,N_7655,N_7714);
xor U8358 (N_8358,N_7875,N_7533);
and U8359 (N_8359,N_7983,N_7757);
and U8360 (N_8360,N_7926,N_7787);
xor U8361 (N_8361,N_7590,N_7736);
and U8362 (N_8362,N_7859,N_7540);
or U8363 (N_8363,N_7982,N_7543);
nand U8364 (N_8364,N_7952,N_7905);
or U8365 (N_8365,N_7607,N_7536);
nand U8366 (N_8366,N_7830,N_7553);
and U8367 (N_8367,N_7725,N_7580);
nor U8368 (N_8368,N_7548,N_7624);
or U8369 (N_8369,N_7505,N_7624);
nand U8370 (N_8370,N_7583,N_7868);
and U8371 (N_8371,N_7646,N_7569);
xnor U8372 (N_8372,N_7716,N_7605);
xor U8373 (N_8373,N_7508,N_7586);
or U8374 (N_8374,N_7705,N_7717);
xnor U8375 (N_8375,N_7673,N_7538);
xnor U8376 (N_8376,N_7964,N_7920);
xor U8377 (N_8377,N_7780,N_7626);
nor U8378 (N_8378,N_7728,N_7588);
xor U8379 (N_8379,N_7719,N_7843);
xor U8380 (N_8380,N_7989,N_7592);
or U8381 (N_8381,N_7823,N_7610);
nand U8382 (N_8382,N_7653,N_7825);
nor U8383 (N_8383,N_7920,N_7546);
xnor U8384 (N_8384,N_7542,N_7578);
or U8385 (N_8385,N_7793,N_7890);
xnor U8386 (N_8386,N_7568,N_7802);
and U8387 (N_8387,N_7542,N_7914);
and U8388 (N_8388,N_7577,N_7842);
nor U8389 (N_8389,N_7684,N_7509);
nor U8390 (N_8390,N_7988,N_7844);
and U8391 (N_8391,N_7603,N_7937);
xor U8392 (N_8392,N_7741,N_7957);
and U8393 (N_8393,N_7614,N_7618);
nor U8394 (N_8394,N_7870,N_7912);
and U8395 (N_8395,N_7894,N_7775);
and U8396 (N_8396,N_7558,N_7906);
or U8397 (N_8397,N_7809,N_7928);
or U8398 (N_8398,N_7604,N_7738);
nand U8399 (N_8399,N_7839,N_7615);
nand U8400 (N_8400,N_7526,N_7667);
nand U8401 (N_8401,N_7618,N_7882);
and U8402 (N_8402,N_7707,N_7543);
and U8403 (N_8403,N_7682,N_7814);
or U8404 (N_8404,N_7558,N_7677);
and U8405 (N_8405,N_7716,N_7995);
xor U8406 (N_8406,N_7649,N_7764);
nor U8407 (N_8407,N_7529,N_7799);
and U8408 (N_8408,N_7653,N_7717);
nor U8409 (N_8409,N_7513,N_7617);
nand U8410 (N_8410,N_7827,N_7782);
or U8411 (N_8411,N_7862,N_7796);
and U8412 (N_8412,N_7545,N_7963);
nand U8413 (N_8413,N_7640,N_7513);
nand U8414 (N_8414,N_7826,N_7852);
and U8415 (N_8415,N_7828,N_7538);
nor U8416 (N_8416,N_7704,N_7902);
nor U8417 (N_8417,N_7924,N_7945);
or U8418 (N_8418,N_7548,N_7551);
nand U8419 (N_8419,N_7772,N_7954);
nand U8420 (N_8420,N_7508,N_7964);
nor U8421 (N_8421,N_7547,N_7913);
and U8422 (N_8422,N_7674,N_7946);
and U8423 (N_8423,N_7805,N_7517);
xor U8424 (N_8424,N_7724,N_7532);
and U8425 (N_8425,N_7596,N_7785);
and U8426 (N_8426,N_7876,N_7875);
and U8427 (N_8427,N_7913,N_7570);
nand U8428 (N_8428,N_7670,N_7856);
xor U8429 (N_8429,N_7590,N_7688);
and U8430 (N_8430,N_7587,N_7689);
and U8431 (N_8431,N_7678,N_7748);
nand U8432 (N_8432,N_7531,N_7895);
nand U8433 (N_8433,N_7952,N_7792);
nand U8434 (N_8434,N_7945,N_7576);
and U8435 (N_8435,N_7565,N_7850);
nor U8436 (N_8436,N_7590,N_7519);
nand U8437 (N_8437,N_7913,N_7870);
or U8438 (N_8438,N_7502,N_7677);
xnor U8439 (N_8439,N_7699,N_7516);
xnor U8440 (N_8440,N_7673,N_7893);
nor U8441 (N_8441,N_7851,N_7511);
nor U8442 (N_8442,N_7657,N_7906);
and U8443 (N_8443,N_7914,N_7669);
xor U8444 (N_8444,N_7981,N_7663);
or U8445 (N_8445,N_7740,N_7638);
nand U8446 (N_8446,N_7779,N_7665);
nor U8447 (N_8447,N_7963,N_7863);
nand U8448 (N_8448,N_7502,N_7838);
and U8449 (N_8449,N_7568,N_7548);
or U8450 (N_8450,N_7944,N_7993);
and U8451 (N_8451,N_7667,N_7789);
nor U8452 (N_8452,N_7636,N_7763);
xnor U8453 (N_8453,N_7971,N_7619);
or U8454 (N_8454,N_7724,N_7728);
xor U8455 (N_8455,N_7967,N_7977);
xnor U8456 (N_8456,N_7537,N_7566);
nor U8457 (N_8457,N_7875,N_7519);
xor U8458 (N_8458,N_7830,N_7661);
or U8459 (N_8459,N_7517,N_7945);
nor U8460 (N_8460,N_7514,N_7900);
xnor U8461 (N_8461,N_7822,N_7703);
or U8462 (N_8462,N_7681,N_7948);
nand U8463 (N_8463,N_7680,N_7548);
xnor U8464 (N_8464,N_7908,N_7792);
or U8465 (N_8465,N_7958,N_7598);
and U8466 (N_8466,N_7504,N_7592);
xor U8467 (N_8467,N_7692,N_7918);
and U8468 (N_8468,N_7773,N_7709);
xor U8469 (N_8469,N_7698,N_7685);
xnor U8470 (N_8470,N_7803,N_7554);
or U8471 (N_8471,N_7983,N_7989);
nand U8472 (N_8472,N_7821,N_7969);
or U8473 (N_8473,N_7560,N_7927);
nand U8474 (N_8474,N_7628,N_7766);
and U8475 (N_8475,N_7534,N_7648);
or U8476 (N_8476,N_7515,N_7524);
and U8477 (N_8477,N_7717,N_7948);
nor U8478 (N_8478,N_7578,N_7716);
nand U8479 (N_8479,N_7730,N_7556);
and U8480 (N_8480,N_7987,N_7671);
or U8481 (N_8481,N_7676,N_7920);
and U8482 (N_8482,N_7795,N_7844);
nor U8483 (N_8483,N_7626,N_7549);
nand U8484 (N_8484,N_7743,N_7742);
or U8485 (N_8485,N_7652,N_7659);
nand U8486 (N_8486,N_7602,N_7768);
nor U8487 (N_8487,N_7501,N_7971);
nand U8488 (N_8488,N_7816,N_7661);
xnor U8489 (N_8489,N_7522,N_7938);
nor U8490 (N_8490,N_7653,N_7952);
xnor U8491 (N_8491,N_7562,N_7858);
and U8492 (N_8492,N_7785,N_7824);
nand U8493 (N_8493,N_7908,N_7523);
and U8494 (N_8494,N_7619,N_7530);
and U8495 (N_8495,N_7500,N_7622);
xnor U8496 (N_8496,N_7609,N_7939);
nor U8497 (N_8497,N_7888,N_7866);
xnor U8498 (N_8498,N_7902,N_7720);
nor U8499 (N_8499,N_7549,N_7727);
and U8500 (N_8500,N_8024,N_8062);
xnor U8501 (N_8501,N_8206,N_8395);
xor U8502 (N_8502,N_8029,N_8084);
or U8503 (N_8503,N_8345,N_8066);
xor U8504 (N_8504,N_8407,N_8163);
xnor U8505 (N_8505,N_8259,N_8362);
or U8506 (N_8506,N_8378,N_8057);
or U8507 (N_8507,N_8482,N_8497);
nor U8508 (N_8508,N_8429,N_8419);
and U8509 (N_8509,N_8307,N_8336);
xnor U8510 (N_8510,N_8221,N_8074);
nand U8511 (N_8511,N_8169,N_8136);
or U8512 (N_8512,N_8243,N_8225);
nor U8513 (N_8513,N_8296,N_8022);
or U8514 (N_8514,N_8071,N_8321);
nor U8515 (N_8515,N_8183,N_8298);
and U8516 (N_8516,N_8190,N_8045);
or U8517 (N_8517,N_8224,N_8073);
nor U8518 (N_8518,N_8116,N_8357);
and U8519 (N_8519,N_8106,N_8326);
xor U8520 (N_8520,N_8317,N_8201);
xor U8521 (N_8521,N_8240,N_8435);
nand U8522 (N_8522,N_8016,N_8314);
and U8523 (N_8523,N_8418,N_8316);
nor U8524 (N_8524,N_8445,N_8196);
xnor U8525 (N_8525,N_8414,N_8396);
nand U8526 (N_8526,N_8188,N_8261);
nand U8527 (N_8527,N_8043,N_8305);
or U8528 (N_8528,N_8175,N_8192);
or U8529 (N_8529,N_8223,N_8454);
nor U8530 (N_8530,N_8064,N_8472);
xnor U8531 (N_8531,N_8462,N_8340);
nor U8532 (N_8532,N_8146,N_8239);
nor U8533 (N_8533,N_8263,N_8214);
and U8534 (N_8534,N_8105,N_8023);
xor U8535 (N_8535,N_8160,N_8095);
nor U8536 (N_8536,N_8274,N_8387);
xnor U8537 (N_8537,N_8158,N_8133);
or U8538 (N_8538,N_8481,N_8000);
and U8539 (N_8539,N_8138,N_8344);
xnor U8540 (N_8540,N_8351,N_8465);
xnor U8541 (N_8541,N_8213,N_8172);
xnor U8542 (N_8542,N_8007,N_8498);
or U8543 (N_8543,N_8083,N_8410);
nor U8544 (N_8544,N_8428,N_8055);
nand U8545 (N_8545,N_8050,N_8255);
nand U8546 (N_8546,N_8207,N_8048);
xor U8547 (N_8547,N_8182,N_8097);
nand U8548 (N_8548,N_8354,N_8186);
and U8549 (N_8549,N_8478,N_8256);
xor U8550 (N_8550,N_8493,N_8438);
nor U8551 (N_8551,N_8211,N_8006);
xor U8552 (N_8552,N_8137,N_8275);
nor U8553 (N_8553,N_8035,N_8003);
nand U8554 (N_8554,N_8315,N_8233);
nor U8555 (N_8555,N_8456,N_8426);
nand U8556 (N_8556,N_8080,N_8290);
and U8557 (N_8557,N_8302,N_8490);
nand U8558 (N_8558,N_8152,N_8331);
xor U8559 (N_8559,N_8355,N_8413);
nor U8560 (N_8560,N_8072,N_8150);
or U8561 (N_8561,N_8432,N_8273);
nand U8562 (N_8562,N_8204,N_8295);
nor U8563 (N_8563,N_8480,N_8085);
xor U8564 (N_8564,N_8185,N_8117);
or U8565 (N_8565,N_8128,N_8360);
or U8566 (N_8566,N_8449,N_8350);
xor U8567 (N_8567,N_8252,N_8087);
nor U8568 (N_8568,N_8247,N_8341);
and U8569 (N_8569,N_8403,N_8191);
nand U8570 (N_8570,N_8184,N_8338);
and U8571 (N_8571,N_8038,N_8492);
or U8572 (N_8572,N_8382,N_8415);
xor U8573 (N_8573,N_8089,N_8384);
and U8574 (N_8574,N_8268,N_8248);
nand U8575 (N_8575,N_8102,N_8303);
xor U8576 (N_8576,N_8283,N_8328);
xnor U8577 (N_8577,N_8494,N_8063);
xor U8578 (N_8578,N_8463,N_8282);
nor U8579 (N_8579,N_8227,N_8078);
or U8580 (N_8580,N_8241,N_8229);
or U8581 (N_8581,N_8455,N_8394);
nor U8582 (N_8582,N_8459,N_8141);
xor U8583 (N_8583,N_8039,N_8200);
xor U8584 (N_8584,N_8004,N_8237);
and U8585 (N_8585,N_8375,N_8260);
nand U8586 (N_8586,N_8156,N_8220);
xnor U8587 (N_8587,N_8193,N_8334);
or U8588 (N_8588,N_8215,N_8297);
nand U8589 (N_8589,N_8070,N_8416);
or U8590 (N_8590,N_8181,N_8325);
or U8591 (N_8591,N_8194,N_8234);
nand U8592 (N_8592,N_8131,N_8242);
or U8593 (N_8593,N_8271,N_8001);
xnor U8594 (N_8594,N_8270,N_8324);
nor U8595 (N_8595,N_8446,N_8244);
nor U8596 (N_8596,N_8470,N_8451);
nand U8597 (N_8597,N_8236,N_8076);
nor U8598 (N_8598,N_8343,N_8028);
nor U8599 (N_8599,N_8369,N_8051);
and U8600 (N_8600,N_8288,N_8139);
xor U8601 (N_8601,N_8042,N_8009);
or U8602 (N_8602,N_8484,N_8420);
nand U8603 (N_8603,N_8232,N_8310);
xnor U8604 (N_8604,N_8319,N_8380);
nand U8605 (N_8605,N_8069,N_8439);
nor U8606 (N_8606,N_8013,N_8230);
nor U8607 (N_8607,N_8312,N_8108);
nand U8608 (N_8608,N_8370,N_8294);
xor U8609 (N_8609,N_8374,N_8311);
nand U8610 (N_8610,N_8276,N_8041);
or U8611 (N_8611,N_8386,N_8499);
xnor U8612 (N_8612,N_8113,N_8166);
nor U8613 (N_8613,N_8352,N_8162);
and U8614 (N_8614,N_8112,N_8301);
or U8615 (N_8615,N_8049,N_8389);
xnor U8616 (N_8616,N_8026,N_8417);
or U8617 (N_8617,N_8266,N_8250);
or U8618 (N_8618,N_8161,N_8176);
xnor U8619 (N_8619,N_8278,N_8358);
and U8620 (N_8620,N_8151,N_8457);
xor U8621 (N_8621,N_8208,N_8329);
xor U8622 (N_8622,N_8281,N_8258);
or U8623 (N_8623,N_8079,N_8460);
nor U8624 (N_8624,N_8412,N_8441);
nand U8625 (N_8625,N_8349,N_8195);
nand U8626 (N_8626,N_8132,N_8167);
nor U8627 (N_8627,N_8202,N_8008);
or U8628 (N_8628,N_8058,N_8199);
xor U8629 (N_8629,N_8265,N_8099);
nand U8630 (N_8630,N_8091,N_8148);
and U8631 (N_8631,N_8385,N_8011);
nor U8632 (N_8632,N_8280,N_8103);
and U8633 (N_8633,N_8368,N_8489);
or U8634 (N_8634,N_8149,N_8450);
xor U8635 (N_8635,N_8020,N_8289);
or U8636 (N_8636,N_8135,N_8123);
nand U8637 (N_8637,N_8306,N_8404);
nand U8638 (N_8638,N_8393,N_8177);
nand U8639 (N_8639,N_8054,N_8322);
xnor U8640 (N_8640,N_8406,N_8052);
nand U8641 (N_8641,N_8264,N_8477);
and U8642 (N_8642,N_8444,N_8381);
nor U8643 (N_8643,N_8122,N_8253);
and U8644 (N_8644,N_8094,N_8143);
xnor U8645 (N_8645,N_8209,N_8483);
nor U8646 (N_8646,N_8238,N_8098);
nor U8647 (N_8647,N_8033,N_8487);
and U8648 (N_8648,N_8053,N_8292);
nand U8649 (N_8649,N_8002,N_8180);
xnor U8650 (N_8650,N_8468,N_8333);
nor U8651 (N_8651,N_8388,N_8170);
or U8652 (N_8652,N_8203,N_8216);
xnor U8653 (N_8653,N_8474,N_8359);
xor U8654 (N_8654,N_8027,N_8473);
nand U8655 (N_8655,N_8347,N_8286);
nor U8656 (N_8656,N_8291,N_8217);
or U8657 (N_8657,N_8452,N_8174);
and U8658 (N_8658,N_8104,N_8372);
nand U8659 (N_8659,N_8440,N_8025);
and U8660 (N_8660,N_8219,N_8017);
xnor U8661 (N_8661,N_8361,N_8005);
nand U8662 (N_8662,N_8115,N_8476);
nor U8663 (N_8663,N_8330,N_8304);
or U8664 (N_8664,N_8390,N_8110);
nor U8665 (N_8665,N_8471,N_8379);
xor U8666 (N_8666,N_8212,N_8399);
xor U8667 (N_8667,N_8398,N_8109);
or U8668 (N_8668,N_8284,N_8145);
or U8669 (N_8669,N_8231,N_8164);
and U8670 (N_8670,N_8431,N_8228);
nand U8671 (N_8671,N_8121,N_8411);
and U8672 (N_8672,N_8165,N_8267);
and U8673 (N_8673,N_8144,N_8142);
xor U8674 (N_8674,N_8218,N_8096);
xor U8675 (N_8675,N_8187,N_8262);
xnor U8676 (N_8676,N_8235,N_8300);
and U8677 (N_8677,N_8125,N_8034);
xor U8678 (N_8678,N_8178,N_8044);
and U8679 (N_8679,N_8434,N_8391);
nor U8680 (N_8680,N_8015,N_8436);
or U8681 (N_8681,N_8285,N_8409);
xnor U8682 (N_8682,N_8111,N_8353);
nand U8683 (N_8683,N_8010,N_8056);
nor U8684 (N_8684,N_8346,N_8040);
nand U8685 (N_8685,N_8100,N_8323);
xor U8686 (N_8686,N_8313,N_8082);
nand U8687 (N_8687,N_8335,N_8342);
and U8688 (N_8688,N_8031,N_8448);
and U8689 (N_8689,N_8422,N_8320);
nand U8690 (N_8690,N_8032,N_8377);
nand U8691 (N_8691,N_8179,N_8447);
nand U8692 (N_8692,N_8257,N_8127);
or U8693 (N_8693,N_8392,N_8383);
or U8694 (N_8694,N_8424,N_8485);
or U8695 (N_8695,N_8293,N_8486);
xor U8696 (N_8696,N_8226,N_8376);
and U8697 (N_8697,N_8437,N_8168);
xor U8698 (N_8698,N_8269,N_8373);
nor U8699 (N_8699,N_8012,N_8060);
nand U8700 (N_8700,N_8205,N_8075);
or U8701 (N_8701,N_8157,N_8086);
or U8702 (N_8702,N_8464,N_8081);
xnor U8703 (N_8703,N_8154,N_8077);
and U8704 (N_8704,N_8332,N_8036);
and U8705 (N_8705,N_8458,N_8400);
nor U8706 (N_8706,N_8118,N_8371);
xor U8707 (N_8707,N_8491,N_8088);
and U8708 (N_8708,N_8065,N_8245);
xnor U8709 (N_8709,N_8129,N_8327);
and U8710 (N_8710,N_8405,N_8363);
xnor U8711 (N_8711,N_8047,N_8249);
xnor U8712 (N_8712,N_8046,N_8272);
nor U8713 (N_8713,N_8356,N_8408);
or U8714 (N_8714,N_8061,N_8014);
and U8715 (N_8715,N_8469,N_8189);
nor U8716 (N_8716,N_8467,N_8495);
nor U8717 (N_8717,N_8308,N_8425);
nor U8718 (N_8718,N_8348,N_8475);
or U8719 (N_8719,N_8130,N_8402);
nor U8720 (N_8720,N_8101,N_8421);
nand U8721 (N_8721,N_8427,N_8153);
nor U8722 (N_8722,N_8246,N_8067);
nand U8723 (N_8723,N_8461,N_8092);
xnor U8724 (N_8724,N_8155,N_8423);
and U8725 (N_8725,N_8037,N_8397);
xor U8726 (N_8726,N_8496,N_8120);
nor U8727 (N_8727,N_8134,N_8299);
or U8728 (N_8728,N_8019,N_8251);
xor U8729 (N_8729,N_8254,N_8366);
xor U8730 (N_8730,N_8318,N_8433);
nand U8731 (N_8731,N_8337,N_8277);
xnor U8732 (N_8732,N_8365,N_8339);
or U8733 (N_8733,N_8488,N_8124);
or U8734 (N_8734,N_8030,N_8197);
or U8735 (N_8735,N_8147,N_8068);
nand U8736 (N_8736,N_8442,N_8021);
xnor U8737 (N_8737,N_8287,N_8114);
nor U8738 (N_8738,N_8126,N_8059);
xor U8739 (N_8739,N_8107,N_8222);
nor U8740 (N_8740,N_8453,N_8198);
and U8741 (N_8741,N_8430,N_8443);
or U8742 (N_8742,N_8171,N_8210);
and U8743 (N_8743,N_8364,N_8018);
or U8744 (N_8744,N_8093,N_8159);
and U8745 (N_8745,N_8090,N_8309);
nor U8746 (N_8746,N_8140,N_8466);
and U8747 (N_8747,N_8479,N_8173);
nor U8748 (N_8748,N_8401,N_8119);
nand U8749 (N_8749,N_8367,N_8279);
nor U8750 (N_8750,N_8208,N_8455);
or U8751 (N_8751,N_8493,N_8412);
nand U8752 (N_8752,N_8298,N_8225);
xnor U8753 (N_8753,N_8173,N_8458);
and U8754 (N_8754,N_8219,N_8368);
xnor U8755 (N_8755,N_8054,N_8329);
nor U8756 (N_8756,N_8197,N_8485);
or U8757 (N_8757,N_8186,N_8092);
and U8758 (N_8758,N_8415,N_8141);
or U8759 (N_8759,N_8279,N_8155);
nand U8760 (N_8760,N_8040,N_8114);
nand U8761 (N_8761,N_8033,N_8468);
xor U8762 (N_8762,N_8343,N_8123);
xnor U8763 (N_8763,N_8050,N_8288);
xor U8764 (N_8764,N_8012,N_8463);
xor U8765 (N_8765,N_8412,N_8046);
xor U8766 (N_8766,N_8115,N_8235);
xnor U8767 (N_8767,N_8476,N_8217);
nor U8768 (N_8768,N_8496,N_8044);
xnor U8769 (N_8769,N_8280,N_8265);
nand U8770 (N_8770,N_8156,N_8425);
nor U8771 (N_8771,N_8243,N_8069);
xnor U8772 (N_8772,N_8219,N_8275);
xor U8773 (N_8773,N_8482,N_8414);
xor U8774 (N_8774,N_8336,N_8031);
nand U8775 (N_8775,N_8188,N_8290);
xor U8776 (N_8776,N_8297,N_8370);
or U8777 (N_8777,N_8387,N_8299);
nand U8778 (N_8778,N_8432,N_8062);
and U8779 (N_8779,N_8384,N_8456);
nor U8780 (N_8780,N_8494,N_8274);
nor U8781 (N_8781,N_8029,N_8477);
and U8782 (N_8782,N_8352,N_8303);
nor U8783 (N_8783,N_8095,N_8266);
and U8784 (N_8784,N_8425,N_8032);
nand U8785 (N_8785,N_8145,N_8290);
and U8786 (N_8786,N_8212,N_8276);
nor U8787 (N_8787,N_8404,N_8249);
nand U8788 (N_8788,N_8155,N_8303);
nor U8789 (N_8789,N_8276,N_8098);
or U8790 (N_8790,N_8009,N_8216);
nand U8791 (N_8791,N_8362,N_8014);
and U8792 (N_8792,N_8474,N_8064);
xor U8793 (N_8793,N_8216,N_8313);
nor U8794 (N_8794,N_8040,N_8270);
nor U8795 (N_8795,N_8423,N_8212);
nand U8796 (N_8796,N_8460,N_8028);
nand U8797 (N_8797,N_8356,N_8484);
nor U8798 (N_8798,N_8112,N_8468);
nor U8799 (N_8799,N_8200,N_8426);
or U8800 (N_8800,N_8340,N_8082);
and U8801 (N_8801,N_8065,N_8492);
or U8802 (N_8802,N_8434,N_8267);
nand U8803 (N_8803,N_8098,N_8329);
nand U8804 (N_8804,N_8466,N_8196);
nand U8805 (N_8805,N_8065,N_8353);
or U8806 (N_8806,N_8281,N_8368);
and U8807 (N_8807,N_8165,N_8406);
or U8808 (N_8808,N_8133,N_8106);
nand U8809 (N_8809,N_8323,N_8003);
and U8810 (N_8810,N_8210,N_8494);
nand U8811 (N_8811,N_8499,N_8142);
nor U8812 (N_8812,N_8284,N_8043);
xor U8813 (N_8813,N_8471,N_8097);
xor U8814 (N_8814,N_8417,N_8124);
or U8815 (N_8815,N_8152,N_8212);
or U8816 (N_8816,N_8047,N_8037);
nand U8817 (N_8817,N_8011,N_8425);
and U8818 (N_8818,N_8101,N_8096);
or U8819 (N_8819,N_8352,N_8070);
nor U8820 (N_8820,N_8159,N_8267);
and U8821 (N_8821,N_8448,N_8140);
and U8822 (N_8822,N_8298,N_8113);
xor U8823 (N_8823,N_8236,N_8240);
nor U8824 (N_8824,N_8153,N_8413);
and U8825 (N_8825,N_8228,N_8038);
and U8826 (N_8826,N_8284,N_8336);
nor U8827 (N_8827,N_8027,N_8026);
nand U8828 (N_8828,N_8451,N_8349);
nor U8829 (N_8829,N_8026,N_8455);
xor U8830 (N_8830,N_8401,N_8142);
xnor U8831 (N_8831,N_8479,N_8285);
or U8832 (N_8832,N_8333,N_8392);
or U8833 (N_8833,N_8400,N_8312);
or U8834 (N_8834,N_8161,N_8400);
xor U8835 (N_8835,N_8215,N_8366);
xnor U8836 (N_8836,N_8381,N_8492);
and U8837 (N_8837,N_8462,N_8232);
and U8838 (N_8838,N_8206,N_8429);
or U8839 (N_8839,N_8265,N_8260);
or U8840 (N_8840,N_8133,N_8006);
nor U8841 (N_8841,N_8112,N_8291);
or U8842 (N_8842,N_8274,N_8049);
or U8843 (N_8843,N_8077,N_8110);
and U8844 (N_8844,N_8115,N_8025);
and U8845 (N_8845,N_8036,N_8433);
and U8846 (N_8846,N_8153,N_8061);
xnor U8847 (N_8847,N_8116,N_8378);
nand U8848 (N_8848,N_8377,N_8133);
nand U8849 (N_8849,N_8473,N_8003);
nor U8850 (N_8850,N_8054,N_8400);
nand U8851 (N_8851,N_8382,N_8341);
xor U8852 (N_8852,N_8414,N_8169);
xor U8853 (N_8853,N_8358,N_8399);
xnor U8854 (N_8854,N_8065,N_8099);
nor U8855 (N_8855,N_8262,N_8003);
nor U8856 (N_8856,N_8006,N_8004);
nor U8857 (N_8857,N_8434,N_8275);
nor U8858 (N_8858,N_8164,N_8249);
nor U8859 (N_8859,N_8248,N_8398);
and U8860 (N_8860,N_8147,N_8362);
nand U8861 (N_8861,N_8275,N_8083);
nand U8862 (N_8862,N_8368,N_8223);
nor U8863 (N_8863,N_8426,N_8255);
xnor U8864 (N_8864,N_8220,N_8350);
or U8865 (N_8865,N_8319,N_8375);
or U8866 (N_8866,N_8026,N_8329);
xnor U8867 (N_8867,N_8404,N_8131);
and U8868 (N_8868,N_8421,N_8137);
nor U8869 (N_8869,N_8323,N_8017);
and U8870 (N_8870,N_8476,N_8039);
or U8871 (N_8871,N_8441,N_8355);
nand U8872 (N_8872,N_8297,N_8174);
nor U8873 (N_8873,N_8228,N_8282);
nor U8874 (N_8874,N_8317,N_8244);
nor U8875 (N_8875,N_8101,N_8261);
and U8876 (N_8876,N_8359,N_8198);
and U8877 (N_8877,N_8304,N_8088);
nand U8878 (N_8878,N_8290,N_8443);
and U8879 (N_8879,N_8289,N_8236);
nand U8880 (N_8880,N_8429,N_8300);
and U8881 (N_8881,N_8424,N_8071);
nor U8882 (N_8882,N_8046,N_8076);
xor U8883 (N_8883,N_8456,N_8272);
or U8884 (N_8884,N_8450,N_8100);
xnor U8885 (N_8885,N_8013,N_8487);
or U8886 (N_8886,N_8357,N_8358);
nor U8887 (N_8887,N_8066,N_8290);
nor U8888 (N_8888,N_8489,N_8097);
or U8889 (N_8889,N_8223,N_8464);
or U8890 (N_8890,N_8392,N_8496);
nor U8891 (N_8891,N_8026,N_8115);
or U8892 (N_8892,N_8336,N_8393);
or U8893 (N_8893,N_8198,N_8079);
and U8894 (N_8894,N_8470,N_8382);
xor U8895 (N_8895,N_8268,N_8138);
nor U8896 (N_8896,N_8024,N_8254);
xor U8897 (N_8897,N_8169,N_8407);
nand U8898 (N_8898,N_8185,N_8227);
and U8899 (N_8899,N_8019,N_8157);
xor U8900 (N_8900,N_8230,N_8229);
and U8901 (N_8901,N_8300,N_8397);
and U8902 (N_8902,N_8054,N_8167);
nor U8903 (N_8903,N_8364,N_8077);
and U8904 (N_8904,N_8307,N_8251);
nor U8905 (N_8905,N_8444,N_8080);
xor U8906 (N_8906,N_8071,N_8054);
nor U8907 (N_8907,N_8007,N_8120);
xnor U8908 (N_8908,N_8143,N_8478);
and U8909 (N_8909,N_8173,N_8280);
nor U8910 (N_8910,N_8075,N_8087);
xor U8911 (N_8911,N_8424,N_8115);
nor U8912 (N_8912,N_8239,N_8219);
xnor U8913 (N_8913,N_8147,N_8159);
xnor U8914 (N_8914,N_8229,N_8365);
and U8915 (N_8915,N_8175,N_8152);
xor U8916 (N_8916,N_8098,N_8355);
or U8917 (N_8917,N_8352,N_8236);
nand U8918 (N_8918,N_8273,N_8485);
nor U8919 (N_8919,N_8290,N_8181);
nor U8920 (N_8920,N_8189,N_8175);
and U8921 (N_8921,N_8498,N_8222);
and U8922 (N_8922,N_8297,N_8229);
xor U8923 (N_8923,N_8067,N_8495);
or U8924 (N_8924,N_8251,N_8009);
or U8925 (N_8925,N_8129,N_8284);
nand U8926 (N_8926,N_8379,N_8355);
or U8927 (N_8927,N_8216,N_8189);
and U8928 (N_8928,N_8114,N_8451);
and U8929 (N_8929,N_8130,N_8126);
and U8930 (N_8930,N_8055,N_8063);
nand U8931 (N_8931,N_8014,N_8160);
and U8932 (N_8932,N_8338,N_8368);
nand U8933 (N_8933,N_8420,N_8026);
nand U8934 (N_8934,N_8132,N_8149);
nand U8935 (N_8935,N_8468,N_8013);
xnor U8936 (N_8936,N_8383,N_8040);
xor U8937 (N_8937,N_8167,N_8494);
and U8938 (N_8938,N_8435,N_8126);
xor U8939 (N_8939,N_8314,N_8347);
and U8940 (N_8940,N_8130,N_8372);
and U8941 (N_8941,N_8099,N_8364);
xnor U8942 (N_8942,N_8079,N_8323);
nor U8943 (N_8943,N_8166,N_8481);
or U8944 (N_8944,N_8065,N_8446);
and U8945 (N_8945,N_8486,N_8033);
nand U8946 (N_8946,N_8033,N_8393);
nor U8947 (N_8947,N_8396,N_8169);
xnor U8948 (N_8948,N_8129,N_8264);
xor U8949 (N_8949,N_8017,N_8178);
nor U8950 (N_8950,N_8314,N_8091);
and U8951 (N_8951,N_8348,N_8127);
xnor U8952 (N_8952,N_8131,N_8264);
or U8953 (N_8953,N_8454,N_8329);
and U8954 (N_8954,N_8394,N_8015);
xor U8955 (N_8955,N_8411,N_8169);
or U8956 (N_8956,N_8440,N_8461);
xnor U8957 (N_8957,N_8135,N_8322);
nor U8958 (N_8958,N_8002,N_8463);
or U8959 (N_8959,N_8007,N_8054);
nor U8960 (N_8960,N_8059,N_8287);
xor U8961 (N_8961,N_8460,N_8414);
xor U8962 (N_8962,N_8123,N_8393);
nor U8963 (N_8963,N_8464,N_8490);
nand U8964 (N_8964,N_8288,N_8022);
or U8965 (N_8965,N_8315,N_8101);
or U8966 (N_8966,N_8148,N_8468);
and U8967 (N_8967,N_8458,N_8197);
nand U8968 (N_8968,N_8147,N_8402);
or U8969 (N_8969,N_8343,N_8456);
and U8970 (N_8970,N_8448,N_8104);
nand U8971 (N_8971,N_8375,N_8437);
or U8972 (N_8972,N_8433,N_8364);
or U8973 (N_8973,N_8000,N_8093);
nand U8974 (N_8974,N_8383,N_8394);
or U8975 (N_8975,N_8358,N_8131);
nand U8976 (N_8976,N_8362,N_8476);
nor U8977 (N_8977,N_8216,N_8390);
xnor U8978 (N_8978,N_8296,N_8274);
xnor U8979 (N_8979,N_8045,N_8168);
and U8980 (N_8980,N_8233,N_8225);
xnor U8981 (N_8981,N_8413,N_8245);
nor U8982 (N_8982,N_8131,N_8185);
or U8983 (N_8983,N_8383,N_8145);
nor U8984 (N_8984,N_8320,N_8358);
and U8985 (N_8985,N_8090,N_8249);
or U8986 (N_8986,N_8465,N_8044);
nor U8987 (N_8987,N_8480,N_8430);
nor U8988 (N_8988,N_8061,N_8082);
nand U8989 (N_8989,N_8330,N_8420);
and U8990 (N_8990,N_8013,N_8284);
nor U8991 (N_8991,N_8454,N_8483);
xnor U8992 (N_8992,N_8025,N_8491);
nor U8993 (N_8993,N_8337,N_8209);
or U8994 (N_8994,N_8306,N_8063);
and U8995 (N_8995,N_8061,N_8026);
or U8996 (N_8996,N_8076,N_8203);
xor U8997 (N_8997,N_8420,N_8193);
nand U8998 (N_8998,N_8132,N_8094);
xnor U8999 (N_8999,N_8169,N_8403);
or U9000 (N_9000,N_8600,N_8956);
and U9001 (N_9001,N_8612,N_8509);
nand U9002 (N_9002,N_8752,N_8959);
nand U9003 (N_9003,N_8503,N_8756);
and U9004 (N_9004,N_8723,N_8868);
and U9005 (N_9005,N_8955,N_8661);
and U9006 (N_9006,N_8584,N_8894);
and U9007 (N_9007,N_8951,N_8987);
nand U9008 (N_9008,N_8844,N_8711);
xnor U9009 (N_9009,N_8765,N_8848);
or U9010 (N_9010,N_8674,N_8950);
nand U9011 (N_9011,N_8753,N_8934);
nor U9012 (N_9012,N_8838,N_8515);
and U9013 (N_9013,N_8738,N_8519);
or U9014 (N_9014,N_8526,N_8918);
and U9015 (N_9015,N_8622,N_8803);
and U9016 (N_9016,N_8912,N_8565);
nand U9017 (N_9017,N_8585,N_8544);
xnor U9018 (N_9018,N_8523,N_8699);
nor U9019 (N_9019,N_8538,N_8801);
or U9020 (N_9020,N_8559,N_8994);
xnor U9021 (N_9021,N_8964,N_8573);
and U9022 (N_9022,N_8802,N_8540);
nand U9023 (N_9023,N_8536,N_8577);
nor U9024 (N_9024,N_8657,N_8676);
xor U9025 (N_9025,N_8599,N_8761);
and U9026 (N_9026,N_8642,N_8804);
xor U9027 (N_9027,N_8941,N_8920);
nor U9028 (N_9028,N_8560,N_8988);
or U9029 (N_9029,N_8973,N_8864);
nand U9030 (N_9030,N_8812,N_8636);
and U9031 (N_9031,N_8703,N_8776);
or U9032 (N_9032,N_8911,N_8645);
xor U9033 (N_9033,N_8879,N_8888);
and U9034 (N_9034,N_8614,N_8827);
nand U9035 (N_9035,N_8714,N_8904);
nand U9036 (N_9036,N_8839,N_8986);
or U9037 (N_9037,N_8913,N_8829);
or U9038 (N_9038,N_8786,N_8579);
nor U9039 (N_9039,N_8866,N_8901);
and U9040 (N_9040,N_8609,N_8917);
nor U9041 (N_9041,N_8887,N_8715);
and U9042 (N_9042,N_8553,N_8795);
xnor U9043 (N_9043,N_8938,N_8834);
nor U9044 (N_9044,N_8905,N_8735);
xnor U9045 (N_9045,N_8744,N_8793);
nor U9046 (N_9046,N_8997,N_8722);
nor U9047 (N_9047,N_8605,N_8851);
or U9048 (N_9048,N_8884,N_8615);
nor U9049 (N_9049,N_8891,N_8800);
and U9050 (N_9050,N_8531,N_8977);
xor U9051 (N_9051,N_8635,N_8721);
or U9052 (N_9052,N_8760,N_8574);
and U9053 (N_9053,N_8820,N_8976);
and U9054 (N_9054,N_8785,N_8683);
and U9055 (N_9055,N_8598,N_8641);
nor U9056 (N_9056,N_8551,N_8548);
and U9057 (N_9057,N_8935,N_8782);
and U9058 (N_9058,N_8880,N_8759);
nand U9059 (N_9059,N_8514,N_8968);
nor U9060 (N_9060,N_8709,N_8885);
nor U9061 (N_9061,N_8613,N_8718);
and U9062 (N_9062,N_8619,N_8936);
or U9063 (N_9063,N_8647,N_8989);
or U9064 (N_9064,N_8773,N_8705);
and U9065 (N_9065,N_8948,N_8652);
nand U9066 (N_9066,N_8763,N_8830);
or U9067 (N_9067,N_8915,N_8807);
xor U9068 (N_9068,N_8682,N_8687);
and U9069 (N_9069,N_8713,N_8638);
or U9070 (N_9070,N_8942,N_8822);
or U9071 (N_9071,N_8798,N_8972);
and U9072 (N_9072,N_8937,N_8805);
xnor U9073 (N_9073,N_8521,N_8589);
xnor U9074 (N_9074,N_8501,N_8766);
nor U9075 (N_9075,N_8663,N_8965);
xnor U9076 (N_9076,N_8762,N_8876);
nor U9077 (N_9077,N_8530,N_8562);
xnor U9078 (N_9078,N_8855,N_8597);
xor U9079 (N_9079,N_8727,N_8872);
or U9080 (N_9080,N_8966,N_8632);
xnor U9081 (N_9081,N_8737,N_8545);
and U9082 (N_9082,N_8960,N_8809);
nand U9083 (N_9083,N_8668,N_8892);
nor U9084 (N_9084,N_8575,N_8555);
or U9085 (N_9085,N_8993,N_8837);
and U9086 (N_9086,N_8666,N_8833);
and U9087 (N_9087,N_8790,N_8607);
xnor U9088 (N_9088,N_8620,N_8821);
and U9089 (N_9089,N_8921,N_8629);
and U9090 (N_9090,N_8750,N_8893);
nor U9091 (N_9091,N_8726,N_8525);
nand U9092 (N_9092,N_8534,N_8845);
and U9093 (N_9093,N_8667,N_8542);
nand U9094 (N_9094,N_8832,N_8507);
xor U9095 (N_9095,N_8724,N_8743);
nand U9096 (N_9096,N_8518,N_8978);
nand U9097 (N_9097,N_8843,N_8995);
and U9098 (N_9098,N_8878,N_8567);
and U9099 (N_9099,N_8967,N_8931);
and U9100 (N_9100,N_8840,N_8811);
or U9101 (N_9101,N_8852,N_8858);
and U9102 (N_9102,N_8586,N_8628);
or U9103 (N_9103,N_8881,N_8546);
nor U9104 (N_9104,N_8588,N_8634);
and U9105 (N_9105,N_8981,N_8857);
or U9106 (N_9106,N_8784,N_8932);
nand U9107 (N_9107,N_8859,N_8982);
nand U9108 (N_9108,N_8949,N_8595);
or U9109 (N_9109,N_8745,N_8922);
nand U9110 (N_9110,N_8617,N_8869);
nor U9111 (N_9111,N_8971,N_8939);
or U9112 (N_9112,N_8513,N_8919);
or U9113 (N_9113,N_8810,N_8865);
and U9114 (N_9114,N_8746,N_8771);
and U9115 (N_9115,N_8680,N_8550);
nor U9116 (N_9116,N_8582,N_8516);
xnor U9117 (N_9117,N_8616,N_8882);
xor U9118 (N_9118,N_8975,N_8849);
or U9119 (N_9119,N_8624,N_8841);
nor U9120 (N_9120,N_8998,N_8506);
or U9121 (N_9121,N_8871,N_8673);
nand U9122 (N_9122,N_8815,N_8603);
xor U9123 (N_9123,N_8946,N_8755);
nand U9124 (N_9124,N_8883,N_8825);
nor U9125 (N_9125,N_8739,N_8954);
nor U9126 (N_9126,N_8625,N_8678);
xor U9127 (N_9127,N_8856,N_8906);
nor U9128 (N_9128,N_8758,N_8899);
xnor U9129 (N_9129,N_8819,N_8779);
or U9130 (N_9130,N_8610,N_8539);
or U9131 (N_9131,N_8929,N_8952);
nand U9132 (N_9132,N_8552,N_8916);
or U9133 (N_9133,N_8863,N_8512);
and U9134 (N_9134,N_8896,N_8770);
and U9135 (N_9135,N_8958,N_8649);
nor U9136 (N_9136,N_8654,N_8716);
and U9137 (N_9137,N_8854,N_8664);
and U9138 (N_9138,N_8653,N_8780);
and U9139 (N_9139,N_8850,N_8842);
nor U9140 (N_9140,N_8626,N_8847);
nand U9141 (N_9141,N_8564,N_8985);
xnor U9142 (N_9142,N_8611,N_8992);
nor U9143 (N_9143,N_8563,N_8731);
nor U9144 (N_9144,N_8720,N_8898);
xnor U9145 (N_9145,N_8940,N_8826);
or U9146 (N_9146,N_8754,N_8717);
xnor U9147 (N_9147,N_8748,N_8510);
xor U9148 (N_9148,N_8511,N_8961);
or U9149 (N_9149,N_8867,N_8658);
nand U9150 (N_9150,N_8925,N_8561);
and U9151 (N_9151,N_8799,N_8873);
and U9152 (N_9152,N_8768,N_8571);
xnor U9153 (N_9153,N_8558,N_8556);
or U9154 (N_9154,N_8631,N_8733);
nor U9155 (N_9155,N_8823,N_8665);
or U9156 (N_9156,N_8902,N_8996);
and U9157 (N_9157,N_8532,N_8816);
nand U9158 (N_9158,N_8914,N_8677);
nor U9159 (N_9159,N_8953,N_8504);
nor U9160 (N_9160,N_8602,N_8923);
nand U9161 (N_9161,N_8728,N_8580);
xnor U9162 (N_9162,N_8907,N_8662);
nand U9163 (N_9163,N_8688,N_8796);
nand U9164 (N_9164,N_8691,N_8508);
or U9165 (N_9165,N_8778,N_8991);
and U9166 (N_9166,N_8643,N_8706);
xor U9167 (N_9167,N_8895,N_8685);
nor U9168 (N_9168,N_8576,N_8660);
nand U9169 (N_9169,N_8983,N_8590);
nand U9170 (N_9170,N_8831,N_8692);
or U9171 (N_9171,N_8529,N_8963);
nor U9172 (N_9172,N_8924,N_8648);
nand U9173 (N_9173,N_8587,N_8690);
xor U9174 (N_9174,N_8569,N_8984);
nor U9175 (N_9175,N_8814,N_8712);
nor U9176 (N_9176,N_8651,N_8694);
nor U9177 (N_9177,N_8862,N_8684);
or U9178 (N_9178,N_8788,N_8719);
nand U9179 (N_9179,N_8775,N_8639);
xnor U9180 (N_9180,N_8897,N_8693);
nand U9181 (N_9181,N_8999,N_8618);
and U9182 (N_9182,N_8772,N_8979);
nor U9183 (N_9183,N_8853,N_8594);
nor U9184 (N_9184,N_8764,N_8926);
nand U9185 (N_9185,N_8945,N_8517);
and U9186 (N_9186,N_8817,N_8524);
xnor U9187 (N_9187,N_8533,N_8974);
nor U9188 (N_9188,N_8543,N_8570);
xor U9189 (N_9189,N_8627,N_8846);
xor U9190 (N_9190,N_8729,N_8725);
nand U9191 (N_9191,N_8608,N_8537);
nor U9192 (N_9192,N_8696,N_8697);
nand U9193 (N_9193,N_8698,N_8623);
and U9194 (N_9194,N_8601,N_8522);
and U9195 (N_9195,N_8704,N_8541);
xor U9196 (N_9196,N_8930,N_8944);
nand U9197 (N_9197,N_8774,N_8943);
and U9198 (N_9198,N_8695,N_8732);
or U9199 (N_9199,N_8679,N_8757);
xor U9200 (N_9200,N_8781,N_8933);
or U9201 (N_9201,N_8908,N_8751);
and U9202 (N_9202,N_8730,N_8910);
xnor U9203 (N_9203,N_8769,N_8630);
xnor U9204 (N_9204,N_8889,N_8606);
nor U9205 (N_9205,N_8500,N_8702);
xnor U9206 (N_9206,N_8672,N_8568);
xnor U9207 (N_9207,N_8836,N_8947);
xor U9208 (N_9208,N_8701,N_8566);
nor U9209 (N_9209,N_8535,N_8797);
and U9210 (N_9210,N_8874,N_8681);
and U9211 (N_9211,N_8783,N_8957);
nand U9212 (N_9212,N_8675,N_8650);
nand U9213 (N_9213,N_8860,N_8813);
and U9214 (N_9214,N_8708,N_8547);
nand U9215 (N_9215,N_8927,N_8794);
xor U9216 (N_9216,N_8669,N_8646);
or U9217 (N_9217,N_8557,N_8604);
nor U9218 (N_9218,N_8824,N_8787);
or U9219 (N_9219,N_8670,N_8791);
nand U9220 (N_9220,N_8789,N_8578);
and U9221 (N_9221,N_8749,N_8520);
or U9222 (N_9222,N_8644,N_8835);
xor U9223 (N_9223,N_8700,N_8740);
or U9224 (N_9224,N_8736,N_8875);
nand U9225 (N_9225,N_8767,N_8808);
nor U9226 (N_9226,N_8710,N_8505);
or U9227 (N_9227,N_8554,N_8792);
and U9228 (N_9228,N_8527,N_8689);
and U9229 (N_9229,N_8962,N_8828);
nor U9230 (N_9230,N_8502,N_8818);
xnor U9231 (N_9231,N_8870,N_8637);
and U9232 (N_9232,N_8671,N_8742);
nor U9233 (N_9233,N_8655,N_8707);
nor U9234 (N_9234,N_8583,N_8980);
nor U9235 (N_9235,N_8581,N_8741);
nor U9236 (N_9236,N_8747,N_8591);
or U9237 (N_9237,N_8990,N_8900);
nand U9238 (N_9238,N_8593,N_8549);
or U9239 (N_9239,N_8806,N_8592);
and U9240 (N_9240,N_8686,N_8886);
and U9241 (N_9241,N_8734,N_8969);
xor U9242 (N_9242,N_8621,N_8970);
xnor U9243 (N_9243,N_8903,N_8633);
or U9244 (N_9244,N_8640,N_8909);
or U9245 (N_9245,N_8572,N_8659);
xor U9246 (N_9246,N_8656,N_8596);
nor U9247 (N_9247,N_8528,N_8928);
and U9248 (N_9248,N_8861,N_8777);
nand U9249 (N_9249,N_8877,N_8890);
and U9250 (N_9250,N_8785,N_8506);
xnor U9251 (N_9251,N_8968,N_8653);
and U9252 (N_9252,N_8712,N_8786);
nor U9253 (N_9253,N_8550,N_8624);
nand U9254 (N_9254,N_8507,N_8583);
and U9255 (N_9255,N_8852,N_8874);
nor U9256 (N_9256,N_8882,N_8975);
nand U9257 (N_9257,N_8597,N_8772);
xor U9258 (N_9258,N_8929,N_8663);
nor U9259 (N_9259,N_8542,N_8583);
nor U9260 (N_9260,N_8585,N_8584);
nor U9261 (N_9261,N_8619,N_8764);
or U9262 (N_9262,N_8779,N_8686);
nor U9263 (N_9263,N_8528,N_8911);
xor U9264 (N_9264,N_8672,N_8644);
and U9265 (N_9265,N_8581,N_8584);
xnor U9266 (N_9266,N_8905,N_8821);
nand U9267 (N_9267,N_8859,N_8735);
or U9268 (N_9268,N_8520,N_8932);
nor U9269 (N_9269,N_8841,N_8899);
nor U9270 (N_9270,N_8934,N_8533);
nand U9271 (N_9271,N_8962,N_8576);
nand U9272 (N_9272,N_8885,N_8749);
nor U9273 (N_9273,N_8524,N_8739);
or U9274 (N_9274,N_8807,N_8516);
nor U9275 (N_9275,N_8964,N_8502);
xor U9276 (N_9276,N_8742,N_8798);
or U9277 (N_9277,N_8676,N_8865);
or U9278 (N_9278,N_8818,N_8878);
nor U9279 (N_9279,N_8843,N_8606);
or U9280 (N_9280,N_8529,N_8569);
nand U9281 (N_9281,N_8662,N_8968);
nand U9282 (N_9282,N_8957,N_8509);
nand U9283 (N_9283,N_8953,N_8554);
nand U9284 (N_9284,N_8907,N_8914);
nor U9285 (N_9285,N_8519,N_8913);
or U9286 (N_9286,N_8708,N_8512);
xor U9287 (N_9287,N_8619,N_8561);
xnor U9288 (N_9288,N_8726,N_8884);
and U9289 (N_9289,N_8535,N_8779);
nand U9290 (N_9290,N_8521,N_8662);
xor U9291 (N_9291,N_8513,N_8537);
nor U9292 (N_9292,N_8533,N_8847);
nor U9293 (N_9293,N_8714,N_8709);
nor U9294 (N_9294,N_8509,N_8581);
and U9295 (N_9295,N_8675,N_8574);
nor U9296 (N_9296,N_8619,N_8954);
xor U9297 (N_9297,N_8682,N_8858);
nor U9298 (N_9298,N_8999,N_8645);
nand U9299 (N_9299,N_8889,N_8670);
nand U9300 (N_9300,N_8940,N_8649);
nor U9301 (N_9301,N_8526,N_8827);
nand U9302 (N_9302,N_8983,N_8651);
and U9303 (N_9303,N_8798,N_8959);
or U9304 (N_9304,N_8934,N_8767);
xnor U9305 (N_9305,N_8870,N_8643);
nand U9306 (N_9306,N_8936,N_8835);
nand U9307 (N_9307,N_8760,N_8781);
nor U9308 (N_9308,N_8504,N_8645);
nand U9309 (N_9309,N_8630,N_8916);
nor U9310 (N_9310,N_8929,N_8617);
xor U9311 (N_9311,N_8820,N_8925);
and U9312 (N_9312,N_8602,N_8766);
nand U9313 (N_9313,N_8995,N_8522);
and U9314 (N_9314,N_8732,N_8904);
nand U9315 (N_9315,N_8896,N_8755);
and U9316 (N_9316,N_8724,N_8783);
xnor U9317 (N_9317,N_8909,N_8523);
xnor U9318 (N_9318,N_8922,N_8819);
and U9319 (N_9319,N_8758,N_8835);
or U9320 (N_9320,N_8850,N_8916);
or U9321 (N_9321,N_8818,N_8912);
or U9322 (N_9322,N_8770,N_8589);
nand U9323 (N_9323,N_8882,N_8854);
xnor U9324 (N_9324,N_8548,N_8525);
xnor U9325 (N_9325,N_8538,N_8822);
xor U9326 (N_9326,N_8829,N_8896);
nor U9327 (N_9327,N_8634,N_8570);
nor U9328 (N_9328,N_8635,N_8513);
xor U9329 (N_9329,N_8548,N_8843);
nor U9330 (N_9330,N_8506,N_8555);
xor U9331 (N_9331,N_8946,N_8677);
or U9332 (N_9332,N_8656,N_8982);
xnor U9333 (N_9333,N_8695,N_8512);
and U9334 (N_9334,N_8932,N_8686);
or U9335 (N_9335,N_8574,N_8558);
xor U9336 (N_9336,N_8650,N_8797);
or U9337 (N_9337,N_8816,N_8707);
nor U9338 (N_9338,N_8815,N_8597);
nand U9339 (N_9339,N_8834,N_8948);
or U9340 (N_9340,N_8811,N_8643);
or U9341 (N_9341,N_8842,N_8973);
and U9342 (N_9342,N_8842,N_8803);
nor U9343 (N_9343,N_8966,N_8627);
nor U9344 (N_9344,N_8719,N_8649);
or U9345 (N_9345,N_8922,N_8591);
and U9346 (N_9346,N_8828,N_8842);
nor U9347 (N_9347,N_8643,N_8923);
xor U9348 (N_9348,N_8770,N_8676);
nor U9349 (N_9349,N_8691,N_8552);
nor U9350 (N_9350,N_8936,N_8512);
and U9351 (N_9351,N_8597,N_8974);
or U9352 (N_9352,N_8709,N_8956);
or U9353 (N_9353,N_8635,N_8631);
or U9354 (N_9354,N_8604,N_8988);
and U9355 (N_9355,N_8823,N_8563);
xnor U9356 (N_9356,N_8555,N_8688);
or U9357 (N_9357,N_8639,N_8547);
or U9358 (N_9358,N_8653,N_8649);
nor U9359 (N_9359,N_8691,N_8786);
nor U9360 (N_9360,N_8875,N_8629);
or U9361 (N_9361,N_8949,N_8657);
or U9362 (N_9362,N_8688,N_8772);
nor U9363 (N_9363,N_8649,N_8963);
or U9364 (N_9364,N_8743,N_8991);
nor U9365 (N_9365,N_8957,N_8813);
or U9366 (N_9366,N_8723,N_8951);
nor U9367 (N_9367,N_8831,N_8977);
or U9368 (N_9368,N_8684,N_8526);
or U9369 (N_9369,N_8555,N_8668);
or U9370 (N_9370,N_8591,N_8759);
nor U9371 (N_9371,N_8833,N_8595);
nor U9372 (N_9372,N_8843,N_8763);
nor U9373 (N_9373,N_8697,N_8765);
and U9374 (N_9374,N_8720,N_8998);
xor U9375 (N_9375,N_8564,N_8632);
xor U9376 (N_9376,N_8610,N_8630);
and U9377 (N_9377,N_8837,N_8652);
or U9378 (N_9378,N_8890,N_8632);
xor U9379 (N_9379,N_8994,N_8723);
or U9380 (N_9380,N_8753,N_8888);
or U9381 (N_9381,N_8847,N_8951);
and U9382 (N_9382,N_8899,N_8677);
nor U9383 (N_9383,N_8710,N_8970);
nor U9384 (N_9384,N_8772,N_8998);
xnor U9385 (N_9385,N_8617,N_8963);
xor U9386 (N_9386,N_8953,N_8587);
nand U9387 (N_9387,N_8914,N_8686);
xor U9388 (N_9388,N_8678,N_8605);
xnor U9389 (N_9389,N_8854,N_8897);
or U9390 (N_9390,N_8694,N_8533);
nand U9391 (N_9391,N_8899,N_8962);
xor U9392 (N_9392,N_8500,N_8845);
or U9393 (N_9393,N_8861,N_8935);
or U9394 (N_9394,N_8995,N_8901);
nand U9395 (N_9395,N_8807,N_8920);
nor U9396 (N_9396,N_8621,N_8915);
and U9397 (N_9397,N_8987,N_8710);
nor U9398 (N_9398,N_8713,N_8998);
nor U9399 (N_9399,N_8688,N_8705);
or U9400 (N_9400,N_8821,N_8780);
and U9401 (N_9401,N_8773,N_8595);
or U9402 (N_9402,N_8913,N_8960);
xnor U9403 (N_9403,N_8660,N_8622);
or U9404 (N_9404,N_8962,N_8865);
and U9405 (N_9405,N_8692,N_8733);
nor U9406 (N_9406,N_8533,N_8540);
or U9407 (N_9407,N_8964,N_8730);
and U9408 (N_9408,N_8989,N_8791);
xnor U9409 (N_9409,N_8709,N_8532);
nor U9410 (N_9410,N_8567,N_8711);
or U9411 (N_9411,N_8848,N_8827);
and U9412 (N_9412,N_8862,N_8936);
and U9413 (N_9413,N_8981,N_8966);
nor U9414 (N_9414,N_8868,N_8737);
xor U9415 (N_9415,N_8882,N_8551);
or U9416 (N_9416,N_8569,N_8992);
xor U9417 (N_9417,N_8928,N_8966);
or U9418 (N_9418,N_8958,N_8857);
and U9419 (N_9419,N_8598,N_8854);
and U9420 (N_9420,N_8850,N_8544);
xor U9421 (N_9421,N_8600,N_8733);
and U9422 (N_9422,N_8916,N_8839);
and U9423 (N_9423,N_8556,N_8588);
nand U9424 (N_9424,N_8517,N_8944);
and U9425 (N_9425,N_8892,N_8641);
nor U9426 (N_9426,N_8990,N_8941);
nand U9427 (N_9427,N_8653,N_8902);
xnor U9428 (N_9428,N_8564,N_8516);
nor U9429 (N_9429,N_8912,N_8629);
nor U9430 (N_9430,N_8656,N_8679);
nor U9431 (N_9431,N_8850,N_8545);
or U9432 (N_9432,N_8940,N_8933);
nor U9433 (N_9433,N_8900,N_8505);
and U9434 (N_9434,N_8658,N_8632);
or U9435 (N_9435,N_8824,N_8845);
nand U9436 (N_9436,N_8707,N_8854);
nand U9437 (N_9437,N_8740,N_8534);
or U9438 (N_9438,N_8751,N_8847);
and U9439 (N_9439,N_8992,N_8997);
or U9440 (N_9440,N_8952,N_8723);
nand U9441 (N_9441,N_8540,N_8731);
xnor U9442 (N_9442,N_8608,N_8725);
nor U9443 (N_9443,N_8697,N_8870);
or U9444 (N_9444,N_8634,N_8650);
xor U9445 (N_9445,N_8691,N_8801);
nor U9446 (N_9446,N_8648,N_8967);
xor U9447 (N_9447,N_8752,N_8837);
nor U9448 (N_9448,N_8997,N_8816);
or U9449 (N_9449,N_8535,N_8634);
or U9450 (N_9450,N_8773,N_8732);
and U9451 (N_9451,N_8549,N_8881);
and U9452 (N_9452,N_8790,N_8842);
nor U9453 (N_9453,N_8913,N_8616);
or U9454 (N_9454,N_8730,N_8560);
or U9455 (N_9455,N_8803,N_8922);
or U9456 (N_9456,N_8532,N_8518);
nand U9457 (N_9457,N_8536,N_8660);
xnor U9458 (N_9458,N_8949,N_8853);
nand U9459 (N_9459,N_8669,N_8832);
xnor U9460 (N_9460,N_8664,N_8966);
nor U9461 (N_9461,N_8866,N_8574);
or U9462 (N_9462,N_8774,N_8604);
nor U9463 (N_9463,N_8740,N_8902);
or U9464 (N_9464,N_8581,N_8648);
xnor U9465 (N_9465,N_8578,N_8798);
nor U9466 (N_9466,N_8777,N_8780);
xor U9467 (N_9467,N_8766,N_8787);
nor U9468 (N_9468,N_8700,N_8534);
nand U9469 (N_9469,N_8774,N_8532);
nand U9470 (N_9470,N_8826,N_8532);
nor U9471 (N_9471,N_8553,N_8675);
xnor U9472 (N_9472,N_8948,N_8787);
and U9473 (N_9473,N_8959,N_8612);
and U9474 (N_9474,N_8934,N_8613);
nor U9475 (N_9475,N_8625,N_8913);
xnor U9476 (N_9476,N_8728,N_8926);
xor U9477 (N_9477,N_8726,N_8761);
or U9478 (N_9478,N_8727,N_8502);
or U9479 (N_9479,N_8919,N_8783);
xor U9480 (N_9480,N_8749,N_8740);
xnor U9481 (N_9481,N_8978,N_8987);
nor U9482 (N_9482,N_8917,N_8824);
or U9483 (N_9483,N_8922,N_8656);
xnor U9484 (N_9484,N_8727,N_8552);
xnor U9485 (N_9485,N_8847,N_8693);
nor U9486 (N_9486,N_8949,N_8715);
and U9487 (N_9487,N_8642,N_8829);
nand U9488 (N_9488,N_8809,N_8683);
or U9489 (N_9489,N_8808,N_8717);
or U9490 (N_9490,N_8758,N_8745);
nor U9491 (N_9491,N_8672,N_8584);
or U9492 (N_9492,N_8826,N_8648);
xnor U9493 (N_9493,N_8606,N_8896);
xnor U9494 (N_9494,N_8934,N_8586);
nor U9495 (N_9495,N_8653,N_8795);
nand U9496 (N_9496,N_8807,N_8949);
nor U9497 (N_9497,N_8886,N_8562);
and U9498 (N_9498,N_8920,N_8780);
nor U9499 (N_9499,N_8553,N_8579);
nand U9500 (N_9500,N_9285,N_9352);
or U9501 (N_9501,N_9320,N_9268);
xnor U9502 (N_9502,N_9478,N_9108);
or U9503 (N_9503,N_9172,N_9357);
and U9504 (N_9504,N_9061,N_9274);
and U9505 (N_9505,N_9000,N_9406);
nor U9506 (N_9506,N_9105,N_9249);
and U9507 (N_9507,N_9411,N_9390);
xor U9508 (N_9508,N_9187,N_9247);
nor U9509 (N_9509,N_9004,N_9388);
and U9510 (N_9510,N_9102,N_9207);
xor U9511 (N_9511,N_9039,N_9259);
and U9512 (N_9512,N_9028,N_9337);
nand U9513 (N_9513,N_9489,N_9446);
xor U9514 (N_9514,N_9188,N_9139);
nand U9515 (N_9515,N_9284,N_9077);
and U9516 (N_9516,N_9303,N_9493);
nand U9517 (N_9517,N_9050,N_9048);
nor U9518 (N_9518,N_9494,N_9286);
and U9519 (N_9519,N_9119,N_9333);
or U9520 (N_9520,N_9385,N_9300);
nand U9521 (N_9521,N_9081,N_9025);
nor U9522 (N_9522,N_9391,N_9047);
nor U9523 (N_9523,N_9323,N_9373);
or U9524 (N_9524,N_9052,N_9153);
or U9525 (N_9525,N_9033,N_9257);
nand U9526 (N_9526,N_9273,N_9218);
and U9527 (N_9527,N_9138,N_9392);
and U9528 (N_9528,N_9194,N_9124);
xor U9529 (N_9529,N_9253,N_9325);
xnor U9530 (N_9530,N_9479,N_9482);
or U9531 (N_9531,N_9023,N_9079);
or U9532 (N_9532,N_9348,N_9024);
or U9533 (N_9533,N_9063,N_9309);
nand U9534 (N_9534,N_9189,N_9227);
nand U9535 (N_9535,N_9184,N_9169);
nor U9536 (N_9536,N_9201,N_9297);
xor U9537 (N_9537,N_9347,N_9476);
nor U9538 (N_9538,N_9318,N_9215);
xor U9539 (N_9539,N_9003,N_9465);
xor U9540 (N_9540,N_9163,N_9487);
xnor U9541 (N_9541,N_9454,N_9130);
and U9542 (N_9542,N_9157,N_9178);
and U9543 (N_9543,N_9020,N_9319);
and U9544 (N_9544,N_9344,N_9151);
xnor U9545 (N_9545,N_9173,N_9426);
nor U9546 (N_9546,N_9302,N_9341);
nor U9547 (N_9547,N_9135,N_9404);
and U9548 (N_9548,N_9382,N_9389);
nand U9549 (N_9549,N_9233,N_9295);
nand U9550 (N_9550,N_9367,N_9156);
nor U9551 (N_9551,N_9304,N_9082);
and U9552 (N_9552,N_9324,N_9013);
nor U9553 (N_9553,N_9236,N_9293);
xnor U9554 (N_9554,N_9275,N_9416);
xor U9555 (N_9555,N_9394,N_9034);
and U9556 (N_9556,N_9093,N_9491);
nor U9557 (N_9557,N_9387,N_9072);
nor U9558 (N_9558,N_9401,N_9451);
xor U9559 (N_9559,N_9434,N_9161);
and U9560 (N_9560,N_9497,N_9095);
and U9561 (N_9561,N_9362,N_9405);
and U9562 (N_9562,N_9204,N_9057);
nor U9563 (N_9563,N_9209,N_9075);
nand U9564 (N_9564,N_9148,N_9179);
xor U9565 (N_9565,N_9042,N_9466);
xnor U9566 (N_9566,N_9355,N_9370);
xnor U9567 (N_9567,N_9035,N_9096);
xnor U9568 (N_9568,N_9398,N_9210);
and U9569 (N_9569,N_9055,N_9089);
xor U9570 (N_9570,N_9032,N_9313);
or U9571 (N_9571,N_9423,N_9384);
and U9572 (N_9572,N_9424,N_9248);
nor U9573 (N_9573,N_9331,N_9483);
or U9574 (N_9574,N_9094,N_9030);
xnor U9575 (N_9575,N_9459,N_9166);
xnor U9576 (N_9576,N_9239,N_9291);
nand U9577 (N_9577,N_9353,N_9338);
nand U9578 (N_9578,N_9164,N_9342);
and U9579 (N_9579,N_9181,N_9321);
nor U9580 (N_9580,N_9059,N_9002);
xnor U9581 (N_9581,N_9414,N_9234);
nand U9582 (N_9582,N_9232,N_9064);
or U9583 (N_9583,N_9141,N_9427);
nand U9584 (N_9584,N_9436,N_9149);
nand U9585 (N_9585,N_9171,N_9073);
and U9586 (N_9586,N_9136,N_9008);
nand U9587 (N_9587,N_9029,N_9216);
xnor U9588 (N_9588,N_9409,N_9441);
and U9589 (N_9589,N_9078,N_9410);
nand U9590 (N_9590,N_9460,N_9018);
or U9591 (N_9591,N_9211,N_9400);
or U9592 (N_9592,N_9340,N_9086);
xor U9593 (N_9593,N_9462,N_9271);
and U9594 (N_9594,N_9174,N_9090);
or U9595 (N_9595,N_9243,N_9343);
nor U9596 (N_9596,N_9241,N_9262);
xor U9597 (N_9597,N_9158,N_9308);
nor U9598 (N_9598,N_9235,N_9246);
nand U9599 (N_9599,N_9397,N_9499);
or U9600 (N_9600,N_9279,N_9069);
xnor U9601 (N_9601,N_9350,N_9422);
nor U9602 (N_9602,N_9365,N_9054);
or U9603 (N_9603,N_9122,N_9457);
nand U9604 (N_9604,N_9464,N_9147);
nand U9605 (N_9605,N_9371,N_9180);
nor U9606 (N_9606,N_9298,N_9165);
and U9607 (N_9607,N_9065,N_9439);
nor U9608 (N_9608,N_9290,N_9126);
nor U9609 (N_9609,N_9408,N_9377);
nand U9610 (N_9610,N_9183,N_9197);
and U9611 (N_9611,N_9175,N_9305);
nor U9612 (N_9612,N_9154,N_9195);
nor U9613 (N_9613,N_9190,N_9244);
nor U9614 (N_9614,N_9425,N_9162);
and U9615 (N_9615,N_9299,N_9440);
and U9616 (N_9616,N_9228,N_9435);
and U9617 (N_9617,N_9229,N_9250);
and U9618 (N_9618,N_9332,N_9326);
and U9619 (N_9619,N_9369,N_9492);
nor U9620 (N_9620,N_9329,N_9134);
and U9621 (N_9621,N_9005,N_9237);
nor U9622 (N_9622,N_9131,N_9038);
xor U9623 (N_9623,N_9264,N_9432);
nand U9624 (N_9624,N_9097,N_9137);
nand U9625 (N_9625,N_9217,N_9354);
or U9626 (N_9626,N_9085,N_9103);
and U9627 (N_9627,N_9222,N_9463);
nand U9628 (N_9628,N_9395,N_9438);
nand U9629 (N_9629,N_9010,N_9027);
xnor U9630 (N_9630,N_9066,N_9345);
and U9631 (N_9631,N_9045,N_9315);
nand U9632 (N_9632,N_9336,N_9402);
nand U9633 (N_9633,N_9040,N_9289);
nand U9634 (N_9634,N_9240,N_9486);
and U9635 (N_9635,N_9037,N_9415);
or U9636 (N_9636,N_9477,N_9068);
xnor U9637 (N_9637,N_9080,N_9220);
xnor U9638 (N_9638,N_9011,N_9144);
nor U9639 (N_9639,N_9112,N_9437);
or U9640 (N_9640,N_9155,N_9396);
nand U9641 (N_9641,N_9001,N_9420);
nand U9642 (N_9642,N_9083,N_9316);
or U9643 (N_9643,N_9356,N_9230);
nor U9644 (N_9644,N_9106,N_9496);
xnor U9645 (N_9645,N_9067,N_9363);
nor U9646 (N_9646,N_9092,N_9480);
or U9647 (N_9647,N_9044,N_9252);
nor U9648 (N_9648,N_9049,N_9288);
nor U9649 (N_9649,N_9242,N_9109);
nor U9650 (N_9650,N_9150,N_9110);
or U9651 (N_9651,N_9191,N_9280);
or U9652 (N_9652,N_9484,N_9115);
and U9653 (N_9653,N_9335,N_9364);
or U9654 (N_9654,N_9260,N_9152);
xor U9655 (N_9655,N_9128,N_9117);
and U9656 (N_9656,N_9430,N_9182);
xor U9657 (N_9657,N_9473,N_9007);
nor U9658 (N_9658,N_9258,N_9413);
or U9659 (N_9659,N_9251,N_9159);
and U9660 (N_9660,N_9375,N_9381);
nand U9661 (N_9661,N_9472,N_9270);
or U9662 (N_9662,N_9403,N_9469);
and U9663 (N_9663,N_9133,N_9121);
xor U9664 (N_9664,N_9084,N_9467);
xor U9665 (N_9665,N_9062,N_9255);
and U9666 (N_9666,N_9100,N_9226);
xnor U9667 (N_9667,N_9202,N_9283);
and U9668 (N_9668,N_9127,N_9143);
nand U9669 (N_9669,N_9186,N_9312);
xor U9670 (N_9670,N_9471,N_9453);
nand U9671 (N_9671,N_9142,N_9417);
and U9672 (N_9672,N_9368,N_9261);
nor U9673 (N_9673,N_9198,N_9118);
and U9674 (N_9674,N_9374,N_9481);
xnor U9675 (N_9675,N_9386,N_9123);
and U9676 (N_9676,N_9287,N_9276);
nor U9677 (N_9677,N_9114,N_9378);
xnor U9678 (N_9678,N_9431,N_9307);
or U9679 (N_9679,N_9495,N_9196);
nand U9680 (N_9680,N_9101,N_9322);
nand U9681 (N_9681,N_9140,N_9455);
nor U9682 (N_9682,N_9224,N_9208);
xor U9683 (N_9683,N_9267,N_9339);
or U9684 (N_9684,N_9301,N_9265);
nor U9685 (N_9685,N_9450,N_9177);
nor U9686 (N_9686,N_9168,N_9419);
or U9687 (N_9687,N_9185,N_9358);
nand U9688 (N_9688,N_9485,N_9263);
nor U9689 (N_9689,N_9372,N_9272);
nand U9690 (N_9690,N_9074,N_9022);
nor U9691 (N_9691,N_9098,N_9266);
xor U9692 (N_9692,N_9418,N_9442);
or U9693 (N_9693,N_9116,N_9311);
or U9694 (N_9694,N_9445,N_9167);
or U9695 (N_9695,N_9379,N_9017);
xor U9696 (N_9696,N_9200,N_9036);
or U9697 (N_9697,N_9129,N_9351);
xnor U9698 (N_9698,N_9015,N_9132);
nor U9699 (N_9699,N_9199,N_9160);
or U9700 (N_9700,N_9328,N_9213);
xnor U9701 (N_9701,N_9366,N_9443);
nand U9702 (N_9702,N_9458,N_9277);
nand U9703 (N_9703,N_9041,N_9359);
nor U9704 (N_9704,N_9125,N_9448);
nor U9705 (N_9705,N_9346,N_9145);
xnor U9706 (N_9706,N_9428,N_9214);
xnor U9707 (N_9707,N_9292,N_9399);
and U9708 (N_9708,N_9053,N_9393);
nor U9709 (N_9709,N_9317,N_9056);
xor U9710 (N_9710,N_9231,N_9021);
nand U9711 (N_9711,N_9349,N_9219);
nor U9712 (N_9712,N_9449,N_9192);
and U9713 (N_9713,N_9281,N_9256);
or U9714 (N_9714,N_9470,N_9444);
nand U9715 (N_9715,N_9314,N_9238);
nor U9716 (N_9716,N_9225,N_9380);
nor U9717 (N_9717,N_9076,N_9310);
nor U9718 (N_9718,N_9203,N_9429);
xnor U9719 (N_9719,N_9334,N_9254);
xor U9720 (N_9720,N_9205,N_9223);
and U9721 (N_9721,N_9245,N_9087);
and U9722 (N_9722,N_9070,N_9488);
and U9723 (N_9723,N_9031,N_9498);
nor U9724 (N_9724,N_9099,N_9206);
nand U9725 (N_9725,N_9058,N_9014);
and U9726 (N_9726,N_9016,N_9412);
nand U9727 (N_9727,N_9327,N_9193);
nand U9728 (N_9728,N_9012,N_9421);
nand U9729 (N_9729,N_9383,N_9104);
xnor U9730 (N_9730,N_9456,N_9269);
nand U9731 (N_9731,N_9407,N_9452);
xnor U9732 (N_9732,N_9330,N_9212);
nor U9733 (N_9733,N_9113,N_9046);
xnor U9734 (N_9734,N_9221,N_9043);
or U9735 (N_9735,N_9009,N_9111);
or U9736 (N_9736,N_9026,N_9170);
xnor U9737 (N_9737,N_9088,N_9306);
nor U9738 (N_9738,N_9060,N_9433);
or U9739 (N_9739,N_9296,N_9468);
nand U9740 (N_9740,N_9006,N_9146);
nor U9741 (N_9741,N_9120,N_9490);
xor U9742 (N_9742,N_9475,N_9294);
xnor U9743 (N_9743,N_9361,N_9019);
nand U9744 (N_9744,N_9376,N_9107);
and U9745 (N_9745,N_9278,N_9071);
nand U9746 (N_9746,N_9282,N_9474);
and U9747 (N_9747,N_9461,N_9091);
xor U9748 (N_9748,N_9447,N_9176);
nand U9749 (N_9749,N_9360,N_9051);
and U9750 (N_9750,N_9085,N_9312);
or U9751 (N_9751,N_9056,N_9362);
nor U9752 (N_9752,N_9042,N_9332);
nor U9753 (N_9753,N_9139,N_9072);
nand U9754 (N_9754,N_9094,N_9420);
nand U9755 (N_9755,N_9476,N_9364);
and U9756 (N_9756,N_9082,N_9246);
nor U9757 (N_9757,N_9010,N_9248);
nor U9758 (N_9758,N_9029,N_9052);
xor U9759 (N_9759,N_9350,N_9029);
or U9760 (N_9760,N_9254,N_9476);
and U9761 (N_9761,N_9364,N_9243);
nand U9762 (N_9762,N_9448,N_9030);
and U9763 (N_9763,N_9450,N_9319);
nand U9764 (N_9764,N_9142,N_9366);
nand U9765 (N_9765,N_9440,N_9384);
and U9766 (N_9766,N_9263,N_9340);
nand U9767 (N_9767,N_9443,N_9266);
and U9768 (N_9768,N_9016,N_9119);
and U9769 (N_9769,N_9325,N_9226);
nor U9770 (N_9770,N_9207,N_9123);
nor U9771 (N_9771,N_9200,N_9126);
nand U9772 (N_9772,N_9337,N_9319);
xor U9773 (N_9773,N_9438,N_9156);
nor U9774 (N_9774,N_9338,N_9027);
or U9775 (N_9775,N_9012,N_9497);
or U9776 (N_9776,N_9059,N_9014);
or U9777 (N_9777,N_9498,N_9185);
and U9778 (N_9778,N_9251,N_9077);
or U9779 (N_9779,N_9492,N_9268);
or U9780 (N_9780,N_9331,N_9268);
or U9781 (N_9781,N_9068,N_9378);
xor U9782 (N_9782,N_9256,N_9107);
nor U9783 (N_9783,N_9236,N_9403);
nor U9784 (N_9784,N_9093,N_9406);
and U9785 (N_9785,N_9102,N_9185);
and U9786 (N_9786,N_9427,N_9027);
nand U9787 (N_9787,N_9444,N_9085);
nor U9788 (N_9788,N_9353,N_9497);
nand U9789 (N_9789,N_9233,N_9256);
xnor U9790 (N_9790,N_9118,N_9366);
or U9791 (N_9791,N_9061,N_9080);
nand U9792 (N_9792,N_9482,N_9288);
nor U9793 (N_9793,N_9033,N_9463);
nand U9794 (N_9794,N_9147,N_9444);
xnor U9795 (N_9795,N_9382,N_9263);
or U9796 (N_9796,N_9499,N_9383);
or U9797 (N_9797,N_9448,N_9282);
nand U9798 (N_9798,N_9342,N_9060);
nor U9799 (N_9799,N_9422,N_9211);
and U9800 (N_9800,N_9294,N_9281);
xnor U9801 (N_9801,N_9226,N_9145);
xor U9802 (N_9802,N_9172,N_9105);
or U9803 (N_9803,N_9231,N_9359);
or U9804 (N_9804,N_9429,N_9178);
nand U9805 (N_9805,N_9403,N_9435);
nand U9806 (N_9806,N_9300,N_9148);
and U9807 (N_9807,N_9346,N_9121);
nor U9808 (N_9808,N_9375,N_9259);
and U9809 (N_9809,N_9072,N_9345);
or U9810 (N_9810,N_9282,N_9445);
xnor U9811 (N_9811,N_9497,N_9453);
or U9812 (N_9812,N_9230,N_9027);
and U9813 (N_9813,N_9289,N_9346);
nor U9814 (N_9814,N_9227,N_9140);
xor U9815 (N_9815,N_9435,N_9094);
and U9816 (N_9816,N_9266,N_9117);
and U9817 (N_9817,N_9261,N_9451);
xor U9818 (N_9818,N_9452,N_9043);
xnor U9819 (N_9819,N_9445,N_9024);
nor U9820 (N_9820,N_9138,N_9189);
and U9821 (N_9821,N_9207,N_9028);
or U9822 (N_9822,N_9169,N_9073);
or U9823 (N_9823,N_9331,N_9340);
xor U9824 (N_9824,N_9368,N_9318);
nand U9825 (N_9825,N_9226,N_9249);
nand U9826 (N_9826,N_9037,N_9330);
or U9827 (N_9827,N_9391,N_9092);
and U9828 (N_9828,N_9194,N_9446);
xnor U9829 (N_9829,N_9416,N_9322);
nand U9830 (N_9830,N_9215,N_9064);
xor U9831 (N_9831,N_9046,N_9029);
nor U9832 (N_9832,N_9428,N_9347);
nor U9833 (N_9833,N_9025,N_9165);
or U9834 (N_9834,N_9348,N_9109);
or U9835 (N_9835,N_9161,N_9331);
and U9836 (N_9836,N_9059,N_9392);
and U9837 (N_9837,N_9150,N_9014);
nand U9838 (N_9838,N_9283,N_9406);
nand U9839 (N_9839,N_9092,N_9413);
nand U9840 (N_9840,N_9277,N_9033);
nor U9841 (N_9841,N_9262,N_9076);
nor U9842 (N_9842,N_9214,N_9263);
and U9843 (N_9843,N_9465,N_9082);
nand U9844 (N_9844,N_9479,N_9308);
or U9845 (N_9845,N_9380,N_9493);
and U9846 (N_9846,N_9036,N_9432);
xor U9847 (N_9847,N_9442,N_9479);
or U9848 (N_9848,N_9430,N_9398);
xor U9849 (N_9849,N_9284,N_9276);
or U9850 (N_9850,N_9351,N_9017);
and U9851 (N_9851,N_9313,N_9191);
nand U9852 (N_9852,N_9351,N_9112);
or U9853 (N_9853,N_9059,N_9258);
or U9854 (N_9854,N_9127,N_9355);
or U9855 (N_9855,N_9296,N_9029);
or U9856 (N_9856,N_9074,N_9251);
nor U9857 (N_9857,N_9358,N_9135);
nor U9858 (N_9858,N_9439,N_9371);
xor U9859 (N_9859,N_9068,N_9450);
or U9860 (N_9860,N_9245,N_9074);
and U9861 (N_9861,N_9087,N_9480);
xnor U9862 (N_9862,N_9058,N_9269);
or U9863 (N_9863,N_9322,N_9305);
nor U9864 (N_9864,N_9308,N_9114);
xnor U9865 (N_9865,N_9174,N_9189);
or U9866 (N_9866,N_9283,N_9266);
or U9867 (N_9867,N_9329,N_9040);
and U9868 (N_9868,N_9403,N_9043);
and U9869 (N_9869,N_9121,N_9492);
or U9870 (N_9870,N_9416,N_9334);
or U9871 (N_9871,N_9421,N_9099);
nand U9872 (N_9872,N_9312,N_9132);
and U9873 (N_9873,N_9021,N_9026);
or U9874 (N_9874,N_9416,N_9177);
and U9875 (N_9875,N_9084,N_9205);
and U9876 (N_9876,N_9426,N_9249);
nor U9877 (N_9877,N_9489,N_9282);
xor U9878 (N_9878,N_9077,N_9351);
or U9879 (N_9879,N_9471,N_9486);
and U9880 (N_9880,N_9022,N_9341);
and U9881 (N_9881,N_9180,N_9434);
xnor U9882 (N_9882,N_9012,N_9373);
nor U9883 (N_9883,N_9328,N_9439);
nand U9884 (N_9884,N_9174,N_9185);
or U9885 (N_9885,N_9335,N_9234);
and U9886 (N_9886,N_9267,N_9153);
and U9887 (N_9887,N_9303,N_9102);
and U9888 (N_9888,N_9444,N_9065);
xor U9889 (N_9889,N_9353,N_9481);
or U9890 (N_9890,N_9410,N_9095);
nor U9891 (N_9891,N_9095,N_9365);
or U9892 (N_9892,N_9342,N_9151);
nor U9893 (N_9893,N_9186,N_9026);
nor U9894 (N_9894,N_9118,N_9228);
xnor U9895 (N_9895,N_9139,N_9165);
nand U9896 (N_9896,N_9004,N_9240);
xor U9897 (N_9897,N_9105,N_9493);
and U9898 (N_9898,N_9055,N_9401);
nand U9899 (N_9899,N_9350,N_9475);
or U9900 (N_9900,N_9281,N_9396);
and U9901 (N_9901,N_9210,N_9277);
xnor U9902 (N_9902,N_9134,N_9114);
nand U9903 (N_9903,N_9240,N_9071);
xnor U9904 (N_9904,N_9494,N_9063);
or U9905 (N_9905,N_9485,N_9419);
or U9906 (N_9906,N_9418,N_9055);
nand U9907 (N_9907,N_9313,N_9426);
nand U9908 (N_9908,N_9019,N_9384);
nor U9909 (N_9909,N_9023,N_9029);
and U9910 (N_9910,N_9339,N_9307);
nor U9911 (N_9911,N_9247,N_9069);
xor U9912 (N_9912,N_9081,N_9374);
nand U9913 (N_9913,N_9184,N_9270);
nor U9914 (N_9914,N_9108,N_9347);
nand U9915 (N_9915,N_9204,N_9403);
and U9916 (N_9916,N_9277,N_9287);
xnor U9917 (N_9917,N_9068,N_9271);
nor U9918 (N_9918,N_9013,N_9331);
xor U9919 (N_9919,N_9033,N_9191);
and U9920 (N_9920,N_9367,N_9250);
xor U9921 (N_9921,N_9324,N_9150);
nor U9922 (N_9922,N_9201,N_9190);
or U9923 (N_9923,N_9224,N_9181);
nor U9924 (N_9924,N_9390,N_9239);
xor U9925 (N_9925,N_9170,N_9017);
nor U9926 (N_9926,N_9007,N_9197);
or U9927 (N_9927,N_9036,N_9407);
nand U9928 (N_9928,N_9049,N_9231);
xnor U9929 (N_9929,N_9401,N_9269);
nor U9930 (N_9930,N_9445,N_9399);
nor U9931 (N_9931,N_9450,N_9055);
nand U9932 (N_9932,N_9446,N_9436);
and U9933 (N_9933,N_9446,N_9078);
xor U9934 (N_9934,N_9332,N_9230);
nand U9935 (N_9935,N_9394,N_9126);
and U9936 (N_9936,N_9301,N_9026);
xor U9937 (N_9937,N_9400,N_9067);
or U9938 (N_9938,N_9108,N_9007);
and U9939 (N_9939,N_9418,N_9106);
xor U9940 (N_9940,N_9033,N_9164);
nand U9941 (N_9941,N_9217,N_9139);
nor U9942 (N_9942,N_9190,N_9382);
nand U9943 (N_9943,N_9137,N_9317);
nand U9944 (N_9944,N_9157,N_9258);
nor U9945 (N_9945,N_9000,N_9368);
nor U9946 (N_9946,N_9095,N_9046);
or U9947 (N_9947,N_9181,N_9320);
xor U9948 (N_9948,N_9078,N_9024);
nor U9949 (N_9949,N_9232,N_9182);
and U9950 (N_9950,N_9292,N_9251);
nand U9951 (N_9951,N_9316,N_9294);
or U9952 (N_9952,N_9221,N_9051);
nand U9953 (N_9953,N_9337,N_9489);
xnor U9954 (N_9954,N_9371,N_9197);
xnor U9955 (N_9955,N_9324,N_9268);
nand U9956 (N_9956,N_9259,N_9171);
or U9957 (N_9957,N_9026,N_9001);
nand U9958 (N_9958,N_9433,N_9125);
or U9959 (N_9959,N_9255,N_9185);
or U9960 (N_9960,N_9312,N_9172);
and U9961 (N_9961,N_9480,N_9402);
or U9962 (N_9962,N_9468,N_9314);
or U9963 (N_9963,N_9347,N_9073);
nand U9964 (N_9964,N_9220,N_9249);
nor U9965 (N_9965,N_9177,N_9146);
nand U9966 (N_9966,N_9109,N_9056);
and U9967 (N_9967,N_9015,N_9294);
xnor U9968 (N_9968,N_9426,N_9139);
and U9969 (N_9969,N_9418,N_9262);
nor U9970 (N_9970,N_9350,N_9445);
and U9971 (N_9971,N_9099,N_9394);
xor U9972 (N_9972,N_9246,N_9349);
or U9973 (N_9973,N_9448,N_9199);
or U9974 (N_9974,N_9313,N_9424);
xor U9975 (N_9975,N_9290,N_9353);
nor U9976 (N_9976,N_9147,N_9251);
nand U9977 (N_9977,N_9068,N_9471);
or U9978 (N_9978,N_9050,N_9030);
nand U9979 (N_9979,N_9283,N_9243);
and U9980 (N_9980,N_9103,N_9411);
or U9981 (N_9981,N_9399,N_9192);
or U9982 (N_9982,N_9038,N_9169);
xnor U9983 (N_9983,N_9418,N_9119);
nand U9984 (N_9984,N_9066,N_9177);
xor U9985 (N_9985,N_9296,N_9059);
nor U9986 (N_9986,N_9035,N_9253);
or U9987 (N_9987,N_9444,N_9318);
and U9988 (N_9988,N_9086,N_9279);
and U9989 (N_9989,N_9034,N_9338);
or U9990 (N_9990,N_9261,N_9002);
xnor U9991 (N_9991,N_9080,N_9344);
xnor U9992 (N_9992,N_9202,N_9159);
and U9993 (N_9993,N_9444,N_9211);
nor U9994 (N_9994,N_9322,N_9160);
nor U9995 (N_9995,N_9136,N_9243);
and U9996 (N_9996,N_9130,N_9479);
xnor U9997 (N_9997,N_9215,N_9249);
or U9998 (N_9998,N_9157,N_9292);
nor U9999 (N_9999,N_9486,N_9289);
nand UO_0 (O_0,N_9780,N_9902);
and UO_1 (O_1,N_9892,N_9698);
nand UO_2 (O_2,N_9757,N_9715);
nor UO_3 (O_3,N_9713,N_9714);
nand UO_4 (O_4,N_9967,N_9838);
xnor UO_5 (O_5,N_9520,N_9742);
or UO_6 (O_6,N_9970,N_9675);
and UO_7 (O_7,N_9626,N_9804);
or UO_8 (O_8,N_9547,N_9997);
nand UO_9 (O_9,N_9894,N_9761);
nand UO_10 (O_10,N_9886,N_9696);
nor UO_11 (O_11,N_9684,N_9994);
and UO_12 (O_12,N_9740,N_9730);
nor UO_13 (O_13,N_9895,N_9922);
nand UO_14 (O_14,N_9578,N_9995);
nand UO_15 (O_15,N_9974,N_9867);
nor UO_16 (O_16,N_9664,N_9975);
nand UO_17 (O_17,N_9687,N_9930);
nand UO_18 (O_18,N_9944,N_9682);
nand UO_19 (O_19,N_9781,N_9782);
or UO_20 (O_20,N_9832,N_9783);
xnor UO_21 (O_21,N_9601,N_9611);
or UO_22 (O_22,N_9795,N_9618);
nand UO_23 (O_23,N_9824,N_9777);
xnor UO_24 (O_24,N_9869,N_9648);
xor UO_25 (O_25,N_9617,N_9670);
nor UO_26 (O_26,N_9656,N_9737);
xnor UO_27 (O_27,N_9848,N_9709);
or UO_28 (O_28,N_9608,N_9548);
nand UO_29 (O_29,N_9645,N_9624);
and UO_30 (O_30,N_9739,N_9514);
nand UO_31 (O_31,N_9841,N_9733);
or UO_32 (O_32,N_9786,N_9502);
nor UO_33 (O_33,N_9529,N_9870);
nor UO_34 (O_34,N_9825,N_9551);
and UO_35 (O_35,N_9985,N_9831);
and UO_36 (O_36,N_9814,N_9758);
xor UO_37 (O_37,N_9691,N_9711);
xnor UO_38 (O_38,N_9999,N_9792);
and UO_39 (O_39,N_9622,N_9968);
xor UO_40 (O_40,N_9508,N_9539);
or UO_41 (O_41,N_9522,N_9540);
nand UO_42 (O_42,N_9532,N_9810);
xor UO_43 (O_43,N_9598,N_9933);
xnor UO_44 (O_44,N_9904,N_9945);
nand UO_45 (O_45,N_9826,N_9557);
and UO_46 (O_46,N_9550,N_9655);
nand UO_47 (O_47,N_9773,N_9785);
and UO_48 (O_48,N_9576,N_9549);
and UO_49 (O_49,N_9596,N_9583);
and UO_50 (O_50,N_9746,N_9720);
xor UO_51 (O_51,N_9573,N_9521);
xor UO_52 (O_52,N_9620,N_9900);
nor UO_53 (O_53,N_9741,N_9574);
and UO_54 (O_54,N_9515,N_9680);
and UO_55 (O_55,N_9558,N_9536);
nor UO_56 (O_56,N_9796,N_9592);
nand UO_57 (O_57,N_9830,N_9669);
xnor UO_58 (O_58,N_9875,N_9585);
or UO_59 (O_59,N_9504,N_9866);
or UO_60 (O_60,N_9602,N_9616);
or UO_61 (O_61,N_9509,N_9523);
or UO_62 (O_62,N_9564,N_9717);
or UO_63 (O_63,N_9980,N_9910);
and UO_64 (O_64,N_9712,N_9914);
xor UO_65 (O_65,N_9543,N_9971);
xnor UO_66 (O_66,N_9513,N_9584);
or UO_67 (O_67,N_9644,N_9978);
xor UO_68 (O_68,N_9721,N_9726);
nand UO_69 (O_69,N_9595,N_9844);
nor UO_70 (O_70,N_9530,N_9766);
xnor UO_71 (O_71,N_9516,N_9633);
and UO_72 (O_72,N_9731,N_9554);
or UO_73 (O_73,N_9984,N_9840);
or UO_74 (O_74,N_9861,N_9525);
and UO_75 (O_75,N_9647,N_9813);
nand UO_76 (O_76,N_9661,N_9623);
or UO_77 (O_77,N_9874,N_9787);
and UO_78 (O_78,N_9562,N_9918);
or UO_79 (O_79,N_9931,N_9628);
or UO_80 (O_80,N_9619,N_9750);
nor UO_81 (O_81,N_9790,N_9560);
and UO_82 (O_82,N_9791,N_9500);
nor UO_83 (O_83,N_9621,N_9969);
or UO_84 (O_84,N_9642,N_9695);
or UO_85 (O_85,N_9986,N_9764);
or UO_86 (O_86,N_9765,N_9754);
nand UO_87 (O_87,N_9565,N_9942);
xnor UO_88 (O_88,N_9939,N_9510);
nand UO_89 (O_89,N_9864,N_9604);
nor UO_90 (O_90,N_9615,N_9660);
xor UO_91 (O_91,N_9819,N_9943);
or UO_92 (O_92,N_9809,N_9563);
and UO_93 (O_93,N_9803,N_9756);
nand UO_94 (O_94,N_9853,N_9883);
or UO_95 (O_95,N_9808,N_9524);
nand UO_96 (O_96,N_9849,N_9772);
nand UO_97 (O_97,N_9950,N_9879);
and UO_98 (O_98,N_9755,N_9991);
and UO_99 (O_99,N_9987,N_9907);
xor UO_100 (O_100,N_9842,N_9799);
or UO_101 (O_101,N_9708,N_9925);
and UO_102 (O_102,N_9589,N_9517);
nor UO_103 (O_103,N_9673,N_9732);
or UO_104 (O_104,N_9724,N_9511);
nand UO_105 (O_105,N_9964,N_9891);
nand UO_106 (O_106,N_9749,N_9581);
nand UO_107 (O_107,N_9685,N_9955);
nand UO_108 (O_108,N_9729,N_9590);
xnor UO_109 (O_109,N_9977,N_9811);
nor UO_110 (O_110,N_9949,N_9863);
and UO_111 (O_111,N_9929,N_9890);
nor UO_112 (O_112,N_9768,N_9896);
and UO_113 (O_113,N_9679,N_9909);
nand UO_114 (O_114,N_9839,N_9632);
xnor UO_115 (O_115,N_9911,N_9920);
nor UO_116 (O_116,N_9659,N_9897);
and UO_117 (O_117,N_9678,N_9747);
nor UO_118 (O_118,N_9802,N_9636);
nor UO_119 (O_119,N_9926,N_9935);
and UO_120 (O_120,N_9881,N_9545);
or UO_121 (O_121,N_9643,N_9940);
xor UO_122 (O_122,N_9658,N_9801);
and UO_123 (O_123,N_9763,N_9577);
nor UO_124 (O_124,N_9899,N_9728);
or UO_125 (O_125,N_9898,N_9917);
nor UO_126 (O_126,N_9976,N_9683);
nand UO_127 (O_127,N_9676,N_9807);
xor UO_128 (O_128,N_9794,N_9889);
or UO_129 (O_129,N_9666,N_9872);
or UO_130 (O_130,N_9805,N_9700);
xor UO_131 (O_131,N_9635,N_9769);
and UO_132 (O_132,N_9927,N_9793);
xnor UO_133 (O_133,N_9921,N_9671);
nor UO_134 (O_134,N_9953,N_9629);
or UO_135 (O_135,N_9934,N_9736);
and UO_136 (O_136,N_9938,N_9851);
nor UO_137 (O_137,N_9871,N_9630);
xor UO_138 (O_138,N_9916,N_9912);
and UO_139 (O_139,N_9653,N_9952);
and UO_140 (O_140,N_9779,N_9705);
nand UO_141 (O_141,N_9996,N_9932);
xnor UO_142 (O_142,N_9963,N_9637);
and UO_143 (O_143,N_9798,N_9770);
and UO_144 (O_144,N_9734,N_9821);
xor UO_145 (O_145,N_9865,N_9690);
nor UO_146 (O_146,N_9778,N_9699);
xnor UO_147 (O_147,N_9552,N_9961);
nand UO_148 (O_148,N_9812,N_9702);
nand UO_149 (O_149,N_9568,N_9582);
nor UO_150 (O_150,N_9919,N_9923);
or UO_151 (O_151,N_9587,N_9639);
and UO_152 (O_152,N_9973,N_9662);
xnor UO_153 (O_153,N_9893,N_9962);
and UO_154 (O_154,N_9519,N_9650);
nand UO_155 (O_155,N_9575,N_9688);
xor UO_156 (O_156,N_9505,N_9860);
xor UO_157 (O_157,N_9579,N_9681);
or UO_158 (O_158,N_9775,N_9607);
or UO_159 (O_159,N_9966,N_9641);
xnor UO_160 (O_160,N_9727,N_9835);
nor UO_161 (O_161,N_9868,N_9905);
xor UO_162 (O_162,N_9706,N_9605);
nand UO_163 (O_163,N_9531,N_9771);
and UO_164 (O_164,N_9836,N_9580);
xor UO_165 (O_165,N_9951,N_9806);
or UO_166 (O_166,N_9906,N_9586);
or UO_167 (O_167,N_9993,N_9937);
xnor UO_168 (O_168,N_9625,N_9846);
xnor UO_169 (O_169,N_9959,N_9957);
or UO_170 (O_170,N_9745,N_9908);
xor UO_171 (O_171,N_9600,N_9816);
nor UO_172 (O_172,N_9990,N_9837);
and UO_173 (O_173,N_9594,N_9762);
nor UO_174 (O_174,N_9834,N_9534);
nor UO_175 (O_175,N_9753,N_9774);
xnor UO_176 (O_176,N_9829,N_9983);
or UO_177 (O_177,N_9913,N_9677);
or UO_178 (O_178,N_9878,N_9651);
and UO_179 (O_179,N_9855,N_9567);
nand UO_180 (O_180,N_9501,N_9631);
or UO_181 (O_181,N_9862,N_9719);
nor UO_182 (O_182,N_9569,N_9668);
nand UO_183 (O_183,N_9704,N_9649);
and UO_184 (O_184,N_9572,N_9760);
xor UO_185 (O_185,N_9689,N_9784);
and UO_186 (O_186,N_9915,N_9946);
nand UO_187 (O_187,N_9665,N_9743);
nor UO_188 (O_188,N_9947,N_9527);
and UO_189 (O_189,N_9697,N_9599);
nand UO_190 (O_190,N_9776,N_9818);
nor UO_191 (O_191,N_9992,N_9627);
or UO_192 (O_192,N_9686,N_9858);
or UO_193 (O_193,N_9887,N_9546);
xor UO_194 (O_194,N_9859,N_9512);
nor UO_195 (O_195,N_9876,N_9960);
or UO_196 (O_196,N_9856,N_9542);
xnor UO_197 (O_197,N_9528,N_9606);
or UO_198 (O_198,N_9748,N_9652);
or UO_199 (O_199,N_9981,N_9537);
nor UO_200 (O_200,N_9877,N_9873);
and UO_201 (O_201,N_9903,N_9610);
and UO_202 (O_202,N_9820,N_9936);
xnor UO_203 (O_203,N_9588,N_9541);
xor UO_204 (O_204,N_9822,N_9710);
nand UO_205 (O_205,N_9634,N_9555);
xnor UO_206 (O_206,N_9956,N_9847);
nor UO_207 (O_207,N_9767,N_9815);
nand UO_208 (O_208,N_9674,N_9998);
and UO_209 (O_209,N_9789,N_9597);
nand UO_210 (O_210,N_9716,N_9751);
or UO_211 (O_211,N_9518,N_9725);
nand UO_212 (O_212,N_9526,N_9718);
or UO_213 (O_213,N_9972,N_9723);
or UO_214 (O_214,N_9566,N_9833);
nand UO_215 (O_215,N_9954,N_9958);
nand UO_216 (O_216,N_9703,N_9735);
xnor UO_217 (O_217,N_9854,N_9928);
nor UO_218 (O_218,N_9857,N_9507);
nor UO_219 (O_219,N_9640,N_9591);
xor UO_220 (O_220,N_9672,N_9800);
or UO_221 (O_221,N_9614,N_9722);
xor UO_222 (O_222,N_9694,N_9657);
nor UO_223 (O_223,N_9752,N_9570);
or UO_224 (O_224,N_9571,N_9982);
nor UO_225 (O_225,N_9603,N_9884);
nand UO_226 (O_226,N_9553,N_9845);
xnor UO_227 (O_227,N_9843,N_9882);
and UO_228 (O_228,N_9759,N_9797);
xnor UO_229 (O_229,N_9593,N_9888);
and UO_230 (O_230,N_9852,N_9559);
nand UO_231 (O_231,N_9988,N_9817);
nor UO_232 (O_232,N_9609,N_9701);
nor UO_233 (O_233,N_9965,N_9646);
or UO_234 (O_234,N_9663,N_9612);
nand UO_235 (O_235,N_9667,N_9613);
nor UO_236 (O_236,N_9561,N_9744);
nand UO_237 (O_237,N_9924,N_9693);
nor UO_238 (O_238,N_9707,N_9828);
nor UO_239 (O_239,N_9788,N_9948);
xnor UO_240 (O_240,N_9506,N_9850);
nand UO_241 (O_241,N_9885,N_9979);
or UO_242 (O_242,N_9544,N_9827);
xnor UO_243 (O_243,N_9738,N_9654);
or UO_244 (O_244,N_9692,N_9533);
or UO_245 (O_245,N_9941,N_9503);
nor UO_246 (O_246,N_9538,N_9638);
nor UO_247 (O_247,N_9535,N_9880);
xnor UO_248 (O_248,N_9901,N_9823);
or UO_249 (O_249,N_9556,N_9989);
nand UO_250 (O_250,N_9572,N_9538);
xnor UO_251 (O_251,N_9915,N_9779);
nor UO_252 (O_252,N_9830,N_9837);
or UO_253 (O_253,N_9825,N_9886);
nor UO_254 (O_254,N_9863,N_9761);
nor UO_255 (O_255,N_9817,N_9767);
nand UO_256 (O_256,N_9871,N_9569);
xnor UO_257 (O_257,N_9964,N_9555);
xor UO_258 (O_258,N_9721,N_9970);
xnor UO_259 (O_259,N_9915,N_9616);
nor UO_260 (O_260,N_9777,N_9675);
xnor UO_261 (O_261,N_9735,N_9847);
nand UO_262 (O_262,N_9789,N_9820);
and UO_263 (O_263,N_9884,N_9879);
nor UO_264 (O_264,N_9502,N_9969);
and UO_265 (O_265,N_9503,N_9883);
and UO_266 (O_266,N_9635,N_9975);
nand UO_267 (O_267,N_9667,N_9661);
nor UO_268 (O_268,N_9957,N_9696);
xor UO_269 (O_269,N_9992,N_9851);
xor UO_270 (O_270,N_9537,N_9766);
or UO_271 (O_271,N_9835,N_9557);
or UO_272 (O_272,N_9979,N_9759);
nand UO_273 (O_273,N_9871,N_9720);
and UO_274 (O_274,N_9958,N_9766);
nor UO_275 (O_275,N_9505,N_9849);
or UO_276 (O_276,N_9845,N_9881);
nor UO_277 (O_277,N_9815,N_9839);
or UO_278 (O_278,N_9887,N_9759);
or UO_279 (O_279,N_9854,N_9520);
xor UO_280 (O_280,N_9780,N_9694);
nor UO_281 (O_281,N_9820,N_9719);
and UO_282 (O_282,N_9545,N_9673);
and UO_283 (O_283,N_9576,N_9916);
and UO_284 (O_284,N_9918,N_9915);
or UO_285 (O_285,N_9920,N_9649);
nor UO_286 (O_286,N_9663,N_9998);
nand UO_287 (O_287,N_9912,N_9825);
nand UO_288 (O_288,N_9612,N_9626);
nor UO_289 (O_289,N_9923,N_9566);
xor UO_290 (O_290,N_9986,N_9658);
nand UO_291 (O_291,N_9816,N_9883);
and UO_292 (O_292,N_9662,N_9525);
nor UO_293 (O_293,N_9654,N_9673);
or UO_294 (O_294,N_9802,N_9502);
and UO_295 (O_295,N_9570,N_9532);
xor UO_296 (O_296,N_9991,N_9537);
or UO_297 (O_297,N_9753,N_9895);
or UO_298 (O_298,N_9900,N_9856);
or UO_299 (O_299,N_9956,N_9931);
or UO_300 (O_300,N_9937,N_9785);
nand UO_301 (O_301,N_9650,N_9703);
xnor UO_302 (O_302,N_9660,N_9748);
xor UO_303 (O_303,N_9657,N_9782);
xnor UO_304 (O_304,N_9511,N_9837);
xor UO_305 (O_305,N_9760,N_9661);
xnor UO_306 (O_306,N_9582,N_9506);
xnor UO_307 (O_307,N_9975,N_9755);
xnor UO_308 (O_308,N_9777,N_9553);
nor UO_309 (O_309,N_9618,N_9883);
and UO_310 (O_310,N_9726,N_9660);
and UO_311 (O_311,N_9706,N_9703);
nor UO_312 (O_312,N_9927,N_9507);
xor UO_313 (O_313,N_9585,N_9674);
nor UO_314 (O_314,N_9689,N_9726);
and UO_315 (O_315,N_9724,N_9700);
or UO_316 (O_316,N_9713,N_9955);
and UO_317 (O_317,N_9897,N_9589);
nand UO_318 (O_318,N_9647,N_9780);
and UO_319 (O_319,N_9939,N_9550);
or UO_320 (O_320,N_9549,N_9685);
nand UO_321 (O_321,N_9871,N_9842);
nor UO_322 (O_322,N_9689,N_9653);
nand UO_323 (O_323,N_9817,N_9822);
nor UO_324 (O_324,N_9577,N_9991);
and UO_325 (O_325,N_9904,N_9544);
or UO_326 (O_326,N_9571,N_9747);
and UO_327 (O_327,N_9963,N_9514);
and UO_328 (O_328,N_9932,N_9694);
or UO_329 (O_329,N_9816,N_9679);
xnor UO_330 (O_330,N_9593,N_9614);
or UO_331 (O_331,N_9700,N_9657);
or UO_332 (O_332,N_9768,N_9583);
xor UO_333 (O_333,N_9729,N_9588);
and UO_334 (O_334,N_9515,N_9733);
nand UO_335 (O_335,N_9609,N_9879);
or UO_336 (O_336,N_9700,N_9705);
and UO_337 (O_337,N_9831,N_9970);
nor UO_338 (O_338,N_9731,N_9598);
nor UO_339 (O_339,N_9615,N_9555);
or UO_340 (O_340,N_9949,N_9634);
nand UO_341 (O_341,N_9562,N_9727);
nand UO_342 (O_342,N_9959,N_9930);
and UO_343 (O_343,N_9744,N_9955);
xnor UO_344 (O_344,N_9592,N_9701);
nor UO_345 (O_345,N_9572,N_9783);
nand UO_346 (O_346,N_9936,N_9894);
nand UO_347 (O_347,N_9934,N_9987);
nor UO_348 (O_348,N_9574,N_9634);
and UO_349 (O_349,N_9627,N_9549);
xor UO_350 (O_350,N_9962,N_9542);
nand UO_351 (O_351,N_9921,N_9579);
nand UO_352 (O_352,N_9722,N_9534);
nand UO_353 (O_353,N_9805,N_9971);
xor UO_354 (O_354,N_9720,N_9556);
nand UO_355 (O_355,N_9796,N_9640);
and UO_356 (O_356,N_9920,N_9642);
nand UO_357 (O_357,N_9613,N_9847);
nand UO_358 (O_358,N_9583,N_9814);
and UO_359 (O_359,N_9980,N_9525);
nand UO_360 (O_360,N_9601,N_9563);
nor UO_361 (O_361,N_9804,N_9602);
nor UO_362 (O_362,N_9538,N_9735);
xor UO_363 (O_363,N_9836,N_9738);
or UO_364 (O_364,N_9884,N_9924);
xor UO_365 (O_365,N_9995,N_9655);
xor UO_366 (O_366,N_9708,N_9518);
and UO_367 (O_367,N_9730,N_9966);
xnor UO_368 (O_368,N_9694,N_9823);
xor UO_369 (O_369,N_9732,N_9623);
or UO_370 (O_370,N_9755,N_9925);
nand UO_371 (O_371,N_9605,N_9792);
and UO_372 (O_372,N_9896,N_9635);
and UO_373 (O_373,N_9538,N_9903);
xnor UO_374 (O_374,N_9599,N_9681);
or UO_375 (O_375,N_9673,N_9603);
and UO_376 (O_376,N_9591,N_9909);
nand UO_377 (O_377,N_9786,N_9908);
and UO_378 (O_378,N_9542,N_9906);
nor UO_379 (O_379,N_9888,N_9856);
nor UO_380 (O_380,N_9722,N_9763);
nor UO_381 (O_381,N_9847,N_9649);
nor UO_382 (O_382,N_9694,N_9769);
and UO_383 (O_383,N_9843,N_9558);
nand UO_384 (O_384,N_9861,N_9713);
or UO_385 (O_385,N_9665,N_9924);
xnor UO_386 (O_386,N_9779,N_9714);
nor UO_387 (O_387,N_9508,N_9613);
and UO_388 (O_388,N_9869,N_9957);
nor UO_389 (O_389,N_9815,N_9588);
and UO_390 (O_390,N_9878,N_9971);
xor UO_391 (O_391,N_9794,N_9555);
xor UO_392 (O_392,N_9842,N_9942);
or UO_393 (O_393,N_9952,N_9821);
and UO_394 (O_394,N_9535,N_9972);
or UO_395 (O_395,N_9852,N_9588);
nand UO_396 (O_396,N_9766,N_9738);
xor UO_397 (O_397,N_9731,N_9505);
and UO_398 (O_398,N_9814,N_9906);
or UO_399 (O_399,N_9694,N_9899);
or UO_400 (O_400,N_9673,N_9725);
and UO_401 (O_401,N_9505,N_9541);
nand UO_402 (O_402,N_9611,N_9624);
nand UO_403 (O_403,N_9690,N_9554);
or UO_404 (O_404,N_9580,N_9920);
xnor UO_405 (O_405,N_9885,N_9884);
nor UO_406 (O_406,N_9581,N_9616);
and UO_407 (O_407,N_9741,N_9546);
xnor UO_408 (O_408,N_9809,N_9582);
and UO_409 (O_409,N_9704,N_9950);
or UO_410 (O_410,N_9792,N_9750);
or UO_411 (O_411,N_9604,N_9539);
nand UO_412 (O_412,N_9923,N_9511);
nor UO_413 (O_413,N_9731,N_9547);
or UO_414 (O_414,N_9500,N_9646);
or UO_415 (O_415,N_9795,N_9808);
nor UO_416 (O_416,N_9617,N_9943);
xor UO_417 (O_417,N_9710,N_9808);
xor UO_418 (O_418,N_9894,N_9812);
nor UO_419 (O_419,N_9595,N_9728);
and UO_420 (O_420,N_9670,N_9946);
nand UO_421 (O_421,N_9885,N_9880);
xor UO_422 (O_422,N_9506,N_9507);
and UO_423 (O_423,N_9835,N_9508);
or UO_424 (O_424,N_9916,N_9641);
nor UO_425 (O_425,N_9775,N_9979);
or UO_426 (O_426,N_9685,N_9787);
or UO_427 (O_427,N_9534,N_9561);
and UO_428 (O_428,N_9537,N_9811);
and UO_429 (O_429,N_9676,N_9581);
nor UO_430 (O_430,N_9557,N_9970);
nand UO_431 (O_431,N_9656,N_9896);
nor UO_432 (O_432,N_9899,N_9591);
or UO_433 (O_433,N_9722,N_9518);
xor UO_434 (O_434,N_9886,N_9535);
xor UO_435 (O_435,N_9665,N_9702);
xnor UO_436 (O_436,N_9853,N_9838);
nand UO_437 (O_437,N_9976,N_9710);
xor UO_438 (O_438,N_9741,N_9931);
and UO_439 (O_439,N_9940,N_9921);
and UO_440 (O_440,N_9532,N_9682);
and UO_441 (O_441,N_9567,N_9929);
nand UO_442 (O_442,N_9911,N_9843);
xor UO_443 (O_443,N_9740,N_9552);
nor UO_444 (O_444,N_9610,N_9754);
nor UO_445 (O_445,N_9598,N_9692);
or UO_446 (O_446,N_9587,N_9696);
or UO_447 (O_447,N_9912,N_9822);
nor UO_448 (O_448,N_9927,N_9751);
or UO_449 (O_449,N_9550,N_9563);
xnor UO_450 (O_450,N_9675,N_9622);
nor UO_451 (O_451,N_9812,N_9720);
and UO_452 (O_452,N_9994,N_9812);
or UO_453 (O_453,N_9668,N_9693);
nor UO_454 (O_454,N_9909,N_9675);
xnor UO_455 (O_455,N_9922,N_9680);
xnor UO_456 (O_456,N_9926,N_9769);
and UO_457 (O_457,N_9809,N_9764);
and UO_458 (O_458,N_9900,N_9548);
xnor UO_459 (O_459,N_9554,N_9641);
nor UO_460 (O_460,N_9896,N_9762);
nor UO_461 (O_461,N_9933,N_9583);
and UO_462 (O_462,N_9546,N_9614);
nor UO_463 (O_463,N_9565,N_9592);
nor UO_464 (O_464,N_9871,N_9549);
nor UO_465 (O_465,N_9894,N_9993);
nand UO_466 (O_466,N_9560,N_9939);
xnor UO_467 (O_467,N_9750,N_9936);
nand UO_468 (O_468,N_9926,N_9593);
or UO_469 (O_469,N_9629,N_9673);
or UO_470 (O_470,N_9905,N_9677);
nor UO_471 (O_471,N_9964,N_9997);
or UO_472 (O_472,N_9529,N_9556);
and UO_473 (O_473,N_9781,N_9674);
and UO_474 (O_474,N_9580,N_9695);
or UO_475 (O_475,N_9902,N_9900);
nand UO_476 (O_476,N_9652,N_9792);
or UO_477 (O_477,N_9870,N_9786);
nor UO_478 (O_478,N_9898,N_9500);
and UO_479 (O_479,N_9720,N_9636);
nand UO_480 (O_480,N_9724,N_9736);
nor UO_481 (O_481,N_9513,N_9789);
nand UO_482 (O_482,N_9810,N_9904);
xor UO_483 (O_483,N_9779,N_9696);
xnor UO_484 (O_484,N_9963,N_9550);
or UO_485 (O_485,N_9834,N_9806);
nor UO_486 (O_486,N_9548,N_9753);
nand UO_487 (O_487,N_9654,N_9638);
or UO_488 (O_488,N_9565,N_9943);
xor UO_489 (O_489,N_9719,N_9752);
or UO_490 (O_490,N_9935,N_9525);
nor UO_491 (O_491,N_9987,N_9902);
xnor UO_492 (O_492,N_9555,N_9887);
and UO_493 (O_493,N_9619,N_9781);
nand UO_494 (O_494,N_9717,N_9834);
or UO_495 (O_495,N_9873,N_9956);
xnor UO_496 (O_496,N_9921,N_9622);
or UO_497 (O_497,N_9592,N_9880);
or UO_498 (O_498,N_9849,N_9592);
xor UO_499 (O_499,N_9769,N_9714);
xor UO_500 (O_500,N_9707,N_9551);
nand UO_501 (O_501,N_9891,N_9523);
or UO_502 (O_502,N_9637,N_9624);
or UO_503 (O_503,N_9553,N_9588);
nor UO_504 (O_504,N_9568,N_9819);
nor UO_505 (O_505,N_9675,N_9738);
xnor UO_506 (O_506,N_9734,N_9918);
xor UO_507 (O_507,N_9573,N_9641);
nand UO_508 (O_508,N_9526,N_9646);
nand UO_509 (O_509,N_9701,N_9953);
or UO_510 (O_510,N_9520,N_9696);
and UO_511 (O_511,N_9863,N_9822);
xnor UO_512 (O_512,N_9642,N_9744);
or UO_513 (O_513,N_9564,N_9575);
or UO_514 (O_514,N_9860,N_9822);
xor UO_515 (O_515,N_9793,N_9584);
or UO_516 (O_516,N_9896,N_9682);
nor UO_517 (O_517,N_9512,N_9867);
or UO_518 (O_518,N_9693,N_9896);
nor UO_519 (O_519,N_9524,N_9989);
or UO_520 (O_520,N_9696,N_9925);
or UO_521 (O_521,N_9883,N_9591);
xor UO_522 (O_522,N_9899,N_9659);
or UO_523 (O_523,N_9563,N_9597);
xor UO_524 (O_524,N_9716,N_9574);
nand UO_525 (O_525,N_9715,N_9530);
xnor UO_526 (O_526,N_9725,N_9682);
nor UO_527 (O_527,N_9699,N_9649);
xnor UO_528 (O_528,N_9789,N_9687);
or UO_529 (O_529,N_9937,N_9764);
nand UO_530 (O_530,N_9999,N_9784);
nand UO_531 (O_531,N_9756,N_9857);
and UO_532 (O_532,N_9910,N_9540);
nand UO_533 (O_533,N_9794,N_9587);
or UO_534 (O_534,N_9667,N_9989);
nor UO_535 (O_535,N_9667,N_9522);
nand UO_536 (O_536,N_9584,N_9919);
nor UO_537 (O_537,N_9893,N_9807);
nand UO_538 (O_538,N_9660,N_9613);
or UO_539 (O_539,N_9639,N_9811);
or UO_540 (O_540,N_9793,N_9693);
nand UO_541 (O_541,N_9805,N_9724);
or UO_542 (O_542,N_9615,N_9970);
nand UO_543 (O_543,N_9830,N_9766);
nor UO_544 (O_544,N_9914,N_9822);
nor UO_545 (O_545,N_9619,N_9884);
nand UO_546 (O_546,N_9694,N_9502);
nand UO_547 (O_547,N_9889,N_9585);
nor UO_548 (O_548,N_9542,N_9563);
nor UO_549 (O_549,N_9950,N_9636);
nor UO_550 (O_550,N_9710,N_9550);
nand UO_551 (O_551,N_9752,N_9821);
nor UO_552 (O_552,N_9898,N_9929);
nand UO_553 (O_553,N_9958,N_9535);
xor UO_554 (O_554,N_9664,N_9981);
or UO_555 (O_555,N_9965,N_9896);
or UO_556 (O_556,N_9625,N_9541);
nor UO_557 (O_557,N_9607,N_9681);
and UO_558 (O_558,N_9837,N_9729);
nand UO_559 (O_559,N_9547,N_9570);
nor UO_560 (O_560,N_9600,N_9847);
xor UO_561 (O_561,N_9614,N_9919);
nand UO_562 (O_562,N_9888,N_9641);
xnor UO_563 (O_563,N_9574,N_9794);
nand UO_564 (O_564,N_9978,N_9836);
and UO_565 (O_565,N_9812,N_9667);
xor UO_566 (O_566,N_9944,N_9670);
nor UO_567 (O_567,N_9855,N_9922);
nor UO_568 (O_568,N_9882,N_9869);
and UO_569 (O_569,N_9731,N_9656);
and UO_570 (O_570,N_9727,N_9649);
or UO_571 (O_571,N_9926,N_9537);
xor UO_572 (O_572,N_9602,N_9948);
xor UO_573 (O_573,N_9570,N_9624);
or UO_574 (O_574,N_9947,N_9889);
nor UO_575 (O_575,N_9955,N_9530);
nor UO_576 (O_576,N_9661,N_9812);
nand UO_577 (O_577,N_9976,N_9860);
nand UO_578 (O_578,N_9953,N_9706);
nand UO_579 (O_579,N_9978,N_9725);
or UO_580 (O_580,N_9619,N_9905);
and UO_581 (O_581,N_9860,N_9768);
nor UO_582 (O_582,N_9744,N_9623);
nor UO_583 (O_583,N_9801,N_9973);
and UO_584 (O_584,N_9704,N_9861);
nand UO_585 (O_585,N_9700,N_9594);
nor UO_586 (O_586,N_9897,N_9512);
and UO_587 (O_587,N_9980,N_9988);
nor UO_588 (O_588,N_9501,N_9735);
nand UO_589 (O_589,N_9866,N_9787);
or UO_590 (O_590,N_9784,N_9846);
xnor UO_591 (O_591,N_9724,N_9978);
xor UO_592 (O_592,N_9807,N_9879);
and UO_593 (O_593,N_9662,N_9899);
nor UO_594 (O_594,N_9527,N_9717);
and UO_595 (O_595,N_9699,N_9998);
nor UO_596 (O_596,N_9728,N_9660);
nand UO_597 (O_597,N_9638,N_9750);
or UO_598 (O_598,N_9746,N_9994);
or UO_599 (O_599,N_9752,N_9745);
and UO_600 (O_600,N_9519,N_9619);
xnor UO_601 (O_601,N_9953,N_9606);
xor UO_602 (O_602,N_9848,N_9841);
or UO_603 (O_603,N_9914,N_9550);
or UO_604 (O_604,N_9872,N_9550);
or UO_605 (O_605,N_9514,N_9702);
or UO_606 (O_606,N_9635,N_9604);
nand UO_607 (O_607,N_9600,N_9721);
nand UO_608 (O_608,N_9984,N_9665);
nand UO_609 (O_609,N_9621,N_9866);
and UO_610 (O_610,N_9558,N_9877);
xnor UO_611 (O_611,N_9654,N_9692);
nor UO_612 (O_612,N_9522,N_9981);
xnor UO_613 (O_613,N_9502,N_9934);
and UO_614 (O_614,N_9716,N_9845);
nand UO_615 (O_615,N_9937,N_9888);
and UO_616 (O_616,N_9534,N_9793);
nand UO_617 (O_617,N_9710,N_9993);
or UO_618 (O_618,N_9735,N_9907);
and UO_619 (O_619,N_9599,N_9559);
and UO_620 (O_620,N_9967,N_9684);
xnor UO_621 (O_621,N_9856,N_9570);
nor UO_622 (O_622,N_9867,N_9892);
nor UO_623 (O_623,N_9942,N_9951);
or UO_624 (O_624,N_9639,N_9967);
and UO_625 (O_625,N_9838,N_9829);
or UO_626 (O_626,N_9729,N_9717);
nand UO_627 (O_627,N_9959,N_9827);
nor UO_628 (O_628,N_9835,N_9544);
nor UO_629 (O_629,N_9927,N_9813);
nand UO_630 (O_630,N_9976,N_9682);
nor UO_631 (O_631,N_9633,N_9604);
or UO_632 (O_632,N_9895,N_9707);
nor UO_633 (O_633,N_9557,N_9939);
xor UO_634 (O_634,N_9720,N_9807);
and UO_635 (O_635,N_9902,N_9744);
nor UO_636 (O_636,N_9770,N_9876);
nand UO_637 (O_637,N_9857,N_9769);
nand UO_638 (O_638,N_9529,N_9566);
and UO_639 (O_639,N_9513,N_9794);
or UO_640 (O_640,N_9959,N_9651);
or UO_641 (O_641,N_9991,N_9953);
nand UO_642 (O_642,N_9850,N_9723);
or UO_643 (O_643,N_9818,N_9808);
nor UO_644 (O_644,N_9982,N_9781);
nand UO_645 (O_645,N_9552,N_9809);
or UO_646 (O_646,N_9892,N_9716);
nor UO_647 (O_647,N_9954,N_9792);
nand UO_648 (O_648,N_9652,N_9771);
and UO_649 (O_649,N_9998,N_9649);
nand UO_650 (O_650,N_9893,N_9563);
nand UO_651 (O_651,N_9507,N_9869);
nand UO_652 (O_652,N_9773,N_9992);
xor UO_653 (O_653,N_9936,N_9577);
nand UO_654 (O_654,N_9817,N_9760);
nor UO_655 (O_655,N_9928,N_9725);
and UO_656 (O_656,N_9904,N_9717);
nor UO_657 (O_657,N_9924,N_9638);
and UO_658 (O_658,N_9529,N_9856);
nor UO_659 (O_659,N_9797,N_9812);
xor UO_660 (O_660,N_9862,N_9789);
nor UO_661 (O_661,N_9930,N_9789);
and UO_662 (O_662,N_9877,N_9532);
and UO_663 (O_663,N_9903,N_9631);
or UO_664 (O_664,N_9517,N_9948);
nor UO_665 (O_665,N_9577,N_9946);
xor UO_666 (O_666,N_9890,N_9983);
and UO_667 (O_667,N_9963,N_9881);
or UO_668 (O_668,N_9957,N_9707);
nor UO_669 (O_669,N_9574,N_9877);
and UO_670 (O_670,N_9823,N_9688);
xor UO_671 (O_671,N_9870,N_9896);
xnor UO_672 (O_672,N_9523,N_9684);
nand UO_673 (O_673,N_9829,N_9566);
nand UO_674 (O_674,N_9751,N_9564);
and UO_675 (O_675,N_9627,N_9651);
nand UO_676 (O_676,N_9968,N_9715);
or UO_677 (O_677,N_9522,N_9929);
or UO_678 (O_678,N_9928,N_9622);
and UO_679 (O_679,N_9653,N_9687);
nand UO_680 (O_680,N_9956,N_9947);
xor UO_681 (O_681,N_9586,N_9536);
and UO_682 (O_682,N_9875,N_9872);
and UO_683 (O_683,N_9879,N_9805);
and UO_684 (O_684,N_9744,N_9503);
nand UO_685 (O_685,N_9961,N_9870);
or UO_686 (O_686,N_9868,N_9596);
nand UO_687 (O_687,N_9986,N_9736);
or UO_688 (O_688,N_9748,N_9536);
xor UO_689 (O_689,N_9978,N_9645);
xnor UO_690 (O_690,N_9742,N_9935);
and UO_691 (O_691,N_9719,N_9628);
and UO_692 (O_692,N_9693,N_9893);
or UO_693 (O_693,N_9769,N_9716);
nor UO_694 (O_694,N_9850,N_9632);
nor UO_695 (O_695,N_9740,N_9968);
nand UO_696 (O_696,N_9951,N_9741);
nand UO_697 (O_697,N_9617,N_9739);
nand UO_698 (O_698,N_9862,N_9706);
nand UO_699 (O_699,N_9883,N_9513);
or UO_700 (O_700,N_9644,N_9602);
nor UO_701 (O_701,N_9880,N_9792);
nor UO_702 (O_702,N_9860,N_9727);
nand UO_703 (O_703,N_9872,N_9992);
nor UO_704 (O_704,N_9728,N_9978);
nor UO_705 (O_705,N_9978,N_9713);
and UO_706 (O_706,N_9616,N_9679);
nor UO_707 (O_707,N_9696,N_9644);
or UO_708 (O_708,N_9838,N_9744);
nor UO_709 (O_709,N_9814,N_9798);
and UO_710 (O_710,N_9646,N_9584);
and UO_711 (O_711,N_9554,N_9837);
and UO_712 (O_712,N_9789,N_9571);
nor UO_713 (O_713,N_9789,N_9902);
or UO_714 (O_714,N_9814,N_9823);
nand UO_715 (O_715,N_9844,N_9812);
or UO_716 (O_716,N_9958,N_9515);
and UO_717 (O_717,N_9544,N_9637);
nor UO_718 (O_718,N_9869,N_9906);
xnor UO_719 (O_719,N_9733,N_9853);
xnor UO_720 (O_720,N_9741,N_9878);
xor UO_721 (O_721,N_9657,N_9945);
nand UO_722 (O_722,N_9778,N_9659);
and UO_723 (O_723,N_9564,N_9740);
nand UO_724 (O_724,N_9927,N_9824);
nor UO_725 (O_725,N_9756,N_9662);
nor UO_726 (O_726,N_9887,N_9530);
xnor UO_727 (O_727,N_9662,N_9704);
xor UO_728 (O_728,N_9688,N_9942);
and UO_729 (O_729,N_9789,N_9593);
nand UO_730 (O_730,N_9671,N_9581);
and UO_731 (O_731,N_9561,N_9749);
and UO_732 (O_732,N_9579,N_9736);
or UO_733 (O_733,N_9855,N_9933);
nand UO_734 (O_734,N_9604,N_9957);
nor UO_735 (O_735,N_9652,N_9902);
nor UO_736 (O_736,N_9687,N_9933);
nand UO_737 (O_737,N_9988,N_9544);
xnor UO_738 (O_738,N_9889,N_9738);
and UO_739 (O_739,N_9529,N_9786);
nor UO_740 (O_740,N_9588,N_9988);
nand UO_741 (O_741,N_9890,N_9871);
xor UO_742 (O_742,N_9677,N_9904);
or UO_743 (O_743,N_9620,N_9919);
xor UO_744 (O_744,N_9828,N_9853);
or UO_745 (O_745,N_9768,N_9780);
xnor UO_746 (O_746,N_9945,N_9899);
or UO_747 (O_747,N_9867,N_9903);
xor UO_748 (O_748,N_9515,N_9686);
xor UO_749 (O_749,N_9946,N_9752);
and UO_750 (O_750,N_9763,N_9858);
nand UO_751 (O_751,N_9583,N_9955);
or UO_752 (O_752,N_9666,N_9531);
xnor UO_753 (O_753,N_9749,N_9918);
xnor UO_754 (O_754,N_9892,N_9694);
and UO_755 (O_755,N_9627,N_9670);
xor UO_756 (O_756,N_9513,N_9615);
nand UO_757 (O_757,N_9912,N_9996);
xor UO_758 (O_758,N_9574,N_9568);
xor UO_759 (O_759,N_9766,N_9802);
or UO_760 (O_760,N_9953,N_9859);
nand UO_761 (O_761,N_9699,N_9755);
xor UO_762 (O_762,N_9975,N_9518);
and UO_763 (O_763,N_9663,N_9529);
and UO_764 (O_764,N_9708,N_9626);
or UO_765 (O_765,N_9940,N_9696);
nand UO_766 (O_766,N_9955,N_9966);
and UO_767 (O_767,N_9569,N_9986);
or UO_768 (O_768,N_9899,N_9767);
nor UO_769 (O_769,N_9723,N_9907);
xnor UO_770 (O_770,N_9946,N_9828);
or UO_771 (O_771,N_9656,N_9672);
nand UO_772 (O_772,N_9652,N_9844);
xor UO_773 (O_773,N_9668,N_9878);
xnor UO_774 (O_774,N_9841,N_9844);
and UO_775 (O_775,N_9500,N_9982);
or UO_776 (O_776,N_9523,N_9762);
nand UO_777 (O_777,N_9514,N_9652);
nand UO_778 (O_778,N_9726,N_9812);
or UO_779 (O_779,N_9861,N_9912);
nand UO_780 (O_780,N_9781,N_9949);
nand UO_781 (O_781,N_9772,N_9792);
or UO_782 (O_782,N_9659,N_9565);
xor UO_783 (O_783,N_9520,N_9868);
or UO_784 (O_784,N_9917,N_9559);
nand UO_785 (O_785,N_9840,N_9857);
nor UO_786 (O_786,N_9865,N_9658);
or UO_787 (O_787,N_9646,N_9842);
xor UO_788 (O_788,N_9587,N_9736);
nand UO_789 (O_789,N_9827,N_9993);
xor UO_790 (O_790,N_9857,N_9624);
nor UO_791 (O_791,N_9821,N_9540);
or UO_792 (O_792,N_9976,N_9915);
or UO_793 (O_793,N_9642,N_9697);
or UO_794 (O_794,N_9930,N_9810);
and UO_795 (O_795,N_9679,N_9694);
xnor UO_796 (O_796,N_9934,N_9690);
and UO_797 (O_797,N_9815,N_9709);
or UO_798 (O_798,N_9710,N_9644);
and UO_799 (O_799,N_9829,N_9966);
xor UO_800 (O_800,N_9956,N_9908);
nand UO_801 (O_801,N_9985,N_9572);
nand UO_802 (O_802,N_9943,N_9684);
xnor UO_803 (O_803,N_9678,N_9645);
xnor UO_804 (O_804,N_9993,N_9695);
xor UO_805 (O_805,N_9698,N_9730);
nor UO_806 (O_806,N_9832,N_9514);
nand UO_807 (O_807,N_9683,N_9618);
or UO_808 (O_808,N_9673,N_9894);
and UO_809 (O_809,N_9632,N_9582);
nand UO_810 (O_810,N_9855,N_9852);
or UO_811 (O_811,N_9590,N_9520);
nand UO_812 (O_812,N_9590,N_9939);
xnor UO_813 (O_813,N_9656,N_9671);
and UO_814 (O_814,N_9957,N_9998);
nor UO_815 (O_815,N_9576,N_9590);
nor UO_816 (O_816,N_9709,N_9842);
xor UO_817 (O_817,N_9955,N_9915);
nand UO_818 (O_818,N_9896,N_9519);
or UO_819 (O_819,N_9757,N_9706);
and UO_820 (O_820,N_9941,N_9928);
and UO_821 (O_821,N_9532,N_9875);
or UO_822 (O_822,N_9575,N_9841);
and UO_823 (O_823,N_9749,N_9877);
or UO_824 (O_824,N_9742,N_9819);
nor UO_825 (O_825,N_9597,N_9649);
nor UO_826 (O_826,N_9731,N_9673);
nor UO_827 (O_827,N_9944,N_9841);
or UO_828 (O_828,N_9962,N_9514);
or UO_829 (O_829,N_9771,N_9911);
nor UO_830 (O_830,N_9850,N_9867);
nand UO_831 (O_831,N_9939,N_9526);
xor UO_832 (O_832,N_9816,N_9844);
or UO_833 (O_833,N_9735,N_9920);
or UO_834 (O_834,N_9531,N_9942);
nand UO_835 (O_835,N_9631,N_9960);
and UO_836 (O_836,N_9819,N_9703);
or UO_837 (O_837,N_9813,N_9585);
xor UO_838 (O_838,N_9515,N_9824);
nor UO_839 (O_839,N_9795,N_9631);
or UO_840 (O_840,N_9615,N_9862);
or UO_841 (O_841,N_9849,N_9907);
xnor UO_842 (O_842,N_9779,N_9849);
or UO_843 (O_843,N_9551,N_9809);
xor UO_844 (O_844,N_9797,N_9902);
nand UO_845 (O_845,N_9779,N_9990);
or UO_846 (O_846,N_9697,N_9960);
or UO_847 (O_847,N_9571,N_9788);
nor UO_848 (O_848,N_9810,N_9658);
nor UO_849 (O_849,N_9633,N_9729);
nand UO_850 (O_850,N_9888,N_9677);
or UO_851 (O_851,N_9651,N_9649);
nand UO_852 (O_852,N_9764,N_9994);
nor UO_853 (O_853,N_9901,N_9527);
nand UO_854 (O_854,N_9502,N_9941);
and UO_855 (O_855,N_9569,N_9900);
nor UO_856 (O_856,N_9797,N_9867);
and UO_857 (O_857,N_9800,N_9559);
nand UO_858 (O_858,N_9606,N_9672);
xor UO_859 (O_859,N_9747,N_9947);
nor UO_860 (O_860,N_9863,N_9795);
nand UO_861 (O_861,N_9806,N_9707);
xnor UO_862 (O_862,N_9740,N_9605);
nand UO_863 (O_863,N_9711,N_9881);
nor UO_864 (O_864,N_9508,N_9655);
nor UO_865 (O_865,N_9964,N_9660);
or UO_866 (O_866,N_9530,N_9941);
nand UO_867 (O_867,N_9678,N_9697);
nor UO_868 (O_868,N_9756,N_9621);
or UO_869 (O_869,N_9755,N_9716);
or UO_870 (O_870,N_9699,N_9987);
xor UO_871 (O_871,N_9691,N_9582);
or UO_872 (O_872,N_9603,N_9830);
and UO_873 (O_873,N_9687,N_9889);
nor UO_874 (O_874,N_9757,N_9707);
and UO_875 (O_875,N_9770,N_9836);
xnor UO_876 (O_876,N_9622,N_9893);
and UO_877 (O_877,N_9679,N_9806);
or UO_878 (O_878,N_9595,N_9541);
xnor UO_879 (O_879,N_9857,N_9972);
xnor UO_880 (O_880,N_9751,N_9531);
nand UO_881 (O_881,N_9701,N_9809);
nor UO_882 (O_882,N_9925,N_9679);
xor UO_883 (O_883,N_9675,N_9644);
nor UO_884 (O_884,N_9662,N_9631);
nand UO_885 (O_885,N_9813,N_9746);
or UO_886 (O_886,N_9801,N_9605);
nor UO_887 (O_887,N_9572,N_9514);
or UO_888 (O_888,N_9948,N_9657);
and UO_889 (O_889,N_9601,N_9888);
or UO_890 (O_890,N_9824,N_9651);
xnor UO_891 (O_891,N_9598,N_9919);
nand UO_892 (O_892,N_9621,N_9840);
xnor UO_893 (O_893,N_9620,N_9873);
and UO_894 (O_894,N_9700,N_9907);
and UO_895 (O_895,N_9898,N_9518);
nor UO_896 (O_896,N_9981,N_9571);
and UO_897 (O_897,N_9693,N_9923);
xnor UO_898 (O_898,N_9658,N_9587);
nand UO_899 (O_899,N_9587,N_9744);
nor UO_900 (O_900,N_9742,N_9890);
nand UO_901 (O_901,N_9522,N_9542);
nand UO_902 (O_902,N_9749,N_9652);
nor UO_903 (O_903,N_9718,N_9540);
and UO_904 (O_904,N_9626,N_9674);
nand UO_905 (O_905,N_9902,N_9704);
or UO_906 (O_906,N_9781,N_9948);
and UO_907 (O_907,N_9656,N_9824);
nand UO_908 (O_908,N_9976,N_9985);
xnor UO_909 (O_909,N_9844,N_9543);
or UO_910 (O_910,N_9661,N_9851);
and UO_911 (O_911,N_9958,N_9982);
xor UO_912 (O_912,N_9901,N_9872);
and UO_913 (O_913,N_9619,N_9651);
nand UO_914 (O_914,N_9717,N_9616);
xor UO_915 (O_915,N_9994,N_9818);
and UO_916 (O_916,N_9716,N_9645);
or UO_917 (O_917,N_9543,N_9582);
xnor UO_918 (O_918,N_9943,N_9698);
nor UO_919 (O_919,N_9787,N_9575);
xor UO_920 (O_920,N_9535,N_9934);
nand UO_921 (O_921,N_9796,N_9845);
nand UO_922 (O_922,N_9982,N_9689);
and UO_923 (O_923,N_9644,N_9896);
xnor UO_924 (O_924,N_9625,N_9888);
and UO_925 (O_925,N_9832,N_9664);
or UO_926 (O_926,N_9606,N_9539);
or UO_927 (O_927,N_9681,N_9811);
nor UO_928 (O_928,N_9944,N_9636);
nor UO_929 (O_929,N_9877,N_9850);
or UO_930 (O_930,N_9957,N_9835);
nand UO_931 (O_931,N_9784,N_9773);
or UO_932 (O_932,N_9766,N_9944);
or UO_933 (O_933,N_9903,N_9553);
xnor UO_934 (O_934,N_9813,N_9726);
nor UO_935 (O_935,N_9757,N_9510);
and UO_936 (O_936,N_9946,N_9874);
and UO_937 (O_937,N_9845,N_9602);
nand UO_938 (O_938,N_9982,N_9619);
or UO_939 (O_939,N_9802,N_9744);
nor UO_940 (O_940,N_9729,N_9955);
nand UO_941 (O_941,N_9638,N_9910);
nand UO_942 (O_942,N_9544,N_9851);
nand UO_943 (O_943,N_9839,N_9737);
xor UO_944 (O_944,N_9764,N_9693);
or UO_945 (O_945,N_9588,N_9930);
or UO_946 (O_946,N_9502,N_9801);
nand UO_947 (O_947,N_9912,N_9903);
xor UO_948 (O_948,N_9651,N_9566);
nand UO_949 (O_949,N_9733,N_9524);
xnor UO_950 (O_950,N_9642,N_9519);
xor UO_951 (O_951,N_9726,N_9751);
or UO_952 (O_952,N_9882,N_9778);
nor UO_953 (O_953,N_9523,N_9648);
nor UO_954 (O_954,N_9587,N_9694);
nor UO_955 (O_955,N_9833,N_9628);
nor UO_956 (O_956,N_9875,N_9845);
or UO_957 (O_957,N_9597,N_9830);
or UO_958 (O_958,N_9585,N_9791);
nand UO_959 (O_959,N_9549,N_9604);
or UO_960 (O_960,N_9537,N_9925);
nand UO_961 (O_961,N_9747,N_9963);
nand UO_962 (O_962,N_9558,N_9512);
nand UO_963 (O_963,N_9723,N_9766);
or UO_964 (O_964,N_9952,N_9520);
xnor UO_965 (O_965,N_9713,N_9546);
and UO_966 (O_966,N_9846,N_9935);
xor UO_967 (O_967,N_9778,N_9987);
and UO_968 (O_968,N_9659,N_9989);
and UO_969 (O_969,N_9670,N_9979);
and UO_970 (O_970,N_9685,N_9541);
nor UO_971 (O_971,N_9884,N_9513);
nor UO_972 (O_972,N_9625,N_9753);
or UO_973 (O_973,N_9991,N_9782);
and UO_974 (O_974,N_9840,N_9732);
xnor UO_975 (O_975,N_9902,N_9699);
nor UO_976 (O_976,N_9673,N_9912);
or UO_977 (O_977,N_9907,N_9514);
and UO_978 (O_978,N_9740,N_9950);
nor UO_979 (O_979,N_9742,N_9599);
nor UO_980 (O_980,N_9764,N_9569);
nand UO_981 (O_981,N_9717,N_9782);
xnor UO_982 (O_982,N_9981,N_9509);
xnor UO_983 (O_983,N_9511,N_9861);
nand UO_984 (O_984,N_9555,N_9504);
nand UO_985 (O_985,N_9728,N_9524);
nand UO_986 (O_986,N_9583,N_9672);
or UO_987 (O_987,N_9949,N_9722);
nor UO_988 (O_988,N_9771,N_9737);
and UO_989 (O_989,N_9775,N_9635);
nor UO_990 (O_990,N_9594,N_9633);
nand UO_991 (O_991,N_9881,N_9899);
and UO_992 (O_992,N_9935,N_9868);
nor UO_993 (O_993,N_9799,N_9980);
nand UO_994 (O_994,N_9516,N_9520);
or UO_995 (O_995,N_9586,N_9664);
nor UO_996 (O_996,N_9640,N_9922);
nor UO_997 (O_997,N_9856,N_9952);
and UO_998 (O_998,N_9620,N_9960);
nor UO_999 (O_999,N_9771,N_9720);
and UO_1000 (O_1000,N_9617,N_9652);
or UO_1001 (O_1001,N_9836,N_9918);
and UO_1002 (O_1002,N_9829,N_9856);
xnor UO_1003 (O_1003,N_9829,N_9590);
nor UO_1004 (O_1004,N_9721,N_9786);
and UO_1005 (O_1005,N_9829,N_9978);
or UO_1006 (O_1006,N_9830,N_9690);
and UO_1007 (O_1007,N_9922,N_9609);
and UO_1008 (O_1008,N_9777,N_9928);
nand UO_1009 (O_1009,N_9911,N_9870);
or UO_1010 (O_1010,N_9811,N_9674);
and UO_1011 (O_1011,N_9511,N_9828);
and UO_1012 (O_1012,N_9563,N_9792);
or UO_1013 (O_1013,N_9670,N_9744);
xnor UO_1014 (O_1014,N_9801,N_9924);
nor UO_1015 (O_1015,N_9773,N_9985);
or UO_1016 (O_1016,N_9952,N_9664);
nand UO_1017 (O_1017,N_9727,N_9623);
nand UO_1018 (O_1018,N_9620,N_9902);
nor UO_1019 (O_1019,N_9743,N_9949);
nand UO_1020 (O_1020,N_9717,N_9889);
or UO_1021 (O_1021,N_9848,N_9585);
xor UO_1022 (O_1022,N_9549,N_9767);
and UO_1023 (O_1023,N_9635,N_9876);
and UO_1024 (O_1024,N_9949,N_9542);
nand UO_1025 (O_1025,N_9591,N_9951);
nor UO_1026 (O_1026,N_9935,N_9877);
nor UO_1027 (O_1027,N_9733,N_9521);
nand UO_1028 (O_1028,N_9912,N_9676);
xnor UO_1029 (O_1029,N_9580,N_9991);
or UO_1030 (O_1030,N_9740,N_9637);
nand UO_1031 (O_1031,N_9942,N_9542);
xor UO_1032 (O_1032,N_9952,N_9702);
nor UO_1033 (O_1033,N_9730,N_9563);
or UO_1034 (O_1034,N_9733,N_9680);
nor UO_1035 (O_1035,N_9556,N_9615);
nand UO_1036 (O_1036,N_9985,N_9904);
xor UO_1037 (O_1037,N_9508,N_9728);
and UO_1038 (O_1038,N_9844,N_9885);
nor UO_1039 (O_1039,N_9703,N_9700);
and UO_1040 (O_1040,N_9939,N_9794);
nor UO_1041 (O_1041,N_9964,N_9541);
xnor UO_1042 (O_1042,N_9546,N_9932);
nand UO_1043 (O_1043,N_9626,N_9638);
nand UO_1044 (O_1044,N_9962,N_9833);
or UO_1045 (O_1045,N_9534,N_9595);
and UO_1046 (O_1046,N_9713,N_9758);
nand UO_1047 (O_1047,N_9626,N_9701);
nand UO_1048 (O_1048,N_9821,N_9958);
xor UO_1049 (O_1049,N_9801,N_9763);
xnor UO_1050 (O_1050,N_9945,N_9519);
xor UO_1051 (O_1051,N_9620,N_9599);
and UO_1052 (O_1052,N_9966,N_9961);
or UO_1053 (O_1053,N_9964,N_9973);
xor UO_1054 (O_1054,N_9699,N_9663);
nand UO_1055 (O_1055,N_9522,N_9836);
xor UO_1056 (O_1056,N_9724,N_9686);
xnor UO_1057 (O_1057,N_9588,N_9938);
nand UO_1058 (O_1058,N_9728,N_9918);
and UO_1059 (O_1059,N_9876,N_9846);
nand UO_1060 (O_1060,N_9783,N_9960);
xor UO_1061 (O_1061,N_9596,N_9783);
or UO_1062 (O_1062,N_9856,N_9783);
nand UO_1063 (O_1063,N_9936,N_9982);
xor UO_1064 (O_1064,N_9577,N_9757);
or UO_1065 (O_1065,N_9504,N_9507);
and UO_1066 (O_1066,N_9981,N_9784);
and UO_1067 (O_1067,N_9805,N_9727);
xor UO_1068 (O_1068,N_9890,N_9633);
nand UO_1069 (O_1069,N_9561,N_9639);
and UO_1070 (O_1070,N_9532,N_9900);
and UO_1071 (O_1071,N_9598,N_9846);
xnor UO_1072 (O_1072,N_9900,N_9822);
or UO_1073 (O_1073,N_9947,N_9972);
and UO_1074 (O_1074,N_9799,N_9674);
and UO_1075 (O_1075,N_9795,N_9737);
or UO_1076 (O_1076,N_9712,N_9691);
xnor UO_1077 (O_1077,N_9761,N_9617);
and UO_1078 (O_1078,N_9570,N_9666);
xnor UO_1079 (O_1079,N_9545,N_9585);
or UO_1080 (O_1080,N_9972,N_9648);
and UO_1081 (O_1081,N_9848,N_9699);
nor UO_1082 (O_1082,N_9667,N_9844);
or UO_1083 (O_1083,N_9802,N_9552);
or UO_1084 (O_1084,N_9925,N_9937);
and UO_1085 (O_1085,N_9932,N_9680);
and UO_1086 (O_1086,N_9970,N_9576);
nor UO_1087 (O_1087,N_9727,N_9903);
xor UO_1088 (O_1088,N_9545,N_9563);
and UO_1089 (O_1089,N_9719,N_9762);
and UO_1090 (O_1090,N_9858,N_9578);
or UO_1091 (O_1091,N_9821,N_9648);
or UO_1092 (O_1092,N_9753,N_9513);
nand UO_1093 (O_1093,N_9605,N_9585);
or UO_1094 (O_1094,N_9789,N_9682);
or UO_1095 (O_1095,N_9664,N_9916);
or UO_1096 (O_1096,N_9769,N_9768);
or UO_1097 (O_1097,N_9792,N_9952);
or UO_1098 (O_1098,N_9688,N_9993);
nor UO_1099 (O_1099,N_9506,N_9657);
and UO_1100 (O_1100,N_9609,N_9631);
xnor UO_1101 (O_1101,N_9970,N_9626);
nor UO_1102 (O_1102,N_9700,N_9748);
or UO_1103 (O_1103,N_9656,N_9995);
nor UO_1104 (O_1104,N_9676,N_9722);
and UO_1105 (O_1105,N_9788,N_9987);
xnor UO_1106 (O_1106,N_9522,N_9529);
and UO_1107 (O_1107,N_9750,N_9757);
xor UO_1108 (O_1108,N_9958,N_9579);
and UO_1109 (O_1109,N_9562,N_9946);
nor UO_1110 (O_1110,N_9837,N_9826);
xnor UO_1111 (O_1111,N_9879,N_9815);
and UO_1112 (O_1112,N_9540,N_9929);
nand UO_1113 (O_1113,N_9706,N_9792);
xnor UO_1114 (O_1114,N_9905,N_9843);
nor UO_1115 (O_1115,N_9965,N_9793);
nor UO_1116 (O_1116,N_9574,N_9802);
and UO_1117 (O_1117,N_9803,N_9714);
or UO_1118 (O_1118,N_9860,N_9783);
xor UO_1119 (O_1119,N_9988,N_9576);
and UO_1120 (O_1120,N_9665,N_9666);
nand UO_1121 (O_1121,N_9867,N_9535);
nor UO_1122 (O_1122,N_9581,N_9632);
nor UO_1123 (O_1123,N_9896,N_9916);
nor UO_1124 (O_1124,N_9776,N_9981);
xnor UO_1125 (O_1125,N_9547,N_9720);
nand UO_1126 (O_1126,N_9886,N_9717);
and UO_1127 (O_1127,N_9872,N_9701);
and UO_1128 (O_1128,N_9794,N_9657);
or UO_1129 (O_1129,N_9994,N_9748);
and UO_1130 (O_1130,N_9637,N_9920);
and UO_1131 (O_1131,N_9941,N_9715);
or UO_1132 (O_1132,N_9740,N_9833);
or UO_1133 (O_1133,N_9760,N_9860);
nor UO_1134 (O_1134,N_9523,N_9799);
and UO_1135 (O_1135,N_9825,N_9670);
and UO_1136 (O_1136,N_9827,N_9775);
or UO_1137 (O_1137,N_9560,N_9626);
and UO_1138 (O_1138,N_9772,N_9718);
xnor UO_1139 (O_1139,N_9505,N_9583);
nor UO_1140 (O_1140,N_9967,N_9531);
xnor UO_1141 (O_1141,N_9735,N_9755);
nor UO_1142 (O_1142,N_9573,N_9823);
xnor UO_1143 (O_1143,N_9964,N_9673);
nor UO_1144 (O_1144,N_9873,N_9852);
nor UO_1145 (O_1145,N_9736,N_9576);
nand UO_1146 (O_1146,N_9513,N_9972);
nor UO_1147 (O_1147,N_9512,N_9800);
xnor UO_1148 (O_1148,N_9816,N_9811);
nand UO_1149 (O_1149,N_9597,N_9617);
nand UO_1150 (O_1150,N_9528,N_9765);
nor UO_1151 (O_1151,N_9970,N_9919);
nand UO_1152 (O_1152,N_9874,N_9899);
and UO_1153 (O_1153,N_9874,N_9937);
or UO_1154 (O_1154,N_9963,N_9794);
nor UO_1155 (O_1155,N_9963,N_9875);
xnor UO_1156 (O_1156,N_9509,N_9719);
nand UO_1157 (O_1157,N_9810,N_9743);
nand UO_1158 (O_1158,N_9853,N_9623);
nand UO_1159 (O_1159,N_9945,N_9806);
or UO_1160 (O_1160,N_9707,N_9642);
nor UO_1161 (O_1161,N_9584,N_9836);
and UO_1162 (O_1162,N_9890,N_9779);
nor UO_1163 (O_1163,N_9685,N_9895);
nand UO_1164 (O_1164,N_9827,N_9931);
xnor UO_1165 (O_1165,N_9904,N_9819);
or UO_1166 (O_1166,N_9831,N_9616);
nand UO_1167 (O_1167,N_9577,N_9939);
xnor UO_1168 (O_1168,N_9693,N_9584);
nand UO_1169 (O_1169,N_9601,N_9887);
nor UO_1170 (O_1170,N_9777,N_9525);
xor UO_1171 (O_1171,N_9551,N_9702);
or UO_1172 (O_1172,N_9729,N_9802);
nor UO_1173 (O_1173,N_9967,N_9569);
nand UO_1174 (O_1174,N_9699,N_9563);
or UO_1175 (O_1175,N_9851,N_9758);
nand UO_1176 (O_1176,N_9806,N_9735);
xor UO_1177 (O_1177,N_9744,N_9637);
nand UO_1178 (O_1178,N_9988,N_9600);
or UO_1179 (O_1179,N_9536,N_9541);
nand UO_1180 (O_1180,N_9835,N_9713);
nor UO_1181 (O_1181,N_9547,N_9949);
nor UO_1182 (O_1182,N_9915,N_9673);
nand UO_1183 (O_1183,N_9879,N_9961);
and UO_1184 (O_1184,N_9623,N_9761);
nor UO_1185 (O_1185,N_9747,N_9697);
xnor UO_1186 (O_1186,N_9886,N_9819);
and UO_1187 (O_1187,N_9952,N_9588);
or UO_1188 (O_1188,N_9982,N_9819);
nor UO_1189 (O_1189,N_9994,N_9708);
xnor UO_1190 (O_1190,N_9547,N_9590);
xor UO_1191 (O_1191,N_9992,N_9534);
or UO_1192 (O_1192,N_9909,N_9857);
or UO_1193 (O_1193,N_9584,N_9891);
nand UO_1194 (O_1194,N_9783,N_9601);
or UO_1195 (O_1195,N_9632,N_9584);
and UO_1196 (O_1196,N_9987,N_9649);
nand UO_1197 (O_1197,N_9909,N_9935);
or UO_1198 (O_1198,N_9850,N_9823);
nand UO_1199 (O_1199,N_9824,N_9796);
xnor UO_1200 (O_1200,N_9554,N_9593);
nor UO_1201 (O_1201,N_9834,N_9697);
nand UO_1202 (O_1202,N_9601,N_9630);
or UO_1203 (O_1203,N_9536,N_9569);
xnor UO_1204 (O_1204,N_9538,N_9508);
and UO_1205 (O_1205,N_9951,N_9720);
or UO_1206 (O_1206,N_9990,N_9836);
nand UO_1207 (O_1207,N_9504,N_9982);
nor UO_1208 (O_1208,N_9541,N_9570);
xnor UO_1209 (O_1209,N_9554,N_9605);
and UO_1210 (O_1210,N_9537,N_9507);
or UO_1211 (O_1211,N_9616,N_9747);
and UO_1212 (O_1212,N_9694,N_9848);
or UO_1213 (O_1213,N_9610,N_9674);
and UO_1214 (O_1214,N_9782,N_9901);
or UO_1215 (O_1215,N_9742,N_9612);
nor UO_1216 (O_1216,N_9652,N_9731);
and UO_1217 (O_1217,N_9785,N_9592);
xnor UO_1218 (O_1218,N_9874,N_9542);
nand UO_1219 (O_1219,N_9713,N_9641);
nor UO_1220 (O_1220,N_9743,N_9513);
nor UO_1221 (O_1221,N_9780,N_9793);
nor UO_1222 (O_1222,N_9805,N_9617);
and UO_1223 (O_1223,N_9929,N_9967);
nand UO_1224 (O_1224,N_9867,N_9849);
xor UO_1225 (O_1225,N_9575,N_9989);
xnor UO_1226 (O_1226,N_9964,N_9664);
xnor UO_1227 (O_1227,N_9803,N_9767);
and UO_1228 (O_1228,N_9658,N_9560);
or UO_1229 (O_1229,N_9967,N_9617);
xnor UO_1230 (O_1230,N_9517,N_9742);
nand UO_1231 (O_1231,N_9913,N_9683);
nor UO_1232 (O_1232,N_9503,N_9957);
xor UO_1233 (O_1233,N_9591,N_9619);
nand UO_1234 (O_1234,N_9944,N_9847);
or UO_1235 (O_1235,N_9521,N_9959);
and UO_1236 (O_1236,N_9761,N_9923);
nor UO_1237 (O_1237,N_9904,N_9752);
nor UO_1238 (O_1238,N_9750,N_9843);
nand UO_1239 (O_1239,N_9912,N_9680);
nand UO_1240 (O_1240,N_9874,N_9835);
nand UO_1241 (O_1241,N_9987,N_9743);
xor UO_1242 (O_1242,N_9896,N_9723);
xnor UO_1243 (O_1243,N_9768,N_9579);
and UO_1244 (O_1244,N_9979,N_9592);
nand UO_1245 (O_1245,N_9534,N_9757);
nand UO_1246 (O_1246,N_9682,N_9737);
nand UO_1247 (O_1247,N_9891,N_9847);
and UO_1248 (O_1248,N_9780,N_9629);
nor UO_1249 (O_1249,N_9897,N_9502);
or UO_1250 (O_1250,N_9743,N_9765);
and UO_1251 (O_1251,N_9923,N_9756);
or UO_1252 (O_1252,N_9710,N_9906);
xnor UO_1253 (O_1253,N_9661,N_9523);
nand UO_1254 (O_1254,N_9976,N_9869);
or UO_1255 (O_1255,N_9803,N_9596);
xor UO_1256 (O_1256,N_9590,N_9885);
nor UO_1257 (O_1257,N_9649,N_9946);
nand UO_1258 (O_1258,N_9877,N_9611);
xnor UO_1259 (O_1259,N_9608,N_9856);
nand UO_1260 (O_1260,N_9815,N_9779);
and UO_1261 (O_1261,N_9639,N_9796);
nand UO_1262 (O_1262,N_9905,N_9536);
nor UO_1263 (O_1263,N_9784,N_9575);
xor UO_1264 (O_1264,N_9789,N_9927);
xnor UO_1265 (O_1265,N_9909,N_9847);
and UO_1266 (O_1266,N_9500,N_9557);
xnor UO_1267 (O_1267,N_9716,N_9994);
nor UO_1268 (O_1268,N_9635,N_9746);
and UO_1269 (O_1269,N_9630,N_9853);
and UO_1270 (O_1270,N_9996,N_9879);
xnor UO_1271 (O_1271,N_9723,N_9614);
xor UO_1272 (O_1272,N_9721,N_9655);
nor UO_1273 (O_1273,N_9928,N_9943);
nand UO_1274 (O_1274,N_9744,N_9727);
and UO_1275 (O_1275,N_9587,N_9950);
xnor UO_1276 (O_1276,N_9547,N_9858);
and UO_1277 (O_1277,N_9788,N_9899);
and UO_1278 (O_1278,N_9993,N_9911);
and UO_1279 (O_1279,N_9566,N_9549);
xnor UO_1280 (O_1280,N_9965,N_9930);
or UO_1281 (O_1281,N_9883,N_9553);
nor UO_1282 (O_1282,N_9904,N_9583);
nand UO_1283 (O_1283,N_9971,N_9981);
nor UO_1284 (O_1284,N_9622,N_9816);
xor UO_1285 (O_1285,N_9837,N_9708);
nand UO_1286 (O_1286,N_9681,N_9967);
or UO_1287 (O_1287,N_9958,N_9835);
xnor UO_1288 (O_1288,N_9674,N_9749);
nand UO_1289 (O_1289,N_9677,N_9824);
and UO_1290 (O_1290,N_9639,N_9744);
xnor UO_1291 (O_1291,N_9763,N_9892);
or UO_1292 (O_1292,N_9593,N_9677);
and UO_1293 (O_1293,N_9683,N_9647);
xor UO_1294 (O_1294,N_9805,N_9838);
or UO_1295 (O_1295,N_9799,N_9720);
or UO_1296 (O_1296,N_9660,N_9716);
or UO_1297 (O_1297,N_9726,N_9915);
or UO_1298 (O_1298,N_9912,N_9568);
and UO_1299 (O_1299,N_9678,N_9939);
or UO_1300 (O_1300,N_9866,N_9793);
xor UO_1301 (O_1301,N_9577,N_9765);
xnor UO_1302 (O_1302,N_9524,N_9991);
nand UO_1303 (O_1303,N_9979,N_9583);
and UO_1304 (O_1304,N_9737,N_9773);
nand UO_1305 (O_1305,N_9572,N_9605);
xnor UO_1306 (O_1306,N_9902,N_9512);
xor UO_1307 (O_1307,N_9832,N_9923);
xnor UO_1308 (O_1308,N_9734,N_9756);
nand UO_1309 (O_1309,N_9597,N_9883);
xnor UO_1310 (O_1310,N_9616,N_9680);
xor UO_1311 (O_1311,N_9742,N_9923);
and UO_1312 (O_1312,N_9571,N_9732);
and UO_1313 (O_1313,N_9519,N_9784);
and UO_1314 (O_1314,N_9807,N_9557);
and UO_1315 (O_1315,N_9924,N_9891);
nor UO_1316 (O_1316,N_9695,N_9709);
and UO_1317 (O_1317,N_9790,N_9670);
or UO_1318 (O_1318,N_9945,N_9601);
xnor UO_1319 (O_1319,N_9967,N_9784);
nor UO_1320 (O_1320,N_9537,N_9960);
nor UO_1321 (O_1321,N_9649,N_9623);
and UO_1322 (O_1322,N_9732,N_9925);
nor UO_1323 (O_1323,N_9757,N_9741);
nor UO_1324 (O_1324,N_9690,N_9649);
nor UO_1325 (O_1325,N_9827,N_9822);
nand UO_1326 (O_1326,N_9710,N_9697);
or UO_1327 (O_1327,N_9946,N_9515);
nand UO_1328 (O_1328,N_9621,N_9892);
nor UO_1329 (O_1329,N_9625,N_9950);
nand UO_1330 (O_1330,N_9980,N_9991);
and UO_1331 (O_1331,N_9667,N_9941);
nor UO_1332 (O_1332,N_9978,N_9753);
nor UO_1333 (O_1333,N_9667,N_9900);
nor UO_1334 (O_1334,N_9826,N_9593);
xnor UO_1335 (O_1335,N_9810,N_9803);
xor UO_1336 (O_1336,N_9668,N_9686);
or UO_1337 (O_1337,N_9554,N_9817);
or UO_1338 (O_1338,N_9934,N_9961);
nor UO_1339 (O_1339,N_9673,N_9569);
and UO_1340 (O_1340,N_9515,N_9684);
nor UO_1341 (O_1341,N_9910,N_9929);
and UO_1342 (O_1342,N_9840,N_9691);
and UO_1343 (O_1343,N_9723,N_9859);
nand UO_1344 (O_1344,N_9819,N_9972);
nand UO_1345 (O_1345,N_9702,N_9697);
nor UO_1346 (O_1346,N_9834,N_9835);
and UO_1347 (O_1347,N_9699,N_9507);
xnor UO_1348 (O_1348,N_9963,N_9570);
or UO_1349 (O_1349,N_9575,N_9806);
nor UO_1350 (O_1350,N_9614,N_9768);
and UO_1351 (O_1351,N_9706,N_9666);
nor UO_1352 (O_1352,N_9626,N_9953);
xnor UO_1353 (O_1353,N_9697,N_9555);
nand UO_1354 (O_1354,N_9636,N_9957);
and UO_1355 (O_1355,N_9649,N_9951);
nand UO_1356 (O_1356,N_9806,N_9730);
nand UO_1357 (O_1357,N_9967,N_9537);
nand UO_1358 (O_1358,N_9942,N_9870);
nand UO_1359 (O_1359,N_9663,N_9895);
xor UO_1360 (O_1360,N_9758,N_9998);
or UO_1361 (O_1361,N_9727,N_9752);
xor UO_1362 (O_1362,N_9703,N_9510);
nor UO_1363 (O_1363,N_9507,N_9827);
and UO_1364 (O_1364,N_9705,N_9862);
and UO_1365 (O_1365,N_9514,N_9724);
xor UO_1366 (O_1366,N_9992,N_9974);
xnor UO_1367 (O_1367,N_9566,N_9637);
or UO_1368 (O_1368,N_9793,N_9595);
and UO_1369 (O_1369,N_9647,N_9934);
nand UO_1370 (O_1370,N_9703,N_9970);
xnor UO_1371 (O_1371,N_9775,N_9634);
nand UO_1372 (O_1372,N_9664,N_9694);
nand UO_1373 (O_1373,N_9538,N_9983);
xnor UO_1374 (O_1374,N_9631,N_9933);
xnor UO_1375 (O_1375,N_9562,N_9743);
xnor UO_1376 (O_1376,N_9777,N_9646);
nand UO_1377 (O_1377,N_9701,N_9552);
xor UO_1378 (O_1378,N_9850,N_9576);
nand UO_1379 (O_1379,N_9872,N_9668);
and UO_1380 (O_1380,N_9762,N_9897);
nand UO_1381 (O_1381,N_9614,N_9900);
and UO_1382 (O_1382,N_9841,N_9909);
and UO_1383 (O_1383,N_9734,N_9617);
nand UO_1384 (O_1384,N_9907,N_9524);
nor UO_1385 (O_1385,N_9773,N_9840);
xor UO_1386 (O_1386,N_9691,N_9536);
nor UO_1387 (O_1387,N_9518,N_9658);
or UO_1388 (O_1388,N_9550,N_9858);
or UO_1389 (O_1389,N_9854,N_9609);
and UO_1390 (O_1390,N_9685,N_9728);
xor UO_1391 (O_1391,N_9537,N_9752);
xnor UO_1392 (O_1392,N_9720,N_9687);
and UO_1393 (O_1393,N_9891,N_9636);
and UO_1394 (O_1394,N_9521,N_9794);
nand UO_1395 (O_1395,N_9854,N_9820);
or UO_1396 (O_1396,N_9519,N_9988);
nor UO_1397 (O_1397,N_9897,N_9563);
nor UO_1398 (O_1398,N_9988,N_9524);
nand UO_1399 (O_1399,N_9731,N_9885);
and UO_1400 (O_1400,N_9706,N_9760);
xnor UO_1401 (O_1401,N_9999,N_9769);
and UO_1402 (O_1402,N_9729,N_9589);
nor UO_1403 (O_1403,N_9580,N_9519);
nor UO_1404 (O_1404,N_9997,N_9526);
xnor UO_1405 (O_1405,N_9636,N_9571);
and UO_1406 (O_1406,N_9705,N_9659);
and UO_1407 (O_1407,N_9971,N_9891);
nor UO_1408 (O_1408,N_9936,N_9843);
nor UO_1409 (O_1409,N_9526,N_9790);
xnor UO_1410 (O_1410,N_9567,N_9830);
xor UO_1411 (O_1411,N_9930,N_9969);
nand UO_1412 (O_1412,N_9564,N_9818);
xor UO_1413 (O_1413,N_9800,N_9726);
and UO_1414 (O_1414,N_9653,N_9918);
xor UO_1415 (O_1415,N_9827,N_9511);
nor UO_1416 (O_1416,N_9667,N_9596);
xor UO_1417 (O_1417,N_9553,N_9882);
or UO_1418 (O_1418,N_9516,N_9776);
xor UO_1419 (O_1419,N_9932,N_9919);
nor UO_1420 (O_1420,N_9702,N_9612);
nand UO_1421 (O_1421,N_9553,N_9916);
nand UO_1422 (O_1422,N_9793,N_9532);
nor UO_1423 (O_1423,N_9551,N_9587);
nand UO_1424 (O_1424,N_9548,N_9623);
nor UO_1425 (O_1425,N_9896,N_9761);
nor UO_1426 (O_1426,N_9698,N_9804);
nor UO_1427 (O_1427,N_9576,N_9723);
and UO_1428 (O_1428,N_9724,N_9541);
and UO_1429 (O_1429,N_9969,N_9537);
nand UO_1430 (O_1430,N_9722,N_9657);
nor UO_1431 (O_1431,N_9864,N_9534);
nand UO_1432 (O_1432,N_9555,N_9798);
nand UO_1433 (O_1433,N_9922,N_9626);
or UO_1434 (O_1434,N_9903,N_9620);
xnor UO_1435 (O_1435,N_9710,N_9640);
nor UO_1436 (O_1436,N_9575,N_9799);
xor UO_1437 (O_1437,N_9882,N_9634);
and UO_1438 (O_1438,N_9692,N_9993);
nand UO_1439 (O_1439,N_9621,N_9520);
nor UO_1440 (O_1440,N_9937,N_9738);
and UO_1441 (O_1441,N_9960,N_9654);
nor UO_1442 (O_1442,N_9646,N_9554);
or UO_1443 (O_1443,N_9594,N_9803);
or UO_1444 (O_1444,N_9749,N_9575);
and UO_1445 (O_1445,N_9713,N_9628);
nand UO_1446 (O_1446,N_9522,N_9976);
xnor UO_1447 (O_1447,N_9701,N_9660);
nor UO_1448 (O_1448,N_9695,N_9975);
and UO_1449 (O_1449,N_9805,N_9900);
or UO_1450 (O_1450,N_9721,N_9830);
nor UO_1451 (O_1451,N_9830,N_9702);
or UO_1452 (O_1452,N_9725,N_9616);
and UO_1453 (O_1453,N_9518,N_9873);
xnor UO_1454 (O_1454,N_9994,N_9887);
xnor UO_1455 (O_1455,N_9894,N_9574);
nor UO_1456 (O_1456,N_9704,N_9791);
xor UO_1457 (O_1457,N_9781,N_9714);
or UO_1458 (O_1458,N_9999,N_9704);
nor UO_1459 (O_1459,N_9502,N_9856);
xor UO_1460 (O_1460,N_9791,N_9575);
xor UO_1461 (O_1461,N_9772,N_9503);
nor UO_1462 (O_1462,N_9617,N_9797);
nor UO_1463 (O_1463,N_9968,N_9913);
and UO_1464 (O_1464,N_9979,N_9657);
nor UO_1465 (O_1465,N_9734,N_9546);
xor UO_1466 (O_1466,N_9606,N_9671);
and UO_1467 (O_1467,N_9583,N_9747);
and UO_1468 (O_1468,N_9755,N_9807);
nand UO_1469 (O_1469,N_9940,N_9532);
or UO_1470 (O_1470,N_9622,N_9789);
and UO_1471 (O_1471,N_9817,N_9586);
xor UO_1472 (O_1472,N_9780,N_9751);
xor UO_1473 (O_1473,N_9911,N_9763);
xnor UO_1474 (O_1474,N_9694,N_9603);
or UO_1475 (O_1475,N_9813,N_9551);
nor UO_1476 (O_1476,N_9790,N_9577);
nor UO_1477 (O_1477,N_9691,N_9898);
nand UO_1478 (O_1478,N_9706,N_9629);
or UO_1479 (O_1479,N_9505,N_9623);
xnor UO_1480 (O_1480,N_9639,N_9667);
nor UO_1481 (O_1481,N_9634,N_9611);
and UO_1482 (O_1482,N_9966,N_9849);
and UO_1483 (O_1483,N_9643,N_9670);
or UO_1484 (O_1484,N_9772,N_9911);
xor UO_1485 (O_1485,N_9602,N_9567);
nor UO_1486 (O_1486,N_9517,N_9868);
or UO_1487 (O_1487,N_9914,N_9865);
nor UO_1488 (O_1488,N_9774,N_9528);
nor UO_1489 (O_1489,N_9710,N_9684);
nor UO_1490 (O_1490,N_9709,N_9562);
and UO_1491 (O_1491,N_9520,N_9632);
xnor UO_1492 (O_1492,N_9594,N_9760);
nor UO_1493 (O_1493,N_9666,N_9688);
or UO_1494 (O_1494,N_9728,N_9529);
xnor UO_1495 (O_1495,N_9700,N_9825);
nand UO_1496 (O_1496,N_9706,N_9816);
and UO_1497 (O_1497,N_9796,N_9948);
xnor UO_1498 (O_1498,N_9673,N_9972);
nor UO_1499 (O_1499,N_9582,N_9850);
endmodule