module basic_2000_20000_2500_20_levels_5xor_9(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999;
and U0 (N_0,In_600,In_1389);
and U1 (N_1,In_1887,In_1307);
or U2 (N_2,In_747,In_239);
xor U3 (N_3,In_1405,In_275);
nand U4 (N_4,In_1404,In_1655);
or U5 (N_5,In_1211,In_436);
nand U6 (N_6,In_1316,In_463);
nor U7 (N_7,In_979,In_458);
and U8 (N_8,In_14,In_723);
nor U9 (N_9,In_1510,In_838);
and U10 (N_10,In_511,In_1977);
nor U11 (N_11,In_1203,In_1707);
nor U12 (N_12,In_1451,In_191);
or U13 (N_13,In_224,In_1525);
nor U14 (N_14,In_1346,In_934);
nor U15 (N_15,In_1670,In_1635);
nand U16 (N_16,In_1287,In_1966);
nand U17 (N_17,In_1234,In_1679);
or U18 (N_18,In_545,In_1607);
xor U19 (N_19,In_1879,In_1233);
nand U20 (N_20,In_1888,In_876);
or U21 (N_21,In_1675,In_356);
nand U22 (N_22,In_118,In_1458);
nor U23 (N_23,In_692,In_1380);
or U24 (N_24,In_1019,In_1944);
and U25 (N_25,In_990,In_1876);
nor U26 (N_26,In_485,In_1120);
nor U27 (N_27,In_1871,In_295);
nand U28 (N_28,In_1087,In_1377);
nand U29 (N_29,In_1927,In_397);
and U30 (N_30,In_999,In_314);
nand U31 (N_31,In_601,In_177);
nand U32 (N_32,In_1273,In_1671);
or U33 (N_33,In_968,In_1833);
xor U34 (N_34,In_1146,In_1547);
and U35 (N_35,In_1256,In_933);
and U36 (N_36,In_281,In_1371);
and U37 (N_37,In_1922,In_1835);
or U38 (N_38,In_716,In_1605);
and U39 (N_39,In_738,In_1765);
and U40 (N_40,In_976,In_1443);
or U41 (N_41,In_160,In_1329);
nand U42 (N_42,In_1946,In_1154);
or U43 (N_43,In_879,In_351);
or U44 (N_44,In_290,In_117);
and U45 (N_45,In_1691,In_613);
or U46 (N_46,In_749,In_928);
nand U47 (N_47,In_384,In_635);
and U48 (N_48,In_1299,In_64);
nor U49 (N_49,In_1207,In_516);
nand U50 (N_50,In_372,In_233);
or U51 (N_51,In_447,In_1272);
and U52 (N_52,In_645,In_273);
nand U53 (N_53,In_1209,In_236);
nor U54 (N_54,In_1846,In_1874);
nand U55 (N_55,In_444,In_88);
and U56 (N_56,In_452,In_854);
nor U57 (N_57,In_1568,In_1028);
nand U58 (N_58,In_1131,In_1258);
and U59 (N_59,In_1192,In_4);
and U60 (N_60,In_1231,In_559);
or U61 (N_61,In_1,In_1771);
xnor U62 (N_62,In_1176,In_1444);
and U63 (N_63,In_468,In_918);
xnor U64 (N_64,In_703,In_1369);
and U65 (N_65,In_1904,In_1000);
nand U66 (N_66,In_503,In_454);
and U67 (N_67,In_1390,In_1261);
nand U68 (N_68,In_693,In_375);
or U69 (N_69,In_1553,In_1683);
and U70 (N_70,In_1873,In_1005);
nor U71 (N_71,In_1807,In_1597);
and U72 (N_72,In_1375,In_1122);
nand U73 (N_73,In_1416,In_1644);
nand U74 (N_74,In_609,In_1106);
nor U75 (N_75,In_1539,In_665);
nand U76 (N_76,In_958,In_38);
and U77 (N_77,In_1354,In_1298);
xor U78 (N_78,In_1698,In_1750);
nand U79 (N_79,In_707,In_1464);
nand U80 (N_80,In_835,In_671);
nand U81 (N_81,In_1733,In_566);
and U82 (N_82,In_1358,In_882);
and U83 (N_83,In_1762,In_1251);
nor U84 (N_84,In_1190,In_970);
nor U85 (N_85,In_1226,In_223);
nand U86 (N_86,In_409,In_941);
nor U87 (N_87,In_333,In_1025);
nand U88 (N_88,In_1681,In_1945);
nor U89 (N_89,In_1002,In_1650);
xor U90 (N_90,In_674,In_914);
or U91 (N_91,In_1401,In_1399);
nand U92 (N_92,In_602,In_1485);
xnor U93 (N_93,In_610,In_346);
and U94 (N_94,In_1570,In_1129);
or U95 (N_95,In_629,In_1950);
and U96 (N_96,In_1069,In_1813);
or U97 (N_97,In_750,In_1712);
nand U98 (N_98,In_994,In_1971);
and U99 (N_99,In_1241,In_1801);
nor U100 (N_100,In_989,In_310);
nor U101 (N_101,In_1237,In_608);
xor U102 (N_102,In_448,In_369);
nor U103 (N_103,In_442,In_1281);
nor U104 (N_104,In_1023,In_949);
or U105 (N_105,In_1284,In_488);
or U106 (N_106,In_1891,In_97);
and U107 (N_107,In_798,In_376);
and U108 (N_108,In_595,In_1587);
or U109 (N_109,In_1892,In_975);
nand U110 (N_110,In_153,In_1688);
and U111 (N_111,In_709,In_418);
nand U112 (N_112,In_45,In_1531);
nor U113 (N_113,In_1572,In_1310);
or U114 (N_114,In_411,In_1214);
nor U115 (N_115,In_124,In_998);
or U116 (N_116,In_134,In_59);
nor U117 (N_117,In_825,In_558);
or U118 (N_118,In_1660,In_1324);
and U119 (N_119,In_966,In_1662);
xor U120 (N_120,In_54,In_345);
and U121 (N_121,In_209,In_410);
and U122 (N_122,In_1884,In_415);
xor U123 (N_123,In_1647,In_1734);
nand U124 (N_124,In_1546,In_1304);
or U125 (N_125,In_348,In_767);
nand U126 (N_126,In_758,In_75);
or U127 (N_127,In_1037,In_1054);
nor U128 (N_128,In_1109,In_626);
nor U129 (N_129,In_977,In_212);
or U130 (N_130,In_12,In_1268);
nand U131 (N_131,In_27,In_257);
nor U132 (N_132,In_89,In_725);
nor U133 (N_133,In_1743,In_752);
nand U134 (N_134,In_457,In_1333);
and U135 (N_135,In_1894,In_107);
or U136 (N_136,In_180,In_823);
and U137 (N_137,In_1787,In_1178);
xor U138 (N_138,In_1540,In_618);
or U139 (N_139,In_1078,In_1973);
xnor U140 (N_140,In_900,In_1244);
nand U141 (N_141,In_1817,In_445);
nor U142 (N_142,In_887,In_1756);
xor U143 (N_143,In_502,In_144);
nand U144 (N_144,In_620,In_695);
and U145 (N_145,In_1561,In_897);
nor U146 (N_146,In_1563,In_1667);
nor U147 (N_147,In_1582,In_9);
nand U148 (N_148,In_221,In_1076);
or U149 (N_149,In_715,In_1940);
nor U150 (N_150,In_687,In_1180);
or U151 (N_151,In_355,In_150);
or U152 (N_152,In_636,In_1355);
and U153 (N_153,In_759,In_782);
nor U154 (N_154,In_663,In_909);
xnor U155 (N_155,In_652,In_788);
or U156 (N_156,In_646,In_612);
nand U157 (N_157,In_1336,In_1665);
nor U158 (N_158,In_896,In_912);
nand U159 (N_159,In_913,In_1737);
and U160 (N_160,In_1452,In_1674);
or U161 (N_161,In_780,In_1278);
or U162 (N_162,In_805,In_541);
or U163 (N_163,In_1749,In_821);
or U164 (N_164,In_1642,In_1091);
xor U165 (N_165,In_971,In_1204);
and U166 (N_166,In_1632,In_1908);
xnor U167 (N_167,In_506,In_1867);
nor U168 (N_168,In_1174,In_1121);
or U169 (N_169,In_43,In_1661);
xnor U170 (N_170,In_342,In_1135);
nor U171 (N_171,In_517,In_1959);
nor U172 (N_172,In_653,In_74);
and U173 (N_173,In_801,In_563);
nor U174 (N_174,In_106,In_438);
and U175 (N_175,In_1323,In_1649);
xnor U176 (N_176,In_1780,In_531);
xor U177 (N_177,In_121,In_1300);
nand U178 (N_178,In_1242,In_812);
nor U179 (N_179,In_455,In_143);
nor U180 (N_180,In_381,In_1509);
nand U181 (N_181,In_1092,In_991);
and U182 (N_182,In_1589,In_1150);
and U183 (N_183,In_8,In_1104);
and U184 (N_184,In_1962,In_967);
nor U185 (N_185,In_858,In_1248);
nand U186 (N_186,In_1314,In_1694);
nand U187 (N_187,In_235,In_382);
or U188 (N_188,In_208,In_917);
nand U189 (N_189,In_1676,In_1555);
and U190 (N_190,In_312,In_286);
and U191 (N_191,In_1045,In_1627);
nor U192 (N_192,In_266,In_1013);
nand U193 (N_193,In_505,In_892);
nand U194 (N_194,In_514,In_885);
and U195 (N_195,In_1511,In_803);
xor U196 (N_196,In_466,In_510);
and U197 (N_197,In_165,In_625);
or U198 (N_198,In_1865,In_787);
xor U199 (N_199,In_568,In_83);
and U200 (N_200,In_1839,In_243);
and U201 (N_201,In_437,In_1090);
and U202 (N_202,In_274,In_1580);
nand U203 (N_203,In_403,In_1437);
or U204 (N_204,In_1987,In_560);
nor U205 (N_205,In_953,In_151);
nand U206 (N_206,In_1890,In_450);
xor U207 (N_207,In_432,In_34);
and U208 (N_208,In_1082,In_1229);
nand U209 (N_209,In_950,In_577);
or U210 (N_210,In_1040,In_816);
nor U211 (N_211,In_844,In_374);
and U212 (N_212,In_301,In_1758);
and U213 (N_213,In_576,In_1421);
and U214 (N_214,In_1680,In_1708);
nand U215 (N_215,In_26,In_1766);
and U216 (N_216,In_1249,In_328);
nand U217 (N_217,In_1169,In_1625);
nand U218 (N_218,In_1476,In_1810);
or U219 (N_219,In_939,In_406);
nor U220 (N_220,In_335,In_1504);
nor U221 (N_221,In_556,In_1498);
nor U222 (N_222,In_1685,In_226);
or U223 (N_223,In_597,In_1978);
nand U224 (N_224,In_954,In_643);
nand U225 (N_225,In_1804,In_269);
nor U226 (N_226,In_596,In_666);
nand U227 (N_227,In_638,In_675);
nand U228 (N_228,In_1710,In_1303);
or U229 (N_229,In_1290,In_255);
nor U230 (N_230,In_512,In_1576);
nand U231 (N_231,In_982,In_929);
and U232 (N_232,In_1085,In_338);
and U233 (N_233,In_845,In_1829);
nor U234 (N_234,In_1334,In_669);
and U235 (N_235,In_158,In_210);
nand U236 (N_236,In_1349,In_1739);
nor U237 (N_237,In_981,In_419);
or U238 (N_238,In_377,In_670);
or U239 (N_239,In_459,In_443);
or U240 (N_240,In_753,In_179);
or U241 (N_241,In_1494,In_1184);
or U242 (N_242,In_82,In_789);
xnor U243 (N_243,In_1432,In_661);
nand U244 (N_244,In_1761,In_1615);
or U245 (N_245,In_589,In_955);
nand U246 (N_246,In_181,In_133);
nand U247 (N_247,In_743,In_1143);
nor U248 (N_248,In_1018,In_537);
and U249 (N_249,In_1984,In_829);
and U250 (N_250,In_1386,In_1056);
xor U251 (N_251,In_334,In_1481);
nand U252 (N_252,In_1538,In_380);
or U253 (N_253,In_1337,In_1191);
or U254 (N_254,In_195,In_1101);
or U255 (N_255,In_478,In_277);
nor U256 (N_256,In_1064,In_1803);
and U257 (N_257,In_1641,In_744);
or U258 (N_258,In_1857,In_607);
xnor U259 (N_259,In_1799,In_867);
xor U260 (N_260,In_1232,In_129);
and U261 (N_261,In_547,In_733);
or U262 (N_262,In_1911,In_776);
and U263 (N_263,In_508,In_1276);
and U264 (N_264,In_174,In_1690);
or U265 (N_265,In_1253,In_1732);
and U266 (N_266,In_399,In_1901);
and U267 (N_267,In_1469,In_116);
nor U268 (N_268,In_416,In_802);
nor U269 (N_269,In_1841,In_1102);
and U270 (N_270,In_688,In_837);
and U271 (N_271,In_549,In_1228);
xnor U272 (N_272,In_146,In_804);
nand U273 (N_273,In_1172,In_1689);
nand U274 (N_274,In_24,In_156);
or U275 (N_275,In_1593,In_1543);
and U276 (N_276,In_1113,In_87);
nor U277 (N_277,In_1083,In_441);
nor U278 (N_278,In_1049,In_891);
xnor U279 (N_279,In_799,In_237);
or U280 (N_280,In_6,In_938);
and U281 (N_281,In_1350,In_718);
nand U282 (N_282,In_1463,In_1628);
and U283 (N_283,In_588,In_1920);
and U284 (N_284,In_852,In_1825);
nand U285 (N_285,In_1439,In_1426);
or U286 (N_286,In_1704,In_42);
nor U287 (N_287,In_1577,In_1201);
or U288 (N_288,In_1021,In_300);
and U289 (N_289,In_1368,In_70);
nand U290 (N_290,In_175,In_1305);
nor U291 (N_291,In_336,In_495);
nand U292 (N_292,In_777,In_579);
or U293 (N_293,In_389,In_396);
or U294 (N_294,In_68,In_757);
nand U295 (N_295,In_572,In_865);
nor U296 (N_296,In_250,In_1133);
and U297 (N_297,In_1425,In_507);
nor U298 (N_298,In_699,In_258);
and U299 (N_299,In_263,In_1484);
and U300 (N_300,In_1721,In_1058);
nand U301 (N_301,In_1493,In_1356);
nand U302 (N_302,In_722,In_717);
or U303 (N_303,In_903,In_745);
and U304 (N_304,In_969,In_352);
or U305 (N_305,In_640,In_1183);
and U306 (N_306,In_905,In_1682);
and U307 (N_307,In_1834,In_1889);
nand U308 (N_308,In_538,In_1949);
or U309 (N_309,In_728,In_1815);
nand U310 (N_310,In_1199,In_360);
and U311 (N_311,In_678,In_498);
or U312 (N_312,In_1473,In_1994);
or U313 (N_313,In_425,In_1594);
nand U314 (N_314,In_119,In_147);
nor U315 (N_315,In_73,In_1265);
xor U316 (N_316,In_1071,In_551);
nand U317 (N_317,In_1312,In_1786);
nor U318 (N_318,In_870,In_1757);
and U319 (N_319,In_472,In_1124);
nor U320 (N_320,In_1210,In_203);
xnor U321 (N_321,In_10,In_99);
and U322 (N_322,In_1055,In_242);
nor U323 (N_323,In_494,In_340);
or U324 (N_324,In_1934,In_272);
nor U325 (N_325,In_93,In_1454);
or U326 (N_326,In_737,In_1322);
nor U327 (N_327,In_1524,In_206);
or U328 (N_328,In_344,In_712);
nand U329 (N_329,In_862,In_1046);
nand U330 (N_330,In_1468,In_1359);
xnor U331 (N_331,In_1247,In_791);
nand U332 (N_332,In_931,In_1447);
nor U333 (N_333,In_1462,In_1882);
or U334 (N_334,In_627,In_766);
and U335 (N_335,In_1467,In_1868);
nand U336 (N_336,In_362,In_713);
nand U337 (N_337,In_1297,In_1391);
or U338 (N_338,In_1522,In_379);
nor U339 (N_339,In_1162,In_846);
or U340 (N_340,In_1792,In_774);
nor U341 (N_341,In_394,In_677);
nand U342 (N_342,In_1910,In_1658);
nand U343 (N_343,In_836,In_1613);
nor U344 (N_344,In_1041,In_408);
nand U345 (N_345,In_199,In_569);
xor U346 (N_346,In_1330,In_983);
or U347 (N_347,In_1042,In_1159);
nand U348 (N_348,In_557,In_947);
nand U349 (N_349,In_435,In_1050);
nand U350 (N_350,In_1744,In_1194);
nand U351 (N_351,In_492,In_960);
nor U352 (N_352,In_139,In_664);
nand U353 (N_353,In_1315,In_1084);
and U354 (N_354,In_1872,In_1086);
nand U355 (N_355,In_1653,In_1808);
and U356 (N_356,In_499,In_102);
or U357 (N_357,In_1866,In_1397);
nor U358 (N_358,In_1279,In_172);
and U359 (N_359,In_1791,In_1429);
xnor U360 (N_360,In_554,In_1789);
xor U361 (N_361,In_1126,In_586);
xor U362 (N_362,In_168,In_1259);
nand U363 (N_363,In_90,In_222);
nor U364 (N_364,In_1151,In_1552);
nand U365 (N_365,In_1038,In_796);
nand U366 (N_366,In_249,In_1626);
nor U367 (N_367,In_111,In_136);
and U368 (N_368,In_986,In_935);
and U369 (N_369,In_1812,In_1581);
nand U370 (N_370,In_1147,In_1805);
xnor U371 (N_371,In_1422,In_851);
nand U372 (N_372,In_114,In_525);
and U373 (N_373,In_240,In_398);
nor U374 (N_374,In_1718,In_292);
nor U375 (N_375,In_730,In_1026);
nor U376 (N_376,In_1983,In_378);
and U377 (N_377,In_1424,In_611);
or U378 (N_378,In_839,In_80);
nor U379 (N_379,In_978,In_1138);
nor U380 (N_380,In_1818,In_591);
nor U381 (N_381,In_1948,In_1383);
nor U382 (N_382,In_1264,In_1497);
or U383 (N_383,In_901,In_1588);
xor U384 (N_384,In_1695,In_1308);
or U385 (N_385,In_878,In_889);
or U386 (N_386,In_857,In_1030);
nor U387 (N_387,In_192,In_1781);
and U388 (N_388,In_1560,In_313);
xnor U389 (N_389,In_50,In_232);
nand U390 (N_390,In_1736,In_278);
or U391 (N_391,In_530,In_673);
xor U392 (N_392,In_1964,In_1573);
and U393 (N_393,In_1755,In_1939);
nor U394 (N_394,In_347,In_1566);
nor U395 (N_395,In_1583,In_1993);
nand U396 (N_396,In_110,In_1379);
nor U397 (N_397,In_642,In_1556);
nand U398 (N_398,In_1802,In_1400);
nor U399 (N_399,In_467,In_552);
nor U400 (N_400,In_0,In_1788);
nor U401 (N_401,In_261,In_482);
nor U402 (N_402,In_1837,In_751);
nand U403 (N_403,In_768,In_946);
xor U404 (N_404,In_440,In_173);
nand U405 (N_405,In_1696,In_1459);
or U406 (N_406,In_1418,In_1981);
and U407 (N_407,In_196,In_872);
or U408 (N_408,In_1483,In_936);
or U409 (N_409,In_1328,In_1535);
or U410 (N_410,In_927,In_270);
and U411 (N_411,In_1932,In_1262);
or U412 (N_412,In_741,In_1544);
xnor U413 (N_413,In_962,In_1823);
nor U414 (N_414,In_262,In_890);
nor U415 (N_415,In_1809,In_1366);
nand U416 (N_416,In_651,In_62);
nor U417 (N_417,In_1185,In_1048);
and U418 (N_418,In_1317,In_349);
and U419 (N_419,In_306,In_327);
or U420 (N_420,In_1206,In_779);
and U421 (N_421,In_1975,In_550);
or U422 (N_422,In_1161,In_60);
or U423 (N_423,In_325,In_621);
nor U424 (N_424,In_1066,In_1119);
xor U425 (N_425,In_1938,In_619);
and U426 (N_426,In_1205,In_1182);
or U427 (N_427,In_1849,In_81);
xor U428 (N_428,In_30,In_1283);
nand U429 (N_429,In_1709,In_18);
nor U430 (N_430,In_1456,In_363);
or U431 (N_431,In_1157,In_658);
nor U432 (N_432,In_1105,In_1434);
and U433 (N_433,In_190,In_1302);
nor U434 (N_434,In_164,In_1601);
nor U435 (N_435,In_1590,In_1850);
and U436 (N_436,In_624,In_1898);
or U437 (N_437,In_1012,In_1020);
and U438 (N_438,In_1035,In_641);
nor U439 (N_439,In_1270,In_1530);
xnor U440 (N_440,In_916,In_1579);
nor U441 (N_441,In_1111,In_341);
xor U442 (N_442,In_1004,In_1164);
nor U443 (N_443,In_1103,In_1387);
nand U444 (N_444,In_504,In_1783);
or U445 (N_445,In_1643,In_686);
and U446 (N_446,In_637,In_1031);
or U447 (N_447,In_320,In_1112);
nor U448 (N_448,In_1398,In_963);
or U449 (N_449,In_1117,In_1830);
or U450 (N_450,In_246,In_1826);
nand U451 (N_451,In_128,In_15);
nor U452 (N_452,In_1461,In_973);
nand U453 (N_453,In_739,In_1595);
nor U454 (N_454,In_784,In_1173);
nor U455 (N_455,In_886,In_1500);
nand U456 (N_456,In_1408,In_1637);
nor U457 (N_457,In_1148,In_1883);
and U458 (N_458,In_1384,In_365);
nor U459 (N_459,In_868,In_1912);
and U460 (N_460,In_305,In_972);
nand U461 (N_461,In_1223,In_724);
nand U462 (N_462,In_1965,In_473);
nor U463 (N_463,In_696,In_52);
nand U464 (N_464,In_296,In_1073);
and U465 (N_465,In_1240,In_1340);
or U466 (N_466,In_390,In_1518);
nor U467 (N_467,In_1089,In_817);
or U468 (N_468,In_1798,In_1598);
nor U469 (N_469,In_1997,In_1428);
xnor U470 (N_470,In_456,In_1853);
xor U471 (N_471,In_373,In_888);
nor U472 (N_472,In_1075,In_1077);
nand U473 (N_473,In_371,In_1748);
and U474 (N_474,In_841,In_1474);
xor U475 (N_475,In_899,In_902);
or U476 (N_476,In_806,In_1811);
nand U477 (N_477,In_881,In_684);
nand U478 (N_478,In_1163,In_1659);
nor U479 (N_479,In_267,In_1238);
and U480 (N_480,In_701,In_1430);
nand U481 (N_481,In_1725,In_706);
and U482 (N_482,In_1928,In_1482);
xor U483 (N_483,In_542,In_765);
and U484 (N_484,In_778,In_1652);
nand U485 (N_485,In_906,In_7);
xor U486 (N_486,In_580,In_259);
nor U487 (N_487,In_1989,In_1186);
and U488 (N_488,In_1008,In_1701);
or U489 (N_489,In_1869,In_383);
nand U490 (N_490,In_1254,In_36);
and U491 (N_491,In_1562,In_1363);
or U492 (N_492,In_1217,In_1925);
or U493 (N_493,In_16,In_1239);
or U494 (N_494,In_439,In_1440);
xnor U495 (N_495,In_1773,In_1980);
and U496 (N_496,In_940,In_1306);
and U497 (N_497,In_56,In_683);
nor U498 (N_498,In_1585,In_319);
nand U499 (N_499,In_475,In_309);
and U500 (N_500,In_1726,In_449);
or U501 (N_501,In_1381,In_1189);
and U502 (N_502,In_47,In_141);
nor U503 (N_503,In_33,In_1784);
nor U504 (N_504,In_698,In_697);
nand U505 (N_505,In_809,In_387);
and U506 (N_506,In_420,In_1724);
and U507 (N_507,In_31,In_1990);
nand U508 (N_508,In_1877,In_200);
nor U509 (N_509,In_1486,In_471);
or U510 (N_510,In_919,In_350);
nor U511 (N_511,In_904,In_339);
or U512 (N_512,In_1847,In_1957);
or U513 (N_513,In_1519,In_1559);
nor U514 (N_514,In_198,In_606);
or U515 (N_515,In_1536,In_1878);
and U516 (N_516,In_660,In_795);
and U517 (N_517,In_1491,In_1554);
or U518 (N_518,In_1294,In_21);
nor U519 (N_519,In_17,In_1108);
or U520 (N_520,In_1702,In_599);
and U521 (N_521,In_1763,In_1664);
nand U522 (N_522,In_1754,In_1700);
xor U523 (N_523,In_1171,In_1961);
nor U524 (N_524,In_329,In_321);
and U525 (N_525,In_1974,In_615);
nand U526 (N_526,In_1852,In_385);
and U527 (N_527,In_654,In_1114);
and U528 (N_528,In_1342,In_1569);
and U529 (N_529,In_197,In_1735);
or U530 (N_530,In_13,In_814);
nor U531 (N_531,In_856,In_1897);
and U532 (N_532,In_543,In_1455);
or U533 (N_533,In_1450,In_1246);
xor U534 (N_534,In_1991,In_708);
nor U535 (N_535,In_930,In_797);
and U536 (N_536,In_145,In_1663);
nand U537 (N_537,In_1548,In_662);
nand U538 (N_538,In_1141,In_461);
and U539 (N_539,In_1557,In_1170);
nand U540 (N_540,In_490,In_483);
nor U541 (N_541,In_1720,In_1863);
xor U542 (N_542,In_1096,In_368);
and U543 (N_543,In_1614,In_1654);
nor U544 (N_544,In_1797,In_1343);
nand U545 (N_545,In_40,In_284);
nand U546 (N_546,In_35,In_29);
or U547 (N_547,In_1723,In_1551);
and U548 (N_548,In_1014,In_137);
or U549 (N_549,In_961,In_79);
nor U550 (N_550,In_1616,In_1730);
and U551 (N_551,In_1620,In_1870);
and U552 (N_552,In_546,In_228);
and U553 (N_553,In_1175,In_1061);
xor U554 (N_554,In_1295,In_460);
nor U555 (N_555,In_268,In_1988);
nor U556 (N_556,In_115,In_875);
or U557 (N_557,In_86,In_205);
or U558 (N_558,In_1168,In_1843);
nand U559 (N_559,In_1604,In_1816);
nand U560 (N_560,In_28,In_1496);
and U561 (N_561,In_1222,In_1779);
nand U562 (N_562,In_280,In_632);
xnor U563 (N_563,In_944,In_1999);
or U564 (N_564,In_1622,In_364);
nor U565 (N_565,In_44,In_1651);
and U566 (N_566,In_170,In_843);
nand U567 (N_567,In_942,In_1052);
xnor U568 (N_568,In_937,In_1022);
nor U569 (N_569,In_109,In_230);
nand U570 (N_570,In_1982,In_561);
or U571 (N_571,In_361,In_1074);
or U572 (N_572,In_734,In_655);
or U573 (N_573,In_446,In_1341);
xnor U574 (N_574,In_1862,In_1070);
and U575 (N_575,In_1969,In_923);
nand U576 (N_576,In_1790,In_1057);
and U577 (N_577,In_1656,In_1360);
nand U578 (N_578,In_1068,In_22);
nand U579 (N_579,In_951,In_307);
nand U580 (N_580,In_159,In_1441);
or U581 (N_581,In_303,In_220);
or U582 (N_582,In_1824,In_1417);
nand U583 (N_583,In_155,In_1527);
nand U584 (N_584,In_20,In_132);
nor U585 (N_585,In_67,In_685);
and U586 (N_586,In_1992,In_140);
and U587 (N_587,In_1574,In_1125);
and U588 (N_588,In_995,In_92);
nand U589 (N_589,In_1475,In_1490);
nor U590 (N_590,In_1845,In_123);
xnor U591 (N_591,In_407,In_1352);
nand U592 (N_592,In_1521,In_1793);
nor U593 (N_593,In_1193,In_1072);
nor U594 (N_594,In_587,In_427);
or U595 (N_595,In_1942,In_590);
and U596 (N_596,In_1095,In_925);
or U597 (N_597,In_1687,In_414);
nand U598 (N_598,In_676,In_659);
nand U599 (N_599,In_1044,In_1918);
and U600 (N_600,In_1320,In_49);
nand U601 (N_601,In_216,In_1036);
nand U602 (N_602,In_711,In_721);
or U603 (N_603,In_1533,In_509);
and U604 (N_604,In_1986,In_1006);
and U605 (N_605,In_1621,In_1624);
and U606 (N_606,In_855,In_1515);
or U607 (N_607,In_126,In_171);
or U608 (N_608,In_540,In_1512);
or U609 (N_609,In_1414,In_592);
nor U610 (N_610,In_1612,In_1778);
nor U611 (N_611,In_1617,In_524);
nor U612 (N_612,In_1213,In_1065);
and U613 (N_613,In_873,In_1378);
nor U614 (N_614,In_1645,In_1321);
or U615 (N_615,In_648,In_649);
or U616 (N_616,In_163,In_331);
nand U617 (N_617,In_465,In_1132);
or U618 (N_618,In_214,In_1692);
nand U619 (N_619,In_1288,In_1309);
or U620 (N_620,In_792,In_952);
xnor U621 (N_621,In_634,In_1431);
nand U622 (N_622,In_1859,In_166);
and U623 (N_623,In_519,In_1196);
or U624 (N_624,In_486,In_1584);
xnor U625 (N_625,In_1996,In_824);
nor U626 (N_626,In_55,In_1094);
and U627 (N_627,In_1137,In_785);
and U628 (N_628,In_322,In_1979);
or U629 (N_629,In_1760,In_769);
or U630 (N_630,In_1130,In_103);
xnor U631 (N_631,In_1367,In_1954);
nor U632 (N_632,In_318,In_480);
nor U633 (N_633,In_451,In_1487);
or U634 (N_634,In_956,In_1706);
xnor U635 (N_635,In_926,In_476);
or U636 (N_636,In_1599,In_924);
nand U637 (N_637,In_1832,In_497);
and U638 (N_638,In_1842,In_748);
nand U639 (N_639,In_783,In_544);
nand U640 (N_640,In_1332,In_1508);
nand U641 (N_641,In_185,In_564);
xor U642 (N_642,In_401,In_1796);
xnor U643 (N_643,In_964,In_1292);
xnor U644 (N_644,In_535,In_1902);
nor U645 (N_645,In_1567,In_1844);
or U646 (N_646,In_430,In_974);
or U647 (N_647,In_1913,In_842);
nor U648 (N_648,In_1998,In_291);
xor U649 (N_649,In_91,In_1591);
nand U650 (N_650,In_1029,In_529);
xor U651 (N_651,In_1470,In_689);
nand U652 (N_652,In_247,In_668);
nand U653 (N_653,In_1449,In_992);
xor U654 (N_654,In_3,In_644);
and U655 (N_655,In_1088,In_1098);
or U656 (N_656,In_1033,In_493);
or U657 (N_657,In_283,In_1931);
or U658 (N_658,In_794,In_1435);
nor U659 (N_659,In_294,In_178);
nor U660 (N_660,In_316,In_691);
and U661 (N_661,In_422,In_1972);
xor U662 (N_662,In_77,In_1123);
and U663 (N_663,In_1906,In_726);
nand U664 (N_664,In_1080,In_1586);
nor U665 (N_665,In_681,In_85);
nand U666 (N_666,In_1423,In_915);
xnor U667 (N_667,In_487,In_1099);
xor U668 (N_668,In_603,In_189);
nand U669 (N_669,In_297,In_631);
and U670 (N_670,In_358,In_1136);
or U671 (N_671,In_1282,In_1678);
nor U672 (N_672,In_819,In_548);
and U673 (N_673,In_521,In_1480);
and U674 (N_674,In_469,In_1202);
and U675 (N_675,In_1564,In_1657);
and U676 (N_676,In_1923,In_1127);
nor U677 (N_677,In_204,In_276);
or U678 (N_678,In_1216,In_1819);
nand U679 (N_679,In_308,In_1167);
nand U680 (N_680,In_215,In_1740);
and U681 (N_681,In_423,In_1139);
nand U682 (N_682,In_1255,In_866);
and U683 (N_683,In_357,In_32);
nand U684 (N_684,In_289,In_279);
nand U685 (N_685,In_332,In_907);
and U686 (N_686,In_562,In_605);
or U687 (N_687,In_1219,In_1361);
or U688 (N_688,In_1728,In_874);
or U689 (N_689,In_1640,In_1703);
and U690 (N_690,In_1446,In_1716);
and U691 (N_691,In_1051,In_705);
and U692 (N_692,In_945,In_1995);
xnor U693 (N_693,In_1752,In_1034);
nand U694 (N_694,In_1705,In_1230);
or U695 (N_695,In_604,In_1603);
and U696 (N_696,In_1930,In_317);
or U697 (N_697,In_1415,In_719);
or U698 (N_698,In_359,In_985);
or U699 (N_699,In_828,In_1402);
and U700 (N_700,In_1840,In_5);
nor U701 (N_701,In_1062,In_1001);
and U702 (N_702,In_1128,In_833);
nand U703 (N_703,In_1218,In_869);
or U704 (N_704,In_1344,In_113);
nor U705 (N_705,In_1501,In_501);
and U706 (N_706,In_1668,In_1177);
xnor U707 (N_707,In_207,In_1465);
and U708 (N_708,In_1260,In_464);
nor U709 (N_709,In_1592,In_1550);
nand U710 (N_710,In_1374,In_421);
or U711 (N_711,In_932,In_1263);
nor U712 (N_712,In_735,In_1745);
nand U713 (N_713,In_1864,In_1097);
nand U714 (N_714,In_391,In_800);
or U715 (N_715,In_1578,In_1746);
and U716 (N_716,In_694,In_593);
nor U717 (N_717,In_108,In_1770);
and U718 (N_718,In_1153,In_1372);
nand U719 (N_719,In_1335,In_520);
nand U720 (N_720,In_176,In_1243);
nand U721 (N_721,In_187,In_617);
xnor U722 (N_722,In_1365,In_1629);
nor U723 (N_723,In_1445,In_1886);
and U724 (N_724,In_1351,In_1776);
xnor U725 (N_725,In_1782,In_84);
nor U726 (N_726,In_324,In_413);
nor U727 (N_727,In_679,In_1406);
and U728 (N_728,In_1854,In_1885);
nand U729 (N_729,In_1188,In_1060);
xnor U730 (N_730,In_1899,In_1686);
nand U731 (N_731,In_453,In_1831);
and U732 (N_732,In_1520,In_764);
and U733 (N_733,In_326,In_581);
or U734 (N_734,In_1919,In_861);
nor U735 (N_735,In_1198,In_702);
or U736 (N_736,In_834,In_1327);
or U737 (N_737,In_898,In_500);
nand U738 (N_738,In_1909,In_433);
nand U739 (N_739,In_1941,In_23);
and U740 (N_740,In_1388,In_1764);
nand U741 (N_741,In_100,In_1684);
or U742 (N_742,In_813,In_1631);
and U743 (N_743,In_853,In_1158);
or U744 (N_744,In_849,In_1252);
and U745 (N_745,In_1362,In_656);
or U746 (N_746,In_1311,In_1433);
and U747 (N_747,In_1738,In_1286);
or U748 (N_748,In_553,In_1855);
and U749 (N_749,In_810,In_1165);
nor U750 (N_750,In_680,In_808);
nor U751 (N_751,In_832,In_948);
and U752 (N_752,In_513,In_1274);
nand U753 (N_753,In_527,In_293);
and U754 (N_754,In_1633,In_58);
nand U755 (N_755,In_1155,In_244);
xor U756 (N_756,In_431,In_1699);
nand U757 (N_757,In_536,In_1373);
nor U758 (N_758,In_217,In_848);
or U759 (N_759,In_1250,In_78);
nor U760 (N_760,In_894,In_183);
nand U761 (N_761,In_1200,In_354);
nor U762 (N_762,In_555,In_1731);
nor U763 (N_763,In_105,In_1741);
or U764 (N_764,In_760,In_1713);
and U765 (N_765,In_1693,In_690);
nor U766 (N_766,In_1729,In_1396);
or U767 (N_767,In_1528,In_1596);
or U768 (N_768,In_1291,In_622);
nor U769 (N_769,In_871,In_811);
nand U770 (N_770,In_1412,In_533);
nor U771 (N_771,In_1419,In_264);
nand U772 (N_772,In_51,In_1924);
or U773 (N_773,In_1296,In_1118);
or U774 (N_774,In_1609,In_130);
or U775 (N_775,In_1623,In_1275);
or U776 (N_776,In_910,In_388);
and U777 (N_777,In_72,In_253);
and U778 (N_778,In_727,In_1149);
or U779 (N_779,In_1630,In_1319);
and U780 (N_780,In_477,In_1505);
nand U781 (N_781,In_426,In_922);
or U782 (N_782,In_772,In_575);
nor U783 (N_783,In_720,In_672);
and U784 (N_784,In_1395,In_1777);
nor U785 (N_785,In_831,In_1212);
nand U786 (N_786,In_1326,In_773);
and U787 (N_787,In_1318,In_1646);
nor U788 (N_788,In_732,In_746);
nor U789 (N_789,In_893,In_1549);
or U790 (N_790,In_234,In_921);
nand U791 (N_791,In_1348,In_1347);
nor U792 (N_792,In_386,In_1943);
and U793 (N_793,In_1489,In_65);
and U794 (N_794,In_1225,In_1382);
nor U795 (N_795,In_1727,In_1717);
nand U796 (N_796,In_496,In_1116);
and U797 (N_797,In_1848,In_194);
and U798 (N_798,In_863,In_104);
and U799 (N_799,In_1903,In_481);
xor U800 (N_800,In_470,In_1385);
and U801 (N_801,In_781,In_1814);
or U802 (N_802,In_1115,In_582);
and U803 (N_803,In_574,In_57);
nor U804 (N_804,In_479,In_1929);
or U805 (N_805,In_167,In_571);
or U806 (N_806,In_1370,In_1900);
or U807 (N_807,In_1513,In_1271);
or U808 (N_808,In_1774,In_218);
nor U809 (N_809,In_112,In_840);
or U810 (N_810,In_793,In_1600);
nand U811 (N_811,In_131,In_1822);
or U812 (N_812,In_1967,In_1187);
nand U813 (N_813,In_1608,In_539);
nor U814 (N_814,In_1331,In_1955);
and U815 (N_815,In_1221,In_1953);
nand U816 (N_816,In_984,In_883);
nand U817 (N_817,In_1926,In_830);
nor U818 (N_818,In_489,In_1677);
nor U819 (N_819,In_161,In_731);
nand U820 (N_820,In_585,In_850);
or U821 (N_821,In_330,In_256);
nor U822 (N_822,In_1916,In_428);
nor U823 (N_823,In_667,In_1227);
and U824 (N_824,In_859,In_1160);
and U825 (N_825,In_260,In_1011);
and U826 (N_826,In_1236,In_370);
or U827 (N_827,In_154,In_298);
and U828 (N_828,In_1144,In_1277);
and U829 (N_829,In_1526,In_1010);
or U830 (N_830,In_135,In_1838);
or U831 (N_831,In_1376,In_628);
and U832 (N_832,In_1722,In_633);
and U833 (N_833,In_19,In_1081);
nand U834 (N_834,In_987,In_76);
or U835 (N_835,In_911,In_248);
and U836 (N_836,In_120,In_238);
and U837 (N_837,In_710,In_1606);
nand U838 (N_838,In_1338,In_1047);
and U839 (N_839,In_366,In_1836);
xnor U840 (N_840,In_988,In_1768);
or U841 (N_841,In_1442,In_231);
nor U842 (N_842,In_1821,In_1407);
nand U843 (N_843,In_1669,In_1110);
nor U844 (N_844,In_1364,In_39);
or U845 (N_845,In_997,In_1220);
or U846 (N_846,In_908,In_827);
or U847 (N_847,In_1339,In_1479);
or U848 (N_848,In_1856,In_69);
nand U849 (N_849,In_1806,In_583);
or U850 (N_850,In_880,In_756);
nand U851 (N_851,In_1963,In_162);
and U852 (N_852,In_714,In_1618);
or U853 (N_853,In_148,In_1905);
and U854 (N_854,In_1970,In_95);
nor U855 (N_855,In_762,In_245);
or U856 (N_856,In_1711,In_965);
or U857 (N_857,In_1769,In_650);
and U858 (N_858,In_996,In_395);
nor U859 (N_859,In_1827,In_251);
and U860 (N_860,In_1800,In_315);
or U861 (N_861,In_1794,In_884);
nand U862 (N_862,In_1015,In_1861);
or U863 (N_863,In_682,In_1453);
nand U864 (N_864,In_367,In_184);
and U865 (N_865,In_1958,In_1759);
nor U866 (N_866,In_125,In_96);
nor U867 (N_867,In_1751,In_567);
nor U868 (N_868,In_518,In_299);
xnor U869 (N_869,In_188,In_1532);
nor U870 (N_870,In_1503,In_1795);
nor U871 (N_871,In_227,In_1639);
nand U872 (N_872,In_66,In_1697);
nor U873 (N_873,In_193,In_818);
nor U874 (N_874,In_1753,In_63);
nand U875 (N_875,In_1881,In_1742);
and U876 (N_876,In_594,In_127);
nor U877 (N_877,In_1747,In_1541);
and U878 (N_878,In_790,In_1951);
or U879 (N_879,In_287,In_94);
nand U880 (N_880,In_1403,In_1393);
and U881 (N_881,In_1289,In_1024);
nand U882 (N_882,In_343,In_532);
nor U883 (N_883,In_142,In_1471);
and U884 (N_884,In_1053,In_1224);
xnor U885 (N_885,In_1875,In_265);
or U886 (N_886,In_771,In_98);
nor U887 (N_887,In_1032,In_474);
nand U888 (N_888,In_1529,In_1215);
nand U889 (N_889,In_1017,In_1514);
or U890 (N_890,In_822,In_169);
or U891 (N_891,In_1915,In_225);
or U892 (N_892,In_775,In_736);
and U893 (N_893,In_1785,In_53);
or U894 (N_894,In_1472,In_630);
and U895 (N_895,In_41,In_1134);
or U896 (N_896,In_565,In_1413);
xor U897 (N_897,In_25,In_288);
xor U898 (N_898,In_1466,In_1672);
xor U899 (N_899,In_1197,In_1960);
or U900 (N_900,In_763,In_807);
xor U901 (N_901,In_1394,In_1495);
or U902 (N_902,In_1947,In_434);
and U903 (N_903,In_1357,In_920);
or U904 (N_904,In_1534,In_1460);
nand U905 (N_905,In_337,In_254);
xnor U906 (N_906,In_304,In_1145);
nand U907 (N_907,In_462,In_826);
xnor U908 (N_908,In_1325,In_1772);
nor U909 (N_909,In_1345,In_1410);
nand U910 (N_910,In_847,In_1851);
or U911 (N_911,In_1917,In_1673);
nor U912 (N_912,In_860,In_1492);
and U913 (N_913,In_1893,In_211);
and U914 (N_914,In_1638,In_1285);
xnor U915 (N_915,In_895,In_1619);
nand U916 (N_916,In_1195,In_957);
nand U917 (N_917,In_271,In_1438);
nor U918 (N_918,In_1507,In_742);
nor U919 (N_919,In_522,In_1610);
or U920 (N_920,In_252,In_400);
xor U921 (N_921,In_37,In_1280);
xor U922 (N_922,In_528,In_1208);
nor U923 (N_923,In_1448,In_1935);
and U924 (N_924,In_424,In_1558);
nor U925 (N_925,In_302,In_1828);
and U926 (N_926,In_404,In_285);
nand U927 (N_927,In_48,In_1936);
or U928 (N_928,In_729,In_1043);
nor U929 (N_929,In_1545,In_1775);
nor U930 (N_930,In_1079,In_149);
or U931 (N_931,In_1516,In_1976);
nor U932 (N_932,In_1502,In_1896);
or U933 (N_933,In_1860,In_761);
or U934 (N_934,In_1499,In_182);
nand U935 (N_935,In_1100,In_598);
nand U936 (N_936,In_1611,In_1714);
nor U937 (N_937,In_1181,In_1565);
nand U938 (N_938,In_1820,In_1142);
nor U939 (N_939,In_1956,In_429);
nor U940 (N_940,In_1420,In_46);
nor U941 (N_941,In_1003,In_138);
or U942 (N_942,In_1571,In_61);
xor U943 (N_943,In_754,In_657);
nor U944 (N_944,In_755,In_740);
nor U945 (N_945,In_353,In_157);
xnor U946 (N_946,In_523,In_1488);
nor U947 (N_947,In_623,In_1968);
or U948 (N_948,In_1921,In_213);
nand U949 (N_949,In_786,In_1537);
or U950 (N_950,In_1266,In_1156);
and U951 (N_951,In_1436,In_1880);
or U952 (N_952,In_1523,In_484);
and U953 (N_953,In_877,In_1634);
xor U954 (N_954,In_980,In_1179);
or U955 (N_955,In_584,In_2);
nor U956 (N_956,In_1409,In_1235);
nand U957 (N_957,In_1027,In_614);
and U958 (N_958,In_1269,In_323);
nor U959 (N_959,In_1478,In_1301);
nor U960 (N_960,In_993,In_1059);
nor U961 (N_961,In_647,In_1293);
nor U962 (N_962,In_534,In_1093);
nand U963 (N_963,In_412,In_1267);
nor U964 (N_964,In_616,In_1392);
nor U965 (N_965,In_1152,In_311);
and U966 (N_966,In_1063,In_202);
and U967 (N_967,In_639,In_1009);
and U968 (N_968,In_101,In_959);
or U969 (N_969,In_122,In_1427);
nor U970 (N_970,In_1636,In_229);
nand U971 (N_971,In_11,In_573);
and U972 (N_972,In_1457,In_700);
nand U973 (N_973,In_1542,In_219);
nor U974 (N_974,In_1937,In_1933);
nor U975 (N_975,In_1107,In_526);
nor U976 (N_976,In_1016,In_402);
nand U977 (N_977,In_282,In_1767);
nor U978 (N_978,In_152,In_1257);
nand U979 (N_979,In_1353,In_820);
and U980 (N_980,In_864,In_1140);
xnor U981 (N_981,In_417,In_1039);
nand U982 (N_982,In_515,In_1411);
nand U983 (N_983,In_186,In_1067);
nand U984 (N_984,In_1648,In_1715);
and U985 (N_985,In_1907,In_943);
nand U986 (N_986,In_491,In_578);
or U987 (N_987,In_1985,In_1245);
and U988 (N_988,In_1858,In_1719);
nand U989 (N_989,In_1575,In_570);
xnor U990 (N_990,In_770,In_1895);
nor U991 (N_991,In_1313,In_1602);
nand U992 (N_992,In_704,In_1477);
nand U993 (N_993,In_1517,In_1952);
nand U994 (N_994,In_392,In_1506);
nand U995 (N_995,In_1166,In_1666);
nor U996 (N_996,In_1914,In_393);
or U997 (N_997,In_405,In_201);
and U998 (N_998,In_1007,In_241);
and U999 (N_999,In_71,In_815);
and U1000 (N_1000,N_728,N_607);
xnor U1001 (N_1001,N_870,N_893);
or U1002 (N_1002,N_213,N_748);
nand U1003 (N_1003,N_152,N_765);
xnor U1004 (N_1004,N_663,N_10);
nor U1005 (N_1005,N_348,N_465);
nand U1006 (N_1006,N_442,N_509);
or U1007 (N_1007,N_744,N_353);
and U1008 (N_1008,N_369,N_515);
and U1009 (N_1009,N_148,N_453);
and U1010 (N_1010,N_492,N_244);
and U1011 (N_1011,N_682,N_814);
or U1012 (N_1012,N_676,N_538);
nor U1013 (N_1013,N_647,N_409);
xor U1014 (N_1014,N_6,N_440);
nor U1015 (N_1015,N_579,N_364);
nand U1016 (N_1016,N_845,N_43);
and U1017 (N_1017,N_424,N_727);
and U1018 (N_1018,N_432,N_464);
nand U1019 (N_1019,N_876,N_127);
and U1020 (N_1020,N_360,N_521);
and U1021 (N_1021,N_762,N_670);
xnor U1022 (N_1022,N_150,N_821);
nor U1023 (N_1023,N_130,N_417);
nor U1024 (N_1024,N_566,N_959);
and U1025 (N_1025,N_236,N_883);
nand U1026 (N_1026,N_71,N_459);
or U1027 (N_1027,N_90,N_486);
nand U1028 (N_1028,N_720,N_422);
or U1029 (N_1029,N_534,N_795);
nand U1030 (N_1030,N_84,N_114);
or U1031 (N_1031,N_927,N_903);
nor U1032 (N_1032,N_366,N_397);
or U1033 (N_1033,N_615,N_441);
and U1034 (N_1034,N_338,N_98);
nor U1035 (N_1035,N_241,N_940);
nor U1036 (N_1036,N_268,N_763);
or U1037 (N_1037,N_574,N_306);
nand U1038 (N_1038,N_643,N_318);
nor U1039 (N_1039,N_507,N_740);
or U1040 (N_1040,N_350,N_828);
or U1041 (N_1041,N_860,N_672);
nor U1042 (N_1042,N_855,N_365);
and U1043 (N_1043,N_657,N_184);
nor U1044 (N_1044,N_550,N_957);
and U1045 (N_1045,N_910,N_882);
nand U1046 (N_1046,N_368,N_645);
or U1047 (N_1047,N_518,N_548);
and U1048 (N_1048,N_337,N_66);
and U1049 (N_1049,N_125,N_841);
or U1050 (N_1050,N_880,N_649);
and U1051 (N_1051,N_951,N_339);
nand U1052 (N_1052,N_864,N_430);
xnor U1053 (N_1053,N_392,N_960);
xnor U1054 (N_1054,N_363,N_954);
nand U1055 (N_1055,N_59,N_609);
nand U1056 (N_1056,N_801,N_810);
and U1057 (N_1057,N_990,N_89);
nand U1058 (N_1058,N_620,N_804);
and U1059 (N_1059,N_5,N_640);
or U1060 (N_1060,N_384,N_275);
or U1061 (N_1061,N_314,N_919);
nand U1062 (N_1062,N_224,N_662);
and U1063 (N_1063,N_242,N_343);
and U1064 (N_1064,N_258,N_310);
nand U1065 (N_1065,N_683,N_264);
nor U1066 (N_1066,N_323,N_266);
nand U1067 (N_1067,N_401,N_939);
or U1068 (N_1068,N_235,N_595);
nand U1069 (N_1069,N_28,N_522);
nand U1070 (N_1070,N_287,N_722);
and U1071 (N_1071,N_375,N_158);
nor U1072 (N_1072,N_109,N_774);
and U1073 (N_1073,N_460,N_161);
nor U1074 (N_1074,N_508,N_93);
nor U1075 (N_1075,N_716,N_496);
nor U1076 (N_1076,N_498,N_450);
xnor U1077 (N_1077,N_965,N_183);
or U1078 (N_1078,N_556,N_379);
and U1079 (N_1079,N_691,N_284);
nand U1080 (N_1080,N_351,N_808);
and U1081 (N_1081,N_151,N_177);
nor U1082 (N_1082,N_833,N_229);
nor U1083 (N_1083,N_978,N_573);
nand U1084 (N_1084,N_112,N_391);
nand U1085 (N_1085,N_584,N_825);
nor U1086 (N_1086,N_793,N_991);
nand U1087 (N_1087,N_488,N_915);
or U1088 (N_1088,N_600,N_297);
and U1089 (N_1089,N_104,N_582);
or U1090 (N_1090,N_688,N_1);
nor U1091 (N_1091,N_525,N_996);
nand U1092 (N_1092,N_116,N_283);
and U1093 (N_1093,N_377,N_106);
nor U1094 (N_1094,N_948,N_862);
nand U1095 (N_1095,N_334,N_160);
or U1096 (N_1096,N_178,N_627);
nand U1097 (N_1097,N_25,N_249);
and U1098 (N_1098,N_8,N_265);
or U1099 (N_1099,N_228,N_324);
nor U1100 (N_1100,N_926,N_270);
nand U1101 (N_1101,N_540,N_24);
nor U1102 (N_1102,N_194,N_868);
and U1103 (N_1103,N_884,N_282);
nand U1104 (N_1104,N_779,N_537);
xnor U1105 (N_1105,N_83,N_513);
xnor U1106 (N_1106,N_9,N_934);
or U1107 (N_1107,N_245,N_239);
nand U1108 (N_1108,N_185,N_588);
nand U1109 (N_1109,N_163,N_555);
and U1110 (N_1110,N_591,N_966);
nor U1111 (N_1111,N_705,N_157);
nor U1112 (N_1112,N_373,N_697);
nand U1113 (N_1113,N_930,N_359);
nor U1114 (N_1114,N_665,N_356);
nor U1115 (N_1115,N_931,N_822);
nand U1116 (N_1116,N_389,N_945);
nand U1117 (N_1117,N_388,N_979);
and U1118 (N_1118,N_427,N_787);
nand U1119 (N_1119,N_520,N_958);
nand U1120 (N_1120,N_302,N_172);
and U1121 (N_1121,N_593,N_802);
xnor U1122 (N_1122,N_803,N_867);
nand U1123 (N_1123,N_374,N_712);
nor U1124 (N_1124,N_501,N_3);
and U1125 (N_1125,N_198,N_526);
nand U1126 (N_1126,N_218,N_973);
nand U1127 (N_1127,N_737,N_431);
and U1128 (N_1128,N_599,N_136);
xnor U1129 (N_1129,N_731,N_552);
nand U1130 (N_1130,N_267,N_659);
nand U1131 (N_1131,N_666,N_576);
or U1132 (N_1132,N_642,N_54);
or U1133 (N_1133,N_820,N_685);
nor U1134 (N_1134,N_942,N_138);
and U1135 (N_1135,N_653,N_468);
nand U1136 (N_1136,N_562,N_704);
xor U1137 (N_1137,N_771,N_72);
or U1138 (N_1138,N_15,N_143);
or U1139 (N_1139,N_110,N_101);
nor U1140 (N_1140,N_625,N_546);
or U1141 (N_1141,N_458,N_211);
and U1142 (N_1142,N_758,N_141);
xnor U1143 (N_1143,N_97,N_896);
and U1144 (N_1144,N_128,N_411);
and U1145 (N_1145,N_517,N_543);
or U1146 (N_1146,N_655,N_840);
or U1147 (N_1147,N_332,N_233);
and U1148 (N_1148,N_289,N_336);
or U1149 (N_1149,N_131,N_524);
or U1150 (N_1150,N_61,N_37);
and U1151 (N_1151,N_73,N_307);
and U1152 (N_1152,N_908,N_901);
or U1153 (N_1153,N_293,N_230);
nand U1154 (N_1154,N_673,N_129);
nand U1155 (N_1155,N_767,N_21);
nor U1156 (N_1156,N_118,N_191);
xor U1157 (N_1157,N_192,N_719);
nand U1158 (N_1158,N_680,N_631);
xor U1159 (N_1159,N_176,N_126);
nor U1160 (N_1160,N_0,N_361);
xor U1161 (N_1161,N_195,N_478);
nor U1162 (N_1162,N_577,N_715);
nand U1163 (N_1163,N_493,N_528);
or U1164 (N_1164,N_756,N_443);
and U1165 (N_1165,N_506,N_564);
nor U1166 (N_1166,N_181,N_541);
nand U1167 (N_1167,N_905,N_906);
nor U1168 (N_1168,N_207,N_637);
xor U1169 (N_1169,N_352,N_120);
nand U1170 (N_1170,N_619,N_405);
or U1171 (N_1171,N_31,N_123);
nand U1172 (N_1172,N_571,N_964);
or U1173 (N_1173,N_45,N_726);
nor U1174 (N_1174,N_829,N_75);
and U1175 (N_1175,N_113,N_22);
nor U1176 (N_1176,N_725,N_234);
and U1177 (N_1177,N_786,N_82);
or U1178 (N_1178,N_18,N_86);
nand U1179 (N_1179,N_572,N_596);
or U1180 (N_1180,N_40,N_985);
nor U1181 (N_1181,N_407,N_861);
nor U1182 (N_1182,N_900,N_987);
nor U1183 (N_1183,N_690,N_357);
nor U1184 (N_1184,N_792,N_830);
or U1185 (N_1185,N_286,N_209);
or U1186 (N_1186,N_156,N_344);
or U1187 (N_1187,N_590,N_606);
nor U1188 (N_1188,N_203,N_300);
or U1189 (N_1189,N_429,N_844);
or U1190 (N_1190,N_408,N_937);
xnor U1191 (N_1191,N_962,N_484);
nor U1192 (N_1192,N_77,N_248);
and U1193 (N_1193,N_39,N_400);
nor U1194 (N_1194,N_404,N_684);
or U1195 (N_1195,N_699,N_916);
nor U1196 (N_1196,N_797,N_50);
nand U1197 (N_1197,N_839,N_479);
nand U1198 (N_1198,N_929,N_633);
nor U1199 (N_1199,N_240,N_626);
or U1200 (N_1200,N_445,N_274);
or U1201 (N_1201,N_581,N_658);
xnor U1202 (N_1202,N_144,N_291);
nor U1203 (N_1203,N_761,N_623);
and U1204 (N_1204,N_886,N_835);
or U1205 (N_1205,N_621,N_617);
or U1206 (N_1206,N_696,N_602);
nor U1207 (N_1207,N_466,N_276);
or U1208 (N_1208,N_542,N_856);
nand U1209 (N_1209,N_674,N_159);
or U1210 (N_1210,N_410,N_372);
or U1211 (N_1211,N_162,N_738);
and U1212 (N_1212,N_199,N_490);
and U1213 (N_1213,N_135,N_523);
nand U1214 (N_1214,N_296,N_333);
and U1215 (N_1215,N_639,N_187);
xnor U1216 (N_1216,N_186,N_694);
and U1217 (N_1217,N_201,N_610);
or U1218 (N_1218,N_817,N_362);
nor U1219 (N_1219,N_656,N_170);
and U1220 (N_1220,N_935,N_438);
nor U1221 (N_1221,N_747,N_76);
nor U1222 (N_1222,N_68,N_335);
xnor U1223 (N_1223,N_798,N_536);
nor U1224 (N_1224,N_706,N_29);
and U1225 (N_1225,N_827,N_980);
xor U1226 (N_1226,N_549,N_371);
and U1227 (N_1227,N_67,N_512);
or U1228 (N_1228,N_741,N_250);
and U1229 (N_1229,N_2,N_132);
or U1230 (N_1230,N_974,N_257);
and U1231 (N_1231,N_46,N_532);
nand U1232 (N_1232,N_586,N_435);
nor U1233 (N_1233,N_853,N_231);
nand U1234 (N_1234,N_452,N_563);
or U1235 (N_1235,N_342,N_601);
and U1236 (N_1236,N_956,N_597);
nand U1237 (N_1237,N_622,N_999);
and U1238 (N_1238,N_122,N_88);
or U1239 (N_1239,N_800,N_225);
nor U1240 (N_1240,N_654,N_754);
xnor U1241 (N_1241,N_341,N_48);
nand U1242 (N_1242,N_354,N_628);
or U1243 (N_1243,N_133,N_834);
nor U1244 (N_1244,N_42,N_475);
xnor U1245 (N_1245,N_847,N_474);
nand U1246 (N_1246,N_585,N_32);
nand U1247 (N_1247,N_85,N_519);
nor U1248 (N_1248,N_155,N_304);
nand U1249 (N_1249,N_885,N_567);
or U1250 (N_1250,N_851,N_646);
and U1251 (N_1251,N_873,N_325);
nor U1252 (N_1252,N_205,N_812);
nand U1253 (N_1253,N_914,N_202);
and U1254 (N_1254,N_277,N_614);
nor U1255 (N_1255,N_482,N_648);
nand U1256 (N_1256,N_416,N_858);
nand U1257 (N_1257,N_843,N_709);
nand U1258 (N_1258,N_587,N_809);
or U1259 (N_1259,N_605,N_922);
and U1260 (N_1260,N_294,N_395);
nand U1261 (N_1261,N_7,N_197);
nand U1262 (N_1262,N_769,N_269);
nor U1263 (N_1263,N_638,N_467);
and U1264 (N_1264,N_477,N_559);
or U1265 (N_1265,N_20,N_819);
nand U1266 (N_1266,N_145,N_938);
and U1267 (N_1267,N_894,N_535);
or U1268 (N_1268,N_315,N_95);
nand U1269 (N_1269,N_944,N_678);
or U1270 (N_1270,N_27,N_23);
nor U1271 (N_1271,N_660,N_871);
or U1272 (N_1272,N_119,N_285);
or U1273 (N_1273,N_742,N_714);
nor U1274 (N_1274,N_383,N_739);
and U1275 (N_1275,N_414,N_390);
nor U1276 (N_1276,N_783,N_428);
and U1277 (N_1277,N_295,N_976);
and U1278 (N_1278,N_79,N_511);
nand U1279 (N_1279,N_51,N_327);
nand U1280 (N_1280,N_251,N_328);
nand U1281 (N_1281,N_986,N_530);
nand U1282 (N_1282,N_838,N_385);
nor U1283 (N_1283,N_92,N_238);
and U1284 (N_1284,N_36,N_381);
xor U1285 (N_1285,N_378,N_669);
and U1286 (N_1286,N_320,N_687);
xor U1287 (N_1287,N_326,N_456);
and U1288 (N_1288,N_613,N_778);
nor U1289 (N_1289,N_358,N_455);
and U1290 (N_1290,N_995,N_949);
or U1291 (N_1291,N_875,N_246);
or U1292 (N_1292,N_107,N_968);
nor U1293 (N_1293,N_529,N_932);
nor U1294 (N_1294,N_263,N_17);
nor U1295 (N_1295,N_396,N_874);
or U1296 (N_1296,N_888,N_329);
nor U1297 (N_1297,N_462,N_811);
xor U1298 (N_1298,N_790,N_997);
and U1299 (N_1299,N_399,N_768);
and U1300 (N_1300,N_992,N_190);
or U1301 (N_1301,N_889,N_636);
and U1302 (N_1302,N_859,N_692);
nor U1303 (N_1303,N_831,N_253);
nor U1304 (N_1304,N_13,N_994);
and U1305 (N_1305,N_451,N_305);
nand U1306 (N_1306,N_953,N_434);
and U1307 (N_1307,N_920,N_904);
nand U1308 (N_1308,N_497,N_255);
xnor U1309 (N_1309,N_299,N_782);
or U1310 (N_1310,N_53,N_698);
xor U1311 (N_1311,N_433,N_412);
or U1312 (N_1312,N_984,N_776);
or U1313 (N_1313,N_818,N_247);
nand U1314 (N_1314,N_100,N_317);
or U1315 (N_1315,N_55,N_387);
nor U1316 (N_1316,N_907,N_899);
and U1317 (N_1317,N_463,N_349);
or U1318 (N_1318,N_309,N_346);
and U1319 (N_1319,N_531,N_206);
or U1320 (N_1320,N_764,N_461);
nor U1321 (N_1321,N_746,N_60);
or U1322 (N_1322,N_760,N_807);
or U1323 (N_1323,N_394,N_243);
or U1324 (N_1324,N_52,N_439);
nor U1325 (N_1325,N_454,N_260);
and U1326 (N_1326,N_925,N_367);
or U1327 (N_1327,N_789,N_921);
and U1328 (N_1328,N_924,N_557);
nor U1329 (N_1329,N_403,N_227);
and U1330 (N_1330,N_167,N_982);
xnor U1331 (N_1331,N_836,N_730);
or U1332 (N_1332,N_402,N_852);
and U1333 (N_1333,N_516,N_721);
nor U1334 (N_1334,N_877,N_651);
and U1335 (N_1335,N_298,N_57);
xor U1336 (N_1336,N_734,N_222);
xor U1337 (N_1337,N_74,N_115);
nand U1338 (N_1338,N_121,N_14);
nor U1339 (N_1339,N_331,N_785);
or U1340 (N_1340,N_603,N_592);
or U1341 (N_1341,N_47,N_480);
or U1342 (N_1342,N_301,N_26);
nor U1343 (N_1343,N_124,N_262);
and U1344 (N_1344,N_311,N_780);
and U1345 (N_1345,N_897,N_69);
and U1346 (N_1346,N_668,N_735);
or U1347 (N_1347,N_70,N_303);
and U1348 (N_1348,N_578,N_226);
nor U1349 (N_1349,N_99,N_418);
nand U1350 (N_1350,N_918,N_256);
or U1351 (N_1351,N_495,N_419);
and U1352 (N_1352,N_558,N_941);
or U1353 (N_1353,N_103,N_909);
or U1354 (N_1354,N_634,N_770);
nand U1355 (N_1355,N_837,N_376);
and U1356 (N_1356,N_554,N_96);
nor U1357 (N_1357,N_272,N_695);
and U1358 (N_1358,N_200,N_718);
nand U1359 (N_1359,N_872,N_560);
nand U1360 (N_1360,N_963,N_707);
nor U1361 (N_1361,N_471,N_12);
nand U1362 (N_1362,N_917,N_168);
xor U1363 (N_1363,N_91,N_689);
or U1364 (N_1364,N_34,N_693);
and U1365 (N_1365,N_664,N_677);
xnor U1366 (N_1366,N_165,N_977);
nor U1367 (N_1367,N_788,N_891);
nor U1368 (N_1368,N_791,N_58);
nand U1369 (N_1369,N_644,N_169);
nor U1370 (N_1370,N_221,N_449);
or U1371 (N_1371,N_308,N_278);
or U1372 (N_1372,N_499,N_641);
xnor U1373 (N_1373,N_164,N_393);
nand U1374 (N_1374,N_4,N_796);
nor U1375 (N_1375,N_140,N_87);
or U1376 (N_1376,N_849,N_80);
nand U1377 (N_1377,N_936,N_193);
and U1378 (N_1378,N_777,N_489);
nand U1379 (N_1379,N_743,N_204);
nand U1380 (N_1380,N_347,N_928);
or U1381 (N_1381,N_16,N_279);
and U1382 (N_1382,N_470,N_446);
nand U1383 (N_1383,N_971,N_970);
nor U1384 (N_1384,N_545,N_611);
or U1385 (N_1385,N_504,N_423);
xor U1386 (N_1386,N_561,N_288);
xnor U1387 (N_1387,N_575,N_632);
or U1388 (N_1388,N_753,N_421);
nor U1389 (N_1389,N_887,N_189);
nand U1390 (N_1390,N_608,N_784);
or U1391 (N_1391,N_950,N_842);
nor U1392 (N_1392,N_667,N_105);
or U1393 (N_1393,N_502,N_166);
or U1394 (N_1394,N_382,N_823);
nand U1395 (N_1395,N_370,N_594);
or U1396 (N_1396,N_710,N_729);
or U1397 (N_1397,N_137,N_196);
or U1398 (N_1398,N_220,N_759);
nand U1399 (N_1399,N_583,N_635);
nand U1400 (N_1400,N_824,N_313);
nor U1401 (N_1401,N_425,N_448);
nand U1402 (N_1402,N_420,N_772);
nand U1403 (N_1403,N_755,N_171);
or U1404 (N_1404,N_65,N_805);
nor U1405 (N_1405,N_436,N_895);
or U1406 (N_1406,N_652,N_898);
nor U1407 (N_1407,N_850,N_911);
or U1408 (N_1408,N_62,N_321);
nand U1409 (N_1409,N_142,N_483);
or U1410 (N_1410,N_174,N_865);
or U1411 (N_1411,N_472,N_879);
or U1412 (N_1412,N_473,N_35);
xnor U1413 (N_1413,N_750,N_533);
nand U1414 (N_1414,N_881,N_413);
or U1415 (N_1415,N_30,N_878);
and U1416 (N_1416,N_612,N_983);
or U1417 (N_1417,N_745,N_94);
nor U1418 (N_1418,N_179,N_943);
nor U1419 (N_1419,N_565,N_866);
or U1420 (N_1420,N_757,N_799);
and U1421 (N_1421,N_598,N_281);
xor U1422 (N_1422,N_514,N_569);
nor U1423 (N_1423,N_271,N_826);
and U1424 (N_1424,N_134,N_752);
nand U1425 (N_1425,N_923,N_216);
nor U1426 (N_1426,N_589,N_437);
nand U1427 (N_1427,N_237,N_469);
nor U1428 (N_1428,N_217,N_700);
nor U1429 (N_1429,N_675,N_153);
nor U1430 (N_1430,N_355,N_679);
nor U1431 (N_1431,N_56,N_212);
nand U1432 (N_1432,N_210,N_998);
and U1433 (N_1433,N_846,N_890);
and U1434 (N_1434,N_500,N_487);
or U1435 (N_1435,N_703,N_322);
xnor U1436 (N_1436,N_33,N_580);
nand U1437 (N_1437,N_223,N_476);
nand U1438 (N_1438,N_913,N_616);
and U1439 (N_1439,N_681,N_215);
nor U1440 (N_1440,N_63,N_848);
nor U1441 (N_1441,N_78,N_989);
nor U1442 (N_1442,N_273,N_975);
nor U1443 (N_1443,N_108,N_139);
nor U1444 (N_1444,N_816,N_481);
or U1445 (N_1445,N_146,N_854);
nor U1446 (N_1446,N_773,N_527);
or U1447 (N_1447,N_175,N_863);
nand U1448 (N_1448,N_147,N_261);
nand U1449 (N_1449,N_316,N_775);
or U1450 (N_1450,N_629,N_806);
xor U1451 (N_1451,N_510,N_280);
and U1452 (N_1452,N_902,N_219);
and U1453 (N_1453,N_708,N_671);
nor U1454 (N_1454,N_981,N_214);
or U1455 (N_1455,N_952,N_618);
nand U1456 (N_1456,N_252,N_539);
nand U1457 (N_1457,N_188,N_149);
nand U1458 (N_1458,N_733,N_857);
and U1459 (N_1459,N_292,N_892);
or U1460 (N_1460,N_312,N_749);
or U1461 (N_1461,N_494,N_38);
nand U1462 (N_1462,N_41,N_711);
nand U1463 (N_1463,N_630,N_398);
nand U1464 (N_1464,N_319,N_604);
and U1465 (N_1465,N_81,N_751);
xor U1466 (N_1466,N_570,N_259);
and U1467 (N_1467,N_485,N_713);
or U1468 (N_1468,N_650,N_701);
nand U1469 (N_1469,N_988,N_180);
nor U1470 (N_1470,N_912,N_815);
and U1471 (N_1471,N_444,N_544);
or U1472 (N_1472,N_345,N_568);
xnor U1473 (N_1473,N_49,N_794);
xor U1474 (N_1474,N_457,N_547);
nor U1475 (N_1475,N_702,N_11);
and U1476 (N_1476,N_946,N_232);
and U1477 (N_1477,N_447,N_624);
or U1478 (N_1478,N_723,N_736);
xnor U1479 (N_1479,N_717,N_380);
or U1480 (N_1480,N_182,N_426);
nor U1481 (N_1481,N_955,N_781);
or U1482 (N_1482,N_406,N_491);
nand U1483 (N_1483,N_415,N_154);
or U1484 (N_1484,N_173,N_832);
nor U1485 (N_1485,N_869,N_553);
nand U1486 (N_1486,N_661,N_967);
and U1487 (N_1487,N_505,N_290);
xor U1488 (N_1488,N_993,N_972);
nand U1489 (N_1489,N_111,N_386);
nor U1490 (N_1490,N_551,N_969);
xnor U1491 (N_1491,N_340,N_64);
nor U1492 (N_1492,N_208,N_766);
and U1493 (N_1493,N_686,N_724);
xor U1494 (N_1494,N_19,N_961);
and U1495 (N_1495,N_330,N_947);
or U1496 (N_1496,N_254,N_117);
nand U1497 (N_1497,N_813,N_102);
nand U1498 (N_1498,N_732,N_44);
and U1499 (N_1499,N_933,N_503);
and U1500 (N_1500,N_843,N_533);
nor U1501 (N_1501,N_209,N_779);
nor U1502 (N_1502,N_283,N_338);
nor U1503 (N_1503,N_284,N_698);
nor U1504 (N_1504,N_827,N_402);
nor U1505 (N_1505,N_425,N_609);
or U1506 (N_1506,N_46,N_260);
or U1507 (N_1507,N_958,N_71);
xnor U1508 (N_1508,N_524,N_62);
nand U1509 (N_1509,N_81,N_748);
and U1510 (N_1510,N_593,N_761);
or U1511 (N_1511,N_447,N_944);
or U1512 (N_1512,N_225,N_77);
and U1513 (N_1513,N_163,N_326);
nor U1514 (N_1514,N_830,N_123);
or U1515 (N_1515,N_865,N_594);
nand U1516 (N_1516,N_832,N_80);
or U1517 (N_1517,N_279,N_889);
or U1518 (N_1518,N_798,N_362);
or U1519 (N_1519,N_947,N_257);
nand U1520 (N_1520,N_693,N_431);
or U1521 (N_1521,N_940,N_339);
nand U1522 (N_1522,N_873,N_417);
or U1523 (N_1523,N_733,N_496);
nand U1524 (N_1524,N_573,N_926);
or U1525 (N_1525,N_492,N_98);
xor U1526 (N_1526,N_541,N_131);
nor U1527 (N_1527,N_945,N_694);
nand U1528 (N_1528,N_419,N_822);
and U1529 (N_1529,N_468,N_447);
or U1530 (N_1530,N_889,N_389);
nor U1531 (N_1531,N_139,N_466);
xnor U1532 (N_1532,N_275,N_436);
nor U1533 (N_1533,N_274,N_403);
or U1534 (N_1534,N_833,N_296);
nor U1535 (N_1535,N_624,N_84);
or U1536 (N_1536,N_45,N_158);
nand U1537 (N_1537,N_414,N_682);
xnor U1538 (N_1538,N_963,N_748);
or U1539 (N_1539,N_880,N_563);
nand U1540 (N_1540,N_865,N_983);
nand U1541 (N_1541,N_391,N_507);
or U1542 (N_1542,N_378,N_492);
nor U1543 (N_1543,N_100,N_56);
or U1544 (N_1544,N_800,N_866);
or U1545 (N_1545,N_992,N_615);
nor U1546 (N_1546,N_661,N_574);
and U1547 (N_1547,N_725,N_155);
nor U1548 (N_1548,N_307,N_114);
or U1549 (N_1549,N_243,N_55);
nand U1550 (N_1550,N_886,N_557);
or U1551 (N_1551,N_951,N_689);
nor U1552 (N_1552,N_367,N_515);
and U1553 (N_1553,N_646,N_635);
and U1554 (N_1554,N_662,N_361);
xor U1555 (N_1555,N_687,N_13);
nand U1556 (N_1556,N_506,N_958);
or U1557 (N_1557,N_691,N_671);
nor U1558 (N_1558,N_662,N_499);
or U1559 (N_1559,N_352,N_941);
nor U1560 (N_1560,N_574,N_866);
and U1561 (N_1561,N_643,N_426);
nor U1562 (N_1562,N_284,N_869);
nand U1563 (N_1563,N_710,N_272);
xor U1564 (N_1564,N_201,N_401);
nand U1565 (N_1565,N_387,N_613);
nand U1566 (N_1566,N_713,N_124);
or U1567 (N_1567,N_719,N_39);
and U1568 (N_1568,N_34,N_23);
nor U1569 (N_1569,N_640,N_156);
nor U1570 (N_1570,N_420,N_183);
or U1571 (N_1571,N_208,N_402);
or U1572 (N_1572,N_699,N_737);
nand U1573 (N_1573,N_47,N_344);
nor U1574 (N_1574,N_212,N_23);
nand U1575 (N_1575,N_765,N_354);
and U1576 (N_1576,N_218,N_117);
and U1577 (N_1577,N_124,N_851);
or U1578 (N_1578,N_780,N_950);
nand U1579 (N_1579,N_288,N_752);
xnor U1580 (N_1580,N_866,N_516);
xnor U1581 (N_1581,N_18,N_824);
or U1582 (N_1582,N_226,N_557);
nand U1583 (N_1583,N_877,N_574);
or U1584 (N_1584,N_468,N_895);
nand U1585 (N_1585,N_507,N_107);
or U1586 (N_1586,N_942,N_998);
nand U1587 (N_1587,N_530,N_553);
xor U1588 (N_1588,N_453,N_649);
or U1589 (N_1589,N_412,N_180);
nand U1590 (N_1590,N_225,N_861);
nor U1591 (N_1591,N_133,N_638);
nand U1592 (N_1592,N_630,N_740);
or U1593 (N_1593,N_7,N_135);
and U1594 (N_1594,N_242,N_116);
nand U1595 (N_1595,N_261,N_279);
nor U1596 (N_1596,N_686,N_253);
and U1597 (N_1597,N_638,N_259);
nor U1598 (N_1598,N_460,N_425);
and U1599 (N_1599,N_598,N_219);
nand U1600 (N_1600,N_743,N_290);
or U1601 (N_1601,N_971,N_72);
and U1602 (N_1602,N_87,N_448);
or U1603 (N_1603,N_990,N_882);
and U1604 (N_1604,N_781,N_615);
and U1605 (N_1605,N_980,N_443);
and U1606 (N_1606,N_221,N_129);
xnor U1607 (N_1607,N_486,N_2);
nand U1608 (N_1608,N_159,N_234);
and U1609 (N_1609,N_816,N_769);
nor U1610 (N_1610,N_904,N_420);
and U1611 (N_1611,N_217,N_272);
nand U1612 (N_1612,N_683,N_788);
xnor U1613 (N_1613,N_976,N_21);
and U1614 (N_1614,N_198,N_959);
nor U1615 (N_1615,N_234,N_853);
or U1616 (N_1616,N_788,N_348);
and U1617 (N_1617,N_147,N_957);
and U1618 (N_1618,N_704,N_292);
or U1619 (N_1619,N_350,N_174);
nand U1620 (N_1620,N_277,N_622);
and U1621 (N_1621,N_266,N_9);
or U1622 (N_1622,N_23,N_315);
nor U1623 (N_1623,N_166,N_512);
or U1624 (N_1624,N_611,N_550);
and U1625 (N_1625,N_247,N_701);
xnor U1626 (N_1626,N_122,N_764);
and U1627 (N_1627,N_517,N_183);
nor U1628 (N_1628,N_281,N_413);
or U1629 (N_1629,N_614,N_256);
or U1630 (N_1630,N_67,N_448);
nand U1631 (N_1631,N_950,N_319);
nand U1632 (N_1632,N_286,N_881);
nand U1633 (N_1633,N_415,N_915);
nor U1634 (N_1634,N_355,N_537);
or U1635 (N_1635,N_872,N_202);
or U1636 (N_1636,N_221,N_136);
and U1637 (N_1637,N_76,N_849);
and U1638 (N_1638,N_415,N_518);
or U1639 (N_1639,N_45,N_227);
nor U1640 (N_1640,N_495,N_194);
nor U1641 (N_1641,N_754,N_409);
xnor U1642 (N_1642,N_343,N_348);
nand U1643 (N_1643,N_37,N_406);
nor U1644 (N_1644,N_439,N_851);
or U1645 (N_1645,N_681,N_255);
and U1646 (N_1646,N_451,N_660);
or U1647 (N_1647,N_899,N_541);
nor U1648 (N_1648,N_33,N_462);
nand U1649 (N_1649,N_162,N_60);
nand U1650 (N_1650,N_161,N_607);
or U1651 (N_1651,N_664,N_367);
nand U1652 (N_1652,N_608,N_633);
nor U1653 (N_1653,N_699,N_321);
and U1654 (N_1654,N_504,N_557);
nand U1655 (N_1655,N_557,N_778);
or U1656 (N_1656,N_352,N_78);
or U1657 (N_1657,N_738,N_966);
xor U1658 (N_1658,N_868,N_792);
nand U1659 (N_1659,N_15,N_233);
and U1660 (N_1660,N_727,N_790);
nand U1661 (N_1661,N_328,N_601);
nand U1662 (N_1662,N_424,N_432);
xnor U1663 (N_1663,N_443,N_21);
and U1664 (N_1664,N_894,N_331);
nor U1665 (N_1665,N_334,N_439);
nor U1666 (N_1666,N_886,N_239);
nor U1667 (N_1667,N_33,N_275);
nand U1668 (N_1668,N_59,N_331);
or U1669 (N_1669,N_42,N_493);
nor U1670 (N_1670,N_675,N_556);
nor U1671 (N_1671,N_971,N_987);
and U1672 (N_1672,N_270,N_209);
nand U1673 (N_1673,N_139,N_494);
nor U1674 (N_1674,N_285,N_497);
nor U1675 (N_1675,N_800,N_258);
and U1676 (N_1676,N_750,N_622);
or U1677 (N_1677,N_755,N_966);
nor U1678 (N_1678,N_114,N_385);
nand U1679 (N_1679,N_567,N_709);
or U1680 (N_1680,N_2,N_872);
and U1681 (N_1681,N_736,N_513);
nor U1682 (N_1682,N_210,N_99);
or U1683 (N_1683,N_449,N_547);
or U1684 (N_1684,N_572,N_617);
or U1685 (N_1685,N_439,N_198);
and U1686 (N_1686,N_409,N_595);
or U1687 (N_1687,N_441,N_800);
nand U1688 (N_1688,N_823,N_452);
nand U1689 (N_1689,N_845,N_345);
and U1690 (N_1690,N_602,N_645);
and U1691 (N_1691,N_613,N_820);
xor U1692 (N_1692,N_280,N_404);
or U1693 (N_1693,N_175,N_80);
nor U1694 (N_1694,N_616,N_682);
or U1695 (N_1695,N_164,N_399);
or U1696 (N_1696,N_708,N_818);
nor U1697 (N_1697,N_180,N_264);
or U1698 (N_1698,N_670,N_100);
and U1699 (N_1699,N_186,N_306);
or U1700 (N_1700,N_734,N_625);
nor U1701 (N_1701,N_475,N_18);
nor U1702 (N_1702,N_552,N_724);
and U1703 (N_1703,N_171,N_218);
nand U1704 (N_1704,N_638,N_16);
and U1705 (N_1705,N_325,N_359);
nand U1706 (N_1706,N_264,N_274);
or U1707 (N_1707,N_413,N_315);
and U1708 (N_1708,N_856,N_768);
or U1709 (N_1709,N_443,N_826);
and U1710 (N_1710,N_189,N_454);
or U1711 (N_1711,N_249,N_803);
nor U1712 (N_1712,N_740,N_320);
nand U1713 (N_1713,N_79,N_578);
and U1714 (N_1714,N_438,N_52);
and U1715 (N_1715,N_124,N_764);
and U1716 (N_1716,N_980,N_45);
and U1717 (N_1717,N_271,N_686);
xor U1718 (N_1718,N_969,N_123);
and U1719 (N_1719,N_905,N_656);
and U1720 (N_1720,N_939,N_58);
nand U1721 (N_1721,N_22,N_705);
nand U1722 (N_1722,N_208,N_83);
nand U1723 (N_1723,N_709,N_921);
nand U1724 (N_1724,N_146,N_787);
nor U1725 (N_1725,N_124,N_946);
nor U1726 (N_1726,N_771,N_314);
nand U1727 (N_1727,N_176,N_204);
or U1728 (N_1728,N_890,N_88);
xor U1729 (N_1729,N_939,N_200);
and U1730 (N_1730,N_678,N_330);
nor U1731 (N_1731,N_693,N_835);
nor U1732 (N_1732,N_775,N_42);
or U1733 (N_1733,N_974,N_958);
nor U1734 (N_1734,N_74,N_493);
nor U1735 (N_1735,N_901,N_435);
nor U1736 (N_1736,N_884,N_608);
nand U1737 (N_1737,N_246,N_313);
and U1738 (N_1738,N_483,N_997);
nand U1739 (N_1739,N_184,N_870);
nor U1740 (N_1740,N_572,N_760);
or U1741 (N_1741,N_561,N_36);
or U1742 (N_1742,N_458,N_141);
xnor U1743 (N_1743,N_270,N_909);
or U1744 (N_1744,N_401,N_470);
or U1745 (N_1745,N_932,N_869);
or U1746 (N_1746,N_596,N_700);
nor U1747 (N_1747,N_777,N_616);
nor U1748 (N_1748,N_84,N_570);
nand U1749 (N_1749,N_474,N_394);
nand U1750 (N_1750,N_330,N_53);
or U1751 (N_1751,N_38,N_215);
xor U1752 (N_1752,N_722,N_792);
and U1753 (N_1753,N_579,N_308);
and U1754 (N_1754,N_400,N_549);
xor U1755 (N_1755,N_929,N_671);
nor U1756 (N_1756,N_198,N_926);
and U1757 (N_1757,N_706,N_499);
xnor U1758 (N_1758,N_533,N_185);
or U1759 (N_1759,N_791,N_910);
xnor U1760 (N_1760,N_489,N_237);
and U1761 (N_1761,N_704,N_303);
nand U1762 (N_1762,N_577,N_691);
or U1763 (N_1763,N_788,N_489);
or U1764 (N_1764,N_927,N_602);
nor U1765 (N_1765,N_756,N_779);
nor U1766 (N_1766,N_72,N_862);
nand U1767 (N_1767,N_618,N_181);
and U1768 (N_1768,N_616,N_754);
or U1769 (N_1769,N_933,N_949);
nand U1770 (N_1770,N_440,N_892);
nand U1771 (N_1771,N_26,N_294);
xor U1772 (N_1772,N_927,N_963);
nor U1773 (N_1773,N_508,N_950);
nand U1774 (N_1774,N_606,N_634);
and U1775 (N_1775,N_555,N_956);
nand U1776 (N_1776,N_911,N_521);
and U1777 (N_1777,N_752,N_901);
nor U1778 (N_1778,N_536,N_695);
or U1779 (N_1779,N_437,N_674);
and U1780 (N_1780,N_989,N_578);
nor U1781 (N_1781,N_529,N_315);
nand U1782 (N_1782,N_609,N_731);
or U1783 (N_1783,N_228,N_925);
nand U1784 (N_1784,N_523,N_99);
nand U1785 (N_1785,N_101,N_974);
and U1786 (N_1786,N_25,N_137);
nor U1787 (N_1787,N_517,N_64);
nand U1788 (N_1788,N_188,N_182);
or U1789 (N_1789,N_672,N_127);
or U1790 (N_1790,N_380,N_650);
nor U1791 (N_1791,N_362,N_245);
nand U1792 (N_1792,N_254,N_804);
and U1793 (N_1793,N_762,N_652);
and U1794 (N_1794,N_873,N_186);
and U1795 (N_1795,N_670,N_3);
and U1796 (N_1796,N_365,N_273);
or U1797 (N_1797,N_671,N_365);
and U1798 (N_1798,N_697,N_116);
nand U1799 (N_1799,N_974,N_532);
nor U1800 (N_1800,N_938,N_49);
and U1801 (N_1801,N_575,N_303);
xor U1802 (N_1802,N_171,N_709);
nor U1803 (N_1803,N_547,N_706);
and U1804 (N_1804,N_370,N_436);
and U1805 (N_1805,N_638,N_613);
nand U1806 (N_1806,N_930,N_968);
xnor U1807 (N_1807,N_786,N_894);
or U1808 (N_1808,N_454,N_963);
or U1809 (N_1809,N_408,N_507);
nor U1810 (N_1810,N_410,N_937);
or U1811 (N_1811,N_868,N_914);
nand U1812 (N_1812,N_257,N_299);
nor U1813 (N_1813,N_561,N_573);
or U1814 (N_1814,N_310,N_841);
nand U1815 (N_1815,N_575,N_29);
and U1816 (N_1816,N_585,N_349);
or U1817 (N_1817,N_33,N_421);
or U1818 (N_1818,N_242,N_249);
and U1819 (N_1819,N_388,N_571);
or U1820 (N_1820,N_386,N_874);
or U1821 (N_1821,N_886,N_667);
nor U1822 (N_1822,N_804,N_26);
nor U1823 (N_1823,N_401,N_755);
and U1824 (N_1824,N_74,N_661);
nand U1825 (N_1825,N_187,N_594);
nand U1826 (N_1826,N_582,N_543);
nand U1827 (N_1827,N_513,N_142);
nor U1828 (N_1828,N_909,N_746);
or U1829 (N_1829,N_516,N_84);
or U1830 (N_1830,N_186,N_203);
xor U1831 (N_1831,N_890,N_52);
nor U1832 (N_1832,N_961,N_363);
and U1833 (N_1833,N_882,N_699);
and U1834 (N_1834,N_686,N_734);
xor U1835 (N_1835,N_69,N_651);
or U1836 (N_1836,N_889,N_338);
and U1837 (N_1837,N_451,N_590);
and U1838 (N_1838,N_245,N_846);
or U1839 (N_1839,N_560,N_33);
and U1840 (N_1840,N_511,N_88);
nand U1841 (N_1841,N_41,N_131);
or U1842 (N_1842,N_523,N_992);
and U1843 (N_1843,N_886,N_104);
and U1844 (N_1844,N_69,N_622);
nand U1845 (N_1845,N_231,N_594);
nand U1846 (N_1846,N_406,N_815);
nor U1847 (N_1847,N_820,N_770);
or U1848 (N_1848,N_823,N_920);
nor U1849 (N_1849,N_158,N_920);
xor U1850 (N_1850,N_760,N_368);
nor U1851 (N_1851,N_517,N_584);
nand U1852 (N_1852,N_510,N_562);
and U1853 (N_1853,N_323,N_117);
and U1854 (N_1854,N_413,N_14);
and U1855 (N_1855,N_621,N_24);
nor U1856 (N_1856,N_502,N_945);
and U1857 (N_1857,N_563,N_862);
nor U1858 (N_1858,N_262,N_205);
or U1859 (N_1859,N_42,N_851);
and U1860 (N_1860,N_454,N_776);
nand U1861 (N_1861,N_636,N_705);
xnor U1862 (N_1862,N_371,N_281);
or U1863 (N_1863,N_912,N_333);
nand U1864 (N_1864,N_709,N_527);
and U1865 (N_1865,N_976,N_766);
or U1866 (N_1866,N_695,N_247);
and U1867 (N_1867,N_767,N_714);
and U1868 (N_1868,N_312,N_213);
or U1869 (N_1869,N_296,N_809);
or U1870 (N_1870,N_460,N_220);
and U1871 (N_1871,N_598,N_804);
nor U1872 (N_1872,N_202,N_624);
or U1873 (N_1873,N_464,N_821);
or U1874 (N_1874,N_49,N_778);
or U1875 (N_1875,N_260,N_122);
nand U1876 (N_1876,N_824,N_133);
or U1877 (N_1877,N_303,N_623);
and U1878 (N_1878,N_680,N_971);
and U1879 (N_1879,N_751,N_54);
and U1880 (N_1880,N_21,N_484);
nand U1881 (N_1881,N_88,N_365);
or U1882 (N_1882,N_920,N_865);
or U1883 (N_1883,N_1,N_510);
nand U1884 (N_1884,N_442,N_864);
nand U1885 (N_1885,N_376,N_75);
or U1886 (N_1886,N_333,N_452);
nor U1887 (N_1887,N_500,N_95);
nor U1888 (N_1888,N_661,N_723);
or U1889 (N_1889,N_983,N_470);
xnor U1890 (N_1890,N_17,N_303);
or U1891 (N_1891,N_905,N_685);
and U1892 (N_1892,N_173,N_478);
nand U1893 (N_1893,N_715,N_584);
nor U1894 (N_1894,N_425,N_389);
and U1895 (N_1895,N_959,N_166);
and U1896 (N_1896,N_571,N_692);
nor U1897 (N_1897,N_830,N_348);
and U1898 (N_1898,N_885,N_966);
and U1899 (N_1899,N_78,N_854);
nand U1900 (N_1900,N_244,N_734);
or U1901 (N_1901,N_63,N_218);
and U1902 (N_1902,N_562,N_123);
xor U1903 (N_1903,N_561,N_53);
nand U1904 (N_1904,N_822,N_845);
nand U1905 (N_1905,N_794,N_565);
or U1906 (N_1906,N_701,N_193);
xnor U1907 (N_1907,N_783,N_518);
nor U1908 (N_1908,N_792,N_137);
or U1909 (N_1909,N_937,N_175);
or U1910 (N_1910,N_771,N_32);
or U1911 (N_1911,N_99,N_656);
nand U1912 (N_1912,N_903,N_152);
xnor U1913 (N_1913,N_978,N_629);
nor U1914 (N_1914,N_664,N_699);
nand U1915 (N_1915,N_671,N_161);
nor U1916 (N_1916,N_336,N_206);
nor U1917 (N_1917,N_226,N_786);
or U1918 (N_1918,N_47,N_598);
nand U1919 (N_1919,N_716,N_117);
nor U1920 (N_1920,N_256,N_125);
nor U1921 (N_1921,N_208,N_77);
nor U1922 (N_1922,N_131,N_642);
nor U1923 (N_1923,N_804,N_504);
nor U1924 (N_1924,N_314,N_20);
and U1925 (N_1925,N_588,N_695);
nand U1926 (N_1926,N_878,N_453);
and U1927 (N_1927,N_727,N_411);
and U1928 (N_1928,N_552,N_986);
or U1929 (N_1929,N_770,N_920);
nand U1930 (N_1930,N_329,N_643);
nor U1931 (N_1931,N_290,N_418);
and U1932 (N_1932,N_479,N_33);
or U1933 (N_1933,N_68,N_410);
nand U1934 (N_1934,N_12,N_285);
nand U1935 (N_1935,N_723,N_431);
and U1936 (N_1936,N_390,N_260);
and U1937 (N_1937,N_805,N_927);
xor U1938 (N_1938,N_289,N_993);
xnor U1939 (N_1939,N_152,N_519);
and U1940 (N_1940,N_521,N_387);
nand U1941 (N_1941,N_302,N_150);
and U1942 (N_1942,N_498,N_380);
and U1943 (N_1943,N_346,N_539);
nand U1944 (N_1944,N_289,N_839);
xor U1945 (N_1945,N_455,N_474);
or U1946 (N_1946,N_388,N_397);
and U1947 (N_1947,N_696,N_971);
nor U1948 (N_1948,N_240,N_162);
or U1949 (N_1949,N_433,N_460);
nand U1950 (N_1950,N_723,N_847);
or U1951 (N_1951,N_922,N_81);
nand U1952 (N_1952,N_847,N_138);
nor U1953 (N_1953,N_624,N_933);
or U1954 (N_1954,N_38,N_564);
nor U1955 (N_1955,N_532,N_37);
or U1956 (N_1956,N_898,N_273);
or U1957 (N_1957,N_274,N_432);
and U1958 (N_1958,N_208,N_654);
xnor U1959 (N_1959,N_442,N_238);
nand U1960 (N_1960,N_703,N_529);
and U1961 (N_1961,N_107,N_224);
nand U1962 (N_1962,N_184,N_931);
or U1963 (N_1963,N_477,N_901);
nor U1964 (N_1964,N_523,N_980);
and U1965 (N_1965,N_450,N_59);
xnor U1966 (N_1966,N_392,N_710);
and U1967 (N_1967,N_449,N_459);
or U1968 (N_1968,N_542,N_453);
nand U1969 (N_1969,N_659,N_586);
nand U1970 (N_1970,N_757,N_481);
and U1971 (N_1971,N_316,N_327);
xnor U1972 (N_1972,N_720,N_974);
or U1973 (N_1973,N_3,N_615);
or U1974 (N_1974,N_320,N_688);
nand U1975 (N_1975,N_627,N_377);
or U1976 (N_1976,N_642,N_484);
and U1977 (N_1977,N_797,N_894);
or U1978 (N_1978,N_458,N_853);
nor U1979 (N_1979,N_534,N_689);
or U1980 (N_1980,N_8,N_570);
nor U1981 (N_1981,N_797,N_565);
xnor U1982 (N_1982,N_986,N_298);
nor U1983 (N_1983,N_239,N_187);
and U1984 (N_1984,N_747,N_751);
and U1985 (N_1985,N_493,N_611);
or U1986 (N_1986,N_730,N_865);
nand U1987 (N_1987,N_970,N_739);
nor U1988 (N_1988,N_520,N_718);
or U1989 (N_1989,N_74,N_949);
or U1990 (N_1990,N_701,N_407);
or U1991 (N_1991,N_945,N_946);
xnor U1992 (N_1992,N_67,N_369);
nand U1993 (N_1993,N_922,N_917);
or U1994 (N_1994,N_409,N_69);
xor U1995 (N_1995,N_279,N_792);
and U1996 (N_1996,N_626,N_313);
nand U1997 (N_1997,N_668,N_430);
and U1998 (N_1998,N_655,N_24);
nand U1999 (N_1999,N_229,N_185);
and U2000 (N_2000,N_1509,N_1660);
nand U2001 (N_2001,N_1214,N_1555);
nor U2002 (N_2002,N_1175,N_1767);
or U2003 (N_2003,N_1096,N_1512);
nand U2004 (N_2004,N_1469,N_1124);
or U2005 (N_2005,N_1447,N_1674);
nand U2006 (N_2006,N_1987,N_1520);
nor U2007 (N_2007,N_1200,N_1911);
xnor U2008 (N_2008,N_1877,N_1100);
and U2009 (N_2009,N_1717,N_1189);
and U2010 (N_2010,N_1890,N_1082);
or U2011 (N_2011,N_1632,N_1549);
nor U2012 (N_2012,N_1445,N_1369);
nand U2013 (N_2013,N_1396,N_1402);
and U2014 (N_2014,N_1944,N_1915);
nor U2015 (N_2015,N_1841,N_1386);
nand U2016 (N_2016,N_1623,N_1655);
nor U2017 (N_2017,N_1011,N_1727);
nor U2018 (N_2018,N_1442,N_1681);
nand U2019 (N_2019,N_1471,N_1785);
xnor U2020 (N_2020,N_1460,N_1163);
nor U2021 (N_2021,N_1181,N_1507);
or U2022 (N_2022,N_1137,N_1734);
or U2023 (N_2023,N_1159,N_1070);
or U2024 (N_2024,N_1346,N_1553);
xor U2025 (N_2025,N_1358,N_1310);
nor U2026 (N_2026,N_1052,N_1781);
nor U2027 (N_2027,N_1943,N_1076);
or U2028 (N_2028,N_1038,N_1769);
nand U2029 (N_2029,N_1609,N_1107);
nor U2030 (N_2030,N_1487,N_1179);
nor U2031 (N_2031,N_1319,N_1295);
or U2032 (N_2032,N_1882,N_1385);
nor U2033 (N_2033,N_1021,N_1782);
nand U2034 (N_2034,N_1049,N_1145);
and U2035 (N_2035,N_1451,N_1851);
nor U2036 (N_2036,N_1739,N_1662);
or U2037 (N_2037,N_1019,N_1054);
nand U2038 (N_2038,N_1653,N_1042);
or U2039 (N_2039,N_1870,N_1673);
xnor U2040 (N_2040,N_1933,N_1462);
or U2041 (N_2041,N_1260,N_1459);
nand U2042 (N_2042,N_1716,N_1786);
nand U2043 (N_2043,N_1363,N_1097);
nor U2044 (N_2044,N_1060,N_1790);
or U2045 (N_2045,N_1055,N_1118);
and U2046 (N_2046,N_1357,N_1616);
or U2047 (N_2047,N_1232,N_1416);
xnor U2048 (N_2048,N_1449,N_1431);
and U2049 (N_2049,N_1132,N_1694);
or U2050 (N_2050,N_1267,N_1773);
nand U2051 (N_2051,N_1069,N_1527);
nand U2052 (N_2052,N_1412,N_1677);
and U2053 (N_2053,N_1091,N_1665);
nand U2054 (N_2054,N_1253,N_1929);
nand U2055 (N_2055,N_1153,N_1765);
nor U2056 (N_2056,N_1088,N_1280);
nor U2057 (N_2057,N_1948,N_1918);
nor U2058 (N_2058,N_1838,N_1365);
or U2059 (N_2059,N_1501,N_1524);
or U2060 (N_2060,N_1411,N_1032);
and U2061 (N_2061,N_1025,N_1580);
and U2062 (N_2062,N_1457,N_1754);
and U2063 (N_2063,N_1992,N_1635);
nor U2064 (N_2064,N_1218,N_1984);
and U2065 (N_2065,N_1066,N_1202);
or U2066 (N_2066,N_1466,N_1233);
or U2067 (N_2067,N_1401,N_1531);
nor U2068 (N_2068,N_1141,N_1843);
and U2069 (N_2069,N_1017,N_1381);
nand U2070 (N_2070,N_1348,N_1906);
or U2071 (N_2071,N_1404,N_1693);
nand U2072 (N_2072,N_1294,N_1910);
nor U2073 (N_2073,N_1110,N_1108);
nand U2074 (N_2074,N_1419,N_1802);
nor U2075 (N_2075,N_1994,N_1043);
and U2076 (N_2076,N_1610,N_1711);
nor U2077 (N_2077,N_1083,N_1747);
nand U2078 (N_2078,N_1429,N_1696);
nand U2079 (N_2079,N_1266,N_1085);
nand U2080 (N_2080,N_1259,N_1892);
nand U2081 (N_2081,N_1756,N_1536);
nand U2082 (N_2082,N_1488,N_1559);
nand U2083 (N_2083,N_1190,N_1116);
or U2084 (N_2084,N_1977,N_1736);
and U2085 (N_2085,N_1165,N_1483);
and U2086 (N_2086,N_1275,N_1226);
and U2087 (N_2087,N_1196,N_1169);
xor U2088 (N_2088,N_1583,N_1669);
nor U2089 (N_2089,N_1486,N_1206);
and U2090 (N_2090,N_1584,N_1596);
or U2091 (N_2091,N_1235,N_1406);
and U2092 (N_2092,N_1277,N_1286);
or U2093 (N_2093,N_1270,N_1177);
or U2094 (N_2094,N_1861,N_1230);
nand U2095 (N_2095,N_1819,N_1515);
and U2096 (N_2096,N_1063,N_1407);
nand U2097 (N_2097,N_1285,N_1245);
nand U2098 (N_2098,N_1899,N_1103);
and U2099 (N_2099,N_1808,N_1680);
or U2100 (N_2100,N_1287,N_1452);
nor U2101 (N_2101,N_1300,N_1258);
and U2102 (N_2102,N_1059,N_1338);
nand U2103 (N_2103,N_1908,N_1852);
and U2104 (N_2104,N_1354,N_1624);
nand U2105 (N_2105,N_1031,N_1119);
nand U2106 (N_2106,N_1435,N_1678);
nand U2107 (N_2107,N_1965,N_1951);
and U2108 (N_2108,N_1384,N_1039);
or U2109 (N_2109,N_1611,N_1254);
or U2110 (N_2110,N_1224,N_1133);
and U2111 (N_2111,N_1242,N_1622);
or U2112 (N_2112,N_1090,N_1774);
nand U2113 (N_2113,N_1383,N_1127);
nor U2114 (N_2114,N_1698,N_1544);
and U2115 (N_2115,N_1697,N_1548);
or U2116 (N_2116,N_1692,N_1249);
nor U2117 (N_2117,N_1092,N_1575);
and U2118 (N_2118,N_1539,N_1814);
and U2119 (N_2119,N_1432,N_1250);
and U2120 (N_2120,N_1582,N_1709);
nor U2121 (N_2121,N_1737,N_1247);
nor U2122 (N_2122,N_1081,N_1554);
nor U2123 (N_2123,N_1523,N_1301);
and U2124 (N_2124,N_1942,N_1872);
nor U2125 (N_2125,N_1009,N_1078);
xnor U2126 (N_2126,N_1847,N_1829);
or U2127 (N_2127,N_1491,N_1903);
nor U2128 (N_2128,N_1298,N_1262);
nor U2129 (N_2129,N_1657,N_1323);
or U2130 (N_2130,N_1506,N_1950);
or U2131 (N_2131,N_1308,N_1114);
nor U2132 (N_2132,N_1125,N_1561);
nand U2133 (N_2133,N_1970,N_1647);
nor U2134 (N_2134,N_1203,N_1683);
xnor U2135 (N_2135,N_1281,N_1307);
and U2136 (N_2136,N_1591,N_1891);
and U2137 (N_2137,N_1728,N_1732);
nor U2138 (N_2138,N_1517,N_1000);
nand U2139 (N_2139,N_1427,N_1322);
and U2140 (N_2140,N_1760,N_1989);
nand U2141 (N_2141,N_1729,N_1593);
xor U2142 (N_2142,N_1008,N_1126);
nand U2143 (N_2143,N_1198,N_1186);
and U2144 (N_2144,N_1188,N_1516);
and U2145 (N_2145,N_1712,N_1390);
nor U2146 (N_2146,N_1542,N_1775);
or U2147 (N_2147,N_1547,N_1821);
or U2148 (N_2148,N_1689,N_1661);
or U2149 (N_2149,N_1271,N_1364);
nor U2150 (N_2150,N_1012,N_1430);
or U2151 (N_2151,N_1378,N_1941);
xnor U2152 (N_2152,N_1156,N_1686);
nor U2153 (N_2153,N_1735,N_1800);
nand U2154 (N_2154,N_1113,N_1441);
and U2155 (N_2155,N_1414,N_1428);
or U2156 (N_2156,N_1492,N_1663);
or U2157 (N_2157,N_1576,N_1848);
or U2158 (N_2158,N_1439,N_1876);
xnor U2159 (N_2159,N_1030,N_1335);
or U2160 (N_2160,N_1556,N_1106);
and U2161 (N_2161,N_1465,N_1444);
or U2162 (N_2162,N_1914,N_1666);
xor U2163 (N_2163,N_1093,N_1649);
or U2164 (N_2164,N_1508,N_1146);
nand U2165 (N_2165,N_1753,N_1574);
nor U2166 (N_2166,N_1636,N_1894);
and U2167 (N_2167,N_1981,N_1881);
nand U2168 (N_2168,N_1751,N_1014);
nand U2169 (N_2169,N_1601,N_1990);
and U2170 (N_2170,N_1150,N_1016);
or U2171 (N_2171,N_1888,N_1764);
nand U2172 (N_2172,N_1541,N_1996);
nor U2173 (N_2173,N_1702,N_1023);
nor U2174 (N_2174,N_1968,N_1426);
xnor U2175 (N_2175,N_1388,N_1740);
xnor U2176 (N_2176,N_1902,N_1268);
or U2177 (N_2177,N_1708,N_1967);
nand U2178 (N_2178,N_1780,N_1244);
nand U2179 (N_2179,N_1885,N_1846);
nand U2180 (N_2180,N_1413,N_1679);
nor U2181 (N_2181,N_1174,N_1639);
and U2182 (N_2182,N_1777,N_1309);
or U2183 (N_2183,N_1535,N_1382);
nand U2184 (N_2184,N_1399,N_1707);
or U2185 (N_2185,N_1652,N_1671);
nand U2186 (N_2186,N_1067,N_1999);
or U2187 (N_2187,N_1068,N_1672);
and U2188 (N_2188,N_1900,N_1571);
and U2189 (N_2189,N_1033,N_1916);
or U2190 (N_2190,N_1592,N_1425);
xor U2191 (N_2191,N_1420,N_1607);
nand U2192 (N_2192,N_1873,N_1857);
xor U2193 (N_2193,N_1131,N_1834);
or U2194 (N_2194,N_1468,N_1788);
nand U2195 (N_2195,N_1599,N_1184);
and U2196 (N_2196,N_1077,N_1952);
nor U2197 (N_2197,N_1567,N_1484);
and U2198 (N_2198,N_1955,N_1518);
nor U2199 (N_2199,N_1745,N_1018);
or U2200 (N_2200,N_1868,N_1884);
nand U2201 (N_2201,N_1072,N_1171);
or U2202 (N_2202,N_1489,N_1495);
nor U2203 (N_2203,N_1194,N_1577);
or U2204 (N_2204,N_1947,N_1646);
nor U2205 (N_2205,N_1878,N_1682);
or U2206 (N_2206,N_1585,N_1654);
nor U2207 (N_2207,N_1762,N_1757);
or U2208 (N_2208,N_1606,N_1409);
or U2209 (N_2209,N_1638,N_1637);
nand U2210 (N_2210,N_1087,N_1629);
xor U2211 (N_2211,N_1768,N_1974);
nand U2212 (N_2212,N_1748,N_1372);
and U2213 (N_2213,N_1143,N_1115);
nor U2214 (N_2214,N_1565,N_1453);
xnor U2215 (N_2215,N_1170,N_1454);
nand U2216 (N_2216,N_1213,N_1853);
nor U2217 (N_2217,N_1744,N_1350);
nand U2218 (N_2218,N_1650,N_1225);
nor U2219 (N_2219,N_1215,N_1809);
or U2220 (N_2220,N_1122,N_1496);
nor U2221 (N_2221,N_1532,N_1216);
nand U2222 (N_2222,N_1315,N_1079);
or U2223 (N_2223,N_1210,N_1252);
or U2224 (N_2224,N_1807,N_1540);
and U2225 (N_2225,N_1563,N_1320);
nand U2226 (N_2226,N_1423,N_1776);
and U2227 (N_2227,N_1208,N_1010);
nand U2228 (N_2228,N_1928,N_1062);
or U2229 (N_2229,N_1341,N_1395);
and U2230 (N_2230,N_1475,N_1109);
and U2231 (N_2231,N_1699,N_1161);
nand U2232 (N_2232,N_1560,N_1869);
nand U2233 (N_2233,N_1424,N_1328);
and U2234 (N_2234,N_1939,N_1600);
nor U2235 (N_2235,N_1504,N_1791);
and U2236 (N_2236,N_1314,N_1719);
xor U2237 (N_2237,N_1236,N_1913);
and U2238 (N_2238,N_1241,N_1581);
xnor U2239 (N_2239,N_1823,N_1332);
nand U2240 (N_2240,N_1936,N_1704);
nand U2241 (N_2241,N_1839,N_1810);
nor U2242 (N_2242,N_1725,N_1771);
nor U2243 (N_2243,N_1227,N_1366);
and U2244 (N_2244,N_1796,N_1620);
or U2245 (N_2245,N_1211,N_1151);
and U2246 (N_2246,N_1687,N_1015);
and U2247 (N_2247,N_1927,N_1050);
or U2248 (N_2248,N_1960,N_1340);
and U2249 (N_2249,N_1130,N_1988);
and U2250 (N_2250,N_1361,N_1789);
nor U2251 (N_2251,N_1074,N_1209);
or U2252 (N_2252,N_1080,N_1587);
or U2253 (N_2253,N_1962,N_1825);
and U2254 (N_2254,N_1051,N_1237);
and U2255 (N_2255,N_1871,N_1343);
nand U2256 (N_2256,N_1590,N_1752);
nor U2257 (N_2257,N_1755,N_1598);
and U2258 (N_2258,N_1034,N_1812);
nand U2259 (N_2259,N_1956,N_1982);
or U2260 (N_2260,N_1519,N_1205);
nand U2261 (N_2261,N_1316,N_1648);
and U2262 (N_2262,N_1979,N_1045);
or U2263 (N_2263,N_1562,N_1797);
and U2264 (N_2264,N_1440,N_1889);
or U2265 (N_2265,N_1530,N_1502);
nor U2266 (N_2266,N_1588,N_1863);
or U2267 (N_2267,N_1879,N_1766);
nor U2268 (N_2268,N_1154,N_1614);
nand U2269 (N_2269,N_1811,N_1972);
or U2270 (N_2270,N_1883,N_1273);
nand U2271 (N_2271,N_1220,N_1026);
or U2272 (N_2272,N_1905,N_1993);
xnor U2273 (N_2273,N_1733,N_1880);
and U2274 (N_2274,N_1302,N_1710);
nor U2275 (N_2275,N_1522,N_1656);
and U2276 (N_2276,N_1276,N_1701);
nand U2277 (N_2277,N_1640,N_1830);
xor U2278 (N_2278,N_1526,N_1120);
and U2279 (N_2279,N_1408,N_1634);
nand U2280 (N_2280,N_1603,N_1255);
nor U2281 (N_2281,N_1136,N_1456);
or U2282 (N_2282,N_1594,N_1498);
nor U2283 (N_2283,N_1257,N_1299);
xor U2284 (N_2284,N_1325,N_1924);
nand U2285 (N_2285,N_1605,N_1651);
and U2286 (N_2286,N_1415,N_1391);
and U2287 (N_2287,N_1180,N_1071);
nand U2288 (N_2288,N_1166,N_1667);
or U2289 (N_2289,N_1670,N_1703);
nor U2290 (N_2290,N_1550,N_1684);
and U2291 (N_2291,N_1898,N_1336);
nand U2292 (N_2292,N_1528,N_1476);
nand U2293 (N_2293,N_1403,N_1705);
nor U2294 (N_2294,N_1101,N_1231);
and U2295 (N_2295,N_1139,N_1613);
nor U2296 (N_2296,N_1907,N_1494);
or U2297 (N_2297,N_1659,N_1351);
nand U2298 (N_2298,N_1305,N_1995);
and U2299 (N_2299,N_1003,N_1028);
xor U2300 (N_2300,N_1772,N_1379);
xnor U2301 (N_2301,N_1713,N_1758);
nor U2302 (N_2302,N_1503,N_1792);
and U2303 (N_2303,N_1730,N_1816);
and U2304 (N_2304,N_1463,N_1685);
and U2305 (N_2305,N_1238,N_1272);
nor U2306 (N_2306,N_1658,N_1443);
nand U2307 (N_2307,N_1618,N_1833);
or U2308 (N_2308,N_1317,N_1630);
or U2309 (N_2309,N_1370,N_1121);
xnor U2310 (N_2310,N_1822,N_1455);
and U2311 (N_2311,N_1438,N_1398);
nor U2312 (N_2312,N_1688,N_1347);
nand U2313 (N_2313,N_1353,N_1246);
nor U2314 (N_2314,N_1595,N_1075);
or U2315 (N_2315,N_1128,N_1356);
or U2316 (N_2316,N_1920,N_1538);
or U2317 (N_2317,N_1065,N_1288);
or U2318 (N_2318,N_1826,N_1633);
and U2319 (N_2319,N_1557,N_1836);
nor U2320 (N_2320,N_1144,N_1264);
and U2321 (N_2321,N_1545,N_1123);
nand U2322 (N_2322,N_1312,N_1155);
nor U2323 (N_2323,N_1828,N_1513);
xor U2324 (N_2324,N_1134,N_1570);
or U2325 (N_2325,N_1448,N_1004);
and U2326 (N_2326,N_1854,N_1221);
nor U2327 (N_2327,N_1589,N_1859);
or U2328 (N_2328,N_1387,N_1784);
nand U2329 (N_2329,N_1958,N_1966);
nand U2330 (N_2330,N_1212,N_1510);
or U2331 (N_2331,N_1217,N_1973);
or U2332 (N_2332,N_1464,N_1690);
and U2333 (N_2333,N_1722,N_1377);
nand U2334 (N_2334,N_1643,N_1434);
and U2335 (N_2335,N_1831,N_1932);
nor U2336 (N_2336,N_1923,N_1473);
and U2337 (N_2337,N_1844,N_1040);
xnor U2338 (N_2338,N_1798,N_1856);
nand U2339 (N_2339,N_1478,N_1371);
xnor U2340 (N_2340,N_1256,N_1006);
nand U2341 (N_2341,N_1248,N_1714);
nand U2342 (N_2342,N_1866,N_1001);
xor U2343 (N_2343,N_1842,N_1183);
and U2344 (N_2344,N_1279,N_1084);
nor U2345 (N_2345,N_1897,N_1865);
nand U2346 (N_2346,N_1105,N_1405);
nand U2347 (N_2347,N_1142,N_1641);
xor U2348 (N_2348,N_1223,N_1723);
and U2349 (N_2349,N_1971,N_1222);
nor U2350 (N_2350,N_1867,N_1835);
nor U2351 (N_2351,N_1837,N_1375);
or U2352 (N_2352,N_1564,N_1437);
nand U2353 (N_2353,N_1537,N_1329);
or U2354 (N_2354,N_1604,N_1858);
or U2355 (N_2355,N_1191,N_1742);
and U2356 (N_2356,N_1389,N_1612);
nand U2357 (N_2357,N_1602,N_1112);
and U2358 (N_2358,N_1787,N_1741);
nand U2359 (N_2359,N_1282,N_1472);
nor U2360 (N_2360,N_1691,N_1041);
nor U2361 (N_2361,N_1534,N_1864);
nand U2362 (N_2362,N_1344,N_1098);
nand U2363 (N_2363,N_1446,N_1036);
and U2364 (N_2364,N_1525,N_1095);
nand U2365 (N_2365,N_1135,N_1311);
nand U2366 (N_2366,N_1645,N_1695);
nor U2367 (N_2367,N_1373,N_1397);
and U2368 (N_2368,N_1514,N_1820);
or U2369 (N_2369,N_1007,N_1860);
xor U2370 (N_2370,N_1073,N_1668);
nor U2371 (N_2371,N_1117,N_1931);
nor U2372 (N_2372,N_1291,N_1976);
nor U2373 (N_2373,N_1228,N_1964);
xor U2374 (N_2374,N_1284,N_1886);
or U2375 (N_2375,N_1761,N_1149);
nor U2376 (N_2376,N_1991,N_1193);
nand U2377 (N_2377,N_1615,N_1355);
and U2378 (N_2378,N_1946,N_1628);
nor U2379 (N_2379,N_1493,N_1706);
and U2380 (N_2380,N_1855,N_1895);
or U2381 (N_2381,N_1485,N_1578);
nor U2382 (N_2382,N_1963,N_1393);
or U2383 (N_2383,N_1922,N_1331);
nor U2384 (N_2384,N_1278,N_1832);
and U2385 (N_2385,N_1197,N_1048);
and U2386 (N_2386,N_1047,N_1978);
xnor U2387 (N_2387,N_1360,N_1569);
and U2388 (N_2388,N_1617,N_1005);
nand U2389 (N_2389,N_1178,N_1497);
nor U2390 (N_2390,N_1631,N_1862);
nand U2391 (N_2391,N_1297,N_1450);
nor U2392 (N_2392,N_1586,N_1953);
or U2393 (N_2393,N_1433,N_1251);
nor U2394 (N_2394,N_1552,N_1056);
xnor U2395 (N_2395,N_1461,N_1436);
nand U2396 (N_2396,N_1313,N_1330);
or U2397 (N_2397,N_1173,N_1339);
nand U2398 (N_2398,N_1195,N_1263);
nand U2399 (N_2399,N_1374,N_1827);
nor U2400 (N_2400,N_1022,N_1718);
nand U2401 (N_2401,N_1417,N_1700);
or U2402 (N_2402,N_1182,N_1199);
nor U2403 (N_2403,N_1572,N_1164);
nor U2404 (N_2404,N_1289,N_1269);
xor U2405 (N_2405,N_1845,N_1874);
nand U2406 (N_2406,N_1949,N_1909);
nor U2407 (N_2407,N_1850,N_1840);
nand U2408 (N_2408,N_1479,N_1763);
nor U2409 (N_2409,N_1240,N_1749);
nand U2410 (N_2410,N_1621,N_1089);
and U2411 (N_2411,N_1321,N_1367);
nand U2412 (N_2412,N_1731,N_1743);
nand U2413 (N_2413,N_1619,N_1458);
or U2414 (N_2414,N_1750,N_1813);
xor U2415 (N_2415,N_1759,N_1793);
xnor U2416 (N_2416,N_1887,N_1334);
and U2417 (N_2417,N_1111,N_1176);
nand U2418 (N_2418,N_1013,N_1376);
nor U2419 (N_2419,N_1934,N_1283);
nand U2420 (N_2420,N_1893,N_1917);
nand U2421 (N_2421,N_1162,N_1783);
nand U2422 (N_2422,N_1805,N_1304);
nand U2423 (N_2423,N_1104,N_1625);
nand U2424 (N_2424,N_1935,N_1035);
nor U2425 (N_2425,N_1362,N_1801);
nand U2426 (N_2426,N_1804,N_1919);
and U2427 (N_2427,N_1152,N_1293);
and U2428 (N_2428,N_1499,N_1925);
or U2429 (N_2429,N_1926,N_1573);
or U2430 (N_2430,N_1568,N_1234);
nand U2431 (N_2431,N_1945,N_1158);
nor U2432 (N_2432,N_1024,N_1477);
nor U2433 (N_2433,N_1037,N_1138);
nand U2434 (N_2434,N_1204,N_1500);
nand U2435 (N_2435,N_1187,N_1147);
nor U2436 (N_2436,N_1306,N_1937);
and U2437 (N_2437,N_1676,N_1207);
and U2438 (N_2438,N_1938,N_1185);
or U2439 (N_2439,N_1986,N_1094);
or U2440 (N_2440,N_1046,N_1511);
or U2441 (N_2441,N_1345,N_1410);
xor U2442 (N_2442,N_1290,N_1148);
nand U2443 (N_2443,N_1664,N_1359);
nor U2444 (N_2444,N_1380,N_1261);
xor U2445 (N_2445,N_1985,N_1474);
or U2446 (N_2446,N_1349,N_1368);
nor U2447 (N_2447,N_1817,N_1608);
or U2448 (N_2448,N_1779,N_1721);
nor U2449 (N_2449,N_1959,N_1418);
or U2450 (N_2450,N_1824,N_1057);
nor U2451 (N_2451,N_1627,N_1229);
nor U2452 (N_2452,N_1481,N_1029);
xor U2453 (N_2453,N_1746,N_1002);
or U2454 (N_2454,N_1644,N_1794);
or U2455 (N_2455,N_1904,N_1770);
and U2456 (N_2456,N_1726,N_1896);
nand U2457 (N_2457,N_1558,N_1053);
or U2458 (N_2458,N_1480,N_1799);
xor U2459 (N_2459,N_1324,N_1274);
or U2460 (N_2460,N_1551,N_1975);
nand U2461 (N_2461,N_1738,N_1265);
nor U2462 (N_2462,N_1818,N_1020);
and U2463 (N_2463,N_1543,N_1930);
or U2464 (N_2464,N_1566,N_1505);
nand U2465 (N_2465,N_1675,N_1521);
xnor U2466 (N_2466,N_1470,N_1061);
and U2467 (N_2467,N_1957,N_1579);
or U2468 (N_2468,N_1157,N_1303);
nand U2469 (N_2469,N_1998,N_1912);
or U2470 (N_2470,N_1467,N_1901);
or U2471 (N_2471,N_1129,N_1086);
nand U2472 (N_2472,N_1219,N_1140);
or U2473 (N_2473,N_1352,N_1961);
and U2474 (N_2474,N_1333,N_1482);
and U2475 (N_2475,N_1597,N_1160);
or U2476 (N_2476,N_1099,N_1529);
nor U2477 (N_2477,N_1167,N_1720);
or U2478 (N_2478,N_1243,N_1296);
nand U2479 (N_2479,N_1327,N_1533);
or U2480 (N_2480,N_1201,N_1318);
and U2481 (N_2481,N_1192,N_1292);
or U2482 (N_2482,N_1921,N_1626);
nor U2483 (N_2483,N_1172,N_1724);
xnor U2484 (N_2484,N_1421,N_1715);
and U2485 (N_2485,N_1546,N_1044);
nand U2486 (N_2486,N_1027,N_1422);
or U2487 (N_2487,N_1815,N_1803);
and U2488 (N_2488,N_1849,N_1342);
nand U2489 (N_2489,N_1940,N_1392);
or U2490 (N_2490,N_1400,N_1642);
nand U2491 (N_2491,N_1326,N_1969);
nand U2492 (N_2492,N_1795,N_1102);
or U2493 (N_2493,N_1983,N_1239);
or U2494 (N_2494,N_1490,N_1875);
or U2495 (N_2495,N_1954,N_1337);
or U2496 (N_2496,N_1168,N_1058);
nand U2497 (N_2497,N_1778,N_1064);
or U2498 (N_2498,N_1394,N_1806);
and U2499 (N_2499,N_1980,N_1997);
and U2500 (N_2500,N_1889,N_1601);
or U2501 (N_2501,N_1286,N_1115);
and U2502 (N_2502,N_1461,N_1365);
xor U2503 (N_2503,N_1788,N_1187);
and U2504 (N_2504,N_1582,N_1777);
nor U2505 (N_2505,N_1651,N_1614);
or U2506 (N_2506,N_1877,N_1205);
nand U2507 (N_2507,N_1488,N_1141);
nand U2508 (N_2508,N_1083,N_1212);
and U2509 (N_2509,N_1693,N_1033);
nand U2510 (N_2510,N_1238,N_1683);
and U2511 (N_2511,N_1361,N_1428);
or U2512 (N_2512,N_1080,N_1883);
or U2513 (N_2513,N_1146,N_1783);
and U2514 (N_2514,N_1709,N_1319);
nand U2515 (N_2515,N_1466,N_1625);
xnor U2516 (N_2516,N_1796,N_1814);
xnor U2517 (N_2517,N_1773,N_1099);
and U2518 (N_2518,N_1416,N_1413);
and U2519 (N_2519,N_1552,N_1342);
or U2520 (N_2520,N_1341,N_1161);
or U2521 (N_2521,N_1996,N_1123);
and U2522 (N_2522,N_1677,N_1020);
nor U2523 (N_2523,N_1179,N_1938);
xor U2524 (N_2524,N_1087,N_1924);
and U2525 (N_2525,N_1463,N_1626);
nand U2526 (N_2526,N_1407,N_1357);
or U2527 (N_2527,N_1513,N_1324);
or U2528 (N_2528,N_1065,N_1090);
nor U2529 (N_2529,N_1524,N_1341);
xnor U2530 (N_2530,N_1545,N_1980);
and U2531 (N_2531,N_1441,N_1171);
xor U2532 (N_2532,N_1961,N_1683);
nand U2533 (N_2533,N_1046,N_1307);
or U2534 (N_2534,N_1671,N_1814);
nand U2535 (N_2535,N_1677,N_1223);
and U2536 (N_2536,N_1083,N_1893);
nor U2537 (N_2537,N_1985,N_1056);
nand U2538 (N_2538,N_1985,N_1918);
nor U2539 (N_2539,N_1083,N_1131);
or U2540 (N_2540,N_1307,N_1862);
xor U2541 (N_2541,N_1489,N_1057);
nor U2542 (N_2542,N_1870,N_1249);
and U2543 (N_2543,N_1732,N_1663);
nand U2544 (N_2544,N_1519,N_1848);
xnor U2545 (N_2545,N_1157,N_1095);
or U2546 (N_2546,N_1318,N_1209);
or U2547 (N_2547,N_1884,N_1693);
nor U2548 (N_2548,N_1739,N_1062);
and U2549 (N_2549,N_1408,N_1560);
and U2550 (N_2550,N_1506,N_1295);
and U2551 (N_2551,N_1656,N_1507);
nor U2552 (N_2552,N_1711,N_1942);
xor U2553 (N_2553,N_1491,N_1022);
or U2554 (N_2554,N_1220,N_1956);
nor U2555 (N_2555,N_1227,N_1312);
and U2556 (N_2556,N_1416,N_1105);
and U2557 (N_2557,N_1936,N_1060);
nor U2558 (N_2558,N_1813,N_1784);
and U2559 (N_2559,N_1721,N_1222);
xnor U2560 (N_2560,N_1340,N_1498);
and U2561 (N_2561,N_1832,N_1557);
and U2562 (N_2562,N_1195,N_1392);
and U2563 (N_2563,N_1632,N_1054);
nand U2564 (N_2564,N_1356,N_1165);
nand U2565 (N_2565,N_1646,N_1600);
nand U2566 (N_2566,N_1902,N_1488);
nand U2567 (N_2567,N_1372,N_1621);
or U2568 (N_2568,N_1310,N_1302);
xnor U2569 (N_2569,N_1410,N_1198);
nor U2570 (N_2570,N_1473,N_1462);
nand U2571 (N_2571,N_1507,N_1695);
nand U2572 (N_2572,N_1458,N_1405);
or U2573 (N_2573,N_1932,N_1402);
nor U2574 (N_2574,N_1219,N_1600);
and U2575 (N_2575,N_1312,N_1013);
and U2576 (N_2576,N_1884,N_1088);
nand U2577 (N_2577,N_1840,N_1238);
and U2578 (N_2578,N_1404,N_1811);
and U2579 (N_2579,N_1975,N_1305);
nor U2580 (N_2580,N_1095,N_1749);
or U2581 (N_2581,N_1979,N_1187);
or U2582 (N_2582,N_1150,N_1821);
nand U2583 (N_2583,N_1677,N_1226);
nor U2584 (N_2584,N_1261,N_1965);
nor U2585 (N_2585,N_1169,N_1191);
nand U2586 (N_2586,N_1795,N_1192);
nand U2587 (N_2587,N_1435,N_1785);
and U2588 (N_2588,N_1846,N_1146);
and U2589 (N_2589,N_1303,N_1364);
and U2590 (N_2590,N_1205,N_1136);
and U2591 (N_2591,N_1332,N_1262);
or U2592 (N_2592,N_1302,N_1995);
and U2593 (N_2593,N_1172,N_1478);
xnor U2594 (N_2594,N_1457,N_1378);
and U2595 (N_2595,N_1060,N_1813);
or U2596 (N_2596,N_1095,N_1619);
and U2597 (N_2597,N_1991,N_1589);
and U2598 (N_2598,N_1092,N_1625);
nand U2599 (N_2599,N_1951,N_1033);
and U2600 (N_2600,N_1468,N_1100);
or U2601 (N_2601,N_1669,N_1205);
and U2602 (N_2602,N_1853,N_1705);
or U2603 (N_2603,N_1040,N_1198);
or U2604 (N_2604,N_1729,N_1052);
nand U2605 (N_2605,N_1414,N_1434);
or U2606 (N_2606,N_1913,N_1549);
nand U2607 (N_2607,N_1211,N_1981);
or U2608 (N_2608,N_1623,N_1752);
or U2609 (N_2609,N_1076,N_1261);
and U2610 (N_2610,N_1283,N_1475);
nor U2611 (N_2611,N_1875,N_1277);
nor U2612 (N_2612,N_1598,N_1382);
xnor U2613 (N_2613,N_1063,N_1983);
nor U2614 (N_2614,N_1109,N_1670);
or U2615 (N_2615,N_1329,N_1703);
nand U2616 (N_2616,N_1289,N_1430);
and U2617 (N_2617,N_1703,N_1652);
nand U2618 (N_2618,N_1857,N_1258);
and U2619 (N_2619,N_1693,N_1271);
and U2620 (N_2620,N_1495,N_1081);
nand U2621 (N_2621,N_1948,N_1783);
nor U2622 (N_2622,N_1594,N_1346);
and U2623 (N_2623,N_1463,N_1221);
nand U2624 (N_2624,N_1652,N_1696);
xnor U2625 (N_2625,N_1832,N_1567);
or U2626 (N_2626,N_1117,N_1578);
xnor U2627 (N_2627,N_1747,N_1789);
or U2628 (N_2628,N_1747,N_1778);
nand U2629 (N_2629,N_1297,N_1546);
xor U2630 (N_2630,N_1799,N_1688);
and U2631 (N_2631,N_1328,N_1256);
xnor U2632 (N_2632,N_1645,N_1273);
nor U2633 (N_2633,N_1781,N_1459);
nand U2634 (N_2634,N_1226,N_1146);
nand U2635 (N_2635,N_1078,N_1520);
nor U2636 (N_2636,N_1553,N_1314);
or U2637 (N_2637,N_1055,N_1839);
or U2638 (N_2638,N_1903,N_1015);
or U2639 (N_2639,N_1183,N_1380);
and U2640 (N_2640,N_1802,N_1716);
nor U2641 (N_2641,N_1504,N_1828);
nor U2642 (N_2642,N_1002,N_1773);
or U2643 (N_2643,N_1828,N_1394);
nand U2644 (N_2644,N_1824,N_1901);
and U2645 (N_2645,N_1404,N_1756);
nand U2646 (N_2646,N_1637,N_1907);
nor U2647 (N_2647,N_1649,N_1429);
nor U2648 (N_2648,N_1043,N_1713);
and U2649 (N_2649,N_1140,N_1090);
or U2650 (N_2650,N_1283,N_1346);
and U2651 (N_2651,N_1037,N_1984);
nand U2652 (N_2652,N_1957,N_1623);
and U2653 (N_2653,N_1674,N_1792);
nor U2654 (N_2654,N_1266,N_1063);
xor U2655 (N_2655,N_1238,N_1884);
or U2656 (N_2656,N_1418,N_1173);
and U2657 (N_2657,N_1842,N_1968);
or U2658 (N_2658,N_1840,N_1303);
or U2659 (N_2659,N_1662,N_1020);
nor U2660 (N_2660,N_1703,N_1759);
and U2661 (N_2661,N_1295,N_1359);
nand U2662 (N_2662,N_1703,N_1766);
or U2663 (N_2663,N_1226,N_1931);
nand U2664 (N_2664,N_1721,N_1163);
or U2665 (N_2665,N_1705,N_1132);
nand U2666 (N_2666,N_1320,N_1028);
nand U2667 (N_2667,N_1816,N_1642);
nor U2668 (N_2668,N_1751,N_1250);
xor U2669 (N_2669,N_1758,N_1893);
xor U2670 (N_2670,N_1363,N_1007);
nand U2671 (N_2671,N_1911,N_1199);
or U2672 (N_2672,N_1046,N_1774);
nor U2673 (N_2673,N_1420,N_1478);
and U2674 (N_2674,N_1690,N_1888);
xor U2675 (N_2675,N_1576,N_1334);
nand U2676 (N_2676,N_1283,N_1003);
nor U2677 (N_2677,N_1090,N_1030);
nor U2678 (N_2678,N_1302,N_1603);
nor U2679 (N_2679,N_1985,N_1529);
nand U2680 (N_2680,N_1277,N_1881);
nor U2681 (N_2681,N_1705,N_1696);
or U2682 (N_2682,N_1441,N_1501);
and U2683 (N_2683,N_1986,N_1459);
and U2684 (N_2684,N_1821,N_1536);
or U2685 (N_2685,N_1269,N_1293);
nand U2686 (N_2686,N_1127,N_1625);
or U2687 (N_2687,N_1271,N_1089);
or U2688 (N_2688,N_1490,N_1366);
xor U2689 (N_2689,N_1293,N_1086);
nor U2690 (N_2690,N_1114,N_1451);
and U2691 (N_2691,N_1739,N_1944);
nand U2692 (N_2692,N_1385,N_1079);
xnor U2693 (N_2693,N_1760,N_1039);
and U2694 (N_2694,N_1795,N_1396);
nor U2695 (N_2695,N_1197,N_1632);
nor U2696 (N_2696,N_1214,N_1116);
or U2697 (N_2697,N_1320,N_1517);
and U2698 (N_2698,N_1460,N_1317);
nand U2699 (N_2699,N_1753,N_1745);
and U2700 (N_2700,N_1344,N_1935);
nor U2701 (N_2701,N_1054,N_1085);
and U2702 (N_2702,N_1574,N_1439);
nand U2703 (N_2703,N_1367,N_1505);
nand U2704 (N_2704,N_1944,N_1616);
nand U2705 (N_2705,N_1821,N_1867);
and U2706 (N_2706,N_1910,N_1336);
nor U2707 (N_2707,N_1525,N_1248);
and U2708 (N_2708,N_1196,N_1806);
or U2709 (N_2709,N_1307,N_1445);
nand U2710 (N_2710,N_1673,N_1735);
nand U2711 (N_2711,N_1798,N_1063);
nor U2712 (N_2712,N_1567,N_1256);
nor U2713 (N_2713,N_1771,N_1250);
nand U2714 (N_2714,N_1689,N_1451);
or U2715 (N_2715,N_1548,N_1347);
or U2716 (N_2716,N_1976,N_1397);
and U2717 (N_2717,N_1365,N_1048);
or U2718 (N_2718,N_1193,N_1822);
and U2719 (N_2719,N_1513,N_1671);
nor U2720 (N_2720,N_1597,N_1611);
and U2721 (N_2721,N_1574,N_1714);
or U2722 (N_2722,N_1302,N_1694);
nor U2723 (N_2723,N_1807,N_1494);
or U2724 (N_2724,N_1175,N_1376);
and U2725 (N_2725,N_1689,N_1874);
nor U2726 (N_2726,N_1598,N_1403);
and U2727 (N_2727,N_1923,N_1403);
or U2728 (N_2728,N_1182,N_1585);
nand U2729 (N_2729,N_1453,N_1223);
nand U2730 (N_2730,N_1216,N_1925);
nand U2731 (N_2731,N_1540,N_1248);
nor U2732 (N_2732,N_1722,N_1396);
nor U2733 (N_2733,N_1168,N_1166);
and U2734 (N_2734,N_1854,N_1826);
nand U2735 (N_2735,N_1875,N_1642);
nand U2736 (N_2736,N_1457,N_1097);
nor U2737 (N_2737,N_1610,N_1096);
nor U2738 (N_2738,N_1672,N_1618);
and U2739 (N_2739,N_1167,N_1746);
nor U2740 (N_2740,N_1037,N_1988);
xnor U2741 (N_2741,N_1687,N_1059);
or U2742 (N_2742,N_1826,N_1089);
nor U2743 (N_2743,N_1191,N_1287);
or U2744 (N_2744,N_1806,N_1318);
xnor U2745 (N_2745,N_1316,N_1029);
and U2746 (N_2746,N_1754,N_1545);
or U2747 (N_2747,N_1217,N_1391);
or U2748 (N_2748,N_1046,N_1656);
and U2749 (N_2749,N_1799,N_1106);
nor U2750 (N_2750,N_1773,N_1427);
nor U2751 (N_2751,N_1801,N_1076);
and U2752 (N_2752,N_1715,N_1072);
nor U2753 (N_2753,N_1650,N_1881);
nand U2754 (N_2754,N_1123,N_1555);
xor U2755 (N_2755,N_1560,N_1826);
and U2756 (N_2756,N_1434,N_1774);
xor U2757 (N_2757,N_1207,N_1689);
nand U2758 (N_2758,N_1035,N_1122);
and U2759 (N_2759,N_1254,N_1467);
nand U2760 (N_2760,N_1496,N_1178);
or U2761 (N_2761,N_1690,N_1416);
and U2762 (N_2762,N_1251,N_1252);
nand U2763 (N_2763,N_1642,N_1324);
and U2764 (N_2764,N_1164,N_1587);
nor U2765 (N_2765,N_1912,N_1982);
or U2766 (N_2766,N_1351,N_1057);
and U2767 (N_2767,N_1948,N_1839);
nand U2768 (N_2768,N_1298,N_1334);
and U2769 (N_2769,N_1224,N_1828);
and U2770 (N_2770,N_1496,N_1447);
xor U2771 (N_2771,N_1775,N_1268);
or U2772 (N_2772,N_1165,N_1858);
xor U2773 (N_2773,N_1712,N_1892);
nor U2774 (N_2774,N_1739,N_1348);
nand U2775 (N_2775,N_1506,N_1052);
nor U2776 (N_2776,N_1544,N_1769);
and U2777 (N_2777,N_1566,N_1278);
or U2778 (N_2778,N_1283,N_1072);
nor U2779 (N_2779,N_1695,N_1758);
xnor U2780 (N_2780,N_1565,N_1418);
nand U2781 (N_2781,N_1475,N_1367);
and U2782 (N_2782,N_1824,N_1208);
or U2783 (N_2783,N_1904,N_1968);
and U2784 (N_2784,N_1791,N_1121);
and U2785 (N_2785,N_1032,N_1973);
nand U2786 (N_2786,N_1909,N_1058);
and U2787 (N_2787,N_1202,N_1768);
or U2788 (N_2788,N_1630,N_1864);
and U2789 (N_2789,N_1703,N_1545);
nor U2790 (N_2790,N_1670,N_1270);
and U2791 (N_2791,N_1813,N_1213);
nand U2792 (N_2792,N_1825,N_1574);
xor U2793 (N_2793,N_1756,N_1799);
nand U2794 (N_2794,N_1717,N_1786);
and U2795 (N_2795,N_1637,N_1780);
and U2796 (N_2796,N_1122,N_1573);
and U2797 (N_2797,N_1060,N_1178);
nand U2798 (N_2798,N_1732,N_1729);
nor U2799 (N_2799,N_1325,N_1792);
nand U2800 (N_2800,N_1171,N_1566);
or U2801 (N_2801,N_1424,N_1069);
nor U2802 (N_2802,N_1072,N_1752);
and U2803 (N_2803,N_1535,N_1217);
or U2804 (N_2804,N_1957,N_1476);
or U2805 (N_2805,N_1077,N_1878);
nor U2806 (N_2806,N_1311,N_1417);
nor U2807 (N_2807,N_1292,N_1807);
or U2808 (N_2808,N_1531,N_1734);
or U2809 (N_2809,N_1838,N_1677);
or U2810 (N_2810,N_1359,N_1107);
nor U2811 (N_2811,N_1256,N_1108);
nor U2812 (N_2812,N_1940,N_1748);
or U2813 (N_2813,N_1371,N_1679);
nor U2814 (N_2814,N_1545,N_1611);
nand U2815 (N_2815,N_1344,N_1966);
xor U2816 (N_2816,N_1398,N_1642);
nand U2817 (N_2817,N_1684,N_1811);
xor U2818 (N_2818,N_1804,N_1770);
nor U2819 (N_2819,N_1777,N_1064);
nor U2820 (N_2820,N_1093,N_1864);
or U2821 (N_2821,N_1657,N_1083);
nor U2822 (N_2822,N_1676,N_1502);
nand U2823 (N_2823,N_1058,N_1593);
nor U2824 (N_2824,N_1875,N_1872);
xnor U2825 (N_2825,N_1986,N_1363);
and U2826 (N_2826,N_1742,N_1730);
and U2827 (N_2827,N_1188,N_1849);
nor U2828 (N_2828,N_1607,N_1283);
nor U2829 (N_2829,N_1589,N_1542);
nand U2830 (N_2830,N_1572,N_1559);
and U2831 (N_2831,N_1270,N_1849);
nor U2832 (N_2832,N_1699,N_1402);
nor U2833 (N_2833,N_1450,N_1626);
nand U2834 (N_2834,N_1665,N_1342);
or U2835 (N_2835,N_1108,N_1696);
nand U2836 (N_2836,N_1924,N_1752);
nand U2837 (N_2837,N_1985,N_1787);
nand U2838 (N_2838,N_1317,N_1047);
nand U2839 (N_2839,N_1737,N_1867);
nor U2840 (N_2840,N_1371,N_1625);
or U2841 (N_2841,N_1700,N_1034);
xor U2842 (N_2842,N_1887,N_1433);
and U2843 (N_2843,N_1802,N_1720);
nor U2844 (N_2844,N_1834,N_1765);
nor U2845 (N_2845,N_1214,N_1687);
xor U2846 (N_2846,N_1042,N_1307);
nor U2847 (N_2847,N_1922,N_1161);
xnor U2848 (N_2848,N_1618,N_1474);
xnor U2849 (N_2849,N_1707,N_1015);
or U2850 (N_2850,N_1190,N_1709);
nand U2851 (N_2851,N_1509,N_1832);
or U2852 (N_2852,N_1337,N_1249);
and U2853 (N_2853,N_1231,N_1720);
or U2854 (N_2854,N_1633,N_1994);
or U2855 (N_2855,N_1218,N_1719);
nand U2856 (N_2856,N_1035,N_1266);
nor U2857 (N_2857,N_1701,N_1198);
and U2858 (N_2858,N_1847,N_1474);
or U2859 (N_2859,N_1927,N_1767);
or U2860 (N_2860,N_1215,N_1926);
xnor U2861 (N_2861,N_1885,N_1050);
xnor U2862 (N_2862,N_1343,N_1852);
or U2863 (N_2863,N_1543,N_1936);
nor U2864 (N_2864,N_1967,N_1426);
nand U2865 (N_2865,N_1934,N_1431);
and U2866 (N_2866,N_1427,N_1580);
or U2867 (N_2867,N_1253,N_1866);
nand U2868 (N_2868,N_1301,N_1748);
nor U2869 (N_2869,N_1435,N_1962);
nand U2870 (N_2870,N_1589,N_1836);
and U2871 (N_2871,N_1118,N_1056);
nand U2872 (N_2872,N_1565,N_1142);
nand U2873 (N_2873,N_1849,N_1384);
and U2874 (N_2874,N_1965,N_1924);
and U2875 (N_2875,N_1167,N_1450);
nor U2876 (N_2876,N_1972,N_1058);
nor U2877 (N_2877,N_1230,N_1504);
or U2878 (N_2878,N_1252,N_1702);
nand U2879 (N_2879,N_1976,N_1446);
or U2880 (N_2880,N_1971,N_1056);
xnor U2881 (N_2881,N_1681,N_1888);
nand U2882 (N_2882,N_1386,N_1276);
and U2883 (N_2883,N_1589,N_1778);
nand U2884 (N_2884,N_1122,N_1584);
nand U2885 (N_2885,N_1162,N_1757);
nand U2886 (N_2886,N_1336,N_1554);
nand U2887 (N_2887,N_1600,N_1376);
or U2888 (N_2888,N_1031,N_1008);
nand U2889 (N_2889,N_1711,N_1162);
and U2890 (N_2890,N_1874,N_1286);
nor U2891 (N_2891,N_1824,N_1188);
nor U2892 (N_2892,N_1984,N_1435);
and U2893 (N_2893,N_1547,N_1019);
nand U2894 (N_2894,N_1535,N_1606);
xnor U2895 (N_2895,N_1173,N_1488);
and U2896 (N_2896,N_1090,N_1710);
nand U2897 (N_2897,N_1607,N_1444);
or U2898 (N_2898,N_1160,N_1203);
or U2899 (N_2899,N_1672,N_1390);
and U2900 (N_2900,N_1202,N_1954);
nand U2901 (N_2901,N_1548,N_1904);
nor U2902 (N_2902,N_1924,N_1252);
or U2903 (N_2903,N_1416,N_1539);
xor U2904 (N_2904,N_1555,N_1210);
xor U2905 (N_2905,N_1559,N_1965);
xor U2906 (N_2906,N_1595,N_1815);
and U2907 (N_2907,N_1886,N_1835);
nor U2908 (N_2908,N_1894,N_1233);
nor U2909 (N_2909,N_1992,N_1908);
or U2910 (N_2910,N_1869,N_1459);
nand U2911 (N_2911,N_1782,N_1354);
or U2912 (N_2912,N_1508,N_1660);
xnor U2913 (N_2913,N_1925,N_1258);
nor U2914 (N_2914,N_1024,N_1677);
and U2915 (N_2915,N_1559,N_1510);
nor U2916 (N_2916,N_1047,N_1852);
or U2917 (N_2917,N_1512,N_1135);
and U2918 (N_2918,N_1052,N_1972);
nor U2919 (N_2919,N_1897,N_1136);
xnor U2920 (N_2920,N_1411,N_1927);
xor U2921 (N_2921,N_1055,N_1162);
or U2922 (N_2922,N_1216,N_1679);
and U2923 (N_2923,N_1124,N_1530);
nor U2924 (N_2924,N_1095,N_1860);
nand U2925 (N_2925,N_1432,N_1539);
xor U2926 (N_2926,N_1858,N_1899);
or U2927 (N_2927,N_1568,N_1496);
xnor U2928 (N_2928,N_1942,N_1087);
and U2929 (N_2929,N_1093,N_1782);
or U2930 (N_2930,N_1170,N_1257);
nand U2931 (N_2931,N_1367,N_1631);
nand U2932 (N_2932,N_1256,N_1228);
and U2933 (N_2933,N_1496,N_1446);
and U2934 (N_2934,N_1851,N_1508);
nand U2935 (N_2935,N_1612,N_1927);
or U2936 (N_2936,N_1610,N_1111);
xor U2937 (N_2937,N_1223,N_1366);
nor U2938 (N_2938,N_1659,N_1952);
xnor U2939 (N_2939,N_1954,N_1793);
nor U2940 (N_2940,N_1141,N_1991);
and U2941 (N_2941,N_1604,N_1062);
nand U2942 (N_2942,N_1773,N_1569);
and U2943 (N_2943,N_1652,N_1291);
or U2944 (N_2944,N_1528,N_1306);
nand U2945 (N_2945,N_1335,N_1265);
nand U2946 (N_2946,N_1605,N_1001);
and U2947 (N_2947,N_1122,N_1531);
xnor U2948 (N_2948,N_1135,N_1422);
or U2949 (N_2949,N_1005,N_1886);
or U2950 (N_2950,N_1904,N_1095);
nor U2951 (N_2951,N_1639,N_1671);
or U2952 (N_2952,N_1242,N_1361);
or U2953 (N_2953,N_1701,N_1417);
or U2954 (N_2954,N_1182,N_1842);
or U2955 (N_2955,N_1461,N_1725);
xor U2956 (N_2956,N_1316,N_1745);
nand U2957 (N_2957,N_1297,N_1742);
or U2958 (N_2958,N_1422,N_1729);
nor U2959 (N_2959,N_1708,N_1376);
nand U2960 (N_2960,N_1577,N_1172);
or U2961 (N_2961,N_1482,N_1983);
nand U2962 (N_2962,N_1882,N_1224);
and U2963 (N_2963,N_1959,N_1027);
xor U2964 (N_2964,N_1592,N_1039);
or U2965 (N_2965,N_1823,N_1862);
xor U2966 (N_2966,N_1727,N_1385);
xor U2967 (N_2967,N_1189,N_1570);
nand U2968 (N_2968,N_1352,N_1459);
nand U2969 (N_2969,N_1524,N_1024);
nor U2970 (N_2970,N_1671,N_1581);
nand U2971 (N_2971,N_1420,N_1521);
nor U2972 (N_2972,N_1257,N_1417);
or U2973 (N_2973,N_1553,N_1578);
or U2974 (N_2974,N_1505,N_1275);
nor U2975 (N_2975,N_1646,N_1066);
and U2976 (N_2976,N_1154,N_1146);
or U2977 (N_2977,N_1133,N_1676);
and U2978 (N_2978,N_1030,N_1598);
and U2979 (N_2979,N_1052,N_1594);
nand U2980 (N_2980,N_1130,N_1923);
or U2981 (N_2981,N_1778,N_1911);
nor U2982 (N_2982,N_1969,N_1574);
and U2983 (N_2983,N_1009,N_1497);
nor U2984 (N_2984,N_1904,N_1627);
nand U2985 (N_2985,N_1553,N_1506);
and U2986 (N_2986,N_1767,N_1906);
and U2987 (N_2987,N_1120,N_1082);
or U2988 (N_2988,N_1385,N_1103);
and U2989 (N_2989,N_1284,N_1410);
or U2990 (N_2990,N_1815,N_1272);
nor U2991 (N_2991,N_1684,N_1235);
nand U2992 (N_2992,N_1828,N_1133);
and U2993 (N_2993,N_1104,N_1188);
and U2994 (N_2994,N_1848,N_1290);
or U2995 (N_2995,N_1053,N_1679);
and U2996 (N_2996,N_1350,N_1811);
or U2997 (N_2997,N_1008,N_1816);
nand U2998 (N_2998,N_1178,N_1521);
or U2999 (N_2999,N_1099,N_1143);
and U3000 (N_3000,N_2351,N_2137);
nand U3001 (N_3001,N_2079,N_2164);
and U3002 (N_3002,N_2167,N_2822);
xor U3003 (N_3003,N_2173,N_2582);
and U3004 (N_3004,N_2465,N_2427);
nand U3005 (N_3005,N_2615,N_2910);
or U3006 (N_3006,N_2852,N_2807);
nor U3007 (N_3007,N_2248,N_2260);
nand U3008 (N_3008,N_2113,N_2255);
nor U3009 (N_3009,N_2107,N_2096);
nor U3010 (N_3010,N_2492,N_2136);
and U3011 (N_3011,N_2784,N_2461);
and U3012 (N_3012,N_2873,N_2140);
nor U3013 (N_3013,N_2854,N_2832);
or U3014 (N_3014,N_2243,N_2944);
nand U3015 (N_3015,N_2808,N_2264);
nand U3016 (N_3016,N_2118,N_2451);
and U3017 (N_3017,N_2604,N_2274);
and U3018 (N_3018,N_2948,N_2573);
or U3019 (N_3019,N_2997,N_2717);
and U3020 (N_3020,N_2631,N_2198);
nand U3021 (N_3021,N_2965,N_2438);
or U3022 (N_3022,N_2031,N_2899);
nor U3023 (N_3023,N_2398,N_2916);
nand U3024 (N_3024,N_2141,N_2077);
nand U3025 (N_3025,N_2320,N_2428);
and U3026 (N_3026,N_2705,N_2287);
and U3027 (N_3027,N_2102,N_2903);
nand U3028 (N_3028,N_2601,N_2953);
and U3029 (N_3029,N_2131,N_2738);
and U3030 (N_3030,N_2922,N_2150);
nand U3031 (N_3031,N_2665,N_2895);
xor U3032 (N_3032,N_2213,N_2824);
nor U3033 (N_3033,N_2078,N_2859);
nor U3034 (N_3034,N_2285,N_2117);
and U3035 (N_3035,N_2012,N_2976);
nor U3036 (N_3036,N_2658,N_2353);
and U3037 (N_3037,N_2553,N_2112);
nand U3038 (N_3038,N_2060,N_2450);
or U3039 (N_3039,N_2099,N_2004);
nor U3040 (N_3040,N_2211,N_2172);
nand U3041 (N_3041,N_2919,N_2844);
xor U3042 (N_3042,N_2623,N_2168);
and U3043 (N_3043,N_2747,N_2086);
and U3044 (N_3044,N_2446,N_2355);
nor U3045 (N_3045,N_2116,N_2769);
xor U3046 (N_3046,N_2605,N_2128);
and U3047 (N_3047,N_2437,N_2933);
and U3048 (N_3048,N_2067,N_2776);
nor U3049 (N_3049,N_2235,N_2265);
nand U3050 (N_3050,N_2232,N_2009);
or U3051 (N_3051,N_2825,N_2126);
and U3052 (N_3052,N_2040,N_2554);
or U3053 (N_3053,N_2845,N_2072);
and U3054 (N_3054,N_2661,N_2098);
or U3055 (N_3055,N_2565,N_2068);
nor U3056 (N_3056,N_2459,N_2360);
nand U3057 (N_3057,N_2151,N_2988);
or U3058 (N_3058,N_2645,N_2901);
and U3059 (N_3059,N_2805,N_2028);
nor U3060 (N_3060,N_2469,N_2357);
or U3061 (N_3061,N_2207,N_2500);
nor U3062 (N_3062,N_2537,N_2075);
or U3063 (N_3063,N_2628,N_2340);
nor U3064 (N_3064,N_2651,N_2810);
and U3065 (N_3065,N_2608,N_2269);
or U3066 (N_3066,N_2379,N_2838);
xor U3067 (N_3067,N_2690,N_2800);
nor U3068 (N_3068,N_2954,N_2829);
nor U3069 (N_3069,N_2687,N_2526);
xor U3070 (N_3070,N_2700,N_2124);
nand U3071 (N_3071,N_2462,N_2331);
and U3072 (N_3072,N_2576,N_2013);
nor U3073 (N_3073,N_2735,N_2335);
or U3074 (N_3074,N_2319,N_2980);
or U3075 (N_3075,N_2505,N_2996);
and U3076 (N_3076,N_2882,N_2667);
xor U3077 (N_3077,N_2962,N_2839);
and U3078 (N_3078,N_2299,N_2448);
or U3079 (N_3079,N_2646,N_2550);
nand U3080 (N_3080,N_2634,N_2236);
and U3081 (N_3081,N_2036,N_2599);
nand U3082 (N_3082,N_2301,N_2404);
or U3083 (N_3083,N_2160,N_2732);
and U3084 (N_3084,N_2951,N_2796);
nor U3085 (N_3085,N_2730,N_2460);
or U3086 (N_3086,N_2445,N_2315);
or U3087 (N_3087,N_2433,N_2278);
and U3088 (N_3088,N_2135,N_2791);
nor U3089 (N_3089,N_2917,N_2836);
or U3090 (N_3090,N_2316,N_2363);
and U3091 (N_3091,N_2397,N_2749);
and U3092 (N_3092,N_2042,N_2372);
or U3093 (N_3093,N_2412,N_2406);
nand U3094 (N_3094,N_2781,N_2080);
nor U3095 (N_3095,N_2212,N_2182);
nor U3096 (N_3096,N_2765,N_2091);
xor U3097 (N_3097,N_2030,N_2921);
or U3098 (N_3098,N_2639,N_2358);
and U3099 (N_3099,N_2435,N_2253);
nand U3100 (N_3100,N_2734,N_2508);
and U3101 (N_3101,N_2386,N_2016);
nor U3102 (N_3102,N_2525,N_2205);
and U3103 (N_3103,N_2673,N_2183);
or U3104 (N_3104,N_2938,N_2345);
and U3105 (N_3105,N_2792,N_2109);
or U3106 (N_3106,N_2069,N_2580);
nor U3107 (N_3107,N_2650,N_2288);
and U3108 (N_3108,N_2929,N_2709);
nand U3109 (N_3109,N_2890,N_2401);
nand U3110 (N_3110,N_2766,N_2385);
nor U3111 (N_3111,N_2737,N_2475);
nor U3112 (N_3112,N_2426,N_2156);
or U3113 (N_3113,N_2755,N_2809);
and U3114 (N_3114,N_2005,N_2620);
nand U3115 (N_3115,N_2621,N_2216);
nand U3116 (N_3116,N_2590,N_2489);
and U3117 (N_3117,N_2330,N_2421);
or U3118 (N_3118,N_2204,N_2354);
xor U3119 (N_3119,N_2159,N_2344);
or U3120 (N_3120,N_2482,N_2498);
or U3121 (N_3121,N_2577,N_2187);
xnor U3122 (N_3122,N_2268,N_2070);
or U3123 (N_3123,N_2878,N_2277);
or U3124 (N_3124,N_2627,N_2066);
nand U3125 (N_3125,N_2991,N_2523);
or U3126 (N_3126,N_2975,N_2926);
and U3127 (N_3127,N_2617,N_2638);
nand U3128 (N_3128,N_2569,N_2990);
nand U3129 (N_3129,N_2480,N_2233);
nand U3130 (N_3130,N_2637,N_2121);
nor U3131 (N_3131,N_2348,N_2097);
or U3132 (N_3132,N_2721,N_2181);
xnor U3133 (N_3133,N_2201,N_2879);
or U3134 (N_3134,N_2564,N_2942);
and U3135 (N_3135,N_2186,N_2964);
or U3136 (N_3136,N_2994,N_2152);
and U3137 (N_3137,N_2228,N_2870);
xor U3138 (N_3138,N_2179,N_2442);
nand U3139 (N_3139,N_2192,N_2476);
or U3140 (N_3140,N_2751,N_2193);
nand U3141 (N_3141,N_2318,N_2613);
and U3142 (N_3142,N_2788,N_2487);
nor U3143 (N_3143,N_2909,N_2485);
and U3144 (N_3144,N_2453,N_2971);
xor U3145 (N_3145,N_2025,N_2297);
and U3146 (N_3146,N_2908,N_2744);
xnor U3147 (N_3147,N_2064,N_2417);
or U3148 (N_3148,N_2946,N_2706);
xor U3149 (N_3149,N_2797,N_2670);
nor U3150 (N_3150,N_2522,N_2396);
or U3151 (N_3151,N_2477,N_2241);
or U3152 (N_3152,N_2868,N_2384);
nor U3153 (N_3153,N_2710,N_2281);
or U3154 (N_3154,N_2995,N_2408);
nor U3155 (N_3155,N_2969,N_2860);
nand U3156 (N_3156,N_2105,N_2783);
nand U3157 (N_3157,N_2680,N_2325);
or U3158 (N_3158,N_2323,N_2983);
nand U3159 (N_3159,N_2444,N_2190);
or U3160 (N_3160,N_2410,N_2263);
and U3161 (N_3161,N_2813,N_2589);
xnor U3162 (N_3162,N_2782,N_2752);
nand U3163 (N_3163,N_2436,N_2468);
or U3164 (N_3164,N_2267,N_2967);
nand U3165 (N_3165,N_2373,N_2885);
nor U3166 (N_3166,N_2777,N_2974);
or U3167 (N_3167,N_2050,N_2496);
or U3168 (N_3168,N_2630,N_2367);
or U3169 (N_3169,N_2409,N_2699);
nor U3170 (N_3170,N_2609,N_2174);
or U3171 (N_3171,N_2957,N_2266);
xnor U3172 (N_3172,N_2225,N_2189);
or U3173 (N_3173,N_2607,N_2147);
and U3174 (N_3174,N_2993,N_2382);
nand U3175 (N_3175,N_2704,N_2308);
or U3176 (N_3176,N_2516,N_2364);
nor U3177 (N_3177,N_2220,N_2689);
nand U3178 (N_3178,N_2578,N_2014);
or U3179 (N_3179,N_2328,N_2332);
or U3180 (N_3180,N_2452,N_2374);
and U3181 (N_3181,N_2506,N_2127);
nand U3182 (N_3182,N_2414,N_2880);
nor U3183 (N_3183,N_2338,N_2778);
and U3184 (N_3184,N_2774,N_2591);
and U3185 (N_3185,N_2780,N_2343);
nor U3186 (N_3186,N_2745,N_2652);
and U3187 (N_3187,N_2304,N_2491);
and U3188 (N_3188,N_2302,N_2440);
or U3189 (N_3189,N_2653,N_2249);
nor U3190 (N_3190,N_2300,N_2712);
nand U3191 (N_3191,N_2146,N_2883);
nor U3192 (N_3192,N_2062,N_2368);
nand U3193 (N_3193,N_2138,N_2943);
and U3194 (N_3194,N_2219,N_2229);
or U3195 (N_3195,N_2519,N_2470);
or U3196 (N_3196,N_2835,N_2884);
and U3197 (N_3197,N_2898,N_2011);
nand U3198 (N_3198,N_2507,N_2337);
nand U3199 (N_3199,N_2855,N_2326);
and U3200 (N_3200,N_2583,N_2720);
and U3201 (N_3201,N_2272,N_2970);
nor U3202 (N_3202,N_2722,N_2043);
and U3203 (N_3203,N_2935,N_2725);
nor U3204 (N_3204,N_2529,N_2688);
nand U3205 (N_3205,N_2356,N_2635);
or U3206 (N_3206,N_2612,N_2934);
or U3207 (N_3207,N_2772,N_2415);
nor U3208 (N_3208,N_2955,N_2510);
nand U3209 (N_3209,N_2170,N_2082);
xor U3210 (N_3210,N_2891,N_2520);
or U3211 (N_3211,N_2544,N_2144);
xnor U3212 (N_3212,N_2336,N_2474);
nor U3213 (N_3213,N_2817,N_2632);
xnor U3214 (N_3214,N_2200,N_2654);
xnor U3215 (N_3215,N_2312,N_2927);
nor U3216 (N_3216,N_2439,N_2432);
nor U3217 (N_3217,N_2416,N_2130);
nor U3218 (N_3218,N_2394,N_2203);
or U3219 (N_3219,N_2940,N_2447);
or U3220 (N_3220,N_2924,N_2321);
nand U3221 (N_3221,N_2930,N_2830);
and U3222 (N_3222,N_2787,N_2913);
and U3223 (N_3223,N_2594,N_2856);
nand U3224 (N_3224,N_2949,N_2915);
nor U3225 (N_3225,N_2828,N_2286);
nor U3226 (N_3226,N_2647,N_2084);
xnor U3227 (N_3227,N_2697,N_2865);
or U3228 (N_3228,N_2618,N_2111);
and U3229 (N_3229,N_2887,N_2763);
nand U3230 (N_3230,N_2333,N_2678);
nand U3231 (N_3231,N_2058,N_2457);
and U3232 (N_3232,N_2642,N_2032);
nor U3233 (N_3233,N_2655,N_2660);
and U3234 (N_3234,N_2317,N_2375);
xnor U3235 (N_3235,N_2585,N_2918);
and U3236 (N_3236,N_2455,N_2503);
and U3237 (N_3237,N_2587,N_2430);
nor U3238 (N_3238,N_2194,N_2133);
nor U3239 (N_3239,N_2261,N_2760);
or U3240 (N_3240,N_2458,N_2244);
and U3241 (N_3241,N_2429,N_2535);
nand U3242 (N_3242,N_2561,N_2359);
nand U3243 (N_3243,N_2403,N_2208);
xor U3244 (N_3244,N_2123,N_2250);
and U3245 (N_3245,N_2958,N_2726);
or U3246 (N_3246,N_2381,N_2039);
nor U3247 (N_3247,N_2081,N_2719);
xnor U3248 (N_3248,N_2463,N_2701);
nor U3249 (N_3249,N_2149,N_2677);
and U3250 (N_3250,N_2464,N_2010);
and U3251 (N_3251,N_2511,N_2196);
nand U3252 (N_3252,N_2513,N_2795);
or U3253 (N_3253,N_2088,N_2657);
nand U3254 (N_3254,N_2346,N_2023);
nand U3255 (N_3255,N_2376,N_2224);
nor U3256 (N_3256,N_2728,N_2692);
nand U3257 (N_3257,N_2380,N_2119);
nand U3258 (N_3258,N_2163,N_2466);
xnor U3259 (N_3259,N_2986,N_2238);
nor U3260 (N_3260,N_2073,N_2662);
or U3261 (N_3261,N_2056,N_2366);
and U3262 (N_3262,N_2659,N_2467);
nor U3263 (N_3263,N_2740,N_2823);
nand U3264 (N_3264,N_2074,N_2925);
nor U3265 (N_3265,N_2104,N_2024);
or U3266 (N_3266,N_2294,N_2847);
nand U3267 (N_3267,N_2831,N_2407);
nand U3268 (N_3268,N_2998,N_2166);
nor U3269 (N_3269,N_2531,N_2682);
nand U3270 (N_3270,N_2085,N_2061);
nand U3271 (N_3271,N_2443,N_2857);
or U3272 (N_3272,N_2812,N_2191);
and U3273 (N_3273,N_2027,N_2388);
or U3274 (N_3274,N_2171,N_2614);
and U3275 (N_3275,N_2021,N_2843);
nand U3276 (N_3276,N_2402,N_2619);
nor U3277 (N_3277,N_2484,N_2158);
and U3278 (N_3278,N_2786,N_2199);
and U3279 (N_3279,N_2020,N_2046);
or U3280 (N_3280,N_2418,N_2142);
nand U3281 (N_3281,N_2252,N_2341);
and U3282 (N_3282,N_2352,N_2672);
nand U3283 (N_3283,N_2371,N_2707);
or U3284 (N_3284,N_2768,N_2675);
xnor U3285 (N_3285,N_2303,N_2959);
nand U3286 (N_3286,N_2092,N_2143);
or U3287 (N_3287,N_2549,N_2479);
nand U3288 (N_3288,N_2122,N_2454);
nor U3289 (N_3289,N_2872,N_2310);
and U3290 (N_3290,N_2848,N_2864);
nand U3291 (N_3291,N_2869,N_2515);
nand U3292 (N_3292,N_2291,N_2851);
and U3293 (N_3293,N_2669,N_2289);
or U3294 (N_3294,N_2509,N_2708);
nand U3295 (N_3295,N_2742,N_2743);
or U3296 (N_3296,N_2390,N_2434);
and U3297 (N_3297,N_2572,N_2392);
or U3298 (N_3298,N_2052,N_2517);
nor U3299 (N_3299,N_2095,N_2307);
or U3300 (N_3300,N_2779,N_2423);
xor U3301 (N_3301,N_2989,N_2888);
nand U3302 (N_3302,N_2616,N_2209);
nand U3303 (N_3303,N_2399,N_2931);
or U3304 (N_3304,N_2767,N_2377);
or U3305 (N_3305,N_2311,N_2683);
or U3306 (N_3306,N_2422,N_2258);
nor U3307 (N_3307,N_2120,N_2861);
or U3308 (N_3308,N_2750,N_2532);
nand U3309 (N_3309,N_2015,N_2110);
nor U3310 (N_3310,N_2853,N_2694);
and U3311 (N_3311,N_2889,N_2598);
nor U3312 (N_3312,N_2019,N_2047);
or U3313 (N_3313,N_2026,N_2065);
xor U3314 (N_3314,N_2862,N_2739);
nand U3315 (N_3315,N_2834,N_2863);
and U3316 (N_3316,N_2273,N_2139);
and U3317 (N_3317,N_2222,N_2696);
or U3318 (N_3318,N_2758,N_2802);
nor U3319 (N_3319,N_2071,N_2871);
or U3320 (N_3320,N_2521,N_2811);
nand U3321 (N_3321,N_2094,N_2973);
or U3322 (N_3322,N_2134,N_2486);
or U3323 (N_3323,N_2668,N_2950);
or U3324 (N_3324,N_2276,N_2488);
or U3325 (N_3325,N_2419,N_2606);
nand U3326 (N_3326,N_2256,N_2982);
nand U3327 (N_3327,N_2499,N_2920);
xor U3328 (N_3328,N_2054,N_2018);
and U3329 (N_3329,N_2902,N_2663);
xor U3330 (N_3330,N_2324,N_2000);
or U3331 (N_3331,N_2757,N_2592);
nand U3332 (N_3332,N_2037,N_2053);
and U3333 (N_3333,N_2570,N_2567);
nor U3334 (N_3334,N_2365,N_2610);
and U3335 (N_3335,N_2494,N_2671);
nand U3336 (N_3336,N_2799,N_2684);
nand U3337 (N_3337,N_2840,N_2875);
nand U3338 (N_3338,N_2257,N_2731);
nand U3339 (N_3339,N_2814,N_2035);
nand U3340 (N_3340,N_2785,N_2695);
and U3341 (N_3341,N_2197,N_2716);
nand U3342 (N_3342,N_2715,N_2034);
nand U3343 (N_3343,N_2999,N_2090);
or U3344 (N_3344,N_2849,N_2649);
or U3345 (N_3345,N_2904,N_2296);
and U3346 (N_3346,N_2533,N_2691);
xnor U3347 (N_3347,N_2478,N_2481);
nor U3348 (N_3348,N_2226,N_2002);
or U3349 (N_3349,N_2846,N_2821);
or U3350 (N_3350,N_2586,N_2383);
or U3351 (N_3351,N_2395,N_2334);
nor U3352 (N_3352,N_2033,N_2185);
nor U3353 (N_3353,N_2221,N_2076);
xor U3354 (N_3354,N_2819,N_2227);
nor U3355 (N_3355,N_2378,N_2770);
and U3356 (N_3356,N_2262,N_2968);
xor U3357 (N_3357,N_2497,N_2527);
or U3358 (N_3358,N_2979,N_2540);
nand U3359 (N_3359,N_2754,N_2771);
nor U3360 (N_3360,N_2282,N_2753);
nand U3361 (N_3361,N_2370,N_2581);
nor U3362 (N_3362,N_2571,N_2247);
or U3363 (N_3363,N_2400,N_2087);
nor U3364 (N_3364,N_2985,N_2575);
nand U3365 (N_3365,N_2275,N_2245);
nand U3366 (N_3366,N_2153,N_2548);
nor U3367 (N_3367,N_2563,N_2798);
and U3368 (N_3368,N_2552,N_2555);
and U3369 (N_3369,N_2293,N_2425);
xor U3370 (N_3370,N_2624,N_2180);
nand U3371 (N_3371,N_2178,N_2633);
nor U3372 (N_3372,N_2309,N_2806);
and U3373 (N_3373,N_2894,N_2214);
nor U3374 (N_3374,N_2937,N_2534);
and U3375 (N_3375,N_2932,N_2006);
nand U3376 (N_3376,N_2947,N_2923);
xnor U3377 (N_3377,N_2886,N_2129);
and U3378 (N_3378,N_2733,N_2698);
nand U3379 (N_3379,N_2703,N_2547);
nand U3380 (N_3380,N_2603,N_2188);
nand U3381 (N_3381,N_2530,N_2342);
nand U3382 (N_3382,N_2471,N_2283);
nand U3383 (N_3383,N_2562,N_2794);
and U3384 (N_3384,N_2055,N_2818);
nor U3385 (N_3385,N_2579,N_2347);
and U3386 (N_3386,N_2718,N_2044);
and U3387 (N_3387,N_2259,N_2231);
nand U3388 (N_3388,N_2161,N_2543);
and U3389 (N_3389,N_2837,N_2625);
nand U3390 (N_3390,N_2556,N_2115);
or U3391 (N_3391,N_2093,N_2827);
and U3392 (N_3392,N_2483,N_2804);
or U3393 (N_3393,N_2693,N_2420);
nor U3394 (N_3394,N_2702,N_2640);
xor U3395 (N_3395,N_2566,N_2905);
nor U3396 (N_3396,N_2584,N_2597);
nor U3397 (N_3397,N_2108,N_2284);
or U3398 (N_3398,N_2896,N_2501);
and U3399 (N_3399,N_2775,N_2038);
and U3400 (N_3400,N_2790,N_2928);
and U3401 (N_3401,N_2103,N_2713);
nand U3402 (N_3402,N_2801,N_2145);
and U3403 (N_3403,N_2114,N_2629);
nand U3404 (N_3404,N_2165,N_2966);
nor U3405 (N_3405,N_2008,N_2051);
nor U3406 (N_3406,N_2313,N_2759);
nor U3407 (N_3407,N_2773,N_2850);
and U3408 (N_3408,N_2685,N_2349);
or U3409 (N_3409,N_2314,N_2290);
or U3410 (N_3410,N_2936,N_2741);
nand U3411 (N_3411,N_2897,N_2559);
or U3412 (N_3412,N_2711,N_2545);
xor U3413 (N_3413,N_2393,N_2512);
xnor U3414 (N_3414,N_2029,N_2714);
xor U3415 (N_3415,N_2322,N_2641);
and U3416 (N_3416,N_2881,N_2017);
nor U3417 (N_3417,N_2254,N_2833);
xor U3418 (N_3418,N_2793,N_2217);
or U3419 (N_3419,N_2636,N_2059);
or U3420 (N_3420,N_2546,N_2912);
or U3421 (N_3421,N_2727,N_2729);
nor U3422 (N_3422,N_2761,N_2723);
nand U3423 (N_3423,N_2148,N_2106);
or U3424 (N_3424,N_2251,N_2963);
and U3425 (N_3425,N_2906,N_2041);
and U3426 (N_3426,N_2490,N_2101);
nor U3427 (N_3427,N_2361,N_2984);
nor U3428 (N_3428,N_2539,N_2648);
or U3429 (N_3429,N_2242,N_2764);
nor U3430 (N_3430,N_2866,N_2472);
nor U3431 (N_3431,N_2724,N_2369);
and U3432 (N_3432,N_2558,N_2643);
and U3433 (N_3433,N_2746,N_2952);
nand U3434 (N_3434,N_2816,N_2125);
nor U3435 (N_3435,N_2234,N_2679);
and U3436 (N_3436,N_2541,N_2280);
or U3437 (N_3437,N_2867,N_2007);
xor U3438 (N_3438,N_2978,N_2210);
and U3439 (N_3439,N_2424,N_2239);
nand U3440 (N_3440,N_2826,N_2820);
nor U3441 (N_3441,N_2387,N_2223);
and U3442 (N_3442,N_2298,N_2674);
nand U3443 (N_3443,N_2956,N_2391);
nand U3444 (N_3444,N_2972,N_2877);
xor U3445 (N_3445,N_2100,N_2939);
nor U3446 (N_3446,N_2063,N_2202);
xnor U3447 (N_3447,N_2279,N_2162);
xor U3448 (N_3448,N_2977,N_2237);
or U3449 (N_3449,N_2538,N_2551);
or U3450 (N_3450,N_2083,N_2600);
nor U3451 (N_3451,N_2132,N_2292);
or U3452 (N_3452,N_2157,N_2736);
and U3453 (N_3453,N_2449,N_2900);
or U3454 (N_3454,N_2596,N_2431);
and U3455 (N_3455,N_2339,N_2169);
nor U3456 (N_3456,N_2049,N_2022);
or U3457 (N_3457,N_2762,N_2177);
nand U3458 (N_3458,N_2175,N_2176);
and U3459 (N_3459,N_2907,N_2518);
nand U3460 (N_3460,N_2914,N_2413);
nand U3461 (N_3461,N_2045,N_2473);
and U3462 (N_3462,N_2626,N_2874);
or U3463 (N_3463,N_2841,N_2911);
or U3464 (N_3464,N_2389,N_2270);
nor U3465 (N_3465,N_2405,N_2789);
nand U3466 (N_3466,N_2504,N_2524);
and U3467 (N_3467,N_2057,N_2941);
and U3468 (N_3468,N_2756,N_2892);
nor U3469 (N_3469,N_2644,N_2441);
or U3470 (N_3470,N_2611,N_2528);
and U3471 (N_3471,N_2656,N_2327);
or U3472 (N_3472,N_2602,N_2622);
and U3473 (N_3473,N_2362,N_2686);
nor U3474 (N_3474,N_2048,N_2666);
xnor U3475 (N_3475,N_2306,N_2981);
nor U3476 (N_3476,N_2502,N_2271);
nand U3477 (N_3477,N_2195,N_2350);
and U3478 (N_3478,N_2493,N_2184);
nand U3479 (N_3479,N_2536,N_2246);
or U3480 (N_3480,N_2329,N_2215);
and U3481 (N_3481,N_2542,N_2495);
nor U3482 (N_3482,N_2295,N_2593);
nor U3483 (N_3483,N_2240,N_2305);
nand U3484 (N_3484,N_2893,N_2154);
or U3485 (N_3485,N_2945,N_2681);
nor U3486 (N_3486,N_2003,N_2568);
nor U3487 (N_3487,N_2514,N_2218);
nor U3488 (N_3488,N_2456,N_2992);
and U3489 (N_3489,N_2858,N_2748);
nand U3490 (N_3490,N_2155,N_2803);
and U3491 (N_3491,N_2206,N_2960);
or U3492 (N_3492,N_2557,N_2815);
or U3493 (N_3493,N_2560,N_2574);
or U3494 (N_3494,N_2842,N_2001);
nand U3495 (N_3495,N_2595,N_2676);
or U3496 (N_3496,N_2664,N_2411);
nand U3497 (N_3497,N_2089,N_2876);
nand U3498 (N_3498,N_2987,N_2230);
nor U3499 (N_3499,N_2961,N_2588);
nand U3500 (N_3500,N_2331,N_2531);
nand U3501 (N_3501,N_2162,N_2211);
and U3502 (N_3502,N_2501,N_2291);
or U3503 (N_3503,N_2576,N_2752);
nor U3504 (N_3504,N_2193,N_2320);
and U3505 (N_3505,N_2308,N_2504);
nand U3506 (N_3506,N_2677,N_2271);
and U3507 (N_3507,N_2406,N_2388);
nand U3508 (N_3508,N_2334,N_2212);
and U3509 (N_3509,N_2431,N_2589);
nand U3510 (N_3510,N_2005,N_2303);
or U3511 (N_3511,N_2808,N_2362);
nor U3512 (N_3512,N_2346,N_2964);
nor U3513 (N_3513,N_2120,N_2605);
nand U3514 (N_3514,N_2183,N_2668);
nand U3515 (N_3515,N_2794,N_2880);
nor U3516 (N_3516,N_2741,N_2369);
nand U3517 (N_3517,N_2173,N_2492);
nand U3518 (N_3518,N_2411,N_2385);
nand U3519 (N_3519,N_2814,N_2971);
nor U3520 (N_3520,N_2233,N_2870);
nor U3521 (N_3521,N_2347,N_2241);
and U3522 (N_3522,N_2340,N_2231);
or U3523 (N_3523,N_2144,N_2657);
or U3524 (N_3524,N_2056,N_2253);
or U3525 (N_3525,N_2380,N_2270);
or U3526 (N_3526,N_2468,N_2023);
and U3527 (N_3527,N_2981,N_2563);
xor U3528 (N_3528,N_2128,N_2313);
and U3529 (N_3529,N_2161,N_2560);
nor U3530 (N_3530,N_2717,N_2100);
and U3531 (N_3531,N_2322,N_2362);
or U3532 (N_3532,N_2774,N_2730);
nand U3533 (N_3533,N_2984,N_2357);
nand U3534 (N_3534,N_2197,N_2070);
nor U3535 (N_3535,N_2044,N_2333);
and U3536 (N_3536,N_2434,N_2508);
or U3537 (N_3537,N_2849,N_2336);
and U3538 (N_3538,N_2084,N_2391);
and U3539 (N_3539,N_2019,N_2482);
nand U3540 (N_3540,N_2280,N_2245);
xor U3541 (N_3541,N_2062,N_2522);
and U3542 (N_3542,N_2130,N_2772);
and U3543 (N_3543,N_2380,N_2111);
and U3544 (N_3544,N_2566,N_2263);
xnor U3545 (N_3545,N_2902,N_2428);
xor U3546 (N_3546,N_2732,N_2963);
and U3547 (N_3547,N_2131,N_2392);
nor U3548 (N_3548,N_2061,N_2296);
or U3549 (N_3549,N_2881,N_2960);
xor U3550 (N_3550,N_2070,N_2954);
nand U3551 (N_3551,N_2417,N_2715);
nor U3552 (N_3552,N_2140,N_2826);
or U3553 (N_3553,N_2029,N_2286);
xnor U3554 (N_3554,N_2253,N_2555);
or U3555 (N_3555,N_2141,N_2693);
and U3556 (N_3556,N_2696,N_2181);
nand U3557 (N_3557,N_2378,N_2063);
and U3558 (N_3558,N_2918,N_2269);
nand U3559 (N_3559,N_2503,N_2917);
nand U3560 (N_3560,N_2433,N_2332);
nand U3561 (N_3561,N_2945,N_2890);
nand U3562 (N_3562,N_2658,N_2100);
nand U3563 (N_3563,N_2334,N_2642);
xor U3564 (N_3564,N_2811,N_2993);
and U3565 (N_3565,N_2991,N_2203);
nand U3566 (N_3566,N_2424,N_2954);
nand U3567 (N_3567,N_2334,N_2942);
nor U3568 (N_3568,N_2595,N_2830);
nor U3569 (N_3569,N_2267,N_2760);
nor U3570 (N_3570,N_2200,N_2579);
or U3571 (N_3571,N_2633,N_2776);
nor U3572 (N_3572,N_2287,N_2595);
or U3573 (N_3573,N_2355,N_2995);
and U3574 (N_3574,N_2844,N_2648);
nand U3575 (N_3575,N_2197,N_2530);
nor U3576 (N_3576,N_2603,N_2632);
and U3577 (N_3577,N_2230,N_2430);
and U3578 (N_3578,N_2012,N_2687);
or U3579 (N_3579,N_2997,N_2929);
xor U3580 (N_3580,N_2080,N_2874);
and U3581 (N_3581,N_2267,N_2574);
nor U3582 (N_3582,N_2314,N_2856);
nor U3583 (N_3583,N_2407,N_2768);
xor U3584 (N_3584,N_2505,N_2512);
or U3585 (N_3585,N_2522,N_2661);
or U3586 (N_3586,N_2730,N_2255);
nor U3587 (N_3587,N_2195,N_2403);
nand U3588 (N_3588,N_2256,N_2720);
nor U3589 (N_3589,N_2801,N_2265);
nor U3590 (N_3590,N_2414,N_2093);
or U3591 (N_3591,N_2311,N_2645);
nor U3592 (N_3592,N_2476,N_2305);
and U3593 (N_3593,N_2093,N_2705);
or U3594 (N_3594,N_2475,N_2833);
nor U3595 (N_3595,N_2212,N_2734);
nor U3596 (N_3596,N_2989,N_2592);
nor U3597 (N_3597,N_2598,N_2961);
xnor U3598 (N_3598,N_2063,N_2587);
xnor U3599 (N_3599,N_2906,N_2715);
or U3600 (N_3600,N_2510,N_2617);
nor U3601 (N_3601,N_2302,N_2275);
nand U3602 (N_3602,N_2224,N_2665);
nand U3603 (N_3603,N_2948,N_2448);
xor U3604 (N_3604,N_2439,N_2910);
nor U3605 (N_3605,N_2325,N_2370);
and U3606 (N_3606,N_2119,N_2774);
and U3607 (N_3607,N_2662,N_2984);
or U3608 (N_3608,N_2292,N_2951);
nand U3609 (N_3609,N_2701,N_2125);
xnor U3610 (N_3610,N_2571,N_2085);
and U3611 (N_3611,N_2159,N_2922);
or U3612 (N_3612,N_2501,N_2339);
or U3613 (N_3613,N_2042,N_2601);
xnor U3614 (N_3614,N_2614,N_2520);
or U3615 (N_3615,N_2893,N_2379);
or U3616 (N_3616,N_2701,N_2393);
or U3617 (N_3617,N_2578,N_2902);
nand U3618 (N_3618,N_2385,N_2974);
nor U3619 (N_3619,N_2384,N_2792);
and U3620 (N_3620,N_2559,N_2339);
nand U3621 (N_3621,N_2981,N_2920);
nand U3622 (N_3622,N_2647,N_2565);
xnor U3623 (N_3623,N_2263,N_2161);
and U3624 (N_3624,N_2420,N_2951);
and U3625 (N_3625,N_2730,N_2258);
xnor U3626 (N_3626,N_2732,N_2577);
nor U3627 (N_3627,N_2394,N_2169);
nor U3628 (N_3628,N_2938,N_2179);
nor U3629 (N_3629,N_2512,N_2173);
or U3630 (N_3630,N_2929,N_2264);
and U3631 (N_3631,N_2784,N_2310);
nand U3632 (N_3632,N_2479,N_2889);
or U3633 (N_3633,N_2608,N_2274);
or U3634 (N_3634,N_2756,N_2736);
nand U3635 (N_3635,N_2137,N_2915);
or U3636 (N_3636,N_2397,N_2657);
nor U3637 (N_3637,N_2022,N_2375);
or U3638 (N_3638,N_2786,N_2956);
and U3639 (N_3639,N_2694,N_2767);
or U3640 (N_3640,N_2011,N_2515);
nand U3641 (N_3641,N_2799,N_2119);
and U3642 (N_3642,N_2210,N_2432);
or U3643 (N_3643,N_2966,N_2662);
and U3644 (N_3644,N_2391,N_2882);
or U3645 (N_3645,N_2201,N_2543);
xor U3646 (N_3646,N_2348,N_2026);
or U3647 (N_3647,N_2200,N_2419);
and U3648 (N_3648,N_2929,N_2020);
nand U3649 (N_3649,N_2431,N_2324);
or U3650 (N_3650,N_2980,N_2345);
or U3651 (N_3651,N_2316,N_2832);
and U3652 (N_3652,N_2836,N_2677);
and U3653 (N_3653,N_2106,N_2387);
and U3654 (N_3654,N_2166,N_2822);
nor U3655 (N_3655,N_2857,N_2152);
nor U3656 (N_3656,N_2115,N_2766);
nor U3657 (N_3657,N_2896,N_2651);
or U3658 (N_3658,N_2664,N_2432);
nor U3659 (N_3659,N_2995,N_2317);
nand U3660 (N_3660,N_2863,N_2190);
xor U3661 (N_3661,N_2737,N_2245);
and U3662 (N_3662,N_2434,N_2211);
or U3663 (N_3663,N_2115,N_2533);
nand U3664 (N_3664,N_2533,N_2135);
nor U3665 (N_3665,N_2997,N_2061);
and U3666 (N_3666,N_2930,N_2600);
nand U3667 (N_3667,N_2689,N_2179);
nand U3668 (N_3668,N_2973,N_2652);
nor U3669 (N_3669,N_2930,N_2004);
and U3670 (N_3670,N_2913,N_2707);
nor U3671 (N_3671,N_2372,N_2633);
and U3672 (N_3672,N_2336,N_2134);
or U3673 (N_3673,N_2500,N_2772);
or U3674 (N_3674,N_2442,N_2608);
and U3675 (N_3675,N_2707,N_2948);
nor U3676 (N_3676,N_2443,N_2981);
or U3677 (N_3677,N_2306,N_2560);
and U3678 (N_3678,N_2483,N_2948);
nand U3679 (N_3679,N_2350,N_2816);
nand U3680 (N_3680,N_2147,N_2385);
nor U3681 (N_3681,N_2332,N_2090);
and U3682 (N_3682,N_2700,N_2767);
nor U3683 (N_3683,N_2347,N_2677);
nand U3684 (N_3684,N_2043,N_2483);
and U3685 (N_3685,N_2238,N_2729);
or U3686 (N_3686,N_2447,N_2507);
and U3687 (N_3687,N_2128,N_2765);
and U3688 (N_3688,N_2589,N_2362);
xor U3689 (N_3689,N_2163,N_2381);
xnor U3690 (N_3690,N_2786,N_2971);
and U3691 (N_3691,N_2719,N_2181);
nand U3692 (N_3692,N_2422,N_2494);
nor U3693 (N_3693,N_2706,N_2429);
nand U3694 (N_3694,N_2836,N_2190);
or U3695 (N_3695,N_2811,N_2606);
and U3696 (N_3696,N_2349,N_2146);
nand U3697 (N_3697,N_2677,N_2459);
nand U3698 (N_3698,N_2120,N_2602);
and U3699 (N_3699,N_2095,N_2561);
nor U3700 (N_3700,N_2547,N_2334);
nand U3701 (N_3701,N_2154,N_2680);
nor U3702 (N_3702,N_2931,N_2817);
nand U3703 (N_3703,N_2302,N_2543);
nand U3704 (N_3704,N_2890,N_2328);
or U3705 (N_3705,N_2669,N_2618);
and U3706 (N_3706,N_2936,N_2833);
nand U3707 (N_3707,N_2067,N_2579);
xnor U3708 (N_3708,N_2192,N_2777);
xor U3709 (N_3709,N_2481,N_2193);
and U3710 (N_3710,N_2664,N_2982);
or U3711 (N_3711,N_2412,N_2443);
nand U3712 (N_3712,N_2485,N_2877);
or U3713 (N_3713,N_2757,N_2970);
and U3714 (N_3714,N_2877,N_2953);
and U3715 (N_3715,N_2846,N_2152);
or U3716 (N_3716,N_2848,N_2509);
xnor U3717 (N_3717,N_2929,N_2289);
nand U3718 (N_3718,N_2116,N_2372);
nand U3719 (N_3719,N_2426,N_2934);
nor U3720 (N_3720,N_2914,N_2171);
nand U3721 (N_3721,N_2826,N_2971);
or U3722 (N_3722,N_2366,N_2963);
nand U3723 (N_3723,N_2995,N_2139);
and U3724 (N_3724,N_2833,N_2133);
and U3725 (N_3725,N_2329,N_2616);
nand U3726 (N_3726,N_2914,N_2938);
and U3727 (N_3727,N_2924,N_2134);
xor U3728 (N_3728,N_2496,N_2210);
nand U3729 (N_3729,N_2142,N_2263);
nand U3730 (N_3730,N_2742,N_2372);
nor U3731 (N_3731,N_2859,N_2543);
nand U3732 (N_3732,N_2118,N_2314);
and U3733 (N_3733,N_2048,N_2427);
nor U3734 (N_3734,N_2854,N_2034);
and U3735 (N_3735,N_2259,N_2648);
nor U3736 (N_3736,N_2515,N_2259);
nor U3737 (N_3737,N_2690,N_2103);
and U3738 (N_3738,N_2366,N_2523);
or U3739 (N_3739,N_2143,N_2405);
or U3740 (N_3740,N_2183,N_2532);
or U3741 (N_3741,N_2086,N_2723);
and U3742 (N_3742,N_2811,N_2643);
nor U3743 (N_3743,N_2781,N_2466);
or U3744 (N_3744,N_2143,N_2475);
and U3745 (N_3745,N_2070,N_2800);
or U3746 (N_3746,N_2368,N_2854);
nor U3747 (N_3747,N_2900,N_2363);
xnor U3748 (N_3748,N_2301,N_2635);
or U3749 (N_3749,N_2640,N_2154);
nor U3750 (N_3750,N_2897,N_2003);
nor U3751 (N_3751,N_2673,N_2489);
nand U3752 (N_3752,N_2901,N_2252);
or U3753 (N_3753,N_2336,N_2346);
xor U3754 (N_3754,N_2606,N_2070);
or U3755 (N_3755,N_2759,N_2214);
or U3756 (N_3756,N_2493,N_2484);
nand U3757 (N_3757,N_2581,N_2484);
or U3758 (N_3758,N_2867,N_2384);
nor U3759 (N_3759,N_2847,N_2511);
nor U3760 (N_3760,N_2355,N_2284);
nor U3761 (N_3761,N_2108,N_2162);
or U3762 (N_3762,N_2778,N_2337);
nor U3763 (N_3763,N_2579,N_2657);
xor U3764 (N_3764,N_2713,N_2182);
or U3765 (N_3765,N_2181,N_2917);
nand U3766 (N_3766,N_2383,N_2661);
nor U3767 (N_3767,N_2274,N_2460);
nand U3768 (N_3768,N_2238,N_2751);
or U3769 (N_3769,N_2546,N_2835);
and U3770 (N_3770,N_2439,N_2614);
xor U3771 (N_3771,N_2116,N_2074);
or U3772 (N_3772,N_2847,N_2347);
and U3773 (N_3773,N_2910,N_2084);
xnor U3774 (N_3774,N_2424,N_2156);
and U3775 (N_3775,N_2756,N_2883);
or U3776 (N_3776,N_2584,N_2207);
and U3777 (N_3777,N_2888,N_2380);
or U3778 (N_3778,N_2644,N_2801);
nand U3779 (N_3779,N_2314,N_2021);
nor U3780 (N_3780,N_2253,N_2868);
nor U3781 (N_3781,N_2152,N_2320);
or U3782 (N_3782,N_2779,N_2361);
nor U3783 (N_3783,N_2975,N_2563);
and U3784 (N_3784,N_2960,N_2909);
xnor U3785 (N_3785,N_2017,N_2401);
and U3786 (N_3786,N_2914,N_2758);
nand U3787 (N_3787,N_2775,N_2271);
xor U3788 (N_3788,N_2095,N_2005);
nand U3789 (N_3789,N_2493,N_2467);
nor U3790 (N_3790,N_2333,N_2708);
nor U3791 (N_3791,N_2149,N_2861);
nor U3792 (N_3792,N_2218,N_2185);
and U3793 (N_3793,N_2350,N_2356);
or U3794 (N_3794,N_2847,N_2769);
nor U3795 (N_3795,N_2640,N_2901);
nor U3796 (N_3796,N_2247,N_2425);
nand U3797 (N_3797,N_2167,N_2051);
and U3798 (N_3798,N_2459,N_2997);
nand U3799 (N_3799,N_2505,N_2717);
nor U3800 (N_3800,N_2375,N_2943);
nor U3801 (N_3801,N_2128,N_2103);
or U3802 (N_3802,N_2948,N_2482);
nor U3803 (N_3803,N_2409,N_2438);
or U3804 (N_3804,N_2823,N_2445);
nor U3805 (N_3805,N_2305,N_2551);
or U3806 (N_3806,N_2508,N_2983);
xor U3807 (N_3807,N_2139,N_2933);
nor U3808 (N_3808,N_2807,N_2926);
nor U3809 (N_3809,N_2208,N_2927);
nor U3810 (N_3810,N_2326,N_2056);
nor U3811 (N_3811,N_2331,N_2951);
or U3812 (N_3812,N_2305,N_2794);
nand U3813 (N_3813,N_2889,N_2886);
or U3814 (N_3814,N_2002,N_2240);
or U3815 (N_3815,N_2970,N_2679);
nor U3816 (N_3816,N_2134,N_2554);
nor U3817 (N_3817,N_2210,N_2229);
nand U3818 (N_3818,N_2303,N_2910);
or U3819 (N_3819,N_2790,N_2403);
or U3820 (N_3820,N_2851,N_2219);
nor U3821 (N_3821,N_2857,N_2044);
or U3822 (N_3822,N_2970,N_2447);
nand U3823 (N_3823,N_2778,N_2149);
and U3824 (N_3824,N_2184,N_2085);
or U3825 (N_3825,N_2834,N_2129);
and U3826 (N_3826,N_2836,N_2706);
nand U3827 (N_3827,N_2100,N_2964);
nand U3828 (N_3828,N_2580,N_2397);
nor U3829 (N_3829,N_2273,N_2522);
and U3830 (N_3830,N_2444,N_2572);
nand U3831 (N_3831,N_2910,N_2062);
and U3832 (N_3832,N_2024,N_2655);
or U3833 (N_3833,N_2242,N_2954);
xor U3834 (N_3834,N_2780,N_2848);
nand U3835 (N_3835,N_2592,N_2487);
and U3836 (N_3836,N_2314,N_2078);
and U3837 (N_3837,N_2461,N_2899);
xnor U3838 (N_3838,N_2584,N_2286);
nor U3839 (N_3839,N_2722,N_2636);
and U3840 (N_3840,N_2073,N_2758);
or U3841 (N_3841,N_2807,N_2359);
nand U3842 (N_3842,N_2056,N_2901);
nor U3843 (N_3843,N_2771,N_2806);
and U3844 (N_3844,N_2710,N_2195);
nand U3845 (N_3845,N_2197,N_2452);
nor U3846 (N_3846,N_2834,N_2774);
nand U3847 (N_3847,N_2647,N_2817);
or U3848 (N_3848,N_2135,N_2638);
nor U3849 (N_3849,N_2561,N_2205);
or U3850 (N_3850,N_2615,N_2135);
nand U3851 (N_3851,N_2073,N_2661);
nand U3852 (N_3852,N_2537,N_2575);
nor U3853 (N_3853,N_2288,N_2220);
and U3854 (N_3854,N_2194,N_2837);
and U3855 (N_3855,N_2242,N_2633);
or U3856 (N_3856,N_2338,N_2203);
nand U3857 (N_3857,N_2186,N_2437);
xnor U3858 (N_3858,N_2547,N_2991);
xnor U3859 (N_3859,N_2216,N_2702);
and U3860 (N_3860,N_2519,N_2640);
nor U3861 (N_3861,N_2924,N_2131);
nand U3862 (N_3862,N_2317,N_2938);
xnor U3863 (N_3863,N_2336,N_2794);
and U3864 (N_3864,N_2418,N_2973);
or U3865 (N_3865,N_2111,N_2795);
xnor U3866 (N_3866,N_2868,N_2845);
and U3867 (N_3867,N_2747,N_2579);
xor U3868 (N_3868,N_2035,N_2117);
xor U3869 (N_3869,N_2164,N_2192);
nand U3870 (N_3870,N_2044,N_2158);
nor U3871 (N_3871,N_2468,N_2975);
xor U3872 (N_3872,N_2738,N_2581);
and U3873 (N_3873,N_2246,N_2906);
nor U3874 (N_3874,N_2923,N_2530);
nand U3875 (N_3875,N_2552,N_2792);
or U3876 (N_3876,N_2002,N_2530);
nor U3877 (N_3877,N_2944,N_2262);
or U3878 (N_3878,N_2931,N_2688);
or U3879 (N_3879,N_2601,N_2584);
or U3880 (N_3880,N_2868,N_2314);
and U3881 (N_3881,N_2025,N_2150);
nor U3882 (N_3882,N_2015,N_2431);
nand U3883 (N_3883,N_2986,N_2535);
and U3884 (N_3884,N_2968,N_2162);
nand U3885 (N_3885,N_2749,N_2888);
nand U3886 (N_3886,N_2513,N_2076);
nor U3887 (N_3887,N_2113,N_2670);
nand U3888 (N_3888,N_2497,N_2949);
and U3889 (N_3889,N_2616,N_2274);
nand U3890 (N_3890,N_2215,N_2908);
xor U3891 (N_3891,N_2228,N_2541);
and U3892 (N_3892,N_2205,N_2117);
xor U3893 (N_3893,N_2304,N_2911);
and U3894 (N_3894,N_2846,N_2909);
or U3895 (N_3895,N_2209,N_2521);
nand U3896 (N_3896,N_2323,N_2615);
xnor U3897 (N_3897,N_2206,N_2094);
and U3898 (N_3898,N_2659,N_2695);
or U3899 (N_3899,N_2400,N_2671);
or U3900 (N_3900,N_2357,N_2534);
nor U3901 (N_3901,N_2747,N_2481);
or U3902 (N_3902,N_2020,N_2845);
and U3903 (N_3903,N_2968,N_2083);
or U3904 (N_3904,N_2233,N_2114);
nand U3905 (N_3905,N_2648,N_2241);
and U3906 (N_3906,N_2261,N_2969);
nor U3907 (N_3907,N_2197,N_2368);
nor U3908 (N_3908,N_2873,N_2529);
nor U3909 (N_3909,N_2453,N_2700);
and U3910 (N_3910,N_2625,N_2862);
or U3911 (N_3911,N_2202,N_2371);
or U3912 (N_3912,N_2799,N_2204);
xor U3913 (N_3913,N_2319,N_2835);
or U3914 (N_3914,N_2549,N_2591);
and U3915 (N_3915,N_2497,N_2743);
and U3916 (N_3916,N_2005,N_2166);
and U3917 (N_3917,N_2295,N_2729);
nor U3918 (N_3918,N_2111,N_2866);
and U3919 (N_3919,N_2403,N_2666);
nor U3920 (N_3920,N_2540,N_2914);
nor U3921 (N_3921,N_2947,N_2373);
or U3922 (N_3922,N_2651,N_2813);
or U3923 (N_3923,N_2736,N_2105);
xor U3924 (N_3924,N_2616,N_2051);
nand U3925 (N_3925,N_2241,N_2781);
or U3926 (N_3926,N_2888,N_2311);
and U3927 (N_3927,N_2060,N_2324);
or U3928 (N_3928,N_2041,N_2904);
nor U3929 (N_3929,N_2631,N_2579);
nor U3930 (N_3930,N_2897,N_2825);
nor U3931 (N_3931,N_2645,N_2193);
nand U3932 (N_3932,N_2032,N_2350);
nand U3933 (N_3933,N_2460,N_2546);
or U3934 (N_3934,N_2399,N_2560);
and U3935 (N_3935,N_2301,N_2253);
or U3936 (N_3936,N_2969,N_2067);
nand U3937 (N_3937,N_2654,N_2667);
and U3938 (N_3938,N_2953,N_2306);
and U3939 (N_3939,N_2568,N_2678);
and U3940 (N_3940,N_2858,N_2579);
xnor U3941 (N_3941,N_2649,N_2278);
xnor U3942 (N_3942,N_2354,N_2871);
nor U3943 (N_3943,N_2596,N_2798);
nor U3944 (N_3944,N_2526,N_2580);
xnor U3945 (N_3945,N_2747,N_2066);
nand U3946 (N_3946,N_2179,N_2796);
nand U3947 (N_3947,N_2606,N_2271);
nor U3948 (N_3948,N_2960,N_2457);
or U3949 (N_3949,N_2187,N_2474);
xnor U3950 (N_3950,N_2601,N_2397);
nor U3951 (N_3951,N_2996,N_2099);
nand U3952 (N_3952,N_2531,N_2074);
and U3953 (N_3953,N_2590,N_2491);
or U3954 (N_3954,N_2811,N_2611);
xor U3955 (N_3955,N_2470,N_2619);
and U3956 (N_3956,N_2105,N_2568);
xor U3957 (N_3957,N_2872,N_2093);
nand U3958 (N_3958,N_2372,N_2679);
nor U3959 (N_3959,N_2630,N_2818);
or U3960 (N_3960,N_2386,N_2402);
nor U3961 (N_3961,N_2476,N_2359);
nor U3962 (N_3962,N_2633,N_2913);
nand U3963 (N_3963,N_2736,N_2826);
and U3964 (N_3964,N_2085,N_2798);
and U3965 (N_3965,N_2905,N_2308);
or U3966 (N_3966,N_2413,N_2351);
and U3967 (N_3967,N_2045,N_2105);
nand U3968 (N_3968,N_2174,N_2707);
and U3969 (N_3969,N_2660,N_2359);
xor U3970 (N_3970,N_2306,N_2171);
nor U3971 (N_3971,N_2908,N_2920);
or U3972 (N_3972,N_2851,N_2779);
nor U3973 (N_3973,N_2078,N_2310);
and U3974 (N_3974,N_2227,N_2192);
nor U3975 (N_3975,N_2081,N_2145);
nand U3976 (N_3976,N_2645,N_2813);
nor U3977 (N_3977,N_2688,N_2497);
nand U3978 (N_3978,N_2617,N_2650);
nand U3979 (N_3979,N_2528,N_2721);
nor U3980 (N_3980,N_2511,N_2424);
and U3981 (N_3981,N_2273,N_2257);
and U3982 (N_3982,N_2643,N_2878);
or U3983 (N_3983,N_2931,N_2028);
and U3984 (N_3984,N_2700,N_2763);
nor U3985 (N_3985,N_2518,N_2602);
and U3986 (N_3986,N_2848,N_2081);
nand U3987 (N_3987,N_2744,N_2188);
nand U3988 (N_3988,N_2381,N_2014);
nand U3989 (N_3989,N_2377,N_2279);
or U3990 (N_3990,N_2979,N_2359);
and U3991 (N_3991,N_2982,N_2404);
nor U3992 (N_3992,N_2251,N_2635);
or U3993 (N_3993,N_2991,N_2498);
and U3994 (N_3994,N_2307,N_2262);
xor U3995 (N_3995,N_2362,N_2022);
nor U3996 (N_3996,N_2636,N_2828);
or U3997 (N_3997,N_2454,N_2818);
or U3998 (N_3998,N_2505,N_2745);
xnor U3999 (N_3999,N_2705,N_2932);
nand U4000 (N_4000,N_3936,N_3420);
nor U4001 (N_4001,N_3690,N_3860);
nor U4002 (N_4002,N_3008,N_3451);
nor U4003 (N_4003,N_3122,N_3150);
nor U4004 (N_4004,N_3842,N_3721);
or U4005 (N_4005,N_3571,N_3095);
nor U4006 (N_4006,N_3823,N_3959);
nor U4007 (N_4007,N_3141,N_3779);
nand U4008 (N_4008,N_3198,N_3203);
or U4009 (N_4009,N_3165,N_3256);
nor U4010 (N_4010,N_3543,N_3263);
nand U4011 (N_4011,N_3989,N_3605);
nor U4012 (N_4012,N_3038,N_3125);
nand U4013 (N_4013,N_3128,N_3152);
and U4014 (N_4014,N_3737,N_3209);
and U4015 (N_4015,N_3376,N_3944);
and U4016 (N_4016,N_3205,N_3522);
and U4017 (N_4017,N_3683,N_3879);
or U4018 (N_4018,N_3770,N_3837);
and U4019 (N_4019,N_3583,N_3418);
xor U4020 (N_4020,N_3354,N_3662);
or U4021 (N_4021,N_3439,N_3600);
or U4022 (N_4022,N_3170,N_3121);
nor U4023 (N_4023,N_3180,N_3063);
or U4024 (N_4024,N_3005,N_3970);
nor U4025 (N_4025,N_3857,N_3328);
and U4026 (N_4026,N_3114,N_3838);
and U4027 (N_4027,N_3753,N_3934);
or U4028 (N_4028,N_3850,N_3361);
xnor U4029 (N_4029,N_3679,N_3937);
nand U4030 (N_4030,N_3100,N_3990);
nand U4031 (N_4031,N_3611,N_3424);
and U4032 (N_4032,N_3493,N_3188);
and U4033 (N_4033,N_3259,N_3289);
or U4034 (N_4034,N_3775,N_3034);
nand U4035 (N_4035,N_3037,N_3137);
nor U4036 (N_4036,N_3680,N_3093);
or U4037 (N_4037,N_3364,N_3469);
nor U4038 (N_4038,N_3254,N_3334);
or U4039 (N_4039,N_3549,N_3978);
nand U4040 (N_4040,N_3131,N_3616);
or U4041 (N_4041,N_3294,N_3278);
nor U4042 (N_4042,N_3658,N_3450);
nor U4043 (N_4043,N_3385,N_3210);
xnor U4044 (N_4044,N_3113,N_3999);
nor U4045 (N_4045,N_3484,N_3781);
nor U4046 (N_4046,N_3962,N_3404);
and U4047 (N_4047,N_3363,N_3515);
and U4048 (N_4048,N_3544,N_3692);
nor U4049 (N_4049,N_3232,N_3175);
nor U4050 (N_4050,N_3297,N_3226);
nor U4051 (N_4051,N_3168,N_3929);
nand U4052 (N_4052,N_3221,N_3715);
and U4053 (N_4053,N_3269,N_3567);
or U4054 (N_4054,N_3598,N_3058);
and U4055 (N_4055,N_3634,N_3280);
nor U4056 (N_4056,N_3824,N_3323);
nor U4057 (N_4057,N_3862,N_3265);
and U4058 (N_4058,N_3649,N_3140);
or U4059 (N_4059,N_3403,N_3446);
nand U4060 (N_4060,N_3873,N_3318);
nor U4061 (N_4061,N_3142,N_3998);
nor U4062 (N_4062,N_3176,N_3985);
nand U4063 (N_4063,N_3836,N_3080);
or U4064 (N_4064,N_3395,N_3725);
or U4065 (N_4065,N_3199,N_3609);
and U4066 (N_4066,N_3160,N_3275);
nor U4067 (N_4067,N_3388,N_3138);
nor U4068 (N_4068,N_3077,N_3052);
nand U4069 (N_4069,N_3468,N_3440);
and U4070 (N_4070,N_3389,N_3988);
nand U4071 (N_4071,N_3072,N_3815);
or U4072 (N_4072,N_3155,N_3143);
or U4073 (N_4073,N_3698,N_3992);
xnor U4074 (N_4074,N_3736,N_3236);
xnor U4075 (N_4075,N_3499,N_3848);
nor U4076 (N_4076,N_3496,N_3261);
nor U4077 (N_4077,N_3082,N_3880);
nand U4078 (N_4078,N_3043,N_3581);
and U4079 (N_4079,N_3467,N_3518);
nor U4080 (N_4080,N_3791,N_3044);
nand U4081 (N_4081,N_3218,N_3716);
nand U4082 (N_4082,N_3246,N_3761);
nand U4083 (N_4083,N_3956,N_3586);
and U4084 (N_4084,N_3964,N_3464);
or U4085 (N_4085,N_3909,N_3103);
nand U4086 (N_4086,N_3902,N_3134);
and U4087 (N_4087,N_3327,N_3671);
nor U4088 (N_4088,N_3454,N_3391);
or U4089 (N_4089,N_3578,N_3763);
and U4090 (N_4090,N_3808,N_3007);
or U4091 (N_4091,N_3248,N_3303);
nor U4092 (N_4092,N_3996,N_3437);
nand U4093 (N_4093,N_3161,N_3979);
or U4094 (N_4094,N_3045,N_3296);
nand U4095 (N_4095,N_3951,N_3587);
nand U4096 (N_4096,N_3215,N_3238);
nand U4097 (N_4097,N_3241,N_3596);
xor U4098 (N_4098,N_3552,N_3745);
nor U4099 (N_4099,N_3928,N_3517);
or U4100 (N_4100,N_3345,N_3426);
nor U4101 (N_4101,N_3379,N_3078);
and U4102 (N_4102,N_3268,N_3738);
and U4103 (N_4103,N_3739,N_3710);
nand U4104 (N_4104,N_3864,N_3251);
nor U4105 (N_4105,N_3833,N_3516);
or U4106 (N_4106,N_3105,N_3333);
nor U4107 (N_4107,N_3235,N_3473);
and U4108 (N_4108,N_3971,N_3788);
and U4109 (N_4109,N_3387,N_3789);
nor U4110 (N_4110,N_3291,N_3491);
nor U4111 (N_4111,N_3352,N_3682);
or U4112 (N_4112,N_3017,N_3868);
nor U4113 (N_4113,N_3640,N_3915);
and U4114 (N_4114,N_3267,N_3346);
nor U4115 (N_4115,N_3025,N_3947);
and U4116 (N_4116,N_3776,N_3503);
and U4117 (N_4117,N_3656,N_3326);
nand U4118 (N_4118,N_3559,N_3109);
nor U4119 (N_4119,N_3347,N_3993);
or U4120 (N_4120,N_3623,N_3801);
nor U4121 (N_4121,N_3191,N_3351);
or U4122 (N_4122,N_3877,N_3432);
and U4123 (N_4123,N_3126,N_3130);
nor U4124 (N_4124,N_3362,N_3633);
and U4125 (N_4125,N_3237,N_3627);
nand U4126 (N_4126,N_3953,N_3967);
xnor U4127 (N_4127,N_3039,N_3691);
xor U4128 (N_4128,N_3494,N_3421);
xor U4129 (N_4129,N_3825,N_3643);
or U4130 (N_4130,N_3146,N_3787);
xnor U4131 (N_4131,N_3281,N_3866);
and U4132 (N_4132,N_3163,N_3270);
nor U4133 (N_4133,N_3807,N_3610);
or U4134 (N_4134,N_3754,N_3921);
xnor U4135 (N_4135,N_3026,N_3485);
xnor U4136 (N_4136,N_3744,N_3054);
or U4137 (N_4137,N_3431,N_3939);
and U4138 (N_4138,N_3615,N_3500);
and U4139 (N_4139,N_3589,N_3065);
nor U4140 (N_4140,N_3523,N_3064);
or U4141 (N_4141,N_3332,N_3531);
and U4142 (N_4142,N_3300,N_3434);
or U4143 (N_4143,N_3478,N_3931);
or U4144 (N_4144,N_3941,N_3288);
xnor U4145 (N_4145,N_3381,N_3952);
nor U4146 (N_4146,N_3250,N_3741);
and U4147 (N_4147,N_3033,N_3782);
or U4148 (N_4148,N_3405,N_3233);
and U4149 (N_4149,N_3092,N_3023);
nor U4150 (N_4150,N_3645,N_3948);
or U4151 (N_4151,N_3365,N_3796);
and U4152 (N_4152,N_3239,N_3747);
nor U4153 (N_4153,N_3704,N_3539);
nor U4154 (N_4154,N_3386,N_3541);
or U4155 (N_4155,N_3081,N_3960);
nand U4156 (N_4156,N_3740,N_3547);
and U4157 (N_4157,N_3231,N_3708);
nand U4158 (N_4158,N_3655,N_3734);
xor U4159 (N_4159,N_3117,N_3301);
or U4160 (N_4160,N_3086,N_3540);
nor U4161 (N_4161,N_3564,N_3339);
nor U4162 (N_4162,N_3219,N_3840);
and U4163 (N_4163,N_3298,N_3094);
and U4164 (N_4164,N_3994,N_3036);
and U4165 (N_4165,N_3317,N_3954);
nand U4166 (N_4166,N_3171,N_3631);
nand U4167 (N_4167,N_3983,N_3356);
nand U4168 (N_4168,N_3678,N_3982);
or U4169 (N_4169,N_3089,N_3487);
and U4170 (N_4170,N_3804,N_3504);
and U4171 (N_4171,N_3012,N_3703);
nor U4172 (N_4172,N_3769,N_3519);
or U4173 (N_4173,N_3553,N_3580);
xnor U4174 (N_4174,N_3475,N_3650);
xnor U4175 (N_4175,N_3695,N_3355);
or U4176 (N_4176,N_3723,N_3187);
nand U4177 (N_4177,N_3729,N_3410);
and U4178 (N_4178,N_3020,N_3858);
and U4179 (N_4179,N_3575,N_3412);
and U4180 (N_4180,N_3509,N_3460);
and U4181 (N_4181,N_3433,N_3652);
nand U4182 (N_4182,N_3972,N_3196);
nor U4183 (N_4183,N_3353,N_3123);
nor U4184 (N_4184,N_3986,N_3133);
and U4185 (N_4185,N_3872,N_3068);
and U4186 (N_4186,N_3202,N_3004);
or U4187 (N_4187,N_3070,N_3375);
nand U4188 (N_4188,N_3922,N_3612);
nor U4189 (N_4189,N_3686,N_3973);
or U4190 (N_4190,N_3147,N_3525);
nor U4191 (N_4191,N_3216,N_3088);
xor U4192 (N_4192,N_3189,N_3844);
or U4193 (N_4193,N_3532,N_3602);
or U4194 (N_4194,N_3335,N_3498);
nand U4195 (N_4195,N_3805,N_3644);
and U4196 (N_4196,N_3456,N_3588);
or U4197 (N_4197,N_3299,N_3041);
or U4198 (N_4198,N_3479,N_3031);
and U4199 (N_4199,N_3661,N_3028);
and U4200 (N_4200,N_3713,N_3204);
or U4201 (N_4201,N_3018,N_3966);
or U4202 (N_4202,N_3794,N_3551);
nand U4203 (N_4203,N_3046,N_3097);
nor U4204 (N_4204,N_3397,N_3413);
xor U4205 (N_4205,N_3200,N_3087);
xor U4206 (N_4206,N_3874,N_3042);
or U4207 (N_4207,N_3359,N_3181);
or U4208 (N_4208,N_3502,N_3980);
nand U4209 (N_4209,N_3730,N_3398);
or U4210 (N_4210,N_3705,N_3950);
and U4211 (N_4211,N_3153,N_3920);
and U4212 (N_4212,N_3030,N_3227);
or U4213 (N_4213,N_3185,N_3774);
or U4214 (N_4214,N_3481,N_3742);
xnor U4215 (N_4215,N_3358,N_3620);
and U4216 (N_4216,N_3336,N_3455);
or U4217 (N_4217,N_3305,N_3178);
nand U4218 (N_4218,N_3124,N_3340);
nor U4219 (N_4219,N_3373,N_3786);
or U4220 (N_4220,N_3257,N_3022);
nor U4221 (N_4221,N_3882,N_3913);
or U4222 (N_4222,N_3795,N_3013);
xor U4223 (N_4223,N_3311,N_3684);
nand U4224 (N_4224,N_3369,N_3442);
xor U4225 (N_4225,N_3622,N_3561);
and U4226 (N_4226,N_3380,N_3597);
xnor U4227 (N_4227,N_3881,N_3115);
or U4228 (N_4228,N_3164,N_3706);
nand U4229 (N_4229,N_3925,N_3797);
or U4230 (N_4230,N_3047,N_3486);
nand U4231 (N_4231,N_3766,N_3696);
or U4232 (N_4232,N_3617,N_3179);
xor U4233 (N_4233,N_3497,N_3530);
nor U4234 (N_4234,N_3918,N_3849);
nor U4235 (N_4235,N_3112,N_3506);
nor U4236 (N_4236,N_3120,N_3669);
and U4237 (N_4237,N_3331,N_3240);
or U4238 (N_4238,N_3430,N_3625);
and U4239 (N_4239,N_3977,N_3748);
nor U4240 (N_4240,N_3073,N_3029);
or U4241 (N_4241,N_3790,N_3834);
nor U4242 (N_4242,N_3482,N_3852);
nand U4243 (N_4243,N_3208,N_3032);
and U4244 (N_4244,N_3129,N_3282);
and U4245 (N_4245,N_3417,N_3524);
nor U4246 (N_4246,N_3702,N_3603);
nor U4247 (N_4247,N_3546,N_3828);
or U4248 (N_4248,N_3400,N_3897);
nor U4249 (N_4249,N_3628,N_3568);
nor U4250 (N_4250,N_3508,N_3987);
nor U4251 (N_4251,N_3995,N_3394);
nor U4252 (N_4252,N_3414,N_3272);
nor U4253 (N_4253,N_3290,N_3701);
nor U4254 (N_4254,N_3957,N_3513);
or U4255 (N_4255,N_3726,N_3908);
and U4256 (N_4256,N_3423,N_3383);
or U4257 (N_4257,N_3694,N_3452);
nand U4258 (N_4258,N_3969,N_3011);
nor U4259 (N_4259,N_3384,N_3878);
nand U4260 (N_4260,N_3222,N_3415);
xnor U4261 (N_4261,N_3832,N_3102);
nand U4262 (N_4262,N_3899,N_3772);
and U4263 (N_4263,N_3449,N_3228);
or U4264 (N_4264,N_3458,N_3511);
and U4265 (N_4265,N_3098,N_3266);
nand U4266 (N_4266,N_3149,N_3407);
nand U4267 (N_4267,N_3157,N_3940);
or U4268 (N_4268,N_3773,N_3071);
nand U4269 (N_4269,N_3718,N_3342);
nor U4270 (N_4270,N_3435,N_3075);
and U4271 (N_4271,N_3074,N_3821);
xor U4272 (N_4272,N_3888,N_3871);
nor U4273 (N_4273,N_3330,N_3116);
nand U4274 (N_4274,N_3006,N_3059);
nor U4275 (N_4275,N_3159,N_3675);
nand U4276 (N_4276,N_3167,N_3906);
or U4277 (N_4277,N_3277,N_3314);
nor U4278 (N_4278,N_3903,N_3810);
and U4279 (N_4279,N_3422,N_3674);
nand U4280 (N_4280,N_3630,N_3554);
and U4281 (N_4281,N_3051,N_3457);
nand U4282 (N_4282,N_3108,N_3341);
nand U4283 (N_4283,N_3308,N_3777);
nand U4284 (N_4284,N_3287,N_3946);
or U4285 (N_4285,N_3416,N_3214);
or U4286 (N_4286,N_3056,N_3963);
nor U4287 (N_4287,N_3390,N_3472);
nor U4288 (N_4288,N_3535,N_3321);
nor U4289 (N_4289,N_3867,N_3447);
and U4290 (N_4290,N_3285,N_3700);
nand U4291 (N_4291,N_3895,N_3111);
xor U4292 (N_4292,N_3595,N_3911);
nand U4293 (N_4293,N_3637,N_3904);
nand U4294 (N_4294,N_3943,N_3016);
nand U4295 (N_4295,N_3193,N_3648);
or U4296 (N_4296,N_3853,N_3639);
xor U4297 (N_4297,N_3854,N_3382);
nor U4298 (N_4298,N_3927,N_3591);
nor U4299 (N_4299,N_3249,N_3593);
or U4300 (N_4300,N_3635,N_3166);
nor U4301 (N_4301,N_3372,N_3091);
nand U4302 (N_4302,N_3154,N_3968);
and U4303 (N_4303,N_3443,N_3014);
and U4304 (N_4304,N_3061,N_3910);
or U4305 (N_4305,N_3192,N_3096);
nor U4306 (N_4306,N_3079,N_3312);
or U4307 (N_4307,N_3760,N_3981);
or U4308 (N_4308,N_3182,N_3846);
nand U4309 (N_4309,N_3893,N_3984);
nor U4310 (N_4310,N_3812,N_3638);
or U4311 (N_4311,N_3247,N_3083);
nor U4312 (N_4312,N_3429,N_3156);
and U4313 (N_4313,N_3641,N_3621);
or U4314 (N_4314,N_3293,N_3276);
or U4315 (N_4315,N_3771,N_3885);
nand U4316 (N_4316,N_3145,N_3264);
nand U4317 (N_4317,N_3090,N_3310);
or U4318 (N_4318,N_3604,N_3759);
nand U4319 (N_4319,N_3802,N_3681);
and U4320 (N_4320,N_3428,N_3732);
xor U4321 (N_4321,N_3545,N_3132);
xor U4322 (N_4322,N_3757,N_3211);
or U4323 (N_4323,N_3320,N_3780);
nor U4324 (N_4324,N_3344,N_3177);
or U4325 (N_4325,N_3002,N_3488);
nand U4326 (N_4326,N_3399,N_3727);
nor U4327 (N_4327,N_3752,N_3629);
or U4328 (N_4328,N_3492,N_3861);
or U4329 (N_4329,N_3712,N_3565);
nor U4330 (N_4330,N_3905,N_3687);
nor U4331 (N_4331,N_3512,N_3378);
or U4332 (N_4332,N_3158,N_3465);
nand U4333 (N_4333,N_3245,N_3914);
xnor U4334 (N_4334,N_3151,N_3229);
and U4335 (N_4335,N_3253,N_3689);
nor U4336 (N_4336,N_3101,N_3783);
nand U4337 (N_4337,N_3548,N_3409);
and U4338 (N_4338,N_3538,N_3190);
nor U4339 (N_4339,N_3784,N_3224);
and U4340 (N_4340,N_3444,N_3894);
xor U4341 (N_4341,N_3912,N_3053);
and U4342 (N_4342,N_3258,N_3830);
or U4343 (N_4343,N_3820,N_3401);
or U4344 (N_4344,N_3217,N_3521);
and U4345 (N_4345,N_3599,N_3377);
xnor U4346 (N_4346,N_3010,N_3060);
or U4347 (N_4347,N_3225,N_3392);
nand U4348 (N_4348,N_3304,N_3490);
nor U4349 (N_4349,N_3040,N_3831);
nand U4350 (N_4350,N_3819,N_3722);
nor U4351 (N_4351,N_3670,N_3212);
or U4352 (N_4352,N_3527,N_3302);
nor U4353 (N_4353,N_3476,N_3896);
xor U4354 (N_4354,N_3436,N_3890);
and U4355 (N_4355,N_3613,N_3021);
and U4356 (N_4356,N_3907,N_3529);
nand U4357 (N_4357,N_3841,N_3919);
and U4358 (N_4358,N_3316,N_3749);
nand U4359 (N_4359,N_3537,N_3550);
and U4360 (N_4360,N_3162,N_3606);
or U4361 (N_4361,N_3338,N_3693);
and U4362 (N_4362,N_3724,N_3876);
and U4363 (N_4363,N_3313,N_3001);
nand U4364 (N_4364,N_3965,N_3107);
xnor U4365 (N_4365,N_3719,N_3889);
nor U4366 (N_4366,N_3916,N_3668);
or U4367 (N_4367,N_3917,N_3720);
and U4368 (N_4368,N_3242,N_3560);
nor U4369 (N_4369,N_3975,N_3533);
or U4370 (N_4370,N_3528,N_3526);
and U4371 (N_4371,N_3514,N_3393);
nand U4372 (N_4372,N_3069,N_3932);
nor U4373 (N_4373,N_3891,N_3000);
nand U4374 (N_4374,N_3955,N_3471);
or U4375 (N_4375,N_3324,N_3839);
nor U4376 (N_4376,N_3197,N_3563);
nor U4377 (N_4377,N_3367,N_3273);
xnor U4378 (N_4378,N_3647,N_3663);
nor U4379 (N_4379,N_3027,N_3817);
nor U4380 (N_4380,N_3746,N_3201);
nor U4381 (N_4381,N_3803,N_3396);
or U4382 (N_4382,N_3213,N_3799);
xor U4383 (N_4383,N_3942,N_3283);
or U4384 (N_4384,N_3019,N_3174);
xor U4385 (N_4385,N_3015,N_3448);
nand U4386 (N_4386,N_3577,N_3349);
nor U4387 (N_4387,N_3348,N_3793);
and U4388 (N_4388,N_3244,N_3624);
or U4389 (N_4389,N_3619,N_3576);
nand U4390 (N_4390,N_3370,N_3295);
nor U4391 (N_4391,N_3735,N_3411);
and U4392 (N_4392,N_3184,N_3651);
or U4393 (N_4393,N_3756,N_3206);
and U4394 (N_4394,N_3127,N_3260);
and U4395 (N_4395,N_3768,N_3558);
nand U4396 (N_4396,N_3262,N_3778);
nor U4397 (N_4397,N_3555,N_3050);
nor U4398 (N_4398,N_3924,N_3665);
nor U4399 (N_4399,N_3750,N_3573);
xnor U4400 (N_4400,N_3672,N_3099);
nor U4401 (N_4401,N_3368,N_3717);
nor U4402 (N_4402,N_3677,N_3360);
and U4403 (N_4403,N_3350,N_3243);
and U4404 (N_4404,N_3697,N_3343);
or U4405 (N_4405,N_3292,N_3510);
or U4406 (N_4406,N_3590,N_3169);
or U4407 (N_4407,N_3207,N_3792);
nor U4408 (N_4408,N_3329,N_3119);
or U4409 (N_4409,N_3856,N_3901);
nor U4410 (N_4410,N_3676,N_3938);
and U4411 (N_4411,N_3085,N_3728);
xnor U4412 (N_4412,N_3286,N_3279);
nand U4413 (N_4413,N_3003,N_3869);
or U4414 (N_4414,N_3307,N_3974);
nor U4415 (N_4415,N_3048,N_3374);
nand U4416 (N_4416,N_3743,N_3570);
nand U4417 (N_4417,N_3762,N_3489);
nand U4418 (N_4418,N_3408,N_3579);
nor U4419 (N_4419,N_3562,N_3751);
or U4420 (N_4420,N_3785,N_3659);
nand U4421 (N_4421,N_3886,N_3062);
nand U4422 (N_4422,N_3632,N_3194);
nor U4423 (N_4423,N_3195,N_3660);
xnor U4424 (N_4424,N_3520,N_3271);
nand U4425 (N_4425,N_3814,N_3319);
and U4426 (N_4426,N_3148,N_3366);
and U4427 (N_4427,N_3664,N_3829);
xor U4428 (N_4428,N_3607,N_3884);
or U4429 (N_4429,N_3425,N_3835);
nor U4430 (N_4430,N_3322,N_3997);
and U4431 (N_4431,N_3767,N_3144);
and U4432 (N_4432,N_3930,N_3594);
or U4433 (N_4433,N_3445,N_3843);
and U4434 (N_4434,N_3325,N_3084);
and U4435 (N_4435,N_3851,N_3223);
nand U4436 (N_4436,N_3667,N_3855);
nor U4437 (N_4437,N_3556,N_3731);
nor U4438 (N_4438,N_3642,N_3711);
or U4439 (N_4439,N_3961,N_3566);
or U4440 (N_4440,N_3765,N_3483);
and U4441 (N_4441,N_3657,N_3306);
nand U4442 (N_4442,N_3536,N_3816);
or U4443 (N_4443,N_3406,N_3892);
nor U4444 (N_4444,N_3234,N_3870);
nor U4445 (N_4445,N_3863,N_3459);
or U4446 (N_4446,N_3709,N_3462);
or U4447 (N_4447,N_3274,N_3357);
xor U4448 (N_4448,N_3255,N_3764);
nand U4449 (N_4449,N_3666,N_3024);
xor U4450 (N_4450,N_3865,N_3654);
nand U4451 (N_4451,N_3900,N_3818);
or U4452 (N_4452,N_3923,N_3608);
nand U4453 (N_4453,N_3811,N_3009);
xor U4454 (N_4454,N_3501,N_3470);
nor U4455 (N_4455,N_3474,N_3441);
nand U4456 (N_4456,N_3847,N_3118);
or U4457 (N_4457,N_3592,N_3495);
xor U4458 (N_4458,N_3614,N_3883);
nor U4459 (N_4459,N_3569,N_3707);
nor U4460 (N_4460,N_3427,N_3136);
xor U4461 (N_4461,N_3636,N_3315);
xnor U4462 (N_4462,N_3875,N_3466);
nand U4463 (N_4463,N_3887,N_3049);
nand U4464 (N_4464,N_3949,N_3582);
nand U4465 (N_4465,N_3173,N_3699);
nand U4466 (N_4466,N_3309,N_3653);
xor U4467 (N_4467,N_3055,N_3618);
nand U4468 (N_4468,N_3135,N_3714);
and U4469 (N_4469,N_3035,N_3673);
xnor U4470 (N_4470,N_3935,N_3534);
xor U4471 (N_4471,N_3845,N_3688);
or U4472 (N_4472,N_3991,N_3220);
or U4473 (N_4473,N_3958,N_3106);
or U4474 (N_4474,N_3809,N_3827);
and U4475 (N_4475,N_3438,N_3453);
or U4476 (N_4476,N_3646,N_3066);
nor U4477 (N_4477,N_3230,N_3480);
nand U4478 (N_4478,N_3584,N_3626);
nand U4479 (N_4479,N_3402,N_3337);
or U4480 (N_4480,N_3172,N_3183);
nor U4481 (N_4481,N_3733,N_3252);
or U4482 (N_4482,N_3806,N_3755);
and U4483 (N_4483,N_3813,N_3104);
or U4484 (N_4484,N_3826,N_3110);
nand U4485 (N_4485,N_3685,N_3557);
or U4486 (N_4486,N_3926,N_3601);
xnor U4487 (N_4487,N_3542,N_3371);
or U4488 (N_4488,N_3463,N_3976);
nand U4489 (N_4489,N_3419,N_3076);
or U4490 (N_4490,N_3933,N_3057);
and U4491 (N_4491,N_3800,N_3585);
nand U4492 (N_4492,N_3461,N_3758);
nor U4493 (N_4493,N_3822,N_3574);
nand U4494 (N_4494,N_3798,N_3505);
nand U4495 (N_4495,N_3139,N_3186);
nand U4496 (N_4496,N_3945,N_3898);
and U4497 (N_4497,N_3507,N_3284);
or U4498 (N_4498,N_3572,N_3477);
nand U4499 (N_4499,N_3859,N_3067);
or U4500 (N_4500,N_3096,N_3514);
and U4501 (N_4501,N_3990,N_3122);
nor U4502 (N_4502,N_3176,N_3682);
or U4503 (N_4503,N_3547,N_3031);
nor U4504 (N_4504,N_3149,N_3329);
and U4505 (N_4505,N_3189,N_3929);
nor U4506 (N_4506,N_3192,N_3844);
and U4507 (N_4507,N_3133,N_3672);
nor U4508 (N_4508,N_3389,N_3277);
and U4509 (N_4509,N_3195,N_3078);
or U4510 (N_4510,N_3357,N_3792);
and U4511 (N_4511,N_3582,N_3291);
nand U4512 (N_4512,N_3328,N_3023);
or U4513 (N_4513,N_3293,N_3348);
or U4514 (N_4514,N_3709,N_3455);
and U4515 (N_4515,N_3454,N_3612);
nor U4516 (N_4516,N_3020,N_3140);
nor U4517 (N_4517,N_3985,N_3593);
nor U4518 (N_4518,N_3779,N_3370);
or U4519 (N_4519,N_3192,N_3399);
and U4520 (N_4520,N_3636,N_3471);
and U4521 (N_4521,N_3766,N_3212);
nor U4522 (N_4522,N_3428,N_3241);
and U4523 (N_4523,N_3855,N_3574);
or U4524 (N_4524,N_3365,N_3582);
nand U4525 (N_4525,N_3212,N_3498);
nand U4526 (N_4526,N_3756,N_3279);
nor U4527 (N_4527,N_3341,N_3019);
or U4528 (N_4528,N_3208,N_3104);
or U4529 (N_4529,N_3938,N_3921);
and U4530 (N_4530,N_3714,N_3615);
nor U4531 (N_4531,N_3989,N_3997);
nor U4532 (N_4532,N_3933,N_3950);
nor U4533 (N_4533,N_3636,N_3434);
nand U4534 (N_4534,N_3622,N_3103);
nor U4535 (N_4535,N_3171,N_3225);
or U4536 (N_4536,N_3312,N_3371);
or U4537 (N_4537,N_3215,N_3483);
nand U4538 (N_4538,N_3320,N_3594);
nor U4539 (N_4539,N_3168,N_3038);
nand U4540 (N_4540,N_3076,N_3129);
nor U4541 (N_4541,N_3414,N_3286);
and U4542 (N_4542,N_3931,N_3572);
and U4543 (N_4543,N_3344,N_3053);
xor U4544 (N_4544,N_3594,N_3056);
or U4545 (N_4545,N_3846,N_3339);
nand U4546 (N_4546,N_3911,N_3138);
nor U4547 (N_4547,N_3839,N_3622);
or U4548 (N_4548,N_3021,N_3593);
and U4549 (N_4549,N_3836,N_3670);
xor U4550 (N_4550,N_3177,N_3053);
and U4551 (N_4551,N_3667,N_3265);
and U4552 (N_4552,N_3036,N_3356);
and U4553 (N_4553,N_3381,N_3375);
and U4554 (N_4554,N_3991,N_3922);
or U4555 (N_4555,N_3974,N_3202);
and U4556 (N_4556,N_3878,N_3589);
or U4557 (N_4557,N_3594,N_3879);
nor U4558 (N_4558,N_3205,N_3274);
nand U4559 (N_4559,N_3902,N_3764);
and U4560 (N_4560,N_3372,N_3358);
or U4561 (N_4561,N_3268,N_3354);
nor U4562 (N_4562,N_3389,N_3316);
and U4563 (N_4563,N_3328,N_3710);
nand U4564 (N_4564,N_3685,N_3282);
nand U4565 (N_4565,N_3241,N_3478);
or U4566 (N_4566,N_3168,N_3021);
nor U4567 (N_4567,N_3416,N_3138);
xor U4568 (N_4568,N_3792,N_3870);
nand U4569 (N_4569,N_3375,N_3800);
or U4570 (N_4570,N_3850,N_3985);
nor U4571 (N_4571,N_3962,N_3730);
and U4572 (N_4572,N_3215,N_3085);
nor U4573 (N_4573,N_3639,N_3764);
and U4574 (N_4574,N_3294,N_3556);
and U4575 (N_4575,N_3860,N_3835);
nor U4576 (N_4576,N_3301,N_3276);
and U4577 (N_4577,N_3227,N_3627);
or U4578 (N_4578,N_3766,N_3878);
or U4579 (N_4579,N_3317,N_3376);
or U4580 (N_4580,N_3889,N_3835);
nand U4581 (N_4581,N_3222,N_3488);
nor U4582 (N_4582,N_3470,N_3474);
and U4583 (N_4583,N_3430,N_3814);
nand U4584 (N_4584,N_3252,N_3827);
nand U4585 (N_4585,N_3798,N_3523);
and U4586 (N_4586,N_3344,N_3201);
nand U4587 (N_4587,N_3806,N_3868);
nor U4588 (N_4588,N_3555,N_3137);
or U4589 (N_4589,N_3985,N_3040);
nand U4590 (N_4590,N_3287,N_3783);
or U4591 (N_4591,N_3651,N_3805);
xnor U4592 (N_4592,N_3533,N_3347);
xor U4593 (N_4593,N_3082,N_3479);
and U4594 (N_4594,N_3256,N_3656);
nor U4595 (N_4595,N_3880,N_3084);
nand U4596 (N_4596,N_3711,N_3103);
nand U4597 (N_4597,N_3304,N_3307);
nand U4598 (N_4598,N_3602,N_3825);
and U4599 (N_4599,N_3080,N_3802);
nor U4600 (N_4600,N_3406,N_3803);
nand U4601 (N_4601,N_3189,N_3390);
nor U4602 (N_4602,N_3753,N_3653);
and U4603 (N_4603,N_3672,N_3922);
nand U4604 (N_4604,N_3046,N_3767);
or U4605 (N_4605,N_3001,N_3770);
nor U4606 (N_4606,N_3619,N_3314);
xnor U4607 (N_4607,N_3445,N_3327);
or U4608 (N_4608,N_3671,N_3922);
and U4609 (N_4609,N_3762,N_3681);
nor U4610 (N_4610,N_3119,N_3437);
and U4611 (N_4611,N_3733,N_3773);
or U4612 (N_4612,N_3441,N_3511);
xor U4613 (N_4613,N_3854,N_3380);
or U4614 (N_4614,N_3931,N_3766);
nor U4615 (N_4615,N_3899,N_3775);
and U4616 (N_4616,N_3473,N_3506);
nor U4617 (N_4617,N_3187,N_3453);
or U4618 (N_4618,N_3191,N_3002);
and U4619 (N_4619,N_3127,N_3137);
and U4620 (N_4620,N_3969,N_3337);
nand U4621 (N_4621,N_3017,N_3873);
and U4622 (N_4622,N_3340,N_3964);
and U4623 (N_4623,N_3560,N_3322);
and U4624 (N_4624,N_3173,N_3337);
xnor U4625 (N_4625,N_3504,N_3509);
nor U4626 (N_4626,N_3310,N_3428);
xnor U4627 (N_4627,N_3425,N_3490);
or U4628 (N_4628,N_3614,N_3780);
nand U4629 (N_4629,N_3553,N_3452);
nor U4630 (N_4630,N_3365,N_3529);
nor U4631 (N_4631,N_3826,N_3698);
nand U4632 (N_4632,N_3080,N_3156);
nand U4633 (N_4633,N_3126,N_3862);
xnor U4634 (N_4634,N_3209,N_3169);
or U4635 (N_4635,N_3015,N_3939);
xnor U4636 (N_4636,N_3592,N_3729);
nor U4637 (N_4637,N_3691,N_3917);
nor U4638 (N_4638,N_3277,N_3285);
and U4639 (N_4639,N_3928,N_3875);
and U4640 (N_4640,N_3198,N_3007);
and U4641 (N_4641,N_3110,N_3589);
xnor U4642 (N_4642,N_3818,N_3821);
and U4643 (N_4643,N_3047,N_3895);
nand U4644 (N_4644,N_3645,N_3733);
nand U4645 (N_4645,N_3069,N_3474);
or U4646 (N_4646,N_3723,N_3411);
or U4647 (N_4647,N_3808,N_3528);
and U4648 (N_4648,N_3853,N_3063);
nand U4649 (N_4649,N_3799,N_3663);
nor U4650 (N_4650,N_3492,N_3513);
xor U4651 (N_4651,N_3473,N_3923);
nand U4652 (N_4652,N_3276,N_3999);
xnor U4653 (N_4653,N_3315,N_3651);
and U4654 (N_4654,N_3752,N_3295);
nor U4655 (N_4655,N_3033,N_3590);
nand U4656 (N_4656,N_3081,N_3615);
or U4657 (N_4657,N_3746,N_3477);
or U4658 (N_4658,N_3890,N_3715);
nand U4659 (N_4659,N_3430,N_3992);
nand U4660 (N_4660,N_3663,N_3279);
or U4661 (N_4661,N_3925,N_3649);
or U4662 (N_4662,N_3981,N_3468);
or U4663 (N_4663,N_3493,N_3696);
xnor U4664 (N_4664,N_3238,N_3801);
nor U4665 (N_4665,N_3005,N_3634);
xnor U4666 (N_4666,N_3732,N_3538);
or U4667 (N_4667,N_3384,N_3035);
or U4668 (N_4668,N_3089,N_3874);
or U4669 (N_4669,N_3683,N_3895);
or U4670 (N_4670,N_3552,N_3975);
nor U4671 (N_4671,N_3187,N_3263);
nand U4672 (N_4672,N_3502,N_3742);
nand U4673 (N_4673,N_3658,N_3643);
nand U4674 (N_4674,N_3356,N_3234);
or U4675 (N_4675,N_3265,N_3933);
xor U4676 (N_4676,N_3616,N_3282);
nor U4677 (N_4677,N_3907,N_3720);
nor U4678 (N_4678,N_3537,N_3829);
and U4679 (N_4679,N_3042,N_3132);
or U4680 (N_4680,N_3159,N_3888);
nand U4681 (N_4681,N_3653,N_3858);
xnor U4682 (N_4682,N_3319,N_3444);
and U4683 (N_4683,N_3780,N_3659);
nand U4684 (N_4684,N_3655,N_3451);
xnor U4685 (N_4685,N_3596,N_3466);
nand U4686 (N_4686,N_3232,N_3823);
and U4687 (N_4687,N_3169,N_3971);
or U4688 (N_4688,N_3324,N_3175);
or U4689 (N_4689,N_3461,N_3588);
nor U4690 (N_4690,N_3068,N_3552);
and U4691 (N_4691,N_3435,N_3999);
nor U4692 (N_4692,N_3328,N_3991);
or U4693 (N_4693,N_3649,N_3094);
nor U4694 (N_4694,N_3863,N_3568);
xnor U4695 (N_4695,N_3667,N_3619);
xor U4696 (N_4696,N_3096,N_3870);
xor U4697 (N_4697,N_3732,N_3093);
nor U4698 (N_4698,N_3835,N_3562);
xnor U4699 (N_4699,N_3317,N_3314);
or U4700 (N_4700,N_3497,N_3683);
and U4701 (N_4701,N_3225,N_3916);
or U4702 (N_4702,N_3361,N_3194);
or U4703 (N_4703,N_3738,N_3162);
nor U4704 (N_4704,N_3009,N_3395);
nand U4705 (N_4705,N_3390,N_3972);
nand U4706 (N_4706,N_3084,N_3286);
nor U4707 (N_4707,N_3893,N_3005);
nand U4708 (N_4708,N_3082,N_3898);
nand U4709 (N_4709,N_3600,N_3717);
nand U4710 (N_4710,N_3856,N_3979);
nor U4711 (N_4711,N_3587,N_3401);
xor U4712 (N_4712,N_3887,N_3272);
and U4713 (N_4713,N_3816,N_3772);
nor U4714 (N_4714,N_3437,N_3978);
and U4715 (N_4715,N_3357,N_3715);
and U4716 (N_4716,N_3477,N_3580);
nand U4717 (N_4717,N_3378,N_3613);
or U4718 (N_4718,N_3839,N_3717);
nand U4719 (N_4719,N_3683,N_3322);
and U4720 (N_4720,N_3260,N_3816);
nor U4721 (N_4721,N_3578,N_3502);
or U4722 (N_4722,N_3093,N_3246);
and U4723 (N_4723,N_3333,N_3434);
or U4724 (N_4724,N_3787,N_3986);
xnor U4725 (N_4725,N_3802,N_3331);
and U4726 (N_4726,N_3658,N_3353);
or U4727 (N_4727,N_3726,N_3862);
or U4728 (N_4728,N_3929,N_3064);
and U4729 (N_4729,N_3309,N_3796);
and U4730 (N_4730,N_3125,N_3266);
xor U4731 (N_4731,N_3095,N_3234);
nand U4732 (N_4732,N_3098,N_3898);
and U4733 (N_4733,N_3027,N_3907);
xor U4734 (N_4734,N_3536,N_3651);
or U4735 (N_4735,N_3595,N_3106);
and U4736 (N_4736,N_3195,N_3020);
and U4737 (N_4737,N_3213,N_3025);
nor U4738 (N_4738,N_3950,N_3720);
xor U4739 (N_4739,N_3841,N_3055);
nand U4740 (N_4740,N_3533,N_3715);
nor U4741 (N_4741,N_3045,N_3997);
nand U4742 (N_4742,N_3325,N_3893);
or U4743 (N_4743,N_3124,N_3439);
nand U4744 (N_4744,N_3374,N_3706);
or U4745 (N_4745,N_3414,N_3437);
nand U4746 (N_4746,N_3884,N_3566);
nand U4747 (N_4747,N_3867,N_3507);
nor U4748 (N_4748,N_3602,N_3696);
and U4749 (N_4749,N_3658,N_3600);
or U4750 (N_4750,N_3995,N_3048);
xor U4751 (N_4751,N_3418,N_3511);
nand U4752 (N_4752,N_3243,N_3088);
nand U4753 (N_4753,N_3810,N_3150);
or U4754 (N_4754,N_3092,N_3854);
xnor U4755 (N_4755,N_3820,N_3499);
or U4756 (N_4756,N_3441,N_3425);
xor U4757 (N_4757,N_3598,N_3724);
nor U4758 (N_4758,N_3802,N_3695);
and U4759 (N_4759,N_3429,N_3498);
and U4760 (N_4760,N_3794,N_3890);
and U4761 (N_4761,N_3692,N_3062);
and U4762 (N_4762,N_3494,N_3901);
nor U4763 (N_4763,N_3657,N_3709);
or U4764 (N_4764,N_3925,N_3296);
xnor U4765 (N_4765,N_3168,N_3476);
nor U4766 (N_4766,N_3367,N_3688);
or U4767 (N_4767,N_3574,N_3609);
and U4768 (N_4768,N_3289,N_3169);
nand U4769 (N_4769,N_3857,N_3956);
nand U4770 (N_4770,N_3764,N_3214);
xnor U4771 (N_4771,N_3529,N_3253);
and U4772 (N_4772,N_3253,N_3452);
nand U4773 (N_4773,N_3829,N_3497);
nand U4774 (N_4774,N_3144,N_3156);
or U4775 (N_4775,N_3406,N_3790);
and U4776 (N_4776,N_3601,N_3227);
and U4777 (N_4777,N_3837,N_3942);
nand U4778 (N_4778,N_3057,N_3405);
nor U4779 (N_4779,N_3047,N_3698);
nor U4780 (N_4780,N_3025,N_3303);
nor U4781 (N_4781,N_3367,N_3583);
and U4782 (N_4782,N_3944,N_3270);
nor U4783 (N_4783,N_3867,N_3395);
or U4784 (N_4784,N_3696,N_3801);
and U4785 (N_4785,N_3343,N_3916);
and U4786 (N_4786,N_3416,N_3030);
or U4787 (N_4787,N_3239,N_3289);
nor U4788 (N_4788,N_3578,N_3623);
or U4789 (N_4789,N_3709,N_3330);
nand U4790 (N_4790,N_3519,N_3974);
and U4791 (N_4791,N_3860,N_3693);
and U4792 (N_4792,N_3346,N_3434);
nand U4793 (N_4793,N_3650,N_3357);
nand U4794 (N_4794,N_3171,N_3667);
or U4795 (N_4795,N_3315,N_3583);
nand U4796 (N_4796,N_3944,N_3161);
nand U4797 (N_4797,N_3311,N_3715);
and U4798 (N_4798,N_3261,N_3373);
and U4799 (N_4799,N_3774,N_3286);
or U4800 (N_4800,N_3126,N_3527);
nand U4801 (N_4801,N_3178,N_3249);
nor U4802 (N_4802,N_3652,N_3337);
nor U4803 (N_4803,N_3245,N_3325);
nor U4804 (N_4804,N_3913,N_3721);
nor U4805 (N_4805,N_3348,N_3562);
xnor U4806 (N_4806,N_3025,N_3247);
and U4807 (N_4807,N_3066,N_3597);
or U4808 (N_4808,N_3397,N_3859);
and U4809 (N_4809,N_3952,N_3096);
nand U4810 (N_4810,N_3204,N_3164);
and U4811 (N_4811,N_3733,N_3894);
nor U4812 (N_4812,N_3896,N_3806);
nand U4813 (N_4813,N_3415,N_3243);
nor U4814 (N_4814,N_3811,N_3561);
xor U4815 (N_4815,N_3838,N_3785);
nor U4816 (N_4816,N_3896,N_3270);
nor U4817 (N_4817,N_3492,N_3977);
nor U4818 (N_4818,N_3849,N_3784);
nor U4819 (N_4819,N_3469,N_3110);
nor U4820 (N_4820,N_3621,N_3832);
and U4821 (N_4821,N_3200,N_3110);
nand U4822 (N_4822,N_3633,N_3750);
xor U4823 (N_4823,N_3979,N_3271);
and U4824 (N_4824,N_3111,N_3257);
xnor U4825 (N_4825,N_3880,N_3086);
xnor U4826 (N_4826,N_3412,N_3037);
or U4827 (N_4827,N_3444,N_3663);
and U4828 (N_4828,N_3518,N_3069);
nor U4829 (N_4829,N_3563,N_3870);
xnor U4830 (N_4830,N_3776,N_3577);
xor U4831 (N_4831,N_3040,N_3961);
nand U4832 (N_4832,N_3721,N_3937);
nor U4833 (N_4833,N_3482,N_3524);
nand U4834 (N_4834,N_3368,N_3079);
nand U4835 (N_4835,N_3110,N_3094);
and U4836 (N_4836,N_3333,N_3525);
or U4837 (N_4837,N_3481,N_3058);
or U4838 (N_4838,N_3915,N_3200);
nor U4839 (N_4839,N_3012,N_3076);
or U4840 (N_4840,N_3822,N_3748);
nand U4841 (N_4841,N_3589,N_3052);
or U4842 (N_4842,N_3970,N_3337);
and U4843 (N_4843,N_3276,N_3881);
nor U4844 (N_4844,N_3446,N_3767);
xnor U4845 (N_4845,N_3287,N_3833);
xnor U4846 (N_4846,N_3182,N_3588);
nand U4847 (N_4847,N_3725,N_3069);
nand U4848 (N_4848,N_3825,N_3199);
and U4849 (N_4849,N_3629,N_3774);
or U4850 (N_4850,N_3235,N_3024);
or U4851 (N_4851,N_3598,N_3817);
or U4852 (N_4852,N_3154,N_3013);
nor U4853 (N_4853,N_3784,N_3109);
or U4854 (N_4854,N_3566,N_3460);
or U4855 (N_4855,N_3224,N_3948);
and U4856 (N_4856,N_3319,N_3816);
nor U4857 (N_4857,N_3123,N_3483);
or U4858 (N_4858,N_3607,N_3569);
nor U4859 (N_4859,N_3949,N_3740);
nand U4860 (N_4860,N_3238,N_3557);
nand U4861 (N_4861,N_3390,N_3572);
xor U4862 (N_4862,N_3310,N_3615);
nand U4863 (N_4863,N_3353,N_3668);
and U4864 (N_4864,N_3440,N_3293);
nand U4865 (N_4865,N_3028,N_3660);
or U4866 (N_4866,N_3726,N_3675);
nand U4867 (N_4867,N_3257,N_3083);
nand U4868 (N_4868,N_3556,N_3167);
or U4869 (N_4869,N_3804,N_3254);
and U4870 (N_4870,N_3538,N_3678);
nor U4871 (N_4871,N_3278,N_3074);
and U4872 (N_4872,N_3478,N_3895);
nor U4873 (N_4873,N_3158,N_3114);
nand U4874 (N_4874,N_3255,N_3278);
nand U4875 (N_4875,N_3999,N_3173);
nor U4876 (N_4876,N_3644,N_3652);
nand U4877 (N_4877,N_3268,N_3110);
nand U4878 (N_4878,N_3237,N_3003);
and U4879 (N_4879,N_3248,N_3245);
nand U4880 (N_4880,N_3542,N_3610);
nor U4881 (N_4881,N_3233,N_3250);
nor U4882 (N_4882,N_3535,N_3376);
xor U4883 (N_4883,N_3951,N_3708);
xnor U4884 (N_4884,N_3325,N_3702);
nand U4885 (N_4885,N_3080,N_3643);
nand U4886 (N_4886,N_3376,N_3493);
and U4887 (N_4887,N_3759,N_3124);
nand U4888 (N_4888,N_3734,N_3871);
nand U4889 (N_4889,N_3714,N_3566);
or U4890 (N_4890,N_3797,N_3627);
and U4891 (N_4891,N_3445,N_3242);
xnor U4892 (N_4892,N_3263,N_3936);
and U4893 (N_4893,N_3621,N_3803);
nand U4894 (N_4894,N_3625,N_3953);
nor U4895 (N_4895,N_3256,N_3257);
or U4896 (N_4896,N_3894,N_3861);
or U4897 (N_4897,N_3293,N_3671);
or U4898 (N_4898,N_3980,N_3569);
xor U4899 (N_4899,N_3014,N_3572);
and U4900 (N_4900,N_3279,N_3197);
or U4901 (N_4901,N_3722,N_3105);
nor U4902 (N_4902,N_3904,N_3885);
xor U4903 (N_4903,N_3166,N_3920);
nor U4904 (N_4904,N_3725,N_3852);
and U4905 (N_4905,N_3984,N_3268);
or U4906 (N_4906,N_3891,N_3231);
and U4907 (N_4907,N_3201,N_3648);
or U4908 (N_4908,N_3438,N_3395);
nand U4909 (N_4909,N_3444,N_3255);
or U4910 (N_4910,N_3112,N_3299);
or U4911 (N_4911,N_3534,N_3715);
and U4912 (N_4912,N_3353,N_3294);
nor U4913 (N_4913,N_3761,N_3557);
nand U4914 (N_4914,N_3543,N_3256);
nand U4915 (N_4915,N_3797,N_3333);
nor U4916 (N_4916,N_3064,N_3280);
nor U4917 (N_4917,N_3598,N_3260);
or U4918 (N_4918,N_3639,N_3631);
nand U4919 (N_4919,N_3877,N_3557);
nor U4920 (N_4920,N_3848,N_3155);
and U4921 (N_4921,N_3696,N_3175);
nor U4922 (N_4922,N_3017,N_3338);
and U4923 (N_4923,N_3950,N_3458);
nor U4924 (N_4924,N_3972,N_3367);
or U4925 (N_4925,N_3399,N_3803);
nor U4926 (N_4926,N_3704,N_3668);
and U4927 (N_4927,N_3740,N_3750);
nand U4928 (N_4928,N_3494,N_3975);
and U4929 (N_4929,N_3919,N_3866);
nor U4930 (N_4930,N_3597,N_3177);
and U4931 (N_4931,N_3212,N_3649);
and U4932 (N_4932,N_3211,N_3443);
and U4933 (N_4933,N_3081,N_3455);
nor U4934 (N_4934,N_3039,N_3603);
nand U4935 (N_4935,N_3736,N_3475);
and U4936 (N_4936,N_3953,N_3719);
nor U4937 (N_4937,N_3148,N_3980);
and U4938 (N_4938,N_3206,N_3396);
nand U4939 (N_4939,N_3611,N_3396);
and U4940 (N_4940,N_3437,N_3256);
or U4941 (N_4941,N_3665,N_3883);
nor U4942 (N_4942,N_3065,N_3128);
or U4943 (N_4943,N_3319,N_3650);
nand U4944 (N_4944,N_3486,N_3561);
and U4945 (N_4945,N_3368,N_3989);
nand U4946 (N_4946,N_3329,N_3917);
or U4947 (N_4947,N_3556,N_3911);
xnor U4948 (N_4948,N_3427,N_3823);
and U4949 (N_4949,N_3682,N_3698);
or U4950 (N_4950,N_3163,N_3709);
or U4951 (N_4951,N_3649,N_3792);
nand U4952 (N_4952,N_3768,N_3527);
xnor U4953 (N_4953,N_3376,N_3974);
and U4954 (N_4954,N_3728,N_3511);
nand U4955 (N_4955,N_3981,N_3927);
nand U4956 (N_4956,N_3178,N_3225);
and U4957 (N_4957,N_3859,N_3005);
nand U4958 (N_4958,N_3841,N_3342);
and U4959 (N_4959,N_3564,N_3793);
and U4960 (N_4960,N_3079,N_3241);
or U4961 (N_4961,N_3803,N_3160);
or U4962 (N_4962,N_3604,N_3986);
nor U4963 (N_4963,N_3798,N_3231);
nor U4964 (N_4964,N_3376,N_3775);
or U4965 (N_4965,N_3484,N_3535);
nor U4966 (N_4966,N_3557,N_3172);
or U4967 (N_4967,N_3502,N_3919);
nand U4968 (N_4968,N_3067,N_3564);
or U4969 (N_4969,N_3168,N_3846);
nand U4970 (N_4970,N_3316,N_3705);
or U4971 (N_4971,N_3330,N_3241);
or U4972 (N_4972,N_3835,N_3994);
nor U4973 (N_4973,N_3993,N_3494);
and U4974 (N_4974,N_3335,N_3386);
and U4975 (N_4975,N_3864,N_3104);
nor U4976 (N_4976,N_3792,N_3877);
xor U4977 (N_4977,N_3811,N_3319);
or U4978 (N_4978,N_3439,N_3180);
nand U4979 (N_4979,N_3176,N_3071);
nor U4980 (N_4980,N_3956,N_3130);
and U4981 (N_4981,N_3264,N_3370);
and U4982 (N_4982,N_3315,N_3290);
nor U4983 (N_4983,N_3740,N_3326);
and U4984 (N_4984,N_3035,N_3571);
or U4985 (N_4985,N_3807,N_3891);
xor U4986 (N_4986,N_3280,N_3617);
nor U4987 (N_4987,N_3948,N_3790);
nand U4988 (N_4988,N_3136,N_3367);
or U4989 (N_4989,N_3670,N_3663);
nand U4990 (N_4990,N_3946,N_3522);
nand U4991 (N_4991,N_3007,N_3995);
nand U4992 (N_4992,N_3239,N_3710);
xnor U4993 (N_4993,N_3364,N_3509);
and U4994 (N_4994,N_3485,N_3010);
xor U4995 (N_4995,N_3971,N_3087);
or U4996 (N_4996,N_3237,N_3946);
or U4997 (N_4997,N_3507,N_3996);
and U4998 (N_4998,N_3633,N_3392);
nor U4999 (N_4999,N_3211,N_3484);
and U5000 (N_5000,N_4414,N_4587);
xor U5001 (N_5001,N_4114,N_4123);
nor U5002 (N_5002,N_4629,N_4199);
nand U5003 (N_5003,N_4084,N_4944);
nand U5004 (N_5004,N_4265,N_4525);
nand U5005 (N_5005,N_4167,N_4656);
nand U5006 (N_5006,N_4027,N_4095);
or U5007 (N_5007,N_4788,N_4166);
nand U5008 (N_5008,N_4042,N_4277);
nor U5009 (N_5009,N_4344,N_4563);
or U5010 (N_5010,N_4016,N_4336);
or U5011 (N_5011,N_4007,N_4418);
or U5012 (N_5012,N_4013,N_4040);
or U5013 (N_5013,N_4358,N_4744);
nor U5014 (N_5014,N_4469,N_4380);
nand U5015 (N_5015,N_4334,N_4090);
and U5016 (N_5016,N_4004,N_4710);
nand U5017 (N_5017,N_4507,N_4850);
and U5018 (N_5018,N_4684,N_4567);
or U5019 (N_5019,N_4089,N_4172);
xor U5020 (N_5020,N_4538,N_4562);
nand U5021 (N_5021,N_4153,N_4681);
or U5022 (N_5022,N_4993,N_4868);
nor U5023 (N_5023,N_4620,N_4981);
or U5024 (N_5024,N_4733,N_4717);
nor U5025 (N_5025,N_4489,N_4616);
nand U5026 (N_5026,N_4386,N_4124);
or U5027 (N_5027,N_4861,N_4400);
xor U5028 (N_5028,N_4964,N_4832);
nand U5029 (N_5029,N_4399,N_4663);
and U5030 (N_5030,N_4549,N_4564);
nand U5031 (N_5031,N_4916,N_4192);
and U5032 (N_5032,N_4838,N_4962);
nand U5033 (N_5033,N_4028,N_4648);
nand U5034 (N_5034,N_4240,N_4968);
xor U5035 (N_5035,N_4643,N_4310);
xor U5036 (N_5036,N_4354,N_4059);
and U5037 (N_5037,N_4675,N_4104);
or U5038 (N_5038,N_4522,N_4718);
or U5039 (N_5039,N_4446,N_4983);
and U5040 (N_5040,N_4075,N_4355);
and U5041 (N_5041,N_4256,N_4992);
or U5042 (N_5042,N_4572,N_4390);
and U5043 (N_5043,N_4700,N_4820);
nor U5044 (N_5044,N_4660,N_4513);
and U5045 (N_5045,N_4279,N_4426);
nand U5046 (N_5046,N_4257,N_4133);
nand U5047 (N_5047,N_4096,N_4183);
nor U5048 (N_5048,N_4917,N_4568);
nand U5049 (N_5049,N_4571,N_4438);
nand U5050 (N_5050,N_4707,N_4407);
or U5051 (N_5051,N_4829,N_4597);
nand U5052 (N_5052,N_4320,N_4604);
and U5053 (N_5053,N_4932,N_4102);
and U5054 (N_5054,N_4530,N_4703);
xor U5055 (N_5055,N_4085,N_4594);
nor U5056 (N_5056,N_4436,N_4593);
or U5057 (N_5057,N_4125,N_4029);
or U5058 (N_5058,N_4931,N_4792);
nand U5059 (N_5059,N_4553,N_4851);
nor U5060 (N_5060,N_4254,N_4785);
xor U5061 (N_5061,N_4221,N_4099);
nand U5062 (N_5062,N_4582,N_4268);
nand U5063 (N_5063,N_4348,N_4319);
nor U5064 (N_5064,N_4904,N_4026);
xor U5065 (N_5065,N_4126,N_4071);
nand U5066 (N_5066,N_4985,N_4152);
nor U5067 (N_5067,N_4474,N_4791);
nor U5068 (N_5068,N_4934,N_4428);
xnor U5069 (N_5069,N_4275,N_4840);
and U5070 (N_5070,N_4862,N_4466);
or U5071 (N_5071,N_4592,N_4843);
nand U5072 (N_5072,N_4163,N_4139);
xnor U5073 (N_5073,N_4999,N_4662);
nand U5074 (N_5074,N_4248,N_4384);
and U5075 (N_5075,N_4879,N_4309);
nand U5076 (N_5076,N_4488,N_4858);
and U5077 (N_5077,N_4869,N_4633);
nand U5078 (N_5078,N_4803,N_4006);
nand U5079 (N_5079,N_4494,N_4263);
nor U5080 (N_5080,N_4994,N_4154);
or U5081 (N_5081,N_4613,N_4450);
or U5082 (N_5082,N_4367,N_4671);
and U5083 (N_5083,N_4545,N_4502);
xnor U5084 (N_5084,N_4989,N_4280);
and U5085 (N_5085,N_4766,N_4382);
or U5086 (N_5086,N_4619,N_4634);
xor U5087 (N_5087,N_4919,N_4325);
xnor U5088 (N_5088,N_4860,N_4548);
or U5089 (N_5089,N_4383,N_4923);
xnor U5090 (N_5090,N_4778,N_4335);
nand U5091 (N_5091,N_4231,N_4926);
nand U5092 (N_5092,N_4030,N_4272);
and U5093 (N_5093,N_4212,N_4053);
nand U5094 (N_5094,N_4284,N_4481);
nand U5095 (N_5095,N_4159,N_4433);
and U5096 (N_5096,N_4782,N_4060);
nor U5097 (N_5097,N_4039,N_4458);
xor U5098 (N_5098,N_4852,N_4554);
and U5099 (N_5099,N_4537,N_4796);
nor U5100 (N_5100,N_4485,N_4132);
nor U5101 (N_5101,N_4500,N_4512);
and U5102 (N_5102,N_4511,N_4445);
or U5103 (N_5103,N_4155,N_4287);
xnor U5104 (N_5104,N_4323,N_4245);
nor U5105 (N_5105,N_4264,N_4061);
xor U5106 (N_5106,N_4559,N_4291);
or U5107 (N_5107,N_4602,N_4241);
and U5108 (N_5108,N_4779,N_4189);
and U5109 (N_5109,N_4317,N_4503);
nand U5110 (N_5110,N_4833,N_4201);
nor U5111 (N_5111,N_4297,N_4252);
or U5112 (N_5112,N_4417,N_4824);
xor U5113 (N_5113,N_4520,N_4220);
xnor U5114 (N_5114,N_4088,N_4091);
nand U5115 (N_5115,N_4557,N_4118);
and U5116 (N_5116,N_4420,N_4455);
nor U5117 (N_5117,N_4872,N_4895);
and U5118 (N_5118,N_4025,N_4746);
and U5119 (N_5119,N_4398,N_4213);
and U5120 (N_5120,N_4750,N_4521);
or U5121 (N_5121,N_4726,N_4610);
nor U5122 (N_5122,N_4262,N_4326);
and U5123 (N_5123,N_4242,N_4544);
nor U5124 (N_5124,N_4122,N_4765);
and U5125 (N_5125,N_4115,N_4516);
and U5126 (N_5126,N_4531,N_4614);
xor U5127 (N_5127,N_4706,N_4724);
nor U5128 (N_5128,N_4318,N_4366);
nand U5129 (N_5129,N_4546,N_4757);
nand U5130 (N_5130,N_4631,N_4289);
nand U5131 (N_5131,N_4477,N_4533);
and U5132 (N_5132,N_4641,N_4147);
or U5133 (N_5133,N_4036,N_4292);
or U5134 (N_5134,N_4041,N_4207);
and U5135 (N_5135,N_4644,N_4471);
and U5136 (N_5136,N_4294,N_4158);
nor U5137 (N_5137,N_4807,N_4727);
or U5138 (N_5138,N_4627,N_4915);
nor U5139 (N_5139,N_4801,N_4736);
or U5140 (N_5140,N_4055,N_4575);
and U5141 (N_5141,N_4628,N_4731);
and U5142 (N_5142,N_4689,N_4527);
nor U5143 (N_5143,N_4753,N_4924);
and U5144 (N_5144,N_4001,N_4774);
nor U5145 (N_5145,N_4720,N_4835);
nand U5146 (N_5146,N_4959,N_4768);
and U5147 (N_5147,N_4705,N_4223);
nor U5148 (N_5148,N_4307,N_4704);
or U5149 (N_5149,N_4342,N_4312);
or U5150 (N_5150,N_4170,N_4187);
or U5151 (N_5151,N_4422,N_4215);
nand U5152 (N_5152,N_4585,N_4330);
nor U5153 (N_5153,N_4800,N_4010);
xnor U5154 (N_5154,N_4440,N_4939);
or U5155 (N_5155,N_4772,N_4712);
nor U5156 (N_5156,N_4763,N_4077);
nand U5157 (N_5157,N_4745,N_4285);
or U5158 (N_5158,N_4211,N_4022);
and U5159 (N_5159,N_4480,N_4823);
or U5160 (N_5160,N_4427,N_4760);
or U5161 (N_5161,N_4106,N_4682);
or U5162 (N_5162,N_4699,N_4729);
nor U5163 (N_5163,N_4035,N_4176);
or U5164 (N_5164,N_4854,N_4160);
nor U5165 (N_5165,N_4395,N_4866);
xnor U5166 (N_5166,N_4584,N_4044);
and U5167 (N_5167,N_4083,N_4739);
nor U5168 (N_5168,N_4863,N_4711);
or U5169 (N_5169,N_4429,N_4119);
nor U5170 (N_5170,N_4270,N_4814);
or U5171 (N_5171,N_4877,N_4408);
and U5172 (N_5172,N_4460,N_4020);
nor U5173 (N_5173,N_4519,N_4828);
nand U5174 (N_5174,N_4658,N_4441);
nand U5175 (N_5175,N_4178,N_4459);
or U5176 (N_5176,N_4974,N_4579);
xor U5177 (N_5177,N_4638,N_4056);
or U5178 (N_5178,N_4299,N_4749);
or U5179 (N_5179,N_4808,N_4817);
and U5180 (N_5180,N_4659,N_4526);
and U5181 (N_5181,N_4278,N_4045);
xnor U5182 (N_5182,N_4327,N_4691);
xnor U5183 (N_5183,N_4424,N_4551);
and U5184 (N_5184,N_4667,N_4702);
nand U5185 (N_5185,N_4595,N_4135);
xnor U5186 (N_5186,N_4352,N_4886);
or U5187 (N_5187,N_4899,N_4226);
or U5188 (N_5188,N_4157,N_4177);
nor U5189 (N_5189,N_4887,N_4875);
xor U5190 (N_5190,N_4723,N_4343);
and U5191 (N_5191,N_4234,N_4642);
or U5192 (N_5192,N_4680,N_4698);
nand U5193 (N_5193,N_4161,N_4837);
or U5194 (N_5194,N_4435,N_4903);
nor U5195 (N_5195,N_4908,N_4473);
nor U5196 (N_5196,N_4518,N_4885);
nand U5197 (N_5197,N_4721,N_4936);
nand U5198 (N_5198,N_4990,N_4871);
nor U5199 (N_5199,N_4216,N_4586);
and U5200 (N_5200,N_4371,N_4009);
and U5201 (N_5201,N_4821,N_4809);
or U5202 (N_5202,N_4333,N_4708);
nand U5203 (N_5203,N_4110,N_4797);
nor U5204 (N_5204,N_4849,N_4515);
or U5205 (N_5205,N_4905,N_4973);
or U5206 (N_5206,N_4780,N_4880);
xor U5207 (N_5207,N_4900,N_4410);
nand U5208 (N_5208,N_4364,N_4332);
nand U5209 (N_5209,N_4014,N_4227);
or U5210 (N_5210,N_4079,N_4238);
nand U5211 (N_5211,N_4784,N_4623);
nor U5212 (N_5212,N_4997,N_4661);
or U5213 (N_5213,N_4305,N_4543);
xor U5214 (N_5214,N_4457,N_4933);
and U5215 (N_5215,N_4491,N_4912);
nand U5216 (N_5216,N_4173,N_4984);
nor U5217 (N_5217,N_4506,N_4771);
xor U5218 (N_5218,N_4683,N_4755);
nand U5219 (N_5219,N_4425,N_4884);
nor U5220 (N_5220,N_4074,N_4730);
and U5221 (N_5221,N_4070,N_4492);
or U5222 (N_5222,N_4058,N_4037);
nand U5223 (N_5223,N_4190,N_4372);
nand U5224 (N_5224,N_4709,N_4409);
nor U5225 (N_5225,N_4467,N_4093);
or U5226 (N_5226,N_4783,N_4393);
nor U5227 (N_5227,N_4635,N_4253);
nand U5228 (N_5228,N_4735,N_4751);
or U5229 (N_5229,N_4969,N_4302);
and U5230 (N_5230,N_4787,N_4357);
nand U5231 (N_5231,N_4909,N_4370);
nor U5232 (N_5232,N_4472,N_4558);
or U5233 (N_5233,N_4756,N_4977);
or U5234 (N_5234,N_4589,N_4636);
nand U5235 (N_5235,N_4591,N_4970);
and U5236 (N_5236,N_4573,N_4376);
nor U5237 (N_5237,N_4770,N_4113);
nand U5238 (N_5238,N_4054,N_4087);
and U5239 (N_5239,N_4368,N_4385);
xor U5240 (N_5240,N_4921,N_4047);
or U5241 (N_5241,N_4836,N_4165);
nor U5242 (N_5242,N_4444,N_4722);
or U5243 (N_5243,N_4987,N_4949);
xor U5244 (N_5244,N_4151,N_4963);
or U5245 (N_5245,N_4322,N_4448);
nor U5246 (N_5246,N_4164,N_4239);
nor U5247 (N_5247,N_4419,N_4387);
nand U5248 (N_5248,N_4894,N_4618);
nand U5249 (N_5249,N_4200,N_4011);
nand U5250 (N_5250,N_4678,N_4228);
and U5251 (N_5251,N_4465,N_4274);
nand U5252 (N_5252,N_4542,N_4626);
nand U5253 (N_5253,N_4742,N_4225);
nor U5254 (N_5254,N_4951,N_4646);
nand U5255 (N_5255,N_4986,N_4191);
xnor U5256 (N_5256,N_4615,N_4937);
nand U5257 (N_5257,N_4655,N_4078);
or U5258 (N_5258,N_4049,N_4209);
or U5259 (N_5259,N_4431,N_4224);
and U5260 (N_5260,N_4893,N_4068);
nand U5261 (N_5261,N_4134,N_4148);
nand U5262 (N_5262,N_4499,N_4108);
and U5263 (N_5263,N_4536,N_4504);
or U5264 (N_5264,N_4452,N_4498);
nand U5265 (N_5265,N_4605,N_4266);
nand U5266 (N_5266,N_4609,N_4954);
nor U5267 (N_5267,N_4131,N_4948);
and U5268 (N_5268,N_4217,N_4421);
xor U5269 (N_5269,N_4598,N_4972);
or U5270 (N_5270,N_4168,N_4901);
or U5271 (N_5271,N_4673,N_4975);
nand U5272 (N_5272,N_4063,N_4560);
or U5273 (N_5273,N_4048,N_4293);
nand U5274 (N_5274,N_4816,N_4066);
and U5275 (N_5275,N_4679,N_4960);
nor U5276 (N_5276,N_4958,N_4911);
nand U5277 (N_5277,N_4142,N_4625);
or U5278 (N_5278,N_4690,N_4490);
or U5279 (N_5279,N_4416,N_4830);
nor U5280 (N_5280,N_4381,N_4639);
nor U5281 (N_5281,N_4906,N_4946);
or U5282 (N_5282,N_4351,N_4486);
xnor U5283 (N_5283,N_4313,N_4574);
or U5284 (N_5284,N_4143,N_4128);
nor U5285 (N_5285,N_4100,N_4260);
or U5286 (N_5286,N_4094,N_4258);
nand U5287 (N_5287,N_4713,N_4107);
or U5288 (N_5288,N_4714,N_4940);
nor U5289 (N_5289,N_4847,N_4082);
nor U5290 (N_5290,N_4140,N_4453);
or U5291 (N_5291,N_4864,N_4261);
nor U5292 (N_5292,N_4012,N_4876);
nor U5293 (N_5293,N_4624,N_4222);
nor U5294 (N_5294,N_4464,N_4630);
nand U5295 (N_5295,N_4608,N_4961);
nand U5296 (N_5296,N_4867,N_4865);
nor U5297 (N_5297,N_4121,N_4194);
xnor U5298 (N_5298,N_4482,N_4813);
and U5299 (N_5299,N_4846,N_4651);
and U5300 (N_5300,N_4316,N_4449);
and U5301 (N_5301,N_4196,N_4423);
and U5302 (N_5302,N_4290,N_4581);
nand U5303 (N_5303,N_4738,N_4988);
nand U5304 (N_5304,N_4966,N_4182);
and U5305 (N_5305,N_4965,N_4758);
and U5306 (N_5306,N_4606,N_4583);
or U5307 (N_5307,N_4617,N_4237);
nand U5308 (N_5308,N_4632,N_4841);
nor U5309 (N_5309,N_4892,N_4669);
nand U5310 (N_5310,N_4031,N_4341);
or U5311 (N_5311,N_4415,N_4953);
xor U5312 (N_5312,N_4046,N_4654);
nor U5313 (N_5313,N_4672,N_4359);
nor U5314 (N_5314,N_4392,N_4184);
nand U5315 (N_5315,N_4080,N_4728);
nand U5316 (N_5316,N_4203,N_4373);
nand U5317 (N_5317,N_4645,N_4769);
nand U5318 (N_5318,N_4649,N_4794);
nand U5319 (N_5319,N_4017,N_4136);
nand U5320 (N_5320,N_4561,N_4127);
xnor U5321 (N_5321,N_4105,N_4790);
nand U5322 (N_5322,N_4269,N_4853);
or U5323 (N_5323,N_4532,N_4483);
nor U5324 (N_5324,N_4204,N_4478);
or U5325 (N_5325,N_4762,N_4913);
nor U5326 (N_5326,N_4795,N_4596);
xnor U5327 (N_5327,N_4379,N_4329);
nor U5328 (N_5328,N_4555,N_4839);
nand U5329 (N_5329,N_4556,N_4300);
or U5330 (N_5330,N_4767,N_4149);
xnor U5331 (N_5331,N_4112,N_4692);
or U5332 (N_5332,N_4405,N_4811);
or U5333 (N_5333,N_4411,N_4111);
nor U5334 (N_5334,N_4236,N_4799);
or U5335 (N_5335,N_4000,N_4514);
or U5336 (N_5336,N_4150,N_4185);
xnor U5337 (N_5337,N_4928,N_4621);
nand U5338 (N_5338,N_4650,N_4523);
nand U5339 (N_5339,N_4377,N_4338);
or U5340 (N_5340,N_4685,N_4505);
nor U5341 (N_5341,N_4676,N_4856);
and U5342 (N_5342,N_4073,N_4747);
nor U5343 (N_5343,N_4064,N_4952);
xnor U5344 (N_5344,N_4295,N_4834);
and U5345 (N_5345,N_4484,N_4777);
nor U5346 (N_5346,N_4324,N_4827);
nor U5347 (N_5347,N_4819,N_4812);
nand U5348 (N_5348,N_4759,N_4802);
and U5349 (N_5349,N_4288,N_4311);
or U5350 (N_5350,N_4804,N_4979);
nor U5351 (N_5351,N_4057,N_4374);
nand U5352 (N_5352,N_4144,N_4023);
and U5353 (N_5353,N_4789,N_4943);
nor U5354 (N_5354,N_4437,N_4547);
nand U5355 (N_5355,N_4391,N_4117);
and U5356 (N_5356,N_4806,N_4461);
xnor U5357 (N_5357,N_4076,N_4443);
nand U5358 (N_5358,N_4818,N_4198);
nand U5359 (N_5359,N_4942,N_4339);
xnor U5360 (N_5360,N_4249,N_4032);
nand U5361 (N_5361,N_4493,N_4998);
nand U5362 (N_5362,N_4668,N_4340);
nor U5363 (N_5363,N_4487,N_4888);
or U5364 (N_5364,N_4328,N_4463);
xnor U5365 (N_5365,N_4362,N_4517);
or U5366 (N_5366,N_4246,N_4403);
nor U5367 (N_5367,N_4695,N_4202);
nor U5368 (N_5368,N_4741,N_4171);
and U5369 (N_5369,N_4232,N_4052);
nand U5370 (N_5370,N_4980,N_4878);
nand U5371 (N_5371,N_4786,N_4550);
or U5372 (N_5372,N_4552,N_4565);
or U5373 (N_5373,N_4003,N_4306);
or U5374 (N_5374,N_4918,N_4622);
nand U5375 (N_5375,N_4496,N_4360);
xor U5376 (N_5376,N_4510,N_4857);
and U5377 (N_5377,N_4897,N_4848);
nor U5378 (N_5378,N_4761,N_4138);
nor U5379 (N_5379,N_4922,N_4267);
nor U5380 (N_5380,N_4401,N_4195);
or U5381 (N_5381,N_4902,N_4688);
nand U5382 (N_5382,N_4982,N_4971);
and U5383 (N_5383,N_4495,N_4101);
or U5384 (N_5384,N_4065,N_4219);
nor U5385 (N_5385,N_4693,N_4508);
nor U5386 (N_5386,N_4955,N_4501);
nor U5387 (N_5387,N_4967,N_4120);
xor U5388 (N_5388,N_4752,N_4337);
or U5389 (N_5389,N_4350,N_4179);
and U5390 (N_5390,N_4637,N_4413);
nor U5391 (N_5391,N_4890,N_4244);
nand U5392 (N_5392,N_4015,N_4652);
and U5393 (N_5393,N_4218,N_4434);
or U5394 (N_5394,N_4169,N_4375);
nand U5395 (N_5395,N_4298,N_4188);
xor U5396 (N_5396,N_4732,N_4208);
and U5397 (N_5397,N_4600,N_4541);
and U5398 (N_5398,N_4186,N_4397);
or U5399 (N_5399,N_4276,N_4855);
or U5400 (N_5400,N_4451,N_4910);
xor U5401 (N_5401,N_4051,N_4734);
nor U5402 (N_5402,N_4881,N_4725);
xnor U5403 (N_5403,N_4907,N_4378);
nor U5404 (N_5404,N_4024,N_4607);
or U5405 (N_5405,N_4303,N_4097);
and U5406 (N_5406,N_4038,N_4456);
nand U5407 (N_5407,N_4034,N_4396);
nand U5408 (N_5408,N_4976,N_4156);
and U5409 (N_5409,N_4920,N_4304);
or U5410 (N_5410,N_4109,N_4670);
or U5411 (N_5411,N_4315,N_4844);
xnor U5412 (N_5412,N_4773,N_4230);
and U5413 (N_5413,N_4406,N_4570);
and U5414 (N_5414,N_4369,N_4447);
or U5415 (N_5415,N_4798,N_4092);
nor U5416 (N_5416,N_4243,N_4308);
and U5417 (N_5417,N_4008,N_4273);
or U5418 (N_5418,N_4930,N_4412);
nand U5419 (N_5419,N_4137,N_4251);
nand U5420 (N_5420,N_4346,N_4402);
or U5421 (N_5421,N_4859,N_4590);
or U5422 (N_5422,N_4404,N_4896);
nor U5423 (N_5423,N_4021,N_4664);
nand U5424 (N_5424,N_4898,N_4611);
or U5425 (N_5425,N_4162,N_4540);
and U5426 (N_5426,N_4874,N_4181);
or U5427 (N_5427,N_4978,N_4229);
nand U5428 (N_5428,N_4282,N_4479);
nor U5429 (N_5429,N_4889,N_4439);
nor U5430 (N_5430,N_4210,N_4529);
or U5431 (N_5431,N_4180,N_4578);
nand U5432 (N_5432,N_4805,N_4193);
or U5433 (N_5433,N_4647,N_4314);
and U5434 (N_5434,N_4018,N_4640);
xor U5435 (N_5435,N_4995,N_4430);
xor U5436 (N_5436,N_4601,N_4259);
nor U5437 (N_5437,N_4891,N_4539);
and U5438 (N_5438,N_4737,N_4247);
and U5439 (N_5439,N_4043,N_4271);
and U5440 (N_5440,N_4941,N_4687);
nand U5441 (N_5441,N_4388,N_4842);
and U5442 (N_5442,N_4822,N_4764);
or U5443 (N_5443,N_4130,N_4255);
nand U5444 (N_5444,N_4033,N_4826);
and U5445 (N_5445,N_4103,N_4454);
nor U5446 (N_5446,N_4250,N_4653);
or U5447 (N_5447,N_4925,N_4141);
nand U5448 (N_5448,N_4086,N_4356);
nor U5449 (N_5449,N_4716,N_4283);
nand U5450 (N_5450,N_4442,N_4081);
xnor U5451 (N_5451,N_4098,N_4349);
nand U5452 (N_5452,N_4938,N_4947);
or U5453 (N_5453,N_4748,N_4365);
nand U5454 (N_5454,N_4286,N_4719);
or U5455 (N_5455,N_4476,N_4991);
or U5456 (N_5456,N_4067,N_4694);
and U5457 (N_5457,N_4588,N_4072);
nand U5458 (N_5458,N_4793,N_4580);
nor U5459 (N_5459,N_4657,N_4666);
and U5460 (N_5460,N_4870,N_4996);
and U5461 (N_5461,N_4686,N_4470);
nor U5462 (N_5462,N_4914,N_4882);
or U5463 (N_5463,N_4715,N_4005);
nor U5464 (N_5464,N_4363,N_4353);
nand U5465 (N_5465,N_4775,N_4815);
nor U5466 (N_5466,N_4296,N_4935);
nor U5467 (N_5467,N_4603,N_4781);
and U5468 (N_5468,N_4576,N_4497);
or U5469 (N_5469,N_4950,N_4831);
or U5470 (N_5470,N_4019,N_4612);
or U5471 (N_5471,N_4677,N_4599);
and U5472 (N_5472,N_4002,N_4776);
nand U5473 (N_5473,N_4740,N_4697);
and U5474 (N_5474,N_4345,N_4475);
and U5475 (N_5475,N_4534,N_4321);
and U5476 (N_5476,N_4394,N_4062);
xor U5477 (N_5477,N_4927,N_4674);
nor U5478 (N_5478,N_4214,N_4432);
nand U5479 (N_5479,N_4569,N_4524);
or U5480 (N_5480,N_4361,N_4175);
nand U5481 (N_5481,N_4929,N_4956);
or U5482 (N_5482,N_4389,N_4301);
nand U5483 (N_5483,N_4468,N_4050);
and U5484 (N_5484,N_4577,N_4825);
or U5485 (N_5485,N_4696,N_4462);
nor U5486 (N_5486,N_4743,N_4331);
or U5487 (N_5487,N_4281,N_4145);
nor U5488 (N_5488,N_4810,N_4528);
and U5489 (N_5489,N_4235,N_4754);
xor U5490 (N_5490,N_4347,N_4873);
or U5491 (N_5491,N_4509,N_4535);
and U5492 (N_5492,N_4206,N_4701);
nand U5493 (N_5493,N_4233,N_4883);
nor U5494 (N_5494,N_4665,N_4845);
nor U5495 (N_5495,N_4129,N_4116);
and U5496 (N_5496,N_4069,N_4945);
or U5497 (N_5497,N_4957,N_4197);
and U5498 (N_5498,N_4174,N_4205);
nand U5499 (N_5499,N_4146,N_4566);
or U5500 (N_5500,N_4060,N_4577);
or U5501 (N_5501,N_4540,N_4665);
xnor U5502 (N_5502,N_4398,N_4421);
nor U5503 (N_5503,N_4469,N_4199);
nor U5504 (N_5504,N_4600,N_4928);
and U5505 (N_5505,N_4587,N_4218);
nor U5506 (N_5506,N_4194,N_4566);
or U5507 (N_5507,N_4001,N_4296);
and U5508 (N_5508,N_4142,N_4410);
xnor U5509 (N_5509,N_4848,N_4984);
and U5510 (N_5510,N_4433,N_4383);
or U5511 (N_5511,N_4088,N_4812);
xor U5512 (N_5512,N_4764,N_4983);
or U5513 (N_5513,N_4758,N_4415);
nand U5514 (N_5514,N_4246,N_4755);
nand U5515 (N_5515,N_4187,N_4511);
or U5516 (N_5516,N_4327,N_4358);
and U5517 (N_5517,N_4076,N_4341);
nand U5518 (N_5518,N_4508,N_4728);
or U5519 (N_5519,N_4448,N_4212);
nand U5520 (N_5520,N_4580,N_4009);
and U5521 (N_5521,N_4576,N_4639);
and U5522 (N_5522,N_4382,N_4453);
and U5523 (N_5523,N_4429,N_4850);
and U5524 (N_5524,N_4180,N_4733);
xnor U5525 (N_5525,N_4905,N_4948);
or U5526 (N_5526,N_4667,N_4768);
and U5527 (N_5527,N_4313,N_4581);
or U5528 (N_5528,N_4956,N_4547);
nor U5529 (N_5529,N_4891,N_4941);
or U5530 (N_5530,N_4354,N_4242);
or U5531 (N_5531,N_4181,N_4187);
nand U5532 (N_5532,N_4508,N_4129);
nand U5533 (N_5533,N_4712,N_4604);
xor U5534 (N_5534,N_4762,N_4445);
nand U5535 (N_5535,N_4978,N_4439);
nor U5536 (N_5536,N_4112,N_4030);
nand U5537 (N_5537,N_4734,N_4759);
or U5538 (N_5538,N_4732,N_4850);
or U5539 (N_5539,N_4348,N_4592);
nand U5540 (N_5540,N_4956,N_4753);
nor U5541 (N_5541,N_4015,N_4298);
nor U5542 (N_5542,N_4309,N_4026);
nor U5543 (N_5543,N_4531,N_4249);
or U5544 (N_5544,N_4614,N_4660);
or U5545 (N_5545,N_4701,N_4108);
nor U5546 (N_5546,N_4018,N_4561);
nor U5547 (N_5547,N_4605,N_4257);
nand U5548 (N_5548,N_4342,N_4430);
nand U5549 (N_5549,N_4017,N_4163);
and U5550 (N_5550,N_4923,N_4366);
nand U5551 (N_5551,N_4364,N_4736);
or U5552 (N_5552,N_4003,N_4944);
xnor U5553 (N_5553,N_4417,N_4277);
nand U5554 (N_5554,N_4621,N_4635);
nor U5555 (N_5555,N_4885,N_4990);
xor U5556 (N_5556,N_4517,N_4050);
and U5557 (N_5557,N_4190,N_4664);
nand U5558 (N_5558,N_4528,N_4551);
nor U5559 (N_5559,N_4248,N_4173);
nand U5560 (N_5560,N_4577,N_4207);
and U5561 (N_5561,N_4545,N_4869);
xor U5562 (N_5562,N_4907,N_4399);
nor U5563 (N_5563,N_4538,N_4117);
nand U5564 (N_5564,N_4418,N_4495);
xnor U5565 (N_5565,N_4183,N_4739);
or U5566 (N_5566,N_4087,N_4179);
and U5567 (N_5567,N_4032,N_4585);
and U5568 (N_5568,N_4772,N_4569);
and U5569 (N_5569,N_4304,N_4641);
nand U5570 (N_5570,N_4704,N_4183);
nand U5571 (N_5571,N_4515,N_4465);
nand U5572 (N_5572,N_4178,N_4610);
and U5573 (N_5573,N_4484,N_4129);
nor U5574 (N_5574,N_4474,N_4547);
or U5575 (N_5575,N_4331,N_4528);
nand U5576 (N_5576,N_4029,N_4158);
or U5577 (N_5577,N_4774,N_4080);
nand U5578 (N_5578,N_4139,N_4475);
nor U5579 (N_5579,N_4208,N_4953);
nor U5580 (N_5580,N_4687,N_4957);
nor U5581 (N_5581,N_4599,N_4252);
nor U5582 (N_5582,N_4880,N_4193);
nand U5583 (N_5583,N_4872,N_4511);
and U5584 (N_5584,N_4483,N_4415);
xnor U5585 (N_5585,N_4251,N_4089);
nor U5586 (N_5586,N_4029,N_4186);
xnor U5587 (N_5587,N_4800,N_4327);
or U5588 (N_5588,N_4338,N_4455);
and U5589 (N_5589,N_4299,N_4088);
nor U5590 (N_5590,N_4593,N_4519);
and U5591 (N_5591,N_4237,N_4907);
nand U5592 (N_5592,N_4330,N_4599);
nand U5593 (N_5593,N_4783,N_4622);
and U5594 (N_5594,N_4232,N_4263);
and U5595 (N_5595,N_4209,N_4613);
nor U5596 (N_5596,N_4454,N_4284);
or U5597 (N_5597,N_4949,N_4249);
or U5598 (N_5598,N_4255,N_4320);
nand U5599 (N_5599,N_4094,N_4363);
nand U5600 (N_5600,N_4995,N_4583);
and U5601 (N_5601,N_4639,N_4890);
nand U5602 (N_5602,N_4349,N_4904);
or U5603 (N_5603,N_4756,N_4507);
nor U5604 (N_5604,N_4092,N_4265);
or U5605 (N_5605,N_4965,N_4917);
nand U5606 (N_5606,N_4359,N_4644);
nand U5607 (N_5607,N_4599,N_4424);
or U5608 (N_5608,N_4794,N_4480);
and U5609 (N_5609,N_4831,N_4238);
xor U5610 (N_5610,N_4392,N_4435);
and U5611 (N_5611,N_4191,N_4536);
nand U5612 (N_5612,N_4953,N_4600);
or U5613 (N_5613,N_4151,N_4087);
and U5614 (N_5614,N_4647,N_4211);
or U5615 (N_5615,N_4608,N_4178);
and U5616 (N_5616,N_4860,N_4534);
nand U5617 (N_5617,N_4929,N_4868);
xnor U5618 (N_5618,N_4967,N_4344);
nand U5619 (N_5619,N_4790,N_4816);
nand U5620 (N_5620,N_4829,N_4725);
or U5621 (N_5621,N_4437,N_4366);
xor U5622 (N_5622,N_4570,N_4471);
xor U5623 (N_5623,N_4441,N_4903);
nor U5624 (N_5624,N_4965,N_4191);
nand U5625 (N_5625,N_4534,N_4235);
and U5626 (N_5626,N_4160,N_4850);
nor U5627 (N_5627,N_4403,N_4667);
or U5628 (N_5628,N_4805,N_4636);
nor U5629 (N_5629,N_4683,N_4066);
nand U5630 (N_5630,N_4885,N_4323);
or U5631 (N_5631,N_4330,N_4683);
and U5632 (N_5632,N_4089,N_4173);
nor U5633 (N_5633,N_4310,N_4201);
or U5634 (N_5634,N_4371,N_4494);
or U5635 (N_5635,N_4675,N_4656);
or U5636 (N_5636,N_4105,N_4142);
nor U5637 (N_5637,N_4353,N_4064);
nor U5638 (N_5638,N_4995,N_4434);
or U5639 (N_5639,N_4945,N_4540);
nand U5640 (N_5640,N_4591,N_4263);
nand U5641 (N_5641,N_4972,N_4051);
nand U5642 (N_5642,N_4422,N_4181);
nand U5643 (N_5643,N_4855,N_4169);
nand U5644 (N_5644,N_4422,N_4289);
nor U5645 (N_5645,N_4422,N_4955);
nand U5646 (N_5646,N_4351,N_4997);
nor U5647 (N_5647,N_4654,N_4847);
or U5648 (N_5648,N_4869,N_4023);
nor U5649 (N_5649,N_4580,N_4977);
or U5650 (N_5650,N_4211,N_4962);
nand U5651 (N_5651,N_4895,N_4190);
or U5652 (N_5652,N_4877,N_4675);
and U5653 (N_5653,N_4251,N_4864);
nor U5654 (N_5654,N_4518,N_4380);
nor U5655 (N_5655,N_4043,N_4213);
nor U5656 (N_5656,N_4937,N_4494);
or U5657 (N_5657,N_4248,N_4174);
or U5658 (N_5658,N_4974,N_4632);
and U5659 (N_5659,N_4158,N_4500);
nor U5660 (N_5660,N_4394,N_4880);
xnor U5661 (N_5661,N_4517,N_4440);
and U5662 (N_5662,N_4266,N_4424);
or U5663 (N_5663,N_4789,N_4210);
nor U5664 (N_5664,N_4924,N_4459);
nand U5665 (N_5665,N_4153,N_4407);
nand U5666 (N_5666,N_4264,N_4187);
and U5667 (N_5667,N_4200,N_4230);
nand U5668 (N_5668,N_4508,N_4719);
nand U5669 (N_5669,N_4186,N_4966);
and U5670 (N_5670,N_4290,N_4302);
nor U5671 (N_5671,N_4304,N_4614);
nor U5672 (N_5672,N_4877,N_4224);
nor U5673 (N_5673,N_4925,N_4978);
or U5674 (N_5674,N_4498,N_4444);
nand U5675 (N_5675,N_4042,N_4512);
nor U5676 (N_5676,N_4116,N_4928);
and U5677 (N_5677,N_4515,N_4864);
and U5678 (N_5678,N_4292,N_4572);
nand U5679 (N_5679,N_4059,N_4857);
nor U5680 (N_5680,N_4790,N_4936);
nor U5681 (N_5681,N_4096,N_4746);
nand U5682 (N_5682,N_4324,N_4547);
and U5683 (N_5683,N_4895,N_4298);
nand U5684 (N_5684,N_4698,N_4886);
or U5685 (N_5685,N_4196,N_4335);
nor U5686 (N_5686,N_4942,N_4625);
or U5687 (N_5687,N_4575,N_4063);
nand U5688 (N_5688,N_4712,N_4244);
nand U5689 (N_5689,N_4523,N_4080);
or U5690 (N_5690,N_4805,N_4336);
or U5691 (N_5691,N_4471,N_4382);
and U5692 (N_5692,N_4072,N_4856);
xnor U5693 (N_5693,N_4092,N_4129);
nand U5694 (N_5694,N_4008,N_4826);
and U5695 (N_5695,N_4299,N_4527);
or U5696 (N_5696,N_4764,N_4515);
nor U5697 (N_5697,N_4321,N_4743);
or U5698 (N_5698,N_4879,N_4095);
nor U5699 (N_5699,N_4445,N_4723);
nand U5700 (N_5700,N_4941,N_4959);
nor U5701 (N_5701,N_4098,N_4839);
and U5702 (N_5702,N_4207,N_4029);
nand U5703 (N_5703,N_4347,N_4390);
nand U5704 (N_5704,N_4901,N_4810);
xor U5705 (N_5705,N_4025,N_4462);
xnor U5706 (N_5706,N_4905,N_4916);
xnor U5707 (N_5707,N_4022,N_4310);
nor U5708 (N_5708,N_4204,N_4290);
nor U5709 (N_5709,N_4400,N_4516);
or U5710 (N_5710,N_4761,N_4928);
or U5711 (N_5711,N_4728,N_4571);
and U5712 (N_5712,N_4746,N_4586);
nand U5713 (N_5713,N_4527,N_4870);
and U5714 (N_5714,N_4233,N_4929);
nor U5715 (N_5715,N_4798,N_4922);
nand U5716 (N_5716,N_4237,N_4456);
or U5717 (N_5717,N_4323,N_4434);
and U5718 (N_5718,N_4897,N_4019);
and U5719 (N_5719,N_4751,N_4440);
or U5720 (N_5720,N_4619,N_4316);
nor U5721 (N_5721,N_4348,N_4536);
or U5722 (N_5722,N_4339,N_4762);
nand U5723 (N_5723,N_4952,N_4268);
nor U5724 (N_5724,N_4527,N_4225);
or U5725 (N_5725,N_4602,N_4714);
and U5726 (N_5726,N_4158,N_4980);
xnor U5727 (N_5727,N_4840,N_4048);
nor U5728 (N_5728,N_4058,N_4290);
nand U5729 (N_5729,N_4935,N_4513);
nand U5730 (N_5730,N_4796,N_4358);
nor U5731 (N_5731,N_4631,N_4085);
or U5732 (N_5732,N_4318,N_4222);
and U5733 (N_5733,N_4103,N_4798);
and U5734 (N_5734,N_4589,N_4879);
and U5735 (N_5735,N_4222,N_4913);
or U5736 (N_5736,N_4081,N_4378);
or U5737 (N_5737,N_4956,N_4466);
or U5738 (N_5738,N_4660,N_4061);
or U5739 (N_5739,N_4115,N_4474);
nand U5740 (N_5740,N_4517,N_4584);
nor U5741 (N_5741,N_4120,N_4050);
xor U5742 (N_5742,N_4109,N_4193);
nor U5743 (N_5743,N_4389,N_4445);
and U5744 (N_5744,N_4473,N_4098);
nor U5745 (N_5745,N_4087,N_4824);
or U5746 (N_5746,N_4385,N_4286);
and U5747 (N_5747,N_4883,N_4591);
or U5748 (N_5748,N_4082,N_4783);
xor U5749 (N_5749,N_4307,N_4773);
xnor U5750 (N_5750,N_4180,N_4232);
and U5751 (N_5751,N_4035,N_4334);
xnor U5752 (N_5752,N_4840,N_4287);
nor U5753 (N_5753,N_4255,N_4315);
xnor U5754 (N_5754,N_4500,N_4115);
or U5755 (N_5755,N_4813,N_4650);
or U5756 (N_5756,N_4371,N_4518);
and U5757 (N_5757,N_4765,N_4552);
nand U5758 (N_5758,N_4445,N_4573);
and U5759 (N_5759,N_4616,N_4720);
nor U5760 (N_5760,N_4493,N_4207);
and U5761 (N_5761,N_4992,N_4855);
xnor U5762 (N_5762,N_4266,N_4916);
and U5763 (N_5763,N_4351,N_4772);
or U5764 (N_5764,N_4045,N_4844);
nand U5765 (N_5765,N_4353,N_4699);
or U5766 (N_5766,N_4886,N_4616);
nor U5767 (N_5767,N_4904,N_4318);
nand U5768 (N_5768,N_4209,N_4242);
nand U5769 (N_5769,N_4600,N_4635);
nor U5770 (N_5770,N_4732,N_4134);
or U5771 (N_5771,N_4935,N_4989);
nor U5772 (N_5772,N_4175,N_4979);
nor U5773 (N_5773,N_4050,N_4548);
nand U5774 (N_5774,N_4640,N_4914);
or U5775 (N_5775,N_4127,N_4435);
or U5776 (N_5776,N_4352,N_4326);
nand U5777 (N_5777,N_4376,N_4056);
nor U5778 (N_5778,N_4456,N_4159);
and U5779 (N_5779,N_4677,N_4216);
or U5780 (N_5780,N_4586,N_4697);
nor U5781 (N_5781,N_4866,N_4497);
nand U5782 (N_5782,N_4365,N_4700);
nand U5783 (N_5783,N_4487,N_4362);
and U5784 (N_5784,N_4669,N_4144);
xnor U5785 (N_5785,N_4093,N_4583);
or U5786 (N_5786,N_4042,N_4568);
nor U5787 (N_5787,N_4695,N_4973);
xnor U5788 (N_5788,N_4161,N_4644);
and U5789 (N_5789,N_4493,N_4190);
nor U5790 (N_5790,N_4382,N_4630);
and U5791 (N_5791,N_4989,N_4598);
nand U5792 (N_5792,N_4282,N_4135);
and U5793 (N_5793,N_4412,N_4249);
nand U5794 (N_5794,N_4229,N_4956);
or U5795 (N_5795,N_4945,N_4870);
and U5796 (N_5796,N_4181,N_4529);
and U5797 (N_5797,N_4796,N_4443);
nand U5798 (N_5798,N_4671,N_4774);
and U5799 (N_5799,N_4161,N_4304);
xnor U5800 (N_5800,N_4306,N_4180);
and U5801 (N_5801,N_4204,N_4702);
xor U5802 (N_5802,N_4688,N_4717);
or U5803 (N_5803,N_4940,N_4761);
nor U5804 (N_5804,N_4956,N_4000);
xnor U5805 (N_5805,N_4103,N_4295);
nor U5806 (N_5806,N_4255,N_4025);
nand U5807 (N_5807,N_4175,N_4878);
nand U5808 (N_5808,N_4428,N_4453);
and U5809 (N_5809,N_4323,N_4471);
nor U5810 (N_5810,N_4437,N_4781);
nand U5811 (N_5811,N_4336,N_4892);
and U5812 (N_5812,N_4402,N_4551);
nor U5813 (N_5813,N_4925,N_4951);
or U5814 (N_5814,N_4819,N_4041);
and U5815 (N_5815,N_4175,N_4343);
nor U5816 (N_5816,N_4410,N_4166);
and U5817 (N_5817,N_4531,N_4220);
nor U5818 (N_5818,N_4872,N_4517);
nand U5819 (N_5819,N_4681,N_4262);
nand U5820 (N_5820,N_4992,N_4589);
nor U5821 (N_5821,N_4635,N_4323);
and U5822 (N_5822,N_4816,N_4192);
or U5823 (N_5823,N_4080,N_4906);
nand U5824 (N_5824,N_4156,N_4839);
nor U5825 (N_5825,N_4044,N_4694);
xor U5826 (N_5826,N_4536,N_4637);
nand U5827 (N_5827,N_4055,N_4047);
nor U5828 (N_5828,N_4431,N_4128);
nand U5829 (N_5829,N_4357,N_4947);
nand U5830 (N_5830,N_4252,N_4115);
or U5831 (N_5831,N_4404,N_4685);
and U5832 (N_5832,N_4531,N_4412);
and U5833 (N_5833,N_4877,N_4762);
nand U5834 (N_5834,N_4391,N_4598);
or U5835 (N_5835,N_4935,N_4954);
or U5836 (N_5836,N_4777,N_4278);
nor U5837 (N_5837,N_4255,N_4679);
and U5838 (N_5838,N_4926,N_4839);
nor U5839 (N_5839,N_4556,N_4856);
and U5840 (N_5840,N_4519,N_4763);
nor U5841 (N_5841,N_4005,N_4544);
nor U5842 (N_5842,N_4696,N_4750);
and U5843 (N_5843,N_4942,N_4535);
or U5844 (N_5844,N_4410,N_4941);
nor U5845 (N_5845,N_4668,N_4242);
or U5846 (N_5846,N_4143,N_4290);
and U5847 (N_5847,N_4572,N_4432);
or U5848 (N_5848,N_4830,N_4194);
nand U5849 (N_5849,N_4687,N_4139);
nor U5850 (N_5850,N_4975,N_4103);
and U5851 (N_5851,N_4566,N_4243);
or U5852 (N_5852,N_4024,N_4696);
and U5853 (N_5853,N_4667,N_4512);
xor U5854 (N_5854,N_4519,N_4620);
nor U5855 (N_5855,N_4800,N_4048);
xor U5856 (N_5856,N_4827,N_4392);
nor U5857 (N_5857,N_4966,N_4454);
or U5858 (N_5858,N_4515,N_4253);
or U5859 (N_5859,N_4583,N_4597);
or U5860 (N_5860,N_4986,N_4979);
nand U5861 (N_5861,N_4005,N_4810);
nor U5862 (N_5862,N_4788,N_4635);
nor U5863 (N_5863,N_4002,N_4833);
or U5864 (N_5864,N_4250,N_4272);
nand U5865 (N_5865,N_4195,N_4734);
and U5866 (N_5866,N_4185,N_4764);
nor U5867 (N_5867,N_4604,N_4929);
or U5868 (N_5868,N_4957,N_4287);
and U5869 (N_5869,N_4229,N_4260);
nor U5870 (N_5870,N_4153,N_4067);
and U5871 (N_5871,N_4510,N_4224);
xnor U5872 (N_5872,N_4453,N_4153);
and U5873 (N_5873,N_4573,N_4909);
and U5874 (N_5874,N_4628,N_4151);
nor U5875 (N_5875,N_4572,N_4031);
nor U5876 (N_5876,N_4923,N_4757);
or U5877 (N_5877,N_4013,N_4769);
or U5878 (N_5878,N_4045,N_4452);
nand U5879 (N_5879,N_4698,N_4235);
nor U5880 (N_5880,N_4107,N_4030);
and U5881 (N_5881,N_4647,N_4005);
or U5882 (N_5882,N_4392,N_4950);
nor U5883 (N_5883,N_4994,N_4776);
and U5884 (N_5884,N_4864,N_4371);
nand U5885 (N_5885,N_4395,N_4913);
or U5886 (N_5886,N_4849,N_4455);
nor U5887 (N_5887,N_4893,N_4486);
and U5888 (N_5888,N_4916,N_4326);
or U5889 (N_5889,N_4293,N_4304);
xor U5890 (N_5890,N_4960,N_4312);
or U5891 (N_5891,N_4444,N_4325);
nor U5892 (N_5892,N_4626,N_4143);
and U5893 (N_5893,N_4576,N_4225);
or U5894 (N_5894,N_4861,N_4641);
or U5895 (N_5895,N_4758,N_4863);
nand U5896 (N_5896,N_4080,N_4274);
nand U5897 (N_5897,N_4727,N_4003);
nor U5898 (N_5898,N_4473,N_4514);
nand U5899 (N_5899,N_4099,N_4607);
xor U5900 (N_5900,N_4949,N_4329);
nor U5901 (N_5901,N_4268,N_4603);
or U5902 (N_5902,N_4986,N_4328);
xor U5903 (N_5903,N_4011,N_4983);
and U5904 (N_5904,N_4051,N_4772);
nor U5905 (N_5905,N_4045,N_4984);
nand U5906 (N_5906,N_4435,N_4363);
and U5907 (N_5907,N_4588,N_4028);
nand U5908 (N_5908,N_4932,N_4953);
and U5909 (N_5909,N_4647,N_4121);
nand U5910 (N_5910,N_4915,N_4138);
or U5911 (N_5911,N_4465,N_4538);
nor U5912 (N_5912,N_4999,N_4183);
nor U5913 (N_5913,N_4519,N_4708);
and U5914 (N_5914,N_4267,N_4704);
nand U5915 (N_5915,N_4212,N_4336);
and U5916 (N_5916,N_4260,N_4841);
nand U5917 (N_5917,N_4269,N_4833);
or U5918 (N_5918,N_4748,N_4643);
nand U5919 (N_5919,N_4958,N_4291);
nand U5920 (N_5920,N_4795,N_4748);
or U5921 (N_5921,N_4586,N_4679);
nand U5922 (N_5922,N_4975,N_4966);
or U5923 (N_5923,N_4851,N_4963);
xnor U5924 (N_5924,N_4407,N_4455);
or U5925 (N_5925,N_4583,N_4283);
or U5926 (N_5926,N_4827,N_4307);
or U5927 (N_5927,N_4375,N_4216);
or U5928 (N_5928,N_4407,N_4039);
and U5929 (N_5929,N_4876,N_4430);
nor U5930 (N_5930,N_4035,N_4669);
nand U5931 (N_5931,N_4448,N_4565);
nor U5932 (N_5932,N_4080,N_4639);
or U5933 (N_5933,N_4584,N_4715);
nor U5934 (N_5934,N_4275,N_4854);
and U5935 (N_5935,N_4290,N_4755);
nor U5936 (N_5936,N_4138,N_4809);
or U5937 (N_5937,N_4236,N_4710);
nand U5938 (N_5938,N_4770,N_4986);
nor U5939 (N_5939,N_4067,N_4062);
nor U5940 (N_5940,N_4590,N_4000);
or U5941 (N_5941,N_4095,N_4402);
or U5942 (N_5942,N_4790,N_4003);
nand U5943 (N_5943,N_4692,N_4917);
nor U5944 (N_5944,N_4091,N_4495);
nand U5945 (N_5945,N_4546,N_4636);
nor U5946 (N_5946,N_4910,N_4295);
nand U5947 (N_5947,N_4978,N_4814);
nor U5948 (N_5948,N_4503,N_4407);
and U5949 (N_5949,N_4484,N_4286);
and U5950 (N_5950,N_4459,N_4608);
nor U5951 (N_5951,N_4200,N_4352);
and U5952 (N_5952,N_4756,N_4002);
nand U5953 (N_5953,N_4978,N_4185);
nand U5954 (N_5954,N_4325,N_4778);
nor U5955 (N_5955,N_4433,N_4331);
or U5956 (N_5956,N_4923,N_4661);
and U5957 (N_5957,N_4402,N_4579);
or U5958 (N_5958,N_4428,N_4909);
xnor U5959 (N_5959,N_4081,N_4280);
nand U5960 (N_5960,N_4658,N_4977);
xor U5961 (N_5961,N_4141,N_4660);
and U5962 (N_5962,N_4377,N_4727);
xor U5963 (N_5963,N_4120,N_4394);
nor U5964 (N_5964,N_4478,N_4143);
nand U5965 (N_5965,N_4621,N_4586);
and U5966 (N_5966,N_4250,N_4936);
or U5967 (N_5967,N_4210,N_4280);
and U5968 (N_5968,N_4704,N_4281);
or U5969 (N_5969,N_4892,N_4056);
and U5970 (N_5970,N_4920,N_4976);
nor U5971 (N_5971,N_4468,N_4776);
or U5972 (N_5972,N_4927,N_4137);
or U5973 (N_5973,N_4990,N_4449);
and U5974 (N_5974,N_4239,N_4552);
and U5975 (N_5975,N_4000,N_4559);
and U5976 (N_5976,N_4435,N_4207);
nor U5977 (N_5977,N_4482,N_4667);
nor U5978 (N_5978,N_4766,N_4955);
and U5979 (N_5979,N_4534,N_4343);
nand U5980 (N_5980,N_4094,N_4946);
or U5981 (N_5981,N_4091,N_4919);
or U5982 (N_5982,N_4346,N_4217);
and U5983 (N_5983,N_4437,N_4976);
nand U5984 (N_5984,N_4845,N_4400);
nand U5985 (N_5985,N_4414,N_4295);
nor U5986 (N_5986,N_4200,N_4248);
nor U5987 (N_5987,N_4943,N_4195);
and U5988 (N_5988,N_4362,N_4919);
xnor U5989 (N_5989,N_4060,N_4679);
nand U5990 (N_5990,N_4378,N_4919);
nand U5991 (N_5991,N_4456,N_4713);
or U5992 (N_5992,N_4748,N_4021);
and U5993 (N_5993,N_4805,N_4882);
or U5994 (N_5994,N_4173,N_4700);
and U5995 (N_5995,N_4587,N_4102);
nor U5996 (N_5996,N_4716,N_4602);
or U5997 (N_5997,N_4726,N_4553);
and U5998 (N_5998,N_4750,N_4081);
and U5999 (N_5999,N_4835,N_4493);
nor U6000 (N_6000,N_5191,N_5597);
and U6001 (N_6001,N_5827,N_5327);
and U6002 (N_6002,N_5808,N_5345);
xnor U6003 (N_6003,N_5602,N_5775);
nor U6004 (N_6004,N_5019,N_5411);
and U6005 (N_6005,N_5279,N_5490);
and U6006 (N_6006,N_5122,N_5944);
nor U6007 (N_6007,N_5621,N_5206);
nor U6008 (N_6008,N_5359,N_5519);
nand U6009 (N_6009,N_5590,N_5509);
xor U6010 (N_6010,N_5097,N_5998);
and U6011 (N_6011,N_5702,N_5055);
nand U6012 (N_6012,N_5347,N_5299);
nor U6013 (N_6013,N_5505,N_5231);
or U6014 (N_6014,N_5009,N_5820);
and U6015 (N_6015,N_5027,N_5050);
nand U6016 (N_6016,N_5170,N_5230);
or U6017 (N_6017,N_5005,N_5907);
nand U6018 (N_6018,N_5551,N_5938);
or U6019 (N_6019,N_5570,N_5884);
xnor U6020 (N_6020,N_5440,N_5840);
and U6021 (N_6021,N_5741,N_5445);
nor U6022 (N_6022,N_5696,N_5360);
and U6023 (N_6023,N_5990,N_5160);
nor U6024 (N_6024,N_5192,N_5951);
nand U6025 (N_6025,N_5633,N_5461);
nor U6026 (N_6026,N_5109,N_5976);
xnor U6027 (N_6027,N_5611,N_5213);
and U6028 (N_6028,N_5473,N_5077);
nor U6029 (N_6029,N_5797,N_5744);
nand U6030 (N_6030,N_5575,N_5755);
xor U6031 (N_6031,N_5225,N_5066);
nand U6032 (N_6032,N_5806,N_5259);
xnor U6033 (N_6033,N_5865,N_5999);
nor U6034 (N_6034,N_5526,N_5662);
and U6035 (N_6035,N_5856,N_5801);
and U6036 (N_6036,N_5614,N_5042);
nor U6037 (N_6037,N_5392,N_5628);
or U6038 (N_6038,N_5914,N_5475);
nor U6039 (N_6039,N_5319,N_5516);
and U6040 (N_6040,N_5261,N_5970);
nand U6041 (N_6041,N_5961,N_5307);
nand U6042 (N_6042,N_5480,N_5555);
and U6043 (N_6043,N_5400,N_5496);
nor U6044 (N_6044,N_5791,N_5150);
nor U6045 (N_6045,N_5011,N_5648);
or U6046 (N_6046,N_5228,N_5442);
xor U6047 (N_6047,N_5935,N_5435);
nor U6048 (N_6048,N_5053,N_5243);
or U6049 (N_6049,N_5926,N_5450);
nor U6050 (N_6050,N_5260,N_5760);
or U6051 (N_6051,N_5098,N_5922);
nand U6052 (N_6052,N_5323,N_5014);
nor U6053 (N_6053,N_5390,N_5304);
and U6054 (N_6054,N_5276,N_5043);
or U6055 (N_6055,N_5069,N_5089);
xor U6056 (N_6056,N_5668,N_5952);
nand U6057 (N_6057,N_5864,N_5193);
nand U6058 (N_6058,N_5444,N_5457);
and U6059 (N_6059,N_5452,N_5068);
and U6060 (N_6060,N_5067,N_5318);
or U6061 (N_6061,N_5655,N_5414);
nor U6062 (N_6062,N_5754,N_5245);
nand U6063 (N_6063,N_5129,N_5572);
nor U6064 (N_6064,N_5402,N_5745);
and U6065 (N_6065,N_5740,N_5131);
or U6066 (N_6066,N_5282,N_5542);
nor U6067 (N_6067,N_5506,N_5479);
and U6068 (N_6068,N_5703,N_5823);
xnor U6069 (N_6069,N_5645,N_5128);
nor U6070 (N_6070,N_5832,N_5691);
xnor U6071 (N_6071,N_5088,N_5091);
or U6072 (N_6072,N_5108,N_5830);
and U6073 (N_6073,N_5185,N_5759);
and U6074 (N_6074,N_5737,N_5373);
nor U6075 (N_6075,N_5449,N_5369);
and U6076 (N_6076,N_5729,N_5671);
and U6077 (N_6077,N_5867,N_5816);
nand U6078 (N_6078,N_5476,N_5749);
and U6079 (N_6079,N_5713,N_5381);
and U6080 (N_6080,N_5266,N_5303);
or U6081 (N_6081,N_5061,N_5636);
and U6082 (N_6082,N_5664,N_5644);
nor U6083 (N_6083,N_5370,N_5924);
xnor U6084 (N_6084,N_5119,N_5874);
xnor U6085 (N_6085,N_5649,N_5796);
or U6086 (N_6086,N_5446,N_5837);
nor U6087 (N_6087,N_5071,N_5658);
nand U6088 (N_6088,N_5888,N_5036);
and U6089 (N_6089,N_5020,N_5571);
and U6090 (N_6090,N_5886,N_5894);
xnor U6091 (N_6091,N_5448,N_5333);
or U6092 (N_6092,N_5424,N_5599);
and U6093 (N_6093,N_5543,N_5157);
and U6094 (N_6094,N_5013,N_5992);
and U6095 (N_6095,N_5210,N_5609);
or U6096 (N_6096,N_5140,N_5877);
xnor U6097 (N_6097,N_5568,N_5289);
nor U6098 (N_6098,N_5681,N_5685);
xnor U6099 (N_6099,N_5637,N_5725);
and U6100 (N_6100,N_5305,N_5386);
and U6101 (N_6101,N_5472,N_5374);
nand U6102 (N_6102,N_5205,N_5394);
nand U6103 (N_6103,N_5474,N_5525);
or U6104 (N_6104,N_5625,N_5781);
nor U6105 (N_6105,N_5463,N_5983);
nand U6106 (N_6106,N_5711,N_5296);
or U6107 (N_6107,N_5149,N_5143);
or U6108 (N_6108,N_5401,N_5382);
or U6109 (N_6109,N_5872,N_5072);
nor U6110 (N_6110,N_5736,N_5675);
nor U6111 (N_6111,N_5340,N_5209);
nand U6112 (N_6112,N_5683,N_5618);
nor U6113 (N_6113,N_5776,N_5470);
or U6114 (N_6114,N_5785,N_5803);
xnor U6115 (N_6115,N_5810,N_5412);
and U6116 (N_6116,N_5849,N_5587);
or U6117 (N_6117,N_5780,N_5226);
nand U6118 (N_6118,N_5393,N_5102);
xor U6119 (N_6119,N_5987,N_5380);
nor U6120 (N_6120,N_5627,N_5742);
or U6121 (N_6121,N_5826,N_5378);
nor U6122 (N_6122,N_5031,N_5447);
and U6123 (N_6123,N_5632,N_5739);
nand U6124 (N_6124,N_5464,N_5025);
nand U6125 (N_6125,N_5168,N_5674);
and U6126 (N_6126,N_5018,N_5265);
nand U6127 (N_6127,N_5631,N_5764);
or U6128 (N_6128,N_5667,N_5134);
and U6129 (N_6129,N_5972,N_5673);
nor U6130 (N_6130,N_5073,N_5881);
xor U6131 (N_6131,N_5166,N_5788);
and U6132 (N_6132,N_5811,N_5385);
and U6133 (N_6133,N_5024,N_5548);
nand U6134 (N_6134,N_5250,N_5107);
nor U6135 (N_6135,N_5301,N_5145);
nor U6136 (N_6136,N_5701,N_5604);
or U6137 (N_6137,N_5178,N_5495);
nor U6138 (N_6138,N_5917,N_5985);
nor U6139 (N_6139,N_5561,N_5203);
xor U6140 (N_6140,N_5275,N_5295);
and U6141 (N_6141,N_5586,N_5286);
nor U6142 (N_6142,N_5873,N_5793);
and U6143 (N_6143,N_5986,N_5251);
nand U6144 (N_6144,N_5123,N_5535);
or U6145 (N_6145,N_5326,N_5167);
and U6146 (N_6146,N_5104,N_5747);
and U6147 (N_6147,N_5771,N_5684);
nor U6148 (N_6148,N_5515,N_5248);
nor U6149 (N_6149,N_5094,N_5404);
xnor U6150 (N_6150,N_5346,N_5866);
or U6151 (N_6151,N_5316,N_5730);
xnor U6152 (N_6152,N_5416,N_5659);
and U6153 (N_6153,N_5851,N_5343);
nand U6154 (N_6154,N_5715,N_5105);
and U6155 (N_6155,N_5117,N_5812);
or U6156 (N_6156,N_5443,N_5748);
or U6157 (N_6157,N_5669,N_5732);
and U6158 (N_6158,N_5844,N_5666);
nor U6159 (N_6159,N_5605,N_5078);
nand U6160 (N_6160,N_5321,N_5798);
nand U6161 (N_6161,N_5906,N_5606);
nand U6162 (N_6162,N_5966,N_5317);
nor U6163 (N_6163,N_5719,N_5254);
nor U6164 (N_6164,N_5152,N_5521);
and U6165 (N_6165,N_5512,N_5728);
or U6166 (N_6166,N_5482,N_5724);
nand U6167 (N_6167,N_5142,N_5647);
and U6168 (N_6168,N_5903,N_5115);
nor U6169 (N_6169,N_5177,N_5549);
and U6170 (N_6170,N_5395,N_5196);
nor U6171 (N_6171,N_5531,N_5032);
nor U6172 (N_6172,N_5908,N_5534);
xor U6173 (N_6173,N_5518,N_5331);
nand U6174 (N_6174,N_5528,N_5086);
and U6175 (N_6175,N_5676,N_5290);
nand U6176 (N_6176,N_5915,N_5132);
nor U6177 (N_6177,N_5436,N_5188);
nor U6178 (N_6178,N_5171,N_5617);
and U6179 (N_6179,N_5106,N_5640);
nand U6180 (N_6180,N_5692,N_5391);
nand U6181 (N_6181,N_5893,N_5697);
nor U6182 (N_6182,N_5984,N_5147);
or U6183 (N_6183,N_5136,N_5639);
nand U6184 (N_6184,N_5629,N_5580);
or U6185 (N_6185,N_5945,N_5410);
nor U6186 (N_6186,N_5767,N_5956);
and U6187 (N_6187,N_5522,N_5680);
or U6188 (N_6188,N_5234,N_5437);
nand U6189 (N_6189,N_5302,N_5332);
nor U6190 (N_6190,N_5799,N_5238);
or U6191 (N_6191,N_5033,N_5179);
nor U6192 (N_6192,N_5194,N_5137);
xnor U6193 (N_6193,N_5557,N_5779);
or U6194 (N_6194,N_5271,N_5267);
nor U6195 (N_6195,N_5379,N_5708);
nand U6196 (N_6196,N_5727,N_5465);
nand U6197 (N_6197,N_5963,N_5315);
or U6198 (N_6198,N_5015,N_5855);
nand U6199 (N_6199,N_5578,N_5284);
nor U6200 (N_6200,N_5172,N_5233);
or U6201 (N_6201,N_5765,N_5070);
nor U6202 (N_6202,N_5207,N_5221);
nor U6203 (N_6203,N_5413,N_5912);
or U6204 (N_6204,N_5573,N_5127);
and U6205 (N_6205,N_5931,N_5320);
xor U6206 (N_6206,N_5901,N_5734);
or U6207 (N_6207,N_5274,N_5537);
xnor U6208 (N_6208,N_5423,N_5634);
nand U6209 (N_6209,N_5037,N_5861);
nand U6210 (N_6210,N_5709,N_5698);
nor U6211 (N_6211,N_5012,N_5195);
and U6212 (N_6212,N_5035,N_5962);
or U6213 (N_6213,N_5199,N_5198);
nor U6214 (N_6214,N_5746,N_5902);
xor U6215 (N_6215,N_5743,N_5536);
nor U6216 (N_6216,N_5052,N_5154);
nand U6217 (N_6217,N_5868,N_5407);
or U6218 (N_6218,N_5778,N_5281);
or U6219 (N_6219,N_5112,N_5163);
or U6220 (N_6220,N_5610,N_5705);
or U6221 (N_6221,N_5859,N_5885);
xnor U6222 (N_6222,N_5264,N_5219);
nor U6223 (N_6223,N_5354,N_5040);
nor U6224 (N_6224,N_5829,N_5690);
or U6225 (N_6225,N_5663,N_5362);
or U6226 (N_6226,N_5039,N_5982);
nor U6227 (N_6227,N_5135,N_5406);
and U6228 (N_6228,N_5022,N_5189);
and U6229 (N_6229,N_5929,N_5314);
nand U6230 (N_6230,N_5898,N_5441);
and U6231 (N_6231,N_5216,N_5419);
nand U6232 (N_6232,N_5624,N_5139);
nor U6233 (N_6233,N_5918,N_5707);
nor U6234 (N_6234,N_5151,N_5766);
nor U6235 (N_6235,N_5467,N_5583);
or U6236 (N_6236,N_5656,N_5242);
nor U6237 (N_6237,N_5925,N_5358);
or U6238 (N_6238,N_5110,N_5298);
or U6239 (N_6239,N_5366,N_5064);
nand U6240 (N_6240,N_5654,N_5116);
nand U6241 (N_6241,N_5991,N_5890);
or U6242 (N_6242,N_5118,N_5857);
and U6243 (N_6243,N_5240,N_5161);
and U6244 (N_6244,N_5026,N_5792);
nand U6245 (N_6245,N_5396,N_5850);
nand U6246 (N_6246,N_5481,N_5761);
nand U6247 (N_6247,N_5054,N_5252);
and U6248 (N_6248,N_5940,N_5076);
and U6249 (N_6249,N_5021,N_5427);
nor U6250 (N_6250,N_5485,N_5834);
and U6251 (N_6251,N_5498,N_5492);
xor U6252 (N_6252,N_5538,N_5312);
nand U6253 (N_6253,N_5501,N_5795);
xor U6254 (N_6254,N_5576,N_5372);
nand U6255 (N_6255,N_5155,N_5126);
nand U6256 (N_6256,N_5477,N_5616);
xor U6257 (N_6257,N_5074,N_5847);
nand U6258 (N_6258,N_5202,N_5060);
nand U6259 (N_6259,N_5959,N_5733);
nor U6260 (N_6260,N_5777,N_5095);
nor U6261 (N_6261,N_5559,N_5581);
and U6262 (N_6262,N_5615,N_5458);
or U6263 (N_6263,N_5397,N_5699);
nor U6264 (N_6264,N_5428,N_5751);
nor U6265 (N_6265,N_5330,N_5566);
or U6266 (N_6266,N_5084,N_5367);
and U6267 (N_6267,N_5297,N_5533);
nand U6268 (N_6268,N_5059,N_5694);
xnor U6269 (N_6269,N_5138,N_5817);
nand U6270 (N_6270,N_5062,N_5080);
and U6271 (N_6271,N_5222,N_5438);
nand U6272 (N_6272,N_5459,N_5075);
or U6273 (N_6273,N_5383,N_5831);
and U6274 (N_6274,N_5603,N_5933);
nor U6275 (N_6275,N_5942,N_5686);
and U6276 (N_6276,N_5208,N_5735);
nand U6277 (N_6277,N_5622,N_5090);
xnor U6278 (N_6278,N_5399,N_5562);
or U6279 (N_6279,N_5153,N_5204);
or U6280 (N_6280,N_5249,N_5565);
nor U6281 (N_6281,N_5247,N_5943);
nand U6282 (N_6282,N_5341,N_5910);
or U6283 (N_6283,N_5688,N_5141);
or U6284 (N_6284,N_5384,N_5967);
nor U6285 (N_6285,N_5169,N_5891);
xor U6286 (N_6286,N_5180,N_5456);
nand U6287 (N_6287,N_5598,N_5594);
and U6288 (N_6288,N_5293,N_5514);
or U6289 (N_6289,N_5946,N_5388);
nand U6290 (N_6290,N_5041,N_5371);
and U6291 (N_6291,N_5882,N_5641);
nand U6292 (N_6292,N_5841,N_5045);
or U6293 (N_6293,N_5977,N_5723);
and U6294 (N_6294,N_5722,N_5964);
and U6295 (N_6295,N_5113,N_5954);
xnor U6296 (N_6296,N_5772,N_5220);
or U6297 (N_6297,N_5883,N_5704);
xor U6298 (N_6298,N_5453,N_5608);
nor U6299 (N_6299,N_5545,N_5941);
and U6300 (N_6300,N_5934,N_5563);
and U6301 (N_6301,N_5805,N_5232);
xor U6302 (N_6302,N_5635,N_5913);
nor U6303 (N_6303,N_5235,N_5835);
xor U6304 (N_6304,N_5786,N_5768);
or U6305 (N_6305,N_5842,N_5409);
or U6306 (N_6306,N_5821,N_5824);
or U6307 (N_6307,N_5661,N_5677);
nor U6308 (N_6308,N_5353,N_5313);
or U6309 (N_6309,N_5229,N_5044);
and U6310 (N_6310,N_5889,N_5130);
nor U6311 (N_6311,N_5556,N_5365);
nor U6312 (N_6312,N_5920,N_5224);
and U6313 (N_6313,N_5978,N_5006);
and U6314 (N_6314,N_5418,N_5101);
nand U6315 (N_6315,N_5981,N_5717);
nand U6316 (N_6316,N_5560,N_5308);
or U6317 (N_6317,N_5726,N_5589);
or U6318 (N_6318,N_5965,N_5968);
and U6319 (N_6319,N_5651,N_5355);
nor U6320 (N_6320,N_5876,N_5994);
nand U6321 (N_6321,N_5591,N_5895);
and U6322 (N_6322,N_5995,N_5752);
and U6323 (N_6323,N_5007,N_5268);
xnor U6324 (N_6324,N_5309,N_5756);
nor U6325 (N_6325,N_5186,N_5344);
or U6326 (N_6326,N_5291,N_5524);
and U6327 (N_6327,N_5283,N_5679);
nand U6328 (N_6328,N_5214,N_5051);
and U6329 (N_6329,N_5949,N_5361);
nand U6330 (N_6330,N_5911,N_5958);
nand U6331 (N_6331,N_5306,N_5652);
nand U6332 (N_6332,N_5494,N_5434);
and U6333 (N_6333,N_5211,N_5769);
and U6334 (N_6334,N_5339,N_5085);
and U6335 (N_6335,N_5974,N_5921);
or U6336 (N_6336,N_5695,N_5612);
nor U6337 (N_6337,N_5335,N_5953);
and U6338 (N_6338,N_5577,N_5415);
nand U6339 (N_6339,N_5493,N_5357);
nor U6340 (N_6340,N_5263,N_5693);
nor U6341 (N_6341,N_5550,N_5356);
nor U6342 (N_6342,N_5646,N_5596);
nand U6343 (N_6343,N_5422,N_5451);
or U6344 (N_6344,N_5016,N_5672);
nand U6345 (N_6345,N_5718,N_5258);
or U6346 (N_6346,N_5499,N_5466);
or U6347 (N_6347,N_5217,N_5818);
nor U6348 (N_6348,N_5774,N_5939);
nor U6349 (N_6349,N_5486,N_5038);
nor U6350 (N_6350,N_5081,N_5593);
or U6351 (N_6351,N_5469,N_5497);
or U6352 (N_6352,N_5517,N_5523);
or U6353 (N_6353,N_5600,N_5969);
nor U6354 (N_6354,N_5763,N_5540);
nor U6355 (N_6355,N_5630,N_5431);
nor U6356 (N_6356,N_5716,N_5770);
or U6357 (N_6357,N_5454,N_5046);
nor U6358 (N_6358,N_5858,N_5004);
nor U6359 (N_6359,N_5433,N_5455);
nor U6360 (N_6360,N_5789,N_5334);
nor U6361 (N_6361,N_5919,N_5133);
and U6362 (N_6362,N_5638,N_5753);
and U6363 (N_6363,N_5687,N_5430);
nand U6364 (N_6364,N_5270,N_5272);
or U6365 (N_6365,N_5028,N_5176);
nor U6366 (N_6366,N_5417,N_5278);
nand U6367 (N_6367,N_5529,N_5121);
and U6368 (N_6368,N_5750,N_5184);
or U6369 (N_6369,N_5955,N_5239);
nor U6370 (N_6370,N_5870,N_5905);
nand U6371 (N_6371,N_5975,N_5862);
xor U6372 (N_6372,N_5324,N_5584);
nor U6373 (N_6373,N_5642,N_5544);
nor U6374 (N_6374,N_5285,N_5403);
or U6375 (N_6375,N_5710,N_5996);
xor U6376 (N_6376,N_5083,N_5338);
nor U6377 (N_6377,N_5350,N_5030);
and U6378 (N_6378,N_5852,N_5223);
nand U6379 (N_6379,N_5825,N_5325);
nand U6380 (N_6380,N_5574,N_5262);
nor U6381 (N_6381,N_5253,N_5504);
nor U6382 (N_6382,N_5714,N_5530);
nand U6383 (N_6383,N_5626,N_5336);
and U6384 (N_6384,N_5124,N_5079);
nor U6385 (N_6385,N_5552,N_5439);
or U6386 (N_6386,N_5706,N_5848);
nor U6387 (N_6387,N_5310,N_5813);
or U6388 (N_6388,N_5569,N_5896);
nand U6389 (N_6389,N_5989,N_5057);
and U6390 (N_6390,N_5553,N_5056);
nand U6391 (N_6391,N_5904,N_5173);
nor U6392 (N_6392,N_5807,N_5513);
or U6393 (N_6393,N_5853,N_5421);
and U6394 (N_6394,N_5782,N_5937);
nor U6395 (N_6395,N_5880,N_5099);
nor U6396 (N_6396,N_5377,N_5280);
nor U6397 (N_6397,N_5507,N_5114);
nor U6398 (N_6398,N_5029,N_5420);
and U6399 (N_6399,N_5197,N_5183);
and U6400 (N_6400,N_5567,N_5815);
and U6401 (N_6401,N_5854,N_5227);
nor U6402 (N_6402,N_5607,N_5120);
nor U6403 (N_6403,N_5348,N_5273);
or U6404 (N_6404,N_5731,N_5546);
or U6405 (N_6405,N_5255,N_5814);
or U6406 (N_6406,N_5843,N_5794);
nor U6407 (N_6407,N_5368,N_5187);
nand U6408 (N_6408,N_5897,N_5181);
or U6409 (N_6409,N_5802,N_5063);
or U6410 (N_6410,N_5471,N_5292);
nor U6411 (N_6411,N_5712,N_5783);
nor U6412 (N_6412,N_5900,N_5980);
nand U6413 (N_6413,N_5948,N_5787);
and U6414 (N_6414,N_5241,N_5375);
or U6415 (N_6415,N_5650,N_5478);
and U6416 (N_6416,N_5916,N_5426);
or U6417 (N_6417,N_5065,N_5988);
and U6418 (N_6418,N_5364,N_5809);
or U6419 (N_6419,N_5483,N_5269);
nand U6420 (N_6420,N_5215,N_5909);
or U6421 (N_6421,N_5846,N_5398);
nor U6422 (N_6422,N_5329,N_5757);
xnor U6423 (N_6423,N_5023,N_5111);
or U6424 (N_6424,N_5585,N_5558);
nand U6425 (N_6425,N_5887,N_5619);
xnor U6426 (N_6426,N_5034,N_5087);
and U6427 (N_6427,N_5363,N_5960);
nor U6428 (N_6428,N_5484,N_5878);
nor U6429 (N_6429,N_5564,N_5508);
nand U6430 (N_6430,N_5790,N_5491);
nand U6431 (N_6431,N_5287,N_5236);
nand U6432 (N_6432,N_5822,N_5588);
and U6433 (N_6433,N_5947,N_5256);
and U6434 (N_6434,N_5670,N_5758);
and U6435 (N_6435,N_5146,N_5277);
nand U6436 (N_6436,N_5294,N_5001);
nand U6437 (N_6437,N_5096,N_5839);
nor U6438 (N_6438,N_5049,N_5376);
or U6439 (N_6439,N_5156,N_5082);
or U6440 (N_6440,N_5971,N_5721);
or U6441 (N_6441,N_5860,N_5541);
nand U6442 (N_6442,N_5973,N_5579);
or U6443 (N_6443,N_5288,N_5502);
nor U6444 (N_6444,N_5869,N_5349);
or U6445 (N_6445,N_5174,N_5657);
xor U6446 (N_6446,N_5158,N_5979);
nor U6447 (N_6447,N_5387,N_5923);
and U6448 (N_6448,N_5017,N_5500);
and U6449 (N_6449,N_5773,N_5468);
or U6450 (N_6450,N_5527,N_5510);
and U6451 (N_6451,N_5212,N_5162);
xnor U6452 (N_6452,N_5892,N_5148);
nand U6453 (N_6453,N_5164,N_5863);
or U6454 (N_6454,N_5845,N_5165);
nand U6455 (N_6455,N_5620,N_5144);
or U6456 (N_6456,N_5432,N_5930);
and U6457 (N_6457,N_5322,N_5048);
nor U6458 (N_6458,N_5246,N_5489);
nand U6459 (N_6459,N_5700,N_5613);
nand U6460 (N_6460,N_5429,N_5093);
nor U6461 (N_6461,N_5405,N_5337);
and U6462 (N_6462,N_5218,N_5003);
and U6463 (N_6463,N_5460,N_5351);
and U6464 (N_6464,N_5993,N_5547);
or U6465 (N_6465,N_5047,N_5008);
or U6466 (N_6466,N_5237,N_5592);
nor U6467 (N_6467,N_5800,N_5899);
nand U6468 (N_6468,N_5503,N_5879);
xor U6469 (N_6469,N_5190,N_5936);
nor U6470 (N_6470,N_5100,N_5408);
nand U6471 (N_6471,N_5957,N_5875);
nor U6472 (N_6472,N_5762,N_5665);
and U6473 (N_6473,N_5300,N_5927);
nand U6474 (N_6474,N_5389,N_5257);
xor U6475 (N_6475,N_5643,N_5804);
and U6476 (N_6476,N_5833,N_5175);
nand U6477 (N_6477,N_5488,N_5819);
and U6478 (N_6478,N_5660,N_5720);
and U6479 (N_6479,N_5539,N_5010);
and U6480 (N_6480,N_5352,N_5311);
nand U6481 (N_6481,N_5784,N_5623);
xnor U6482 (N_6482,N_5328,N_5682);
or U6483 (N_6483,N_5092,N_5342);
nand U6484 (N_6484,N_5511,N_5595);
nor U6485 (N_6485,N_5653,N_5058);
or U6486 (N_6486,N_5838,N_5244);
nand U6487 (N_6487,N_5462,N_5103);
nor U6488 (N_6488,N_5678,N_5928);
nor U6489 (N_6489,N_5182,N_5871);
nand U6490 (N_6490,N_5487,N_5828);
nor U6491 (N_6491,N_5000,N_5200);
nand U6492 (N_6492,N_5554,N_5532);
xor U6493 (N_6493,N_5689,N_5125);
nor U6494 (N_6494,N_5201,N_5836);
xnor U6495 (N_6495,N_5950,N_5601);
nand U6496 (N_6496,N_5582,N_5738);
nor U6497 (N_6497,N_5997,N_5159);
or U6498 (N_6498,N_5520,N_5932);
or U6499 (N_6499,N_5425,N_5002);
or U6500 (N_6500,N_5331,N_5738);
and U6501 (N_6501,N_5120,N_5652);
nor U6502 (N_6502,N_5499,N_5378);
or U6503 (N_6503,N_5362,N_5574);
or U6504 (N_6504,N_5142,N_5298);
or U6505 (N_6505,N_5181,N_5463);
or U6506 (N_6506,N_5580,N_5816);
nand U6507 (N_6507,N_5860,N_5126);
and U6508 (N_6508,N_5851,N_5512);
xnor U6509 (N_6509,N_5579,N_5626);
xnor U6510 (N_6510,N_5457,N_5523);
nand U6511 (N_6511,N_5015,N_5204);
or U6512 (N_6512,N_5509,N_5533);
and U6513 (N_6513,N_5678,N_5632);
or U6514 (N_6514,N_5178,N_5688);
and U6515 (N_6515,N_5501,N_5506);
and U6516 (N_6516,N_5830,N_5542);
nor U6517 (N_6517,N_5337,N_5963);
nor U6518 (N_6518,N_5650,N_5608);
or U6519 (N_6519,N_5307,N_5299);
or U6520 (N_6520,N_5017,N_5029);
or U6521 (N_6521,N_5191,N_5989);
xor U6522 (N_6522,N_5500,N_5206);
or U6523 (N_6523,N_5038,N_5307);
or U6524 (N_6524,N_5537,N_5533);
nand U6525 (N_6525,N_5131,N_5759);
nor U6526 (N_6526,N_5995,N_5704);
xnor U6527 (N_6527,N_5157,N_5099);
and U6528 (N_6528,N_5678,N_5962);
and U6529 (N_6529,N_5048,N_5927);
nand U6530 (N_6530,N_5708,N_5227);
and U6531 (N_6531,N_5667,N_5774);
xor U6532 (N_6532,N_5354,N_5731);
and U6533 (N_6533,N_5483,N_5362);
nand U6534 (N_6534,N_5606,N_5890);
nand U6535 (N_6535,N_5997,N_5923);
xnor U6536 (N_6536,N_5726,N_5321);
nor U6537 (N_6537,N_5031,N_5988);
or U6538 (N_6538,N_5230,N_5831);
nand U6539 (N_6539,N_5263,N_5638);
nor U6540 (N_6540,N_5242,N_5253);
nor U6541 (N_6541,N_5688,N_5152);
and U6542 (N_6542,N_5903,N_5637);
and U6543 (N_6543,N_5661,N_5114);
and U6544 (N_6544,N_5420,N_5783);
or U6545 (N_6545,N_5266,N_5430);
or U6546 (N_6546,N_5886,N_5373);
or U6547 (N_6547,N_5839,N_5499);
xor U6548 (N_6548,N_5827,N_5048);
nand U6549 (N_6549,N_5449,N_5642);
nor U6550 (N_6550,N_5030,N_5931);
nand U6551 (N_6551,N_5527,N_5931);
xnor U6552 (N_6552,N_5273,N_5388);
or U6553 (N_6553,N_5944,N_5069);
and U6554 (N_6554,N_5278,N_5090);
nand U6555 (N_6555,N_5984,N_5031);
xor U6556 (N_6556,N_5244,N_5551);
nand U6557 (N_6557,N_5581,N_5927);
and U6558 (N_6558,N_5372,N_5278);
and U6559 (N_6559,N_5011,N_5569);
and U6560 (N_6560,N_5516,N_5155);
nand U6561 (N_6561,N_5631,N_5300);
or U6562 (N_6562,N_5614,N_5334);
nor U6563 (N_6563,N_5971,N_5869);
nand U6564 (N_6564,N_5307,N_5929);
or U6565 (N_6565,N_5598,N_5491);
nand U6566 (N_6566,N_5945,N_5540);
or U6567 (N_6567,N_5320,N_5183);
nor U6568 (N_6568,N_5791,N_5533);
and U6569 (N_6569,N_5544,N_5030);
nand U6570 (N_6570,N_5219,N_5296);
or U6571 (N_6571,N_5331,N_5200);
or U6572 (N_6572,N_5623,N_5767);
nor U6573 (N_6573,N_5577,N_5268);
or U6574 (N_6574,N_5947,N_5074);
nand U6575 (N_6575,N_5329,N_5043);
or U6576 (N_6576,N_5437,N_5293);
nand U6577 (N_6577,N_5093,N_5554);
nand U6578 (N_6578,N_5434,N_5115);
or U6579 (N_6579,N_5186,N_5383);
or U6580 (N_6580,N_5638,N_5500);
and U6581 (N_6581,N_5691,N_5405);
nor U6582 (N_6582,N_5038,N_5698);
or U6583 (N_6583,N_5077,N_5031);
nand U6584 (N_6584,N_5668,N_5600);
and U6585 (N_6585,N_5628,N_5006);
xnor U6586 (N_6586,N_5477,N_5288);
and U6587 (N_6587,N_5233,N_5440);
nor U6588 (N_6588,N_5884,N_5041);
or U6589 (N_6589,N_5990,N_5882);
nand U6590 (N_6590,N_5114,N_5014);
xor U6591 (N_6591,N_5697,N_5988);
nand U6592 (N_6592,N_5882,N_5493);
and U6593 (N_6593,N_5571,N_5900);
nor U6594 (N_6594,N_5857,N_5722);
or U6595 (N_6595,N_5237,N_5735);
nor U6596 (N_6596,N_5536,N_5989);
nor U6597 (N_6597,N_5492,N_5897);
nor U6598 (N_6598,N_5734,N_5168);
and U6599 (N_6599,N_5867,N_5356);
and U6600 (N_6600,N_5716,N_5644);
and U6601 (N_6601,N_5478,N_5391);
and U6602 (N_6602,N_5824,N_5949);
nand U6603 (N_6603,N_5954,N_5121);
nor U6604 (N_6604,N_5453,N_5389);
and U6605 (N_6605,N_5970,N_5870);
and U6606 (N_6606,N_5966,N_5115);
and U6607 (N_6607,N_5835,N_5039);
nand U6608 (N_6608,N_5604,N_5833);
nor U6609 (N_6609,N_5238,N_5384);
xor U6610 (N_6610,N_5590,N_5738);
nor U6611 (N_6611,N_5329,N_5091);
nand U6612 (N_6612,N_5672,N_5544);
or U6613 (N_6613,N_5794,N_5482);
or U6614 (N_6614,N_5437,N_5148);
nand U6615 (N_6615,N_5982,N_5880);
xor U6616 (N_6616,N_5237,N_5692);
xor U6617 (N_6617,N_5099,N_5109);
nand U6618 (N_6618,N_5662,N_5215);
or U6619 (N_6619,N_5056,N_5778);
nor U6620 (N_6620,N_5454,N_5700);
nor U6621 (N_6621,N_5464,N_5777);
nand U6622 (N_6622,N_5862,N_5055);
or U6623 (N_6623,N_5794,N_5151);
xor U6624 (N_6624,N_5211,N_5954);
and U6625 (N_6625,N_5343,N_5324);
or U6626 (N_6626,N_5860,N_5049);
or U6627 (N_6627,N_5648,N_5054);
nand U6628 (N_6628,N_5908,N_5207);
nor U6629 (N_6629,N_5475,N_5625);
or U6630 (N_6630,N_5175,N_5158);
and U6631 (N_6631,N_5314,N_5182);
nor U6632 (N_6632,N_5078,N_5106);
and U6633 (N_6633,N_5996,N_5872);
or U6634 (N_6634,N_5180,N_5340);
or U6635 (N_6635,N_5670,N_5904);
and U6636 (N_6636,N_5330,N_5311);
and U6637 (N_6637,N_5518,N_5818);
nor U6638 (N_6638,N_5392,N_5422);
nand U6639 (N_6639,N_5843,N_5202);
and U6640 (N_6640,N_5402,N_5567);
or U6641 (N_6641,N_5714,N_5384);
nor U6642 (N_6642,N_5041,N_5612);
or U6643 (N_6643,N_5277,N_5157);
xnor U6644 (N_6644,N_5706,N_5346);
nand U6645 (N_6645,N_5957,N_5577);
nor U6646 (N_6646,N_5631,N_5608);
or U6647 (N_6647,N_5198,N_5343);
or U6648 (N_6648,N_5068,N_5483);
and U6649 (N_6649,N_5508,N_5266);
nand U6650 (N_6650,N_5155,N_5645);
nand U6651 (N_6651,N_5488,N_5638);
or U6652 (N_6652,N_5140,N_5234);
and U6653 (N_6653,N_5732,N_5389);
or U6654 (N_6654,N_5943,N_5828);
xnor U6655 (N_6655,N_5984,N_5512);
nand U6656 (N_6656,N_5585,N_5803);
and U6657 (N_6657,N_5152,N_5087);
nand U6658 (N_6658,N_5054,N_5463);
nand U6659 (N_6659,N_5629,N_5060);
xor U6660 (N_6660,N_5327,N_5594);
nand U6661 (N_6661,N_5251,N_5004);
nand U6662 (N_6662,N_5300,N_5221);
nor U6663 (N_6663,N_5436,N_5340);
nor U6664 (N_6664,N_5447,N_5432);
and U6665 (N_6665,N_5204,N_5268);
nand U6666 (N_6666,N_5013,N_5541);
nand U6667 (N_6667,N_5531,N_5935);
nand U6668 (N_6668,N_5547,N_5989);
nand U6669 (N_6669,N_5120,N_5263);
xnor U6670 (N_6670,N_5775,N_5712);
and U6671 (N_6671,N_5894,N_5209);
xnor U6672 (N_6672,N_5052,N_5573);
xor U6673 (N_6673,N_5546,N_5278);
or U6674 (N_6674,N_5264,N_5591);
nor U6675 (N_6675,N_5055,N_5363);
and U6676 (N_6676,N_5834,N_5739);
nand U6677 (N_6677,N_5056,N_5829);
and U6678 (N_6678,N_5082,N_5328);
or U6679 (N_6679,N_5707,N_5429);
or U6680 (N_6680,N_5545,N_5765);
nand U6681 (N_6681,N_5335,N_5311);
xnor U6682 (N_6682,N_5223,N_5051);
or U6683 (N_6683,N_5149,N_5789);
nand U6684 (N_6684,N_5715,N_5525);
or U6685 (N_6685,N_5442,N_5768);
xnor U6686 (N_6686,N_5693,N_5217);
nor U6687 (N_6687,N_5067,N_5922);
or U6688 (N_6688,N_5286,N_5563);
nor U6689 (N_6689,N_5333,N_5221);
or U6690 (N_6690,N_5647,N_5015);
and U6691 (N_6691,N_5489,N_5838);
or U6692 (N_6692,N_5541,N_5054);
and U6693 (N_6693,N_5819,N_5920);
xor U6694 (N_6694,N_5711,N_5885);
nand U6695 (N_6695,N_5546,N_5552);
nor U6696 (N_6696,N_5992,N_5899);
nand U6697 (N_6697,N_5733,N_5615);
nand U6698 (N_6698,N_5181,N_5657);
and U6699 (N_6699,N_5424,N_5161);
nor U6700 (N_6700,N_5798,N_5989);
and U6701 (N_6701,N_5725,N_5636);
and U6702 (N_6702,N_5461,N_5717);
nand U6703 (N_6703,N_5464,N_5999);
nand U6704 (N_6704,N_5985,N_5309);
nor U6705 (N_6705,N_5427,N_5759);
nand U6706 (N_6706,N_5407,N_5461);
or U6707 (N_6707,N_5733,N_5222);
nor U6708 (N_6708,N_5860,N_5630);
and U6709 (N_6709,N_5727,N_5190);
nor U6710 (N_6710,N_5924,N_5700);
nand U6711 (N_6711,N_5845,N_5946);
nand U6712 (N_6712,N_5845,N_5369);
or U6713 (N_6713,N_5517,N_5778);
nand U6714 (N_6714,N_5400,N_5719);
nand U6715 (N_6715,N_5834,N_5249);
or U6716 (N_6716,N_5383,N_5410);
and U6717 (N_6717,N_5185,N_5534);
or U6718 (N_6718,N_5566,N_5971);
nand U6719 (N_6719,N_5047,N_5983);
and U6720 (N_6720,N_5734,N_5860);
or U6721 (N_6721,N_5647,N_5451);
or U6722 (N_6722,N_5557,N_5095);
or U6723 (N_6723,N_5121,N_5370);
xor U6724 (N_6724,N_5414,N_5244);
and U6725 (N_6725,N_5493,N_5844);
and U6726 (N_6726,N_5952,N_5479);
and U6727 (N_6727,N_5550,N_5843);
xnor U6728 (N_6728,N_5302,N_5173);
nand U6729 (N_6729,N_5403,N_5423);
or U6730 (N_6730,N_5769,N_5827);
nand U6731 (N_6731,N_5569,N_5683);
xor U6732 (N_6732,N_5349,N_5957);
nand U6733 (N_6733,N_5630,N_5837);
or U6734 (N_6734,N_5144,N_5877);
nor U6735 (N_6735,N_5913,N_5325);
nand U6736 (N_6736,N_5759,N_5304);
or U6737 (N_6737,N_5236,N_5333);
and U6738 (N_6738,N_5214,N_5043);
nor U6739 (N_6739,N_5504,N_5590);
nand U6740 (N_6740,N_5946,N_5172);
and U6741 (N_6741,N_5704,N_5121);
or U6742 (N_6742,N_5515,N_5664);
nor U6743 (N_6743,N_5237,N_5230);
xnor U6744 (N_6744,N_5918,N_5856);
nor U6745 (N_6745,N_5150,N_5056);
and U6746 (N_6746,N_5559,N_5557);
or U6747 (N_6747,N_5381,N_5987);
nand U6748 (N_6748,N_5094,N_5231);
and U6749 (N_6749,N_5390,N_5984);
and U6750 (N_6750,N_5695,N_5197);
nand U6751 (N_6751,N_5900,N_5211);
nor U6752 (N_6752,N_5336,N_5860);
or U6753 (N_6753,N_5589,N_5342);
nor U6754 (N_6754,N_5190,N_5620);
or U6755 (N_6755,N_5296,N_5811);
xor U6756 (N_6756,N_5929,N_5060);
or U6757 (N_6757,N_5230,N_5459);
xnor U6758 (N_6758,N_5849,N_5276);
nand U6759 (N_6759,N_5652,N_5858);
nand U6760 (N_6760,N_5556,N_5292);
nor U6761 (N_6761,N_5941,N_5268);
and U6762 (N_6762,N_5564,N_5434);
or U6763 (N_6763,N_5451,N_5590);
or U6764 (N_6764,N_5702,N_5073);
nor U6765 (N_6765,N_5767,N_5373);
nor U6766 (N_6766,N_5127,N_5447);
and U6767 (N_6767,N_5221,N_5165);
nand U6768 (N_6768,N_5130,N_5445);
or U6769 (N_6769,N_5704,N_5181);
nor U6770 (N_6770,N_5115,N_5907);
nor U6771 (N_6771,N_5301,N_5384);
and U6772 (N_6772,N_5297,N_5232);
nand U6773 (N_6773,N_5946,N_5455);
or U6774 (N_6774,N_5936,N_5069);
or U6775 (N_6775,N_5845,N_5041);
nand U6776 (N_6776,N_5872,N_5820);
nand U6777 (N_6777,N_5501,N_5661);
xnor U6778 (N_6778,N_5977,N_5749);
nor U6779 (N_6779,N_5441,N_5300);
or U6780 (N_6780,N_5640,N_5599);
nand U6781 (N_6781,N_5954,N_5341);
nand U6782 (N_6782,N_5757,N_5856);
nor U6783 (N_6783,N_5977,N_5330);
nand U6784 (N_6784,N_5182,N_5537);
and U6785 (N_6785,N_5406,N_5820);
and U6786 (N_6786,N_5065,N_5008);
nor U6787 (N_6787,N_5673,N_5105);
nor U6788 (N_6788,N_5877,N_5191);
xnor U6789 (N_6789,N_5993,N_5965);
nand U6790 (N_6790,N_5787,N_5327);
xnor U6791 (N_6791,N_5059,N_5284);
nor U6792 (N_6792,N_5153,N_5464);
nand U6793 (N_6793,N_5600,N_5971);
xnor U6794 (N_6794,N_5054,N_5446);
and U6795 (N_6795,N_5665,N_5234);
nand U6796 (N_6796,N_5438,N_5268);
nand U6797 (N_6797,N_5953,N_5460);
and U6798 (N_6798,N_5997,N_5661);
nand U6799 (N_6799,N_5842,N_5436);
nand U6800 (N_6800,N_5204,N_5788);
nor U6801 (N_6801,N_5611,N_5100);
nor U6802 (N_6802,N_5906,N_5281);
xnor U6803 (N_6803,N_5476,N_5171);
and U6804 (N_6804,N_5413,N_5294);
nor U6805 (N_6805,N_5406,N_5364);
nand U6806 (N_6806,N_5911,N_5688);
or U6807 (N_6807,N_5066,N_5277);
nand U6808 (N_6808,N_5728,N_5261);
and U6809 (N_6809,N_5160,N_5851);
nor U6810 (N_6810,N_5717,N_5168);
or U6811 (N_6811,N_5418,N_5537);
or U6812 (N_6812,N_5256,N_5879);
or U6813 (N_6813,N_5524,N_5050);
nand U6814 (N_6814,N_5792,N_5546);
nand U6815 (N_6815,N_5775,N_5570);
nor U6816 (N_6816,N_5742,N_5570);
or U6817 (N_6817,N_5508,N_5037);
and U6818 (N_6818,N_5660,N_5651);
nor U6819 (N_6819,N_5550,N_5028);
or U6820 (N_6820,N_5181,N_5498);
nor U6821 (N_6821,N_5028,N_5313);
and U6822 (N_6822,N_5424,N_5258);
nand U6823 (N_6823,N_5692,N_5523);
nor U6824 (N_6824,N_5899,N_5658);
and U6825 (N_6825,N_5713,N_5238);
and U6826 (N_6826,N_5689,N_5926);
xnor U6827 (N_6827,N_5296,N_5864);
nand U6828 (N_6828,N_5273,N_5457);
or U6829 (N_6829,N_5405,N_5042);
and U6830 (N_6830,N_5173,N_5495);
nor U6831 (N_6831,N_5935,N_5125);
nor U6832 (N_6832,N_5859,N_5593);
xnor U6833 (N_6833,N_5737,N_5669);
xnor U6834 (N_6834,N_5194,N_5170);
nand U6835 (N_6835,N_5094,N_5586);
xnor U6836 (N_6836,N_5442,N_5681);
nor U6837 (N_6837,N_5282,N_5539);
and U6838 (N_6838,N_5073,N_5097);
and U6839 (N_6839,N_5488,N_5779);
or U6840 (N_6840,N_5810,N_5310);
and U6841 (N_6841,N_5666,N_5125);
and U6842 (N_6842,N_5788,N_5249);
nand U6843 (N_6843,N_5600,N_5626);
or U6844 (N_6844,N_5880,N_5419);
nor U6845 (N_6845,N_5509,N_5024);
xor U6846 (N_6846,N_5712,N_5315);
nand U6847 (N_6847,N_5387,N_5764);
nand U6848 (N_6848,N_5104,N_5787);
nand U6849 (N_6849,N_5400,N_5144);
and U6850 (N_6850,N_5484,N_5079);
or U6851 (N_6851,N_5321,N_5172);
nor U6852 (N_6852,N_5600,N_5642);
or U6853 (N_6853,N_5350,N_5612);
and U6854 (N_6854,N_5216,N_5492);
and U6855 (N_6855,N_5796,N_5471);
xor U6856 (N_6856,N_5776,N_5799);
and U6857 (N_6857,N_5720,N_5227);
or U6858 (N_6858,N_5579,N_5518);
or U6859 (N_6859,N_5377,N_5320);
nor U6860 (N_6860,N_5474,N_5718);
and U6861 (N_6861,N_5584,N_5264);
nand U6862 (N_6862,N_5075,N_5687);
and U6863 (N_6863,N_5094,N_5547);
and U6864 (N_6864,N_5336,N_5474);
and U6865 (N_6865,N_5960,N_5115);
or U6866 (N_6866,N_5063,N_5935);
xor U6867 (N_6867,N_5776,N_5329);
and U6868 (N_6868,N_5437,N_5365);
nor U6869 (N_6869,N_5055,N_5416);
nand U6870 (N_6870,N_5770,N_5528);
or U6871 (N_6871,N_5400,N_5851);
nor U6872 (N_6872,N_5883,N_5912);
and U6873 (N_6873,N_5704,N_5144);
and U6874 (N_6874,N_5886,N_5468);
and U6875 (N_6875,N_5903,N_5616);
nand U6876 (N_6876,N_5234,N_5536);
nor U6877 (N_6877,N_5019,N_5809);
nor U6878 (N_6878,N_5160,N_5294);
or U6879 (N_6879,N_5874,N_5048);
and U6880 (N_6880,N_5649,N_5578);
or U6881 (N_6881,N_5382,N_5978);
xnor U6882 (N_6882,N_5381,N_5295);
xnor U6883 (N_6883,N_5124,N_5753);
or U6884 (N_6884,N_5058,N_5928);
nor U6885 (N_6885,N_5736,N_5295);
nor U6886 (N_6886,N_5130,N_5312);
or U6887 (N_6887,N_5775,N_5609);
nor U6888 (N_6888,N_5036,N_5444);
and U6889 (N_6889,N_5690,N_5530);
nand U6890 (N_6890,N_5457,N_5558);
or U6891 (N_6891,N_5768,N_5867);
nand U6892 (N_6892,N_5602,N_5538);
or U6893 (N_6893,N_5851,N_5673);
or U6894 (N_6894,N_5597,N_5001);
xor U6895 (N_6895,N_5031,N_5081);
nand U6896 (N_6896,N_5844,N_5016);
or U6897 (N_6897,N_5422,N_5265);
nand U6898 (N_6898,N_5635,N_5232);
nand U6899 (N_6899,N_5696,N_5685);
or U6900 (N_6900,N_5882,N_5224);
nor U6901 (N_6901,N_5559,N_5172);
and U6902 (N_6902,N_5206,N_5208);
nand U6903 (N_6903,N_5912,N_5111);
nand U6904 (N_6904,N_5641,N_5544);
nand U6905 (N_6905,N_5311,N_5552);
nand U6906 (N_6906,N_5443,N_5516);
nor U6907 (N_6907,N_5657,N_5451);
nor U6908 (N_6908,N_5961,N_5156);
nor U6909 (N_6909,N_5374,N_5271);
nand U6910 (N_6910,N_5095,N_5650);
or U6911 (N_6911,N_5638,N_5856);
and U6912 (N_6912,N_5826,N_5788);
or U6913 (N_6913,N_5146,N_5965);
xnor U6914 (N_6914,N_5886,N_5753);
or U6915 (N_6915,N_5968,N_5195);
nor U6916 (N_6916,N_5621,N_5604);
nor U6917 (N_6917,N_5868,N_5152);
nor U6918 (N_6918,N_5525,N_5577);
or U6919 (N_6919,N_5140,N_5604);
nand U6920 (N_6920,N_5322,N_5277);
nor U6921 (N_6921,N_5371,N_5784);
or U6922 (N_6922,N_5308,N_5649);
or U6923 (N_6923,N_5294,N_5816);
or U6924 (N_6924,N_5975,N_5259);
nand U6925 (N_6925,N_5312,N_5417);
nand U6926 (N_6926,N_5008,N_5195);
or U6927 (N_6927,N_5481,N_5755);
or U6928 (N_6928,N_5993,N_5052);
nor U6929 (N_6929,N_5108,N_5201);
nor U6930 (N_6930,N_5241,N_5424);
or U6931 (N_6931,N_5331,N_5775);
and U6932 (N_6932,N_5788,N_5512);
or U6933 (N_6933,N_5731,N_5803);
nand U6934 (N_6934,N_5732,N_5818);
or U6935 (N_6935,N_5541,N_5958);
and U6936 (N_6936,N_5723,N_5261);
and U6937 (N_6937,N_5802,N_5739);
and U6938 (N_6938,N_5523,N_5066);
nand U6939 (N_6939,N_5348,N_5484);
xor U6940 (N_6940,N_5128,N_5104);
xnor U6941 (N_6941,N_5959,N_5991);
and U6942 (N_6942,N_5672,N_5700);
and U6943 (N_6943,N_5705,N_5061);
nand U6944 (N_6944,N_5833,N_5324);
nand U6945 (N_6945,N_5535,N_5530);
or U6946 (N_6946,N_5503,N_5267);
xor U6947 (N_6947,N_5557,N_5486);
nor U6948 (N_6948,N_5353,N_5032);
or U6949 (N_6949,N_5561,N_5116);
xnor U6950 (N_6950,N_5567,N_5485);
nor U6951 (N_6951,N_5928,N_5031);
or U6952 (N_6952,N_5162,N_5387);
nand U6953 (N_6953,N_5749,N_5128);
and U6954 (N_6954,N_5069,N_5456);
or U6955 (N_6955,N_5989,N_5896);
or U6956 (N_6956,N_5083,N_5555);
and U6957 (N_6957,N_5954,N_5484);
or U6958 (N_6958,N_5278,N_5296);
nand U6959 (N_6959,N_5329,N_5536);
nand U6960 (N_6960,N_5595,N_5515);
nand U6961 (N_6961,N_5258,N_5955);
nand U6962 (N_6962,N_5409,N_5837);
and U6963 (N_6963,N_5438,N_5718);
or U6964 (N_6964,N_5090,N_5744);
nor U6965 (N_6965,N_5545,N_5485);
or U6966 (N_6966,N_5221,N_5838);
nor U6967 (N_6967,N_5000,N_5453);
xor U6968 (N_6968,N_5115,N_5788);
nor U6969 (N_6969,N_5745,N_5209);
xor U6970 (N_6970,N_5748,N_5550);
nand U6971 (N_6971,N_5574,N_5524);
or U6972 (N_6972,N_5040,N_5858);
nand U6973 (N_6973,N_5136,N_5375);
xnor U6974 (N_6974,N_5160,N_5771);
or U6975 (N_6975,N_5507,N_5603);
and U6976 (N_6976,N_5991,N_5033);
and U6977 (N_6977,N_5206,N_5590);
nor U6978 (N_6978,N_5172,N_5460);
nand U6979 (N_6979,N_5763,N_5617);
or U6980 (N_6980,N_5961,N_5708);
and U6981 (N_6981,N_5594,N_5718);
or U6982 (N_6982,N_5352,N_5054);
nor U6983 (N_6983,N_5465,N_5608);
or U6984 (N_6984,N_5693,N_5536);
or U6985 (N_6985,N_5544,N_5441);
and U6986 (N_6986,N_5886,N_5955);
nand U6987 (N_6987,N_5951,N_5028);
or U6988 (N_6988,N_5516,N_5147);
and U6989 (N_6989,N_5967,N_5888);
nor U6990 (N_6990,N_5949,N_5034);
or U6991 (N_6991,N_5752,N_5585);
xor U6992 (N_6992,N_5112,N_5382);
or U6993 (N_6993,N_5904,N_5037);
nor U6994 (N_6994,N_5037,N_5583);
nor U6995 (N_6995,N_5645,N_5867);
nand U6996 (N_6996,N_5676,N_5193);
xor U6997 (N_6997,N_5398,N_5993);
nand U6998 (N_6998,N_5109,N_5609);
nand U6999 (N_6999,N_5375,N_5317);
or U7000 (N_7000,N_6577,N_6284);
and U7001 (N_7001,N_6571,N_6775);
nand U7002 (N_7002,N_6424,N_6715);
nand U7003 (N_7003,N_6903,N_6902);
or U7004 (N_7004,N_6745,N_6847);
nor U7005 (N_7005,N_6696,N_6261);
nor U7006 (N_7006,N_6033,N_6385);
or U7007 (N_7007,N_6782,N_6206);
nand U7008 (N_7008,N_6429,N_6087);
nor U7009 (N_7009,N_6014,N_6403);
or U7010 (N_7010,N_6949,N_6938);
or U7011 (N_7011,N_6232,N_6740);
nor U7012 (N_7012,N_6107,N_6088);
or U7013 (N_7013,N_6720,N_6807);
or U7014 (N_7014,N_6305,N_6558);
or U7015 (N_7015,N_6130,N_6515);
nor U7016 (N_7016,N_6254,N_6115);
or U7017 (N_7017,N_6164,N_6648);
nor U7018 (N_7018,N_6564,N_6679);
nor U7019 (N_7019,N_6652,N_6205);
or U7020 (N_7020,N_6849,N_6327);
xor U7021 (N_7021,N_6478,N_6230);
and U7022 (N_7022,N_6127,N_6494);
or U7023 (N_7023,N_6560,N_6905);
nand U7024 (N_7024,N_6279,N_6591);
xnor U7025 (N_7025,N_6021,N_6645);
and U7026 (N_7026,N_6883,N_6774);
and U7027 (N_7027,N_6855,N_6813);
nor U7028 (N_7028,N_6104,N_6751);
and U7029 (N_7029,N_6147,N_6910);
or U7030 (N_7030,N_6935,N_6892);
nor U7031 (N_7031,N_6603,N_6208);
nand U7032 (N_7032,N_6395,N_6341);
nand U7033 (N_7033,N_6166,N_6349);
and U7034 (N_7034,N_6729,N_6983);
xnor U7035 (N_7035,N_6225,N_6643);
nand U7036 (N_7036,N_6201,N_6943);
nor U7037 (N_7037,N_6476,N_6725);
or U7038 (N_7038,N_6499,N_6960);
and U7039 (N_7039,N_6777,N_6522);
and U7040 (N_7040,N_6997,N_6796);
and U7041 (N_7041,N_6037,N_6992);
nand U7042 (N_7042,N_6797,N_6419);
or U7043 (N_7043,N_6788,N_6831);
and U7044 (N_7044,N_6452,N_6183);
and U7045 (N_7045,N_6704,N_6714);
and U7046 (N_7046,N_6890,N_6680);
nand U7047 (N_7047,N_6133,N_6152);
nand U7048 (N_7048,N_6787,N_6393);
and U7049 (N_7049,N_6302,N_6095);
nand U7050 (N_7050,N_6283,N_6271);
and U7051 (N_7051,N_6655,N_6574);
xor U7052 (N_7052,N_6102,N_6042);
or U7053 (N_7053,N_6776,N_6894);
or U7054 (N_7054,N_6288,N_6337);
and U7055 (N_7055,N_6212,N_6243);
and U7056 (N_7056,N_6396,N_6218);
or U7057 (N_7057,N_6669,N_6540);
or U7058 (N_7058,N_6402,N_6688);
nand U7059 (N_7059,N_6245,N_6372);
and U7060 (N_7060,N_6580,N_6052);
or U7061 (N_7061,N_6320,N_6398);
or U7062 (N_7062,N_6013,N_6599);
nand U7063 (N_7063,N_6015,N_6238);
and U7064 (N_7064,N_6755,N_6300);
nor U7065 (N_7065,N_6982,N_6771);
and U7066 (N_7066,N_6213,N_6623);
and U7067 (N_7067,N_6597,N_6695);
nand U7068 (N_7068,N_6416,N_6074);
nand U7069 (N_7069,N_6163,N_6445);
xnor U7070 (N_7070,N_6518,N_6073);
nand U7071 (N_7071,N_6672,N_6861);
nor U7072 (N_7072,N_6301,N_6091);
and U7073 (N_7073,N_6140,N_6195);
and U7074 (N_7074,N_6611,N_6519);
nand U7075 (N_7075,N_6219,N_6584);
xnor U7076 (N_7076,N_6871,N_6743);
xnor U7077 (N_7077,N_6008,N_6728);
xnor U7078 (N_7078,N_6646,N_6931);
or U7079 (N_7079,N_6204,N_6589);
or U7080 (N_7080,N_6532,N_6523);
nand U7081 (N_7081,N_6985,N_6436);
and U7082 (N_7082,N_6870,N_6733);
and U7083 (N_7083,N_6827,N_6474);
and U7084 (N_7084,N_6785,N_6566);
and U7085 (N_7085,N_6613,N_6790);
or U7086 (N_7086,N_6826,N_6141);
nand U7087 (N_7087,N_6348,N_6925);
nor U7088 (N_7088,N_6984,N_6318);
nand U7089 (N_7089,N_6241,N_6820);
nand U7090 (N_7090,N_6904,N_6131);
xor U7091 (N_7091,N_6634,N_6585);
nand U7092 (N_7092,N_6717,N_6362);
or U7093 (N_7093,N_6530,N_6723);
and U7094 (N_7094,N_6379,N_6897);
nand U7095 (N_7095,N_6350,N_6588);
and U7096 (N_7096,N_6959,N_6307);
or U7097 (N_7097,N_6422,N_6628);
or U7098 (N_7098,N_6525,N_6375);
and U7099 (N_7099,N_6442,N_6490);
and U7100 (N_7100,N_6946,N_6435);
xor U7101 (N_7101,N_6587,N_6317);
xnor U7102 (N_7102,N_6411,N_6630);
or U7103 (N_7103,N_6291,N_6251);
and U7104 (N_7104,N_6962,N_6330);
or U7105 (N_7105,N_6868,N_6413);
nand U7106 (N_7106,N_6917,N_6150);
nor U7107 (N_7107,N_6760,N_6712);
nand U7108 (N_7108,N_6080,N_6296);
and U7109 (N_7109,N_6889,N_6814);
or U7110 (N_7110,N_6576,N_6344);
or U7111 (N_7111,N_6865,N_6686);
nand U7112 (N_7112,N_6404,N_6573);
nor U7113 (N_7113,N_6101,N_6980);
xnor U7114 (N_7114,N_6867,N_6108);
and U7115 (N_7115,N_6508,N_6612);
nor U7116 (N_7116,N_6399,N_6031);
and U7117 (N_7117,N_6321,N_6227);
and U7118 (N_7118,N_6264,N_6465);
and U7119 (N_7119,N_6900,N_6893);
and U7120 (N_7120,N_6338,N_6516);
and U7121 (N_7121,N_6778,N_6840);
nand U7122 (N_7122,N_6352,N_6124);
or U7123 (N_7123,N_6637,N_6884);
and U7124 (N_7124,N_6551,N_6644);
or U7125 (N_7125,N_6501,N_6114);
or U7126 (N_7126,N_6026,N_6081);
nor U7127 (N_7127,N_6622,N_6561);
or U7128 (N_7128,N_6666,N_6376);
or U7129 (N_7129,N_6640,N_6565);
nand U7130 (N_7130,N_6387,N_6038);
and U7131 (N_7131,N_6810,N_6981);
or U7132 (N_7132,N_6449,N_6872);
or U7133 (N_7133,N_6312,N_6194);
or U7134 (N_7134,N_6484,N_6651);
and U7135 (N_7135,N_6016,N_6632);
xnor U7136 (N_7136,N_6489,N_6151);
nor U7137 (N_7137,N_6702,N_6443);
xnor U7138 (N_7138,N_6400,N_6236);
nand U7139 (N_7139,N_6899,N_6239);
nor U7140 (N_7140,N_6873,N_6996);
xor U7141 (N_7141,N_6991,N_6039);
or U7142 (N_7142,N_6267,N_6001);
nand U7143 (N_7143,N_6964,N_6846);
nor U7144 (N_7144,N_6377,N_6477);
or U7145 (N_7145,N_6405,N_6950);
and U7146 (N_7146,N_6111,N_6196);
or U7147 (N_7147,N_6380,N_6117);
nand U7148 (N_7148,N_6223,N_6093);
and U7149 (N_7149,N_6731,N_6426);
or U7150 (N_7150,N_6019,N_6944);
xor U7151 (N_7151,N_6285,N_6216);
nand U7152 (N_7152,N_6521,N_6410);
nor U7153 (N_7153,N_6756,N_6542);
or U7154 (N_7154,N_6830,N_6520);
and U7155 (N_7155,N_6467,N_6973);
nor U7156 (N_7156,N_6248,N_6649);
xor U7157 (N_7157,N_6010,N_6783);
nor U7158 (N_7158,N_6311,N_6050);
nor U7159 (N_7159,N_6674,N_6915);
nor U7160 (N_7160,N_6498,N_6392);
nand U7161 (N_7161,N_6553,N_6535);
and U7162 (N_7162,N_6441,N_6358);
nor U7163 (N_7163,N_6907,N_6684);
nor U7164 (N_7164,N_6631,N_6313);
or U7165 (N_7165,N_6281,N_6968);
nor U7166 (N_7166,N_6186,N_6444);
nor U7167 (N_7167,N_6616,N_6138);
or U7168 (N_7168,N_6541,N_6382);
and U7169 (N_7169,N_6058,N_6838);
xnor U7170 (N_7170,N_6466,N_6180);
xor U7171 (N_7171,N_6278,N_6149);
nand U7172 (N_7172,N_6823,N_6062);
nand U7173 (N_7173,N_6852,N_6664);
nor U7174 (N_7174,N_6993,N_6594);
nor U7175 (N_7175,N_6537,N_6182);
nand U7176 (N_7176,N_6389,N_6303);
nor U7177 (N_7177,N_6753,N_6076);
and U7178 (N_7178,N_6043,N_6425);
nand U7179 (N_7179,N_6965,N_6974);
and U7180 (N_7180,N_6896,N_6171);
nor U7181 (N_7181,N_6675,N_6447);
nor U7182 (N_7182,N_6136,N_6512);
nor U7183 (N_7183,N_6825,N_6579);
and U7184 (N_7184,N_6332,N_6682);
xnor U7185 (N_7185,N_6713,N_6668);
nand U7186 (N_7186,N_6134,N_6233);
or U7187 (N_7187,N_6657,N_6257);
nand U7188 (N_7188,N_6707,N_6086);
nand U7189 (N_7189,N_6027,N_6761);
and U7190 (N_7190,N_6005,N_6249);
nor U7191 (N_7191,N_6878,N_6568);
and U7192 (N_7192,N_6507,N_6608);
and U7193 (N_7193,N_6642,N_6315);
xnor U7194 (N_7194,N_6011,N_6698);
nand U7195 (N_7195,N_6866,N_6534);
nor U7196 (N_7196,N_6070,N_6921);
nor U7197 (N_7197,N_6650,N_6420);
or U7198 (N_7198,N_6110,N_6699);
nor U7199 (N_7199,N_6654,N_6364);
nor U7200 (N_7200,N_6978,N_6527);
nor U7201 (N_7201,N_6482,N_6408);
and U7202 (N_7202,N_6353,N_6770);
or U7203 (N_7203,N_6839,N_6132);
and U7204 (N_7204,N_6609,N_6809);
and U7205 (N_7205,N_6113,N_6298);
and U7206 (N_7206,N_6438,N_6924);
nand U7207 (N_7207,N_6295,N_6750);
nand U7208 (N_7208,N_6843,N_6224);
or U7209 (N_7209,N_6184,N_6463);
or U7210 (N_7210,N_6817,N_6805);
nor U7211 (N_7211,N_6605,N_6162);
and U7212 (N_7212,N_6531,N_6667);
nand U7213 (N_7213,N_6383,N_6635);
and U7214 (N_7214,N_6493,N_6898);
nand U7215 (N_7215,N_6369,N_6895);
nand U7216 (N_7216,N_6055,N_6240);
nand U7217 (N_7217,N_6044,N_6386);
or U7218 (N_7218,N_6880,N_6693);
nand U7219 (N_7219,N_6173,N_6144);
nor U7220 (N_7220,N_6203,N_6148);
and U7221 (N_7221,N_6409,N_6908);
or U7222 (N_7222,N_6316,N_6459);
or U7223 (N_7223,N_6671,N_6549);
nand U7224 (N_7224,N_6097,N_6112);
nand U7225 (N_7225,N_6948,N_6262);
and U7226 (N_7226,N_6781,N_6911);
and U7227 (N_7227,N_6954,N_6069);
and U7228 (N_7228,N_6933,N_6828);
nand U7229 (N_7229,N_6263,N_6439);
nand U7230 (N_7230,N_6177,N_6546);
xnor U7231 (N_7231,N_6990,N_6373);
or U7232 (N_7232,N_6887,N_6100);
and U7233 (N_7233,N_6582,N_6142);
and U7234 (N_7234,N_6617,N_6638);
nand U7235 (N_7235,N_6235,N_6129);
and U7236 (N_7236,N_6876,N_6356);
nor U7237 (N_7237,N_6421,N_6747);
and U7238 (N_7238,N_6381,N_6256);
and U7239 (N_7239,N_6446,N_6034);
nand U7240 (N_7240,N_6060,N_6246);
nand U7241 (N_7241,N_6673,N_6615);
xor U7242 (N_7242,N_6461,N_6290);
and U7243 (N_7243,N_6504,N_6601);
nor U7244 (N_7244,N_6165,N_6816);
or U7245 (N_7245,N_6388,N_6976);
nor U7246 (N_7246,N_6139,N_6986);
nand U7247 (N_7247,N_6346,N_6685);
or U7248 (N_7248,N_6928,N_6094);
and U7249 (N_7249,N_6539,N_6071);
nor U7250 (N_7250,N_6106,N_6934);
and U7251 (N_7251,N_6047,N_6691);
and U7252 (N_7252,N_6853,N_6629);
nor U7253 (N_7253,N_6914,N_6727);
xnor U7254 (N_7254,N_6122,N_6319);
nor U7255 (N_7255,N_6120,N_6118);
or U7256 (N_7256,N_6592,N_6187);
nand U7257 (N_7257,N_6475,N_6123);
or U7258 (N_7258,N_6175,N_6423);
and U7259 (N_7259,N_6090,N_6741);
or U7260 (N_7260,N_6503,N_6193);
nor U7261 (N_7261,N_6277,N_6406);
nor U7262 (N_7262,N_6456,N_6524);
or U7263 (N_7263,N_6683,N_6735);
nor U7264 (N_7264,N_6333,N_6738);
nand U7265 (N_7265,N_6412,N_6430);
or U7266 (N_7266,N_6951,N_6862);
nand U7267 (N_7267,N_6331,N_6252);
nand U7268 (N_7268,N_6222,N_6082);
or U7269 (N_7269,N_6431,N_6721);
nor U7270 (N_7270,N_6701,N_6098);
nor U7271 (N_7271,N_6460,N_6567);
or U7272 (N_7272,N_6719,N_6229);
and U7273 (N_7273,N_6266,N_6936);
nand U7274 (N_7274,N_6197,N_6875);
nand U7275 (N_7275,N_6939,N_6084);
or U7276 (N_7276,N_6153,N_6178);
nor U7277 (N_7277,N_6029,N_6024);
and U7278 (N_7278,N_6326,N_6660);
nor U7279 (N_7279,N_6586,N_6784);
or U7280 (N_7280,N_6077,N_6795);
xnor U7281 (N_7281,N_6168,N_6665);
or U7282 (N_7282,N_6545,N_6414);
and U7283 (N_7283,N_6979,N_6506);
or U7284 (N_7284,N_6351,N_6786);
and U7285 (N_7285,N_6590,N_6803);
and U7286 (N_7286,N_6607,N_6920);
nand U7287 (N_7287,N_6842,N_6036);
nand U7288 (N_7288,N_6470,N_6121);
nand U7289 (N_7289,N_6211,N_6103);
nor U7290 (N_7290,N_6970,N_6995);
or U7291 (N_7291,N_6496,N_6157);
xor U7292 (N_7292,N_6799,N_6517);
xor U7293 (N_7293,N_6502,N_6200);
nand U7294 (N_7294,N_6835,N_6739);
or U7295 (N_7295,N_6054,N_6155);
and U7296 (N_7296,N_6538,N_6472);
and U7297 (N_7297,N_6918,N_6763);
or U7298 (N_7298,N_6032,N_6972);
nor U7299 (N_7299,N_6837,N_6017);
or U7300 (N_7300,N_6730,N_6068);
nand U7301 (N_7301,N_6336,N_6174);
xnor U7302 (N_7302,N_6209,N_6045);
nand U7303 (N_7303,N_6947,N_6602);
nand U7304 (N_7304,N_6215,N_6806);
and U7305 (N_7305,N_6793,N_6007);
nand U7306 (N_7306,N_6022,N_6916);
nand U7307 (N_7307,N_6929,N_6237);
nand U7308 (N_7308,N_6250,N_6244);
and U7309 (N_7309,N_6334,N_6772);
nand U7310 (N_7310,N_6692,N_6955);
nand U7311 (N_7311,N_6716,N_6457);
nor U7312 (N_7312,N_6641,N_6159);
nor U7313 (N_7313,N_6626,N_6768);
and U7314 (N_7314,N_6766,N_6304);
or U7315 (N_7315,N_6308,N_6614);
nor U7316 (N_7316,N_6354,N_6879);
nand U7317 (N_7317,N_6083,N_6548);
and U7318 (N_7318,N_6006,N_6374);
and U7319 (N_7319,N_6427,N_6802);
and U7320 (N_7320,N_6670,N_6000);
nor U7321 (N_7321,N_6309,N_6002);
and U7322 (N_7322,N_6048,N_6176);
nor U7323 (N_7323,N_6851,N_6273);
nand U7324 (N_7324,N_6046,N_6618);
and U7325 (N_7325,N_6289,N_6845);
nand U7326 (N_7326,N_6736,N_6468);
nand U7327 (N_7327,N_6848,N_6505);
nor U7328 (N_7328,N_6051,N_6335);
xnor U7329 (N_7329,N_6957,N_6578);
nor U7330 (N_7330,N_6694,N_6479);
or U7331 (N_7331,N_6247,N_6690);
xnor U7332 (N_7332,N_6119,N_6368);
and U7333 (N_7333,N_6292,N_6661);
nand U7334 (N_7334,N_6495,N_6156);
nand U7335 (N_7335,N_6804,N_6299);
nand U7336 (N_7336,N_6562,N_6625);
nor U7337 (N_7337,N_6759,N_6025);
nor U7338 (N_7338,N_6528,N_6179);
nand U7339 (N_7339,N_6663,N_6620);
nand U7340 (N_7340,N_6836,N_6514);
nor U7341 (N_7341,N_6886,N_6869);
and U7342 (N_7342,N_6481,N_6035);
or U7343 (N_7343,N_6882,N_6480);
nand U7344 (N_7344,N_6259,N_6780);
nor U7345 (N_7345,N_6658,N_6742);
and U7346 (N_7346,N_6529,N_6994);
and U7347 (N_7347,N_6687,N_6293);
nor U7348 (N_7348,N_6606,N_6390);
nor U7349 (N_7349,N_6509,N_6863);
xnor U7350 (N_7350,N_6619,N_6555);
nor U7351 (N_7351,N_6056,N_6483);
nand U7352 (N_7352,N_6202,N_6627);
nand U7353 (N_7353,N_6394,N_6199);
or U7354 (N_7354,N_6487,N_6593);
nand U7355 (N_7355,N_6563,N_6343);
nand U7356 (N_7356,N_6064,N_6049);
and U7357 (N_7357,N_6231,N_6109);
nor U7358 (N_7358,N_6340,N_6988);
and U7359 (N_7359,N_6513,N_6407);
nand U7360 (N_7360,N_6569,N_6057);
and U7361 (N_7361,N_6361,N_6966);
nor U7362 (N_7362,N_6536,N_6473);
xor U7363 (N_7363,N_6217,N_6434);
or U7364 (N_7364,N_6072,N_6912);
nand U7365 (N_7365,N_6061,N_6856);
and U7366 (N_7366,N_6734,N_6488);
and U7367 (N_7367,N_6418,N_6926);
nand U7368 (N_7368,N_6556,N_6089);
nand U7369 (N_7369,N_6927,N_6595);
xor U7370 (N_7370,N_6137,N_6314);
and U7371 (N_7371,N_6794,N_6697);
xor U7372 (N_7372,N_6749,N_6877);
nand U7373 (N_7373,N_6276,N_6711);
or U7374 (N_7374,N_6722,N_6269);
and U7375 (N_7375,N_6339,N_6167);
nand U7376 (N_7376,N_6226,N_6812);
and U7377 (N_7377,N_6919,N_6428);
nand U7378 (N_7378,N_6365,N_6030);
nor U7379 (N_7379,N_6758,N_6829);
nand U7380 (N_7380,N_6710,N_6066);
xnor U7381 (N_7381,N_6700,N_6891);
xor U7382 (N_7382,N_6359,N_6708);
nor U7383 (N_7383,N_6448,N_6018);
nand U7384 (N_7384,N_6681,N_6085);
xor U7385 (N_7385,N_6961,N_6450);
and U7386 (N_7386,N_6078,N_6258);
or U7387 (N_7387,N_6306,N_6378);
or U7388 (N_7388,N_6347,N_6185);
nor U7389 (N_7389,N_6922,N_6440);
nor U7390 (N_7390,N_6366,N_6188);
or U7391 (N_7391,N_6371,N_6345);
and U7392 (N_7392,N_6492,N_6547);
or U7393 (N_7393,N_6329,N_6706);
nor U7394 (N_7394,N_6647,N_6971);
and U7395 (N_7395,N_6397,N_6937);
or U7396 (N_7396,N_6901,N_6987);
nand U7397 (N_7397,N_6063,N_6989);
nand U7398 (N_7398,N_6275,N_6214);
nand U7399 (N_7399,N_6952,N_6821);
nand U7400 (N_7400,N_6822,N_6059);
and U7401 (N_7401,N_6497,N_6065);
and U7402 (N_7402,N_6486,N_6909);
or U7403 (N_7403,N_6105,N_6287);
or U7404 (N_7404,N_6570,N_6041);
nor U7405 (N_7405,N_6432,N_6881);
nor U7406 (N_7406,N_6181,N_6945);
nor U7407 (N_7407,N_6092,N_6834);
xor U7408 (N_7408,N_6621,N_6415);
or U7409 (N_7409,N_6930,N_6145);
nand U7410 (N_7410,N_6533,N_6744);
and U7411 (N_7411,N_6575,N_6940);
and U7412 (N_7412,N_6004,N_6757);
and U7413 (N_7413,N_6659,N_6454);
nor U7414 (N_7414,N_6557,N_6458);
nand U7415 (N_7415,N_6913,N_6818);
nor U7416 (N_7416,N_6732,N_6737);
nor U7417 (N_7417,N_6748,N_6769);
nor U7418 (N_7418,N_6864,N_6135);
nand U7419 (N_7419,N_6656,N_6453);
and U7420 (N_7420,N_6255,N_6850);
and U7421 (N_7421,N_6128,N_6154);
or U7422 (N_7422,N_6357,N_6272);
and U7423 (N_7423,N_6462,N_6554);
and U7424 (N_7424,N_6328,N_6469);
or U7425 (N_7425,N_6800,N_6234);
nor U7426 (N_7426,N_6798,N_6689);
or U7427 (N_7427,N_6511,N_6819);
and U7428 (N_7428,N_6367,N_6324);
nand U7429 (N_7429,N_6491,N_6859);
nand U7430 (N_7430,N_6792,N_6815);
and U7431 (N_7431,N_6791,N_6040);
nor U7432 (N_7432,N_6762,N_6274);
nor U7433 (N_7433,N_6779,N_6221);
or U7434 (N_7434,N_6999,N_6242);
and U7435 (N_7435,N_6633,N_6752);
nor U7436 (N_7436,N_6636,N_6604);
and U7437 (N_7437,N_6801,N_6764);
and U7438 (N_7438,N_6464,N_6009);
and U7439 (N_7439,N_6220,N_6559);
xnor U7440 (N_7440,N_6360,N_6370);
and U7441 (N_7441,N_6550,N_6485);
nand U7442 (N_7442,N_6260,N_6923);
and U7443 (N_7443,N_6500,N_6012);
or U7444 (N_7444,N_6941,N_6169);
nand U7445 (N_7445,N_6191,N_6280);
nor U7446 (N_7446,N_6726,N_6526);
or U7447 (N_7447,N_6906,N_6265);
nor U7448 (N_7448,N_6653,N_6583);
nor U7449 (N_7449,N_6437,N_6958);
and U7450 (N_7450,N_6841,N_6355);
nor U7451 (N_7451,N_6967,N_6067);
nor U7452 (N_7452,N_6170,N_6746);
nand U7453 (N_7453,N_6451,N_6857);
nand U7454 (N_7454,N_6833,N_6192);
and U7455 (N_7455,N_6600,N_6172);
nand U7456 (N_7456,N_6767,N_6297);
nand U7457 (N_7457,N_6322,N_6754);
nand U7458 (N_7458,N_6718,N_6096);
nor U7459 (N_7459,N_6323,N_6189);
or U7460 (N_7460,N_6789,N_6268);
nor U7461 (N_7461,N_6510,N_6932);
or U7462 (N_7462,N_6342,N_6858);
nor U7463 (N_7463,N_6676,N_6126);
nand U7464 (N_7464,N_6003,N_6998);
and U7465 (N_7465,N_6270,N_6190);
nand U7466 (N_7466,N_6610,N_6158);
or U7467 (N_7467,N_6099,N_6854);
nor U7468 (N_7468,N_6956,N_6160);
and U7469 (N_7469,N_6662,N_6384);
or U7470 (N_7470,N_6310,N_6028);
xor U7471 (N_7471,N_6765,N_6210);
xor U7472 (N_7472,N_6860,N_6598);
or U7473 (N_7473,N_6709,N_6143);
or U7474 (N_7474,N_6401,N_6161);
nor U7475 (N_7475,N_6953,N_6844);
nand U7476 (N_7476,N_6417,N_6596);
nand U7477 (N_7477,N_6773,N_6677);
nor U7478 (N_7478,N_6079,N_6207);
nand U7479 (N_7479,N_6053,N_6294);
and U7480 (N_7480,N_6471,N_6724);
or U7481 (N_7481,N_6146,N_6228);
xor U7482 (N_7482,N_6639,N_6116);
xnor U7483 (N_7483,N_6433,N_6286);
nor U7484 (N_7484,N_6543,N_6125);
xnor U7485 (N_7485,N_6391,N_6581);
and U7486 (N_7486,N_6325,N_6703);
or U7487 (N_7487,N_6020,N_6808);
and U7488 (N_7488,N_6705,N_6552);
or U7489 (N_7489,N_6678,N_6075);
or U7490 (N_7490,N_6363,N_6963);
and U7491 (N_7491,N_6969,N_6455);
or U7492 (N_7492,N_6811,N_6977);
nand U7493 (N_7493,N_6832,N_6885);
nor U7494 (N_7494,N_6874,N_6824);
nand U7495 (N_7495,N_6572,N_6624);
and U7496 (N_7496,N_6975,N_6253);
and U7497 (N_7497,N_6023,N_6544);
nor U7498 (N_7498,N_6942,N_6282);
and U7499 (N_7499,N_6888,N_6198);
and U7500 (N_7500,N_6361,N_6415);
and U7501 (N_7501,N_6707,N_6640);
nand U7502 (N_7502,N_6996,N_6481);
nor U7503 (N_7503,N_6351,N_6502);
or U7504 (N_7504,N_6022,N_6874);
nand U7505 (N_7505,N_6351,N_6749);
xor U7506 (N_7506,N_6424,N_6657);
and U7507 (N_7507,N_6159,N_6830);
nand U7508 (N_7508,N_6428,N_6887);
nand U7509 (N_7509,N_6696,N_6657);
nor U7510 (N_7510,N_6858,N_6580);
nand U7511 (N_7511,N_6865,N_6932);
or U7512 (N_7512,N_6358,N_6123);
xor U7513 (N_7513,N_6690,N_6710);
nand U7514 (N_7514,N_6949,N_6372);
or U7515 (N_7515,N_6364,N_6147);
nor U7516 (N_7516,N_6096,N_6336);
or U7517 (N_7517,N_6243,N_6994);
and U7518 (N_7518,N_6904,N_6311);
xor U7519 (N_7519,N_6123,N_6762);
nor U7520 (N_7520,N_6693,N_6780);
and U7521 (N_7521,N_6266,N_6709);
or U7522 (N_7522,N_6646,N_6590);
and U7523 (N_7523,N_6061,N_6902);
and U7524 (N_7524,N_6290,N_6465);
nor U7525 (N_7525,N_6044,N_6665);
and U7526 (N_7526,N_6094,N_6250);
and U7527 (N_7527,N_6129,N_6185);
and U7528 (N_7528,N_6679,N_6308);
nor U7529 (N_7529,N_6760,N_6104);
xnor U7530 (N_7530,N_6162,N_6252);
and U7531 (N_7531,N_6379,N_6414);
xnor U7532 (N_7532,N_6065,N_6725);
and U7533 (N_7533,N_6805,N_6961);
and U7534 (N_7534,N_6068,N_6251);
nand U7535 (N_7535,N_6195,N_6328);
nor U7536 (N_7536,N_6435,N_6064);
nand U7537 (N_7537,N_6172,N_6991);
xor U7538 (N_7538,N_6117,N_6812);
or U7539 (N_7539,N_6723,N_6482);
and U7540 (N_7540,N_6469,N_6571);
nor U7541 (N_7541,N_6073,N_6547);
and U7542 (N_7542,N_6776,N_6841);
and U7543 (N_7543,N_6839,N_6042);
nand U7544 (N_7544,N_6699,N_6369);
nor U7545 (N_7545,N_6416,N_6752);
or U7546 (N_7546,N_6388,N_6959);
or U7547 (N_7547,N_6845,N_6796);
nand U7548 (N_7548,N_6276,N_6946);
or U7549 (N_7549,N_6760,N_6788);
nor U7550 (N_7550,N_6815,N_6781);
or U7551 (N_7551,N_6146,N_6865);
nor U7552 (N_7552,N_6226,N_6527);
xnor U7553 (N_7553,N_6256,N_6394);
nor U7554 (N_7554,N_6476,N_6478);
and U7555 (N_7555,N_6387,N_6198);
and U7556 (N_7556,N_6542,N_6106);
nor U7557 (N_7557,N_6521,N_6313);
and U7558 (N_7558,N_6587,N_6740);
nand U7559 (N_7559,N_6706,N_6070);
and U7560 (N_7560,N_6151,N_6252);
nand U7561 (N_7561,N_6178,N_6383);
nand U7562 (N_7562,N_6911,N_6058);
nand U7563 (N_7563,N_6627,N_6735);
nand U7564 (N_7564,N_6180,N_6746);
nor U7565 (N_7565,N_6805,N_6819);
or U7566 (N_7566,N_6439,N_6863);
or U7567 (N_7567,N_6703,N_6023);
xnor U7568 (N_7568,N_6857,N_6991);
and U7569 (N_7569,N_6790,N_6751);
nor U7570 (N_7570,N_6209,N_6118);
and U7571 (N_7571,N_6954,N_6141);
nand U7572 (N_7572,N_6844,N_6312);
and U7573 (N_7573,N_6166,N_6377);
nand U7574 (N_7574,N_6199,N_6437);
nand U7575 (N_7575,N_6191,N_6349);
and U7576 (N_7576,N_6136,N_6181);
nand U7577 (N_7577,N_6095,N_6922);
nor U7578 (N_7578,N_6874,N_6336);
xor U7579 (N_7579,N_6718,N_6120);
nor U7580 (N_7580,N_6882,N_6777);
nand U7581 (N_7581,N_6840,N_6754);
nor U7582 (N_7582,N_6056,N_6800);
nor U7583 (N_7583,N_6059,N_6283);
xor U7584 (N_7584,N_6468,N_6702);
and U7585 (N_7585,N_6903,N_6819);
nor U7586 (N_7586,N_6236,N_6238);
or U7587 (N_7587,N_6993,N_6784);
nor U7588 (N_7588,N_6933,N_6810);
nor U7589 (N_7589,N_6416,N_6640);
and U7590 (N_7590,N_6178,N_6680);
nand U7591 (N_7591,N_6181,N_6027);
nand U7592 (N_7592,N_6696,N_6042);
nor U7593 (N_7593,N_6814,N_6625);
nand U7594 (N_7594,N_6035,N_6927);
xor U7595 (N_7595,N_6668,N_6264);
nand U7596 (N_7596,N_6299,N_6281);
xor U7597 (N_7597,N_6440,N_6772);
or U7598 (N_7598,N_6883,N_6621);
and U7599 (N_7599,N_6791,N_6178);
nor U7600 (N_7600,N_6256,N_6578);
or U7601 (N_7601,N_6522,N_6889);
or U7602 (N_7602,N_6182,N_6315);
nor U7603 (N_7603,N_6388,N_6600);
and U7604 (N_7604,N_6221,N_6021);
xor U7605 (N_7605,N_6883,N_6416);
or U7606 (N_7606,N_6114,N_6357);
and U7607 (N_7607,N_6480,N_6692);
or U7608 (N_7608,N_6310,N_6807);
nand U7609 (N_7609,N_6233,N_6974);
xnor U7610 (N_7610,N_6324,N_6614);
nand U7611 (N_7611,N_6913,N_6743);
nand U7612 (N_7612,N_6116,N_6695);
nor U7613 (N_7613,N_6167,N_6126);
or U7614 (N_7614,N_6787,N_6228);
and U7615 (N_7615,N_6391,N_6717);
or U7616 (N_7616,N_6259,N_6858);
nor U7617 (N_7617,N_6428,N_6220);
or U7618 (N_7618,N_6081,N_6926);
or U7619 (N_7619,N_6904,N_6536);
nand U7620 (N_7620,N_6415,N_6618);
or U7621 (N_7621,N_6202,N_6249);
nand U7622 (N_7622,N_6046,N_6341);
nor U7623 (N_7623,N_6141,N_6824);
and U7624 (N_7624,N_6012,N_6625);
or U7625 (N_7625,N_6202,N_6534);
nand U7626 (N_7626,N_6435,N_6957);
nand U7627 (N_7627,N_6771,N_6452);
nor U7628 (N_7628,N_6120,N_6341);
nor U7629 (N_7629,N_6280,N_6563);
nor U7630 (N_7630,N_6732,N_6183);
nand U7631 (N_7631,N_6858,N_6630);
nand U7632 (N_7632,N_6536,N_6520);
or U7633 (N_7633,N_6590,N_6898);
or U7634 (N_7634,N_6875,N_6909);
nand U7635 (N_7635,N_6547,N_6465);
or U7636 (N_7636,N_6074,N_6743);
nand U7637 (N_7637,N_6878,N_6687);
and U7638 (N_7638,N_6196,N_6645);
and U7639 (N_7639,N_6684,N_6390);
or U7640 (N_7640,N_6817,N_6349);
and U7641 (N_7641,N_6087,N_6060);
nor U7642 (N_7642,N_6857,N_6426);
and U7643 (N_7643,N_6621,N_6499);
nor U7644 (N_7644,N_6971,N_6841);
xnor U7645 (N_7645,N_6166,N_6369);
or U7646 (N_7646,N_6124,N_6616);
nor U7647 (N_7647,N_6520,N_6729);
nor U7648 (N_7648,N_6666,N_6026);
and U7649 (N_7649,N_6905,N_6540);
and U7650 (N_7650,N_6161,N_6145);
nor U7651 (N_7651,N_6760,N_6766);
and U7652 (N_7652,N_6870,N_6867);
nor U7653 (N_7653,N_6460,N_6340);
nand U7654 (N_7654,N_6851,N_6371);
nand U7655 (N_7655,N_6317,N_6332);
and U7656 (N_7656,N_6475,N_6210);
nor U7657 (N_7657,N_6373,N_6564);
or U7658 (N_7658,N_6172,N_6224);
and U7659 (N_7659,N_6195,N_6060);
nor U7660 (N_7660,N_6341,N_6472);
nor U7661 (N_7661,N_6047,N_6964);
xor U7662 (N_7662,N_6398,N_6423);
nor U7663 (N_7663,N_6997,N_6076);
or U7664 (N_7664,N_6769,N_6890);
or U7665 (N_7665,N_6230,N_6956);
nor U7666 (N_7666,N_6531,N_6031);
and U7667 (N_7667,N_6993,N_6734);
or U7668 (N_7668,N_6567,N_6932);
xor U7669 (N_7669,N_6941,N_6753);
xor U7670 (N_7670,N_6123,N_6183);
and U7671 (N_7671,N_6814,N_6199);
and U7672 (N_7672,N_6781,N_6410);
and U7673 (N_7673,N_6811,N_6353);
and U7674 (N_7674,N_6909,N_6033);
nand U7675 (N_7675,N_6634,N_6584);
nand U7676 (N_7676,N_6518,N_6438);
nor U7677 (N_7677,N_6390,N_6649);
and U7678 (N_7678,N_6180,N_6005);
nand U7679 (N_7679,N_6709,N_6120);
or U7680 (N_7680,N_6769,N_6615);
or U7681 (N_7681,N_6463,N_6883);
nand U7682 (N_7682,N_6522,N_6695);
or U7683 (N_7683,N_6140,N_6924);
nand U7684 (N_7684,N_6640,N_6757);
and U7685 (N_7685,N_6656,N_6666);
nor U7686 (N_7686,N_6684,N_6746);
and U7687 (N_7687,N_6160,N_6986);
and U7688 (N_7688,N_6681,N_6001);
nor U7689 (N_7689,N_6594,N_6824);
and U7690 (N_7690,N_6380,N_6818);
and U7691 (N_7691,N_6210,N_6382);
nor U7692 (N_7692,N_6900,N_6459);
xnor U7693 (N_7693,N_6300,N_6120);
nand U7694 (N_7694,N_6388,N_6058);
nand U7695 (N_7695,N_6223,N_6645);
or U7696 (N_7696,N_6012,N_6807);
nand U7697 (N_7697,N_6289,N_6825);
or U7698 (N_7698,N_6905,N_6051);
nor U7699 (N_7699,N_6635,N_6340);
or U7700 (N_7700,N_6536,N_6807);
nor U7701 (N_7701,N_6339,N_6659);
nand U7702 (N_7702,N_6055,N_6232);
or U7703 (N_7703,N_6198,N_6200);
and U7704 (N_7704,N_6790,N_6926);
nor U7705 (N_7705,N_6847,N_6117);
nand U7706 (N_7706,N_6045,N_6061);
nor U7707 (N_7707,N_6267,N_6464);
or U7708 (N_7708,N_6667,N_6978);
nor U7709 (N_7709,N_6912,N_6761);
or U7710 (N_7710,N_6066,N_6723);
nor U7711 (N_7711,N_6209,N_6571);
or U7712 (N_7712,N_6651,N_6402);
xor U7713 (N_7713,N_6767,N_6658);
and U7714 (N_7714,N_6787,N_6621);
and U7715 (N_7715,N_6587,N_6286);
or U7716 (N_7716,N_6903,N_6938);
and U7717 (N_7717,N_6499,N_6596);
or U7718 (N_7718,N_6036,N_6363);
nor U7719 (N_7719,N_6866,N_6004);
nand U7720 (N_7720,N_6161,N_6737);
and U7721 (N_7721,N_6392,N_6254);
and U7722 (N_7722,N_6176,N_6002);
nor U7723 (N_7723,N_6778,N_6150);
or U7724 (N_7724,N_6862,N_6055);
nor U7725 (N_7725,N_6790,N_6729);
or U7726 (N_7726,N_6244,N_6064);
nand U7727 (N_7727,N_6746,N_6585);
and U7728 (N_7728,N_6518,N_6012);
nand U7729 (N_7729,N_6479,N_6598);
and U7730 (N_7730,N_6170,N_6580);
or U7731 (N_7731,N_6906,N_6992);
and U7732 (N_7732,N_6530,N_6680);
xor U7733 (N_7733,N_6275,N_6081);
nor U7734 (N_7734,N_6957,N_6098);
nor U7735 (N_7735,N_6462,N_6044);
and U7736 (N_7736,N_6151,N_6612);
and U7737 (N_7737,N_6557,N_6556);
nand U7738 (N_7738,N_6421,N_6438);
and U7739 (N_7739,N_6836,N_6463);
nand U7740 (N_7740,N_6859,N_6187);
xor U7741 (N_7741,N_6795,N_6589);
nand U7742 (N_7742,N_6028,N_6951);
nand U7743 (N_7743,N_6043,N_6729);
xnor U7744 (N_7744,N_6327,N_6299);
or U7745 (N_7745,N_6395,N_6985);
or U7746 (N_7746,N_6557,N_6684);
nand U7747 (N_7747,N_6195,N_6104);
and U7748 (N_7748,N_6408,N_6955);
nand U7749 (N_7749,N_6721,N_6561);
and U7750 (N_7750,N_6959,N_6224);
and U7751 (N_7751,N_6041,N_6837);
or U7752 (N_7752,N_6151,N_6431);
or U7753 (N_7753,N_6880,N_6973);
xor U7754 (N_7754,N_6306,N_6097);
nand U7755 (N_7755,N_6501,N_6667);
and U7756 (N_7756,N_6335,N_6947);
nor U7757 (N_7757,N_6114,N_6737);
and U7758 (N_7758,N_6101,N_6962);
or U7759 (N_7759,N_6234,N_6100);
or U7760 (N_7760,N_6961,N_6885);
nand U7761 (N_7761,N_6340,N_6662);
and U7762 (N_7762,N_6028,N_6236);
or U7763 (N_7763,N_6153,N_6354);
or U7764 (N_7764,N_6467,N_6979);
nand U7765 (N_7765,N_6590,N_6778);
and U7766 (N_7766,N_6014,N_6934);
nor U7767 (N_7767,N_6864,N_6560);
and U7768 (N_7768,N_6784,N_6357);
and U7769 (N_7769,N_6674,N_6104);
nor U7770 (N_7770,N_6451,N_6443);
nand U7771 (N_7771,N_6876,N_6919);
nand U7772 (N_7772,N_6432,N_6529);
and U7773 (N_7773,N_6671,N_6466);
and U7774 (N_7774,N_6758,N_6448);
nand U7775 (N_7775,N_6680,N_6737);
nand U7776 (N_7776,N_6888,N_6044);
or U7777 (N_7777,N_6764,N_6291);
nand U7778 (N_7778,N_6639,N_6881);
nor U7779 (N_7779,N_6507,N_6478);
nand U7780 (N_7780,N_6814,N_6849);
and U7781 (N_7781,N_6640,N_6506);
and U7782 (N_7782,N_6521,N_6145);
nand U7783 (N_7783,N_6225,N_6485);
or U7784 (N_7784,N_6406,N_6405);
nand U7785 (N_7785,N_6635,N_6764);
or U7786 (N_7786,N_6855,N_6944);
nand U7787 (N_7787,N_6379,N_6131);
nand U7788 (N_7788,N_6294,N_6507);
nor U7789 (N_7789,N_6174,N_6243);
nand U7790 (N_7790,N_6816,N_6571);
nand U7791 (N_7791,N_6400,N_6280);
or U7792 (N_7792,N_6081,N_6295);
nor U7793 (N_7793,N_6259,N_6495);
and U7794 (N_7794,N_6348,N_6472);
nor U7795 (N_7795,N_6318,N_6241);
nor U7796 (N_7796,N_6562,N_6556);
and U7797 (N_7797,N_6166,N_6632);
nand U7798 (N_7798,N_6614,N_6600);
xnor U7799 (N_7799,N_6416,N_6313);
xnor U7800 (N_7800,N_6414,N_6370);
nand U7801 (N_7801,N_6462,N_6296);
and U7802 (N_7802,N_6341,N_6254);
and U7803 (N_7803,N_6275,N_6239);
or U7804 (N_7804,N_6223,N_6778);
nor U7805 (N_7805,N_6215,N_6324);
nand U7806 (N_7806,N_6007,N_6621);
and U7807 (N_7807,N_6447,N_6011);
nor U7808 (N_7808,N_6587,N_6037);
or U7809 (N_7809,N_6315,N_6989);
and U7810 (N_7810,N_6516,N_6410);
and U7811 (N_7811,N_6623,N_6879);
nand U7812 (N_7812,N_6658,N_6948);
nor U7813 (N_7813,N_6551,N_6178);
nor U7814 (N_7814,N_6113,N_6766);
nor U7815 (N_7815,N_6503,N_6989);
and U7816 (N_7816,N_6047,N_6504);
nand U7817 (N_7817,N_6506,N_6920);
nor U7818 (N_7818,N_6033,N_6283);
nor U7819 (N_7819,N_6773,N_6318);
or U7820 (N_7820,N_6966,N_6667);
and U7821 (N_7821,N_6113,N_6284);
or U7822 (N_7822,N_6243,N_6784);
and U7823 (N_7823,N_6196,N_6424);
or U7824 (N_7824,N_6804,N_6108);
and U7825 (N_7825,N_6309,N_6012);
nand U7826 (N_7826,N_6937,N_6271);
xor U7827 (N_7827,N_6223,N_6203);
or U7828 (N_7828,N_6163,N_6446);
xor U7829 (N_7829,N_6436,N_6898);
and U7830 (N_7830,N_6150,N_6346);
nand U7831 (N_7831,N_6258,N_6815);
or U7832 (N_7832,N_6534,N_6881);
and U7833 (N_7833,N_6734,N_6194);
nor U7834 (N_7834,N_6484,N_6281);
nand U7835 (N_7835,N_6647,N_6631);
nand U7836 (N_7836,N_6265,N_6091);
and U7837 (N_7837,N_6780,N_6171);
or U7838 (N_7838,N_6949,N_6802);
xor U7839 (N_7839,N_6216,N_6094);
nor U7840 (N_7840,N_6234,N_6315);
and U7841 (N_7841,N_6963,N_6283);
nor U7842 (N_7842,N_6490,N_6032);
nand U7843 (N_7843,N_6421,N_6243);
xor U7844 (N_7844,N_6071,N_6872);
and U7845 (N_7845,N_6771,N_6018);
or U7846 (N_7846,N_6849,N_6999);
and U7847 (N_7847,N_6132,N_6947);
nor U7848 (N_7848,N_6572,N_6638);
nor U7849 (N_7849,N_6336,N_6497);
or U7850 (N_7850,N_6396,N_6071);
and U7851 (N_7851,N_6788,N_6809);
xnor U7852 (N_7852,N_6770,N_6118);
or U7853 (N_7853,N_6960,N_6773);
xnor U7854 (N_7854,N_6028,N_6079);
and U7855 (N_7855,N_6937,N_6115);
and U7856 (N_7856,N_6303,N_6220);
nor U7857 (N_7857,N_6971,N_6792);
and U7858 (N_7858,N_6818,N_6666);
and U7859 (N_7859,N_6742,N_6779);
and U7860 (N_7860,N_6389,N_6477);
nor U7861 (N_7861,N_6814,N_6091);
or U7862 (N_7862,N_6428,N_6545);
and U7863 (N_7863,N_6066,N_6401);
and U7864 (N_7864,N_6409,N_6219);
and U7865 (N_7865,N_6794,N_6896);
or U7866 (N_7866,N_6905,N_6396);
nand U7867 (N_7867,N_6440,N_6694);
and U7868 (N_7868,N_6470,N_6414);
nand U7869 (N_7869,N_6326,N_6049);
or U7870 (N_7870,N_6837,N_6029);
nor U7871 (N_7871,N_6663,N_6598);
nand U7872 (N_7872,N_6319,N_6179);
or U7873 (N_7873,N_6206,N_6818);
nand U7874 (N_7874,N_6334,N_6396);
xor U7875 (N_7875,N_6282,N_6964);
or U7876 (N_7876,N_6479,N_6106);
nor U7877 (N_7877,N_6650,N_6597);
and U7878 (N_7878,N_6038,N_6892);
or U7879 (N_7879,N_6847,N_6312);
and U7880 (N_7880,N_6993,N_6143);
or U7881 (N_7881,N_6946,N_6361);
nand U7882 (N_7882,N_6679,N_6685);
and U7883 (N_7883,N_6749,N_6785);
and U7884 (N_7884,N_6887,N_6089);
nor U7885 (N_7885,N_6493,N_6614);
nand U7886 (N_7886,N_6924,N_6222);
and U7887 (N_7887,N_6681,N_6939);
nand U7888 (N_7888,N_6136,N_6116);
nor U7889 (N_7889,N_6769,N_6968);
nor U7890 (N_7890,N_6878,N_6223);
nor U7891 (N_7891,N_6421,N_6997);
or U7892 (N_7892,N_6792,N_6464);
nand U7893 (N_7893,N_6817,N_6072);
or U7894 (N_7894,N_6212,N_6437);
xor U7895 (N_7895,N_6565,N_6969);
and U7896 (N_7896,N_6799,N_6022);
nand U7897 (N_7897,N_6343,N_6970);
nand U7898 (N_7898,N_6532,N_6654);
nor U7899 (N_7899,N_6731,N_6224);
or U7900 (N_7900,N_6915,N_6125);
nand U7901 (N_7901,N_6824,N_6981);
or U7902 (N_7902,N_6598,N_6148);
nor U7903 (N_7903,N_6424,N_6525);
and U7904 (N_7904,N_6364,N_6693);
and U7905 (N_7905,N_6842,N_6746);
and U7906 (N_7906,N_6128,N_6635);
or U7907 (N_7907,N_6691,N_6439);
and U7908 (N_7908,N_6840,N_6338);
xor U7909 (N_7909,N_6052,N_6626);
nor U7910 (N_7910,N_6707,N_6200);
xnor U7911 (N_7911,N_6203,N_6430);
and U7912 (N_7912,N_6669,N_6922);
and U7913 (N_7913,N_6615,N_6572);
and U7914 (N_7914,N_6163,N_6086);
and U7915 (N_7915,N_6081,N_6059);
xnor U7916 (N_7916,N_6622,N_6440);
and U7917 (N_7917,N_6300,N_6093);
nor U7918 (N_7918,N_6776,N_6834);
or U7919 (N_7919,N_6382,N_6718);
nor U7920 (N_7920,N_6953,N_6156);
nand U7921 (N_7921,N_6662,N_6658);
nor U7922 (N_7922,N_6482,N_6281);
xor U7923 (N_7923,N_6197,N_6506);
nor U7924 (N_7924,N_6143,N_6987);
nand U7925 (N_7925,N_6694,N_6822);
or U7926 (N_7926,N_6480,N_6922);
and U7927 (N_7927,N_6759,N_6376);
and U7928 (N_7928,N_6403,N_6965);
xor U7929 (N_7929,N_6128,N_6682);
xor U7930 (N_7930,N_6689,N_6758);
xnor U7931 (N_7931,N_6969,N_6647);
and U7932 (N_7932,N_6000,N_6046);
nand U7933 (N_7933,N_6025,N_6532);
or U7934 (N_7934,N_6100,N_6813);
or U7935 (N_7935,N_6499,N_6075);
and U7936 (N_7936,N_6797,N_6544);
nor U7937 (N_7937,N_6264,N_6832);
nor U7938 (N_7938,N_6019,N_6704);
nand U7939 (N_7939,N_6415,N_6929);
or U7940 (N_7940,N_6298,N_6874);
or U7941 (N_7941,N_6677,N_6508);
nand U7942 (N_7942,N_6367,N_6272);
nor U7943 (N_7943,N_6862,N_6359);
or U7944 (N_7944,N_6407,N_6859);
xor U7945 (N_7945,N_6871,N_6708);
nor U7946 (N_7946,N_6475,N_6143);
and U7947 (N_7947,N_6160,N_6554);
nor U7948 (N_7948,N_6447,N_6634);
nor U7949 (N_7949,N_6896,N_6429);
nor U7950 (N_7950,N_6972,N_6041);
xnor U7951 (N_7951,N_6310,N_6587);
and U7952 (N_7952,N_6744,N_6831);
and U7953 (N_7953,N_6190,N_6999);
and U7954 (N_7954,N_6232,N_6522);
and U7955 (N_7955,N_6030,N_6939);
nor U7956 (N_7956,N_6728,N_6425);
and U7957 (N_7957,N_6211,N_6679);
nand U7958 (N_7958,N_6952,N_6461);
nor U7959 (N_7959,N_6030,N_6011);
or U7960 (N_7960,N_6099,N_6670);
or U7961 (N_7961,N_6879,N_6777);
and U7962 (N_7962,N_6856,N_6639);
or U7963 (N_7963,N_6431,N_6103);
or U7964 (N_7964,N_6362,N_6335);
nor U7965 (N_7965,N_6694,N_6688);
nand U7966 (N_7966,N_6176,N_6455);
nand U7967 (N_7967,N_6985,N_6225);
nor U7968 (N_7968,N_6721,N_6403);
nand U7969 (N_7969,N_6900,N_6162);
and U7970 (N_7970,N_6019,N_6498);
or U7971 (N_7971,N_6607,N_6441);
nor U7972 (N_7972,N_6556,N_6602);
nor U7973 (N_7973,N_6325,N_6898);
and U7974 (N_7974,N_6877,N_6882);
nor U7975 (N_7975,N_6834,N_6991);
nor U7976 (N_7976,N_6196,N_6662);
or U7977 (N_7977,N_6733,N_6375);
or U7978 (N_7978,N_6904,N_6911);
and U7979 (N_7979,N_6276,N_6171);
and U7980 (N_7980,N_6341,N_6376);
nor U7981 (N_7981,N_6795,N_6914);
or U7982 (N_7982,N_6803,N_6317);
and U7983 (N_7983,N_6136,N_6019);
nand U7984 (N_7984,N_6315,N_6920);
nand U7985 (N_7985,N_6227,N_6403);
nor U7986 (N_7986,N_6204,N_6510);
and U7987 (N_7987,N_6565,N_6613);
nand U7988 (N_7988,N_6674,N_6099);
xor U7989 (N_7989,N_6212,N_6382);
and U7990 (N_7990,N_6894,N_6588);
xnor U7991 (N_7991,N_6422,N_6561);
nand U7992 (N_7992,N_6546,N_6155);
and U7993 (N_7993,N_6599,N_6783);
xor U7994 (N_7994,N_6421,N_6483);
and U7995 (N_7995,N_6982,N_6206);
and U7996 (N_7996,N_6251,N_6362);
nand U7997 (N_7997,N_6629,N_6268);
nor U7998 (N_7998,N_6402,N_6254);
nand U7999 (N_7999,N_6358,N_6432);
or U8000 (N_8000,N_7309,N_7004);
or U8001 (N_8001,N_7364,N_7612);
nand U8002 (N_8002,N_7100,N_7091);
nor U8003 (N_8003,N_7257,N_7930);
and U8004 (N_8004,N_7263,N_7692);
or U8005 (N_8005,N_7881,N_7926);
nor U8006 (N_8006,N_7474,N_7492);
or U8007 (N_8007,N_7621,N_7062);
nand U8008 (N_8008,N_7082,N_7054);
xor U8009 (N_8009,N_7316,N_7246);
and U8010 (N_8010,N_7842,N_7835);
nand U8011 (N_8011,N_7590,N_7884);
nor U8012 (N_8012,N_7851,N_7404);
nand U8013 (N_8013,N_7837,N_7941);
nor U8014 (N_8014,N_7391,N_7682);
and U8015 (N_8015,N_7102,N_7997);
and U8016 (N_8016,N_7751,N_7301);
and U8017 (N_8017,N_7581,N_7708);
and U8018 (N_8018,N_7186,N_7457);
and U8019 (N_8019,N_7768,N_7323);
or U8020 (N_8020,N_7470,N_7182);
nor U8021 (N_8021,N_7256,N_7018);
nor U8022 (N_8022,N_7880,N_7329);
or U8023 (N_8023,N_7295,N_7615);
nor U8024 (N_8024,N_7414,N_7703);
or U8025 (N_8025,N_7764,N_7347);
nand U8026 (N_8026,N_7467,N_7523);
nor U8027 (N_8027,N_7962,N_7187);
nor U8028 (N_8028,N_7285,N_7326);
nor U8029 (N_8029,N_7743,N_7800);
nand U8030 (N_8030,N_7732,N_7903);
nand U8031 (N_8031,N_7971,N_7373);
nor U8032 (N_8032,N_7169,N_7225);
nor U8033 (N_8033,N_7524,N_7741);
and U8034 (N_8034,N_7509,N_7180);
nand U8035 (N_8035,N_7385,N_7072);
or U8036 (N_8036,N_7589,N_7033);
nor U8037 (N_8037,N_7411,N_7689);
nand U8038 (N_8038,N_7977,N_7325);
nand U8039 (N_8039,N_7924,N_7558);
or U8040 (N_8040,N_7773,N_7296);
and U8041 (N_8041,N_7633,N_7080);
nand U8042 (N_8042,N_7655,N_7731);
nor U8043 (N_8043,N_7950,N_7912);
nor U8044 (N_8044,N_7852,N_7630);
nand U8045 (N_8045,N_7552,N_7118);
nor U8046 (N_8046,N_7405,N_7964);
nand U8047 (N_8047,N_7146,N_7090);
or U8048 (N_8048,N_7324,N_7674);
nand U8049 (N_8049,N_7554,N_7846);
nor U8050 (N_8050,N_7020,N_7645);
xnor U8051 (N_8051,N_7602,N_7679);
or U8052 (N_8052,N_7663,N_7916);
nand U8053 (N_8053,N_7588,N_7879);
nand U8054 (N_8054,N_7642,N_7580);
and U8055 (N_8055,N_7436,N_7586);
and U8056 (N_8056,N_7793,N_7268);
nor U8057 (N_8057,N_7440,N_7421);
and U8058 (N_8058,N_7332,N_7306);
nand U8059 (N_8059,N_7643,N_7745);
nor U8060 (N_8060,N_7279,N_7949);
nor U8061 (N_8061,N_7623,N_7855);
nand U8062 (N_8062,N_7006,N_7401);
nor U8063 (N_8063,N_7841,N_7055);
or U8064 (N_8064,N_7810,N_7951);
or U8065 (N_8065,N_7752,N_7357);
nor U8066 (N_8066,N_7957,N_7857);
and U8067 (N_8067,N_7668,N_7025);
or U8068 (N_8068,N_7925,N_7906);
nand U8069 (N_8069,N_7736,N_7089);
nor U8070 (N_8070,N_7008,N_7378);
nand U8071 (N_8071,N_7922,N_7486);
nand U8072 (N_8072,N_7678,N_7733);
and U8073 (N_8073,N_7226,N_7730);
and U8074 (N_8074,N_7988,N_7711);
and U8075 (N_8075,N_7178,N_7734);
xor U8076 (N_8076,N_7009,N_7371);
nand U8077 (N_8077,N_7656,N_7041);
and U8078 (N_8078,N_7005,N_7681);
nor U8079 (N_8079,N_7893,N_7998);
or U8080 (N_8080,N_7699,N_7471);
nand U8081 (N_8081,N_7044,N_7836);
and U8082 (N_8082,N_7850,N_7048);
and U8083 (N_8083,N_7431,N_7874);
and U8084 (N_8084,N_7389,N_7978);
xor U8085 (N_8085,N_7770,N_7298);
xnor U8086 (N_8086,N_7153,N_7042);
nand U8087 (N_8087,N_7076,N_7993);
nor U8088 (N_8088,N_7046,N_7334);
or U8089 (N_8089,N_7662,N_7777);
nand U8090 (N_8090,N_7819,N_7218);
nand U8091 (N_8091,N_7567,N_7490);
nor U8092 (N_8092,N_7706,N_7454);
and U8093 (N_8093,N_7255,N_7318);
and U8094 (N_8094,N_7130,N_7904);
nand U8095 (N_8095,N_7863,N_7198);
nor U8096 (N_8096,N_7902,N_7578);
or U8097 (N_8097,N_7849,N_7231);
nor U8098 (N_8098,N_7463,N_7038);
nor U8099 (N_8099,N_7680,N_7189);
and U8100 (N_8100,N_7227,N_7070);
nor U8101 (N_8101,N_7654,N_7002);
or U8102 (N_8102,N_7936,N_7345);
nor U8103 (N_8103,N_7876,N_7501);
and U8104 (N_8104,N_7536,N_7363);
nor U8105 (N_8105,N_7196,N_7079);
nand U8106 (N_8106,N_7016,N_7212);
or U8107 (N_8107,N_7735,N_7195);
or U8108 (N_8108,N_7336,N_7388);
or U8109 (N_8109,N_7183,N_7720);
and U8110 (N_8110,N_7300,N_7099);
xnor U8111 (N_8111,N_7783,N_7223);
or U8112 (N_8112,N_7286,N_7366);
nor U8113 (N_8113,N_7015,N_7619);
and U8114 (N_8114,N_7119,N_7980);
and U8115 (N_8115,N_7175,N_7353);
and U8116 (N_8116,N_7972,N_7249);
nor U8117 (N_8117,N_7131,N_7392);
nor U8118 (N_8118,N_7505,N_7785);
nand U8119 (N_8119,N_7503,N_7460);
nand U8120 (N_8120,N_7224,N_7968);
nand U8121 (N_8121,N_7928,N_7817);
and U8122 (N_8122,N_7381,N_7862);
or U8123 (N_8123,N_7833,N_7894);
or U8124 (N_8124,N_7540,N_7164);
and U8125 (N_8125,N_7715,N_7379);
or U8126 (N_8126,N_7151,N_7024);
or U8127 (N_8127,N_7278,N_7466);
nand U8128 (N_8128,N_7609,N_7696);
or U8129 (N_8129,N_7487,N_7160);
and U8130 (N_8130,N_7010,N_7648);
nor U8131 (N_8131,N_7050,N_7291);
xnor U8132 (N_8132,N_7425,N_7308);
nor U8133 (N_8133,N_7613,N_7780);
and U8134 (N_8134,N_7631,N_7843);
nor U8135 (N_8135,N_7337,N_7999);
and U8136 (N_8136,N_7142,N_7267);
nor U8137 (N_8137,N_7791,N_7254);
nor U8138 (N_8138,N_7823,N_7493);
or U8139 (N_8139,N_7485,N_7701);
nor U8140 (N_8140,N_7600,N_7116);
nor U8141 (N_8141,N_7495,N_7756);
nor U8142 (N_8142,N_7352,N_7313);
nor U8143 (N_8143,N_7779,N_7684);
xnor U8144 (N_8144,N_7700,N_7955);
xor U8145 (N_8145,N_7737,N_7694);
nand U8146 (N_8146,N_7331,N_7284);
nor U8147 (N_8147,N_7349,N_7420);
or U8148 (N_8148,N_7830,N_7141);
nor U8149 (N_8149,N_7302,N_7832);
nand U8150 (N_8150,N_7104,N_7443);
or U8151 (N_8151,N_7543,N_7624);
or U8152 (N_8152,N_7801,N_7799);
and U8153 (N_8153,N_7891,N_7686);
nor U8154 (N_8154,N_7270,N_7551);
nand U8155 (N_8155,N_7166,N_7013);
and U8156 (N_8156,N_7790,N_7568);
nand U8157 (N_8157,N_7387,N_7125);
nor U8158 (N_8158,N_7652,N_7803);
nor U8159 (N_8159,N_7190,N_7521);
nand U8160 (N_8160,N_7864,N_7776);
or U8161 (N_8161,N_7539,N_7909);
and U8162 (N_8162,N_7872,N_7370);
xor U8163 (N_8163,N_7671,N_7611);
xnor U8164 (N_8164,N_7135,N_7165);
and U8165 (N_8165,N_7570,N_7188);
nand U8166 (N_8166,N_7593,N_7123);
nor U8167 (N_8167,N_7144,N_7320);
or U8168 (N_8168,N_7563,N_7986);
xor U8169 (N_8169,N_7264,N_7883);
and U8170 (N_8170,N_7746,N_7172);
nand U8171 (N_8171,N_7210,N_7533);
or U8172 (N_8172,N_7214,N_7825);
nand U8173 (N_8173,N_7106,N_7606);
nand U8174 (N_8174,N_7544,N_7281);
nor U8175 (N_8175,N_7519,N_7510);
or U8176 (N_8176,N_7161,N_7209);
nand U8177 (N_8177,N_7342,N_7506);
and U8178 (N_8178,N_7572,N_7078);
nand U8179 (N_8179,N_7895,N_7838);
xor U8180 (N_8180,N_7139,N_7649);
and U8181 (N_8181,N_7233,N_7339);
nor U8182 (N_8182,N_7987,N_7494);
nor U8183 (N_8183,N_7721,N_7150);
nor U8184 (N_8184,N_7896,N_7758);
nand U8185 (N_8185,N_7028,N_7739);
or U8186 (N_8186,N_7573,N_7557);
xor U8187 (N_8187,N_7488,N_7087);
nor U8188 (N_8188,N_7637,N_7806);
or U8189 (N_8189,N_7661,N_7243);
or U8190 (N_8190,N_7512,N_7133);
nand U8191 (N_8191,N_7386,N_7629);
nor U8192 (N_8192,N_7238,N_7356);
nor U8193 (N_8193,N_7556,N_7582);
or U8194 (N_8194,N_7763,N_7945);
and U8195 (N_8195,N_7887,N_7577);
nor U8196 (N_8196,N_7695,N_7113);
nor U8197 (N_8197,N_7333,N_7958);
and U8198 (N_8198,N_7075,N_7083);
nand U8199 (N_8199,N_7650,N_7412);
or U8200 (N_8200,N_7596,N_7129);
nor U8201 (N_8201,N_7128,N_7375);
or U8202 (N_8202,N_7597,N_7697);
nor U8203 (N_8203,N_7618,N_7625);
xnor U8204 (N_8204,N_7712,N_7240);
and U8205 (N_8205,N_7416,N_7134);
or U8206 (N_8206,N_7826,N_7380);
or U8207 (N_8207,N_7867,N_7458);
xor U8208 (N_8208,N_7344,N_7241);
or U8209 (N_8209,N_7060,N_7418);
or U8210 (N_8210,N_7262,N_7340);
nor U8211 (N_8211,N_7795,N_7515);
and U8212 (N_8212,N_7750,N_7628);
nor U8213 (N_8213,N_7946,N_7766);
and U8214 (N_8214,N_7289,N_7651);
xor U8215 (N_8215,N_7448,N_7937);
nor U8216 (N_8216,N_7927,N_7096);
nand U8217 (N_8217,N_7396,N_7744);
or U8218 (N_8218,N_7499,N_7472);
or U8219 (N_8219,N_7067,N_7234);
and U8220 (N_8220,N_7818,N_7383);
or U8221 (N_8221,N_7415,N_7000);
and U8222 (N_8222,N_7056,N_7029);
and U8223 (N_8223,N_7136,N_7673);
or U8224 (N_8224,N_7138,N_7394);
nand U8225 (N_8225,N_7157,N_7878);
and U8226 (N_8226,N_7839,N_7959);
nand U8227 (N_8227,N_7579,N_7030);
or U8228 (N_8228,N_7147,N_7868);
nor U8229 (N_8229,N_7346,N_7402);
and U8230 (N_8230,N_7395,N_7753);
and U8231 (N_8231,N_7538,N_7963);
nand U8232 (N_8232,N_7669,N_7504);
or U8233 (N_8233,N_7702,N_7114);
or U8234 (N_8234,N_7564,N_7107);
xnor U8235 (N_8235,N_7798,N_7635);
xor U8236 (N_8236,N_7479,N_7239);
xor U8237 (N_8237,N_7315,N_7176);
nor U8238 (N_8238,N_7489,N_7307);
and U8239 (N_8239,N_7498,N_7944);
and U8240 (N_8240,N_7451,N_7714);
or U8241 (N_8241,N_7426,N_7638);
xnor U8242 (N_8242,N_7769,N_7181);
nand U8243 (N_8243,N_7815,N_7261);
and U8244 (N_8244,N_7283,N_7321);
or U8245 (N_8245,N_7250,N_7541);
xor U8246 (N_8246,N_7858,N_7974);
nor U8247 (N_8247,N_7667,N_7603);
nor U8248 (N_8248,N_7634,N_7253);
and U8249 (N_8249,N_7031,N_7954);
and U8250 (N_8250,N_7742,N_7917);
xor U8251 (N_8251,N_7410,N_7870);
xor U8252 (N_8252,N_7991,N_7774);
or U8253 (N_8253,N_7216,N_7417);
nand U8254 (N_8254,N_7975,N_7052);
or U8255 (N_8255,N_7456,N_7011);
nor U8256 (N_8256,N_7036,N_7861);
and U8257 (N_8257,N_7772,N_7057);
nor U8258 (N_8258,N_7814,N_7549);
or U8259 (N_8259,N_7531,N_7996);
or U8260 (N_8260,N_7704,N_7093);
nand U8261 (N_8261,N_7423,N_7914);
nor U8262 (N_8262,N_7368,N_7088);
and U8263 (N_8263,N_7901,N_7361);
xor U8264 (N_8264,N_7317,N_7095);
nand U8265 (N_8265,N_7132,N_7259);
nor U8266 (N_8266,N_7413,N_7705);
or U8267 (N_8267,N_7707,N_7351);
xnor U8268 (N_8268,N_7502,N_7251);
nor U8269 (N_8269,N_7845,N_7709);
nand U8270 (N_8270,N_7314,N_7156);
or U8271 (N_8271,N_7081,N_7856);
or U8272 (N_8272,N_7873,N_7328);
and U8273 (N_8273,N_7976,N_7021);
nor U8274 (N_8274,N_7518,N_7127);
xnor U8275 (N_8275,N_7910,N_7084);
or U8276 (N_8276,N_7913,N_7529);
and U8277 (N_8277,N_7358,N_7517);
and U8278 (N_8278,N_7585,N_7532);
nor U8279 (N_8279,N_7433,N_7061);
nor U8280 (N_8280,N_7108,N_7280);
nand U8281 (N_8281,N_7397,N_7235);
nor U8282 (N_8282,N_7059,N_7882);
xor U8283 (N_8283,N_7859,N_7807);
and U8284 (N_8284,N_7237,N_7527);
nand U8285 (N_8285,N_7110,N_7897);
nor U8286 (N_8286,N_7754,N_7449);
nor U8287 (N_8287,N_7691,N_7848);
xor U8288 (N_8288,N_7865,N_7407);
nand U8289 (N_8289,N_7229,N_7595);
nand U8290 (N_8290,N_7507,N_7014);
nand U8291 (N_8291,N_7583,N_7120);
and U8292 (N_8292,N_7001,N_7875);
nand U8293 (N_8293,N_7561,N_7967);
nand U8294 (N_8294,N_7724,N_7468);
and U8295 (N_8295,N_7022,N_7117);
and U8296 (N_8296,N_7690,N_7162);
nor U8297 (N_8297,N_7242,N_7462);
nand U8298 (N_8298,N_7382,N_7427);
nor U8299 (N_8299,N_7399,N_7007);
nand U8300 (N_8300,N_7647,N_7698);
or U8301 (N_8301,N_7207,N_7159);
nand U8302 (N_8302,N_7670,N_7824);
and U8303 (N_8303,N_7604,N_7481);
xnor U8304 (N_8304,N_7534,N_7408);
xor U8305 (N_8305,N_7137,N_7171);
and U8306 (N_8306,N_7074,N_7660);
or U8307 (N_8307,N_7476,N_7728);
or U8308 (N_8308,N_7071,N_7933);
and U8309 (N_8309,N_7947,N_7525);
nand U8310 (N_8310,N_7453,N_7455);
and U8311 (N_8311,N_7767,N_7553);
xnor U8312 (N_8312,N_7445,N_7437);
and U8313 (N_8313,N_7866,N_7086);
or U8314 (N_8314,N_7961,N_7956);
or U8315 (N_8315,N_7204,N_7860);
and U8316 (N_8316,N_7441,N_7693);
xnor U8317 (N_8317,N_7429,N_7886);
nand U8318 (N_8318,N_7778,N_7526);
nor U8319 (N_8319,N_7215,N_7994);
nor U8320 (N_8320,N_7584,N_7571);
nand U8321 (N_8321,N_7012,N_7938);
nand U8322 (N_8322,N_7464,N_7748);
nand U8323 (N_8323,N_7040,N_7688);
nand U8324 (N_8324,N_7636,N_7177);
or U8325 (N_8325,N_7816,N_7522);
or U8326 (N_8326,N_7710,N_7676);
xnor U8327 (N_8327,N_7155,N_7892);
and U8328 (N_8328,N_7304,N_7219);
nand U8329 (N_8329,N_7452,N_7335);
and U8330 (N_8330,N_7197,N_7788);
nor U8331 (N_8331,N_7664,N_7723);
xnor U8332 (N_8332,N_7354,N_7569);
or U8333 (N_8333,N_7066,N_7992);
xor U8334 (N_8334,N_7065,N_7666);
nor U8335 (N_8335,N_7199,N_7252);
xnor U8336 (N_8336,N_7247,N_7899);
nor U8337 (N_8337,N_7970,N_7948);
and U8338 (N_8338,N_7222,N_7771);
nor U8339 (N_8339,N_7469,N_7154);
nand U8340 (N_8340,N_7528,N_7786);
and U8341 (N_8341,N_7173,N_7943);
and U8342 (N_8342,N_7068,N_7034);
nand U8343 (N_8343,N_7966,N_7657);
nand U8344 (N_8344,N_7989,N_7276);
or U8345 (N_8345,N_7592,N_7713);
nor U8346 (N_8346,N_7442,N_7167);
and U8347 (N_8347,N_7822,N_7101);
nor U8348 (N_8348,N_7761,N_7475);
nand U8349 (N_8349,N_7828,N_7905);
and U8350 (N_8350,N_7362,N_7174);
or U8351 (N_8351,N_7367,N_7729);
nor U8352 (N_8352,N_7400,N_7047);
or U8353 (N_8353,N_7871,N_7221);
or U8354 (N_8354,N_7685,N_7665);
xor U8355 (N_8355,N_7935,N_7312);
and U8356 (N_8356,N_7658,N_7508);
or U8357 (N_8357,N_7726,N_7853);
and U8358 (N_8358,N_7145,N_7069);
xor U8359 (N_8359,N_7244,N_7717);
or U8360 (N_8360,N_7434,N_7112);
nand U8361 (N_8361,N_7939,N_7447);
nand U8362 (N_8362,N_7184,N_7794);
or U8363 (N_8363,N_7749,N_7537);
and U8364 (N_8364,N_7045,N_7311);
or U8365 (N_8365,N_7804,N_7043);
nor U8366 (N_8366,N_7430,N_7480);
nand U8367 (N_8367,N_7152,N_7105);
xor U8368 (N_8368,N_7126,N_7360);
nand U8369 (N_8369,N_7158,N_7220);
nor U8370 (N_8370,N_7796,N_7432);
and U8371 (N_8371,N_7566,N_7587);
nor U8372 (N_8372,N_7802,N_7271);
or U8373 (N_8373,N_7406,N_7511);
or U8374 (N_8374,N_7542,N_7960);
and U8375 (N_8375,N_7759,N_7051);
nor U8376 (N_8376,N_7201,N_7419);
and U8377 (N_8377,N_7918,N_7622);
or U8378 (N_8378,N_7439,N_7393);
xor U8379 (N_8379,N_7821,N_7844);
and U8380 (N_8380,N_7103,N_7122);
and U8381 (N_8381,N_7607,N_7919);
nand U8382 (N_8382,N_7027,N_7109);
nand U8383 (N_8383,N_7359,N_7591);
nor U8384 (N_8384,N_7716,N_7185);
or U8385 (N_8385,N_7626,N_7111);
nand U8386 (N_8386,N_7598,N_7760);
and U8387 (N_8387,N_7438,N_7322);
nor U8388 (N_8388,N_7725,N_7934);
nand U8389 (N_8389,N_7288,N_7273);
and U8390 (N_8390,N_7341,N_7124);
nand U8391 (N_8391,N_7847,N_7203);
nor U8392 (N_8392,N_7535,N_7374);
nand U8393 (N_8393,N_7547,N_7459);
nor U8394 (N_8394,N_7245,N_7921);
xor U8395 (N_8395,N_7200,N_7484);
nand U8396 (N_8396,N_7377,N_7202);
nand U8397 (N_8397,N_7548,N_7019);
xor U8398 (N_8398,N_7266,N_7565);
nand U8399 (N_8399,N_7514,N_7064);
nand U8400 (N_8400,N_7740,N_7940);
and U8401 (N_8401,N_7639,N_7984);
or U8402 (N_8402,N_7319,N_7403);
nor U8403 (N_8403,N_7272,N_7775);
nor U8404 (N_8404,N_7275,N_7915);
and U8405 (N_8405,N_7755,N_7115);
or U8406 (N_8406,N_7026,N_7888);
nand U8407 (N_8407,N_7605,N_7911);
nand U8408 (N_8408,N_7170,N_7576);
nor U8409 (N_8409,N_7907,N_7632);
nor U8410 (N_8410,N_7230,N_7877);
xnor U8411 (N_8411,N_7931,N_7781);
nand U8412 (N_8412,N_7620,N_7343);
nor U8413 (N_8413,N_7477,N_7831);
or U8414 (N_8414,N_7599,N_7898);
nand U8415 (N_8415,N_7820,N_7981);
nor U8416 (N_8416,N_7675,N_7149);
nor U8417 (N_8417,N_7274,N_7829);
nor U8418 (N_8418,N_7265,N_7369);
or U8419 (N_8419,N_7092,N_7348);
or U8420 (N_8420,N_7834,N_7969);
and U8421 (N_8421,N_7640,N_7236);
or U8422 (N_8422,N_7809,N_7208);
nor U8423 (N_8423,N_7390,N_7789);
nor U8424 (N_8424,N_7757,N_7646);
and U8425 (N_8425,N_7797,N_7398);
and U8426 (N_8426,N_7500,N_7516);
nand U8427 (N_8427,N_7953,N_7659);
nor U8428 (N_8428,N_7805,N_7677);
or U8429 (N_8429,N_7653,N_7747);
and U8430 (N_8430,N_7428,N_7073);
nor U8431 (N_8431,N_7929,N_7520);
and U8432 (N_8432,N_7491,N_7032);
and U8433 (N_8433,N_7497,N_7424);
or U8434 (N_8434,N_7465,N_7496);
or U8435 (N_8435,N_7277,N_7384);
or U8436 (N_8436,N_7297,N_7035);
nand U8437 (N_8437,N_7942,N_7217);
or U8438 (N_8438,N_7601,N_7952);
nand U8439 (N_8439,N_7854,N_7473);
xnor U8440 (N_8440,N_7973,N_7545);
xor U8441 (N_8441,N_7719,N_7784);
and U8442 (N_8442,N_7827,N_7258);
and U8443 (N_8443,N_7722,N_7094);
nand U8444 (N_8444,N_7097,N_7979);
nand U8445 (N_8445,N_7148,N_7017);
nand U8446 (N_8446,N_7299,N_7513);
nor U8447 (N_8447,N_7191,N_7098);
xor U8448 (N_8448,N_7327,N_7478);
and U8449 (N_8449,N_7672,N_7575);
or U8450 (N_8450,N_7330,N_7687);
nor U8451 (N_8451,N_7192,N_7530);
nor U8452 (N_8452,N_7762,N_7574);
nand U8453 (N_8453,N_7811,N_7211);
nand U8454 (N_8454,N_7985,N_7409);
xnor U8455 (N_8455,N_7765,N_7206);
and U8456 (N_8456,N_7450,N_7983);
nor U8457 (N_8457,N_7037,N_7248);
or U8458 (N_8458,N_7179,N_7435);
nor U8459 (N_8459,N_7965,N_7058);
nand U8460 (N_8460,N_7163,N_7228);
and U8461 (N_8461,N_7049,N_7355);
and U8462 (N_8462,N_7085,N_7287);
and U8463 (N_8463,N_7121,N_7644);
and U8464 (N_8464,N_7023,N_7140);
or U8465 (N_8465,N_7594,N_7260);
xnor U8466 (N_8466,N_7727,N_7444);
nand U8467 (N_8467,N_7290,N_7338);
or U8468 (N_8468,N_7294,N_7303);
or U8469 (N_8469,N_7990,N_7482);
or U8470 (N_8470,N_7446,N_7995);
and U8471 (N_8471,N_7461,N_7143);
and U8472 (N_8472,N_7559,N_7792);
or U8473 (N_8473,N_7885,N_7923);
or U8474 (N_8474,N_7641,N_7365);
and U8475 (N_8475,N_7562,N_7908);
xor U8476 (N_8476,N_7168,N_7813);
and U8477 (N_8477,N_7610,N_7205);
and U8478 (N_8478,N_7683,N_7808);
xor U8479 (N_8479,N_7053,N_7077);
and U8480 (N_8480,N_7310,N_7982);
xnor U8481 (N_8481,N_7812,N_7292);
nand U8482 (N_8482,N_7213,N_7718);
nor U8483 (N_8483,N_7269,N_7738);
nand U8484 (N_8484,N_7840,N_7560);
and U8485 (N_8485,N_7900,N_7920);
or U8486 (N_8486,N_7305,N_7627);
xor U8487 (N_8487,N_7193,N_7890);
and U8488 (N_8488,N_7003,N_7293);
nand U8489 (N_8489,N_7232,N_7376);
and U8490 (N_8490,N_7889,N_7063);
nand U8491 (N_8491,N_7782,N_7483);
nor U8492 (N_8492,N_7787,N_7608);
and U8493 (N_8493,N_7869,N_7616);
and U8494 (N_8494,N_7550,N_7039);
or U8495 (N_8495,N_7422,N_7546);
or U8496 (N_8496,N_7350,N_7614);
and U8497 (N_8497,N_7282,N_7372);
and U8498 (N_8498,N_7617,N_7932);
or U8499 (N_8499,N_7555,N_7194);
nand U8500 (N_8500,N_7324,N_7819);
or U8501 (N_8501,N_7982,N_7520);
and U8502 (N_8502,N_7175,N_7285);
nand U8503 (N_8503,N_7701,N_7192);
and U8504 (N_8504,N_7577,N_7982);
and U8505 (N_8505,N_7499,N_7982);
nand U8506 (N_8506,N_7405,N_7864);
nor U8507 (N_8507,N_7746,N_7361);
nand U8508 (N_8508,N_7312,N_7121);
xor U8509 (N_8509,N_7119,N_7784);
xnor U8510 (N_8510,N_7104,N_7730);
and U8511 (N_8511,N_7093,N_7020);
or U8512 (N_8512,N_7318,N_7566);
nor U8513 (N_8513,N_7145,N_7546);
nor U8514 (N_8514,N_7402,N_7643);
nor U8515 (N_8515,N_7214,N_7579);
nand U8516 (N_8516,N_7676,N_7491);
and U8517 (N_8517,N_7254,N_7377);
and U8518 (N_8518,N_7123,N_7161);
nand U8519 (N_8519,N_7481,N_7074);
nor U8520 (N_8520,N_7607,N_7533);
nand U8521 (N_8521,N_7538,N_7496);
nand U8522 (N_8522,N_7222,N_7109);
nor U8523 (N_8523,N_7221,N_7702);
xor U8524 (N_8524,N_7779,N_7258);
and U8525 (N_8525,N_7089,N_7447);
or U8526 (N_8526,N_7650,N_7921);
and U8527 (N_8527,N_7080,N_7032);
xnor U8528 (N_8528,N_7211,N_7527);
nand U8529 (N_8529,N_7057,N_7191);
nand U8530 (N_8530,N_7767,N_7981);
xnor U8531 (N_8531,N_7191,N_7083);
or U8532 (N_8532,N_7773,N_7027);
nor U8533 (N_8533,N_7272,N_7715);
nand U8534 (N_8534,N_7228,N_7947);
nand U8535 (N_8535,N_7477,N_7368);
or U8536 (N_8536,N_7553,N_7739);
and U8537 (N_8537,N_7414,N_7196);
xor U8538 (N_8538,N_7658,N_7832);
and U8539 (N_8539,N_7503,N_7337);
nand U8540 (N_8540,N_7713,N_7489);
nor U8541 (N_8541,N_7099,N_7761);
nor U8542 (N_8542,N_7926,N_7887);
and U8543 (N_8543,N_7230,N_7328);
and U8544 (N_8544,N_7837,N_7165);
or U8545 (N_8545,N_7152,N_7998);
and U8546 (N_8546,N_7407,N_7044);
nor U8547 (N_8547,N_7463,N_7794);
nand U8548 (N_8548,N_7127,N_7995);
nor U8549 (N_8549,N_7587,N_7162);
or U8550 (N_8550,N_7358,N_7831);
and U8551 (N_8551,N_7284,N_7730);
or U8552 (N_8552,N_7830,N_7326);
nor U8553 (N_8553,N_7385,N_7765);
nand U8554 (N_8554,N_7772,N_7737);
nor U8555 (N_8555,N_7148,N_7890);
nand U8556 (N_8556,N_7558,N_7794);
or U8557 (N_8557,N_7289,N_7010);
and U8558 (N_8558,N_7150,N_7578);
xnor U8559 (N_8559,N_7046,N_7077);
nor U8560 (N_8560,N_7969,N_7587);
or U8561 (N_8561,N_7773,N_7708);
and U8562 (N_8562,N_7377,N_7789);
nand U8563 (N_8563,N_7644,N_7330);
or U8564 (N_8564,N_7630,N_7651);
and U8565 (N_8565,N_7593,N_7475);
xnor U8566 (N_8566,N_7551,N_7811);
nand U8567 (N_8567,N_7671,N_7320);
and U8568 (N_8568,N_7517,N_7226);
nor U8569 (N_8569,N_7526,N_7387);
or U8570 (N_8570,N_7161,N_7898);
and U8571 (N_8571,N_7822,N_7650);
nor U8572 (N_8572,N_7246,N_7464);
nor U8573 (N_8573,N_7792,N_7781);
nor U8574 (N_8574,N_7075,N_7273);
and U8575 (N_8575,N_7453,N_7416);
xnor U8576 (N_8576,N_7940,N_7642);
and U8577 (N_8577,N_7924,N_7041);
or U8578 (N_8578,N_7467,N_7098);
and U8579 (N_8579,N_7452,N_7659);
or U8580 (N_8580,N_7482,N_7093);
nand U8581 (N_8581,N_7586,N_7244);
nor U8582 (N_8582,N_7568,N_7844);
xor U8583 (N_8583,N_7708,N_7074);
nor U8584 (N_8584,N_7491,N_7286);
nor U8585 (N_8585,N_7404,N_7739);
nor U8586 (N_8586,N_7206,N_7756);
and U8587 (N_8587,N_7045,N_7111);
or U8588 (N_8588,N_7566,N_7805);
or U8589 (N_8589,N_7497,N_7996);
nand U8590 (N_8590,N_7379,N_7253);
xnor U8591 (N_8591,N_7714,N_7325);
nand U8592 (N_8592,N_7179,N_7466);
xor U8593 (N_8593,N_7210,N_7339);
nor U8594 (N_8594,N_7354,N_7683);
nand U8595 (N_8595,N_7397,N_7360);
xnor U8596 (N_8596,N_7111,N_7148);
or U8597 (N_8597,N_7702,N_7557);
and U8598 (N_8598,N_7167,N_7501);
nor U8599 (N_8599,N_7122,N_7108);
xor U8600 (N_8600,N_7600,N_7003);
nor U8601 (N_8601,N_7229,N_7247);
xnor U8602 (N_8602,N_7195,N_7312);
and U8603 (N_8603,N_7725,N_7927);
and U8604 (N_8604,N_7626,N_7606);
xnor U8605 (N_8605,N_7646,N_7824);
and U8606 (N_8606,N_7324,N_7077);
xor U8607 (N_8607,N_7871,N_7009);
and U8608 (N_8608,N_7709,N_7088);
and U8609 (N_8609,N_7010,N_7896);
and U8610 (N_8610,N_7494,N_7705);
or U8611 (N_8611,N_7344,N_7264);
nand U8612 (N_8612,N_7897,N_7763);
nand U8613 (N_8613,N_7200,N_7280);
nand U8614 (N_8614,N_7564,N_7283);
xnor U8615 (N_8615,N_7842,N_7576);
xor U8616 (N_8616,N_7289,N_7210);
nand U8617 (N_8617,N_7327,N_7088);
nor U8618 (N_8618,N_7066,N_7319);
nand U8619 (N_8619,N_7596,N_7879);
and U8620 (N_8620,N_7799,N_7505);
xor U8621 (N_8621,N_7804,N_7148);
and U8622 (N_8622,N_7549,N_7109);
nand U8623 (N_8623,N_7132,N_7049);
and U8624 (N_8624,N_7691,N_7286);
nand U8625 (N_8625,N_7839,N_7761);
nor U8626 (N_8626,N_7525,N_7078);
or U8627 (N_8627,N_7762,N_7125);
or U8628 (N_8628,N_7009,N_7839);
and U8629 (N_8629,N_7754,N_7843);
and U8630 (N_8630,N_7777,N_7159);
nand U8631 (N_8631,N_7079,N_7387);
nand U8632 (N_8632,N_7982,N_7345);
and U8633 (N_8633,N_7342,N_7255);
nand U8634 (N_8634,N_7320,N_7407);
nor U8635 (N_8635,N_7203,N_7104);
and U8636 (N_8636,N_7897,N_7326);
nand U8637 (N_8637,N_7600,N_7072);
and U8638 (N_8638,N_7593,N_7006);
xor U8639 (N_8639,N_7816,N_7252);
nor U8640 (N_8640,N_7725,N_7690);
or U8641 (N_8641,N_7287,N_7306);
nand U8642 (N_8642,N_7056,N_7756);
nor U8643 (N_8643,N_7129,N_7425);
nand U8644 (N_8644,N_7539,N_7617);
nand U8645 (N_8645,N_7323,N_7369);
and U8646 (N_8646,N_7205,N_7640);
nor U8647 (N_8647,N_7168,N_7332);
or U8648 (N_8648,N_7927,N_7617);
or U8649 (N_8649,N_7430,N_7233);
nand U8650 (N_8650,N_7502,N_7454);
nor U8651 (N_8651,N_7828,N_7260);
nor U8652 (N_8652,N_7927,N_7460);
xor U8653 (N_8653,N_7478,N_7319);
or U8654 (N_8654,N_7340,N_7176);
nand U8655 (N_8655,N_7027,N_7820);
nand U8656 (N_8656,N_7022,N_7445);
xor U8657 (N_8657,N_7683,N_7949);
nand U8658 (N_8658,N_7323,N_7279);
nand U8659 (N_8659,N_7859,N_7801);
nor U8660 (N_8660,N_7848,N_7001);
and U8661 (N_8661,N_7844,N_7741);
nand U8662 (N_8662,N_7483,N_7497);
and U8663 (N_8663,N_7613,N_7210);
nor U8664 (N_8664,N_7396,N_7652);
and U8665 (N_8665,N_7431,N_7901);
and U8666 (N_8666,N_7630,N_7895);
or U8667 (N_8667,N_7532,N_7701);
or U8668 (N_8668,N_7504,N_7678);
and U8669 (N_8669,N_7142,N_7622);
or U8670 (N_8670,N_7320,N_7083);
or U8671 (N_8671,N_7015,N_7758);
or U8672 (N_8672,N_7879,N_7474);
xor U8673 (N_8673,N_7999,N_7544);
or U8674 (N_8674,N_7952,N_7511);
nand U8675 (N_8675,N_7839,N_7354);
nor U8676 (N_8676,N_7855,N_7411);
nor U8677 (N_8677,N_7516,N_7568);
and U8678 (N_8678,N_7199,N_7881);
or U8679 (N_8679,N_7059,N_7307);
and U8680 (N_8680,N_7752,N_7635);
or U8681 (N_8681,N_7463,N_7939);
or U8682 (N_8682,N_7763,N_7361);
nor U8683 (N_8683,N_7199,N_7819);
nand U8684 (N_8684,N_7861,N_7171);
nor U8685 (N_8685,N_7558,N_7370);
and U8686 (N_8686,N_7530,N_7592);
xor U8687 (N_8687,N_7520,N_7780);
xnor U8688 (N_8688,N_7178,N_7078);
xor U8689 (N_8689,N_7608,N_7553);
nor U8690 (N_8690,N_7802,N_7691);
nand U8691 (N_8691,N_7174,N_7991);
nor U8692 (N_8692,N_7289,N_7309);
nor U8693 (N_8693,N_7918,N_7541);
and U8694 (N_8694,N_7073,N_7882);
and U8695 (N_8695,N_7144,N_7954);
xor U8696 (N_8696,N_7590,N_7516);
nor U8697 (N_8697,N_7117,N_7879);
xnor U8698 (N_8698,N_7376,N_7022);
or U8699 (N_8699,N_7232,N_7766);
and U8700 (N_8700,N_7484,N_7719);
or U8701 (N_8701,N_7133,N_7357);
nand U8702 (N_8702,N_7002,N_7907);
nand U8703 (N_8703,N_7619,N_7360);
nor U8704 (N_8704,N_7271,N_7270);
and U8705 (N_8705,N_7516,N_7842);
nor U8706 (N_8706,N_7217,N_7292);
and U8707 (N_8707,N_7732,N_7704);
nand U8708 (N_8708,N_7315,N_7355);
or U8709 (N_8709,N_7237,N_7737);
xnor U8710 (N_8710,N_7049,N_7676);
or U8711 (N_8711,N_7062,N_7448);
or U8712 (N_8712,N_7853,N_7507);
nand U8713 (N_8713,N_7036,N_7496);
or U8714 (N_8714,N_7543,N_7696);
nand U8715 (N_8715,N_7923,N_7156);
nor U8716 (N_8716,N_7574,N_7609);
nand U8717 (N_8717,N_7470,N_7661);
nor U8718 (N_8718,N_7280,N_7729);
or U8719 (N_8719,N_7455,N_7293);
or U8720 (N_8720,N_7219,N_7046);
xnor U8721 (N_8721,N_7973,N_7953);
and U8722 (N_8722,N_7381,N_7624);
nor U8723 (N_8723,N_7727,N_7544);
and U8724 (N_8724,N_7208,N_7045);
xnor U8725 (N_8725,N_7958,N_7718);
nand U8726 (N_8726,N_7457,N_7791);
xnor U8727 (N_8727,N_7211,N_7052);
and U8728 (N_8728,N_7599,N_7267);
xor U8729 (N_8729,N_7954,N_7949);
nor U8730 (N_8730,N_7822,N_7803);
nand U8731 (N_8731,N_7966,N_7279);
and U8732 (N_8732,N_7296,N_7170);
nand U8733 (N_8733,N_7579,N_7109);
nor U8734 (N_8734,N_7395,N_7997);
xor U8735 (N_8735,N_7072,N_7345);
nand U8736 (N_8736,N_7226,N_7932);
and U8737 (N_8737,N_7178,N_7853);
and U8738 (N_8738,N_7661,N_7246);
nand U8739 (N_8739,N_7363,N_7295);
and U8740 (N_8740,N_7579,N_7608);
and U8741 (N_8741,N_7831,N_7422);
nand U8742 (N_8742,N_7925,N_7709);
or U8743 (N_8743,N_7583,N_7357);
or U8744 (N_8744,N_7519,N_7201);
or U8745 (N_8745,N_7945,N_7936);
nand U8746 (N_8746,N_7296,N_7466);
nor U8747 (N_8747,N_7715,N_7471);
nand U8748 (N_8748,N_7333,N_7997);
and U8749 (N_8749,N_7760,N_7985);
nand U8750 (N_8750,N_7319,N_7666);
xnor U8751 (N_8751,N_7860,N_7920);
and U8752 (N_8752,N_7057,N_7725);
or U8753 (N_8753,N_7624,N_7265);
and U8754 (N_8754,N_7831,N_7373);
nor U8755 (N_8755,N_7162,N_7935);
nor U8756 (N_8756,N_7377,N_7673);
nor U8757 (N_8757,N_7032,N_7605);
nor U8758 (N_8758,N_7561,N_7332);
xor U8759 (N_8759,N_7477,N_7579);
or U8760 (N_8760,N_7094,N_7580);
nor U8761 (N_8761,N_7127,N_7529);
or U8762 (N_8762,N_7456,N_7431);
and U8763 (N_8763,N_7112,N_7738);
nand U8764 (N_8764,N_7720,N_7437);
nor U8765 (N_8765,N_7900,N_7442);
nand U8766 (N_8766,N_7386,N_7096);
and U8767 (N_8767,N_7864,N_7808);
nor U8768 (N_8768,N_7204,N_7384);
nand U8769 (N_8769,N_7802,N_7811);
or U8770 (N_8770,N_7209,N_7223);
and U8771 (N_8771,N_7678,N_7018);
nand U8772 (N_8772,N_7430,N_7159);
or U8773 (N_8773,N_7206,N_7474);
nor U8774 (N_8774,N_7145,N_7366);
nor U8775 (N_8775,N_7884,N_7471);
and U8776 (N_8776,N_7210,N_7923);
and U8777 (N_8777,N_7433,N_7813);
or U8778 (N_8778,N_7714,N_7369);
nor U8779 (N_8779,N_7678,N_7728);
or U8780 (N_8780,N_7823,N_7773);
or U8781 (N_8781,N_7212,N_7495);
nor U8782 (N_8782,N_7937,N_7008);
xnor U8783 (N_8783,N_7299,N_7372);
and U8784 (N_8784,N_7729,N_7668);
and U8785 (N_8785,N_7016,N_7518);
and U8786 (N_8786,N_7193,N_7205);
xnor U8787 (N_8787,N_7410,N_7477);
nand U8788 (N_8788,N_7394,N_7549);
nand U8789 (N_8789,N_7039,N_7122);
nand U8790 (N_8790,N_7931,N_7471);
xnor U8791 (N_8791,N_7701,N_7997);
nand U8792 (N_8792,N_7703,N_7479);
or U8793 (N_8793,N_7988,N_7385);
and U8794 (N_8794,N_7494,N_7897);
xnor U8795 (N_8795,N_7338,N_7289);
nor U8796 (N_8796,N_7240,N_7741);
or U8797 (N_8797,N_7268,N_7324);
nand U8798 (N_8798,N_7767,N_7642);
nor U8799 (N_8799,N_7867,N_7760);
xor U8800 (N_8800,N_7505,N_7568);
nor U8801 (N_8801,N_7422,N_7184);
nand U8802 (N_8802,N_7992,N_7139);
and U8803 (N_8803,N_7461,N_7928);
and U8804 (N_8804,N_7629,N_7393);
and U8805 (N_8805,N_7220,N_7234);
xnor U8806 (N_8806,N_7814,N_7135);
nor U8807 (N_8807,N_7051,N_7757);
nand U8808 (N_8808,N_7899,N_7196);
xnor U8809 (N_8809,N_7322,N_7302);
and U8810 (N_8810,N_7333,N_7973);
or U8811 (N_8811,N_7786,N_7879);
nand U8812 (N_8812,N_7631,N_7294);
nor U8813 (N_8813,N_7365,N_7323);
nor U8814 (N_8814,N_7124,N_7828);
or U8815 (N_8815,N_7741,N_7026);
nor U8816 (N_8816,N_7752,N_7721);
nand U8817 (N_8817,N_7010,N_7378);
nand U8818 (N_8818,N_7391,N_7423);
nand U8819 (N_8819,N_7769,N_7790);
and U8820 (N_8820,N_7402,N_7796);
or U8821 (N_8821,N_7031,N_7861);
nand U8822 (N_8822,N_7785,N_7519);
nor U8823 (N_8823,N_7916,N_7989);
or U8824 (N_8824,N_7859,N_7280);
and U8825 (N_8825,N_7634,N_7227);
nand U8826 (N_8826,N_7300,N_7279);
or U8827 (N_8827,N_7455,N_7487);
and U8828 (N_8828,N_7398,N_7063);
nor U8829 (N_8829,N_7278,N_7960);
nor U8830 (N_8830,N_7599,N_7914);
nand U8831 (N_8831,N_7710,N_7713);
and U8832 (N_8832,N_7973,N_7436);
nor U8833 (N_8833,N_7675,N_7382);
nor U8834 (N_8834,N_7912,N_7657);
nand U8835 (N_8835,N_7535,N_7229);
nor U8836 (N_8836,N_7347,N_7245);
nor U8837 (N_8837,N_7154,N_7484);
nand U8838 (N_8838,N_7997,N_7166);
and U8839 (N_8839,N_7190,N_7324);
nor U8840 (N_8840,N_7624,N_7021);
or U8841 (N_8841,N_7203,N_7607);
or U8842 (N_8842,N_7674,N_7571);
nor U8843 (N_8843,N_7272,N_7378);
nand U8844 (N_8844,N_7978,N_7512);
or U8845 (N_8845,N_7261,N_7473);
nor U8846 (N_8846,N_7411,N_7500);
nor U8847 (N_8847,N_7999,N_7749);
and U8848 (N_8848,N_7282,N_7990);
and U8849 (N_8849,N_7322,N_7847);
nor U8850 (N_8850,N_7166,N_7871);
xor U8851 (N_8851,N_7687,N_7610);
or U8852 (N_8852,N_7516,N_7915);
and U8853 (N_8853,N_7388,N_7048);
xor U8854 (N_8854,N_7321,N_7181);
and U8855 (N_8855,N_7212,N_7064);
and U8856 (N_8856,N_7122,N_7350);
nand U8857 (N_8857,N_7692,N_7914);
and U8858 (N_8858,N_7095,N_7672);
nor U8859 (N_8859,N_7571,N_7946);
xor U8860 (N_8860,N_7736,N_7583);
and U8861 (N_8861,N_7428,N_7450);
xor U8862 (N_8862,N_7521,N_7454);
or U8863 (N_8863,N_7204,N_7940);
nor U8864 (N_8864,N_7987,N_7779);
nor U8865 (N_8865,N_7135,N_7610);
xnor U8866 (N_8866,N_7251,N_7515);
nor U8867 (N_8867,N_7755,N_7722);
nand U8868 (N_8868,N_7277,N_7049);
or U8869 (N_8869,N_7806,N_7064);
xor U8870 (N_8870,N_7054,N_7458);
xnor U8871 (N_8871,N_7619,N_7610);
nor U8872 (N_8872,N_7665,N_7562);
and U8873 (N_8873,N_7960,N_7723);
xnor U8874 (N_8874,N_7815,N_7125);
and U8875 (N_8875,N_7484,N_7869);
xnor U8876 (N_8876,N_7386,N_7824);
xnor U8877 (N_8877,N_7386,N_7184);
nand U8878 (N_8878,N_7432,N_7719);
and U8879 (N_8879,N_7801,N_7797);
nor U8880 (N_8880,N_7494,N_7459);
or U8881 (N_8881,N_7433,N_7496);
nor U8882 (N_8882,N_7656,N_7628);
nand U8883 (N_8883,N_7439,N_7021);
nor U8884 (N_8884,N_7057,N_7107);
nand U8885 (N_8885,N_7001,N_7775);
nor U8886 (N_8886,N_7997,N_7493);
and U8887 (N_8887,N_7756,N_7505);
or U8888 (N_8888,N_7876,N_7146);
xnor U8889 (N_8889,N_7624,N_7886);
and U8890 (N_8890,N_7449,N_7045);
nand U8891 (N_8891,N_7347,N_7830);
nor U8892 (N_8892,N_7957,N_7511);
nor U8893 (N_8893,N_7900,N_7919);
nor U8894 (N_8894,N_7922,N_7490);
and U8895 (N_8895,N_7705,N_7498);
or U8896 (N_8896,N_7471,N_7283);
nor U8897 (N_8897,N_7725,N_7534);
or U8898 (N_8898,N_7794,N_7386);
nor U8899 (N_8899,N_7109,N_7149);
nor U8900 (N_8900,N_7783,N_7447);
or U8901 (N_8901,N_7294,N_7731);
or U8902 (N_8902,N_7567,N_7911);
nor U8903 (N_8903,N_7615,N_7028);
or U8904 (N_8904,N_7614,N_7212);
nor U8905 (N_8905,N_7345,N_7435);
nor U8906 (N_8906,N_7382,N_7666);
and U8907 (N_8907,N_7201,N_7428);
nand U8908 (N_8908,N_7006,N_7465);
or U8909 (N_8909,N_7261,N_7317);
or U8910 (N_8910,N_7726,N_7286);
nand U8911 (N_8911,N_7499,N_7246);
or U8912 (N_8912,N_7053,N_7048);
nand U8913 (N_8913,N_7304,N_7278);
and U8914 (N_8914,N_7356,N_7898);
nand U8915 (N_8915,N_7409,N_7752);
nand U8916 (N_8916,N_7269,N_7137);
and U8917 (N_8917,N_7302,N_7117);
nand U8918 (N_8918,N_7534,N_7650);
and U8919 (N_8919,N_7233,N_7448);
nor U8920 (N_8920,N_7556,N_7086);
and U8921 (N_8921,N_7821,N_7419);
nand U8922 (N_8922,N_7476,N_7905);
nor U8923 (N_8923,N_7484,N_7428);
and U8924 (N_8924,N_7582,N_7210);
and U8925 (N_8925,N_7823,N_7890);
nor U8926 (N_8926,N_7402,N_7503);
or U8927 (N_8927,N_7336,N_7467);
xnor U8928 (N_8928,N_7372,N_7426);
or U8929 (N_8929,N_7580,N_7278);
nor U8930 (N_8930,N_7635,N_7369);
or U8931 (N_8931,N_7863,N_7896);
nand U8932 (N_8932,N_7692,N_7427);
nand U8933 (N_8933,N_7555,N_7629);
nand U8934 (N_8934,N_7922,N_7844);
nand U8935 (N_8935,N_7067,N_7059);
nor U8936 (N_8936,N_7821,N_7387);
nor U8937 (N_8937,N_7914,N_7392);
nor U8938 (N_8938,N_7090,N_7332);
nand U8939 (N_8939,N_7769,N_7044);
nor U8940 (N_8940,N_7489,N_7954);
or U8941 (N_8941,N_7819,N_7502);
nand U8942 (N_8942,N_7948,N_7856);
nor U8943 (N_8943,N_7699,N_7325);
nor U8944 (N_8944,N_7429,N_7594);
and U8945 (N_8945,N_7421,N_7299);
or U8946 (N_8946,N_7096,N_7649);
nand U8947 (N_8947,N_7280,N_7387);
nand U8948 (N_8948,N_7801,N_7649);
nand U8949 (N_8949,N_7438,N_7557);
nand U8950 (N_8950,N_7070,N_7348);
and U8951 (N_8951,N_7618,N_7208);
nand U8952 (N_8952,N_7529,N_7365);
xor U8953 (N_8953,N_7808,N_7195);
nor U8954 (N_8954,N_7152,N_7025);
xor U8955 (N_8955,N_7211,N_7924);
nand U8956 (N_8956,N_7450,N_7619);
nand U8957 (N_8957,N_7368,N_7703);
and U8958 (N_8958,N_7382,N_7600);
xor U8959 (N_8959,N_7488,N_7912);
nor U8960 (N_8960,N_7121,N_7036);
or U8961 (N_8961,N_7521,N_7672);
nor U8962 (N_8962,N_7955,N_7841);
or U8963 (N_8963,N_7773,N_7372);
nand U8964 (N_8964,N_7340,N_7253);
nor U8965 (N_8965,N_7742,N_7223);
nand U8966 (N_8966,N_7295,N_7829);
or U8967 (N_8967,N_7739,N_7266);
and U8968 (N_8968,N_7779,N_7874);
xnor U8969 (N_8969,N_7249,N_7961);
nor U8970 (N_8970,N_7614,N_7510);
xnor U8971 (N_8971,N_7396,N_7887);
nor U8972 (N_8972,N_7712,N_7388);
or U8973 (N_8973,N_7415,N_7302);
and U8974 (N_8974,N_7765,N_7836);
nor U8975 (N_8975,N_7343,N_7595);
nor U8976 (N_8976,N_7029,N_7248);
and U8977 (N_8977,N_7821,N_7512);
or U8978 (N_8978,N_7208,N_7124);
or U8979 (N_8979,N_7964,N_7536);
or U8980 (N_8980,N_7113,N_7428);
nand U8981 (N_8981,N_7063,N_7180);
nor U8982 (N_8982,N_7284,N_7344);
nand U8983 (N_8983,N_7604,N_7293);
nand U8984 (N_8984,N_7830,N_7181);
nor U8985 (N_8985,N_7966,N_7709);
or U8986 (N_8986,N_7722,N_7946);
nor U8987 (N_8987,N_7443,N_7374);
nor U8988 (N_8988,N_7161,N_7336);
nor U8989 (N_8989,N_7267,N_7046);
xor U8990 (N_8990,N_7780,N_7717);
nand U8991 (N_8991,N_7034,N_7917);
and U8992 (N_8992,N_7668,N_7466);
xnor U8993 (N_8993,N_7690,N_7875);
xnor U8994 (N_8994,N_7715,N_7226);
nor U8995 (N_8995,N_7324,N_7073);
or U8996 (N_8996,N_7159,N_7338);
nor U8997 (N_8997,N_7033,N_7007);
or U8998 (N_8998,N_7538,N_7037);
and U8999 (N_8999,N_7004,N_7313);
xor U9000 (N_9000,N_8832,N_8190);
and U9001 (N_9001,N_8641,N_8514);
and U9002 (N_9002,N_8588,N_8792);
or U9003 (N_9003,N_8130,N_8167);
nor U9004 (N_9004,N_8137,N_8296);
or U9005 (N_9005,N_8444,N_8540);
nand U9006 (N_9006,N_8652,N_8688);
xnor U9007 (N_9007,N_8060,N_8681);
nand U9008 (N_9008,N_8191,N_8057);
nor U9009 (N_9009,N_8156,N_8772);
nand U9010 (N_9010,N_8303,N_8608);
or U9011 (N_9011,N_8555,N_8087);
or U9012 (N_9012,N_8454,N_8751);
and U9013 (N_9013,N_8706,N_8918);
and U9014 (N_9014,N_8682,N_8865);
xor U9015 (N_9015,N_8725,N_8850);
nor U9016 (N_9016,N_8929,N_8013);
nand U9017 (N_9017,N_8058,N_8789);
xor U9018 (N_9018,N_8234,N_8068);
xor U9019 (N_9019,N_8487,N_8337);
nor U9020 (N_9020,N_8081,N_8469);
nor U9021 (N_9021,N_8025,N_8007);
xnor U9022 (N_9022,N_8204,N_8536);
or U9023 (N_9023,N_8127,N_8786);
or U9024 (N_9024,N_8312,N_8619);
nor U9025 (N_9025,N_8072,N_8959);
or U9026 (N_9026,N_8745,N_8175);
xor U9027 (N_9027,N_8217,N_8197);
nor U9028 (N_9028,N_8790,N_8675);
nor U9029 (N_9029,N_8853,N_8680);
nor U9030 (N_9030,N_8339,N_8036);
and U9031 (N_9031,N_8991,N_8542);
and U9032 (N_9032,N_8676,N_8791);
and U9033 (N_9033,N_8027,N_8898);
or U9034 (N_9034,N_8620,N_8963);
and U9035 (N_9035,N_8402,N_8131);
nor U9036 (N_9036,N_8064,N_8823);
nand U9037 (N_9037,N_8075,N_8389);
or U9038 (N_9038,N_8358,N_8295);
and U9039 (N_9039,N_8925,N_8494);
nor U9040 (N_9040,N_8951,N_8926);
nand U9041 (N_9041,N_8315,N_8924);
or U9042 (N_9042,N_8121,N_8887);
xor U9043 (N_9043,N_8096,N_8777);
and U9044 (N_9044,N_8435,N_8573);
or U9045 (N_9045,N_8908,N_8106);
and U9046 (N_9046,N_8883,N_8592);
or U9047 (N_9047,N_8351,N_8231);
or U9048 (N_9048,N_8211,N_8802);
and U9049 (N_9049,N_8507,N_8974);
or U9050 (N_9050,N_8519,N_8289);
nand U9051 (N_9051,N_8903,N_8492);
and U9052 (N_9052,N_8896,N_8525);
nor U9053 (N_9053,N_8173,N_8817);
nor U9054 (N_9054,N_8660,N_8651);
and U9055 (N_9055,N_8687,N_8664);
or U9056 (N_9056,N_8272,N_8366);
nor U9057 (N_9057,N_8223,N_8143);
and U9058 (N_9058,N_8799,N_8214);
and U9059 (N_9059,N_8819,N_8014);
or U9060 (N_9060,N_8711,N_8856);
nand U9061 (N_9061,N_8637,N_8810);
nand U9062 (N_9062,N_8804,N_8553);
nor U9063 (N_9063,N_8931,N_8394);
or U9064 (N_9064,N_8348,N_8370);
or U9065 (N_9065,N_8615,N_8414);
and U9066 (N_9066,N_8873,N_8093);
and U9067 (N_9067,N_8142,N_8026);
or U9068 (N_9068,N_8294,N_8219);
nor U9069 (N_9069,N_8482,N_8771);
or U9070 (N_9070,N_8645,N_8779);
nand U9071 (N_9071,N_8415,N_8362);
or U9072 (N_9072,N_8486,N_8806);
and U9073 (N_9073,N_8907,N_8445);
and U9074 (N_9074,N_8811,N_8686);
or U9075 (N_9075,N_8148,N_8077);
nand U9076 (N_9076,N_8201,N_8511);
or U9077 (N_9077,N_8422,N_8760);
nand U9078 (N_9078,N_8404,N_8338);
or U9079 (N_9079,N_8446,N_8563);
xnor U9080 (N_9080,N_8943,N_8580);
nand U9081 (N_9081,N_8576,N_8083);
or U9082 (N_9082,N_8617,N_8203);
xor U9083 (N_9083,N_8374,N_8601);
nor U9084 (N_9084,N_8528,N_8015);
and U9085 (N_9085,N_8185,N_8129);
and U9086 (N_9086,N_8597,N_8793);
nor U9087 (N_9087,N_8766,N_8661);
or U9088 (N_9088,N_8040,N_8120);
nand U9089 (N_9089,N_8632,N_8248);
nand U9090 (N_9090,N_8677,N_8202);
nor U9091 (N_9091,N_8852,N_8816);
or U9092 (N_9092,N_8221,N_8023);
nand U9093 (N_9093,N_8070,N_8471);
or U9094 (N_9094,N_8421,N_8773);
and U9095 (N_9095,N_8569,N_8470);
or U9096 (N_9096,N_8061,N_8610);
xnor U9097 (N_9097,N_8624,N_8979);
nand U9098 (N_9098,N_8562,N_8603);
nor U9099 (N_9099,N_8043,N_8798);
xor U9100 (N_9100,N_8073,N_8813);
nor U9101 (N_9101,N_8183,N_8359);
and U9102 (N_9102,N_8177,N_8721);
xor U9103 (N_9103,N_8133,N_8674);
xor U9104 (N_9104,N_8892,N_8334);
or U9105 (N_9105,N_8376,N_8499);
nand U9106 (N_9106,N_8824,N_8483);
nor U9107 (N_9107,N_8350,N_8265);
and U9108 (N_9108,N_8094,N_8554);
and U9109 (N_9109,N_8559,N_8988);
nand U9110 (N_9110,N_8179,N_8548);
xnor U9111 (N_9111,N_8273,N_8134);
nor U9112 (N_9112,N_8982,N_8886);
nand U9113 (N_9113,N_8089,N_8700);
nor U9114 (N_9114,N_8616,N_8729);
or U9115 (N_9115,N_8938,N_8801);
nor U9116 (N_9116,N_8961,N_8270);
nand U9117 (N_9117,N_8010,N_8168);
nand U9118 (N_9118,N_8233,N_8648);
nor U9119 (N_9119,N_8037,N_8478);
or U9120 (N_9120,N_8349,N_8847);
or U9121 (N_9121,N_8080,N_8556);
nand U9122 (N_9122,N_8385,N_8047);
xor U9123 (N_9123,N_8479,N_8713);
or U9124 (N_9124,N_8984,N_8837);
or U9125 (N_9125,N_8689,N_8267);
xnor U9126 (N_9126,N_8715,N_8112);
and U9127 (N_9127,N_8243,N_8218);
or U9128 (N_9128,N_8612,N_8602);
or U9129 (N_9129,N_8298,N_8780);
and U9130 (N_9130,N_8379,N_8972);
nor U9131 (N_9131,N_8305,N_8508);
or U9132 (N_9132,N_8044,N_8291);
nor U9133 (N_9133,N_8405,N_8574);
xor U9134 (N_9134,N_8503,N_8899);
or U9135 (N_9135,N_8720,N_8498);
nand U9136 (N_9136,N_8363,N_8105);
nor U9137 (N_9137,N_8212,N_8467);
nand U9138 (N_9138,N_8252,N_8322);
and U9139 (N_9139,N_8744,N_8008);
and U9140 (N_9140,N_8095,N_8749);
and U9141 (N_9141,N_8333,N_8730);
and U9142 (N_9142,N_8258,N_8942);
and U9143 (N_9143,N_8284,N_8532);
nand U9144 (N_9144,N_8262,N_8182);
and U9145 (N_9145,N_8826,N_8572);
or U9146 (N_9146,N_8079,N_8714);
nor U9147 (N_9147,N_8885,N_8048);
nor U9148 (N_9148,N_8424,N_8859);
and U9149 (N_9149,N_8066,N_8902);
nor U9150 (N_9150,N_8236,N_8210);
and U9151 (N_9151,N_8353,N_8582);
and U9152 (N_9152,N_8022,N_8287);
nor U9153 (N_9153,N_8906,N_8945);
and U9154 (N_9154,N_8875,N_8957);
and U9155 (N_9155,N_8250,N_8631);
xor U9156 (N_9156,N_8895,N_8088);
nand U9157 (N_9157,N_8172,N_8855);
nor U9158 (N_9158,N_8516,N_8276);
nor U9159 (N_9159,N_8719,N_8384);
nor U9160 (N_9160,N_8980,N_8805);
nand U9161 (N_9161,N_8230,N_8831);
nand U9162 (N_9162,N_8456,N_8227);
nor U9163 (N_9163,N_8736,N_8235);
nand U9164 (N_9164,N_8481,N_8990);
and U9165 (N_9165,N_8878,N_8987);
or U9166 (N_9166,N_8785,N_8975);
or U9167 (N_9167,N_8994,N_8739);
xnor U9168 (N_9168,N_8319,N_8141);
and U9169 (N_9169,N_8858,N_8473);
nor U9170 (N_9170,N_8364,N_8417);
and U9171 (N_9171,N_8992,N_8288);
or U9172 (N_9172,N_8413,N_8433);
nor U9173 (N_9173,N_8625,N_8577);
nor U9174 (N_9174,N_8600,N_8151);
and U9175 (N_9175,N_8090,N_8844);
or U9176 (N_9176,N_8448,N_8327);
nor U9177 (N_9177,N_8455,N_8623);
and U9178 (N_9178,N_8189,N_8461);
or U9179 (N_9179,N_8253,N_8472);
nor U9180 (N_9180,N_8357,N_8225);
or U9181 (N_9181,N_8004,N_8005);
xnor U9182 (N_9182,N_8419,N_8505);
and U9183 (N_9183,N_8439,N_8849);
nor U9184 (N_9184,N_8378,N_8782);
or U9185 (N_9185,N_8176,N_8956);
and U9186 (N_9186,N_8642,N_8520);
nand U9187 (N_9187,N_8398,N_8738);
nor U9188 (N_9188,N_8981,N_8937);
nor U9189 (N_9189,N_8775,N_8740);
or U9190 (N_9190,N_8857,N_8800);
nand U9191 (N_9191,N_8006,N_8890);
nand U9192 (N_9192,N_8116,N_8474);
nand U9193 (N_9193,N_8476,N_8071);
or U9194 (N_9194,N_8587,N_8867);
and U9195 (N_9195,N_8368,N_8581);
nand U9196 (N_9196,N_8659,N_8283);
and U9197 (N_9197,N_8955,N_8281);
or U9198 (N_9198,N_8764,N_8643);
nand U9199 (N_9199,N_8526,N_8716);
or U9200 (N_9200,N_8663,N_8242);
or U9201 (N_9201,N_8369,N_8840);
xnor U9202 (N_9202,N_8449,N_8732);
nor U9203 (N_9203,N_8578,N_8459);
or U9204 (N_9204,N_8690,N_8078);
nand U9205 (N_9205,N_8174,N_8407);
and U9206 (N_9206,N_8484,N_8488);
nor U9207 (N_9207,N_8579,N_8551);
nor U9208 (N_9208,N_8451,N_8159);
and U9209 (N_9209,N_8052,N_8535);
nand U9210 (N_9210,N_8564,N_8460);
nor U9211 (N_9211,N_8967,N_8640);
and U9212 (N_9212,N_8397,N_8746);
and U9213 (N_9213,N_8101,N_8808);
and U9214 (N_9214,N_8029,N_8846);
or U9215 (N_9215,N_8973,N_8051);
nor U9216 (N_9216,N_8868,N_8910);
nor U9217 (N_9217,N_8316,N_8544);
nand U9218 (N_9218,N_8876,N_8392);
nand U9219 (N_9219,N_8821,N_8621);
xor U9220 (N_9220,N_8927,N_8274);
and U9221 (N_9221,N_8718,N_8110);
nor U9222 (N_9222,N_8122,N_8011);
and U9223 (N_9223,N_8879,N_8263);
or U9224 (N_9224,N_8067,N_8438);
and U9225 (N_9225,N_8709,N_8205);
nor U9226 (N_9226,N_8665,N_8904);
or U9227 (N_9227,N_8033,N_8053);
or U9228 (N_9228,N_8627,N_8325);
nand U9229 (N_9229,N_8426,N_8605);
and U9230 (N_9230,N_8125,N_8136);
nand U9231 (N_9231,N_8935,N_8107);
nand U9232 (N_9232,N_8039,N_8443);
and U9233 (N_9233,N_8765,N_8226);
and U9234 (N_9234,N_8045,N_8939);
or U9235 (N_9235,N_8517,N_8543);
or U9236 (N_9236,N_8518,N_8649);
and U9237 (N_9237,N_8796,N_8871);
or U9238 (N_9238,N_8123,N_8054);
or U9239 (N_9239,N_8373,N_8560);
nand U9240 (N_9240,N_8703,N_8475);
and U9241 (N_9241,N_8377,N_8157);
nand U9242 (N_9242,N_8031,N_8237);
and U9243 (N_9243,N_8038,N_8271);
and U9244 (N_9244,N_8671,N_8309);
nor U9245 (N_9245,N_8318,N_8021);
nor U9246 (N_9246,N_8001,N_8256);
nor U9247 (N_9247,N_8758,N_8198);
or U9248 (N_9248,N_8386,N_8229);
or U9249 (N_9249,N_8457,N_8825);
or U9250 (N_9250,N_8917,N_8523);
and U9251 (N_9251,N_8841,N_8091);
nor U9252 (N_9252,N_8418,N_8894);
or U9253 (N_9253,N_8335,N_8650);
and U9254 (N_9254,N_8874,N_8585);
nand U9255 (N_9255,N_8017,N_8900);
or U9256 (N_9256,N_8084,N_8261);
or U9257 (N_9257,N_8326,N_8538);
or U9258 (N_9258,N_8332,N_8797);
or U9259 (N_9259,N_8440,N_8646);
nand U9260 (N_9260,N_8341,N_8647);
and U9261 (N_9261,N_8656,N_8814);
or U9262 (N_9262,N_8016,N_8035);
xor U9263 (N_9263,N_8864,N_8324);
xor U9264 (N_9264,N_8727,N_8835);
nand U9265 (N_9265,N_8952,N_8195);
nor U9266 (N_9266,N_8977,N_8639);
or U9267 (N_9267,N_8609,N_8742);
or U9268 (N_9268,N_8493,N_8161);
xor U9269 (N_9269,N_8187,N_8254);
nand U9270 (N_9270,N_8784,N_8403);
or U9271 (N_9271,N_8770,N_8200);
and U9272 (N_9272,N_8845,N_8126);
nor U9273 (N_9273,N_8763,N_8442);
nor U9274 (N_9274,N_8290,N_8117);
nand U9275 (N_9275,N_8178,N_8683);
nor U9276 (N_9276,N_8372,N_8300);
and U9277 (N_9277,N_8521,N_8224);
nor U9278 (N_9278,N_8111,N_8003);
and U9279 (N_9279,N_8983,N_8192);
xor U9280 (N_9280,N_8590,N_8583);
or U9281 (N_9281,N_8065,N_8976);
xor U9282 (N_9282,N_8969,N_8566);
or U9283 (N_9283,N_8812,N_8728);
nor U9284 (N_9284,N_8997,N_8251);
and U9285 (N_9285,N_8153,N_8400);
or U9286 (N_9286,N_8306,N_8541);
or U9287 (N_9287,N_8795,N_8589);
and U9288 (N_9288,N_8074,N_8940);
nor U9289 (N_9289,N_8346,N_8128);
nand U9290 (N_9290,N_8416,N_8496);
or U9291 (N_9291,N_8032,N_8345);
or U9292 (N_9292,N_8781,N_8552);
xnor U9293 (N_9293,N_8815,N_8870);
or U9294 (N_9294,N_8743,N_8794);
and U9295 (N_9295,N_8410,N_8667);
nand U9296 (N_9296,N_8998,N_8034);
xnor U9297 (N_9297,N_8238,N_8666);
and U9298 (N_9298,N_8750,N_8776);
nor U9299 (N_9299,N_8558,N_8606);
and U9300 (N_9300,N_8186,N_8654);
and U9301 (N_9301,N_8302,N_8921);
and U9302 (N_9302,N_8299,N_8170);
nand U9303 (N_9303,N_8266,N_8930);
nor U9304 (N_9304,N_8365,N_8063);
and U9305 (N_9305,N_8247,N_8042);
and U9306 (N_9306,N_8323,N_8028);
and U9307 (N_9307,N_8055,N_8644);
and U9308 (N_9308,N_8999,N_8568);
or U9309 (N_9309,N_8638,N_8628);
xor U9310 (N_9310,N_8390,N_8259);
nand U9311 (N_9311,N_8428,N_8731);
nand U9312 (N_9312,N_8452,N_8836);
xor U9313 (N_9313,N_8901,N_8391);
nand U9314 (N_9314,N_8171,N_8916);
and U9315 (N_9315,N_8704,N_8082);
nand U9316 (N_9316,N_8249,N_8950);
nand U9317 (N_9317,N_8881,N_8000);
or U9318 (N_9318,N_8759,N_8480);
nor U9319 (N_9319,N_8539,N_8513);
nand U9320 (N_9320,N_8747,N_8947);
nand U9321 (N_9321,N_8355,N_8504);
nor U9322 (N_9322,N_8018,N_8944);
nor U9323 (N_9323,N_8375,N_8685);
xor U9324 (N_9324,N_8423,N_8477);
nand U9325 (N_9325,N_8872,N_8336);
or U9326 (N_9326,N_8458,N_8207);
and U9327 (N_9327,N_8599,N_8100);
and U9328 (N_9328,N_8510,N_8436);
or U9329 (N_9329,N_8260,N_8549);
nor U9330 (N_9330,N_8596,N_8147);
nor U9331 (N_9331,N_8672,N_8367);
nor U9332 (N_9332,N_8277,N_8395);
xor U9333 (N_9333,N_8245,N_8705);
and U9334 (N_9334,N_8124,N_8684);
nor U9335 (N_9335,N_8860,N_8630);
or U9336 (N_9336,N_8635,N_8618);
nor U9337 (N_9337,N_8432,N_8188);
nand U9338 (N_9338,N_8320,N_8669);
and U9339 (N_9339,N_8928,N_8429);
nor U9340 (N_9340,N_8607,N_8138);
nand U9341 (N_9341,N_8464,N_8030);
nand U9342 (N_9342,N_8614,N_8862);
xor U9343 (N_9343,N_8557,N_8206);
or U9344 (N_9344,N_8149,N_8912);
nor U9345 (N_9345,N_8968,N_8531);
nand U9346 (N_9346,N_8570,N_8949);
or U9347 (N_9347,N_8527,N_8502);
nor U9348 (N_9348,N_8411,N_8024);
nand U9349 (N_9349,N_8293,N_8232);
or U9350 (N_9350,N_8059,N_8501);
nor U9351 (N_9351,N_8604,N_8241);
xor U9352 (N_9352,N_8803,N_8098);
nand U9353 (N_9353,N_8522,N_8104);
or U9354 (N_9354,N_8915,N_8753);
and U9355 (N_9355,N_8196,N_8297);
xor U9356 (N_9356,N_8882,N_8833);
nor U9357 (N_9357,N_8113,N_8936);
nor U9358 (N_9358,N_8160,N_8702);
or U9359 (N_9359,N_8768,N_8971);
and U9360 (N_9360,N_8118,N_8893);
nand U9361 (N_9361,N_8228,N_8960);
nand U9362 (N_9362,N_8958,N_8565);
xor U9363 (N_9363,N_8550,N_8877);
or U9364 (N_9364,N_8809,N_8489);
or U9365 (N_9365,N_8655,N_8807);
and U9366 (N_9366,N_8437,N_8537);
xor U9367 (N_9367,N_8158,N_8985);
xnor U9368 (N_9368,N_8453,N_8280);
nand U9369 (N_9369,N_8450,N_8629);
nand U9370 (N_9370,N_8839,N_8425);
and U9371 (N_9371,N_8653,N_8076);
nand U9372 (N_9372,N_8636,N_8115);
and U9373 (N_9373,N_8056,N_8757);
and U9374 (N_9374,N_8275,N_8490);
and U9375 (N_9375,N_8408,N_8679);
and U9376 (N_9376,N_8530,N_8342);
xnor U9377 (N_9377,N_8818,N_8279);
nor U9378 (N_9378,N_8571,N_8184);
or U9379 (N_9379,N_8344,N_8880);
nor U9380 (N_9380,N_8891,N_8140);
nand U9381 (N_9381,N_8012,N_8097);
xor U9382 (N_9382,N_8748,N_8723);
or U9383 (N_9383,N_8466,N_8662);
and U9384 (N_9384,N_8694,N_8500);
and U9385 (N_9385,N_8381,N_8388);
and U9386 (N_9386,N_8953,N_8310);
or U9387 (N_9387,N_8257,N_8282);
nor U9388 (N_9388,N_8354,N_8180);
or U9389 (N_9389,N_8595,N_8162);
and U9390 (N_9390,N_8626,N_8062);
or U9391 (N_9391,N_8695,N_8427);
and U9392 (N_9392,N_8215,N_8752);
and U9393 (N_9393,N_8163,N_8829);
xor U9394 (N_9394,N_8146,N_8888);
nor U9395 (N_9395,N_8524,N_8092);
or U9396 (N_9396,N_8827,N_8668);
or U9397 (N_9397,N_8399,N_8409);
or U9398 (N_9398,N_8099,N_8986);
nand U9399 (N_9399,N_8380,N_8495);
or U9400 (N_9400,N_8246,N_8382);
nand U9401 (N_9401,N_8737,N_8307);
nand U9402 (N_9402,N_8598,N_8547);
nand U9403 (N_9403,N_8164,N_8165);
and U9404 (N_9404,N_8948,N_8707);
nand U9405 (N_9405,N_8889,N_8993);
nand U9406 (N_9406,N_8828,N_8561);
and U9407 (N_9407,N_8697,N_8468);
xor U9408 (N_9408,N_8778,N_8869);
or U9409 (N_9409,N_8329,N_8995);
nor U9410 (N_9410,N_8155,N_8774);
and U9411 (N_9411,N_8041,N_8584);
or U9412 (N_9412,N_8002,N_8866);
xnor U9413 (N_9413,N_8360,N_8788);
nor U9414 (N_9414,N_8678,N_8966);
nor U9415 (N_9415,N_8199,N_8691);
xnor U9416 (N_9416,N_8301,N_8069);
nand U9417 (N_9417,N_8670,N_8328);
nor U9418 (N_9418,N_8304,N_8311);
xor U9419 (N_9419,N_8401,N_8135);
or U9420 (N_9420,N_8923,N_8086);
nor U9421 (N_9421,N_8352,N_8420);
and U9422 (N_9422,N_8657,N_8208);
xor U9423 (N_9423,N_8497,N_8108);
nand U9424 (N_9424,N_8506,N_8330);
nor U9425 (N_9425,N_8244,N_8314);
and U9426 (N_9426,N_8693,N_8181);
and U9427 (N_9427,N_8139,N_8696);
nand U9428 (N_9428,N_8383,N_8533);
nor U9429 (N_9429,N_8019,N_8361);
nand U9430 (N_9430,N_8269,N_8613);
nor U9431 (N_9431,N_8989,N_8848);
and U9432 (N_9432,N_8712,N_8692);
nand U9433 (N_9433,N_8546,N_8726);
nor U9434 (N_9434,N_8634,N_8240);
and U9435 (N_9435,N_8050,N_8529);
and U9436 (N_9436,N_8913,N_8762);
nand U9437 (N_9437,N_8049,N_8434);
nor U9438 (N_9438,N_8462,N_8114);
xor U9439 (N_9439,N_8340,N_8854);
or U9440 (N_9440,N_8193,N_8996);
and U9441 (N_9441,N_8756,N_8843);
xor U9442 (N_9442,N_8863,N_8264);
nor U9443 (N_9443,N_8343,N_8658);
or U9444 (N_9444,N_8255,N_8046);
and U9445 (N_9445,N_8145,N_8321);
xnor U9446 (N_9446,N_8308,N_8717);
and U9447 (N_9447,N_8393,N_8209);
and U9448 (N_9448,N_8509,N_8194);
and U9449 (N_9449,N_8946,N_8216);
nand U9450 (N_9450,N_8734,N_8964);
or U9451 (N_9451,N_8861,N_8586);
nor U9452 (N_9452,N_8922,N_8905);
xnor U9453 (N_9453,N_8965,N_8754);
nor U9454 (N_9454,N_8396,N_8673);
nand U9455 (N_9455,N_8842,N_8701);
and U9456 (N_9456,N_8169,N_8755);
and U9457 (N_9457,N_8594,N_8278);
nor U9458 (N_9458,N_8708,N_8769);
xor U9459 (N_9459,N_8285,N_8783);
or U9460 (N_9460,N_8699,N_8724);
nand U9461 (N_9461,N_8591,N_8109);
nand U9462 (N_9462,N_8710,N_8911);
or U9463 (N_9463,N_8698,N_8933);
nand U9464 (N_9464,N_8430,N_8102);
nand U9465 (N_9465,N_8932,N_8622);
or U9466 (N_9466,N_8633,N_8970);
xnor U9467 (N_9467,N_8962,N_8431);
or U9468 (N_9468,N_8220,N_8593);
or U9469 (N_9469,N_8914,N_8735);
and U9470 (N_9470,N_8838,N_8465);
nand U9471 (N_9471,N_8834,N_8347);
and U9472 (N_9472,N_8515,N_8761);
nand U9473 (N_9473,N_8213,N_8317);
nor U9474 (N_9474,N_8512,N_8441);
or U9475 (N_9475,N_8820,N_8741);
or U9476 (N_9476,N_8897,N_8150);
nor U9477 (N_9477,N_8239,N_8103);
nand U9478 (N_9478,N_8292,N_8406);
nand U9479 (N_9479,N_8222,N_8934);
and U9480 (N_9480,N_8767,N_8412);
nand U9481 (N_9481,N_8387,N_8491);
nand U9482 (N_9482,N_8463,N_8020);
or U9483 (N_9483,N_8909,N_8009);
or U9484 (N_9484,N_8722,N_8447);
nor U9485 (N_9485,N_8822,N_8567);
or U9486 (N_9486,N_8851,N_8534);
nor U9487 (N_9487,N_8144,N_8919);
nand U9488 (N_9488,N_8884,N_8152);
nor U9489 (N_9489,N_8545,N_8978);
or U9490 (N_9490,N_8371,N_8941);
xnor U9491 (N_9491,N_8787,N_8166);
nand U9492 (N_9492,N_8119,N_8954);
or U9493 (N_9493,N_8313,N_8575);
and U9494 (N_9494,N_8331,N_8611);
nand U9495 (N_9495,N_8485,N_8356);
and U9496 (N_9496,N_8154,N_8286);
nand U9497 (N_9497,N_8268,N_8085);
nand U9498 (N_9498,N_8920,N_8132);
or U9499 (N_9499,N_8830,N_8733);
nor U9500 (N_9500,N_8402,N_8801);
and U9501 (N_9501,N_8453,N_8959);
nor U9502 (N_9502,N_8929,N_8928);
or U9503 (N_9503,N_8000,N_8915);
nor U9504 (N_9504,N_8307,N_8823);
and U9505 (N_9505,N_8708,N_8838);
nand U9506 (N_9506,N_8230,N_8240);
nand U9507 (N_9507,N_8019,N_8237);
nor U9508 (N_9508,N_8068,N_8391);
nor U9509 (N_9509,N_8038,N_8507);
nand U9510 (N_9510,N_8885,N_8732);
and U9511 (N_9511,N_8000,N_8226);
or U9512 (N_9512,N_8829,N_8260);
or U9513 (N_9513,N_8738,N_8299);
and U9514 (N_9514,N_8597,N_8533);
nand U9515 (N_9515,N_8642,N_8316);
nand U9516 (N_9516,N_8435,N_8624);
or U9517 (N_9517,N_8955,N_8614);
or U9518 (N_9518,N_8280,N_8795);
xnor U9519 (N_9519,N_8735,N_8201);
nand U9520 (N_9520,N_8596,N_8295);
and U9521 (N_9521,N_8114,N_8353);
nor U9522 (N_9522,N_8769,N_8954);
or U9523 (N_9523,N_8800,N_8215);
and U9524 (N_9524,N_8373,N_8251);
or U9525 (N_9525,N_8921,N_8437);
nand U9526 (N_9526,N_8198,N_8214);
nor U9527 (N_9527,N_8408,N_8905);
or U9528 (N_9528,N_8238,N_8211);
or U9529 (N_9529,N_8167,N_8669);
nand U9530 (N_9530,N_8326,N_8047);
or U9531 (N_9531,N_8377,N_8562);
and U9532 (N_9532,N_8699,N_8284);
nor U9533 (N_9533,N_8856,N_8683);
xnor U9534 (N_9534,N_8915,N_8748);
and U9535 (N_9535,N_8980,N_8607);
xor U9536 (N_9536,N_8131,N_8310);
nand U9537 (N_9537,N_8575,N_8102);
nand U9538 (N_9538,N_8147,N_8271);
or U9539 (N_9539,N_8260,N_8998);
nand U9540 (N_9540,N_8651,N_8729);
or U9541 (N_9541,N_8890,N_8547);
nor U9542 (N_9542,N_8549,N_8867);
nor U9543 (N_9543,N_8163,N_8851);
and U9544 (N_9544,N_8324,N_8145);
xnor U9545 (N_9545,N_8081,N_8604);
and U9546 (N_9546,N_8505,N_8571);
nor U9547 (N_9547,N_8602,N_8231);
or U9548 (N_9548,N_8756,N_8990);
nor U9549 (N_9549,N_8316,N_8110);
or U9550 (N_9550,N_8325,N_8862);
nand U9551 (N_9551,N_8742,N_8996);
and U9552 (N_9552,N_8209,N_8047);
nand U9553 (N_9553,N_8929,N_8768);
or U9554 (N_9554,N_8472,N_8917);
or U9555 (N_9555,N_8381,N_8199);
and U9556 (N_9556,N_8947,N_8598);
and U9557 (N_9557,N_8328,N_8697);
nor U9558 (N_9558,N_8331,N_8258);
and U9559 (N_9559,N_8551,N_8630);
nor U9560 (N_9560,N_8928,N_8310);
or U9561 (N_9561,N_8148,N_8682);
nand U9562 (N_9562,N_8048,N_8112);
nand U9563 (N_9563,N_8442,N_8891);
and U9564 (N_9564,N_8247,N_8641);
and U9565 (N_9565,N_8382,N_8802);
nor U9566 (N_9566,N_8936,N_8528);
and U9567 (N_9567,N_8542,N_8891);
nand U9568 (N_9568,N_8492,N_8992);
nor U9569 (N_9569,N_8879,N_8428);
or U9570 (N_9570,N_8628,N_8539);
and U9571 (N_9571,N_8167,N_8834);
and U9572 (N_9572,N_8203,N_8412);
nand U9573 (N_9573,N_8118,N_8127);
nor U9574 (N_9574,N_8239,N_8620);
and U9575 (N_9575,N_8715,N_8041);
nand U9576 (N_9576,N_8471,N_8869);
nand U9577 (N_9577,N_8944,N_8779);
xnor U9578 (N_9578,N_8309,N_8630);
nand U9579 (N_9579,N_8869,N_8329);
and U9580 (N_9580,N_8461,N_8820);
nor U9581 (N_9581,N_8982,N_8622);
and U9582 (N_9582,N_8614,N_8578);
and U9583 (N_9583,N_8062,N_8215);
nor U9584 (N_9584,N_8021,N_8478);
or U9585 (N_9585,N_8537,N_8785);
xor U9586 (N_9586,N_8247,N_8970);
and U9587 (N_9587,N_8715,N_8447);
or U9588 (N_9588,N_8588,N_8274);
or U9589 (N_9589,N_8379,N_8824);
nor U9590 (N_9590,N_8276,N_8903);
or U9591 (N_9591,N_8509,N_8097);
nor U9592 (N_9592,N_8503,N_8488);
and U9593 (N_9593,N_8179,N_8214);
and U9594 (N_9594,N_8062,N_8776);
and U9595 (N_9595,N_8833,N_8003);
and U9596 (N_9596,N_8907,N_8962);
nor U9597 (N_9597,N_8407,N_8797);
or U9598 (N_9598,N_8821,N_8192);
and U9599 (N_9599,N_8618,N_8214);
and U9600 (N_9600,N_8221,N_8369);
nor U9601 (N_9601,N_8305,N_8352);
nor U9602 (N_9602,N_8331,N_8334);
nand U9603 (N_9603,N_8328,N_8623);
and U9604 (N_9604,N_8415,N_8596);
xor U9605 (N_9605,N_8961,N_8463);
nor U9606 (N_9606,N_8019,N_8168);
xnor U9607 (N_9607,N_8788,N_8177);
and U9608 (N_9608,N_8394,N_8393);
and U9609 (N_9609,N_8409,N_8014);
or U9610 (N_9610,N_8565,N_8243);
and U9611 (N_9611,N_8265,N_8247);
or U9612 (N_9612,N_8718,N_8032);
xor U9613 (N_9613,N_8466,N_8392);
or U9614 (N_9614,N_8187,N_8197);
xor U9615 (N_9615,N_8133,N_8122);
nand U9616 (N_9616,N_8078,N_8981);
xnor U9617 (N_9617,N_8352,N_8796);
and U9618 (N_9618,N_8247,N_8489);
nand U9619 (N_9619,N_8903,N_8404);
or U9620 (N_9620,N_8588,N_8477);
nor U9621 (N_9621,N_8778,N_8861);
and U9622 (N_9622,N_8437,N_8678);
and U9623 (N_9623,N_8612,N_8808);
nand U9624 (N_9624,N_8046,N_8630);
and U9625 (N_9625,N_8306,N_8114);
or U9626 (N_9626,N_8718,N_8324);
and U9627 (N_9627,N_8552,N_8112);
nand U9628 (N_9628,N_8815,N_8257);
and U9629 (N_9629,N_8315,N_8516);
nor U9630 (N_9630,N_8982,N_8361);
or U9631 (N_9631,N_8245,N_8935);
nor U9632 (N_9632,N_8392,N_8936);
or U9633 (N_9633,N_8694,N_8019);
and U9634 (N_9634,N_8189,N_8283);
and U9635 (N_9635,N_8203,N_8757);
or U9636 (N_9636,N_8225,N_8135);
xor U9637 (N_9637,N_8492,N_8429);
nor U9638 (N_9638,N_8064,N_8466);
and U9639 (N_9639,N_8127,N_8056);
nand U9640 (N_9640,N_8395,N_8280);
nor U9641 (N_9641,N_8978,N_8347);
nand U9642 (N_9642,N_8131,N_8987);
nor U9643 (N_9643,N_8366,N_8948);
nand U9644 (N_9644,N_8898,N_8008);
and U9645 (N_9645,N_8042,N_8129);
nand U9646 (N_9646,N_8167,N_8490);
nor U9647 (N_9647,N_8794,N_8285);
nor U9648 (N_9648,N_8276,N_8941);
nor U9649 (N_9649,N_8856,N_8452);
xor U9650 (N_9650,N_8353,N_8064);
and U9651 (N_9651,N_8871,N_8022);
nor U9652 (N_9652,N_8100,N_8217);
or U9653 (N_9653,N_8460,N_8630);
nor U9654 (N_9654,N_8607,N_8006);
and U9655 (N_9655,N_8954,N_8808);
and U9656 (N_9656,N_8742,N_8919);
xnor U9657 (N_9657,N_8854,N_8388);
nor U9658 (N_9658,N_8832,N_8019);
nor U9659 (N_9659,N_8816,N_8124);
nand U9660 (N_9660,N_8683,N_8858);
nor U9661 (N_9661,N_8244,N_8064);
and U9662 (N_9662,N_8106,N_8578);
xor U9663 (N_9663,N_8471,N_8494);
nor U9664 (N_9664,N_8580,N_8703);
nor U9665 (N_9665,N_8044,N_8208);
xor U9666 (N_9666,N_8621,N_8432);
nand U9667 (N_9667,N_8288,N_8021);
nand U9668 (N_9668,N_8413,N_8247);
nor U9669 (N_9669,N_8092,N_8881);
nor U9670 (N_9670,N_8090,N_8738);
nor U9671 (N_9671,N_8010,N_8876);
nor U9672 (N_9672,N_8077,N_8280);
or U9673 (N_9673,N_8318,N_8395);
and U9674 (N_9674,N_8519,N_8564);
xor U9675 (N_9675,N_8846,N_8899);
nand U9676 (N_9676,N_8656,N_8182);
or U9677 (N_9677,N_8357,N_8154);
nand U9678 (N_9678,N_8470,N_8444);
nor U9679 (N_9679,N_8442,N_8434);
nor U9680 (N_9680,N_8798,N_8221);
or U9681 (N_9681,N_8738,N_8570);
and U9682 (N_9682,N_8190,N_8202);
nor U9683 (N_9683,N_8815,N_8767);
or U9684 (N_9684,N_8350,N_8565);
or U9685 (N_9685,N_8317,N_8554);
nor U9686 (N_9686,N_8458,N_8133);
and U9687 (N_9687,N_8411,N_8742);
and U9688 (N_9688,N_8117,N_8439);
or U9689 (N_9689,N_8422,N_8831);
or U9690 (N_9690,N_8488,N_8332);
and U9691 (N_9691,N_8724,N_8807);
and U9692 (N_9692,N_8165,N_8981);
nand U9693 (N_9693,N_8630,N_8299);
nor U9694 (N_9694,N_8529,N_8577);
xor U9695 (N_9695,N_8240,N_8299);
or U9696 (N_9696,N_8478,N_8960);
nand U9697 (N_9697,N_8781,N_8214);
or U9698 (N_9698,N_8978,N_8859);
nand U9699 (N_9699,N_8753,N_8742);
and U9700 (N_9700,N_8111,N_8408);
and U9701 (N_9701,N_8889,N_8043);
nand U9702 (N_9702,N_8887,N_8762);
xor U9703 (N_9703,N_8841,N_8628);
and U9704 (N_9704,N_8062,N_8298);
nor U9705 (N_9705,N_8072,N_8502);
xor U9706 (N_9706,N_8685,N_8261);
and U9707 (N_9707,N_8290,N_8757);
nor U9708 (N_9708,N_8185,N_8448);
and U9709 (N_9709,N_8355,N_8719);
nor U9710 (N_9710,N_8330,N_8507);
xor U9711 (N_9711,N_8380,N_8221);
and U9712 (N_9712,N_8827,N_8330);
nand U9713 (N_9713,N_8307,N_8833);
and U9714 (N_9714,N_8944,N_8052);
nand U9715 (N_9715,N_8669,N_8513);
or U9716 (N_9716,N_8221,N_8112);
or U9717 (N_9717,N_8605,N_8091);
and U9718 (N_9718,N_8964,N_8613);
and U9719 (N_9719,N_8826,N_8416);
nand U9720 (N_9720,N_8272,N_8460);
nor U9721 (N_9721,N_8211,N_8226);
or U9722 (N_9722,N_8654,N_8963);
or U9723 (N_9723,N_8430,N_8601);
and U9724 (N_9724,N_8055,N_8808);
nor U9725 (N_9725,N_8397,N_8840);
nand U9726 (N_9726,N_8176,N_8796);
nor U9727 (N_9727,N_8471,N_8486);
xor U9728 (N_9728,N_8859,N_8514);
nand U9729 (N_9729,N_8132,N_8655);
nor U9730 (N_9730,N_8467,N_8050);
xnor U9731 (N_9731,N_8157,N_8704);
xor U9732 (N_9732,N_8620,N_8003);
nand U9733 (N_9733,N_8041,N_8792);
and U9734 (N_9734,N_8875,N_8832);
or U9735 (N_9735,N_8233,N_8534);
nand U9736 (N_9736,N_8684,N_8049);
nor U9737 (N_9737,N_8251,N_8215);
nor U9738 (N_9738,N_8342,N_8203);
and U9739 (N_9739,N_8400,N_8175);
or U9740 (N_9740,N_8802,N_8535);
nand U9741 (N_9741,N_8581,N_8951);
nor U9742 (N_9742,N_8363,N_8522);
nand U9743 (N_9743,N_8843,N_8352);
nand U9744 (N_9744,N_8310,N_8355);
nor U9745 (N_9745,N_8402,N_8983);
or U9746 (N_9746,N_8071,N_8241);
nand U9747 (N_9747,N_8786,N_8818);
nor U9748 (N_9748,N_8241,N_8008);
or U9749 (N_9749,N_8129,N_8648);
nor U9750 (N_9750,N_8898,N_8453);
or U9751 (N_9751,N_8118,N_8425);
nand U9752 (N_9752,N_8562,N_8302);
nand U9753 (N_9753,N_8606,N_8228);
or U9754 (N_9754,N_8822,N_8103);
xnor U9755 (N_9755,N_8076,N_8788);
xnor U9756 (N_9756,N_8121,N_8051);
and U9757 (N_9757,N_8286,N_8942);
nand U9758 (N_9758,N_8962,N_8833);
nand U9759 (N_9759,N_8091,N_8581);
or U9760 (N_9760,N_8717,N_8976);
xnor U9761 (N_9761,N_8512,N_8171);
or U9762 (N_9762,N_8798,N_8860);
or U9763 (N_9763,N_8050,N_8771);
and U9764 (N_9764,N_8513,N_8349);
nor U9765 (N_9765,N_8560,N_8603);
nand U9766 (N_9766,N_8531,N_8366);
nand U9767 (N_9767,N_8339,N_8315);
and U9768 (N_9768,N_8667,N_8092);
and U9769 (N_9769,N_8926,N_8353);
or U9770 (N_9770,N_8843,N_8379);
and U9771 (N_9771,N_8082,N_8455);
nor U9772 (N_9772,N_8723,N_8898);
and U9773 (N_9773,N_8937,N_8854);
xnor U9774 (N_9774,N_8775,N_8892);
nand U9775 (N_9775,N_8265,N_8436);
nor U9776 (N_9776,N_8863,N_8583);
nand U9777 (N_9777,N_8755,N_8314);
xnor U9778 (N_9778,N_8302,N_8601);
nand U9779 (N_9779,N_8824,N_8015);
nand U9780 (N_9780,N_8684,N_8921);
and U9781 (N_9781,N_8754,N_8599);
xor U9782 (N_9782,N_8829,N_8460);
and U9783 (N_9783,N_8901,N_8768);
nor U9784 (N_9784,N_8663,N_8668);
and U9785 (N_9785,N_8647,N_8810);
nand U9786 (N_9786,N_8504,N_8250);
nand U9787 (N_9787,N_8559,N_8164);
nor U9788 (N_9788,N_8261,N_8232);
nand U9789 (N_9789,N_8858,N_8931);
or U9790 (N_9790,N_8089,N_8218);
nand U9791 (N_9791,N_8370,N_8168);
or U9792 (N_9792,N_8258,N_8528);
nor U9793 (N_9793,N_8267,N_8290);
or U9794 (N_9794,N_8502,N_8775);
and U9795 (N_9795,N_8001,N_8027);
nand U9796 (N_9796,N_8577,N_8885);
or U9797 (N_9797,N_8581,N_8834);
and U9798 (N_9798,N_8745,N_8203);
and U9799 (N_9799,N_8597,N_8741);
xor U9800 (N_9800,N_8321,N_8934);
and U9801 (N_9801,N_8508,N_8610);
xnor U9802 (N_9802,N_8126,N_8296);
xor U9803 (N_9803,N_8335,N_8825);
nand U9804 (N_9804,N_8613,N_8334);
nand U9805 (N_9805,N_8269,N_8523);
and U9806 (N_9806,N_8633,N_8956);
nand U9807 (N_9807,N_8816,N_8791);
nor U9808 (N_9808,N_8490,N_8747);
or U9809 (N_9809,N_8532,N_8059);
xnor U9810 (N_9810,N_8950,N_8518);
and U9811 (N_9811,N_8410,N_8188);
and U9812 (N_9812,N_8316,N_8075);
and U9813 (N_9813,N_8698,N_8204);
nor U9814 (N_9814,N_8248,N_8189);
nor U9815 (N_9815,N_8893,N_8711);
or U9816 (N_9816,N_8696,N_8541);
xnor U9817 (N_9817,N_8863,N_8062);
nand U9818 (N_9818,N_8822,N_8991);
or U9819 (N_9819,N_8470,N_8049);
nor U9820 (N_9820,N_8926,N_8735);
xor U9821 (N_9821,N_8377,N_8498);
or U9822 (N_9822,N_8123,N_8261);
and U9823 (N_9823,N_8425,N_8095);
or U9824 (N_9824,N_8598,N_8817);
nor U9825 (N_9825,N_8969,N_8304);
nand U9826 (N_9826,N_8561,N_8379);
and U9827 (N_9827,N_8031,N_8029);
or U9828 (N_9828,N_8275,N_8689);
nand U9829 (N_9829,N_8330,N_8832);
nor U9830 (N_9830,N_8882,N_8702);
nor U9831 (N_9831,N_8900,N_8212);
and U9832 (N_9832,N_8081,N_8385);
nand U9833 (N_9833,N_8830,N_8658);
nor U9834 (N_9834,N_8199,N_8451);
xor U9835 (N_9835,N_8868,N_8681);
nor U9836 (N_9836,N_8834,N_8782);
or U9837 (N_9837,N_8756,N_8191);
nor U9838 (N_9838,N_8554,N_8250);
or U9839 (N_9839,N_8917,N_8743);
nor U9840 (N_9840,N_8832,N_8590);
nor U9841 (N_9841,N_8758,N_8375);
or U9842 (N_9842,N_8651,N_8932);
nor U9843 (N_9843,N_8369,N_8195);
nor U9844 (N_9844,N_8088,N_8134);
nand U9845 (N_9845,N_8214,N_8682);
nor U9846 (N_9846,N_8097,N_8769);
and U9847 (N_9847,N_8719,N_8800);
and U9848 (N_9848,N_8434,N_8154);
nor U9849 (N_9849,N_8718,N_8609);
nor U9850 (N_9850,N_8181,N_8282);
nand U9851 (N_9851,N_8807,N_8887);
and U9852 (N_9852,N_8296,N_8180);
or U9853 (N_9853,N_8588,N_8170);
nand U9854 (N_9854,N_8774,N_8244);
nor U9855 (N_9855,N_8663,N_8904);
nor U9856 (N_9856,N_8749,N_8351);
or U9857 (N_9857,N_8061,N_8907);
nand U9858 (N_9858,N_8289,N_8908);
nor U9859 (N_9859,N_8518,N_8010);
nor U9860 (N_9860,N_8061,N_8615);
nand U9861 (N_9861,N_8610,N_8309);
xnor U9862 (N_9862,N_8991,N_8398);
nand U9863 (N_9863,N_8514,N_8665);
and U9864 (N_9864,N_8668,N_8870);
or U9865 (N_9865,N_8045,N_8337);
nand U9866 (N_9866,N_8977,N_8139);
nor U9867 (N_9867,N_8689,N_8727);
nor U9868 (N_9868,N_8830,N_8798);
and U9869 (N_9869,N_8838,N_8006);
nand U9870 (N_9870,N_8130,N_8273);
xor U9871 (N_9871,N_8668,N_8333);
and U9872 (N_9872,N_8100,N_8916);
or U9873 (N_9873,N_8530,N_8999);
and U9874 (N_9874,N_8672,N_8092);
nand U9875 (N_9875,N_8399,N_8686);
and U9876 (N_9876,N_8336,N_8391);
and U9877 (N_9877,N_8504,N_8874);
or U9878 (N_9878,N_8689,N_8728);
and U9879 (N_9879,N_8200,N_8540);
or U9880 (N_9880,N_8246,N_8392);
or U9881 (N_9881,N_8108,N_8820);
and U9882 (N_9882,N_8375,N_8155);
or U9883 (N_9883,N_8856,N_8199);
or U9884 (N_9884,N_8345,N_8720);
or U9885 (N_9885,N_8965,N_8532);
nor U9886 (N_9886,N_8757,N_8053);
nor U9887 (N_9887,N_8147,N_8068);
nand U9888 (N_9888,N_8396,N_8871);
or U9889 (N_9889,N_8409,N_8682);
nand U9890 (N_9890,N_8002,N_8440);
and U9891 (N_9891,N_8397,N_8100);
or U9892 (N_9892,N_8853,N_8511);
nor U9893 (N_9893,N_8872,N_8425);
nand U9894 (N_9894,N_8103,N_8511);
or U9895 (N_9895,N_8448,N_8637);
nand U9896 (N_9896,N_8924,N_8673);
nand U9897 (N_9897,N_8910,N_8586);
nand U9898 (N_9898,N_8235,N_8758);
or U9899 (N_9899,N_8993,N_8318);
or U9900 (N_9900,N_8186,N_8785);
xnor U9901 (N_9901,N_8821,N_8680);
nand U9902 (N_9902,N_8438,N_8486);
nand U9903 (N_9903,N_8864,N_8001);
nor U9904 (N_9904,N_8929,N_8410);
nand U9905 (N_9905,N_8934,N_8420);
nor U9906 (N_9906,N_8880,N_8773);
or U9907 (N_9907,N_8325,N_8734);
nand U9908 (N_9908,N_8485,N_8360);
or U9909 (N_9909,N_8759,N_8370);
and U9910 (N_9910,N_8211,N_8822);
nor U9911 (N_9911,N_8769,N_8763);
or U9912 (N_9912,N_8636,N_8704);
or U9913 (N_9913,N_8525,N_8756);
nor U9914 (N_9914,N_8143,N_8803);
and U9915 (N_9915,N_8741,N_8348);
nand U9916 (N_9916,N_8135,N_8056);
and U9917 (N_9917,N_8427,N_8662);
nand U9918 (N_9918,N_8785,N_8478);
nand U9919 (N_9919,N_8248,N_8242);
nand U9920 (N_9920,N_8572,N_8675);
and U9921 (N_9921,N_8560,N_8302);
and U9922 (N_9922,N_8516,N_8008);
and U9923 (N_9923,N_8496,N_8783);
nand U9924 (N_9924,N_8625,N_8415);
and U9925 (N_9925,N_8776,N_8764);
and U9926 (N_9926,N_8689,N_8583);
nor U9927 (N_9927,N_8750,N_8358);
and U9928 (N_9928,N_8174,N_8497);
and U9929 (N_9929,N_8767,N_8704);
or U9930 (N_9930,N_8608,N_8233);
xnor U9931 (N_9931,N_8296,N_8713);
and U9932 (N_9932,N_8413,N_8192);
and U9933 (N_9933,N_8481,N_8379);
and U9934 (N_9934,N_8301,N_8159);
nand U9935 (N_9935,N_8481,N_8563);
nand U9936 (N_9936,N_8046,N_8342);
xor U9937 (N_9937,N_8532,N_8901);
or U9938 (N_9938,N_8607,N_8804);
and U9939 (N_9939,N_8490,N_8042);
xnor U9940 (N_9940,N_8216,N_8301);
and U9941 (N_9941,N_8378,N_8212);
nor U9942 (N_9942,N_8589,N_8025);
xnor U9943 (N_9943,N_8639,N_8716);
xnor U9944 (N_9944,N_8788,N_8988);
nor U9945 (N_9945,N_8951,N_8404);
nand U9946 (N_9946,N_8974,N_8151);
nor U9947 (N_9947,N_8209,N_8515);
nand U9948 (N_9948,N_8528,N_8524);
and U9949 (N_9949,N_8385,N_8095);
xnor U9950 (N_9950,N_8428,N_8985);
and U9951 (N_9951,N_8197,N_8004);
nor U9952 (N_9952,N_8059,N_8666);
xnor U9953 (N_9953,N_8221,N_8192);
and U9954 (N_9954,N_8390,N_8143);
nor U9955 (N_9955,N_8765,N_8507);
xnor U9956 (N_9956,N_8256,N_8633);
nor U9957 (N_9957,N_8362,N_8721);
nand U9958 (N_9958,N_8846,N_8535);
nor U9959 (N_9959,N_8303,N_8018);
and U9960 (N_9960,N_8644,N_8839);
nand U9961 (N_9961,N_8110,N_8116);
and U9962 (N_9962,N_8241,N_8151);
or U9963 (N_9963,N_8736,N_8200);
or U9964 (N_9964,N_8598,N_8403);
or U9965 (N_9965,N_8568,N_8505);
nor U9966 (N_9966,N_8326,N_8474);
xor U9967 (N_9967,N_8094,N_8157);
nand U9968 (N_9968,N_8873,N_8920);
nand U9969 (N_9969,N_8006,N_8082);
xor U9970 (N_9970,N_8563,N_8268);
or U9971 (N_9971,N_8826,N_8776);
and U9972 (N_9972,N_8603,N_8166);
xor U9973 (N_9973,N_8891,N_8692);
nor U9974 (N_9974,N_8022,N_8670);
nand U9975 (N_9975,N_8405,N_8701);
xnor U9976 (N_9976,N_8693,N_8952);
or U9977 (N_9977,N_8953,N_8267);
nor U9978 (N_9978,N_8208,N_8270);
or U9979 (N_9979,N_8094,N_8816);
and U9980 (N_9980,N_8218,N_8197);
or U9981 (N_9981,N_8952,N_8461);
nor U9982 (N_9982,N_8267,N_8019);
nor U9983 (N_9983,N_8340,N_8475);
nand U9984 (N_9984,N_8949,N_8924);
nor U9985 (N_9985,N_8693,N_8461);
and U9986 (N_9986,N_8784,N_8124);
nand U9987 (N_9987,N_8778,N_8439);
nand U9988 (N_9988,N_8971,N_8963);
nand U9989 (N_9989,N_8230,N_8430);
and U9990 (N_9990,N_8235,N_8678);
and U9991 (N_9991,N_8755,N_8568);
or U9992 (N_9992,N_8423,N_8327);
or U9993 (N_9993,N_8049,N_8963);
nand U9994 (N_9994,N_8670,N_8693);
or U9995 (N_9995,N_8245,N_8997);
nand U9996 (N_9996,N_8803,N_8790);
and U9997 (N_9997,N_8707,N_8419);
and U9998 (N_9998,N_8604,N_8359);
nor U9999 (N_9999,N_8387,N_8030);
nand U10000 (N_10000,N_9673,N_9485);
nor U10001 (N_10001,N_9581,N_9349);
or U10002 (N_10002,N_9802,N_9133);
nand U10003 (N_10003,N_9708,N_9936);
and U10004 (N_10004,N_9305,N_9624);
and U10005 (N_10005,N_9403,N_9049);
xor U10006 (N_10006,N_9202,N_9979);
or U10007 (N_10007,N_9442,N_9881);
nor U10008 (N_10008,N_9385,N_9353);
nor U10009 (N_10009,N_9718,N_9505);
nand U10010 (N_10010,N_9509,N_9529);
nand U10011 (N_10011,N_9228,N_9625);
nor U10012 (N_10012,N_9914,N_9953);
nand U10013 (N_10013,N_9332,N_9294);
or U10014 (N_10014,N_9768,N_9942);
nand U10015 (N_10015,N_9514,N_9666);
and U10016 (N_10016,N_9838,N_9033);
nor U10017 (N_10017,N_9097,N_9705);
nor U10018 (N_10018,N_9498,N_9905);
nor U10019 (N_10019,N_9947,N_9085);
nor U10020 (N_10020,N_9820,N_9396);
nor U10021 (N_10021,N_9036,N_9676);
or U10022 (N_10022,N_9343,N_9408);
or U10023 (N_10023,N_9525,N_9751);
xor U10024 (N_10024,N_9621,N_9369);
nor U10025 (N_10025,N_9523,N_9703);
nand U10026 (N_10026,N_9064,N_9288);
and U10027 (N_10027,N_9100,N_9304);
or U10028 (N_10028,N_9563,N_9913);
nor U10029 (N_10029,N_9484,N_9561);
or U10030 (N_10030,N_9285,N_9730);
nor U10031 (N_10031,N_9334,N_9531);
nand U10032 (N_10032,N_9083,N_9140);
xnor U10033 (N_10033,N_9923,N_9930);
nor U10034 (N_10034,N_9082,N_9990);
and U10035 (N_10035,N_9207,N_9231);
or U10036 (N_10036,N_9185,N_9495);
nor U10037 (N_10037,N_9190,N_9964);
and U10038 (N_10038,N_9599,N_9892);
nand U10039 (N_10039,N_9093,N_9917);
and U10040 (N_10040,N_9131,N_9874);
nor U10041 (N_10041,N_9926,N_9585);
and U10042 (N_10042,N_9669,N_9073);
or U10043 (N_10043,N_9181,N_9216);
xnor U10044 (N_10044,N_9389,N_9859);
nor U10045 (N_10045,N_9124,N_9754);
nand U10046 (N_10046,N_9086,N_9316);
xor U10047 (N_10047,N_9595,N_9588);
xor U10048 (N_10048,N_9478,N_9031);
or U10049 (N_10049,N_9088,N_9213);
nand U10050 (N_10050,N_9989,N_9186);
and U10051 (N_10051,N_9032,N_9924);
or U10052 (N_10052,N_9507,N_9861);
nor U10053 (N_10053,N_9402,N_9192);
and U10054 (N_10054,N_9643,N_9896);
or U10055 (N_10055,N_9569,N_9035);
xnor U10056 (N_10056,N_9797,N_9863);
and U10057 (N_10057,N_9919,N_9842);
nand U10058 (N_10058,N_9274,N_9125);
xnor U10059 (N_10059,N_9998,N_9452);
and U10060 (N_10060,N_9882,N_9799);
nor U10061 (N_10061,N_9240,N_9806);
and U10062 (N_10062,N_9577,N_9114);
or U10063 (N_10063,N_9620,N_9675);
and U10064 (N_10064,N_9107,N_9096);
or U10065 (N_10065,N_9571,N_9547);
xor U10066 (N_10066,N_9262,N_9184);
and U10067 (N_10067,N_9350,N_9464);
and U10068 (N_10068,N_9215,N_9511);
nor U10069 (N_10069,N_9938,N_9579);
nand U10070 (N_10070,N_9263,N_9432);
nor U10071 (N_10071,N_9732,N_9607);
nor U10072 (N_10072,N_9287,N_9250);
nor U10073 (N_10073,N_9441,N_9182);
or U10074 (N_10074,N_9986,N_9677);
nand U10075 (N_10075,N_9277,N_9612);
xor U10076 (N_10076,N_9940,N_9494);
nor U10077 (N_10077,N_9671,N_9860);
or U10078 (N_10078,N_9273,N_9741);
nand U10079 (N_10079,N_9771,N_9243);
and U10080 (N_10080,N_9999,N_9760);
and U10081 (N_10081,N_9841,N_9183);
and U10082 (N_10082,N_9050,N_9428);
nor U10083 (N_10083,N_9493,N_9283);
nand U10084 (N_10084,N_9380,N_9707);
and U10085 (N_10085,N_9112,N_9003);
or U10086 (N_10086,N_9617,N_9413);
nand U10087 (N_10087,N_9309,N_9813);
nand U10088 (N_10088,N_9312,N_9709);
or U10089 (N_10089,N_9686,N_9536);
and U10090 (N_10090,N_9632,N_9412);
xor U10091 (N_10091,N_9743,N_9652);
nand U10092 (N_10092,N_9174,N_9555);
or U10093 (N_10093,N_9013,N_9598);
and U10094 (N_10094,N_9694,N_9382);
or U10095 (N_10095,N_9067,N_9904);
nor U10096 (N_10096,N_9356,N_9483);
and U10097 (N_10097,N_9526,N_9266);
and U10098 (N_10098,N_9368,N_9109);
or U10099 (N_10099,N_9846,N_9340);
and U10100 (N_10100,N_9293,N_9487);
nand U10101 (N_10101,N_9360,N_9706);
and U10102 (N_10102,N_9257,N_9715);
nor U10103 (N_10103,N_9341,N_9435);
nand U10104 (N_10104,N_9911,N_9681);
nand U10105 (N_10105,N_9609,N_9546);
nand U10106 (N_10106,N_9766,N_9450);
nor U10107 (N_10107,N_9533,N_9918);
nand U10108 (N_10108,N_9299,N_9142);
or U10109 (N_10109,N_9761,N_9091);
nor U10110 (N_10110,N_9858,N_9967);
nor U10111 (N_10111,N_9866,N_9572);
nand U10112 (N_10112,N_9395,N_9587);
or U10113 (N_10113,N_9017,N_9653);
xor U10114 (N_10114,N_9254,N_9795);
nand U10115 (N_10115,N_9994,N_9138);
and U10116 (N_10116,N_9524,N_9455);
nor U10117 (N_10117,N_9251,N_9638);
and U10118 (N_10118,N_9649,N_9727);
and U10119 (N_10119,N_9935,N_9249);
nor U10120 (N_10120,N_9749,N_9463);
nand U10121 (N_10121,N_9027,N_9451);
nand U10122 (N_10122,N_9233,N_9070);
and U10123 (N_10123,N_9225,N_9034);
nor U10124 (N_10124,N_9414,N_9252);
xnor U10125 (N_10125,N_9622,N_9457);
xnor U10126 (N_10126,N_9674,N_9672);
nor U10127 (N_10127,N_9748,N_9634);
or U10128 (N_10128,N_9223,N_9246);
nor U10129 (N_10129,N_9869,N_9370);
nand U10130 (N_10130,N_9982,N_9823);
and U10131 (N_10131,N_9684,N_9603);
and U10132 (N_10132,N_9218,N_9129);
or U10133 (N_10133,N_9245,N_9520);
nand U10134 (N_10134,N_9700,N_9591);
nor U10135 (N_10135,N_9566,N_9358);
and U10136 (N_10136,N_9220,N_9880);
or U10137 (N_10137,N_9884,N_9016);
and U10138 (N_10138,N_9560,N_9470);
or U10139 (N_10139,N_9416,N_9697);
and U10140 (N_10140,N_9026,N_9302);
and U10141 (N_10141,N_9835,N_9122);
and U10142 (N_10142,N_9168,N_9055);
and U10143 (N_10143,N_9264,N_9196);
or U10144 (N_10144,N_9957,N_9152);
nand U10145 (N_10145,N_9557,N_9628);
nand U10146 (N_10146,N_9508,N_9044);
and U10147 (N_10147,N_9646,N_9059);
or U10148 (N_10148,N_9871,N_9931);
xnor U10149 (N_10149,N_9271,N_9499);
or U10150 (N_10150,N_9038,N_9636);
or U10151 (N_10151,N_9807,N_9012);
nand U10152 (N_10152,N_9849,N_9039);
nand U10153 (N_10153,N_9770,N_9386);
nand U10154 (N_10154,N_9907,N_9401);
xor U10155 (N_10155,N_9641,N_9651);
xnor U10156 (N_10156,N_9654,N_9565);
nor U10157 (N_10157,N_9278,N_9247);
or U10158 (N_10158,N_9980,N_9545);
nor U10159 (N_10159,N_9750,N_9532);
nand U10160 (N_10160,N_9147,N_9699);
nor U10161 (N_10161,N_9659,N_9118);
nor U10162 (N_10162,N_9567,N_9199);
nand U10163 (N_10163,N_9586,N_9438);
xnor U10164 (N_10164,N_9375,N_9205);
and U10165 (N_10165,N_9130,N_9388);
or U10166 (N_10166,N_9968,N_9877);
nor U10167 (N_10167,N_9418,N_9738);
xor U10168 (N_10168,N_9217,N_9374);
or U10169 (N_10169,N_9279,N_9976);
nor U10170 (N_10170,N_9790,N_9993);
xor U10171 (N_10171,N_9972,N_9430);
xor U10172 (N_10172,N_9746,N_9724);
nand U10173 (N_10173,N_9466,N_9095);
and U10174 (N_10174,N_9791,N_9721);
xnor U10175 (N_10175,N_9387,N_9134);
nor U10176 (N_10176,N_9966,N_9977);
nand U10177 (N_10177,N_9851,N_9803);
or U10178 (N_10178,N_9473,N_9680);
nor U10179 (N_10179,N_9108,N_9132);
or U10180 (N_10180,N_9420,N_9324);
xnor U10181 (N_10181,N_9745,N_9178);
nand U10182 (N_10182,N_9594,N_9175);
xnor U10183 (N_10183,N_9153,N_9757);
nand U10184 (N_10184,N_9145,N_9203);
nor U10185 (N_10185,N_9023,N_9297);
and U10186 (N_10186,N_9166,N_9090);
xor U10187 (N_10187,N_9482,N_9501);
and U10188 (N_10188,N_9137,N_9020);
or U10189 (N_10189,N_9883,N_9782);
xor U10190 (N_10190,N_9048,N_9978);
and U10191 (N_10191,N_9206,N_9394);
and U10192 (N_10192,N_9837,N_9729);
and U10193 (N_10193,N_9965,N_9845);
xnor U10194 (N_10194,N_9758,N_9519);
nand U10195 (N_10195,N_9656,N_9764);
nand U10196 (N_10196,N_9901,N_9822);
and U10197 (N_10197,N_9080,N_9028);
xor U10198 (N_10198,N_9698,N_9135);
and U10199 (N_10199,N_9322,N_9633);
or U10200 (N_10200,N_9510,N_9513);
or U10201 (N_10201,N_9261,N_9619);
and U10202 (N_10202,N_9069,N_9679);
and U10203 (N_10203,N_9197,N_9504);
nand U10204 (N_10204,N_9150,N_9308);
xnor U10205 (N_10205,N_9722,N_9406);
nor U10206 (N_10206,N_9248,N_9253);
xnor U10207 (N_10207,N_9736,N_9188);
xnor U10208 (N_10208,N_9425,N_9005);
and U10209 (N_10209,N_9830,N_9479);
and U10210 (N_10210,N_9945,N_9068);
nor U10211 (N_10211,N_9126,N_9007);
xor U10212 (N_10212,N_9956,N_9265);
or U10213 (N_10213,N_9839,N_9713);
or U10214 (N_10214,N_9436,N_9241);
nor U10215 (N_10215,N_9065,N_9584);
and U10216 (N_10216,N_9958,N_9983);
nor U10217 (N_10217,N_9827,N_9981);
or U10218 (N_10218,N_9787,N_9578);
nor U10219 (N_10219,N_9204,N_9716);
or U10220 (N_10220,N_9548,N_9336);
and U10221 (N_10221,N_9201,N_9717);
nor U10222 (N_10222,N_9025,N_9276);
nand U10223 (N_10223,N_9422,N_9480);
nand U10224 (N_10224,N_9844,N_9163);
or U10225 (N_10225,N_9431,N_9735);
or U10226 (N_10226,N_9377,N_9310);
nand U10227 (N_10227,N_9991,N_9339);
or U10228 (N_10228,N_9921,N_9879);
nand U10229 (N_10229,N_9209,N_9602);
and U10230 (N_10230,N_9384,N_9773);
or U10231 (N_10231,N_9345,N_9973);
and U10232 (N_10232,N_9922,N_9057);
nand U10233 (N_10233,N_9361,N_9856);
nand U10234 (N_10234,N_9221,N_9933);
and U10235 (N_10235,N_9392,N_9898);
and U10236 (N_10236,N_9793,N_9191);
nand U10237 (N_10237,N_9326,N_9194);
nor U10238 (N_10238,N_9852,N_9502);
xor U10239 (N_10239,N_9331,N_9576);
and U10240 (N_10240,N_9895,N_9066);
or U10241 (N_10241,N_9834,N_9954);
nor U10242 (N_10242,N_9959,N_9235);
nor U10243 (N_10243,N_9559,N_9600);
nor U10244 (N_10244,N_9714,N_9840);
and U10245 (N_10245,N_9267,N_9890);
and U10246 (N_10246,N_9497,N_9378);
nor U10247 (N_10247,N_9056,N_9614);
or U10248 (N_10248,N_9063,N_9338);
nand U10249 (N_10249,N_9992,N_9828);
or U10250 (N_10250,N_9164,N_9704);
and U10251 (N_10251,N_9290,N_9259);
xor U10252 (N_10252,N_9021,N_9342);
nor U10253 (N_10253,N_9885,N_9329);
nand U10254 (N_10254,N_9219,N_9029);
xor U10255 (N_10255,N_9516,N_9214);
nand U10256 (N_10256,N_9469,N_9540);
or U10257 (N_10257,N_9461,N_9444);
nand U10258 (N_10258,N_9702,N_9149);
nor U10259 (N_10259,N_9562,N_9521);
nor U10260 (N_10260,N_9593,N_9597);
and U10261 (N_10261,N_9465,N_9426);
and U10262 (N_10262,N_9106,N_9004);
nand U10263 (N_10263,N_9001,N_9535);
nand U10264 (N_10264,N_9755,N_9682);
or U10265 (N_10265,N_9291,N_9725);
and U10266 (N_10266,N_9237,N_9058);
xnor U10267 (N_10267,N_9988,N_9558);
or U10268 (N_10268,N_9503,N_9136);
or U10269 (N_10269,N_9117,N_9325);
xnor U10270 (N_10270,N_9024,N_9011);
nand U10271 (N_10271,N_9542,N_9330);
or U10272 (N_10272,N_9155,N_9071);
or U10273 (N_10273,N_9951,N_9631);
nor U10274 (N_10274,N_9037,N_9712);
xor U10275 (N_10275,N_9670,N_9543);
and U10276 (N_10276,N_9678,N_9928);
or U10277 (N_10277,N_9969,N_9658);
xor U10278 (N_10278,N_9886,N_9832);
and U10279 (N_10279,N_9417,N_9078);
nor U10280 (N_10280,N_9275,N_9492);
nand U10281 (N_10281,N_9644,N_9286);
and U10282 (N_10282,N_9995,N_9648);
or U10283 (N_10283,N_9788,N_9052);
or U10284 (N_10284,N_9177,N_9195);
nand U10285 (N_10285,N_9113,N_9333);
nor U10286 (N_10286,N_9517,N_9101);
nor U10287 (N_10287,N_9728,N_9045);
xnor U10288 (N_10288,N_9236,N_9808);
or U10289 (N_10289,N_9894,N_9857);
or U10290 (N_10290,N_9888,N_9355);
xor U10291 (N_10291,N_9047,N_9912);
nor U10292 (N_10292,N_9552,N_9512);
and U10293 (N_10293,N_9372,N_9475);
nor U10294 (N_10294,N_9317,N_9775);
nand U10295 (N_10295,N_9893,N_9847);
and U10296 (N_10296,N_9887,N_9723);
xor U10297 (N_10297,N_9015,N_9800);
nor U10298 (N_10298,N_9590,N_9637);
nor U10299 (N_10299,N_9371,N_9193);
nor U10300 (N_10300,N_9210,N_9159);
xnor U10301 (N_10301,N_9937,N_9635);
and U10302 (N_10302,N_9367,N_9903);
nor U10303 (N_10303,N_9689,N_9601);
xor U10304 (N_10304,N_9076,N_9925);
nand U10305 (N_10305,N_9061,N_9819);
and U10306 (N_10306,N_9315,N_9604);
xnor U10307 (N_10307,N_9810,N_9574);
and U10308 (N_10308,N_9087,N_9300);
or U10309 (N_10309,N_9962,N_9123);
and U10310 (N_10310,N_9351,N_9391);
nor U10311 (N_10311,N_9752,N_9929);
xnor U10312 (N_10312,N_9110,N_9891);
nand U10313 (N_10313,N_9971,N_9939);
or U10314 (N_10314,N_9415,N_9363);
or U10315 (N_10315,N_9655,N_9008);
nor U10316 (N_10316,N_9640,N_9941);
xnor U10317 (N_10317,N_9997,N_9102);
nand U10318 (N_10318,N_9139,N_9908);
nor U10319 (N_10319,N_9753,N_9870);
xnor U10320 (N_10320,N_9796,N_9379);
nor U10321 (N_10321,N_9701,N_9019);
nand U10322 (N_10322,N_9311,N_9961);
or U10323 (N_10323,N_9934,N_9344);
and U10324 (N_10324,N_9774,N_9270);
xor U10325 (N_10325,N_9948,N_9605);
nand U10326 (N_10326,N_9843,N_9824);
nand U10327 (N_10327,N_9833,N_9148);
nand U10328 (N_10328,N_9623,N_9060);
nor U10329 (N_10329,N_9429,N_9556);
nand U10330 (N_10330,N_9688,N_9411);
xor U10331 (N_10331,N_9295,N_9365);
and U10332 (N_10332,N_9121,N_9440);
nor U10333 (N_10333,N_9352,N_9439);
nand U10334 (N_10334,N_9878,N_9613);
nor U10335 (N_10335,N_9539,N_9410);
nor U10336 (N_10336,N_9281,N_9639);
nand U10337 (N_10337,N_9119,N_9282);
nor U10338 (N_10338,N_9811,N_9528);
and U10339 (N_10339,N_9167,N_9734);
or U10340 (N_10340,N_9608,N_9784);
nand U10341 (N_10341,N_9301,N_9272);
nor U10342 (N_10342,N_9779,N_9230);
nor U10343 (N_10343,N_9906,N_9875);
nor U10344 (N_10344,N_9496,N_9446);
nand U10345 (N_10345,N_9116,N_9224);
nor U10346 (N_10346,N_9872,N_9084);
nand U10347 (N_10347,N_9711,N_9018);
and U10348 (N_10348,N_9269,N_9002);
nor U10349 (N_10349,N_9260,N_9868);
nor U10350 (N_10350,N_9695,N_9647);
nand U10351 (N_10351,N_9081,N_9500);
nor U10352 (N_10352,N_9098,N_9792);
xor U10353 (N_10353,N_9160,N_9783);
nand U10354 (N_10354,N_9042,N_9474);
nor U10355 (N_10355,N_9865,N_9337);
nand U10356 (N_10356,N_9459,N_9970);
or U10357 (N_10357,N_9296,N_9335);
nor U10358 (N_10358,N_9685,N_9952);
nand U10359 (N_10359,N_9897,N_9383);
nor U10360 (N_10360,N_9229,N_9950);
nand U10361 (N_10361,N_9433,N_9234);
or U10362 (N_10362,N_9357,N_9393);
nand U10363 (N_10363,N_9850,N_9143);
xnor U10364 (N_10364,N_9550,N_9158);
nand U10365 (N_10365,N_9364,N_9815);
and U10366 (N_10366,N_9359,N_9902);
and U10367 (N_10367,N_9855,N_9876);
nand U10368 (N_10368,N_9161,N_9405);
or U10369 (N_10369,N_9362,N_9580);
nand U10370 (N_10370,N_9169,N_9915);
and U10371 (N_10371,N_9280,N_9772);
nor U10372 (N_10372,N_9289,N_9544);
and U10373 (N_10373,N_9105,N_9458);
nand U10374 (N_10374,N_9873,N_9006);
or U10375 (N_10375,N_9256,N_9814);
or U10376 (N_10376,N_9805,N_9780);
nand U10377 (N_10377,N_9541,N_9354);
nand U10378 (N_10378,N_9568,N_9984);
nand U10379 (N_10379,N_9051,N_9737);
or U10380 (N_10380,N_9974,N_9211);
xnor U10381 (N_10381,N_9212,N_9836);
nor U10382 (N_10382,N_9157,N_9477);
nand U10383 (N_10383,N_9258,N_9127);
or U10384 (N_10384,N_9404,N_9089);
nor U10385 (N_10385,N_9955,N_9156);
nand U10386 (N_10386,N_9443,N_9610);
or U10387 (N_10387,N_9592,N_9744);
nand U10388 (N_10388,N_9103,N_9400);
and U10389 (N_10389,N_9665,N_9319);
xor U10390 (N_10390,N_9927,N_9645);
nand U10391 (N_10391,N_9996,N_9664);
nor U10392 (N_10392,N_9151,N_9407);
nand U10393 (N_10393,N_9486,N_9762);
and U10394 (N_10394,N_9128,N_9767);
and U10395 (N_10395,N_9009,N_9573);
or U10396 (N_10396,N_9825,N_9094);
nand U10397 (N_10397,N_9074,N_9611);
and U10398 (N_10398,N_9693,N_9522);
and U10399 (N_10399,N_9570,N_9077);
nor U10400 (N_10400,N_9348,N_9899);
nor U10401 (N_10401,N_9690,N_9471);
nor U10402 (N_10402,N_9226,N_9687);
nor U10403 (N_10403,N_9255,N_9314);
nor U10404 (N_10404,N_9376,N_9120);
or U10405 (N_10405,N_9818,N_9650);
or U10406 (N_10406,N_9238,N_9900);
nand U10407 (N_10407,N_9176,N_9014);
nor U10408 (N_10408,N_9423,N_9642);
or U10409 (N_10409,N_9946,N_9030);
nand U10410 (N_10410,N_9826,N_9072);
nor U10411 (N_10411,N_9985,N_9812);
and U10412 (N_10412,N_9115,N_9615);
nand U10413 (N_10413,N_9794,N_9589);
nor U10414 (N_10414,N_9853,N_9862);
and U10415 (N_10415,N_9583,N_9447);
nand U10416 (N_10416,N_9848,N_9733);
nand U10417 (N_10417,N_9949,N_9437);
and U10418 (N_10418,N_9710,N_9831);
or U10419 (N_10419,N_9975,N_9920);
nand U10420 (N_10420,N_9373,N_9909);
and U10421 (N_10421,N_9244,N_9816);
nor U10422 (N_10422,N_9551,N_9538);
nand U10423 (N_10423,N_9777,N_9456);
xnor U10424 (N_10424,N_9141,N_9165);
nand U10425 (N_10425,N_9381,N_9798);
and U10426 (N_10426,N_9910,N_9667);
nor U10427 (N_10427,N_9756,N_9144);
nand U10428 (N_10428,N_9944,N_9306);
or U10429 (N_10429,N_9448,N_9720);
nand U10430 (N_10430,N_9731,N_9769);
nand U10431 (N_10431,N_9663,N_9419);
and U10432 (N_10432,N_9691,N_9427);
nor U10433 (N_10433,N_9683,N_9173);
nand U10434 (N_10434,N_9747,N_9445);
or U10435 (N_10435,N_9696,N_9328);
nor U10436 (N_10436,N_9227,N_9726);
nand U10437 (N_10437,N_9434,N_9170);
nand U10438 (N_10438,N_9618,N_9453);
xnor U10439 (N_10439,N_9318,N_9489);
and U10440 (N_10440,N_9657,N_9307);
or U10441 (N_10441,N_9390,N_9763);
xnor U10442 (N_10442,N_9321,N_9022);
or U10443 (N_10443,N_9960,N_9399);
xor U10444 (N_10444,N_9104,N_9626);
nor U10445 (N_10445,N_9943,N_9629);
nand U10446 (N_10446,N_9963,N_9462);
nor U10447 (N_10447,N_9467,N_9449);
and U10448 (N_10448,N_9146,N_9046);
xnor U10449 (N_10449,N_9692,N_9111);
nand U10450 (N_10450,N_9232,N_9916);
nand U10451 (N_10451,N_9398,N_9179);
nand U10452 (N_10452,N_9189,N_9454);
or U10453 (N_10453,N_9506,N_9518);
nor U10454 (N_10454,N_9515,N_9200);
nand U10455 (N_10455,N_9421,N_9187);
xnor U10456 (N_10456,N_9062,N_9778);
nor U10457 (N_10457,N_9476,N_9864);
nand U10458 (N_10458,N_9630,N_9549);
nand U10459 (N_10459,N_9180,N_9010);
xnor U10460 (N_10460,N_9075,N_9616);
nand U10461 (N_10461,N_9298,N_9564);
xnor U10462 (N_10462,N_9662,N_9079);
nor U10463 (N_10463,N_9242,N_9472);
nand U10464 (N_10464,N_9460,N_9303);
or U10465 (N_10465,N_9627,N_9154);
nor U10466 (N_10466,N_9668,N_9323);
nor U10467 (N_10467,N_9829,N_9534);
or U10468 (N_10468,N_9397,N_9987);
nor U10469 (N_10469,N_9099,N_9040);
or U10470 (N_10470,N_9239,N_9596);
and U10471 (N_10471,N_9785,N_9582);
or U10472 (N_10472,N_9347,N_9759);
nand U10473 (N_10473,N_9740,N_9781);
nor U10474 (N_10474,N_9409,N_9327);
and U10475 (N_10475,N_9488,N_9092);
and U10476 (N_10476,N_9606,N_9742);
and U10477 (N_10477,N_9268,N_9491);
and U10478 (N_10478,N_9172,N_9801);
xor U10479 (N_10479,N_9313,N_9171);
xor U10480 (N_10480,N_9817,N_9854);
and U10481 (N_10481,N_9366,N_9424);
nor U10482 (N_10482,N_9932,N_9804);
nor U10483 (N_10483,N_9660,N_9222);
and U10484 (N_10484,N_9821,N_9789);
nor U10485 (N_10485,N_9809,N_9490);
nand U10486 (N_10486,N_9537,N_9553);
nand U10487 (N_10487,N_9776,N_9162);
xor U10488 (N_10488,N_9867,N_9575);
or U10489 (N_10489,N_9765,N_9719);
nor U10490 (N_10490,N_9530,N_9284);
nand U10491 (N_10491,N_9043,N_9054);
nand U10492 (N_10492,N_9739,N_9053);
or U10493 (N_10493,N_9481,N_9554);
nor U10494 (N_10494,N_9208,N_9198);
and U10495 (N_10495,N_9346,N_9000);
xor U10496 (N_10496,N_9292,N_9889);
or U10497 (N_10497,N_9527,N_9786);
or U10498 (N_10498,N_9468,N_9320);
and U10499 (N_10499,N_9661,N_9041);
or U10500 (N_10500,N_9031,N_9160);
nor U10501 (N_10501,N_9026,N_9135);
nor U10502 (N_10502,N_9052,N_9279);
nor U10503 (N_10503,N_9045,N_9893);
or U10504 (N_10504,N_9368,N_9105);
and U10505 (N_10505,N_9819,N_9570);
and U10506 (N_10506,N_9332,N_9279);
or U10507 (N_10507,N_9719,N_9926);
nand U10508 (N_10508,N_9815,N_9385);
xor U10509 (N_10509,N_9939,N_9924);
xor U10510 (N_10510,N_9581,N_9423);
xor U10511 (N_10511,N_9260,N_9477);
and U10512 (N_10512,N_9800,N_9230);
or U10513 (N_10513,N_9508,N_9792);
nor U10514 (N_10514,N_9064,N_9511);
or U10515 (N_10515,N_9919,N_9547);
or U10516 (N_10516,N_9361,N_9145);
nand U10517 (N_10517,N_9131,N_9724);
or U10518 (N_10518,N_9433,N_9018);
or U10519 (N_10519,N_9738,N_9505);
nor U10520 (N_10520,N_9682,N_9389);
or U10521 (N_10521,N_9039,N_9070);
nand U10522 (N_10522,N_9967,N_9653);
nand U10523 (N_10523,N_9157,N_9861);
or U10524 (N_10524,N_9230,N_9202);
nor U10525 (N_10525,N_9211,N_9885);
and U10526 (N_10526,N_9811,N_9456);
nand U10527 (N_10527,N_9006,N_9890);
and U10528 (N_10528,N_9852,N_9194);
nor U10529 (N_10529,N_9491,N_9791);
and U10530 (N_10530,N_9934,N_9428);
xnor U10531 (N_10531,N_9818,N_9551);
nand U10532 (N_10532,N_9474,N_9446);
and U10533 (N_10533,N_9624,N_9051);
and U10534 (N_10534,N_9135,N_9202);
nand U10535 (N_10535,N_9593,N_9814);
nand U10536 (N_10536,N_9292,N_9692);
xnor U10537 (N_10537,N_9412,N_9399);
or U10538 (N_10538,N_9438,N_9735);
and U10539 (N_10539,N_9768,N_9472);
or U10540 (N_10540,N_9607,N_9201);
nand U10541 (N_10541,N_9843,N_9903);
or U10542 (N_10542,N_9804,N_9451);
or U10543 (N_10543,N_9971,N_9238);
and U10544 (N_10544,N_9763,N_9985);
or U10545 (N_10545,N_9661,N_9561);
nor U10546 (N_10546,N_9192,N_9440);
nand U10547 (N_10547,N_9253,N_9724);
xnor U10548 (N_10548,N_9002,N_9556);
nand U10549 (N_10549,N_9315,N_9825);
and U10550 (N_10550,N_9580,N_9848);
xor U10551 (N_10551,N_9686,N_9403);
and U10552 (N_10552,N_9851,N_9742);
xor U10553 (N_10553,N_9665,N_9913);
and U10554 (N_10554,N_9373,N_9205);
or U10555 (N_10555,N_9075,N_9156);
and U10556 (N_10556,N_9812,N_9965);
nor U10557 (N_10557,N_9100,N_9608);
xor U10558 (N_10558,N_9493,N_9495);
or U10559 (N_10559,N_9295,N_9098);
nor U10560 (N_10560,N_9862,N_9001);
and U10561 (N_10561,N_9767,N_9595);
and U10562 (N_10562,N_9742,N_9070);
and U10563 (N_10563,N_9242,N_9224);
and U10564 (N_10564,N_9052,N_9410);
or U10565 (N_10565,N_9885,N_9107);
xnor U10566 (N_10566,N_9526,N_9301);
or U10567 (N_10567,N_9166,N_9048);
or U10568 (N_10568,N_9724,N_9339);
nand U10569 (N_10569,N_9902,N_9078);
nor U10570 (N_10570,N_9252,N_9384);
or U10571 (N_10571,N_9267,N_9498);
nor U10572 (N_10572,N_9801,N_9097);
or U10573 (N_10573,N_9242,N_9209);
nor U10574 (N_10574,N_9057,N_9441);
xnor U10575 (N_10575,N_9940,N_9616);
or U10576 (N_10576,N_9131,N_9107);
nand U10577 (N_10577,N_9513,N_9884);
nor U10578 (N_10578,N_9682,N_9304);
nand U10579 (N_10579,N_9346,N_9707);
nand U10580 (N_10580,N_9755,N_9009);
and U10581 (N_10581,N_9924,N_9709);
nand U10582 (N_10582,N_9477,N_9714);
xnor U10583 (N_10583,N_9740,N_9329);
xnor U10584 (N_10584,N_9554,N_9787);
nand U10585 (N_10585,N_9727,N_9053);
nand U10586 (N_10586,N_9558,N_9896);
nand U10587 (N_10587,N_9603,N_9114);
nor U10588 (N_10588,N_9934,N_9438);
xor U10589 (N_10589,N_9277,N_9939);
nand U10590 (N_10590,N_9330,N_9466);
and U10591 (N_10591,N_9474,N_9720);
and U10592 (N_10592,N_9781,N_9136);
nor U10593 (N_10593,N_9246,N_9396);
nand U10594 (N_10594,N_9570,N_9149);
nor U10595 (N_10595,N_9939,N_9426);
or U10596 (N_10596,N_9680,N_9464);
nor U10597 (N_10597,N_9310,N_9465);
or U10598 (N_10598,N_9028,N_9762);
or U10599 (N_10599,N_9490,N_9850);
nor U10600 (N_10600,N_9941,N_9446);
and U10601 (N_10601,N_9022,N_9108);
or U10602 (N_10602,N_9588,N_9382);
nor U10603 (N_10603,N_9048,N_9950);
and U10604 (N_10604,N_9810,N_9072);
nand U10605 (N_10605,N_9021,N_9541);
nor U10606 (N_10606,N_9880,N_9263);
nor U10607 (N_10607,N_9298,N_9143);
or U10608 (N_10608,N_9297,N_9531);
nand U10609 (N_10609,N_9614,N_9303);
or U10610 (N_10610,N_9776,N_9129);
nand U10611 (N_10611,N_9136,N_9406);
or U10612 (N_10612,N_9544,N_9064);
xor U10613 (N_10613,N_9018,N_9286);
nand U10614 (N_10614,N_9442,N_9770);
nand U10615 (N_10615,N_9169,N_9613);
nand U10616 (N_10616,N_9180,N_9216);
and U10617 (N_10617,N_9110,N_9994);
xor U10618 (N_10618,N_9814,N_9810);
nand U10619 (N_10619,N_9069,N_9651);
nand U10620 (N_10620,N_9298,N_9033);
or U10621 (N_10621,N_9485,N_9176);
or U10622 (N_10622,N_9785,N_9021);
or U10623 (N_10623,N_9845,N_9962);
nand U10624 (N_10624,N_9483,N_9800);
and U10625 (N_10625,N_9120,N_9596);
nand U10626 (N_10626,N_9293,N_9366);
xor U10627 (N_10627,N_9623,N_9289);
nor U10628 (N_10628,N_9436,N_9253);
nand U10629 (N_10629,N_9594,N_9396);
xor U10630 (N_10630,N_9798,N_9179);
or U10631 (N_10631,N_9379,N_9964);
nor U10632 (N_10632,N_9417,N_9164);
or U10633 (N_10633,N_9025,N_9485);
or U10634 (N_10634,N_9633,N_9493);
xnor U10635 (N_10635,N_9810,N_9940);
nor U10636 (N_10636,N_9422,N_9450);
nand U10637 (N_10637,N_9677,N_9513);
xnor U10638 (N_10638,N_9153,N_9784);
nor U10639 (N_10639,N_9337,N_9950);
nand U10640 (N_10640,N_9064,N_9339);
nand U10641 (N_10641,N_9536,N_9660);
xnor U10642 (N_10642,N_9832,N_9588);
nand U10643 (N_10643,N_9139,N_9486);
or U10644 (N_10644,N_9017,N_9008);
and U10645 (N_10645,N_9147,N_9252);
and U10646 (N_10646,N_9407,N_9216);
or U10647 (N_10647,N_9538,N_9031);
or U10648 (N_10648,N_9515,N_9801);
nand U10649 (N_10649,N_9425,N_9959);
or U10650 (N_10650,N_9850,N_9386);
or U10651 (N_10651,N_9944,N_9187);
xor U10652 (N_10652,N_9412,N_9249);
and U10653 (N_10653,N_9447,N_9662);
nor U10654 (N_10654,N_9031,N_9095);
nand U10655 (N_10655,N_9113,N_9552);
nor U10656 (N_10656,N_9995,N_9772);
or U10657 (N_10657,N_9193,N_9265);
and U10658 (N_10658,N_9281,N_9678);
and U10659 (N_10659,N_9222,N_9094);
and U10660 (N_10660,N_9325,N_9020);
and U10661 (N_10661,N_9104,N_9403);
nand U10662 (N_10662,N_9598,N_9326);
and U10663 (N_10663,N_9863,N_9754);
or U10664 (N_10664,N_9718,N_9220);
nor U10665 (N_10665,N_9791,N_9481);
or U10666 (N_10666,N_9348,N_9564);
and U10667 (N_10667,N_9446,N_9727);
xor U10668 (N_10668,N_9663,N_9890);
nor U10669 (N_10669,N_9128,N_9215);
or U10670 (N_10670,N_9830,N_9269);
and U10671 (N_10671,N_9432,N_9163);
nand U10672 (N_10672,N_9124,N_9232);
nor U10673 (N_10673,N_9458,N_9839);
nand U10674 (N_10674,N_9444,N_9217);
xnor U10675 (N_10675,N_9022,N_9028);
and U10676 (N_10676,N_9249,N_9949);
and U10677 (N_10677,N_9503,N_9715);
xor U10678 (N_10678,N_9482,N_9668);
or U10679 (N_10679,N_9039,N_9902);
or U10680 (N_10680,N_9753,N_9331);
nor U10681 (N_10681,N_9687,N_9236);
and U10682 (N_10682,N_9225,N_9871);
nor U10683 (N_10683,N_9237,N_9144);
or U10684 (N_10684,N_9163,N_9002);
or U10685 (N_10685,N_9543,N_9593);
or U10686 (N_10686,N_9786,N_9257);
or U10687 (N_10687,N_9099,N_9565);
nand U10688 (N_10688,N_9457,N_9906);
nor U10689 (N_10689,N_9587,N_9750);
nor U10690 (N_10690,N_9838,N_9302);
and U10691 (N_10691,N_9658,N_9330);
nand U10692 (N_10692,N_9025,N_9390);
or U10693 (N_10693,N_9560,N_9975);
and U10694 (N_10694,N_9939,N_9225);
nor U10695 (N_10695,N_9549,N_9599);
and U10696 (N_10696,N_9595,N_9386);
nor U10697 (N_10697,N_9391,N_9991);
nand U10698 (N_10698,N_9034,N_9441);
nor U10699 (N_10699,N_9271,N_9395);
and U10700 (N_10700,N_9178,N_9892);
nor U10701 (N_10701,N_9337,N_9820);
or U10702 (N_10702,N_9709,N_9154);
nor U10703 (N_10703,N_9533,N_9746);
nor U10704 (N_10704,N_9583,N_9485);
or U10705 (N_10705,N_9554,N_9636);
nor U10706 (N_10706,N_9533,N_9568);
xor U10707 (N_10707,N_9803,N_9807);
or U10708 (N_10708,N_9110,N_9374);
nor U10709 (N_10709,N_9387,N_9143);
or U10710 (N_10710,N_9637,N_9470);
and U10711 (N_10711,N_9960,N_9390);
or U10712 (N_10712,N_9056,N_9734);
nor U10713 (N_10713,N_9331,N_9672);
nand U10714 (N_10714,N_9445,N_9508);
and U10715 (N_10715,N_9849,N_9351);
and U10716 (N_10716,N_9261,N_9085);
nor U10717 (N_10717,N_9591,N_9220);
and U10718 (N_10718,N_9745,N_9669);
xnor U10719 (N_10719,N_9082,N_9643);
nor U10720 (N_10720,N_9640,N_9296);
nor U10721 (N_10721,N_9177,N_9474);
nor U10722 (N_10722,N_9259,N_9734);
nand U10723 (N_10723,N_9814,N_9021);
or U10724 (N_10724,N_9369,N_9470);
and U10725 (N_10725,N_9314,N_9156);
nand U10726 (N_10726,N_9368,N_9015);
nor U10727 (N_10727,N_9427,N_9054);
and U10728 (N_10728,N_9954,N_9462);
xor U10729 (N_10729,N_9867,N_9963);
or U10730 (N_10730,N_9001,N_9012);
or U10731 (N_10731,N_9497,N_9867);
or U10732 (N_10732,N_9054,N_9049);
nor U10733 (N_10733,N_9510,N_9267);
nor U10734 (N_10734,N_9989,N_9492);
and U10735 (N_10735,N_9474,N_9917);
and U10736 (N_10736,N_9662,N_9950);
xnor U10737 (N_10737,N_9012,N_9094);
nor U10738 (N_10738,N_9563,N_9279);
nor U10739 (N_10739,N_9613,N_9358);
or U10740 (N_10740,N_9676,N_9620);
xor U10741 (N_10741,N_9971,N_9846);
xor U10742 (N_10742,N_9571,N_9873);
or U10743 (N_10743,N_9007,N_9185);
xor U10744 (N_10744,N_9871,N_9066);
nor U10745 (N_10745,N_9197,N_9483);
or U10746 (N_10746,N_9464,N_9097);
or U10747 (N_10747,N_9864,N_9189);
nand U10748 (N_10748,N_9707,N_9053);
nand U10749 (N_10749,N_9669,N_9853);
nand U10750 (N_10750,N_9832,N_9266);
and U10751 (N_10751,N_9493,N_9678);
nand U10752 (N_10752,N_9459,N_9872);
nor U10753 (N_10753,N_9139,N_9078);
nand U10754 (N_10754,N_9391,N_9047);
nand U10755 (N_10755,N_9147,N_9473);
nor U10756 (N_10756,N_9107,N_9288);
and U10757 (N_10757,N_9599,N_9678);
xnor U10758 (N_10758,N_9550,N_9706);
and U10759 (N_10759,N_9298,N_9169);
nand U10760 (N_10760,N_9838,N_9767);
or U10761 (N_10761,N_9900,N_9380);
nand U10762 (N_10762,N_9897,N_9520);
nand U10763 (N_10763,N_9790,N_9313);
or U10764 (N_10764,N_9386,N_9514);
and U10765 (N_10765,N_9782,N_9505);
or U10766 (N_10766,N_9844,N_9401);
or U10767 (N_10767,N_9906,N_9826);
and U10768 (N_10768,N_9802,N_9666);
and U10769 (N_10769,N_9036,N_9179);
nor U10770 (N_10770,N_9230,N_9777);
or U10771 (N_10771,N_9338,N_9942);
nand U10772 (N_10772,N_9525,N_9787);
nor U10773 (N_10773,N_9444,N_9893);
or U10774 (N_10774,N_9500,N_9528);
nand U10775 (N_10775,N_9642,N_9270);
nand U10776 (N_10776,N_9888,N_9795);
and U10777 (N_10777,N_9091,N_9558);
and U10778 (N_10778,N_9021,N_9728);
or U10779 (N_10779,N_9929,N_9677);
nand U10780 (N_10780,N_9228,N_9825);
nor U10781 (N_10781,N_9292,N_9569);
nand U10782 (N_10782,N_9633,N_9848);
and U10783 (N_10783,N_9402,N_9606);
and U10784 (N_10784,N_9647,N_9434);
or U10785 (N_10785,N_9612,N_9381);
and U10786 (N_10786,N_9714,N_9102);
or U10787 (N_10787,N_9213,N_9477);
nand U10788 (N_10788,N_9195,N_9331);
nor U10789 (N_10789,N_9632,N_9282);
or U10790 (N_10790,N_9274,N_9216);
or U10791 (N_10791,N_9730,N_9670);
nand U10792 (N_10792,N_9750,N_9639);
nand U10793 (N_10793,N_9308,N_9447);
and U10794 (N_10794,N_9540,N_9684);
xor U10795 (N_10795,N_9671,N_9717);
xnor U10796 (N_10796,N_9541,N_9754);
and U10797 (N_10797,N_9465,N_9437);
nor U10798 (N_10798,N_9781,N_9489);
xor U10799 (N_10799,N_9130,N_9829);
nand U10800 (N_10800,N_9823,N_9058);
xnor U10801 (N_10801,N_9505,N_9590);
nor U10802 (N_10802,N_9007,N_9276);
and U10803 (N_10803,N_9039,N_9010);
nand U10804 (N_10804,N_9915,N_9851);
xnor U10805 (N_10805,N_9245,N_9677);
nand U10806 (N_10806,N_9016,N_9874);
and U10807 (N_10807,N_9053,N_9890);
nor U10808 (N_10808,N_9922,N_9864);
and U10809 (N_10809,N_9780,N_9440);
nand U10810 (N_10810,N_9009,N_9338);
and U10811 (N_10811,N_9513,N_9895);
and U10812 (N_10812,N_9801,N_9163);
and U10813 (N_10813,N_9415,N_9281);
nor U10814 (N_10814,N_9472,N_9597);
nor U10815 (N_10815,N_9150,N_9985);
or U10816 (N_10816,N_9721,N_9690);
nor U10817 (N_10817,N_9220,N_9335);
nand U10818 (N_10818,N_9726,N_9008);
nand U10819 (N_10819,N_9404,N_9486);
nand U10820 (N_10820,N_9197,N_9771);
nand U10821 (N_10821,N_9275,N_9712);
nand U10822 (N_10822,N_9843,N_9136);
nand U10823 (N_10823,N_9234,N_9292);
nor U10824 (N_10824,N_9662,N_9168);
and U10825 (N_10825,N_9196,N_9869);
nor U10826 (N_10826,N_9475,N_9095);
and U10827 (N_10827,N_9883,N_9576);
nand U10828 (N_10828,N_9602,N_9321);
nand U10829 (N_10829,N_9080,N_9981);
nand U10830 (N_10830,N_9766,N_9602);
and U10831 (N_10831,N_9932,N_9354);
nand U10832 (N_10832,N_9150,N_9728);
nand U10833 (N_10833,N_9442,N_9934);
xor U10834 (N_10834,N_9866,N_9788);
and U10835 (N_10835,N_9259,N_9815);
nand U10836 (N_10836,N_9401,N_9094);
nor U10837 (N_10837,N_9663,N_9223);
or U10838 (N_10838,N_9467,N_9191);
or U10839 (N_10839,N_9529,N_9638);
xor U10840 (N_10840,N_9378,N_9853);
or U10841 (N_10841,N_9369,N_9899);
nand U10842 (N_10842,N_9678,N_9189);
xnor U10843 (N_10843,N_9230,N_9836);
and U10844 (N_10844,N_9648,N_9042);
and U10845 (N_10845,N_9530,N_9482);
or U10846 (N_10846,N_9810,N_9783);
or U10847 (N_10847,N_9801,N_9052);
and U10848 (N_10848,N_9579,N_9219);
or U10849 (N_10849,N_9282,N_9647);
xnor U10850 (N_10850,N_9926,N_9485);
nand U10851 (N_10851,N_9867,N_9778);
and U10852 (N_10852,N_9018,N_9490);
and U10853 (N_10853,N_9614,N_9237);
and U10854 (N_10854,N_9440,N_9838);
or U10855 (N_10855,N_9248,N_9362);
or U10856 (N_10856,N_9719,N_9319);
or U10857 (N_10857,N_9408,N_9929);
nand U10858 (N_10858,N_9055,N_9315);
nor U10859 (N_10859,N_9213,N_9941);
or U10860 (N_10860,N_9302,N_9906);
nand U10861 (N_10861,N_9508,N_9886);
nand U10862 (N_10862,N_9143,N_9430);
nand U10863 (N_10863,N_9892,N_9079);
nor U10864 (N_10864,N_9132,N_9509);
and U10865 (N_10865,N_9650,N_9369);
and U10866 (N_10866,N_9765,N_9241);
nand U10867 (N_10867,N_9646,N_9618);
nand U10868 (N_10868,N_9722,N_9636);
nor U10869 (N_10869,N_9245,N_9624);
nand U10870 (N_10870,N_9692,N_9606);
nor U10871 (N_10871,N_9257,N_9471);
nand U10872 (N_10872,N_9829,N_9661);
or U10873 (N_10873,N_9250,N_9192);
nand U10874 (N_10874,N_9470,N_9120);
or U10875 (N_10875,N_9385,N_9752);
xor U10876 (N_10876,N_9069,N_9140);
and U10877 (N_10877,N_9494,N_9229);
xor U10878 (N_10878,N_9006,N_9596);
nand U10879 (N_10879,N_9014,N_9042);
xor U10880 (N_10880,N_9886,N_9871);
or U10881 (N_10881,N_9474,N_9806);
xnor U10882 (N_10882,N_9878,N_9002);
xnor U10883 (N_10883,N_9722,N_9981);
nor U10884 (N_10884,N_9865,N_9210);
xnor U10885 (N_10885,N_9157,N_9669);
or U10886 (N_10886,N_9204,N_9844);
nor U10887 (N_10887,N_9044,N_9864);
nor U10888 (N_10888,N_9810,N_9380);
nand U10889 (N_10889,N_9106,N_9131);
nor U10890 (N_10890,N_9873,N_9037);
nor U10891 (N_10891,N_9911,N_9828);
xor U10892 (N_10892,N_9423,N_9644);
nor U10893 (N_10893,N_9867,N_9204);
nand U10894 (N_10894,N_9539,N_9682);
nor U10895 (N_10895,N_9317,N_9508);
xor U10896 (N_10896,N_9438,N_9589);
nor U10897 (N_10897,N_9880,N_9168);
or U10898 (N_10898,N_9262,N_9773);
nand U10899 (N_10899,N_9992,N_9124);
or U10900 (N_10900,N_9500,N_9529);
and U10901 (N_10901,N_9657,N_9802);
and U10902 (N_10902,N_9105,N_9365);
xnor U10903 (N_10903,N_9808,N_9614);
xor U10904 (N_10904,N_9679,N_9138);
nor U10905 (N_10905,N_9345,N_9656);
and U10906 (N_10906,N_9882,N_9953);
nand U10907 (N_10907,N_9915,N_9712);
xnor U10908 (N_10908,N_9031,N_9629);
or U10909 (N_10909,N_9800,N_9569);
and U10910 (N_10910,N_9191,N_9729);
nand U10911 (N_10911,N_9745,N_9248);
nand U10912 (N_10912,N_9075,N_9354);
and U10913 (N_10913,N_9257,N_9588);
nor U10914 (N_10914,N_9805,N_9065);
nand U10915 (N_10915,N_9904,N_9773);
nand U10916 (N_10916,N_9887,N_9536);
nand U10917 (N_10917,N_9128,N_9735);
and U10918 (N_10918,N_9800,N_9588);
or U10919 (N_10919,N_9852,N_9702);
and U10920 (N_10920,N_9667,N_9127);
and U10921 (N_10921,N_9584,N_9262);
or U10922 (N_10922,N_9068,N_9095);
nor U10923 (N_10923,N_9778,N_9137);
nand U10924 (N_10924,N_9029,N_9235);
xnor U10925 (N_10925,N_9531,N_9971);
nand U10926 (N_10926,N_9145,N_9100);
or U10927 (N_10927,N_9210,N_9459);
nand U10928 (N_10928,N_9334,N_9894);
nor U10929 (N_10929,N_9592,N_9505);
nand U10930 (N_10930,N_9296,N_9290);
nor U10931 (N_10931,N_9341,N_9584);
nand U10932 (N_10932,N_9689,N_9434);
nand U10933 (N_10933,N_9446,N_9743);
or U10934 (N_10934,N_9259,N_9973);
xor U10935 (N_10935,N_9335,N_9852);
xor U10936 (N_10936,N_9436,N_9987);
or U10937 (N_10937,N_9013,N_9037);
nor U10938 (N_10938,N_9085,N_9378);
or U10939 (N_10939,N_9841,N_9537);
nand U10940 (N_10940,N_9783,N_9064);
and U10941 (N_10941,N_9267,N_9776);
and U10942 (N_10942,N_9647,N_9206);
nor U10943 (N_10943,N_9092,N_9523);
and U10944 (N_10944,N_9303,N_9119);
nand U10945 (N_10945,N_9222,N_9158);
or U10946 (N_10946,N_9056,N_9279);
nor U10947 (N_10947,N_9815,N_9091);
nor U10948 (N_10948,N_9159,N_9905);
xnor U10949 (N_10949,N_9086,N_9530);
nand U10950 (N_10950,N_9554,N_9539);
or U10951 (N_10951,N_9965,N_9773);
nor U10952 (N_10952,N_9602,N_9545);
nor U10953 (N_10953,N_9569,N_9402);
and U10954 (N_10954,N_9131,N_9599);
and U10955 (N_10955,N_9272,N_9401);
nor U10956 (N_10956,N_9258,N_9585);
nor U10957 (N_10957,N_9773,N_9912);
nor U10958 (N_10958,N_9311,N_9061);
nand U10959 (N_10959,N_9609,N_9978);
xor U10960 (N_10960,N_9222,N_9178);
and U10961 (N_10961,N_9873,N_9961);
or U10962 (N_10962,N_9254,N_9441);
nor U10963 (N_10963,N_9896,N_9439);
nor U10964 (N_10964,N_9089,N_9864);
and U10965 (N_10965,N_9651,N_9276);
or U10966 (N_10966,N_9430,N_9545);
or U10967 (N_10967,N_9996,N_9034);
or U10968 (N_10968,N_9864,N_9701);
nand U10969 (N_10969,N_9265,N_9724);
xnor U10970 (N_10970,N_9290,N_9391);
or U10971 (N_10971,N_9390,N_9917);
or U10972 (N_10972,N_9768,N_9145);
and U10973 (N_10973,N_9686,N_9274);
and U10974 (N_10974,N_9769,N_9646);
nand U10975 (N_10975,N_9791,N_9862);
and U10976 (N_10976,N_9239,N_9232);
or U10977 (N_10977,N_9222,N_9712);
nand U10978 (N_10978,N_9523,N_9484);
nand U10979 (N_10979,N_9418,N_9326);
and U10980 (N_10980,N_9220,N_9914);
or U10981 (N_10981,N_9705,N_9962);
xnor U10982 (N_10982,N_9951,N_9667);
nand U10983 (N_10983,N_9485,N_9886);
nor U10984 (N_10984,N_9054,N_9771);
nand U10985 (N_10985,N_9951,N_9715);
nor U10986 (N_10986,N_9533,N_9921);
and U10987 (N_10987,N_9474,N_9829);
xor U10988 (N_10988,N_9257,N_9153);
nand U10989 (N_10989,N_9414,N_9076);
and U10990 (N_10990,N_9088,N_9198);
nor U10991 (N_10991,N_9817,N_9286);
or U10992 (N_10992,N_9869,N_9703);
and U10993 (N_10993,N_9562,N_9737);
and U10994 (N_10994,N_9781,N_9954);
xnor U10995 (N_10995,N_9644,N_9310);
and U10996 (N_10996,N_9625,N_9266);
xnor U10997 (N_10997,N_9407,N_9246);
nand U10998 (N_10998,N_9233,N_9660);
nor U10999 (N_10999,N_9308,N_9414);
nor U11000 (N_11000,N_10172,N_10980);
nor U11001 (N_11001,N_10716,N_10624);
or U11002 (N_11002,N_10938,N_10569);
or U11003 (N_11003,N_10465,N_10259);
or U11004 (N_11004,N_10018,N_10575);
or U11005 (N_11005,N_10255,N_10698);
nor U11006 (N_11006,N_10142,N_10444);
nor U11007 (N_11007,N_10615,N_10048);
nand U11008 (N_11008,N_10801,N_10198);
or U11009 (N_11009,N_10295,N_10217);
nand U11010 (N_11010,N_10260,N_10239);
and U11011 (N_11011,N_10301,N_10655);
nor U11012 (N_11012,N_10755,N_10478);
nor U11013 (N_11013,N_10505,N_10925);
nand U11014 (N_11014,N_10396,N_10237);
nand U11015 (N_11015,N_10376,N_10857);
nor U11016 (N_11016,N_10009,N_10571);
and U11017 (N_11017,N_10795,N_10016);
and U11018 (N_11018,N_10041,N_10882);
nor U11019 (N_11019,N_10401,N_10119);
nand U11020 (N_11020,N_10178,N_10727);
and U11021 (N_11021,N_10865,N_10961);
and U11022 (N_11022,N_10513,N_10429);
or U11023 (N_11023,N_10752,N_10274);
and U11024 (N_11024,N_10231,N_10621);
nand U11025 (N_11025,N_10032,N_10663);
xnor U11026 (N_11026,N_10361,N_10993);
nand U11027 (N_11027,N_10304,N_10927);
and U11028 (N_11028,N_10856,N_10890);
and U11029 (N_11029,N_10717,N_10699);
or U11030 (N_11030,N_10149,N_10991);
xnor U11031 (N_11031,N_10736,N_10166);
or U11032 (N_11032,N_10597,N_10601);
or U11033 (N_11033,N_10103,N_10303);
nand U11034 (N_11034,N_10293,N_10090);
nand U11035 (N_11035,N_10386,N_10483);
nand U11036 (N_11036,N_10824,N_10999);
nand U11037 (N_11037,N_10776,N_10711);
or U11038 (N_11038,N_10940,N_10366);
or U11039 (N_11039,N_10443,N_10430);
xnor U11040 (N_11040,N_10768,N_10964);
nor U11041 (N_11041,N_10791,N_10334);
nor U11042 (N_11042,N_10249,N_10404);
and U11043 (N_11043,N_10760,N_10447);
nand U11044 (N_11044,N_10081,N_10657);
and U11045 (N_11045,N_10855,N_10536);
xnor U11046 (N_11046,N_10286,N_10683);
nand U11047 (N_11047,N_10313,N_10127);
xnor U11048 (N_11048,N_10561,N_10472);
or U11049 (N_11049,N_10549,N_10954);
and U11050 (N_11050,N_10547,N_10137);
nand U11051 (N_11051,N_10029,N_10317);
nand U11052 (N_11052,N_10641,N_10735);
and U11053 (N_11053,N_10634,N_10240);
and U11054 (N_11054,N_10230,N_10794);
or U11055 (N_11055,N_10947,N_10086);
nand U11056 (N_11056,N_10011,N_10061);
nor U11057 (N_11057,N_10963,N_10729);
nand U11058 (N_11058,N_10251,N_10777);
or U11059 (N_11059,N_10374,N_10704);
nand U11060 (N_11060,N_10728,N_10682);
nor U11061 (N_11061,N_10510,N_10707);
or U11062 (N_11062,N_10144,N_10842);
or U11063 (N_11063,N_10025,N_10992);
nand U11064 (N_11064,N_10299,N_10676);
xor U11065 (N_11065,N_10382,N_10343);
and U11066 (N_11066,N_10845,N_10452);
or U11067 (N_11067,N_10461,N_10858);
or U11068 (N_11068,N_10246,N_10241);
and U11069 (N_11069,N_10347,N_10455);
xor U11070 (N_11070,N_10123,N_10407);
and U11071 (N_11071,N_10079,N_10595);
or U11072 (N_11072,N_10527,N_10170);
nand U11073 (N_11073,N_10941,N_10365);
nand U11074 (N_11074,N_10434,N_10418);
nor U11075 (N_11075,N_10248,N_10796);
nor U11076 (N_11076,N_10692,N_10083);
or U11077 (N_11077,N_10821,N_10490);
or U11078 (N_11078,N_10691,N_10793);
and U11079 (N_11079,N_10179,N_10305);
and U11080 (N_11080,N_10417,N_10633);
nor U11081 (N_11081,N_10713,N_10405);
and U11082 (N_11082,N_10587,N_10651);
nand U11083 (N_11083,N_10918,N_10630);
or U11084 (N_11084,N_10010,N_10610);
nand U11085 (N_11085,N_10757,N_10785);
or U11086 (N_11086,N_10849,N_10403);
or U11087 (N_11087,N_10390,N_10371);
xnor U11088 (N_11088,N_10470,N_10631);
nand U11089 (N_11089,N_10213,N_10649);
nand U11090 (N_11090,N_10422,N_10021);
and U11091 (N_11091,N_10773,N_10071);
or U11092 (N_11092,N_10135,N_10830);
and U11093 (N_11093,N_10911,N_10111);
xor U11094 (N_11094,N_10360,N_10700);
or U11095 (N_11095,N_10618,N_10158);
nor U11096 (N_11096,N_10632,N_10994);
or U11097 (N_11097,N_10955,N_10074);
nor U11098 (N_11098,N_10840,N_10296);
nor U11099 (N_11099,N_10531,N_10266);
and U11100 (N_11100,N_10984,N_10550);
nand U11101 (N_11101,N_10096,N_10620);
nand U11102 (N_11102,N_10533,N_10590);
or U11103 (N_11103,N_10194,N_10015);
and U11104 (N_11104,N_10945,N_10221);
nor U11105 (N_11105,N_10362,N_10986);
nor U11106 (N_11106,N_10863,N_10236);
or U11107 (N_11107,N_10934,N_10888);
xor U11108 (N_11108,N_10501,N_10432);
or U11109 (N_11109,N_10666,N_10391);
nand U11110 (N_11110,N_10280,N_10530);
and U11111 (N_11111,N_10572,N_10839);
and U11112 (N_11112,N_10114,N_10315);
or U11113 (N_11113,N_10415,N_10869);
nor U11114 (N_11114,N_10492,N_10147);
or U11115 (N_11115,N_10007,N_10148);
and U11116 (N_11116,N_10891,N_10277);
or U11117 (N_11117,N_10051,N_10364);
nor U11118 (N_11118,N_10215,N_10953);
nor U11119 (N_11119,N_10662,N_10759);
nor U11120 (N_11120,N_10060,N_10384);
or U11121 (N_11121,N_10827,N_10988);
and U11122 (N_11122,N_10431,N_10859);
nor U11123 (N_11123,N_10762,N_10106);
xnor U11124 (N_11124,N_10093,N_10720);
or U11125 (N_11125,N_10926,N_10851);
nand U11126 (N_11126,N_10502,N_10087);
or U11127 (N_11127,N_10958,N_10639);
or U11128 (N_11128,N_10543,N_10970);
nand U11129 (N_11129,N_10529,N_10562);
xnor U11130 (N_11130,N_10555,N_10837);
or U11131 (N_11131,N_10073,N_10541);
or U11132 (N_11132,N_10544,N_10894);
nand U11133 (N_11133,N_10145,N_10834);
and U11134 (N_11134,N_10576,N_10514);
nor U11135 (N_11135,N_10050,N_10458);
nand U11136 (N_11136,N_10611,N_10772);
and U11137 (N_11137,N_10748,N_10730);
nor U11138 (N_11138,N_10696,N_10878);
nor U11139 (N_11139,N_10302,N_10121);
nand U11140 (N_11140,N_10151,N_10416);
nand U11141 (N_11141,N_10804,N_10424);
nand U11142 (N_11142,N_10314,N_10598);
or U11143 (N_11143,N_10517,N_10936);
and U11144 (N_11144,N_10136,N_10578);
and U11145 (N_11145,N_10281,N_10512);
and U11146 (N_11146,N_10603,N_10116);
or U11147 (N_11147,N_10614,N_10175);
nor U11148 (N_11148,N_10053,N_10037);
nand U11149 (N_11149,N_10921,N_10905);
and U11150 (N_11150,N_10881,N_10250);
and U11151 (N_11151,N_10895,N_10697);
or U11152 (N_11152,N_10781,N_10627);
nor U11153 (N_11153,N_10625,N_10787);
nor U11154 (N_11154,N_10216,N_10181);
nor U11155 (N_11155,N_10565,N_10798);
and U11156 (N_11156,N_10409,N_10400);
nor U11157 (N_11157,N_10721,N_10256);
or U11158 (N_11158,N_10423,N_10650);
nor U11159 (N_11159,N_10695,N_10414);
nand U11160 (N_11160,N_10703,N_10171);
nand U11161 (N_11161,N_10024,N_10321);
nand U11162 (N_11162,N_10002,N_10352);
or U11163 (N_11163,N_10033,N_10591);
nand U11164 (N_11164,N_10893,N_10998);
or U11165 (N_11165,N_10677,N_10885);
nand U11166 (N_11166,N_10104,N_10658);
and U11167 (N_11167,N_10130,N_10197);
and U11168 (N_11168,N_10671,N_10069);
nand U11169 (N_11169,N_10039,N_10107);
nor U11170 (N_11170,N_10460,N_10319);
nor U11171 (N_11171,N_10066,N_10402);
nand U11172 (N_11172,N_10826,N_10968);
nor U11173 (N_11173,N_10232,N_10388);
nand U11174 (N_11174,N_10645,N_10264);
nor U11175 (N_11175,N_10504,N_10210);
and U11176 (N_11176,N_10348,N_10099);
nand U11177 (N_11177,N_10628,N_10901);
and U11178 (N_11178,N_10582,N_10883);
nor U11179 (N_11179,N_10389,N_10908);
and U11180 (N_11180,N_10880,N_10814);
or U11181 (N_11181,N_10258,N_10316);
nand U11182 (N_11182,N_10267,N_10588);
or U11183 (N_11183,N_10556,N_10976);
and U11184 (N_11184,N_10548,N_10291);
or U11185 (N_11185,N_10327,N_10480);
or U11186 (N_11186,N_10937,N_10740);
nor U11187 (N_11187,N_10643,N_10006);
or U11188 (N_11188,N_10346,N_10511);
nand U11189 (N_11189,N_10674,N_10503);
xor U11190 (N_11190,N_10488,N_10325);
and U11191 (N_11191,N_10373,N_10584);
and U11192 (N_11192,N_10479,N_10208);
or U11193 (N_11193,N_10448,N_10499);
xnor U11194 (N_11194,N_10623,N_10219);
or U11195 (N_11195,N_10163,N_10214);
nor U11196 (N_11196,N_10358,N_10985);
or U11197 (N_11197,N_10846,N_10898);
xnor U11198 (N_11198,N_10949,N_10309);
nand U11199 (N_11199,N_10900,N_10084);
nor U11200 (N_11200,N_10693,N_10741);
nand U11201 (N_11201,N_10951,N_10323);
or U11202 (N_11202,N_10000,N_10800);
nor U11203 (N_11203,N_10355,N_10310);
nor U11204 (N_11204,N_10743,N_10224);
or U11205 (N_11205,N_10385,N_10056);
and U11206 (N_11206,N_10031,N_10195);
nand U11207 (N_11207,N_10477,N_10844);
or U11208 (N_11208,N_10177,N_10290);
and U11209 (N_11209,N_10924,N_10944);
nand U11210 (N_11210,N_10660,N_10899);
or U11211 (N_11211,N_10468,N_10471);
nor U11212 (N_11212,N_10235,N_10742);
nor U11213 (N_11213,N_10738,N_10819);
or U11214 (N_11214,N_10435,N_10823);
nand U11215 (N_11215,N_10218,N_10694);
and U11216 (N_11216,N_10320,N_10126);
or U11217 (N_11217,N_10068,N_10661);
nor U11218 (N_11218,N_10876,N_10825);
and U11219 (N_11219,N_10872,N_10943);
or U11220 (N_11220,N_10581,N_10124);
nand U11221 (N_11221,N_10012,N_10690);
or U11222 (N_11222,N_10515,N_10560);
nand U11223 (N_11223,N_10853,N_10831);
and U11224 (N_11224,N_10270,N_10324);
nand U11225 (N_11225,N_10629,N_10211);
or U11226 (N_11226,N_10586,N_10428);
nor U11227 (N_11227,N_10257,N_10356);
xor U11228 (N_11228,N_10585,N_10678);
nand U11229 (N_11229,N_10102,N_10120);
and U11230 (N_11230,N_10558,N_10363);
or U11231 (N_11231,N_10017,N_10318);
nand U11232 (N_11232,N_10962,N_10289);
and U11233 (N_11233,N_10987,N_10808);
xor U11234 (N_11234,N_10912,N_10688);
or U11235 (N_11235,N_10708,N_10080);
and U11236 (N_11236,N_10854,N_10566);
and U11237 (N_11237,N_10298,N_10487);
or U11238 (N_11238,N_10058,N_10750);
xor U11239 (N_11239,N_10563,N_10372);
nor U11240 (N_11240,N_10836,N_10220);
and U11241 (N_11241,N_10522,N_10702);
nor U11242 (N_11242,N_10790,N_10705);
or U11243 (N_11243,N_10023,N_10718);
or U11244 (N_11244,N_10841,N_10493);
and U11245 (N_11245,N_10710,N_10684);
and U11246 (N_11246,N_10916,N_10605);
xor U11247 (N_11247,N_10331,N_10254);
or U11248 (N_11248,N_10817,N_10134);
xor U11249 (N_11249,N_10789,N_10019);
nor U11250 (N_11250,N_10832,N_10336);
and U11251 (N_11251,N_10734,N_10689);
or U11252 (N_11252,N_10764,N_10110);
nand U11253 (N_11253,N_10180,N_10408);
nand U11254 (N_11254,N_10063,N_10067);
or U11255 (N_11255,N_10542,N_10654);
nor U11256 (N_11256,N_10199,N_10196);
and U11257 (N_11257,N_10187,N_10338);
or U11258 (N_11258,N_10108,N_10227);
nor U11259 (N_11259,N_10481,N_10269);
xnor U11260 (N_11260,N_10835,N_10131);
or U11261 (N_11261,N_10820,N_10969);
nand U11262 (N_11262,N_10636,N_10456);
nand U11263 (N_11263,N_10829,N_10739);
nor U11264 (N_11264,N_10112,N_10770);
nor U11265 (N_11265,N_10775,N_10959);
and U11266 (N_11266,N_10604,N_10028);
nor U11267 (N_11267,N_10642,N_10329);
xnor U11268 (N_11268,N_10972,N_10904);
xor U11269 (N_11269,N_10557,N_10525);
nor U11270 (N_11270,N_10341,N_10202);
nand U11271 (N_11271,N_10780,N_10744);
or U11272 (N_11272,N_10173,N_10647);
and U11273 (N_11273,N_10152,N_10767);
and U11274 (N_11274,N_10877,N_10375);
nor U11275 (N_11275,N_10109,N_10380);
nand U11276 (N_11276,N_10207,N_10635);
and U11277 (N_11277,N_10370,N_10105);
nor U11278 (N_11278,N_10507,N_10013);
nand U11279 (N_11279,N_10065,N_10769);
and U11280 (N_11280,N_10852,N_10439);
nor U11281 (N_11281,N_10279,N_10129);
nor U11282 (N_11282,N_10225,N_10995);
nor U11283 (N_11283,N_10973,N_10378);
or U11284 (N_11284,N_10589,N_10498);
and U11285 (N_11285,N_10810,N_10681);
or U11286 (N_11286,N_10935,N_10828);
nor U11287 (N_11287,N_10054,N_10003);
or U11288 (N_11288,N_10540,N_10297);
or U11289 (N_11289,N_10640,N_10005);
xor U11290 (N_11290,N_10596,N_10545);
xor U11291 (N_11291,N_10866,N_10273);
nor U11292 (N_11292,N_10245,N_10141);
xor U11293 (N_11293,N_10608,N_10359);
nor U11294 (N_11294,N_10622,N_10164);
and U11295 (N_11295,N_10607,N_10047);
nand U11296 (N_11296,N_10797,N_10395);
or U11297 (N_11297,N_10599,N_10523);
nand U11298 (N_11298,N_10043,N_10648);
nor U11299 (N_11299,N_10537,N_10433);
and U11300 (N_11300,N_10156,N_10082);
nand U11301 (N_11301,N_10485,N_10484);
xor U11302 (N_11302,N_10191,N_10884);
or U11303 (N_11303,N_10095,N_10307);
and U11304 (N_11304,N_10754,N_10075);
xor U11305 (N_11305,N_10150,N_10466);
and U11306 (N_11306,N_10115,N_10766);
or U11307 (N_11307,N_10722,N_10871);
or U11308 (N_11308,N_10157,N_10606);
nor U11309 (N_11309,N_10592,N_10387);
nand U11310 (N_11310,N_10494,N_10807);
or U11311 (N_11311,N_10714,N_10816);
and U11312 (N_11312,N_10538,N_10097);
or U11313 (N_11313,N_10806,N_10091);
nor U11314 (N_11314,N_10539,N_10726);
nor U11315 (N_11315,N_10756,N_10686);
xor U11316 (N_11316,N_10931,N_10209);
nand U11317 (N_11317,N_10903,N_10638);
nor U11318 (N_11318,N_10920,N_10753);
nand U11319 (N_11319,N_10185,N_10344);
or U11320 (N_11320,N_10244,N_10763);
nor U11321 (N_11321,N_10919,N_10410);
and U11322 (N_11322,N_10300,N_10799);
nand U11323 (N_11323,N_10950,N_10783);
or U11324 (N_11324,N_10875,N_10613);
xor U11325 (N_11325,N_10008,N_10906);
xnor U11326 (N_11326,N_10887,N_10860);
nand U11327 (N_11327,N_10519,N_10474);
nand U11328 (N_11328,N_10496,N_10778);
xor U11329 (N_11329,N_10026,N_10965);
or U11330 (N_11330,N_10437,N_10521);
and U11331 (N_11331,N_10282,N_10328);
xor U11332 (N_11332,N_10974,N_10377);
nor U11333 (N_11333,N_10553,N_10271);
nor U11334 (N_11334,N_10929,N_10100);
nand U11335 (N_11335,N_10574,N_10275);
and U11336 (N_11336,N_10670,N_10774);
nor U11337 (N_11337,N_10602,N_10265);
nor U11338 (N_11338,N_10724,N_10983);
and U11339 (N_11339,N_10161,N_10917);
xor U11340 (N_11340,N_10311,N_10247);
nor U11341 (N_11341,N_10782,N_10914);
or U11342 (N_11342,N_10982,N_10679);
nand U11343 (N_11343,N_10233,N_10731);
or U11344 (N_11344,N_10189,N_10709);
nand U11345 (N_11345,N_10712,N_10526);
or U11346 (N_11346,N_10680,N_10870);
and U11347 (N_11347,N_10577,N_10457);
or U11348 (N_11348,N_10652,N_10222);
nor U11349 (N_11349,N_10646,N_10838);
xnor U11350 (N_11350,N_10340,N_10140);
xor U11351 (N_11351,N_10500,N_10125);
or U11352 (N_11352,N_10438,N_10552);
nor U11353 (N_11353,N_10534,N_10188);
or U11354 (N_11354,N_10508,N_10867);
and U11355 (N_11355,N_10672,N_10491);
and U11356 (N_11356,N_10788,N_10292);
nor U11357 (N_11357,N_10568,N_10229);
or U11358 (N_11358,N_10203,N_10659);
and U11359 (N_11359,N_10128,N_10354);
nand U11360 (N_11360,N_10205,N_10809);
and U11361 (N_11361,N_10668,N_10101);
nor U11362 (N_11362,N_10892,N_10412);
and U11363 (N_11363,N_10847,N_10052);
or U11364 (N_11364,N_10656,N_10922);
and U11365 (N_11365,N_10312,N_10368);
and U11366 (N_11366,N_10383,N_10886);
or U11367 (N_11367,N_10057,N_10154);
or U11368 (N_11368,N_10546,N_10706);
or U11369 (N_11369,N_10879,N_10139);
nor U11370 (N_11370,N_10996,N_10072);
or U11371 (N_11371,N_10459,N_10913);
or U11372 (N_11372,N_10284,N_10669);
and U11373 (N_11373,N_10242,N_10786);
nand U11374 (N_11374,N_10909,N_10436);
xnor U11375 (N_11375,N_10176,N_10528);
nor U11376 (N_11376,N_10805,N_10326);
xnor U11377 (N_11377,N_10520,N_10524);
and U11378 (N_11378,N_10088,N_10896);
nand U11379 (N_11379,N_10966,N_10077);
nand U11380 (N_11380,N_10392,N_10948);
nand U11381 (N_11381,N_10813,N_10200);
and U11382 (N_11382,N_10567,N_10206);
nor U11383 (N_11383,N_10667,N_10771);
or U11384 (N_11384,N_10420,N_10153);
xor U11385 (N_11385,N_10322,N_10287);
nor U11386 (N_11386,N_10579,N_10022);
or U11387 (N_11387,N_10915,N_10978);
or U11388 (N_11388,N_10035,N_10308);
nand U11389 (N_11389,N_10283,N_10049);
or U11390 (N_11390,N_10653,N_10942);
and U11391 (N_11391,N_10160,N_10143);
nand U11392 (N_11392,N_10045,N_10559);
and U11393 (N_11393,N_10473,N_10272);
or U11394 (N_11394,N_10042,N_10070);
and U11395 (N_11395,N_10843,N_10850);
xor U11396 (N_11396,N_10746,N_10803);
nand U11397 (N_11397,N_10454,N_10059);
nor U11398 (N_11398,N_10747,N_10989);
and U11399 (N_11399,N_10394,N_10467);
nand U11400 (N_11400,N_10333,N_10441);
nor U11401 (N_11401,N_10446,N_10593);
and U11402 (N_11402,N_10497,N_10902);
or U11403 (N_11403,N_10779,N_10268);
or U11404 (N_11404,N_10910,N_10113);
or U11405 (N_11405,N_10737,N_10535);
nor U11406 (N_11406,N_10122,N_10092);
and U11407 (N_11407,N_10462,N_10811);
and U11408 (N_11408,N_10085,N_10078);
or U11409 (N_11409,N_10001,N_10133);
nand U11410 (N_11410,N_10398,N_10367);
or U11411 (N_11411,N_10223,N_10971);
and U11412 (N_11412,N_10228,N_10288);
or U11413 (N_11413,N_10040,N_10294);
nand U11414 (N_11414,N_10076,N_10184);
xor U11415 (N_11415,N_10226,N_10014);
nand U11416 (N_11416,N_10723,N_10673);
or U11417 (N_11417,N_10204,N_10862);
and U11418 (N_11418,N_10476,N_10960);
and U11419 (N_11419,N_10263,N_10345);
nor U11420 (N_11420,N_10977,N_10238);
nand U11421 (N_11421,N_10617,N_10532);
or U11422 (N_11422,N_10815,N_10637);
nor U11423 (N_11423,N_10165,N_10733);
or U11424 (N_11424,N_10118,N_10933);
nand U11425 (N_11425,N_10353,N_10406);
and U11426 (N_11426,N_10253,N_10193);
nand U11427 (N_11427,N_10411,N_10337);
and U11428 (N_11428,N_10725,N_10952);
nor U11429 (N_11429,N_10609,N_10046);
xnor U11430 (N_11430,N_10034,N_10981);
nand U11431 (N_11431,N_10551,N_10956);
nand U11432 (N_11432,N_10138,N_10168);
and U11433 (N_11433,N_10463,N_10749);
nand U11434 (N_11434,N_10475,N_10201);
xor U11435 (N_11435,N_10427,N_10393);
xnor U11436 (N_11436,N_10020,N_10278);
and U11437 (N_11437,N_10687,N_10453);
and U11438 (N_11438,N_10594,N_10818);
or U11439 (N_11439,N_10469,N_10167);
nor U11440 (N_11440,N_10030,N_10132);
and U11441 (N_11441,N_10907,N_10413);
and U11442 (N_11442,N_10451,N_10350);
and U11443 (N_11443,N_10330,N_10261);
nand U11444 (N_11444,N_10812,N_10967);
and U11445 (N_11445,N_10745,N_10044);
and U11446 (N_11446,N_10833,N_10306);
or U11447 (N_11447,N_10159,N_10186);
nand U11448 (N_11448,N_10062,N_10445);
nor U11449 (N_11449,N_10162,N_10094);
or U11450 (N_11450,N_10155,N_10685);
or U11451 (N_11451,N_10234,N_10064);
nor U11452 (N_11452,N_10212,N_10861);
nand U11453 (N_11453,N_10923,N_10506);
nand U11454 (N_11454,N_10252,N_10421);
xor U11455 (N_11455,N_10399,N_10616);
xnor U11456 (N_11456,N_10285,N_10675);
or U11457 (N_11457,N_10339,N_10975);
nand U11458 (N_11458,N_10486,N_10719);
and U11459 (N_11459,N_10516,N_10440);
or U11460 (N_11460,N_10644,N_10379);
and U11461 (N_11461,N_10027,N_10276);
or U11462 (N_11462,N_10939,N_10038);
nand U11463 (N_11463,N_10117,N_10357);
nand U11464 (N_11464,N_10419,N_10848);
xor U11465 (N_11465,N_10089,N_10174);
and U11466 (N_11466,N_10715,N_10802);
nor U11467 (N_11467,N_10619,N_10946);
xnor U11468 (N_11468,N_10489,N_10751);
and U11469 (N_11469,N_10182,N_10928);
xor U11470 (N_11470,N_10997,N_10868);
xor U11471 (N_11471,N_10495,N_10442);
nand U11472 (N_11472,N_10450,N_10874);
xnor U11473 (N_11473,N_10957,N_10701);
and U11474 (N_11474,N_10564,N_10765);
nand U11475 (N_11475,N_10381,N_10192);
or U11476 (N_11476,N_10873,N_10889);
and U11477 (N_11477,N_10146,N_10518);
nor U11478 (N_11478,N_10784,N_10897);
or U11479 (N_11479,N_10335,N_10397);
nor U11480 (N_11480,N_10612,N_10570);
or U11481 (N_11481,N_10580,N_10600);
and U11482 (N_11482,N_10369,N_10190);
or U11483 (N_11483,N_10732,N_10664);
and U11484 (N_11484,N_10262,N_10098);
nand U11485 (N_11485,N_10758,N_10979);
nand U11486 (N_11486,N_10349,N_10990);
or U11487 (N_11487,N_10449,N_10509);
or U11488 (N_11488,N_10573,N_10792);
nand U11489 (N_11489,N_10425,N_10004);
or U11490 (N_11490,N_10036,N_10426);
or U11491 (N_11491,N_10626,N_10342);
nor U11492 (N_11492,N_10351,N_10864);
and U11493 (N_11493,N_10932,N_10583);
xor U11494 (N_11494,N_10482,N_10464);
xnor U11495 (N_11495,N_10665,N_10554);
xor U11496 (N_11496,N_10930,N_10183);
nor U11497 (N_11497,N_10169,N_10332);
nand U11498 (N_11498,N_10761,N_10822);
or U11499 (N_11499,N_10055,N_10243);
or U11500 (N_11500,N_10891,N_10297);
and U11501 (N_11501,N_10395,N_10245);
nor U11502 (N_11502,N_10584,N_10247);
nand U11503 (N_11503,N_10459,N_10038);
and U11504 (N_11504,N_10180,N_10560);
nand U11505 (N_11505,N_10115,N_10062);
or U11506 (N_11506,N_10155,N_10410);
nor U11507 (N_11507,N_10831,N_10286);
nor U11508 (N_11508,N_10860,N_10764);
or U11509 (N_11509,N_10936,N_10498);
nand U11510 (N_11510,N_10437,N_10979);
nor U11511 (N_11511,N_10435,N_10582);
nor U11512 (N_11512,N_10135,N_10396);
or U11513 (N_11513,N_10461,N_10049);
nand U11514 (N_11514,N_10933,N_10712);
nor U11515 (N_11515,N_10704,N_10306);
and U11516 (N_11516,N_10769,N_10188);
nor U11517 (N_11517,N_10357,N_10338);
nand U11518 (N_11518,N_10394,N_10881);
or U11519 (N_11519,N_10985,N_10301);
and U11520 (N_11520,N_10763,N_10543);
and U11521 (N_11521,N_10612,N_10870);
nor U11522 (N_11522,N_10106,N_10301);
nor U11523 (N_11523,N_10830,N_10266);
nor U11524 (N_11524,N_10384,N_10523);
and U11525 (N_11525,N_10485,N_10875);
nor U11526 (N_11526,N_10977,N_10430);
and U11527 (N_11527,N_10111,N_10242);
nand U11528 (N_11528,N_10911,N_10960);
nor U11529 (N_11529,N_10177,N_10902);
xnor U11530 (N_11530,N_10746,N_10353);
nand U11531 (N_11531,N_10956,N_10050);
and U11532 (N_11532,N_10601,N_10028);
or U11533 (N_11533,N_10246,N_10826);
or U11534 (N_11534,N_10100,N_10082);
nor U11535 (N_11535,N_10699,N_10187);
and U11536 (N_11536,N_10105,N_10369);
and U11537 (N_11537,N_10042,N_10097);
nor U11538 (N_11538,N_10170,N_10707);
nor U11539 (N_11539,N_10596,N_10746);
nand U11540 (N_11540,N_10357,N_10290);
or U11541 (N_11541,N_10732,N_10837);
xnor U11542 (N_11542,N_10412,N_10426);
xor U11543 (N_11543,N_10233,N_10736);
nor U11544 (N_11544,N_10278,N_10053);
nor U11545 (N_11545,N_10523,N_10676);
xnor U11546 (N_11546,N_10939,N_10164);
nand U11547 (N_11547,N_10175,N_10160);
nand U11548 (N_11548,N_10558,N_10001);
nand U11549 (N_11549,N_10408,N_10101);
nor U11550 (N_11550,N_10259,N_10734);
or U11551 (N_11551,N_10818,N_10338);
nor U11552 (N_11552,N_10246,N_10456);
and U11553 (N_11553,N_10757,N_10129);
nand U11554 (N_11554,N_10127,N_10965);
xnor U11555 (N_11555,N_10694,N_10363);
or U11556 (N_11556,N_10346,N_10499);
and U11557 (N_11557,N_10967,N_10425);
nand U11558 (N_11558,N_10656,N_10328);
and U11559 (N_11559,N_10382,N_10918);
xor U11560 (N_11560,N_10038,N_10829);
and U11561 (N_11561,N_10042,N_10301);
nand U11562 (N_11562,N_10816,N_10887);
and U11563 (N_11563,N_10043,N_10362);
and U11564 (N_11564,N_10055,N_10271);
or U11565 (N_11565,N_10105,N_10714);
nor U11566 (N_11566,N_10064,N_10807);
or U11567 (N_11567,N_10722,N_10440);
nand U11568 (N_11568,N_10352,N_10487);
nand U11569 (N_11569,N_10049,N_10831);
or U11570 (N_11570,N_10470,N_10174);
nor U11571 (N_11571,N_10118,N_10270);
or U11572 (N_11572,N_10523,N_10585);
or U11573 (N_11573,N_10495,N_10261);
or U11574 (N_11574,N_10840,N_10458);
nand U11575 (N_11575,N_10442,N_10890);
xor U11576 (N_11576,N_10394,N_10278);
and U11577 (N_11577,N_10237,N_10336);
or U11578 (N_11578,N_10039,N_10374);
or U11579 (N_11579,N_10725,N_10020);
xor U11580 (N_11580,N_10181,N_10036);
and U11581 (N_11581,N_10468,N_10495);
nand U11582 (N_11582,N_10201,N_10435);
and U11583 (N_11583,N_10258,N_10560);
nand U11584 (N_11584,N_10298,N_10752);
nor U11585 (N_11585,N_10713,N_10795);
and U11586 (N_11586,N_10173,N_10134);
and U11587 (N_11587,N_10896,N_10806);
nor U11588 (N_11588,N_10464,N_10620);
and U11589 (N_11589,N_10081,N_10880);
and U11590 (N_11590,N_10344,N_10570);
nor U11591 (N_11591,N_10128,N_10014);
or U11592 (N_11592,N_10364,N_10859);
and U11593 (N_11593,N_10752,N_10930);
nor U11594 (N_11594,N_10799,N_10586);
nor U11595 (N_11595,N_10201,N_10266);
nand U11596 (N_11596,N_10582,N_10603);
xor U11597 (N_11597,N_10642,N_10606);
nor U11598 (N_11598,N_10982,N_10055);
or U11599 (N_11599,N_10449,N_10379);
or U11600 (N_11600,N_10429,N_10254);
or U11601 (N_11601,N_10385,N_10718);
or U11602 (N_11602,N_10236,N_10079);
or U11603 (N_11603,N_10361,N_10896);
nand U11604 (N_11604,N_10468,N_10349);
nand U11605 (N_11605,N_10509,N_10721);
nor U11606 (N_11606,N_10852,N_10295);
nand U11607 (N_11607,N_10698,N_10987);
or U11608 (N_11608,N_10448,N_10876);
and U11609 (N_11609,N_10013,N_10949);
or U11610 (N_11610,N_10407,N_10928);
and U11611 (N_11611,N_10767,N_10157);
and U11612 (N_11612,N_10978,N_10747);
or U11613 (N_11613,N_10458,N_10875);
nand U11614 (N_11614,N_10797,N_10547);
nor U11615 (N_11615,N_10400,N_10323);
nor U11616 (N_11616,N_10378,N_10250);
and U11617 (N_11617,N_10886,N_10904);
xnor U11618 (N_11618,N_10885,N_10595);
xnor U11619 (N_11619,N_10716,N_10410);
nand U11620 (N_11620,N_10210,N_10187);
nor U11621 (N_11621,N_10291,N_10762);
or U11622 (N_11622,N_10919,N_10050);
or U11623 (N_11623,N_10998,N_10657);
nand U11624 (N_11624,N_10550,N_10029);
or U11625 (N_11625,N_10043,N_10932);
and U11626 (N_11626,N_10914,N_10279);
or U11627 (N_11627,N_10375,N_10947);
nor U11628 (N_11628,N_10829,N_10246);
or U11629 (N_11629,N_10719,N_10897);
nor U11630 (N_11630,N_10337,N_10665);
or U11631 (N_11631,N_10873,N_10534);
and U11632 (N_11632,N_10711,N_10820);
nand U11633 (N_11633,N_10620,N_10993);
nor U11634 (N_11634,N_10952,N_10440);
nand U11635 (N_11635,N_10666,N_10502);
or U11636 (N_11636,N_10560,N_10462);
nor U11637 (N_11637,N_10436,N_10177);
nand U11638 (N_11638,N_10949,N_10231);
or U11639 (N_11639,N_10851,N_10912);
nor U11640 (N_11640,N_10080,N_10081);
nor U11641 (N_11641,N_10660,N_10104);
nand U11642 (N_11642,N_10684,N_10149);
or U11643 (N_11643,N_10237,N_10034);
nor U11644 (N_11644,N_10548,N_10049);
nand U11645 (N_11645,N_10616,N_10821);
or U11646 (N_11646,N_10105,N_10978);
nor U11647 (N_11647,N_10853,N_10597);
nand U11648 (N_11648,N_10476,N_10267);
or U11649 (N_11649,N_10175,N_10497);
and U11650 (N_11650,N_10387,N_10338);
and U11651 (N_11651,N_10499,N_10934);
and U11652 (N_11652,N_10907,N_10722);
nand U11653 (N_11653,N_10888,N_10140);
nor U11654 (N_11654,N_10128,N_10438);
and U11655 (N_11655,N_10692,N_10700);
nor U11656 (N_11656,N_10113,N_10227);
or U11657 (N_11657,N_10092,N_10658);
nor U11658 (N_11658,N_10331,N_10262);
and U11659 (N_11659,N_10667,N_10027);
xnor U11660 (N_11660,N_10515,N_10935);
and U11661 (N_11661,N_10509,N_10675);
nand U11662 (N_11662,N_10919,N_10046);
or U11663 (N_11663,N_10436,N_10798);
nor U11664 (N_11664,N_10657,N_10491);
nand U11665 (N_11665,N_10826,N_10936);
and U11666 (N_11666,N_10200,N_10060);
nand U11667 (N_11667,N_10184,N_10309);
nand U11668 (N_11668,N_10839,N_10506);
or U11669 (N_11669,N_10206,N_10173);
or U11670 (N_11670,N_10992,N_10028);
nand U11671 (N_11671,N_10039,N_10539);
or U11672 (N_11672,N_10986,N_10507);
or U11673 (N_11673,N_10043,N_10058);
nand U11674 (N_11674,N_10149,N_10895);
xor U11675 (N_11675,N_10380,N_10644);
nand U11676 (N_11676,N_10158,N_10952);
and U11677 (N_11677,N_10298,N_10445);
and U11678 (N_11678,N_10005,N_10737);
nand U11679 (N_11679,N_10283,N_10707);
nor U11680 (N_11680,N_10861,N_10052);
nand U11681 (N_11681,N_10212,N_10904);
nor U11682 (N_11682,N_10301,N_10092);
nand U11683 (N_11683,N_10375,N_10401);
nor U11684 (N_11684,N_10614,N_10461);
nor U11685 (N_11685,N_10791,N_10195);
nor U11686 (N_11686,N_10014,N_10277);
and U11687 (N_11687,N_10330,N_10106);
nor U11688 (N_11688,N_10734,N_10017);
xnor U11689 (N_11689,N_10748,N_10545);
nand U11690 (N_11690,N_10950,N_10938);
nand U11691 (N_11691,N_10930,N_10251);
or U11692 (N_11692,N_10524,N_10526);
or U11693 (N_11693,N_10500,N_10965);
nor U11694 (N_11694,N_10715,N_10781);
or U11695 (N_11695,N_10019,N_10269);
nor U11696 (N_11696,N_10553,N_10252);
and U11697 (N_11697,N_10226,N_10130);
nand U11698 (N_11698,N_10945,N_10079);
nor U11699 (N_11699,N_10704,N_10154);
xor U11700 (N_11700,N_10108,N_10812);
xor U11701 (N_11701,N_10713,N_10005);
and U11702 (N_11702,N_10588,N_10486);
or U11703 (N_11703,N_10248,N_10854);
and U11704 (N_11704,N_10667,N_10188);
nand U11705 (N_11705,N_10333,N_10794);
and U11706 (N_11706,N_10170,N_10906);
and U11707 (N_11707,N_10287,N_10771);
nor U11708 (N_11708,N_10185,N_10250);
nor U11709 (N_11709,N_10188,N_10102);
and U11710 (N_11710,N_10538,N_10014);
or U11711 (N_11711,N_10254,N_10549);
nand U11712 (N_11712,N_10713,N_10583);
and U11713 (N_11713,N_10288,N_10990);
nand U11714 (N_11714,N_10323,N_10689);
xor U11715 (N_11715,N_10921,N_10964);
nor U11716 (N_11716,N_10134,N_10684);
nand U11717 (N_11717,N_10527,N_10196);
nor U11718 (N_11718,N_10031,N_10860);
nand U11719 (N_11719,N_10881,N_10732);
nor U11720 (N_11720,N_10711,N_10181);
or U11721 (N_11721,N_10453,N_10094);
and U11722 (N_11722,N_10944,N_10818);
nor U11723 (N_11723,N_10807,N_10203);
xnor U11724 (N_11724,N_10818,N_10022);
xor U11725 (N_11725,N_10986,N_10269);
xnor U11726 (N_11726,N_10758,N_10888);
or U11727 (N_11727,N_10927,N_10908);
nor U11728 (N_11728,N_10028,N_10795);
nand U11729 (N_11729,N_10361,N_10224);
nand U11730 (N_11730,N_10063,N_10059);
and U11731 (N_11731,N_10178,N_10033);
nor U11732 (N_11732,N_10528,N_10813);
xor U11733 (N_11733,N_10301,N_10273);
nand U11734 (N_11734,N_10250,N_10107);
or U11735 (N_11735,N_10778,N_10753);
xor U11736 (N_11736,N_10473,N_10178);
nor U11737 (N_11737,N_10424,N_10104);
or U11738 (N_11738,N_10340,N_10017);
or U11739 (N_11739,N_10407,N_10024);
or U11740 (N_11740,N_10862,N_10214);
and U11741 (N_11741,N_10706,N_10121);
xnor U11742 (N_11742,N_10625,N_10928);
nor U11743 (N_11743,N_10053,N_10002);
nor U11744 (N_11744,N_10521,N_10316);
nand U11745 (N_11745,N_10779,N_10095);
or U11746 (N_11746,N_10003,N_10146);
and U11747 (N_11747,N_10423,N_10089);
and U11748 (N_11748,N_10924,N_10989);
nor U11749 (N_11749,N_10261,N_10275);
or U11750 (N_11750,N_10442,N_10990);
and U11751 (N_11751,N_10497,N_10207);
and U11752 (N_11752,N_10667,N_10373);
or U11753 (N_11753,N_10702,N_10392);
nor U11754 (N_11754,N_10145,N_10071);
nor U11755 (N_11755,N_10533,N_10810);
and U11756 (N_11756,N_10406,N_10943);
nand U11757 (N_11757,N_10506,N_10932);
or U11758 (N_11758,N_10257,N_10057);
or U11759 (N_11759,N_10934,N_10337);
nand U11760 (N_11760,N_10278,N_10743);
or U11761 (N_11761,N_10361,N_10769);
nor U11762 (N_11762,N_10768,N_10390);
or U11763 (N_11763,N_10664,N_10747);
xor U11764 (N_11764,N_10454,N_10841);
and U11765 (N_11765,N_10971,N_10001);
nor U11766 (N_11766,N_10227,N_10725);
or U11767 (N_11767,N_10373,N_10281);
or U11768 (N_11768,N_10396,N_10176);
xnor U11769 (N_11769,N_10100,N_10454);
nand U11770 (N_11770,N_10918,N_10115);
nor U11771 (N_11771,N_10212,N_10167);
nor U11772 (N_11772,N_10234,N_10757);
nor U11773 (N_11773,N_10987,N_10413);
or U11774 (N_11774,N_10628,N_10641);
nor U11775 (N_11775,N_10460,N_10138);
and U11776 (N_11776,N_10109,N_10717);
nand U11777 (N_11777,N_10668,N_10561);
nor U11778 (N_11778,N_10435,N_10377);
or U11779 (N_11779,N_10379,N_10002);
and U11780 (N_11780,N_10057,N_10414);
and U11781 (N_11781,N_10667,N_10409);
nor U11782 (N_11782,N_10463,N_10513);
and U11783 (N_11783,N_10210,N_10713);
or U11784 (N_11784,N_10404,N_10837);
nand U11785 (N_11785,N_10810,N_10527);
xnor U11786 (N_11786,N_10696,N_10674);
nand U11787 (N_11787,N_10458,N_10491);
nand U11788 (N_11788,N_10650,N_10874);
nor U11789 (N_11789,N_10013,N_10434);
nor U11790 (N_11790,N_10647,N_10011);
xnor U11791 (N_11791,N_10300,N_10127);
or U11792 (N_11792,N_10104,N_10784);
xnor U11793 (N_11793,N_10716,N_10658);
and U11794 (N_11794,N_10288,N_10777);
or U11795 (N_11795,N_10169,N_10228);
or U11796 (N_11796,N_10519,N_10651);
and U11797 (N_11797,N_10422,N_10837);
and U11798 (N_11798,N_10691,N_10564);
nor U11799 (N_11799,N_10737,N_10266);
nand U11800 (N_11800,N_10762,N_10590);
nor U11801 (N_11801,N_10760,N_10883);
and U11802 (N_11802,N_10562,N_10433);
nand U11803 (N_11803,N_10380,N_10676);
xnor U11804 (N_11804,N_10236,N_10644);
xor U11805 (N_11805,N_10553,N_10346);
xor U11806 (N_11806,N_10283,N_10340);
or U11807 (N_11807,N_10863,N_10219);
or U11808 (N_11808,N_10415,N_10614);
nor U11809 (N_11809,N_10534,N_10327);
or U11810 (N_11810,N_10616,N_10120);
xor U11811 (N_11811,N_10573,N_10499);
nand U11812 (N_11812,N_10883,N_10509);
and U11813 (N_11813,N_10862,N_10109);
and U11814 (N_11814,N_10684,N_10482);
nand U11815 (N_11815,N_10502,N_10808);
or U11816 (N_11816,N_10259,N_10601);
or U11817 (N_11817,N_10918,N_10604);
nand U11818 (N_11818,N_10885,N_10527);
nor U11819 (N_11819,N_10030,N_10139);
nor U11820 (N_11820,N_10837,N_10806);
xor U11821 (N_11821,N_10200,N_10161);
xnor U11822 (N_11822,N_10411,N_10815);
or U11823 (N_11823,N_10982,N_10601);
xor U11824 (N_11824,N_10629,N_10908);
or U11825 (N_11825,N_10638,N_10564);
nand U11826 (N_11826,N_10403,N_10276);
nand U11827 (N_11827,N_10316,N_10458);
and U11828 (N_11828,N_10797,N_10901);
nand U11829 (N_11829,N_10872,N_10665);
nand U11830 (N_11830,N_10619,N_10894);
or U11831 (N_11831,N_10720,N_10210);
or U11832 (N_11832,N_10990,N_10247);
and U11833 (N_11833,N_10603,N_10279);
and U11834 (N_11834,N_10314,N_10939);
xor U11835 (N_11835,N_10303,N_10078);
xor U11836 (N_11836,N_10543,N_10579);
nand U11837 (N_11837,N_10433,N_10563);
and U11838 (N_11838,N_10078,N_10216);
nand U11839 (N_11839,N_10065,N_10339);
nand U11840 (N_11840,N_10183,N_10512);
nor U11841 (N_11841,N_10968,N_10514);
nand U11842 (N_11842,N_10957,N_10321);
nor U11843 (N_11843,N_10241,N_10526);
nor U11844 (N_11844,N_10244,N_10687);
nand U11845 (N_11845,N_10536,N_10577);
xnor U11846 (N_11846,N_10478,N_10952);
xor U11847 (N_11847,N_10378,N_10737);
nand U11848 (N_11848,N_10609,N_10839);
or U11849 (N_11849,N_10827,N_10109);
or U11850 (N_11850,N_10377,N_10325);
or U11851 (N_11851,N_10810,N_10847);
nand U11852 (N_11852,N_10505,N_10909);
nor U11853 (N_11853,N_10546,N_10379);
nor U11854 (N_11854,N_10325,N_10980);
nor U11855 (N_11855,N_10180,N_10826);
or U11856 (N_11856,N_10323,N_10916);
or U11857 (N_11857,N_10569,N_10776);
nor U11858 (N_11858,N_10422,N_10709);
or U11859 (N_11859,N_10927,N_10789);
nor U11860 (N_11860,N_10205,N_10200);
nor U11861 (N_11861,N_10240,N_10102);
nor U11862 (N_11862,N_10659,N_10630);
or U11863 (N_11863,N_10072,N_10764);
and U11864 (N_11864,N_10208,N_10108);
xnor U11865 (N_11865,N_10127,N_10642);
nand U11866 (N_11866,N_10648,N_10838);
or U11867 (N_11867,N_10181,N_10895);
and U11868 (N_11868,N_10544,N_10647);
or U11869 (N_11869,N_10155,N_10418);
and U11870 (N_11870,N_10807,N_10986);
nor U11871 (N_11871,N_10536,N_10604);
or U11872 (N_11872,N_10391,N_10811);
or U11873 (N_11873,N_10037,N_10760);
nor U11874 (N_11874,N_10590,N_10324);
nor U11875 (N_11875,N_10092,N_10852);
and U11876 (N_11876,N_10988,N_10549);
or U11877 (N_11877,N_10241,N_10907);
nor U11878 (N_11878,N_10281,N_10925);
nand U11879 (N_11879,N_10986,N_10139);
nor U11880 (N_11880,N_10605,N_10153);
or U11881 (N_11881,N_10358,N_10870);
nor U11882 (N_11882,N_10067,N_10215);
nor U11883 (N_11883,N_10648,N_10474);
or U11884 (N_11884,N_10460,N_10524);
or U11885 (N_11885,N_10805,N_10768);
nand U11886 (N_11886,N_10570,N_10746);
and U11887 (N_11887,N_10855,N_10407);
nor U11888 (N_11888,N_10898,N_10559);
nor U11889 (N_11889,N_10405,N_10615);
nand U11890 (N_11890,N_10627,N_10322);
and U11891 (N_11891,N_10840,N_10003);
or U11892 (N_11892,N_10555,N_10905);
nand U11893 (N_11893,N_10213,N_10478);
nand U11894 (N_11894,N_10689,N_10276);
nor U11895 (N_11895,N_10625,N_10612);
xor U11896 (N_11896,N_10184,N_10287);
and U11897 (N_11897,N_10620,N_10296);
and U11898 (N_11898,N_10137,N_10177);
or U11899 (N_11899,N_10264,N_10845);
and U11900 (N_11900,N_10893,N_10204);
or U11901 (N_11901,N_10993,N_10073);
and U11902 (N_11902,N_10752,N_10259);
nor U11903 (N_11903,N_10995,N_10516);
nand U11904 (N_11904,N_10129,N_10554);
and U11905 (N_11905,N_10746,N_10400);
nor U11906 (N_11906,N_10422,N_10077);
nand U11907 (N_11907,N_10228,N_10059);
nand U11908 (N_11908,N_10817,N_10961);
nand U11909 (N_11909,N_10959,N_10689);
nor U11910 (N_11910,N_10757,N_10572);
nand U11911 (N_11911,N_10914,N_10580);
and U11912 (N_11912,N_10155,N_10841);
nand U11913 (N_11913,N_10028,N_10730);
and U11914 (N_11914,N_10571,N_10668);
xor U11915 (N_11915,N_10435,N_10621);
xor U11916 (N_11916,N_10497,N_10908);
nand U11917 (N_11917,N_10704,N_10581);
nand U11918 (N_11918,N_10088,N_10078);
and U11919 (N_11919,N_10838,N_10382);
nor U11920 (N_11920,N_10104,N_10252);
nand U11921 (N_11921,N_10035,N_10144);
and U11922 (N_11922,N_10705,N_10375);
or U11923 (N_11923,N_10884,N_10576);
or U11924 (N_11924,N_10178,N_10164);
or U11925 (N_11925,N_10636,N_10374);
or U11926 (N_11926,N_10029,N_10825);
nor U11927 (N_11927,N_10086,N_10451);
nor U11928 (N_11928,N_10587,N_10063);
and U11929 (N_11929,N_10198,N_10886);
or U11930 (N_11930,N_10617,N_10033);
nor U11931 (N_11931,N_10015,N_10859);
xnor U11932 (N_11932,N_10708,N_10573);
nand U11933 (N_11933,N_10253,N_10156);
and U11934 (N_11934,N_10827,N_10580);
nand U11935 (N_11935,N_10076,N_10470);
nand U11936 (N_11936,N_10923,N_10170);
or U11937 (N_11937,N_10893,N_10323);
and U11938 (N_11938,N_10373,N_10349);
and U11939 (N_11939,N_10096,N_10538);
and U11940 (N_11940,N_10295,N_10123);
nand U11941 (N_11941,N_10489,N_10889);
nand U11942 (N_11942,N_10304,N_10008);
nor U11943 (N_11943,N_10986,N_10597);
and U11944 (N_11944,N_10664,N_10391);
nor U11945 (N_11945,N_10932,N_10656);
and U11946 (N_11946,N_10655,N_10434);
or U11947 (N_11947,N_10729,N_10680);
nor U11948 (N_11948,N_10410,N_10053);
nand U11949 (N_11949,N_10581,N_10925);
or U11950 (N_11950,N_10341,N_10280);
or U11951 (N_11951,N_10058,N_10921);
and U11952 (N_11952,N_10350,N_10549);
nor U11953 (N_11953,N_10601,N_10022);
or U11954 (N_11954,N_10539,N_10486);
nor U11955 (N_11955,N_10664,N_10653);
or U11956 (N_11956,N_10440,N_10114);
or U11957 (N_11957,N_10591,N_10211);
nor U11958 (N_11958,N_10674,N_10357);
or U11959 (N_11959,N_10936,N_10910);
nor U11960 (N_11960,N_10066,N_10346);
nor U11961 (N_11961,N_10908,N_10107);
xnor U11962 (N_11962,N_10255,N_10413);
nand U11963 (N_11963,N_10339,N_10037);
nor U11964 (N_11964,N_10861,N_10362);
and U11965 (N_11965,N_10830,N_10959);
nor U11966 (N_11966,N_10243,N_10429);
nor U11967 (N_11967,N_10244,N_10150);
and U11968 (N_11968,N_10573,N_10732);
nand U11969 (N_11969,N_10143,N_10614);
and U11970 (N_11970,N_10006,N_10391);
and U11971 (N_11971,N_10444,N_10003);
xnor U11972 (N_11972,N_10638,N_10968);
nand U11973 (N_11973,N_10328,N_10638);
or U11974 (N_11974,N_10320,N_10440);
or U11975 (N_11975,N_10631,N_10480);
nor U11976 (N_11976,N_10794,N_10353);
and U11977 (N_11977,N_10722,N_10830);
or U11978 (N_11978,N_10600,N_10496);
nor U11979 (N_11979,N_10015,N_10695);
or U11980 (N_11980,N_10667,N_10104);
and U11981 (N_11981,N_10237,N_10667);
or U11982 (N_11982,N_10597,N_10935);
or U11983 (N_11983,N_10668,N_10497);
nand U11984 (N_11984,N_10741,N_10538);
nand U11985 (N_11985,N_10059,N_10916);
nor U11986 (N_11986,N_10404,N_10970);
and U11987 (N_11987,N_10737,N_10884);
nand U11988 (N_11988,N_10760,N_10820);
nor U11989 (N_11989,N_10563,N_10592);
or U11990 (N_11990,N_10392,N_10202);
and U11991 (N_11991,N_10406,N_10851);
nor U11992 (N_11992,N_10189,N_10901);
xnor U11993 (N_11993,N_10693,N_10349);
nor U11994 (N_11994,N_10647,N_10581);
nor U11995 (N_11995,N_10675,N_10315);
nor U11996 (N_11996,N_10102,N_10223);
or U11997 (N_11997,N_10078,N_10420);
nand U11998 (N_11998,N_10004,N_10259);
and U11999 (N_11999,N_10165,N_10380);
xor U12000 (N_12000,N_11533,N_11656);
and U12001 (N_12001,N_11760,N_11486);
nor U12002 (N_12002,N_11095,N_11127);
nor U12003 (N_12003,N_11988,N_11493);
or U12004 (N_12004,N_11488,N_11061);
nor U12005 (N_12005,N_11932,N_11016);
nor U12006 (N_12006,N_11597,N_11151);
nor U12007 (N_12007,N_11429,N_11200);
nand U12008 (N_12008,N_11909,N_11706);
and U12009 (N_12009,N_11783,N_11096);
and U12010 (N_12010,N_11718,N_11693);
and U12011 (N_12011,N_11641,N_11337);
and U12012 (N_12012,N_11088,N_11809);
and U12013 (N_12013,N_11444,N_11619);
or U12014 (N_12014,N_11567,N_11307);
or U12015 (N_12015,N_11209,N_11997);
nor U12016 (N_12016,N_11038,N_11058);
or U12017 (N_12017,N_11366,N_11328);
or U12018 (N_12018,N_11230,N_11348);
and U12019 (N_12019,N_11880,N_11271);
xor U12020 (N_12020,N_11412,N_11859);
nor U12021 (N_12021,N_11196,N_11367);
nor U12022 (N_12022,N_11144,N_11379);
or U12023 (N_12023,N_11084,N_11423);
nor U12024 (N_12024,N_11319,N_11664);
nand U12025 (N_12025,N_11150,N_11229);
and U12026 (N_12026,N_11466,N_11532);
nand U12027 (N_12027,N_11278,N_11076);
nor U12028 (N_12028,N_11382,N_11138);
xor U12029 (N_12029,N_11836,N_11164);
nor U12030 (N_12030,N_11049,N_11373);
and U12031 (N_12031,N_11947,N_11945);
nand U12032 (N_12032,N_11637,N_11985);
nor U12033 (N_12033,N_11601,N_11147);
xnor U12034 (N_12034,N_11941,N_11006);
nor U12035 (N_12035,N_11251,N_11030);
or U12036 (N_12036,N_11413,N_11811);
nor U12037 (N_12037,N_11161,N_11701);
and U12038 (N_12038,N_11329,N_11846);
and U12039 (N_12039,N_11370,N_11876);
and U12040 (N_12040,N_11363,N_11600);
nand U12041 (N_12041,N_11044,N_11132);
or U12042 (N_12042,N_11331,N_11757);
nor U12043 (N_12043,N_11079,N_11008);
nor U12044 (N_12044,N_11820,N_11626);
and U12045 (N_12045,N_11697,N_11189);
and U12046 (N_12046,N_11046,N_11910);
or U12047 (N_12047,N_11677,N_11216);
or U12048 (N_12048,N_11159,N_11724);
and U12049 (N_12049,N_11395,N_11793);
nand U12050 (N_12050,N_11901,N_11220);
nand U12051 (N_12051,N_11661,N_11123);
and U12052 (N_12052,N_11145,N_11416);
nor U12053 (N_12053,N_11443,N_11921);
nand U12054 (N_12054,N_11628,N_11037);
or U12055 (N_12055,N_11835,N_11935);
nand U12056 (N_12056,N_11447,N_11696);
nand U12057 (N_12057,N_11440,N_11420);
nor U12058 (N_12058,N_11344,N_11356);
nor U12059 (N_12059,N_11109,N_11093);
nand U12060 (N_12060,N_11173,N_11680);
nor U12061 (N_12061,N_11430,N_11971);
and U12062 (N_12062,N_11998,N_11911);
nor U12063 (N_12063,N_11678,N_11224);
or U12064 (N_12064,N_11866,N_11133);
and U12065 (N_12065,N_11618,N_11643);
xnor U12066 (N_12066,N_11839,N_11769);
nor U12067 (N_12067,N_11290,N_11804);
nand U12068 (N_12068,N_11943,N_11075);
or U12069 (N_12069,N_11270,N_11887);
nand U12070 (N_12070,N_11891,N_11338);
or U12071 (N_12071,N_11474,N_11591);
nor U12072 (N_12072,N_11882,N_11540);
and U12073 (N_12073,N_11573,N_11512);
or U12074 (N_12074,N_11436,N_11824);
xnor U12075 (N_12075,N_11286,N_11722);
nor U12076 (N_12076,N_11665,N_11993);
nor U12077 (N_12077,N_11915,N_11020);
and U12078 (N_12078,N_11865,N_11396);
nor U12079 (N_12079,N_11875,N_11136);
nand U12080 (N_12080,N_11203,N_11922);
nor U12081 (N_12081,N_11742,N_11633);
and U12082 (N_12082,N_11130,N_11924);
or U12083 (N_12083,N_11148,N_11146);
nand U12084 (N_12084,N_11113,N_11383);
xor U12085 (N_12085,N_11424,N_11794);
and U12086 (N_12086,N_11013,N_11798);
nand U12087 (N_12087,N_11640,N_11106);
and U12088 (N_12088,N_11805,N_11566);
or U12089 (N_12089,N_11776,N_11105);
nand U12090 (N_12090,N_11761,N_11828);
and U12091 (N_12091,N_11978,N_11931);
nand U12092 (N_12092,N_11647,N_11874);
nand U12093 (N_12093,N_11873,N_11381);
and U12094 (N_12094,N_11631,N_11558);
xnor U12095 (N_12095,N_11180,N_11861);
nand U12096 (N_12096,N_11260,N_11497);
or U12097 (N_12097,N_11767,N_11187);
nand U12098 (N_12098,N_11682,N_11245);
nor U12099 (N_12099,N_11923,N_11546);
nand U12100 (N_12100,N_11670,N_11895);
xor U12101 (N_12101,N_11578,N_11545);
and U12102 (N_12102,N_11306,N_11314);
nor U12103 (N_12103,N_11082,N_11362);
nor U12104 (N_12104,N_11575,N_11483);
and U12105 (N_12105,N_11397,N_11855);
nor U12106 (N_12106,N_11886,N_11465);
xnor U12107 (N_12107,N_11730,N_11142);
nand U12108 (N_12108,N_11221,N_11199);
or U12109 (N_12109,N_11459,N_11639);
or U12110 (N_12110,N_11283,N_11360);
or U12111 (N_12111,N_11428,N_11657);
nand U12112 (N_12112,N_11983,N_11871);
or U12113 (N_12113,N_11791,N_11154);
nor U12114 (N_12114,N_11893,N_11821);
nand U12115 (N_12115,N_11765,N_11115);
and U12116 (N_12116,N_11916,N_11606);
nand U12117 (N_12117,N_11070,N_11490);
and U12118 (N_12118,N_11559,N_11713);
nand U12119 (N_12119,N_11375,N_11234);
or U12120 (N_12120,N_11255,N_11374);
nand U12121 (N_12121,N_11691,N_11040);
and U12122 (N_12122,N_11389,N_11981);
or U12123 (N_12123,N_11334,N_11748);
or U12124 (N_12124,N_11499,N_11045);
xnor U12125 (N_12125,N_11295,N_11966);
nand U12126 (N_12126,N_11257,N_11913);
nand U12127 (N_12127,N_11675,N_11621);
or U12128 (N_12128,N_11226,N_11433);
nor U12129 (N_12129,N_11128,N_11725);
nor U12130 (N_12130,N_11303,N_11609);
nand U12131 (N_12131,N_11312,N_11168);
nand U12132 (N_12132,N_11071,N_11946);
and U12133 (N_12133,N_11894,N_11974);
and U12134 (N_12134,N_11027,N_11408);
and U12135 (N_12135,N_11717,N_11349);
xor U12136 (N_12136,N_11309,N_11059);
nor U12137 (N_12137,N_11281,N_11788);
nor U12138 (N_12138,N_11250,N_11405);
and U12139 (N_12139,N_11651,N_11970);
nor U12140 (N_12140,N_11995,N_11852);
or U12141 (N_12141,N_11249,N_11077);
or U12142 (N_12142,N_11623,N_11014);
xor U12143 (N_12143,N_11755,N_11456);
and U12144 (N_12144,N_11743,N_11376);
nand U12145 (N_12145,N_11962,N_11979);
or U12146 (N_12146,N_11509,N_11228);
nand U12147 (N_12147,N_11720,N_11799);
or U12148 (N_12148,N_11273,N_11065);
and U12149 (N_12149,N_11442,N_11646);
nand U12150 (N_12150,N_11476,N_11984);
nand U12151 (N_12151,N_11241,N_11630);
nand U12152 (N_12152,N_11026,N_11043);
or U12153 (N_12153,N_11425,N_11683);
nor U12154 (N_12154,N_11638,N_11898);
or U12155 (N_12155,N_11118,N_11515);
or U12156 (N_12156,N_11684,N_11751);
nand U12157 (N_12157,N_11243,N_11564);
nor U12158 (N_12158,N_11897,N_11291);
and U12159 (N_12159,N_11489,N_11523);
nand U12160 (N_12160,N_11698,N_11218);
nand U12161 (N_12161,N_11634,N_11977);
and U12162 (N_12162,N_11569,N_11885);
nor U12163 (N_12163,N_11137,N_11345);
nand U12164 (N_12164,N_11908,N_11458);
or U12165 (N_12165,N_11192,N_11426);
and U12166 (N_12166,N_11587,N_11299);
and U12167 (N_12167,N_11529,N_11169);
nand U12168 (N_12168,N_11032,N_11053);
nor U12169 (N_12169,N_11590,N_11593);
nand U12170 (N_12170,N_11961,N_11134);
nand U12171 (N_12171,N_11510,N_11400);
or U12172 (N_12172,N_11479,N_11942);
and U12173 (N_12173,N_11266,N_11611);
or U12174 (N_12174,N_11632,N_11949);
nor U12175 (N_12175,N_11581,N_11589);
nor U12176 (N_12176,N_11481,N_11103);
xnor U12177 (N_12177,N_11104,N_11500);
nor U12178 (N_12178,N_11948,N_11539);
or U12179 (N_12179,N_11627,N_11726);
or U12180 (N_12180,N_11141,N_11648);
nand U12181 (N_12181,N_11193,N_11582);
nor U12182 (N_12182,N_11156,N_11881);
xnor U12183 (N_12183,N_11789,N_11610);
nand U12184 (N_12184,N_11064,N_11108);
nor U12185 (N_12185,N_11845,N_11603);
nand U12186 (N_12186,N_11553,N_11732);
nor U12187 (N_12187,N_11750,N_11004);
nor U12188 (N_12188,N_11853,N_11555);
nand U12189 (N_12189,N_11432,N_11666);
or U12190 (N_12190,N_11153,N_11635);
nand U12191 (N_12191,N_11892,N_11779);
nand U12192 (N_12192,N_11129,N_11222);
nor U12193 (N_12193,N_11987,N_11676);
nor U12194 (N_12194,N_11741,N_11302);
nor U12195 (N_12195,N_11517,N_11749);
xnor U12196 (N_12196,N_11120,N_11066);
xnor U12197 (N_12197,N_11073,N_11326);
or U12198 (N_12198,N_11736,N_11506);
nor U12199 (N_12199,N_11803,N_11364);
or U12200 (N_12200,N_11808,N_11048);
or U12201 (N_12201,N_11832,N_11354);
nor U12202 (N_12202,N_11796,N_11795);
or U12203 (N_12203,N_11175,N_11311);
and U12204 (N_12204,N_11502,N_11386);
or U12205 (N_12205,N_11361,N_11300);
nor U12206 (N_12206,N_11957,N_11936);
nand U12207 (N_12207,N_11797,N_11090);
nor U12208 (N_12208,N_11872,N_11912);
nand U12209 (N_12209,N_11588,N_11878);
and U12210 (N_12210,N_11455,N_11178);
and U12211 (N_12211,N_11403,N_11800);
nand U12212 (N_12212,N_11191,N_11181);
or U12213 (N_12213,N_11507,N_11658);
xor U12214 (N_12214,N_11900,N_11771);
or U12215 (N_12215,N_11530,N_11205);
and U12216 (N_12216,N_11155,N_11359);
and U12217 (N_12217,N_11157,N_11753);
or U12218 (N_12218,N_11541,N_11078);
nand U12219 (N_12219,N_11663,N_11484);
xnor U12220 (N_12220,N_11451,N_11737);
nand U12221 (N_12221,N_11904,N_11607);
nand U12222 (N_12222,N_11340,N_11116);
or U12223 (N_12223,N_11653,N_11491);
or U12224 (N_12224,N_11111,N_11525);
nor U12225 (N_12225,N_11527,N_11210);
or U12226 (N_12226,N_11819,N_11215);
and U12227 (N_12227,N_11940,N_11131);
nand U12228 (N_12228,N_11369,N_11034);
nand U12229 (N_12229,N_11959,N_11399);
nor U12230 (N_12230,N_11446,N_11518);
and U12231 (N_12231,N_11327,N_11163);
xor U12232 (N_12232,N_11135,N_11204);
or U12233 (N_12233,N_11551,N_11960);
nor U12234 (N_12234,N_11896,N_11568);
xnor U12235 (N_12235,N_11785,N_11469);
and U12236 (N_12236,N_11035,N_11087);
or U12237 (N_12237,N_11033,N_11160);
nor U12238 (N_12238,N_11669,N_11315);
and U12239 (N_12239,N_11398,N_11801);
or U12240 (N_12240,N_11528,N_11232);
and U12241 (N_12241,N_11535,N_11263);
xnor U12242 (N_12242,N_11010,N_11950);
or U12243 (N_12243,N_11877,N_11615);
nor U12244 (N_12244,N_11256,N_11671);
and U12245 (N_12245,N_11667,N_11705);
and U12246 (N_12246,N_11213,N_11051);
or U12247 (N_12247,N_11023,N_11715);
or U12248 (N_12248,N_11752,N_11831);
nor U12249 (N_12249,N_11316,N_11025);
and U12250 (N_12250,N_11919,N_11235);
or U12251 (N_12251,N_11171,N_11384);
nand U12252 (N_12252,N_11738,N_11417);
xor U12253 (N_12253,N_11511,N_11332);
xnor U12254 (N_12254,N_11339,N_11850);
xnor U12255 (N_12255,N_11437,N_11028);
xor U12256 (N_12256,N_11052,N_11834);
nand U12257 (N_12257,N_11143,N_11091);
and U12258 (N_12258,N_11351,N_11790);
or U12259 (N_12259,N_11862,N_11556);
and U12260 (N_12260,N_11847,N_11787);
xnor U12261 (N_12261,N_11268,N_11390);
or U12262 (N_12262,N_11756,N_11099);
and U12263 (N_12263,N_11557,N_11662);
or U12264 (N_12264,N_11700,N_11195);
and U12265 (N_12265,N_11461,N_11907);
nand U12266 (N_12266,N_11057,N_11542);
nor U12267 (N_12267,N_11259,N_11728);
nand U12268 (N_12268,N_11172,N_11094);
and U12269 (N_12269,N_11242,N_11325);
nor U12270 (N_12270,N_11297,N_11547);
nand U12271 (N_12271,N_11584,N_11604);
or U12272 (N_12272,N_11644,N_11121);
or U12273 (N_12273,N_11980,N_11264);
and U12274 (N_12274,N_11560,N_11454);
xor U12275 (N_12275,N_11571,N_11524);
nand U12276 (N_12276,N_11284,N_11577);
or U12277 (N_12277,N_11650,N_11237);
and U12278 (N_12278,N_11183,N_11434);
or U12279 (N_12279,N_11830,N_11357);
and U12280 (N_12280,N_11421,N_11955);
and U12281 (N_12281,N_11543,N_11276);
nor U12282 (N_12282,N_11703,N_11406);
xor U12283 (N_12283,N_11007,N_11414);
or U12284 (N_12284,N_11176,N_11239);
nand U12285 (N_12285,N_11544,N_11704);
nor U12286 (N_12286,N_11857,N_11746);
nor U12287 (N_12287,N_11925,N_11072);
nor U12288 (N_12288,N_11687,N_11478);
nor U12289 (N_12289,N_11672,N_11485);
or U12290 (N_12290,N_11906,N_11179);
nand U12291 (N_12291,N_11758,N_11652);
nand U12292 (N_12292,N_11762,N_11184);
or U12293 (N_12293,N_11822,N_11620);
and U12294 (N_12294,N_11402,N_11009);
or U12295 (N_12295,N_11448,N_11692);
and U12296 (N_12296,N_11233,N_11838);
xnor U12297 (N_12297,N_11534,N_11177);
or U12298 (N_12298,N_11438,N_11505);
nor U12299 (N_12299,N_11770,N_11343);
nand U12300 (N_12300,N_11565,N_11688);
xnor U12301 (N_12301,N_11333,N_11280);
nor U12302 (N_12302,N_11735,N_11063);
and U12303 (N_12303,N_11937,N_11825);
or U12304 (N_12304,N_11310,N_11719);
xor U12305 (N_12305,N_11552,N_11659);
nand U12306 (N_12306,N_11868,N_11068);
nor U12307 (N_12307,N_11365,N_11165);
xnor U12308 (N_12308,N_11973,N_11681);
xnor U12309 (N_12309,N_11012,N_11114);
nand U12310 (N_12310,N_11764,N_11371);
and U12311 (N_12311,N_11707,N_11188);
nor U12312 (N_12312,N_11080,N_11214);
xor U12313 (N_12313,N_11645,N_11994);
and U12314 (N_12314,N_11207,N_11807);
and U12315 (N_12315,N_11521,N_11740);
and U12316 (N_12316,N_11201,N_11083);
nand U12317 (N_12317,N_11347,N_11810);
nand U12318 (N_12318,N_11212,N_11914);
or U12319 (N_12319,N_11258,N_11392);
or U12320 (N_12320,N_11335,N_11102);
or U12321 (N_12321,N_11225,N_11968);
nand U12322 (N_12322,N_11554,N_11453);
and U12323 (N_12323,N_11689,N_11269);
nand U12324 (N_12324,N_11378,N_11975);
nor U12325 (N_12325,N_11990,N_11562);
nor U12326 (N_12326,N_11279,N_11122);
xor U12327 (N_12327,N_11092,N_11733);
and U12328 (N_12328,N_11393,N_11410);
or U12329 (N_12329,N_11902,N_11636);
and U12330 (N_12330,N_11254,N_11470);
and U12331 (N_12331,N_11777,N_11353);
and U12332 (N_12332,N_11001,N_11449);
or U12333 (N_12333,N_11967,N_11890);
nor U12334 (N_12334,N_11464,N_11951);
xnor U12335 (N_12335,N_11827,N_11813);
nand U12336 (N_12336,N_11774,N_11101);
nor U12337 (N_12337,N_11870,N_11323);
or U12338 (N_12338,N_11784,N_11391);
nand U12339 (N_12339,N_11289,N_11206);
nand U12340 (N_12340,N_11842,N_11823);
nand U12341 (N_12341,N_11956,N_11867);
xnor U12342 (N_12342,N_11712,N_11039);
and U12343 (N_12343,N_11586,N_11883);
nor U12344 (N_12344,N_11321,N_11926);
or U12345 (N_12345,N_11576,N_11954);
xor U12346 (N_12346,N_11248,N_11158);
and U12347 (N_12347,N_11198,N_11772);
or U12348 (N_12348,N_11763,N_11240);
nor U12349 (N_12349,N_11537,N_11976);
nand U12350 (N_12350,N_11185,N_11744);
or U12351 (N_12351,N_11431,N_11595);
xnor U12352 (N_12352,N_11388,N_11531);
xnor U12353 (N_12353,N_11654,N_11247);
nand U12354 (N_12354,N_11387,N_11739);
nor U12355 (N_12355,N_11296,N_11503);
nand U12356 (N_12356,N_11152,N_11274);
nand U12357 (N_12357,N_11580,N_11986);
or U12358 (N_12358,N_11814,N_11782);
nor U12359 (N_12359,N_11018,N_11275);
and U12360 (N_12360,N_11298,N_11320);
or U12361 (N_12361,N_11287,N_11294);
or U12362 (N_12362,N_11067,N_11649);
nand U12363 (N_12363,N_11317,N_11494);
nand U12364 (N_12364,N_11526,N_11514);
and U12365 (N_12365,N_11999,N_11686);
xnor U12366 (N_12366,N_11944,N_11100);
nand U12367 (N_12367,N_11538,N_11427);
or U12368 (N_12368,N_11843,N_11081);
xnor U12369 (N_12369,N_11342,N_11612);
or U12370 (N_12370,N_11599,N_11561);
or U12371 (N_12371,N_11170,N_11734);
nand U12372 (N_12372,N_11244,N_11711);
or U12373 (N_12373,N_11404,N_11047);
or U12374 (N_12374,N_11934,N_11322);
nand U12375 (N_12375,N_11419,N_11024);
and U12376 (N_12376,N_11149,N_11000);
xor U12377 (N_12377,N_11731,N_11930);
nand U12378 (N_12378,N_11699,N_11021);
nand U12379 (N_12379,N_11952,N_11826);
nand U12380 (N_12380,N_11265,N_11308);
nor U12381 (N_12381,N_11889,N_11418);
nand U12382 (N_12382,N_11754,N_11655);
nor U12383 (N_12383,N_11679,N_11017);
xor U12384 (N_12384,N_11710,N_11817);
and U12385 (N_12385,N_11938,N_11450);
and U12386 (N_12386,N_11812,N_11267);
or U12387 (N_12387,N_11992,N_11953);
xor U12388 (N_12388,N_11714,N_11112);
and U12389 (N_12389,N_11492,N_11854);
or U12390 (N_12390,N_11837,N_11602);
or U12391 (N_12391,N_11031,N_11721);
or U12392 (N_12392,N_11833,N_11480);
xnor U12393 (N_12393,N_11487,N_11860);
and U12394 (N_12394,N_11140,N_11457);
nor U12395 (N_12395,N_11462,N_11708);
and U12396 (N_12396,N_11802,N_11504);
nand U12397 (N_12397,N_11208,N_11062);
or U12398 (N_12398,N_11252,N_11261);
and U12399 (N_12399,N_11745,N_11330);
nor U12400 (N_12400,N_11508,N_11918);
nor U12401 (N_12401,N_11781,N_11969);
or U12402 (N_12402,N_11253,N_11313);
or U12403 (N_12403,N_11608,N_11227);
xor U12404 (N_12404,N_11996,N_11288);
xnor U12405 (N_12405,N_11928,N_11592);
and U12406 (N_12406,N_11840,N_11549);
or U12407 (N_12407,N_11098,N_11501);
nor U12408 (N_12408,N_11522,N_11864);
nor U12409 (N_12409,N_11879,N_11792);
xnor U12410 (N_12410,N_11238,N_11019);
or U12411 (N_12411,N_11579,N_11965);
nand U12412 (N_12412,N_11614,N_11989);
nand U12413 (N_12413,N_11598,N_11352);
xor U12414 (N_12414,N_11617,N_11211);
nor U12415 (N_12415,N_11848,N_11441);
xor U12416 (N_12416,N_11685,N_11119);
nor U12417 (N_12417,N_11041,N_11629);
nor U12418 (N_12418,N_11729,N_11613);
nand U12419 (N_12419,N_11884,N_11668);
or U12420 (N_12420,N_11415,N_11336);
or U12421 (N_12421,N_11806,N_11888);
nor U12422 (N_12422,N_11085,N_11920);
xnor U12423 (N_12423,N_11460,N_11851);
nor U12424 (N_12424,N_11747,N_11385);
nor U12425 (N_12425,N_11219,N_11574);
nand U12426 (N_12426,N_11060,N_11411);
xnor U12427 (N_12427,N_11816,N_11422);
nor U12428 (N_12428,N_11858,N_11174);
nor U12429 (N_12429,N_11285,N_11162);
nand U12430 (N_12430,N_11126,N_11829);
or U12431 (N_12431,N_11318,N_11394);
nor U12432 (N_12432,N_11572,N_11563);
nor U12433 (N_12433,N_11972,N_11002);
xor U12434 (N_12434,N_11089,N_11818);
nand U12435 (N_12435,N_11759,N_11125);
and U12436 (N_12436,N_11029,N_11022);
and U12437 (N_12437,N_11355,N_11863);
xnor U12438 (N_12438,N_11495,N_11475);
xnor U12439 (N_12439,N_11709,N_11056);
xor U12440 (N_12440,N_11856,N_11054);
nand U12441 (N_12441,N_11358,N_11585);
and U12442 (N_12442,N_11477,N_11292);
nand U12443 (N_12443,N_11766,N_11844);
nor U12444 (N_12444,N_11350,N_11223);
or U12445 (N_12445,N_11439,N_11069);
and U12446 (N_12446,N_11472,N_11482);
nand U12447 (N_12447,N_11786,N_11727);
or U12448 (N_12448,N_11282,N_11695);
and U12449 (N_12449,N_11036,N_11305);
nand U12450 (N_12450,N_11516,N_11377);
xnor U12451 (N_12451,N_11939,N_11217);
nand U12452 (N_12452,N_11991,N_11780);
nor U12453 (N_12453,N_11660,N_11015);
nand U12454 (N_12454,N_11778,N_11380);
nand U12455 (N_12455,N_11272,N_11194);
nor U12456 (N_12456,N_11086,N_11473);
nand U12457 (N_12457,N_11011,N_11074);
or U12458 (N_12458,N_11346,N_11513);
nor U12459 (N_12459,N_11050,N_11042);
nor U12460 (N_12460,N_11167,N_11594);
and U12461 (N_12461,N_11190,N_11139);
nor U12462 (N_12462,N_11236,N_11899);
nor U12463 (N_12463,N_11674,N_11372);
nor U12464 (N_12464,N_11723,N_11231);
nor U12465 (N_12465,N_11815,N_11673);
and U12466 (N_12466,N_11982,N_11202);
or U12467 (N_12467,N_11166,N_11905);
or U12468 (N_12468,N_11548,N_11841);
nand U12469 (N_12469,N_11293,N_11622);
and U12470 (N_12470,N_11596,N_11768);
nor U12471 (N_12471,N_11702,N_11498);
or U12472 (N_12472,N_11583,N_11694);
or U12473 (N_12473,N_11452,N_11401);
nand U12474 (N_12474,N_11903,N_11055);
and U12475 (N_12475,N_11471,N_11642);
xnor U12476 (N_12476,N_11003,N_11107);
nand U12477 (N_12477,N_11775,N_11605);
nor U12478 (N_12478,N_11964,N_11624);
nor U12479 (N_12479,N_11849,N_11929);
nor U12480 (N_12480,N_11616,N_11301);
nor U12481 (N_12481,N_11368,N_11110);
nor U12482 (N_12482,N_11246,N_11445);
and U12483 (N_12483,N_11625,N_11467);
or U12484 (N_12484,N_11182,N_11536);
and U12485 (N_12485,N_11409,N_11570);
nor U12486 (N_12486,N_11716,N_11869);
and U12487 (N_12487,N_11277,N_11690);
nand U12488 (N_12488,N_11186,N_11407);
nand U12489 (N_12489,N_11933,N_11117);
or U12490 (N_12490,N_11963,N_11463);
nand U12491 (N_12491,N_11124,N_11917);
xor U12492 (N_12492,N_11958,N_11341);
nor U12493 (N_12493,N_11097,N_11519);
or U12494 (N_12494,N_11468,N_11435);
or U12495 (N_12495,N_11324,N_11927);
nor U12496 (N_12496,N_11496,N_11005);
nor U12497 (N_12497,N_11197,N_11520);
or U12498 (N_12498,N_11262,N_11773);
xor U12499 (N_12499,N_11304,N_11550);
xnor U12500 (N_12500,N_11640,N_11193);
nand U12501 (N_12501,N_11547,N_11831);
nand U12502 (N_12502,N_11884,N_11372);
and U12503 (N_12503,N_11838,N_11566);
or U12504 (N_12504,N_11138,N_11353);
and U12505 (N_12505,N_11407,N_11415);
and U12506 (N_12506,N_11908,N_11593);
or U12507 (N_12507,N_11203,N_11963);
or U12508 (N_12508,N_11255,N_11386);
nand U12509 (N_12509,N_11390,N_11822);
xnor U12510 (N_12510,N_11540,N_11139);
or U12511 (N_12511,N_11286,N_11643);
xor U12512 (N_12512,N_11595,N_11407);
nand U12513 (N_12513,N_11979,N_11786);
nand U12514 (N_12514,N_11331,N_11939);
nand U12515 (N_12515,N_11548,N_11074);
nor U12516 (N_12516,N_11638,N_11024);
and U12517 (N_12517,N_11878,N_11479);
nor U12518 (N_12518,N_11811,N_11861);
xor U12519 (N_12519,N_11071,N_11035);
nor U12520 (N_12520,N_11798,N_11906);
or U12521 (N_12521,N_11680,N_11852);
or U12522 (N_12522,N_11844,N_11959);
nand U12523 (N_12523,N_11928,N_11418);
and U12524 (N_12524,N_11666,N_11413);
and U12525 (N_12525,N_11549,N_11098);
nor U12526 (N_12526,N_11677,N_11445);
and U12527 (N_12527,N_11609,N_11007);
nand U12528 (N_12528,N_11126,N_11742);
or U12529 (N_12529,N_11347,N_11828);
and U12530 (N_12530,N_11465,N_11591);
or U12531 (N_12531,N_11164,N_11821);
and U12532 (N_12532,N_11548,N_11024);
and U12533 (N_12533,N_11616,N_11145);
or U12534 (N_12534,N_11683,N_11154);
nand U12535 (N_12535,N_11033,N_11647);
nor U12536 (N_12536,N_11068,N_11296);
nand U12537 (N_12537,N_11979,N_11800);
and U12538 (N_12538,N_11206,N_11824);
nand U12539 (N_12539,N_11075,N_11005);
and U12540 (N_12540,N_11251,N_11724);
nand U12541 (N_12541,N_11745,N_11768);
or U12542 (N_12542,N_11697,N_11718);
nor U12543 (N_12543,N_11613,N_11108);
nor U12544 (N_12544,N_11798,N_11745);
and U12545 (N_12545,N_11390,N_11284);
xor U12546 (N_12546,N_11506,N_11159);
and U12547 (N_12547,N_11053,N_11156);
xor U12548 (N_12548,N_11088,N_11227);
or U12549 (N_12549,N_11513,N_11811);
or U12550 (N_12550,N_11647,N_11732);
and U12551 (N_12551,N_11842,N_11406);
and U12552 (N_12552,N_11881,N_11664);
xnor U12553 (N_12553,N_11984,N_11756);
xor U12554 (N_12554,N_11856,N_11478);
nand U12555 (N_12555,N_11235,N_11785);
and U12556 (N_12556,N_11986,N_11576);
and U12557 (N_12557,N_11929,N_11629);
nor U12558 (N_12558,N_11157,N_11575);
nand U12559 (N_12559,N_11989,N_11570);
or U12560 (N_12560,N_11434,N_11407);
and U12561 (N_12561,N_11349,N_11461);
nor U12562 (N_12562,N_11101,N_11953);
or U12563 (N_12563,N_11615,N_11362);
nand U12564 (N_12564,N_11212,N_11540);
nor U12565 (N_12565,N_11082,N_11688);
nor U12566 (N_12566,N_11070,N_11396);
or U12567 (N_12567,N_11726,N_11044);
nand U12568 (N_12568,N_11951,N_11186);
xnor U12569 (N_12569,N_11590,N_11379);
or U12570 (N_12570,N_11571,N_11094);
nand U12571 (N_12571,N_11660,N_11997);
nor U12572 (N_12572,N_11553,N_11327);
nand U12573 (N_12573,N_11317,N_11158);
and U12574 (N_12574,N_11243,N_11898);
or U12575 (N_12575,N_11073,N_11508);
nand U12576 (N_12576,N_11332,N_11899);
or U12577 (N_12577,N_11281,N_11099);
and U12578 (N_12578,N_11414,N_11986);
and U12579 (N_12579,N_11546,N_11199);
or U12580 (N_12580,N_11767,N_11382);
nor U12581 (N_12581,N_11059,N_11565);
nor U12582 (N_12582,N_11485,N_11551);
or U12583 (N_12583,N_11701,N_11415);
and U12584 (N_12584,N_11212,N_11677);
nand U12585 (N_12585,N_11917,N_11693);
or U12586 (N_12586,N_11750,N_11761);
nor U12587 (N_12587,N_11823,N_11014);
or U12588 (N_12588,N_11026,N_11157);
or U12589 (N_12589,N_11854,N_11629);
and U12590 (N_12590,N_11686,N_11498);
nor U12591 (N_12591,N_11201,N_11569);
or U12592 (N_12592,N_11807,N_11478);
nand U12593 (N_12593,N_11830,N_11843);
nor U12594 (N_12594,N_11003,N_11330);
or U12595 (N_12595,N_11862,N_11572);
nand U12596 (N_12596,N_11177,N_11155);
or U12597 (N_12597,N_11226,N_11491);
or U12598 (N_12598,N_11232,N_11381);
nor U12599 (N_12599,N_11264,N_11414);
or U12600 (N_12600,N_11863,N_11337);
xor U12601 (N_12601,N_11652,N_11465);
nand U12602 (N_12602,N_11946,N_11302);
or U12603 (N_12603,N_11355,N_11379);
xor U12604 (N_12604,N_11281,N_11102);
nor U12605 (N_12605,N_11891,N_11592);
or U12606 (N_12606,N_11602,N_11105);
or U12607 (N_12607,N_11653,N_11820);
nand U12608 (N_12608,N_11930,N_11302);
nand U12609 (N_12609,N_11549,N_11634);
nor U12610 (N_12610,N_11431,N_11416);
nand U12611 (N_12611,N_11212,N_11525);
nand U12612 (N_12612,N_11977,N_11616);
and U12613 (N_12613,N_11098,N_11038);
xor U12614 (N_12614,N_11378,N_11461);
nand U12615 (N_12615,N_11828,N_11125);
or U12616 (N_12616,N_11093,N_11078);
or U12617 (N_12617,N_11847,N_11804);
nand U12618 (N_12618,N_11668,N_11483);
nor U12619 (N_12619,N_11810,N_11033);
nor U12620 (N_12620,N_11617,N_11195);
or U12621 (N_12621,N_11212,N_11707);
xor U12622 (N_12622,N_11798,N_11763);
and U12623 (N_12623,N_11059,N_11969);
or U12624 (N_12624,N_11810,N_11265);
nor U12625 (N_12625,N_11468,N_11589);
and U12626 (N_12626,N_11022,N_11927);
and U12627 (N_12627,N_11055,N_11629);
or U12628 (N_12628,N_11959,N_11164);
nand U12629 (N_12629,N_11675,N_11486);
and U12630 (N_12630,N_11689,N_11237);
or U12631 (N_12631,N_11621,N_11898);
xnor U12632 (N_12632,N_11198,N_11681);
or U12633 (N_12633,N_11178,N_11126);
and U12634 (N_12634,N_11103,N_11725);
nand U12635 (N_12635,N_11752,N_11459);
xnor U12636 (N_12636,N_11265,N_11824);
nor U12637 (N_12637,N_11724,N_11317);
nor U12638 (N_12638,N_11614,N_11888);
and U12639 (N_12639,N_11608,N_11640);
and U12640 (N_12640,N_11629,N_11547);
nor U12641 (N_12641,N_11797,N_11508);
nor U12642 (N_12642,N_11600,N_11082);
nor U12643 (N_12643,N_11029,N_11818);
nand U12644 (N_12644,N_11866,N_11920);
and U12645 (N_12645,N_11067,N_11745);
xnor U12646 (N_12646,N_11119,N_11150);
xor U12647 (N_12647,N_11120,N_11047);
and U12648 (N_12648,N_11859,N_11949);
xor U12649 (N_12649,N_11078,N_11151);
nand U12650 (N_12650,N_11431,N_11584);
or U12651 (N_12651,N_11336,N_11159);
nand U12652 (N_12652,N_11358,N_11813);
xor U12653 (N_12653,N_11557,N_11193);
and U12654 (N_12654,N_11297,N_11996);
and U12655 (N_12655,N_11749,N_11702);
nand U12656 (N_12656,N_11775,N_11816);
or U12657 (N_12657,N_11659,N_11529);
xnor U12658 (N_12658,N_11893,N_11959);
and U12659 (N_12659,N_11676,N_11969);
nand U12660 (N_12660,N_11947,N_11602);
or U12661 (N_12661,N_11256,N_11209);
nor U12662 (N_12662,N_11474,N_11225);
nor U12663 (N_12663,N_11499,N_11573);
and U12664 (N_12664,N_11969,N_11005);
xor U12665 (N_12665,N_11613,N_11312);
nand U12666 (N_12666,N_11890,N_11408);
nor U12667 (N_12667,N_11318,N_11547);
or U12668 (N_12668,N_11744,N_11153);
and U12669 (N_12669,N_11801,N_11750);
or U12670 (N_12670,N_11548,N_11909);
nor U12671 (N_12671,N_11503,N_11017);
or U12672 (N_12672,N_11070,N_11945);
nand U12673 (N_12673,N_11000,N_11058);
nor U12674 (N_12674,N_11262,N_11200);
or U12675 (N_12675,N_11614,N_11809);
nor U12676 (N_12676,N_11771,N_11106);
nor U12677 (N_12677,N_11826,N_11204);
nor U12678 (N_12678,N_11147,N_11667);
or U12679 (N_12679,N_11058,N_11342);
nand U12680 (N_12680,N_11099,N_11914);
xor U12681 (N_12681,N_11866,N_11078);
nor U12682 (N_12682,N_11982,N_11100);
or U12683 (N_12683,N_11221,N_11842);
and U12684 (N_12684,N_11219,N_11949);
nand U12685 (N_12685,N_11465,N_11264);
nor U12686 (N_12686,N_11576,N_11561);
nor U12687 (N_12687,N_11505,N_11043);
and U12688 (N_12688,N_11056,N_11976);
nand U12689 (N_12689,N_11018,N_11691);
nor U12690 (N_12690,N_11645,N_11208);
nor U12691 (N_12691,N_11829,N_11671);
or U12692 (N_12692,N_11087,N_11603);
or U12693 (N_12693,N_11558,N_11954);
nand U12694 (N_12694,N_11062,N_11027);
nand U12695 (N_12695,N_11306,N_11647);
and U12696 (N_12696,N_11149,N_11097);
nor U12697 (N_12697,N_11645,N_11560);
nand U12698 (N_12698,N_11057,N_11857);
xnor U12699 (N_12699,N_11565,N_11391);
or U12700 (N_12700,N_11901,N_11241);
and U12701 (N_12701,N_11135,N_11584);
nand U12702 (N_12702,N_11789,N_11408);
and U12703 (N_12703,N_11242,N_11364);
or U12704 (N_12704,N_11414,N_11446);
nor U12705 (N_12705,N_11106,N_11954);
nor U12706 (N_12706,N_11462,N_11671);
and U12707 (N_12707,N_11047,N_11342);
nor U12708 (N_12708,N_11773,N_11594);
or U12709 (N_12709,N_11090,N_11258);
nor U12710 (N_12710,N_11417,N_11306);
and U12711 (N_12711,N_11570,N_11898);
xor U12712 (N_12712,N_11581,N_11296);
or U12713 (N_12713,N_11398,N_11807);
or U12714 (N_12714,N_11341,N_11834);
nor U12715 (N_12715,N_11899,N_11493);
nor U12716 (N_12716,N_11371,N_11191);
or U12717 (N_12717,N_11725,N_11174);
nand U12718 (N_12718,N_11437,N_11093);
and U12719 (N_12719,N_11338,N_11245);
nor U12720 (N_12720,N_11083,N_11731);
and U12721 (N_12721,N_11326,N_11163);
nor U12722 (N_12722,N_11649,N_11098);
and U12723 (N_12723,N_11165,N_11474);
nor U12724 (N_12724,N_11327,N_11762);
xor U12725 (N_12725,N_11757,N_11295);
or U12726 (N_12726,N_11624,N_11958);
nand U12727 (N_12727,N_11120,N_11891);
nor U12728 (N_12728,N_11502,N_11108);
and U12729 (N_12729,N_11221,N_11890);
or U12730 (N_12730,N_11622,N_11204);
and U12731 (N_12731,N_11980,N_11903);
nand U12732 (N_12732,N_11510,N_11800);
and U12733 (N_12733,N_11596,N_11760);
nor U12734 (N_12734,N_11997,N_11287);
and U12735 (N_12735,N_11879,N_11051);
nor U12736 (N_12736,N_11670,N_11888);
xnor U12737 (N_12737,N_11181,N_11725);
or U12738 (N_12738,N_11228,N_11444);
nor U12739 (N_12739,N_11776,N_11232);
or U12740 (N_12740,N_11077,N_11186);
xor U12741 (N_12741,N_11911,N_11869);
nand U12742 (N_12742,N_11737,N_11838);
and U12743 (N_12743,N_11061,N_11123);
nand U12744 (N_12744,N_11748,N_11709);
xor U12745 (N_12745,N_11734,N_11279);
and U12746 (N_12746,N_11026,N_11431);
nor U12747 (N_12747,N_11734,N_11699);
nor U12748 (N_12748,N_11707,N_11561);
or U12749 (N_12749,N_11740,N_11608);
or U12750 (N_12750,N_11882,N_11021);
nor U12751 (N_12751,N_11888,N_11323);
or U12752 (N_12752,N_11087,N_11047);
and U12753 (N_12753,N_11130,N_11903);
nand U12754 (N_12754,N_11757,N_11376);
nand U12755 (N_12755,N_11984,N_11251);
nor U12756 (N_12756,N_11155,N_11916);
and U12757 (N_12757,N_11717,N_11948);
nand U12758 (N_12758,N_11304,N_11795);
nor U12759 (N_12759,N_11849,N_11674);
nor U12760 (N_12760,N_11553,N_11124);
or U12761 (N_12761,N_11319,N_11929);
or U12762 (N_12762,N_11751,N_11916);
and U12763 (N_12763,N_11414,N_11764);
nand U12764 (N_12764,N_11432,N_11863);
or U12765 (N_12765,N_11205,N_11117);
nor U12766 (N_12766,N_11775,N_11393);
or U12767 (N_12767,N_11018,N_11632);
nand U12768 (N_12768,N_11736,N_11975);
xnor U12769 (N_12769,N_11556,N_11373);
and U12770 (N_12770,N_11797,N_11292);
and U12771 (N_12771,N_11255,N_11767);
nand U12772 (N_12772,N_11624,N_11815);
nand U12773 (N_12773,N_11443,N_11517);
or U12774 (N_12774,N_11110,N_11191);
or U12775 (N_12775,N_11788,N_11167);
or U12776 (N_12776,N_11292,N_11072);
nand U12777 (N_12777,N_11030,N_11467);
nand U12778 (N_12778,N_11099,N_11229);
or U12779 (N_12779,N_11951,N_11147);
or U12780 (N_12780,N_11013,N_11903);
and U12781 (N_12781,N_11346,N_11271);
nor U12782 (N_12782,N_11121,N_11573);
nor U12783 (N_12783,N_11594,N_11122);
xor U12784 (N_12784,N_11818,N_11375);
nand U12785 (N_12785,N_11690,N_11342);
or U12786 (N_12786,N_11604,N_11882);
and U12787 (N_12787,N_11949,N_11622);
nor U12788 (N_12788,N_11875,N_11924);
nor U12789 (N_12789,N_11739,N_11335);
and U12790 (N_12790,N_11186,N_11543);
or U12791 (N_12791,N_11924,N_11998);
and U12792 (N_12792,N_11748,N_11298);
nor U12793 (N_12793,N_11282,N_11528);
nand U12794 (N_12794,N_11507,N_11505);
or U12795 (N_12795,N_11875,N_11259);
or U12796 (N_12796,N_11153,N_11489);
or U12797 (N_12797,N_11522,N_11616);
nand U12798 (N_12798,N_11539,N_11290);
and U12799 (N_12799,N_11148,N_11323);
nor U12800 (N_12800,N_11546,N_11574);
and U12801 (N_12801,N_11321,N_11467);
xor U12802 (N_12802,N_11037,N_11642);
nor U12803 (N_12803,N_11963,N_11526);
nor U12804 (N_12804,N_11676,N_11732);
or U12805 (N_12805,N_11672,N_11945);
and U12806 (N_12806,N_11534,N_11446);
and U12807 (N_12807,N_11699,N_11716);
nand U12808 (N_12808,N_11166,N_11925);
nand U12809 (N_12809,N_11939,N_11982);
and U12810 (N_12810,N_11913,N_11753);
nand U12811 (N_12811,N_11232,N_11166);
nand U12812 (N_12812,N_11698,N_11407);
and U12813 (N_12813,N_11816,N_11758);
or U12814 (N_12814,N_11204,N_11775);
nand U12815 (N_12815,N_11041,N_11418);
and U12816 (N_12816,N_11289,N_11761);
nor U12817 (N_12817,N_11512,N_11110);
or U12818 (N_12818,N_11451,N_11952);
or U12819 (N_12819,N_11051,N_11188);
and U12820 (N_12820,N_11467,N_11130);
nand U12821 (N_12821,N_11387,N_11767);
and U12822 (N_12822,N_11417,N_11232);
nand U12823 (N_12823,N_11226,N_11218);
and U12824 (N_12824,N_11205,N_11040);
and U12825 (N_12825,N_11404,N_11958);
and U12826 (N_12826,N_11318,N_11550);
nand U12827 (N_12827,N_11572,N_11228);
nor U12828 (N_12828,N_11939,N_11786);
and U12829 (N_12829,N_11100,N_11189);
nor U12830 (N_12830,N_11255,N_11108);
nand U12831 (N_12831,N_11730,N_11915);
nor U12832 (N_12832,N_11058,N_11590);
nand U12833 (N_12833,N_11074,N_11825);
nor U12834 (N_12834,N_11121,N_11376);
nand U12835 (N_12835,N_11079,N_11218);
xnor U12836 (N_12836,N_11641,N_11973);
nor U12837 (N_12837,N_11702,N_11281);
nand U12838 (N_12838,N_11676,N_11926);
or U12839 (N_12839,N_11787,N_11241);
and U12840 (N_12840,N_11960,N_11630);
nand U12841 (N_12841,N_11781,N_11589);
nor U12842 (N_12842,N_11337,N_11255);
nand U12843 (N_12843,N_11031,N_11460);
nand U12844 (N_12844,N_11306,N_11196);
or U12845 (N_12845,N_11640,N_11580);
and U12846 (N_12846,N_11668,N_11219);
xnor U12847 (N_12847,N_11295,N_11535);
or U12848 (N_12848,N_11675,N_11089);
and U12849 (N_12849,N_11720,N_11707);
nor U12850 (N_12850,N_11710,N_11728);
nand U12851 (N_12851,N_11956,N_11989);
nand U12852 (N_12852,N_11387,N_11611);
nor U12853 (N_12853,N_11913,N_11184);
nand U12854 (N_12854,N_11223,N_11365);
and U12855 (N_12855,N_11846,N_11242);
nand U12856 (N_12856,N_11662,N_11754);
or U12857 (N_12857,N_11838,N_11854);
nand U12858 (N_12858,N_11681,N_11643);
nor U12859 (N_12859,N_11450,N_11197);
nor U12860 (N_12860,N_11592,N_11639);
and U12861 (N_12861,N_11554,N_11754);
and U12862 (N_12862,N_11340,N_11693);
nand U12863 (N_12863,N_11858,N_11488);
nor U12864 (N_12864,N_11182,N_11744);
nand U12865 (N_12865,N_11222,N_11350);
nor U12866 (N_12866,N_11340,N_11234);
nor U12867 (N_12867,N_11655,N_11136);
nand U12868 (N_12868,N_11789,N_11441);
nor U12869 (N_12869,N_11526,N_11180);
or U12870 (N_12870,N_11259,N_11900);
nor U12871 (N_12871,N_11964,N_11108);
nand U12872 (N_12872,N_11971,N_11751);
and U12873 (N_12873,N_11885,N_11916);
nand U12874 (N_12874,N_11581,N_11964);
or U12875 (N_12875,N_11365,N_11175);
nor U12876 (N_12876,N_11162,N_11319);
nor U12877 (N_12877,N_11222,N_11130);
nand U12878 (N_12878,N_11847,N_11119);
and U12879 (N_12879,N_11938,N_11044);
and U12880 (N_12880,N_11966,N_11330);
nand U12881 (N_12881,N_11295,N_11567);
xor U12882 (N_12882,N_11968,N_11759);
nor U12883 (N_12883,N_11302,N_11271);
nor U12884 (N_12884,N_11236,N_11904);
or U12885 (N_12885,N_11478,N_11253);
or U12886 (N_12886,N_11079,N_11455);
nor U12887 (N_12887,N_11457,N_11055);
nor U12888 (N_12888,N_11840,N_11202);
xor U12889 (N_12889,N_11822,N_11759);
nand U12890 (N_12890,N_11283,N_11030);
or U12891 (N_12891,N_11870,N_11206);
and U12892 (N_12892,N_11997,N_11302);
xor U12893 (N_12893,N_11214,N_11395);
or U12894 (N_12894,N_11253,N_11788);
nand U12895 (N_12895,N_11050,N_11323);
xnor U12896 (N_12896,N_11011,N_11430);
nand U12897 (N_12897,N_11255,N_11050);
nor U12898 (N_12898,N_11773,N_11369);
or U12899 (N_12899,N_11320,N_11263);
or U12900 (N_12900,N_11012,N_11548);
nand U12901 (N_12901,N_11297,N_11392);
nor U12902 (N_12902,N_11908,N_11145);
nand U12903 (N_12903,N_11736,N_11965);
nor U12904 (N_12904,N_11415,N_11391);
and U12905 (N_12905,N_11329,N_11071);
nor U12906 (N_12906,N_11145,N_11816);
and U12907 (N_12907,N_11901,N_11320);
or U12908 (N_12908,N_11964,N_11954);
and U12909 (N_12909,N_11918,N_11208);
nand U12910 (N_12910,N_11998,N_11554);
nand U12911 (N_12911,N_11019,N_11907);
nor U12912 (N_12912,N_11157,N_11288);
or U12913 (N_12913,N_11374,N_11725);
and U12914 (N_12914,N_11030,N_11890);
or U12915 (N_12915,N_11756,N_11341);
nand U12916 (N_12916,N_11719,N_11829);
xor U12917 (N_12917,N_11508,N_11132);
nor U12918 (N_12918,N_11304,N_11207);
and U12919 (N_12919,N_11317,N_11015);
or U12920 (N_12920,N_11230,N_11900);
nor U12921 (N_12921,N_11496,N_11444);
and U12922 (N_12922,N_11000,N_11224);
or U12923 (N_12923,N_11078,N_11468);
and U12924 (N_12924,N_11847,N_11639);
or U12925 (N_12925,N_11562,N_11258);
nand U12926 (N_12926,N_11184,N_11715);
and U12927 (N_12927,N_11527,N_11598);
nor U12928 (N_12928,N_11371,N_11175);
nor U12929 (N_12929,N_11411,N_11081);
nor U12930 (N_12930,N_11944,N_11570);
nand U12931 (N_12931,N_11185,N_11493);
nor U12932 (N_12932,N_11936,N_11229);
nand U12933 (N_12933,N_11624,N_11448);
or U12934 (N_12934,N_11489,N_11120);
or U12935 (N_12935,N_11379,N_11819);
xnor U12936 (N_12936,N_11725,N_11477);
and U12937 (N_12937,N_11905,N_11972);
nor U12938 (N_12938,N_11398,N_11387);
nor U12939 (N_12939,N_11881,N_11249);
nand U12940 (N_12940,N_11748,N_11389);
nand U12941 (N_12941,N_11048,N_11270);
or U12942 (N_12942,N_11582,N_11873);
or U12943 (N_12943,N_11216,N_11530);
or U12944 (N_12944,N_11100,N_11152);
nand U12945 (N_12945,N_11688,N_11214);
nor U12946 (N_12946,N_11098,N_11925);
nand U12947 (N_12947,N_11550,N_11911);
and U12948 (N_12948,N_11078,N_11058);
nor U12949 (N_12949,N_11322,N_11624);
nand U12950 (N_12950,N_11452,N_11408);
or U12951 (N_12951,N_11895,N_11314);
nand U12952 (N_12952,N_11374,N_11313);
nand U12953 (N_12953,N_11358,N_11065);
xor U12954 (N_12954,N_11850,N_11605);
nor U12955 (N_12955,N_11362,N_11020);
nand U12956 (N_12956,N_11661,N_11747);
nand U12957 (N_12957,N_11504,N_11247);
nor U12958 (N_12958,N_11146,N_11504);
or U12959 (N_12959,N_11214,N_11095);
nand U12960 (N_12960,N_11354,N_11940);
or U12961 (N_12961,N_11771,N_11417);
nand U12962 (N_12962,N_11160,N_11848);
xnor U12963 (N_12963,N_11725,N_11974);
xor U12964 (N_12964,N_11547,N_11435);
nand U12965 (N_12965,N_11434,N_11849);
or U12966 (N_12966,N_11207,N_11123);
nor U12967 (N_12967,N_11025,N_11978);
nand U12968 (N_12968,N_11028,N_11244);
nand U12969 (N_12969,N_11749,N_11003);
xor U12970 (N_12970,N_11831,N_11992);
nand U12971 (N_12971,N_11648,N_11026);
nor U12972 (N_12972,N_11047,N_11930);
xor U12973 (N_12973,N_11209,N_11444);
nand U12974 (N_12974,N_11442,N_11899);
or U12975 (N_12975,N_11169,N_11187);
or U12976 (N_12976,N_11209,N_11930);
nand U12977 (N_12977,N_11495,N_11465);
and U12978 (N_12978,N_11447,N_11774);
and U12979 (N_12979,N_11623,N_11208);
and U12980 (N_12980,N_11409,N_11951);
or U12981 (N_12981,N_11790,N_11567);
nor U12982 (N_12982,N_11687,N_11074);
nand U12983 (N_12983,N_11281,N_11158);
nand U12984 (N_12984,N_11261,N_11766);
xor U12985 (N_12985,N_11322,N_11538);
or U12986 (N_12986,N_11979,N_11000);
or U12987 (N_12987,N_11015,N_11997);
nor U12988 (N_12988,N_11728,N_11811);
or U12989 (N_12989,N_11769,N_11365);
nand U12990 (N_12990,N_11553,N_11837);
nand U12991 (N_12991,N_11199,N_11878);
or U12992 (N_12992,N_11157,N_11967);
nand U12993 (N_12993,N_11287,N_11925);
nand U12994 (N_12994,N_11750,N_11040);
nor U12995 (N_12995,N_11530,N_11755);
and U12996 (N_12996,N_11854,N_11131);
or U12997 (N_12997,N_11616,N_11906);
or U12998 (N_12998,N_11299,N_11435);
nand U12999 (N_12999,N_11485,N_11702);
nor U13000 (N_13000,N_12624,N_12848);
nand U13001 (N_13001,N_12393,N_12042);
and U13002 (N_13002,N_12509,N_12784);
or U13003 (N_13003,N_12902,N_12401);
nor U13004 (N_13004,N_12482,N_12626);
or U13005 (N_13005,N_12919,N_12027);
xnor U13006 (N_13006,N_12828,N_12849);
and U13007 (N_13007,N_12392,N_12181);
nor U13008 (N_13008,N_12557,N_12255);
nand U13009 (N_13009,N_12096,N_12763);
xor U13010 (N_13010,N_12861,N_12313);
nor U13011 (N_13011,N_12333,N_12842);
nand U13012 (N_13012,N_12185,N_12057);
or U13013 (N_13013,N_12868,N_12007);
or U13014 (N_13014,N_12951,N_12693);
or U13015 (N_13015,N_12550,N_12862);
nand U13016 (N_13016,N_12111,N_12016);
and U13017 (N_13017,N_12934,N_12238);
xor U13018 (N_13018,N_12399,N_12069);
and U13019 (N_13019,N_12450,N_12499);
nand U13020 (N_13020,N_12944,N_12014);
nor U13021 (N_13021,N_12968,N_12692);
and U13022 (N_13022,N_12438,N_12706);
nor U13023 (N_13023,N_12101,N_12044);
nor U13024 (N_13024,N_12725,N_12325);
xor U13025 (N_13025,N_12252,N_12371);
nand U13026 (N_13026,N_12491,N_12261);
or U13027 (N_13027,N_12166,N_12493);
and U13028 (N_13028,N_12687,N_12200);
nor U13029 (N_13029,N_12078,N_12616);
and U13030 (N_13030,N_12536,N_12378);
or U13031 (N_13031,N_12584,N_12956);
nand U13032 (N_13032,N_12782,N_12742);
xnor U13033 (N_13033,N_12983,N_12955);
nand U13034 (N_13034,N_12685,N_12085);
or U13035 (N_13035,N_12795,N_12530);
or U13036 (N_13036,N_12937,N_12437);
nand U13037 (N_13037,N_12946,N_12816);
nand U13038 (N_13038,N_12621,N_12760);
and U13039 (N_13039,N_12328,N_12113);
nor U13040 (N_13040,N_12143,N_12641);
nand U13041 (N_13041,N_12202,N_12984);
or U13042 (N_13042,N_12406,N_12194);
nor U13043 (N_13043,N_12971,N_12239);
and U13044 (N_13044,N_12894,N_12290);
or U13045 (N_13045,N_12589,N_12368);
and U13046 (N_13046,N_12236,N_12998);
or U13047 (N_13047,N_12957,N_12366);
and U13048 (N_13048,N_12344,N_12746);
nand U13049 (N_13049,N_12941,N_12588);
or U13050 (N_13050,N_12758,N_12337);
and U13051 (N_13051,N_12248,N_12443);
nand U13052 (N_13052,N_12822,N_12100);
and U13053 (N_13053,N_12191,N_12581);
nor U13054 (N_13054,N_12487,N_12628);
and U13055 (N_13055,N_12153,N_12747);
nor U13056 (N_13056,N_12182,N_12470);
xor U13057 (N_13057,N_12764,N_12989);
or U13058 (N_13058,N_12282,N_12750);
nand U13059 (N_13059,N_12323,N_12400);
nor U13060 (N_13060,N_12089,N_12835);
nor U13061 (N_13061,N_12730,N_12217);
nand U13062 (N_13062,N_12208,N_12529);
nand U13063 (N_13063,N_12108,N_12121);
nand U13064 (N_13064,N_12295,N_12434);
nand U13065 (N_13065,N_12966,N_12321);
nand U13066 (N_13066,N_12579,N_12504);
or U13067 (N_13067,N_12990,N_12445);
and U13068 (N_13068,N_12637,N_12526);
nor U13069 (N_13069,N_12080,N_12312);
nor U13070 (N_13070,N_12864,N_12379);
nand U13071 (N_13071,N_12205,N_12396);
or U13072 (N_13072,N_12954,N_12347);
and U13073 (N_13073,N_12767,N_12674);
nand U13074 (N_13074,N_12876,N_12712);
and U13075 (N_13075,N_12840,N_12924);
nor U13076 (N_13076,N_12053,N_12022);
and U13077 (N_13077,N_12225,N_12117);
or U13078 (N_13078,N_12247,N_12353);
or U13079 (N_13079,N_12918,N_12883);
nor U13080 (N_13080,N_12150,N_12943);
and U13081 (N_13081,N_12890,N_12729);
nor U13082 (N_13082,N_12308,N_12420);
or U13083 (N_13083,N_12567,N_12939);
nor U13084 (N_13084,N_12723,N_12133);
nand U13085 (N_13085,N_12190,N_12935);
nand U13086 (N_13086,N_12929,N_12696);
and U13087 (N_13087,N_12600,N_12008);
or U13088 (N_13088,N_12978,N_12967);
xor U13089 (N_13089,N_12229,N_12005);
xnor U13090 (N_13090,N_12518,N_12301);
or U13091 (N_13091,N_12115,N_12235);
nor U13092 (N_13092,N_12300,N_12775);
nand U13093 (N_13093,N_12187,N_12291);
nor U13094 (N_13094,N_12461,N_12768);
nand U13095 (N_13095,N_12000,N_12718);
nand U13096 (N_13096,N_12218,N_12360);
and U13097 (N_13097,N_12836,N_12852);
nor U13098 (N_13098,N_12908,N_12374);
and U13099 (N_13099,N_12413,N_12986);
nand U13100 (N_13100,N_12538,N_12112);
nand U13101 (N_13101,N_12036,N_12352);
nand U13102 (N_13102,N_12549,N_12260);
nor U13103 (N_13103,N_12179,N_12761);
and U13104 (N_13104,N_12613,N_12972);
or U13105 (N_13105,N_12907,N_12365);
and U13106 (N_13106,N_12433,N_12256);
and U13107 (N_13107,N_12201,N_12534);
and U13108 (N_13108,N_12815,N_12316);
nor U13109 (N_13109,N_12915,N_12077);
or U13110 (N_13110,N_12863,N_12394);
nor U13111 (N_13111,N_12601,N_12029);
nand U13112 (N_13112,N_12359,N_12219);
or U13113 (N_13113,N_12326,N_12369);
and U13114 (N_13114,N_12683,N_12426);
or U13115 (N_13115,N_12796,N_12783);
or U13116 (N_13116,N_12031,N_12129);
xnor U13117 (N_13117,N_12410,N_12668);
xnor U13118 (N_13118,N_12342,N_12855);
nor U13119 (N_13119,N_12574,N_12521);
nand U13120 (N_13120,N_12040,N_12009);
nor U13121 (N_13121,N_12331,N_12982);
nand U13122 (N_13122,N_12858,N_12748);
or U13123 (N_13123,N_12933,N_12074);
nor U13124 (N_13124,N_12168,N_12072);
or U13125 (N_13125,N_12421,N_12043);
nor U13126 (N_13126,N_12932,N_12887);
nor U13127 (N_13127,N_12576,N_12528);
xor U13128 (N_13128,N_12411,N_12165);
or U13129 (N_13129,N_12173,N_12498);
and U13130 (N_13130,N_12423,N_12432);
and U13131 (N_13131,N_12176,N_12987);
nor U13132 (N_13132,N_12599,N_12854);
or U13133 (N_13133,N_12464,N_12569);
nand U13134 (N_13134,N_12304,N_12682);
or U13135 (N_13135,N_12094,N_12644);
or U13136 (N_13136,N_12677,N_12083);
and U13137 (N_13137,N_12032,N_12759);
nor U13138 (N_13138,N_12339,N_12170);
or U13139 (N_13139,N_12812,N_12542);
and U13140 (N_13140,N_12596,N_12125);
or U13141 (N_13141,N_12517,N_12422);
or U13142 (N_13142,N_12947,N_12778);
or U13143 (N_13143,N_12048,N_12669);
and U13144 (N_13144,N_12329,N_12506);
xnor U13145 (N_13145,N_12361,N_12676);
nor U13146 (N_13146,N_12899,N_12702);
nor U13147 (N_13147,N_12192,N_12382);
and U13148 (N_13148,N_12772,N_12926);
and U13149 (N_13149,N_12212,N_12925);
and U13150 (N_13150,N_12597,N_12116);
nand U13151 (N_13151,N_12324,N_12348);
and U13152 (N_13152,N_12631,N_12271);
nor U13153 (N_13153,N_12996,N_12246);
nand U13154 (N_13154,N_12037,N_12152);
nand U13155 (N_13155,N_12351,N_12653);
xor U13156 (N_13156,N_12846,N_12727);
nor U13157 (N_13157,N_12976,N_12198);
or U13158 (N_13158,N_12390,N_12845);
and U13159 (N_13159,N_12994,N_12086);
xor U13160 (N_13160,N_12771,N_12817);
and U13161 (N_13161,N_12573,N_12566);
or U13162 (N_13162,N_12804,N_12741);
nor U13163 (N_13163,N_12395,N_12879);
and U13164 (N_13164,N_12448,N_12684);
and U13165 (N_13165,N_12178,N_12265);
and U13166 (N_13166,N_12250,N_12928);
or U13167 (N_13167,N_12722,N_12444);
xnor U13168 (N_13168,N_12708,N_12473);
nand U13169 (N_13169,N_12656,N_12690);
nand U13170 (N_13170,N_12226,N_12633);
nand U13171 (N_13171,N_12895,N_12012);
or U13172 (N_13172,N_12640,N_12026);
nand U13173 (N_13173,N_12507,N_12713);
and U13174 (N_13174,N_12732,N_12647);
nor U13175 (N_13175,N_12385,N_12652);
or U13176 (N_13176,N_12267,N_12680);
nor U13177 (N_13177,N_12992,N_12885);
and U13178 (N_13178,N_12535,N_12617);
nand U13179 (N_13179,N_12346,N_12625);
and U13180 (N_13180,N_12338,N_12439);
nand U13181 (N_13181,N_12552,N_12303);
or U13182 (N_13182,N_12131,N_12866);
nor U13183 (N_13183,N_12277,N_12427);
nor U13184 (N_13184,N_12950,N_12160);
or U13185 (N_13185,N_12296,N_12468);
or U13186 (N_13186,N_12857,N_12503);
and U13187 (N_13187,N_12788,N_12577);
nor U13188 (N_13188,N_12013,N_12765);
nor U13189 (N_13189,N_12466,N_12561);
xor U13190 (N_13190,N_12824,N_12478);
xor U13191 (N_13191,N_12435,N_12974);
and U13192 (N_13192,N_12233,N_12122);
nor U13193 (N_13193,N_12716,N_12310);
xor U13194 (N_13194,N_12480,N_12797);
nor U13195 (N_13195,N_12903,N_12106);
nor U13196 (N_13196,N_12222,N_12632);
nor U13197 (N_13197,N_12293,N_12847);
nor U13198 (N_13198,N_12490,N_12388);
nand U13199 (N_13199,N_12556,N_12288);
nor U13200 (N_13200,N_12622,N_12207);
nor U13201 (N_13201,N_12524,N_12402);
xor U13202 (N_13202,N_12414,N_12999);
nand U13203 (N_13203,N_12384,N_12523);
and U13204 (N_13204,N_12512,N_12193);
xor U13205 (N_13205,N_12896,N_12881);
nor U13206 (N_13206,N_12901,N_12243);
and U13207 (N_13207,N_12560,N_12472);
xnor U13208 (N_13208,N_12062,N_12398);
or U13209 (N_13209,N_12496,N_12403);
nand U13210 (N_13210,N_12808,N_12594);
nor U13211 (N_13211,N_12638,N_12098);
nor U13212 (N_13212,N_12958,N_12463);
and U13213 (N_13213,N_12520,N_12734);
xnor U13214 (N_13214,N_12270,N_12372);
or U13215 (N_13215,N_12407,N_12068);
or U13216 (N_13216,N_12010,N_12714);
and U13217 (N_13217,N_12969,N_12021);
and U13218 (N_13218,N_12436,N_12041);
xnor U13219 (N_13219,N_12819,N_12017);
or U13220 (N_13220,N_12921,N_12287);
nor U13221 (N_13221,N_12284,N_12412);
or U13222 (N_13222,N_12389,N_12878);
xor U13223 (N_13223,N_12602,N_12033);
or U13224 (N_13224,N_12244,N_12162);
and U13225 (N_13225,N_12744,N_12649);
nor U13226 (N_13226,N_12608,N_12704);
nand U13227 (N_13227,N_12405,N_12709);
nor U13228 (N_13228,N_12501,N_12335);
or U13229 (N_13229,N_12736,N_12237);
nor U13230 (N_13230,N_12663,N_12047);
or U13231 (N_13231,N_12157,N_12306);
xor U13232 (N_13232,N_12320,N_12197);
nand U13233 (N_13233,N_12672,N_12497);
nor U13234 (N_13234,N_12871,N_12457);
nor U13235 (N_13235,N_12332,N_12505);
nand U13236 (N_13236,N_12780,N_12721);
or U13237 (N_13237,N_12770,N_12701);
or U13238 (N_13238,N_12158,N_12280);
and U13239 (N_13239,N_12206,N_12964);
nand U13240 (N_13240,N_12268,N_12532);
nand U13241 (N_13241,N_12651,N_12350);
or U13242 (N_13242,N_12686,N_12059);
nor U13243 (N_13243,N_12163,N_12234);
xnor U13244 (N_13244,N_12615,N_12906);
and U13245 (N_13245,N_12429,N_12144);
xnor U13246 (N_13246,N_12965,N_12773);
and U13247 (N_13247,N_12809,N_12880);
or U13248 (N_13248,N_12298,N_12859);
and U13249 (N_13249,N_12645,N_12790);
nand U13250 (N_13250,N_12024,N_12130);
or U13251 (N_13251,N_12114,N_12850);
nor U13252 (N_13252,N_12109,N_12161);
and U13253 (N_13253,N_12897,N_12263);
and U13254 (N_13254,N_12458,N_12756);
xnor U13255 (N_13255,N_12662,N_12164);
and U13256 (N_13256,N_12962,N_12643);
xor U13257 (N_13257,N_12830,N_12084);
or U13258 (N_13258,N_12107,N_12533);
nor U13259 (N_13259,N_12035,N_12650);
and U13260 (N_13260,N_12807,N_12126);
nand U13261 (N_13261,N_12948,N_12699);
nand U13262 (N_13262,N_12038,N_12299);
xnor U13263 (N_13263,N_12180,N_12249);
nor U13264 (N_13264,N_12343,N_12664);
nand U13265 (N_13265,N_12909,N_12060);
nor U13266 (N_13266,N_12737,N_12891);
or U13267 (N_13267,N_12777,N_12541);
nand U13268 (N_13268,N_12720,N_12110);
nor U13269 (N_13269,N_12140,N_12474);
or U13270 (N_13270,N_12648,N_12373);
or U13271 (N_13271,N_12203,N_12922);
and U13272 (N_13272,N_12095,N_12051);
and U13273 (N_13273,N_12492,N_12869);
and U13274 (N_13274,N_12514,N_12075);
nand U13275 (N_13275,N_12548,N_12431);
or U13276 (N_13276,N_12305,N_12050);
and U13277 (N_13277,N_12171,N_12483);
nand U13278 (N_13278,N_12156,N_12386);
and U13279 (N_13279,N_12266,N_12104);
nand U13280 (N_13280,N_12551,N_12091);
nor U13281 (N_13281,N_12449,N_12079);
nand U13282 (N_13282,N_12877,N_12066);
nor U13283 (N_13283,N_12120,N_12565);
xor U13284 (N_13284,N_12169,N_12015);
and U13285 (N_13285,N_12446,N_12149);
nor U13286 (N_13286,N_12274,N_12991);
nor U13287 (N_13287,N_12397,N_12341);
nor U13288 (N_13288,N_12317,N_12619);
nor U13289 (N_13289,N_12054,N_12465);
and U13290 (N_13290,N_12264,N_12058);
nor U13291 (N_13291,N_12330,N_12802);
and U13292 (N_13292,N_12949,N_12214);
or U13293 (N_13293,N_12322,N_12315);
nor U13294 (N_13294,N_12930,N_12019);
nand U13295 (N_13295,N_12189,N_12916);
or U13296 (N_13296,N_12884,N_12911);
nand U13297 (N_13297,N_12592,N_12774);
and U13298 (N_13298,N_12289,N_12279);
and U13299 (N_13299,N_12914,N_12242);
or U13300 (N_13300,N_12415,N_12598);
or U13301 (N_13301,N_12367,N_12961);
and U13302 (N_13302,N_12245,N_12227);
or U13303 (N_13303,N_12064,N_12665);
and U13304 (N_13304,N_12654,N_12417);
xor U13305 (N_13305,N_12297,N_12061);
and U13306 (N_13306,N_12997,N_12319);
and U13307 (N_13307,N_12011,N_12105);
and U13308 (N_13308,N_12381,N_12791);
and U13309 (N_13309,N_12540,N_12476);
nand U13310 (N_13310,N_12585,N_12762);
xor U13311 (N_13311,N_12988,N_12612);
nor U13312 (N_13312,N_12658,N_12408);
or U13313 (N_13313,N_12695,N_12258);
and U13314 (N_13314,N_12087,N_12134);
nand U13315 (N_13315,N_12151,N_12065);
and U13316 (N_13316,N_12798,N_12092);
nand U13317 (N_13317,N_12975,N_12872);
nand U13318 (N_13318,N_12519,N_12831);
nor U13319 (N_13319,N_12580,N_12546);
or U13320 (N_13320,N_12749,N_12071);
or U13321 (N_13321,N_12841,N_12159);
or U13322 (N_13322,N_12609,N_12082);
xnor U13323 (N_13323,N_12927,N_12023);
or U13324 (N_13324,N_12981,N_12726);
and U13325 (N_13325,N_12132,N_12118);
nand U13326 (N_13326,N_12302,N_12155);
or U13327 (N_13327,N_12428,N_12562);
nor U13328 (N_13328,N_12874,N_12525);
nor U13329 (N_13329,N_12275,N_12088);
or U13330 (N_13330,N_12820,N_12823);
xor U13331 (N_13331,N_12670,N_12860);
and U13332 (N_13332,N_12294,N_12188);
nor U13333 (N_13333,N_12634,N_12826);
or U13334 (N_13334,N_12004,N_12667);
nand U13335 (N_13335,N_12442,N_12177);
and U13336 (N_13336,N_12856,N_12694);
nand U13337 (N_13337,N_12779,N_12886);
or U13338 (N_13338,N_12454,N_12142);
nor U13339 (N_13339,N_12545,N_12418);
and U13340 (N_13340,N_12605,N_12278);
or U13341 (N_13341,N_12851,N_12728);
and U13342 (N_13342,N_12138,N_12210);
nor U13343 (N_13343,N_12500,N_12232);
nor U13344 (N_13344,N_12655,N_12660);
or U13345 (N_13345,N_12931,N_12595);
nor U13346 (N_13346,N_12568,N_12495);
nand U13347 (N_13347,N_12103,N_12776);
or U13348 (N_13348,N_12618,N_12554);
or U13349 (N_13349,N_12707,N_12073);
and U13350 (N_13350,N_12920,N_12827);
and U13351 (N_13351,N_12544,N_12515);
nand U13352 (N_13352,N_12357,N_12710);
or U13353 (N_13353,N_12183,N_12636);
nand U13354 (N_13354,N_12553,N_12285);
nor U13355 (N_13355,N_12508,N_12953);
or U13356 (N_13356,N_12629,N_12067);
or U13357 (N_13357,N_12898,N_12471);
and U13358 (N_13358,N_12485,N_12838);
and U13359 (N_13359,N_12785,N_12810);
nor U13360 (N_13360,N_12698,N_12805);
nor U13361 (N_13361,N_12383,N_12980);
and U13362 (N_13362,N_12547,N_12558);
nor U13363 (N_13363,N_12829,N_12211);
nor U13364 (N_13364,N_12416,N_12006);
and U13365 (N_13365,N_12757,N_12711);
xor U13366 (N_13366,N_12754,N_12952);
and U13367 (N_13367,N_12889,N_12570);
and U13368 (N_13368,N_12063,N_12221);
and U13369 (N_13369,N_12590,N_12583);
nand U13370 (N_13370,N_12787,N_12821);
nor U13371 (N_13371,N_12184,N_12052);
nor U13372 (N_13372,N_12527,N_12362);
and U13373 (N_13373,N_12689,N_12241);
nand U13374 (N_13374,N_12910,N_12799);
nand U13375 (N_13375,N_12970,N_12705);
nand U13376 (N_13376,N_12124,N_12314);
nor U13377 (N_13377,N_12257,N_12766);
nand U13378 (N_13378,N_12963,N_12912);
xnor U13379 (N_13379,N_12995,N_12469);
and U13380 (N_13380,N_12959,N_12145);
nor U13381 (N_13381,N_12404,N_12681);
and U13382 (N_13382,N_12380,N_12635);
xnor U13383 (N_13383,N_12196,N_12803);
nor U13384 (N_13384,N_12452,N_12093);
nor U13385 (N_13385,N_12049,N_12659);
or U13386 (N_13386,N_12657,N_12494);
nor U13387 (N_13387,N_12174,N_12940);
nor U13388 (N_13388,N_12070,N_12703);
and U13389 (N_13389,N_12844,N_12571);
nor U13390 (N_13390,N_12440,N_12905);
nor U13391 (N_13391,N_12055,N_12003);
or U13392 (N_13392,N_12195,N_12630);
nand U13393 (N_13393,N_12376,N_12801);
nand U13394 (N_13394,N_12673,N_12484);
nand U13395 (N_13395,N_12276,N_12985);
and U13396 (N_13396,N_12539,N_12455);
and U13397 (N_13397,N_12025,N_12419);
nor U13398 (N_13398,N_12309,N_12018);
and U13399 (N_13399,N_12642,N_12215);
and U13400 (N_13400,N_12475,N_12893);
nand U13401 (N_13401,N_12186,N_12942);
and U13402 (N_13402,N_12076,N_12811);
nand U13403 (N_13403,N_12479,N_12979);
and U13404 (N_13404,N_12724,N_12020);
nor U13405 (N_13405,N_12141,N_12262);
nor U13406 (N_13406,N_12254,N_12230);
or U13407 (N_13407,N_12833,N_12447);
nor U13408 (N_13408,N_12700,N_12209);
and U13409 (N_13409,N_12888,N_12090);
and U13410 (N_13410,N_12307,N_12391);
or U13411 (N_13411,N_12843,N_12738);
and U13412 (N_13412,N_12814,N_12611);
nor U13413 (N_13413,N_12719,N_12513);
nand U13414 (N_13414,N_12510,N_12269);
nor U13415 (N_13415,N_12224,N_12792);
nor U13416 (N_13416,N_12753,N_12001);
nand U13417 (N_13417,N_12993,N_12867);
nand U13418 (N_13418,N_12837,N_12128);
and U13419 (N_13419,N_12318,N_12904);
nand U13420 (N_13420,N_12136,N_12697);
and U13421 (N_13421,N_12977,N_12620);
nor U13422 (N_13422,N_12752,N_12477);
nand U13423 (N_13423,N_12900,N_12559);
nand U13424 (N_13424,N_12030,N_12387);
xnor U13425 (N_13425,N_12148,N_12356);
nor U13426 (N_13426,N_12870,N_12167);
xnor U13427 (N_13427,N_12639,N_12818);
nor U13428 (N_13428,N_12502,N_12781);
nand U13429 (N_13429,N_12354,N_12960);
nand U13430 (N_13430,N_12675,N_12733);
and U13431 (N_13431,N_12789,N_12220);
nand U13432 (N_13432,N_12671,N_12610);
nand U13433 (N_13433,N_12614,N_12204);
xor U13434 (N_13434,N_12481,N_12028);
nor U13435 (N_13435,N_12459,N_12800);
or U13436 (N_13436,N_12358,N_12606);
xor U13437 (N_13437,N_12039,N_12623);
and U13438 (N_13438,N_12199,N_12240);
nand U13439 (N_13439,N_12661,N_12216);
xnor U13440 (N_13440,N_12739,N_12147);
nand U13441 (N_13441,N_12715,N_12228);
or U13442 (N_13442,N_12587,N_12172);
nor U13443 (N_13443,N_12213,N_12586);
nand U13444 (N_13444,N_12137,N_12002);
nand U13445 (N_13445,N_12045,N_12865);
or U13446 (N_13446,N_12127,N_12441);
or U13447 (N_13447,N_12832,N_12769);
nor U13448 (N_13448,N_12462,N_12794);
or U13449 (N_13449,N_12231,N_12355);
nor U13450 (N_13450,N_12292,N_12489);
xor U13451 (N_13451,N_12460,N_12751);
nor U13452 (N_13452,N_12451,N_12575);
or U13453 (N_13453,N_12253,N_12679);
nand U13454 (N_13454,N_12456,N_12511);
or U13455 (N_13455,N_12488,N_12875);
nand U13456 (N_13456,N_12516,N_12572);
and U13457 (N_13457,N_12813,N_12409);
nand U13458 (N_13458,N_12731,N_12146);
xor U13459 (N_13459,N_12537,N_12873);
nor U13460 (N_13460,N_12123,N_12563);
nor U13461 (N_13461,N_12097,N_12467);
or U13462 (N_13462,N_12283,N_12375);
and U13463 (N_13463,N_12046,N_12119);
and U13464 (N_13464,N_12056,N_12717);
nor U13465 (N_13465,N_12281,N_12735);
and U13466 (N_13466,N_12593,N_12364);
nor U13467 (N_13467,N_12892,N_12430);
and U13468 (N_13468,N_12377,N_12603);
nand U13469 (N_13469,N_12745,N_12607);
xnor U13470 (N_13470,N_12543,N_12917);
or U13471 (N_13471,N_12425,N_12834);
nand U13472 (N_13472,N_12691,N_12154);
and U13473 (N_13473,N_12522,N_12688);
nor U13474 (N_13474,N_12825,N_12882);
nand U13475 (N_13475,N_12251,N_12336);
or U13476 (N_13476,N_12340,N_12135);
or U13477 (N_13477,N_12853,N_12666);
nor U13478 (N_13478,N_12743,N_12311);
and U13479 (N_13479,N_12740,N_12604);
or U13480 (N_13480,N_12945,N_12793);
or U13481 (N_13481,N_12034,N_12139);
or U13482 (N_13482,N_12486,N_12627);
nor U13483 (N_13483,N_12938,N_12272);
and U13484 (N_13484,N_12175,N_12363);
nor U13485 (N_13485,N_12578,N_12327);
nand U13486 (N_13486,N_12973,N_12936);
nand U13487 (N_13487,N_12102,N_12678);
or U13488 (N_13488,N_12424,N_12646);
or U13489 (N_13489,N_12755,N_12081);
xor U13490 (N_13490,N_12582,N_12349);
and U13491 (N_13491,N_12334,N_12913);
nand U13492 (N_13492,N_12286,N_12531);
or U13493 (N_13493,N_12099,N_12453);
or U13494 (N_13494,N_12370,N_12564);
nor U13495 (N_13495,N_12923,N_12591);
nor U13496 (N_13496,N_12806,N_12223);
and U13497 (N_13497,N_12555,N_12259);
or U13498 (N_13498,N_12786,N_12273);
or U13499 (N_13499,N_12839,N_12345);
or U13500 (N_13500,N_12938,N_12368);
nor U13501 (N_13501,N_12680,N_12481);
or U13502 (N_13502,N_12795,N_12439);
and U13503 (N_13503,N_12760,N_12518);
nor U13504 (N_13504,N_12074,N_12404);
or U13505 (N_13505,N_12146,N_12786);
xnor U13506 (N_13506,N_12616,N_12588);
or U13507 (N_13507,N_12070,N_12167);
and U13508 (N_13508,N_12733,N_12905);
nand U13509 (N_13509,N_12498,N_12495);
nand U13510 (N_13510,N_12016,N_12579);
xor U13511 (N_13511,N_12429,N_12932);
or U13512 (N_13512,N_12446,N_12547);
or U13513 (N_13513,N_12118,N_12223);
nand U13514 (N_13514,N_12159,N_12016);
nand U13515 (N_13515,N_12027,N_12664);
or U13516 (N_13516,N_12748,N_12726);
nand U13517 (N_13517,N_12245,N_12104);
nand U13518 (N_13518,N_12557,N_12621);
and U13519 (N_13519,N_12659,N_12451);
nand U13520 (N_13520,N_12128,N_12771);
and U13521 (N_13521,N_12492,N_12288);
nor U13522 (N_13522,N_12943,N_12817);
nand U13523 (N_13523,N_12036,N_12214);
nand U13524 (N_13524,N_12361,N_12966);
or U13525 (N_13525,N_12117,N_12717);
and U13526 (N_13526,N_12568,N_12335);
nor U13527 (N_13527,N_12945,N_12265);
and U13528 (N_13528,N_12115,N_12492);
nor U13529 (N_13529,N_12333,N_12769);
or U13530 (N_13530,N_12057,N_12264);
nor U13531 (N_13531,N_12245,N_12619);
nor U13532 (N_13532,N_12937,N_12617);
xor U13533 (N_13533,N_12192,N_12666);
nor U13534 (N_13534,N_12229,N_12624);
xor U13535 (N_13535,N_12159,N_12710);
nand U13536 (N_13536,N_12538,N_12913);
nor U13537 (N_13537,N_12269,N_12747);
xnor U13538 (N_13538,N_12509,N_12326);
or U13539 (N_13539,N_12269,N_12048);
and U13540 (N_13540,N_12934,N_12338);
nand U13541 (N_13541,N_12508,N_12805);
nand U13542 (N_13542,N_12226,N_12542);
nor U13543 (N_13543,N_12592,N_12689);
or U13544 (N_13544,N_12773,N_12788);
or U13545 (N_13545,N_12369,N_12431);
and U13546 (N_13546,N_12483,N_12583);
or U13547 (N_13547,N_12894,N_12180);
nand U13548 (N_13548,N_12499,N_12092);
nor U13549 (N_13549,N_12216,N_12780);
or U13550 (N_13550,N_12022,N_12082);
nor U13551 (N_13551,N_12201,N_12287);
xor U13552 (N_13552,N_12928,N_12973);
nor U13553 (N_13553,N_12686,N_12065);
or U13554 (N_13554,N_12975,N_12108);
nor U13555 (N_13555,N_12422,N_12681);
and U13556 (N_13556,N_12415,N_12728);
nand U13557 (N_13557,N_12099,N_12780);
and U13558 (N_13558,N_12571,N_12070);
and U13559 (N_13559,N_12985,N_12559);
and U13560 (N_13560,N_12622,N_12103);
nand U13561 (N_13561,N_12626,N_12672);
or U13562 (N_13562,N_12238,N_12458);
nand U13563 (N_13563,N_12910,N_12156);
xnor U13564 (N_13564,N_12514,N_12613);
or U13565 (N_13565,N_12936,N_12952);
xnor U13566 (N_13566,N_12987,N_12661);
nor U13567 (N_13567,N_12751,N_12088);
or U13568 (N_13568,N_12935,N_12140);
nand U13569 (N_13569,N_12214,N_12724);
and U13570 (N_13570,N_12100,N_12622);
or U13571 (N_13571,N_12233,N_12249);
nand U13572 (N_13572,N_12898,N_12939);
or U13573 (N_13573,N_12321,N_12970);
and U13574 (N_13574,N_12355,N_12771);
and U13575 (N_13575,N_12282,N_12570);
and U13576 (N_13576,N_12901,N_12317);
or U13577 (N_13577,N_12098,N_12785);
xnor U13578 (N_13578,N_12031,N_12800);
and U13579 (N_13579,N_12107,N_12404);
and U13580 (N_13580,N_12358,N_12501);
nand U13581 (N_13581,N_12601,N_12637);
or U13582 (N_13582,N_12607,N_12766);
and U13583 (N_13583,N_12490,N_12432);
xor U13584 (N_13584,N_12045,N_12072);
nand U13585 (N_13585,N_12053,N_12153);
nand U13586 (N_13586,N_12353,N_12260);
and U13587 (N_13587,N_12109,N_12461);
and U13588 (N_13588,N_12928,N_12637);
nor U13589 (N_13589,N_12415,N_12758);
and U13590 (N_13590,N_12175,N_12793);
nand U13591 (N_13591,N_12700,N_12801);
nor U13592 (N_13592,N_12225,N_12930);
nor U13593 (N_13593,N_12842,N_12453);
nand U13594 (N_13594,N_12315,N_12390);
xnor U13595 (N_13595,N_12047,N_12455);
xor U13596 (N_13596,N_12087,N_12819);
nand U13597 (N_13597,N_12924,N_12109);
and U13598 (N_13598,N_12557,N_12490);
and U13599 (N_13599,N_12750,N_12153);
or U13600 (N_13600,N_12920,N_12983);
or U13601 (N_13601,N_12143,N_12899);
xnor U13602 (N_13602,N_12008,N_12210);
xnor U13603 (N_13603,N_12462,N_12997);
or U13604 (N_13604,N_12339,N_12225);
or U13605 (N_13605,N_12191,N_12197);
nand U13606 (N_13606,N_12880,N_12565);
or U13607 (N_13607,N_12401,N_12066);
or U13608 (N_13608,N_12883,N_12413);
or U13609 (N_13609,N_12709,N_12976);
nand U13610 (N_13610,N_12269,N_12293);
nand U13611 (N_13611,N_12332,N_12945);
nor U13612 (N_13612,N_12804,N_12935);
nor U13613 (N_13613,N_12929,N_12099);
nand U13614 (N_13614,N_12636,N_12584);
nor U13615 (N_13615,N_12034,N_12445);
or U13616 (N_13616,N_12564,N_12141);
nand U13617 (N_13617,N_12579,N_12693);
and U13618 (N_13618,N_12699,N_12068);
or U13619 (N_13619,N_12724,N_12432);
xor U13620 (N_13620,N_12281,N_12732);
nor U13621 (N_13621,N_12383,N_12138);
nand U13622 (N_13622,N_12776,N_12041);
nor U13623 (N_13623,N_12022,N_12694);
nor U13624 (N_13624,N_12823,N_12516);
nand U13625 (N_13625,N_12955,N_12382);
nor U13626 (N_13626,N_12777,N_12351);
nand U13627 (N_13627,N_12863,N_12975);
and U13628 (N_13628,N_12436,N_12249);
or U13629 (N_13629,N_12090,N_12405);
or U13630 (N_13630,N_12153,N_12408);
nor U13631 (N_13631,N_12237,N_12021);
nor U13632 (N_13632,N_12269,N_12338);
nor U13633 (N_13633,N_12917,N_12880);
xor U13634 (N_13634,N_12174,N_12781);
nand U13635 (N_13635,N_12561,N_12460);
nand U13636 (N_13636,N_12525,N_12445);
xor U13637 (N_13637,N_12341,N_12906);
xnor U13638 (N_13638,N_12930,N_12709);
xnor U13639 (N_13639,N_12813,N_12407);
nor U13640 (N_13640,N_12052,N_12126);
xnor U13641 (N_13641,N_12864,N_12565);
or U13642 (N_13642,N_12833,N_12981);
nand U13643 (N_13643,N_12373,N_12695);
or U13644 (N_13644,N_12966,N_12194);
nor U13645 (N_13645,N_12086,N_12859);
or U13646 (N_13646,N_12349,N_12697);
nor U13647 (N_13647,N_12777,N_12478);
and U13648 (N_13648,N_12134,N_12972);
and U13649 (N_13649,N_12821,N_12311);
or U13650 (N_13650,N_12631,N_12602);
or U13651 (N_13651,N_12944,N_12300);
xnor U13652 (N_13652,N_12949,N_12717);
and U13653 (N_13653,N_12924,N_12559);
and U13654 (N_13654,N_12510,N_12798);
or U13655 (N_13655,N_12971,N_12920);
nor U13656 (N_13656,N_12444,N_12174);
or U13657 (N_13657,N_12934,N_12114);
xnor U13658 (N_13658,N_12391,N_12356);
nor U13659 (N_13659,N_12342,N_12225);
nand U13660 (N_13660,N_12336,N_12226);
nand U13661 (N_13661,N_12757,N_12087);
xor U13662 (N_13662,N_12708,N_12595);
xnor U13663 (N_13663,N_12649,N_12536);
nor U13664 (N_13664,N_12487,N_12645);
nand U13665 (N_13665,N_12025,N_12618);
nand U13666 (N_13666,N_12136,N_12184);
nor U13667 (N_13667,N_12777,N_12717);
or U13668 (N_13668,N_12070,N_12340);
nor U13669 (N_13669,N_12131,N_12517);
nand U13670 (N_13670,N_12769,N_12239);
or U13671 (N_13671,N_12933,N_12566);
or U13672 (N_13672,N_12233,N_12730);
nor U13673 (N_13673,N_12531,N_12696);
nor U13674 (N_13674,N_12649,N_12714);
xor U13675 (N_13675,N_12334,N_12883);
nor U13676 (N_13676,N_12563,N_12411);
and U13677 (N_13677,N_12372,N_12775);
or U13678 (N_13678,N_12483,N_12069);
and U13679 (N_13679,N_12641,N_12758);
or U13680 (N_13680,N_12401,N_12041);
xnor U13681 (N_13681,N_12899,N_12940);
nand U13682 (N_13682,N_12654,N_12484);
or U13683 (N_13683,N_12405,N_12482);
or U13684 (N_13684,N_12930,N_12598);
nand U13685 (N_13685,N_12599,N_12622);
nand U13686 (N_13686,N_12957,N_12016);
nand U13687 (N_13687,N_12457,N_12866);
or U13688 (N_13688,N_12014,N_12048);
and U13689 (N_13689,N_12203,N_12494);
or U13690 (N_13690,N_12420,N_12296);
nor U13691 (N_13691,N_12131,N_12214);
nor U13692 (N_13692,N_12983,N_12249);
nand U13693 (N_13693,N_12578,N_12021);
and U13694 (N_13694,N_12026,N_12698);
or U13695 (N_13695,N_12831,N_12854);
nand U13696 (N_13696,N_12052,N_12384);
and U13697 (N_13697,N_12311,N_12805);
nand U13698 (N_13698,N_12953,N_12451);
and U13699 (N_13699,N_12877,N_12841);
nand U13700 (N_13700,N_12056,N_12168);
nand U13701 (N_13701,N_12425,N_12332);
and U13702 (N_13702,N_12696,N_12312);
nor U13703 (N_13703,N_12786,N_12977);
or U13704 (N_13704,N_12806,N_12723);
xor U13705 (N_13705,N_12452,N_12240);
and U13706 (N_13706,N_12558,N_12240);
or U13707 (N_13707,N_12589,N_12014);
nor U13708 (N_13708,N_12593,N_12354);
or U13709 (N_13709,N_12352,N_12383);
and U13710 (N_13710,N_12914,N_12110);
and U13711 (N_13711,N_12646,N_12356);
xor U13712 (N_13712,N_12279,N_12196);
nor U13713 (N_13713,N_12646,N_12068);
and U13714 (N_13714,N_12133,N_12322);
nand U13715 (N_13715,N_12423,N_12853);
nand U13716 (N_13716,N_12313,N_12565);
or U13717 (N_13717,N_12854,N_12560);
and U13718 (N_13718,N_12871,N_12686);
or U13719 (N_13719,N_12285,N_12629);
or U13720 (N_13720,N_12370,N_12950);
nor U13721 (N_13721,N_12517,N_12400);
nand U13722 (N_13722,N_12075,N_12109);
nor U13723 (N_13723,N_12725,N_12002);
and U13724 (N_13724,N_12895,N_12531);
and U13725 (N_13725,N_12723,N_12841);
or U13726 (N_13726,N_12032,N_12007);
nor U13727 (N_13727,N_12451,N_12356);
or U13728 (N_13728,N_12052,N_12210);
and U13729 (N_13729,N_12558,N_12019);
nand U13730 (N_13730,N_12086,N_12617);
nand U13731 (N_13731,N_12287,N_12989);
and U13732 (N_13732,N_12696,N_12666);
and U13733 (N_13733,N_12061,N_12525);
or U13734 (N_13734,N_12983,N_12586);
or U13735 (N_13735,N_12519,N_12033);
nor U13736 (N_13736,N_12202,N_12735);
and U13737 (N_13737,N_12461,N_12932);
xnor U13738 (N_13738,N_12495,N_12534);
xnor U13739 (N_13739,N_12207,N_12107);
nand U13740 (N_13740,N_12468,N_12760);
nand U13741 (N_13741,N_12367,N_12026);
or U13742 (N_13742,N_12824,N_12215);
or U13743 (N_13743,N_12112,N_12476);
nand U13744 (N_13744,N_12914,N_12627);
or U13745 (N_13745,N_12068,N_12384);
or U13746 (N_13746,N_12198,N_12749);
xor U13747 (N_13747,N_12845,N_12936);
nor U13748 (N_13748,N_12293,N_12137);
or U13749 (N_13749,N_12392,N_12647);
or U13750 (N_13750,N_12455,N_12981);
xor U13751 (N_13751,N_12222,N_12630);
nand U13752 (N_13752,N_12739,N_12898);
nand U13753 (N_13753,N_12132,N_12370);
or U13754 (N_13754,N_12266,N_12384);
and U13755 (N_13755,N_12033,N_12786);
or U13756 (N_13756,N_12781,N_12284);
nand U13757 (N_13757,N_12302,N_12181);
and U13758 (N_13758,N_12600,N_12737);
nor U13759 (N_13759,N_12617,N_12595);
nor U13760 (N_13760,N_12186,N_12590);
and U13761 (N_13761,N_12536,N_12360);
nor U13762 (N_13762,N_12981,N_12303);
nand U13763 (N_13763,N_12809,N_12096);
xor U13764 (N_13764,N_12915,N_12232);
or U13765 (N_13765,N_12443,N_12417);
xor U13766 (N_13766,N_12675,N_12288);
nor U13767 (N_13767,N_12840,N_12359);
and U13768 (N_13768,N_12046,N_12823);
or U13769 (N_13769,N_12046,N_12639);
or U13770 (N_13770,N_12255,N_12978);
nor U13771 (N_13771,N_12141,N_12750);
and U13772 (N_13772,N_12435,N_12055);
or U13773 (N_13773,N_12706,N_12560);
and U13774 (N_13774,N_12384,N_12314);
or U13775 (N_13775,N_12800,N_12904);
xor U13776 (N_13776,N_12181,N_12674);
and U13777 (N_13777,N_12781,N_12192);
nor U13778 (N_13778,N_12904,N_12846);
or U13779 (N_13779,N_12377,N_12418);
and U13780 (N_13780,N_12948,N_12059);
or U13781 (N_13781,N_12274,N_12627);
nor U13782 (N_13782,N_12402,N_12901);
nor U13783 (N_13783,N_12203,N_12337);
xor U13784 (N_13784,N_12594,N_12973);
nor U13785 (N_13785,N_12844,N_12228);
xor U13786 (N_13786,N_12495,N_12547);
nor U13787 (N_13787,N_12190,N_12791);
xor U13788 (N_13788,N_12464,N_12705);
or U13789 (N_13789,N_12412,N_12837);
and U13790 (N_13790,N_12777,N_12211);
xor U13791 (N_13791,N_12861,N_12634);
and U13792 (N_13792,N_12964,N_12343);
nand U13793 (N_13793,N_12514,N_12237);
and U13794 (N_13794,N_12251,N_12298);
or U13795 (N_13795,N_12131,N_12437);
and U13796 (N_13796,N_12785,N_12724);
or U13797 (N_13797,N_12959,N_12307);
nor U13798 (N_13798,N_12007,N_12691);
or U13799 (N_13799,N_12257,N_12649);
or U13800 (N_13800,N_12974,N_12965);
and U13801 (N_13801,N_12937,N_12839);
and U13802 (N_13802,N_12250,N_12696);
or U13803 (N_13803,N_12148,N_12223);
and U13804 (N_13804,N_12971,N_12158);
nor U13805 (N_13805,N_12014,N_12815);
or U13806 (N_13806,N_12722,N_12731);
nor U13807 (N_13807,N_12143,N_12259);
and U13808 (N_13808,N_12834,N_12347);
nand U13809 (N_13809,N_12205,N_12848);
or U13810 (N_13810,N_12849,N_12566);
or U13811 (N_13811,N_12883,N_12135);
and U13812 (N_13812,N_12897,N_12059);
or U13813 (N_13813,N_12468,N_12071);
or U13814 (N_13814,N_12828,N_12774);
and U13815 (N_13815,N_12628,N_12202);
nand U13816 (N_13816,N_12986,N_12063);
nor U13817 (N_13817,N_12886,N_12850);
nand U13818 (N_13818,N_12004,N_12699);
or U13819 (N_13819,N_12507,N_12202);
or U13820 (N_13820,N_12275,N_12467);
and U13821 (N_13821,N_12136,N_12117);
nor U13822 (N_13822,N_12027,N_12111);
nor U13823 (N_13823,N_12894,N_12069);
nor U13824 (N_13824,N_12391,N_12372);
xor U13825 (N_13825,N_12892,N_12312);
nand U13826 (N_13826,N_12192,N_12435);
nor U13827 (N_13827,N_12669,N_12371);
xor U13828 (N_13828,N_12264,N_12664);
and U13829 (N_13829,N_12779,N_12614);
xor U13830 (N_13830,N_12948,N_12021);
nand U13831 (N_13831,N_12518,N_12951);
nor U13832 (N_13832,N_12113,N_12790);
nand U13833 (N_13833,N_12164,N_12552);
xor U13834 (N_13834,N_12125,N_12068);
and U13835 (N_13835,N_12781,N_12787);
nand U13836 (N_13836,N_12179,N_12208);
or U13837 (N_13837,N_12393,N_12483);
nor U13838 (N_13838,N_12639,N_12395);
xnor U13839 (N_13839,N_12403,N_12712);
or U13840 (N_13840,N_12567,N_12812);
or U13841 (N_13841,N_12544,N_12103);
nor U13842 (N_13842,N_12767,N_12035);
xor U13843 (N_13843,N_12310,N_12799);
or U13844 (N_13844,N_12013,N_12344);
nand U13845 (N_13845,N_12263,N_12158);
and U13846 (N_13846,N_12033,N_12043);
or U13847 (N_13847,N_12572,N_12192);
or U13848 (N_13848,N_12747,N_12435);
or U13849 (N_13849,N_12296,N_12598);
or U13850 (N_13850,N_12381,N_12868);
or U13851 (N_13851,N_12620,N_12745);
nor U13852 (N_13852,N_12412,N_12406);
nand U13853 (N_13853,N_12463,N_12121);
nor U13854 (N_13854,N_12451,N_12529);
or U13855 (N_13855,N_12544,N_12292);
nand U13856 (N_13856,N_12270,N_12592);
nand U13857 (N_13857,N_12829,N_12526);
nor U13858 (N_13858,N_12878,N_12291);
and U13859 (N_13859,N_12268,N_12415);
and U13860 (N_13860,N_12762,N_12700);
or U13861 (N_13861,N_12558,N_12815);
or U13862 (N_13862,N_12556,N_12365);
or U13863 (N_13863,N_12049,N_12128);
and U13864 (N_13864,N_12425,N_12460);
nand U13865 (N_13865,N_12641,N_12555);
nor U13866 (N_13866,N_12639,N_12919);
or U13867 (N_13867,N_12034,N_12323);
and U13868 (N_13868,N_12219,N_12035);
and U13869 (N_13869,N_12975,N_12516);
and U13870 (N_13870,N_12163,N_12407);
nor U13871 (N_13871,N_12775,N_12999);
or U13872 (N_13872,N_12393,N_12044);
nor U13873 (N_13873,N_12567,N_12482);
nand U13874 (N_13874,N_12985,N_12197);
xnor U13875 (N_13875,N_12752,N_12343);
nand U13876 (N_13876,N_12076,N_12616);
nor U13877 (N_13877,N_12994,N_12687);
nand U13878 (N_13878,N_12310,N_12262);
xor U13879 (N_13879,N_12158,N_12541);
and U13880 (N_13880,N_12309,N_12477);
xnor U13881 (N_13881,N_12526,N_12407);
nor U13882 (N_13882,N_12049,N_12960);
nor U13883 (N_13883,N_12530,N_12793);
nor U13884 (N_13884,N_12169,N_12838);
nor U13885 (N_13885,N_12409,N_12779);
nand U13886 (N_13886,N_12281,N_12668);
or U13887 (N_13887,N_12872,N_12669);
and U13888 (N_13888,N_12967,N_12872);
nand U13889 (N_13889,N_12475,N_12234);
nor U13890 (N_13890,N_12162,N_12818);
nor U13891 (N_13891,N_12494,N_12741);
nor U13892 (N_13892,N_12495,N_12834);
and U13893 (N_13893,N_12732,N_12719);
or U13894 (N_13894,N_12390,N_12964);
nand U13895 (N_13895,N_12195,N_12806);
and U13896 (N_13896,N_12956,N_12055);
nor U13897 (N_13897,N_12973,N_12872);
xnor U13898 (N_13898,N_12524,N_12575);
or U13899 (N_13899,N_12971,N_12967);
nor U13900 (N_13900,N_12218,N_12907);
and U13901 (N_13901,N_12194,N_12130);
or U13902 (N_13902,N_12836,N_12270);
or U13903 (N_13903,N_12227,N_12801);
or U13904 (N_13904,N_12194,N_12283);
nor U13905 (N_13905,N_12095,N_12059);
or U13906 (N_13906,N_12136,N_12016);
or U13907 (N_13907,N_12663,N_12706);
nand U13908 (N_13908,N_12973,N_12708);
nor U13909 (N_13909,N_12184,N_12068);
nand U13910 (N_13910,N_12654,N_12763);
nand U13911 (N_13911,N_12494,N_12622);
and U13912 (N_13912,N_12706,N_12766);
and U13913 (N_13913,N_12354,N_12518);
or U13914 (N_13914,N_12289,N_12151);
or U13915 (N_13915,N_12665,N_12412);
or U13916 (N_13916,N_12646,N_12142);
xnor U13917 (N_13917,N_12875,N_12275);
nand U13918 (N_13918,N_12911,N_12916);
nand U13919 (N_13919,N_12883,N_12938);
xor U13920 (N_13920,N_12663,N_12521);
nand U13921 (N_13921,N_12869,N_12615);
and U13922 (N_13922,N_12416,N_12294);
or U13923 (N_13923,N_12417,N_12546);
and U13924 (N_13924,N_12650,N_12361);
xor U13925 (N_13925,N_12925,N_12692);
and U13926 (N_13926,N_12094,N_12307);
or U13927 (N_13927,N_12990,N_12163);
xor U13928 (N_13928,N_12084,N_12760);
and U13929 (N_13929,N_12743,N_12977);
and U13930 (N_13930,N_12579,N_12827);
nor U13931 (N_13931,N_12257,N_12504);
nor U13932 (N_13932,N_12164,N_12099);
nor U13933 (N_13933,N_12721,N_12928);
or U13934 (N_13934,N_12694,N_12602);
nand U13935 (N_13935,N_12665,N_12601);
or U13936 (N_13936,N_12078,N_12206);
nor U13937 (N_13937,N_12911,N_12852);
nand U13938 (N_13938,N_12405,N_12686);
nand U13939 (N_13939,N_12124,N_12996);
nor U13940 (N_13940,N_12051,N_12251);
nor U13941 (N_13941,N_12114,N_12093);
nand U13942 (N_13942,N_12184,N_12134);
nand U13943 (N_13943,N_12554,N_12485);
xnor U13944 (N_13944,N_12158,N_12258);
nand U13945 (N_13945,N_12877,N_12723);
and U13946 (N_13946,N_12207,N_12266);
nor U13947 (N_13947,N_12731,N_12974);
nand U13948 (N_13948,N_12074,N_12561);
and U13949 (N_13949,N_12058,N_12424);
and U13950 (N_13950,N_12053,N_12787);
nor U13951 (N_13951,N_12325,N_12292);
or U13952 (N_13952,N_12226,N_12229);
or U13953 (N_13953,N_12666,N_12942);
xnor U13954 (N_13954,N_12573,N_12224);
or U13955 (N_13955,N_12620,N_12093);
nor U13956 (N_13956,N_12552,N_12080);
and U13957 (N_13957,N_12493,N_12944);
nand U13958 (N_13958,N_12399,N_12638);
nand U13959 (N_13959,N_12387,N_12843);
and U13960 (N_13960,N_12841,N_12135);
and U13961 (N_13961,N_12067,N_12547);
nor U13962 (N_13962,N_12587,N_12643);
or U13963 (N_13963,N_12998,N_12053);
and U13964 (N_13964,N_12653,N_12034);
or U13965 (N_13965,N_12359,N_12151);
or U13966 (N_13966,N_12702,N_12655);
or U13967 (N_13967,N_12433,N_12711);
nor U13968 (N_13968,N_12523,N_12275);
and U13969 (N_13969,N_12307,N_12983);
nor U13970 (N_13970,N_12344,N_12329);
nand U13971 (N_13971,N_12227,N_12189);
and U13972 (N_13972,N_12621,N_12987);
nor U13973 (N_13973,N_12303,N_12597);
nor U13974 (N_13974,N_12304,N_12995);
nor U13975 (N_13975,N_12541,N_12227);
or U13976 (N_13976,N_12776,N_12795);
and U13977 (N_13977,N_12635,N_12512);
nor U13978 (N_13978,N_12032,N_12936);
or U13979 (N_13979,N_12893,N_12996);
xor U13980 (N_13980,N_12921,N_12797);
nor U13981 (N_13981,N_12412,N_12325);
or U13982 (N_13982,N_12500,N_12327);
and U13983 (N_13983,N_12811,N_12588);
or U13984 (N_13984,N_12497,N_12900);
nand U13985 (N_13985,N_12873,N_12622);
nand U13986 (N_13986,N_12080,N_12133);
nand U13987 (N_13987,N_12916,N_12560);
nand U13988 (N_13988,N_12740,N_12263);
or U13989 (N_13989,N_12554,N_12591);
nand U13990 (N_13990,N_12187,N_12890);
and U13991 (N_13991,N_12283,N_12156);
or U13992 (N_13992,N_12417,N_12548);
and U13993 (N_13993,N_12387,N_12121);
and U13994 (N_13994,N_12865,N_12329);
xnor U13995 (N_13995,N_12524,N_12742);
nand U13996 (N_13996,N_12949,N_12118);
nand U13997 (N_13997,N_12080,N_12009);
xor U13998 (N_13998,N_12930,N_12991);
nor U13999 (N_13999,N_12630,N_12363);
nand U14000 (N_14000,N_13189,N_13628);
xor U14001 (N_14001,N_13792,N_13315);
or U14002 (N_14002,N_13049,N_13329);
or U14003 (N_14003,N_13778,N_13129);
or U14004 (N_14004,N_13516,N_13241);
and U14005 (N_14005,N_13784,N_13080);
nand U14006 (N_14006,N_13703,N_13376);
and U14007 (N_14007,N_13742,N_13253);
and U14008 (N_14008,N_13344,N_13065);
xor U14009 (N_14009,N_13437,N_13165);
and U14010 (N_14010,N_13215,N_13918);
nand U14011 (N_14011,N_13860,N_13578);
and U14012 (N_14012,N_13306,N_13675);
nand U14013 (N_14013,N_13947,N_13436);
nor U14014 (N_14014,N_13530,N_13214);
nor U14015 (N_14015,N_13713,N_13973);
nand U14016 (N_14016,N_13369,N_13154);
nand U14017 (N_14017,N_13445,N_13804);
or U14018 (N_14018,N_13280,N_13272);
and U14019 (N_14019,N_13757,N_13115);
nand U14020 (N_14020,N_13011,N_13102);
xor U14021 (N_14021,N_13554,N_13967);
or U14022 (N_14022,N_13624,N_13463);
nor U14023 (N_14023,N_13796,N_13111);
nand U14024 (N_14024,N_13782,N_13701);
nor U14025 (N_14025,N_13911,N_13205);
xor U14026 (N_14026,N_13119,N_13546);
nand U14027 (N_14027,N_13599,N_13263);
or U14028 (N_14028,N_13970,N_13181);
nor U14029 (N_14029,N_13831,N_13311);
xor U14030 (N_14030,N_13120,N_13723);
nand U14031 (N_14031,N_13951,N_13396);
or U14032 (N_14032,N_13432,N_13333);
nand U14033 (N_14033,N_13319,N_13525);
and U14034 (N_14034,N_13219,N_13190);
xor U14035 (N_14035,N_13191,N_13460);
or U14036 (N_14036,N_13686,N_13337);
nor U14037 (N_14037,N_13922,N_13455);
or U14038 (N_14038,N_13575,N_13729);
nand U14039 (N_14039,N_13381,N_13441);
or U14040 (N_14040,N_13134,N_13290);
and U14041 (N_14041,N_13481,N_13569);
or U14042 (N_14042,N_13946,N_13880);
xor U14043 (N_14043,N_13475,N_13687);
xnor U14044 (N_14044,N_13122,N_13852);
and U14045 (N_14045,N_13987,N_13171);
nand U14046 (N_14046,N_13935,N_13028);
xor U14047 (N_14047,N_13330,N_13461);
nand U14048 (N_14048,N_13513,N_13601);
xor U14049 (N_14049,N_13895,N_13738);
xor U14050 (N_14050,N_13244,N_13885);
and U14051 (N_14051,N_13641,N_13053);
and U14052 (N_14052,N_13638,N_13142);
nand U14053 (N_14053,N_13781,N_13602);
nor U14054 (N_14054,N_13283,N_13303);
nor U14055 (N_14055,N_13137,N_13022);
xnor U14056 (N_14056,N_13741,N_13822);
nor U14057 (N_14057,N_13535,N_13590);
and U14058 (N_14058,N_13487,N_13024);
nor U14059 (N_14059,N_13503,N_13453);
or U14060 (N_14060,N_13767,N_13538);
nand U14061 (N_14061,N_13479,N_13071);
nor U14062 (N_14062,N_13084,N_13281);
xnor U14063 (N_14063,N_13655,N_13710);
nor U14064 (N_14064,N_13013,N_13643);
and U14065 (N_14065,N_13623,N_13884);
nand U14066 (N_14066,N_13220,N_13772);
nand U14067 (N_14067,N_13294,N_13770);
or U14068 (N_14068,N_13609,N_13185);
or U14069 (N_14069,N_13036,N_13667);
or U14070 (N_14070,N_13000,N_13175);
xor U14071 (N_14071,N_13801,N_13485);
or U14072 (N_14072,N_13331,N_13780);
nor U14073 (N_14073,N_13825,N_13360);
nand U14074 (N_14074,N_13188,N_13737);
xnor U14075 (N_14075,N_13228,N_13731);
or U14076 (N_14076,N_13705,N_13978);
or U14077 (N_14077,N_13265,N_13630);
nand U14078 (N_14078,N_13187,N_13876);
and U14079 (N_14079,N_13679,N_13926);
or U14080 (N_14080,N_13902,N_13562);
nand U14081 (N_14081,N_13997,N_13199);
or U14082 (N_14082,N_13786,N_13339);
and U14083 (N_14083,N_13510,N_13894);
nand U14084 (N_14084,N_13541,N_13478);
xor U14085 (N_14085,N_13576,N_13553);
nand U14086 (N_14086,N_13023,N_13358);
nand U14087 (N_14087,N_13332,N_13151);
and U14088 (N_14088,N_13821,N_13979);
xnor U14089 (N_14089,N_13074,N_13431);
nor U14090 (N_14090,N_13616,N_13775);
or U14091 (N_14091,N_13055,N_13100);
nor U14092 (N_14092,N_13140,N_13939);
xor U14093 (N_14093,N_13818,N_13309);
nand U14094 (N_14094,N_13061,N_13328);
and U14095 (N_14095,N_13318,N_13960);
nor U14096 (N_14096,N_13514,N_13052);
xnor U14097 (N_14097,N_13669,N_13813);
or U14098 (N_14098,N_13598,N_13676);
or U14099 (N_14099,N_13378,N_13260);
nor U14100 (N_14100,N_13150,N_13484);
and U14101 (N_14101,N_13982,N_13106);
xor U14102 (N_14102,N_13898,N_13755);
nand U14103 (N_14103,N_13278,N_13949);
and U14104 (N_14104,N_13934,N_13999);
nor U14105 (N_14105,N_13548,N_13744);
nand U14106 (N_14106,N_13101,N_13889);
xnor U14107 (N_14107,N_13844,N_13210);
and U14108 (N_14108,N_13573,N_13783);
nor U14109 (N_14109,N_13537,N_13958);
and U14110 (N_14110,N_13403,N_13651);
or U14111 (N_14111,N_13653,N_13863);
nor U14112 (N_14112,N_13920,N_13501);
or U14113 (N_14113,N_13008,N_13234);
and U14114 (N_14114,N_13787,N_13352);
nor U14115 (N_14115,N_13660,N_13254);
nand U14116 (N_14116,N_13143,N_13625);
nand U14117 (N_14117,N_13005,N_13622);
nand U14118 (N_14118,N_13697,N_13823);
or U14119 (N_14119,N_13093,N_13149);
nand U14120 (N_14120,N_13515,N_13492);
nand U14121 (N_14121,N_13699,N_13502);
and U14122 (N_14122,N_13010,N_13216);
nor U14123 (N_14123,N_13247,N_13488);
and U14124 (N_14124,N_13928,N_13635);
and U14125 (N_14125,N_13275,N_13314);
nand U14126 (N_14126,N_13913,N_13883);
nand U14127 (N_14127,N_13736,N_13159);
nor U14128 (N_14128,N_13932,N_13568);
nand U14129 (N_14129,N_13145,N_13680);
xnor U14130 (N_14130,N_13647,N_13615);
xor U14131 (N_14131,N_13689,N_13419);
and U14132 (N_14132,N_13504,N_13652);
and U14133 (N_14133,N_13245,N_13700);
and U14134 (N_14134,N_13584,N_13449);
nand U14135 (N_14135,N_13843,N_13560);
nand U14136 (N_14136,N_13287,N_13135);
nor U14137 (N_14137,N_13060,N_13415);
nor U14138 (N_14138,N_13972,N_13486);
nor U14139 (N_14139,N_13029,N_13649);
and U14140 (N_14140,N_13961,N_13048);
nor U14141 (N_14141,N_13851,N_13083);
and U14142 (N_14142,N_13289,N_13671);
xor U14143 (N_14143,N_13607,N_13202);
nand U14144 (N_14144,N_13075,N_13917);
xor U14145 (N_14145,N_13046,N_13929);
or U14146 (N_14146,N_13322,N_13659);
and U14147 (N_14147,N_13434,N_13948);
and U14148 (N_14148,N_13092,N_13511);
nand U14149 (N_14149,N_13325,N_13761);
and U14150 (N_14150,N_13520,N_13448);
nor U14151 (N_14151,N_13147,N_13959);
or U14152 (N_14152,N_13994,N_13820);
nand U14153 (N_14153,N_13766,N_13239);
nand U14154 (N_14154,N_13428,N_13802);
or U14155 (N_14155,N_13126,N_13370);
or U14156 (N_14156,N_13062,N_13886);
or U14157 (N_14157,N_13565,N_13237);
or U14158 (N_14158,N_13279,N_13916);
and U14159 (N_14159,N_13853,N_13421);
nand U14160 (N_14160,N_13161,N_13570);
xor U14161 (N_14161,N_13123,N_13809);
nand U14162 (N_14162,N_13042,N_13409);
nand U14163 (N_14163,N_13897,N_13596);
nand U14164 (N_14164,N_13217,N_13855);
or U14165 (N_14165,N_13577,N_13636);
xnor U14166 (N_14166,N_13589,N_13662);
nor U14167 (N_14167,N_13629,N_13976);
or U14168 (N_14168,N_13533,N_13564);
and U14169 (N_14169,N_13079,N_13915);
nor U14170 (N_14170,N_13412,N_13706);
and U14171 (N_14171,N_13580,N_13020);
or U14172 (N_14172,N_13404,N_13373);
or U14173 (N_14173,N_13218,N_13316);
nand U14174 (N_14174,N_13899,N_13238);
nand U14175 (N_14175,N_13176,N_13971);
and U14176 (N_14176,N_13732,N_13034);
nor U14177 (N_14177,N_13206,N_13483);
xnor U14178 (N_14178,N_13387,N_13256);
xnor U14179 (N_14179,N_13534,N_13438);
and U14180 (N_14180,N_13435,N_13201);
and U14181 (N_14181,N_13341,N_13193);
and U14182 (N_14182,N_13167,N_13637);
xor U14183 (N_14183,N_13608,N_13025);
or U14184 (N_14184,N_13940,N_13004);
or U14185 (N_14185,N_13733,N_13019);
nor U14186 (N_14186,N_13800,N_13859);
nor U14187 (N_14187,N_13385,N_13118);
or U14188 (N_14188,N_13454,N_13197);
nor U14189 (N_14189,N_13942,N_13222);
xor U14190 (N_14190,N_13719,N_13849);
nand U14191 (N_14191,N_13944,N_13726);
nand U14192 (N_14192,N_13566,N_13517);
and U14193 (N_14193,N_13743,N_13099);
nor U14194 (N_14194,N_13364,N_13012);
nor U14195 (N_14195,N_13808,N_13847);
and U14196 (N_14196,N_13491,N_13196);
xnor U14197 (N_14197,N_13868,N_13451);
and U14198 (N_14198,N_13368,N_13160);
xnor U14199 (N_14199,N_13021,N_13058);
nor U14200 (N_14200,N_13721,N_13921);
nand U14201 (N_14201,N_13300,N_13054);
nor U14202 (N_14202,N_13184,N_13270);
xnor U14203 (N_14203,N_13712,N_13839);
nor U14204 (N_14204,N_13410,N_13192);
nand U14205 (N_14205,N_13727,N_13108);
and U14206 (N_14206,N_13977,N_13774);
xor U14207 (N_14207,N_13842,N_13871);
nor U14208 (N_14208,N_13363,N_13477);
and U14209 (N_14209,N_13612,N_13420);
or U14210 (N_14210,N_13657,N_13232);
nand U14211 (N_14211,N_13914,N_13925);
nor U14212 (N_14212,N_13026,N_13350);
and U14213 (N_14213,N_13722,N_13696);
nand U14214 (N_14214,N_13450,N_13128);
and U14215 (N_14215,N_13178,N_13704);
and U14216 (N_14216,N_13764,N_13874);
and U14217 (N_14217,N_13073,N_13496);
nand U14218 (N_14218,N_13896,N_13439);
or U14219 (N_14219,N_13776,N_13634);
and U14220 (N_14220,N_13670,N_13457);
or U14221 (N_14221,N_13685,N_13327);
nor U14222 (N_14222,N_13208,N_13295);
or U14223 (N_14223,N_13654,N_13805);
or U14224 (N_14224,N_13811,N_13499);
nand U14225 (N_14225,N_13936,N_13297);
nand U14226 (N_14226,N_13984,N_13963);
nand U14227 (N_14227,N_13398,N_13989);
nor U14228 (N_14228,N_13072,N_13945);
nand U14229 (N_14229,N_13051,N_13550);
or U14230 (N_14230,N_13248,N_13665);
xnor U14231 (N_14231,N_13542,N_13250);
nand U14232 (N_14232,N_13114,N_13267);
xnor U14233 (N_14233,N_13045,N_13257);
xor U14234 (N_14234,N_13347,N_13271);
or U14235 (N_14235,N_13355,N_13954);
nand U14236 (N_14236,N_13169,N_13284);
nand U14237 (N_14237,N_13221,N_13528);
nand U14238 (N_14238,N_13714,N_13383);
nor U14239 (N_14239,N_13644,N_13268);
nand U14240 (N_14240,N_13246,N_13888);
or U14241 (N_14241,N_13207,N_13030);
and U14242 (N_14242,N_13173,N_13837);
nand U14243 (N_14243,N_13305,N_13482);
xnor U14244 (N_14244,N_13240,N_13124);
nand U14245 (N_14245,N_13473,N_13819);
nand U14246 (N_14246,N_13966,N_13224);
nor U14247 (N_14247,N_13139,N_13829);
xnor U14248 (N_14248,N_13050,N_13746);
nand U14249 (N_14249,N_13968,N_13259);
and U14250 (N_14250,N_13426,N_13040);
xor U14251 (N_14251,N_13795,N_13125);
and U14252 (N_14252,N_13867,N_13585);
xor U14253 (N_14253,N_13446,N_13832);
xor U14254 (N_14254,N_13231,N_13090);
and U14255 (N_14255,N_13956,N_13522);
nor U14256 (N_14256,N_13827,N_13291);
and U14257 (N_14257,N_13225,N_13349);
nand U14258 (N_14258,N_13440,N_13172);
or U14259 (N_14259,N_13113,N_13321);
xor U14260 (N_14260,N_13572,N_13198);
and U14261 (N_14261,N_13489,N_13536);
nor U14262 (N_14262,N_13715,N_13174);
and U14263 (N_14263,N_13032,N_13266);
and U14264 (N_14264,N_13866,N_13877);
nor U14265 (N_14265,N_13462,N_13063);
or U14266 (N_14266,N_13433,N_13459);
and U14267 (N_14267,N_13286,N_13262);
xor U14268 (N_14268,N_13312,N_13807);
nand U14269 (N_14269,N_13717,N_13725);
xor U14270 (N_14270,N_13927,N_13027);
and U14271 (N_14271,N_13826,N_13508);
nor U14272 (N_14272,N_13758,N_13393);
and U14273 (N_14273,N_13390,N_13583);
nor U14274 (N_14274,N_13249,N_13044);
nor U14275 (N_14275,N_13518,N_13740);
nor U14276 (N_14276,N_13324,N_13779);
and U14277 (N_14277,N_13177,N_13474);
or U14278 (N_14278,N_13812,N_13739);
or U14279 (N_14279,N_13561,N_13497);
nand U14280 (N_14280,N_13127,N_13116);
nand U14281 (N_14281,N_13833,N_13955);
xnor U14282 (N_14282,N_13226,N_13059);
nor U14283 (N_14283,N_13425,N_13089);
nand U14284 (N_14284,N_13148,N_13632);
or U14285 (N_14285,N_13146,N_13777);
and U14286 (N_14286,N_13892,N_13017);
or U14287 (N_14287,N_13170,N_13708);
xnor U14288 (N_14288,N_13724,N_13552);
and U14289 (N_14289,N_13865,N_13974);
nand U14290 (N_14290,N_13668,N_13557);
nand U14291 (N_14291,N_13138,N_13908);
and U14292 (N_14292,N_13957,N_13422);
nor U14293 (N_14293,N_13862,N_13493);
or U14294 (N_14294,N_13688,N_13941);
nand U14295 (N_14295,N_13698,N_13830);
nor U14296 (N_14296,N_13323,N_13790);
or U14297 (N_14297,N_13748,N_13498);
nor U14298 (N_14298,N_13320,N_13605);
and U14299 (N_14299,N_13338,N_13003);
nor U14300 (N_14300,N_13371,N_13904);
or U14301 (N_14301,N_13751,N_13591);
or U14302 (N_14302,N_13870,N_13788);
nand U14303 (N_14303,N_13069,N_13621);
and U14304 (N_14304,N_13252,N_13658);
nand U14305 (N_14305,N_13693,N_13334);
nor U14306 (N_14306,N_13374,N_13799);
or U14307 (N_14307,N_13543,N_13683);
nor U14308 (N_14308,N_13603,N_13407);
nor U14309 (N_14309,N_13157,N_13563);
nand U14310 (N_14310,N_13836,N_13523);
and U14311 (N_14311,N_13512,N_13179);
and U14312 (N_14312,N_13965,N_13549);
nand U14313 (N_14313,N_13141,N_13233);
xor U14314 (N_14314,N_13923,N_13117);
and U14315 (N_14315,N_13745,N_13472);
and U14316 (N_14316,N_13430,N_13183);
nor U14317 (N_14317,N_13413,N_13351);
or U14318 (N_14318,N_13995,N_13304);
or U14319 (N_14319,N_13586,N_13991);
and U14320 (N_14320,N_13288,N_13136);
nor U14321 (N_14321,N_13937,N_13707);
and U14322 (N_14322,N_13285,N_13856);
and U14323 (N_14323,N_13296,N_13905);
xor U14324 (N_14324,N_13070,N_13845);
nand U14325 (N_14325,N_13131,N_13620);
nand U14326 (N_14326,N_13213,N_13834);
or U14327 (N_14327,N_13105,N_13869);
nand U14328 (N_14328,N_13588,N_13992);
nand U14329 (N_14329,N_13753,N_13469);
or U14330 (N_14330,N_13962,N_13047);
or U14331 (N_14331,N_13597,N_13039);
nand U14332 (N_14332,N_13759,N_13524);
or U14333 (N_14333,N_13816,N_13909);
and U14334 (N_14334,N_13639,N_13919);
and U14335 (N_14335,N_13633,N_13308);
or U14336 (N_14336,N_13640,N_13838);
nor U14337 (N_14337,N_13674,N_13785);
nor U14338 (N_14338,N_13041,N_13365);
or U14339 (N_14339,N_13156,N_13619);
nand U14340 (N_14340,N_13336,N_13545);
nor U14341 (N_14341,N_13692,N_13121);
or U14342 (N_14342,N_13841,N_13529);
and U14343 (N_14343,N_13392,N_13163);
nor U14344 (N_14344,N_13067,N_13212);
nand U14345 (N_14345,N_13002,N_13342);
nor U14346 (N_14346,N_13377,N_13081);
or U14347 (N_14347,N_13646,N_13104);
or U14348 (N_14348,N_13251,N_13112);
nand U14349 (N_14349,N_13875,N_13085);
xor U14350 (N_14350,N_13414,N_13500);
nor U14351 (N_14351,N_13427,N_13153);
nand U14352 (N_14352,N_13872,N_13760);
nor U14353 (N_14353,N_13611,N_13681);
or U14354 (N_14354,N_13155,N_13858);
nor U14355 (N_14355,N_13064,N_13943);
or U14356 (N_14356,N_13815,N_13031);
or U14357 (N_14357,N_13594,N_13677);
nor U14358 (N_14358,N_13879,N_13367);
nor U14359 (N_14359,N_13953,N_13765);
or U14360 (N_14360,N_13107,N_13539);
xor U14361 (N_14361,N_13166,N_13990);
nor U14362 (N_14362,N_13794,N_13702);
nor U14363 (N_14363,N_13103,N_13930);
nand U14364 (N_14364,N_13379,N_13587);
and U14365 (N_14365,N_13521,N_13527);
or U14366 (N_14366,N_13581,N_13035);
or U14367 (N_14367,N_13709,N_13182);
and U14368 (N_14368,N_13903,N_13988);
or U14369 (N_14369,N_13087,N_13227);
xor U14370 (N_14370,N_13718,N_13519);
and U14371 (N_14371,N_13168,N_13993);
nand U14372 (N_14372,N_13292,N_13470);
or U14373 (N_14373,N_13626,N_13223);
nor U14374 (N_14374,N_13933,N_13720);
nor U14375 (N_14375,N_13068,N_13711);
or U14376 (N_14376,N_13400,N_13384);
and U14377 (N_14377,N_13912,N_13057);
nand U14378 (N_14378,N_13195,N_13531);
and U14379 (N_14379,N_13098,N_13269);
nand U14380 (N_14380,N_13204,N_13109);
nand U14381 (N_14381,N_13353,N_13416);
or U14382 (N_14382,N_13797,N_13773);
xnor U14383 (N_14383,N_13684,N_13873);
or U14384 (N_14384,N_13526,N_13540);
xnor U14385 (N_14385,N_13015,N_13273);
and U14386 (N_14386,N_13200,N_13507);
nor U14387 (N_14387,N_13356,N_13018);
nor U14388 (N_14388,N_13411,N_13480);
and U14389 (N_14389,N_13229,N_13924);
or U14390 (N_14390,N_13996,N_13906);
and U14391 (N_14391,N_13769,N_13386);
and U14392 (N_14392,N_13747,N_13734);
nand U14393 (N_14393,N_13037,N_13980);
nor U14394 (N_14394,N_13656,N_13097);
nor U14395 (N_14395,N_13950,N_13985);
nand U14396 (N_14396,N_13394,N_13211);
xor U14397 (N_14397,N_13691,N_13406);
or U14398 (N_14398,N_13354,N_13604);
xnor U14399 (N_14399,N_13806,N_13397);
nand U14400 (N_14400,N_13362,N_13835);
and U14401 (N_14401,N_13900,N_13975);
and U14402 (N_14402,N_13682,N_13828);
or U14403 (N_14403,N_13375,N_13645);
or U14404 (N_14404,N_13348,N_13194);
or U14405 (N_14405,N_13694,N_13133);
nor U14406 (N_14406,N_13673,N_13606);
or U14407 (N_14407,N_13798,N_13763);
or U14408 (N_14408,N_13592,N_13506);
or U14409 (N_14409,N_13901,N_13810);
or U14410 (N_14410,N_13695,N_13361);
nor U14411 (N_14411,N_13261,N_13110);
nand U14412 (N_14412,N_13610,N_13983);
or U14413 (N_14413,N_13094,N_13443);
or U14414 (N_14414,N_13088,N_13582);
and U14415 (N_14415,N_13130,N_13716);
xnor U14416 (N_14416,N_13551,N_13555);
xor U14417 (N_14417,N_13547,N_13310);
nor U14418 (N_14418,N_13840,N_13158);
nor U14419 (N_14419,N_13180,N_13264);
nand U14420 (N_14420,N_13505,N_13299);
and U14421 (N_14421,N_13752,N_13793);
nand U14422 (N_14422,N_13846,N_13490);
xnor U14423 (N_14423,N_13754,N_13442);
and U14424 (N_14424,N_13452,N_13236);
or U14425 (N_14425,N_13335,N_13750);
nand U14426 (N_14426,N_13418,N_13405);
nand U14427 (N_14427,N_13447,N_13007);
nand U14428 (N_14428,N_13313,N_13009);
or U14429 (N_14429,N_13043,N_13399);
and U14430 (N_14430,N_13298,N_13791);
and U14431 (N_14431,N_13476,N_13789);
nand U14432 (N_14432,N_13056,N_13618);
and U14433 (N_14433,N_13817,N_13077);
or U14434 (N_14434,N_13382,N_13952);
or U14435 (N_14435,N_13372,N_13824);
nand U14436 (N_14436,N_13230,N_13209);
nand U14437 (N_14437,N_13650,N_13307);
nor U14438 (N_14438,N_13408,N_13814);
and U14439 (N_14439,N_13661,N_13235);
nand U14440 (N_14440,N_13664,N_13558);
and U14441 (N_14441,N_13891,N_13910);
nor U14442 (N_14442,N_13803,N_13456);
nor U14443 (N_14443,N_13144,N_13850);
xnor U14444 (N_14444,N_13302,N_13340);
and U14445 (N_14445,N_13388,N_13038);
nor U14446 (N_14446,N_13907,N_13465);
nor U14447 (N_14447,N_13678,N_13882);
nand U14448 (N_14448,N_13571,N_13595);
nor U14449 (N_14449,N_13893,N_13878);
or U14450 (N_14450,N_13762,N_13293);
or U14451 (N_14451,N_13672,N_13617);
or U14452 (N_14452,N_13066,N_13986);
or U14453 (N_14453,N_13164,N_13346);
and U14454 (N_14454,N_13642,N_13735);
or U14455 (N_14455,N_13964,N_13544);
nor U14456 (N_14456,N_13317,N_13864);
and U14457 (N_14457,N_13076,N_13391);
or U14458 (N_14458,N_13768,N_13931);
or U14459 (N_14459,N_13468,N_13014);
and U14460 (N_14460,N_13532,N_13969);
and U14461 (N_14461,N_13016,N_13366);
nor U14462 (N_14462,N_13423,N_13756);
and U14463 (N_14463,N_13690,N_13471);
nand U14464 (N_14464,N_13086,N_13091);
or U14465 (N_14465,N_13326,N_13132);
nand U14466 (N_14466,N_13771,N_13359);
xor U14467 (N_14467,N_13495,N_13887);
nor U14468 (N_14468,N_13593,N_13417);
or U14469 (N_14469,N_13627,N_13749);
nand U14470 (N_14470,N_13274,N_13402);
or U14471 (N_14471,N_13401,N_13579);
nand U14472 (N_14472,N_13890,N_13666);
or U14473 (N_14473,N_13881,N_13203);
nand U14474 (N_14474,N_13728,N_13981);
nor U14475 (N_14475,N_13277,N_13600);
nand U14476 (N_14476,N_13006,N_13464);
and U14477 (N_14477,N_13574,N_13648);
nand U14478 (N_14478,N_13082,N_13078);
nand U14479 (N_14479,N_13357,N_13096);
and U14480 (N_14480,N_13395,N_13938);
nand U14481 (N_14481,N_13614,N_13095);
or U14482 (N_14482,N_13631,N_13276);
or U14483 (N_14483,N_13162,N_13255);
or U14484 (N_14484,N_13258,N_13509);
and U14485 (N_14485,N_13857,N_13389);
nand U14486 (N_14486,N_13301,N_13458);
nand U14487 (N_14487,N_13848,N_13282);
or U14488 (N_14488,N_13429,N_13242);
or U14489 (N_14489,N_13001,N_13186);
nor U14490 (N_14490,N_13243,N_13998);
nand U14491 (N_14491,N_13345,N_13033);
nand U14492 (N_14492,N_13424,N_13556);
or U14493 (N_14493,N_13861,N_13494);
nand U14494 (N_14494,N_13567,N_13152);
nand U14495 (N_14495,N_13380,N_13730);
nand U14496 (N_14496,N_13613,N_13467);
and U14497 (N_14497,N_13854,N_13444);
and U14498 (N_14498,N_13663,N_13559);
nand U14499 (N_14499,N_13343,N_13466);
and U14500 (N_14500,N_13961,N_13055);
and U14501 (N_14501,N_13326,N_13003);
and U14502 (N_14502,N_13880,N_13852);
nor U14503 (N_14503,N_13561,N_13836);
xor U14504 (N_14504,N_13482,N_13087);
and U14505 (N_14505,N_13958,N_13405);
and U14506 (N_14506,N_13356,N_13442);
and U14507 (N_14507,N_13937,N_13899);
nor U14508 (N_14508,N_13551,N_13138);
nor U14509 (N_14509,N_13864,N_13933);
or U14510 (N_14510,N_13880,N_13587);
or U14511 (N_14511,N_13971,N_13222);
xor U14512 (N_14512,N_13896,N_13120);
xor U14513 (N_14513,N_13167,N_13584);
and U14514 (N_14514,N_13961,N_13202);
or U14515 (N_14515,N_13610,N_13848);
xnor U14516 (N_14516,N_13943,N_13571);
or U14517 (N_14517,N_13039,N_13767);
or U14518 (N_14518,N_13711,N_13777);
nand U14519 (N_14519,N_13677,N_13380);
nor U14520 (N_14520,N_13955,N_13382);
nand U14521 (N_14521,N_13397,N_13655);
or U14522 (N_14522,N_13176,N_13427);
nand U14523 (N_14523,N_13242,N_13449);
xnor U14524 (N_14524,N_13040,N_13412);
nand U14525 (N_14525,N_13937,N_13210);
and U14526 (N_14526,N_13853,N_13154);
nor U14527 (N_14527,N_13440,N_13785);
xnor U14528 (N_14528,N_13825,N_13408);
nand U14529 (N_14529,N_13862,N_13233);
xor U14530 (N_14530,N_13568,N_13709);
and U14531 (N_14531,N_13539,N_13189);
nor U14532 (N_14532,N_13641,N_13850);
and U14533 (N_14533,N_13083,N_13204);
and U14534 (N_14534,N_13420,N_13725);
nor U14535 (N_14535,N_13413,N_13273);
or U14536 (N_14536,N_13166,N_13279);
and U14537 (N_14537,N_13872,N_13810);
nand U14538 (N_14538,N_13750,N_13278);
xnor U14539 (N_14539,N_13237,N_13873);
or U14540 (N_14540,N_13026,N_13600);
nand U14541 (N_14541,N_13416,N_13522);
nand U14542 (N_14542,N_13101,N_13555);
and U14543 (N_14543,N_13647,N_13707);
nor U14544 (N_14544,N_13459,N_13043);
nand U14545 (N_14545,N_13074,N_13343);
or U14546 (N_14546,N_13684,N_13730);
xnor U14547 (N_14547,N_13432,N_13716);
or U14548 (N_14548,N_13969,N_13010);
and U14549 (N_14549,N_13216,N_13013);
nand U14550 (N_14550,N_13289,N_13811);
nand U14551 (N_14551,N_13495,N_13066);
nor U14552 (N_14552,N_13072,N_13388);
nand U14553 (N_14553,N_13575,N_13274);
xnor U14554 (N_14554,N_13025,N_13452);
nor U14555 (N_14555,N_13679,N_13810);
and U14556 (N_14556,N_13872,N_13942);
or U14557 (N_14557,N_13942,N_13409);
nand U14558 (N_14558,N_13891,N_13269);
or U14559 (N_14559,N_13440,N_13047);
nand U14560 (N_14560,N_13893,N_13320);
xor U14561 (N_14561,N_13527,N_13754);
nor U14562 (N_14562,N_13821,N_13971);
nor U14563 (N_14563,N_13680,N_13942);
and U14564 (N_14564,N_13283,N_13247);
and U14565 (N_14565,N_13153,N_13933);
or U14566 (N_14566,N_13441,N_13969);
or U14567 (N_14567,N_13998,N_13519);
and U14568 (N_14568,N_13971,N_13508);
and U14569 (N_14569,N_13367,N_13489);
nand U14570 (N_14570,N_13915,N_13768);
or U14571 (N_14571,N_13705,N_13519);
or U14572 (N_14572,N_13434,N_13079);
and U14573 (N_14573,N_13647,N_13062);
or U14574 (N_14574,N_13439,N_13224);
nor U14575 (N_14575,N_13118,N_13569);
nand U14576 (N_14576,N_13554,N_13819);
xor U14577 (N_14577,N_13485,N_13911);
nand U14578 (N_14578,N_13255,N_13439);
nand U14579 (N_14579,N_13855,N_13831);
and U14580 (N_14580,N_13586,N_13652);
nand U14581 (N_14581,N_13832,N_13152);
or U14582 (N_14582,N_13936,N_13793);
xor U14583 (N_14583,N_13386,N_13480);
or U14584 (N_14584,N_13782,N_13075);
and U14585 (N_14585,N_13616,N_13030);
and U14586 (N_14586,N_13122,N_13178);
or U14587 (N_14587,N_13439,N_13999);
or U14588 (N_14588,N_13366,N_13663);
and U14589 (N_14589,N_13638,N_13721);
nor U14590 (N_14590,N_13716,N_13554);
and U14591 (N_14591,N_13530,N_13347);
and U14592 (N_14592,N_13666,N_13833);
or U14593 (N_14593,N_13169,N_13546);
or U14594 (N_14594,N_13140,N_13196);
nand U14595 (N_14595,N_13517,N_13500);
and U14596 (N_14596,N_13557,N_13704);
or U14597 (N_14597,N_13565,N_13236);
or U14598 (N_14598,N_13154,N_13764);
nor U14599 (N_14599,N_13819,N_13250);
and U14600 (N_14600,N_13797,N_13025);
nand U14601 (N_14601,N_13697,N_13158);
or U14602 (N_14602,N_13501,N_13993);
nor U14603 (N_14603,N_13273,N_13706);
nor U14604 (N_14604,N_13574,N_13311);
nor U14605 (N_14605,N_13330,N_13798);
or U14606 (N_14606,N_13581,N_13119);
nand U14607 (N_14607,N_13258,N_13172);
or U14608 (N_14608,N_13495,N_13733);
or U14609 (N_14609,N_13613,N_13953);
xor U14610 (N_14610,N_13325,N_13123);
and U14611 (N_14611,N_13044,N_13589);
or U14612 (N_14612,N_13105,N_13480);
and U14613 (N_14613,N_13994,N_13596);
and U14614 (N_14614,N_13617,N_13905);
nor U14615 (N_14615,N_13157,N_13452);
or U14616 (N_14616,N_13738,N_13251);
nor U14617 (N_14617,N_13690,N_13791);
and U14618 (N_14618,N_13492,N_13895);
and U14619 (N_14619,N_13479,N_13765);
or U14620 (N_14620,N_13918,N_13406);
nand U14621 (N_14621,N_13352,N_13950);
and U14622 (N_14622,N_13392,N_13657);
or U14623 (N_14623,N_13142,N_13280);
nand U14624 (N_14624,N_13688,N_13581);
nand U14625 (N_14625,N_13658,N_13701);
nor U14626 (N_14626,N_13112,N_13174);
or U14627 (N_14627,N_13821,N_13326);
nand U14628 (N_14628,N_13417,N_13899);
nand U14629 (N_14629,N_13473,N_13818);
nand U14630 (N_14630,N_13630,N_13354);
nor U14631 (N_14631,N_13919,N_13802);
nand U14632 (N_14632,N_13632,N_13296);
and U14633 (N_14633,N_13046,N_13693);
nand U14634 (N_14634,N_13357,N_13532);
or U14635 (N_14635,N_13690,N_13334);
nand U14636 (N_14636,N_13223,N_13387);
xor U14637 (N_14637,N_13724,N_13075);
and U14638 (N_14638,N_13986,N_13987);
and U14639 (N_14639,N_13013,N_13063);
nor U14640 (N_14640,N_13004,N_13315);
and U14641 (N_14641,N_13037,N_13213);
nor U14642 (N_14642,N_13860,N_13517);
nor U14643 (N_14643,N_13978,N_13316);
xor U14644 (N_14644,N_13049,N_13223);
nor U14645 (N_14645,N_13046,N_13161);
or U14646 (N_14646,N_13464,N_13260);
or U14647 (N_14647,N_13068,N_13647);
and U14648 (N_14648,N_13561,N_13892);
xor U14649 (N_14649,N_13997,N_13805);
and U14650 (N_14650,N_13577,N_13022);
nand U14651 (N_14651,N_13141,N_13831);
nor U14652 (N_14652,N_13089,N_13533);
nor U14653 (N_14653,N_13756,N_13816);
or U14654 (N_14654,N_13573,N_13441);
nor U14655 (N_14655,N_13677,N_13910);
and U14656 (N_14656,N_13819,N_13640);
nor U14657 (N_14657,N_13459,N_13492);
or U14658 (N_14658,N_13763,N_13469);
nand U14659 (N_14659,N_13798,N_13434);
nand U14660 (N_14660,N_13106,N_13354);
and U14661 (N_14661,N_13583,N_13517);
nor U14662 (N_14662,N_13204,N_13893);
nand U14663 (N_14663,N_13604,N_13073);
nor U14664 (N_14664,N_13652,N_13001);
nand U14665 (N_14665,N_13924,N_13210);
and U14666 (N_14666,N_13279,N_13887);
or U14667 (N_14667,N_13484,N_13757);
or U14668 (N_14668,N_13056,N_13778);
or U14669 (N_14669,N_13993,N_13161);
xor U14670 (N_14670,N_13399,N_13607);
or U14671 (N_14671,N_13435,N_13140);
or U14672 (N_14672,N_13394,N_13048);
or U14673 (N_14673,N_13342,N_13707);
nand U14674 (N_14674,N_13330,N_13088);
nor U14675 (N_14675,N_13351,N_13299);
nand U14676 (N_14676,N_13425,N_13630);
and U14677 (N_14677,N_13774,N_13826);
and U14678 (N_14678,N_13450,N_13771);
and U14679 (N_14679,N_13175,N_13685);
or U14680 (N_14680,N_13401,N_13286);
nand U14681 (N_14681,N_13513,N_13987);
or U14682 (N_14682,N_13470,N_13596);
and U14683 (N_14683,N_13157,N_13741);
nand U14684 (N_14684,N_13439,N_13871);
nand U14685 (N_14685,N_13626,N_13988);
nand U14686 (N_14686,N_13650,N_13131);
or U14687 (N_14687,N_13645,N_13825);
and U14688 (N_14688,N_13137,N_13842);
and U14689 (N_14689,N_13639,N_13404);
and U14690 (N_14690,N_13135,N_13413);
nor U14691 (N_14691,N_13810,N_13856);
nand U14692 (N_14692,N_13277,N_13038);
or U14693 (N_14693,N_13574,N_13909);
nand U14694 (N_14694,N_13848,N_13488);
nand U14695 (N_14695,N_13317,N_13368);
or U14696 (N_14696,N_13606,N_13581);
nor U14697 (N_14697,N_13494,N_13446);
or U14698 (N_14698,N_13224,N_13848);
nor U14699 (N_14699,N_13233,N_13966);
and U14700 (N_14700,N_13149,N_13581);
xnor U14701 (N_14701,N_13861,N_13367);
and U14702 (N_14702,N_13151,N_13397);
and U14703 (N_14703,N_13097,N_13014);
and U14704 (N_14704,N_13992,N_13449);
nand U14705 (N_14705,N_13016,N_13561);
nand U14706 (N_14706,N_13506,N_13122);
and U14707 (N_14707,N_13052,N_13447);
and U14708 (N_14708,N_13013,N_13934);
nand U14709 (N_14709,N_13319,N_13420);
nor U14710 (N_14710,N_13151,N_13242);
nor U14711 (N_14711,N_13880,N_13172);
nor U14712 (N_14712,N_13791,N_13110);
or U14713 (N_14713,N_13059,N_13596);
or U14714 (N_14714,N_13511,N_13121);
nand U14715 (N_14715,N_13736,N_13629);
nor U14716 (N_14716,N_13880,N_13559);
and U14717 (N_14717,N_13740,N_13998);
and U14718 (N_14718,N_13475,N_13446);
nor U14719 (N_14719,N_13339,N_13226);
nor U14720 (N_14720,N_13087,N_13221);
nand U14721 (N_14721,N_13480,N_13540);
and U14722 (N_14722,N_13499,N_13187);
nor U14723 (N_14723,N_13283,N_13232);
and U14724 (N_14724,N_13616,N_13895);
nand U14725 (N_14725,N_13413,N_13368);
and U14726 (N_14726,N_13545,N_13618);
and U14727 (N_14727,N_13012,N_13391);
or U14728 (N_14728,N_13000,N_13636);
nand U14729 (N_14729,N_13435,N_13543);
nand U14730 (N_14730,N_13169,N_13562);
nand U14731 (N_14731,N_13929,N_13828);
nor U14732 (N_14732,N_13457,N_13451);
nand U14733 (N_14733,N_13989,N_13331);
or U14734 (N_14734,N_13991,N_13526);
or U14735 (N_14735,N_13752,N_13697);
or U14736 (N_14736,N_13944,N_13861);
and U14737 (N_14737,N_13456,N_13657);
nor U14738 (N_14738,N_13727,N_13976);
xor U14739 (N_14739,N_13021,N_13280);
and U14740 (N_14740,N_13370,N_13071);
or U14741 (N_14741,N_13221,N_13545);
nor U14742 (N_14742,N_13846,N_13965);
and U14743 (N_14743,N_13411,N_13639);
or U14744 (N_14744,N_13163,N_13617);
nor U14745 (N_14745,N_13586,N_13703);
or U14746 (N_14746,N_13820,N_13856);
nand U14747 (N_14747,N_13736,N_13532);
xnor U14748 (N_14748,N_13166,N_13604);
nand U14749 (N_14749,N_13341,N_13075);
nand U14750 (N_14750,N_13555,N_13939);
or U14751 (N_14751,N_13119,N_13284);
nand U14752 (N_14752,N_13953,N_13961);
or U14753 (N_14753,N_13061,N_13561);
nor U14754 (N_14754,N_13143,N_13315);
and U14755 (N_14755,N_13017,N_13475);
and U14756 (N_14756,N_13090,N_13350);
or U14757 (N_14757,N_13091,N_13672);
nand U14758 (N_14758,N_13087,N_13674);
or U14759 (N_14759,N_13464,N_13820);
nand U14760 (N_14760,N_13032,N_13602);
xor U14761 (N_14761,N_13482,N_13265);
and U14762 (N_14762,N_13325,N_13104);
or U14763 (N_14763,N_13047,N_13728);
xor U14764 (N_14764,N_13169,N_13229);
nor U14765 (N_14765,N_13066,N_13106);
nand U14766 (N_14766,N_13925,N_13186);
and U14767 (N_14767,N_13227,N_13190);
nor U14768 (N_14768,N_13089,N_13883);
nor U14769 (N_14769,N_13147,N_13878);
or U14770 (N_14770,N_13072,N_13956);
and U14771 (N_14771,N_13351,N_13711);
and U14772 (N_14772,N_13102,N_13092);
nand U14773 (N_14773,N_13434,N_13577);
nor U14774 (N_14774,N_13062,N_13463);
and U14775 (N_14775,N_13905,N_13574);
and U14776 (N_14776,N_13919,N_13669);
nor U14777 (N_14777,N_13766,N_13670);
or U14778 (N_14778,N_13153,N_13770);
nor U14779 (N_14779,N_13177,N_13129);
nor U14780 (N_14780,N_13251,N_13877);
or U14781 (N_14781,N_13164,N_13404);
and U14782 (N_14782,N_13312,N_13064);
or U14783 (N_14783,N_13627,N_13957);
nor U14784 (N_14784,N_13912,N_13205);
nand U14785 (N_14785,N_13749,N_13842);
nor U14786 (N_14786,N_13699,N_13601);
nand U14787 (N_14787,N_13290,N_13817);
and U14788 (N_14788,N_13749,N_13191);
xor U14789 (N_14789,N_13676,N_13753);
xnor U14790 (N_14790,N_13717,N_13138);
and U14791 (N_14791,N_13919,N_13281);
or U14792 (N_14792,N_13004,N_13869);
xor U14793 (N_14793,N_13430,N_13982);
or U14794 (N_14794,N_13431,N_13455);
nor U14795 (N_14795,N_13211,N_13418);
nand U14796 (N_14796,N_13471,N_13234);
and U14797 (N_14797,N_13716,N_13219);
or U14798 (N_14798,N_13368,N_13470);
or U14799 (N_14799,N_13141,N_13797);
or U14800 (N_14800,N_13666,N_13727);
or U14801 (N_14801,N_13087,N_13374);
nor U14802 (N_14802,N_13231,N_13215);
or U14803 (N_14803,N_13288,N_13235);
and U14804 (N_14804,N_13625,N_13513);
nand U14805 (N_14805,N_13748,N_13685);
and U14806 (N_14806,N_13246,N_13448);
nor U14807 (N_14807,N_13929,N_13708);
or U14808 (N_14808,N_13460,N_13340);
nor U14809 (N_14809,N_13975,N_13804);
or U14810 (N_14810,N_13078,N_13532);
nand U14811 (N_14811,N_13852,N_13340);
nor U14812 (N_14812,N_13305,N_13536);
nor U14813 (N_14813,N_13182,N_13990);
nand U14814 (N_14814,N_13383,N_13444);
nor U14815 (N_14815,N_13358,N_13986);
nand U14816 (N_14816,N_13752,N_13416);
nand U14817 (N_14817,N_13037,N_13185);
xnor U14818 (N_14818,N_13779,N_13036);
nand U14819 (N_14819,N_13323,N_13727);
xnor U14820 (N_14820,N_13984,N_13385);
nor U14821 (N_14821,N_13141,N_13404);
nor U14822 (N_14822,N_13306,N_13757);
and U14823 (N_14823,N_13575,N_13413);
or U14824 (N_14824,N_13771,N_13476);
xnor U14825 (N_14825,N_13715,N_13315);
and U14826 (N_14826,N_13425,N_13485);
or U14827 (N_14827,N_13189,N_13414);
and U14828 (N_14828,N_13767,N_13641);
or U14829 (N_14829,N_13930,N_13544);
or U14830 (N_14830,N_13968,N_13497);
or U14831 (N_14831,N_13990,N_13043);
nand U14832 (N_14832,N_13112,N_13039);
and U14833 (N_14833,N_13388,N_13441);
and U14834 (N_14834,N_13423,N_13521);
or U14835 (N_14835,N_13164,N_13683);
xor U14836 (N_14836,N_13371,N_13430);
and U14837 (N_14837,N_13271,N_13590);
nor U14838 (N_14838,N_13554,N_13941);
or U14839 (N_14839,N_13599,N_13163);
or U14840 (N_14840,N_13655,N_13362);
or U14841 (N_14841,N_13025,N_13724);
or U14842 (N_14842,N_13673,N_13866);
nor U14843 (N_14843,N_13598,N_13378);
or U14844 (N_14844,N_13823,N_13190);
and U14845 (N_14845,N_13940,N_13745);
nand U14846 (N_14846,N_13316,N_13308);
nor U14847 (N_14847,N_13841,N_13198);
xor U14848 (N_14848,N_13959,N_13423);
or U14849 (N_14849,N_13238,N_13012);
nand U14850 (N_14850,N_13180,N_13044);
or U14851 (N_14851,N_13558,N_13441);
and U14852 (N_14852,N_13972,N_13639);
and U14853 (N_14853,N_13789,N_13644);
and U14854 (N_14854,N_13296,N_13982);
nor U14855 (N_14855,N_13937,N_13927);
nor U14856 (N_14856,N_13613,N_13639);
and U14857 (N_14857,N_13301,N_13335);
and U14858 (N_14858,N_13420,N_13614);
nor U14859 (N_14859,N_13911,N_13220);
or U14860 (N_14860,N_13587,N_13603);
or U14861 (N_14861,N_13674,N_13567);
nor U14862 (N_14862,N_13837,N_13916);
or U14863 (N_14863,N_13959,N_13712);
nor U14864 (N_14864,N_13473,N_13972);
or U14865 (N_14865,N_13046,N_13417);
xnor U14866 (N_14866,N_13837,N_13689);
nand U14867 (N_14867,N_13972,N_13009);
and U14868 (N_14868,N_13978,N_13120);
nand U14869 (N_14869,N_13297,N_13864);
and U14870 (N_14870,N_13060,N_13713);
nor U14871 (N_14871,N_13310,N_13500);
nor U14872 (N_14872,N_13515,N_13587);
nor U14873 (N_14873,N_13984,N_13476);
or U14874 (N_14874,N_13186,N_13376);
nor U14875 (N_14875,N_13753,N_13258);
nand U14876 (N_14876,N_13662,N_13957);
xor U14877 (N_14877,N_13149,N_13567);
nand U14878 (N_14878,N_13031,N_13665);
and U14879 (N_14879,N_13585,N_13260);
nand U14880 (N_14880,N_13399,N_13736);
nor U14881 (N_14881,N_13748,N_13433);
xor U14882 (N_14882,N_13805,N_13209);
nor U14883 (N_14883,N_13293,N_13967);
or U14884 (N_14884,N_13742,N_13657);
or U14885 (N_14885,N_13392,N_13725);
nand U14886 (N_14886,N_13741,N_13519);
or U14887 (N_14887,N_13333,N_13687);
nor U14888 (N_14888,N_13237,N_13255);
nand U14889 (N_14889,N_13043,N_13085);
nand U14890 (N_14890,N_13550,N_13960);
nor U14891 (N_14891,N_13809,N_13604);
nor U14892 (N_14892,N_13714,N_13283);
nand U14893 (N_14893,N_13107,N_13728);
nand U14894 (N_14894,N_13903,N_13691);
nor U14895 (N_14895,N_13399,N_13135);
and U14896 (N_14896,N_13526,N_13223);
nand U14897 (N_14897,N_13714,N_13440);
and U14898 (N_14898,N_13382,N_13465);
nor U14899 (N_14899,N_13783,N_13942);
or U14900 (N_14900,N_13203,N_13237);
xnor U14901 (N_14901,N_13806,N_13906);
nand U14902 (N_14902,N_13524,N_13178);
or U14903 (N_14903,N_13668,N_13111);
and U14904 (N_14904,N_13395,N_13345);
or U14905 (N_14905,N_13167,N_13604);
nor U14906 (N_14906,N_13855,N_13893);
and U14907 (N_14907,N_13882,N_13884);
nor U14908 (N_14908,N_13410,N_13399);
nor U14909 (N_14909,N_13792,N_13255);
or U14910 (N_14910,N_13838,N_13645);
nand U14911 (N_14911,N_13109,N_13230);
xor U14912 (N_14912,N_13721,N_13580);
nor U14913 (N_14913,N_13038,N_13292);
or U14914 (N_14914,N_13156,N_13456);
nand U14915 (N_14915,N_13371,N_13325);
nand U14916 (N_14916,N_13039,N_13010);
nor U14917 (N_14917,N_13913,N_13569);
and U14918 (N_14918,N_13818,N_13648);
nor U14919 (N_14919,N_13588,N_13154);
xnor U14920 (N_14920,N_13731,N_13304);
or U14921 (N_14921,N_13481,N_13997);
and U14922 (N_14922,N_13674,N_13224);
xnor U14923 (N_14923,N_13042,N_13349);
and U14924 (N_14924,N_13633,N_13870);
or U14925 (N_14925,N_13102,N_13563);
or U14926 (N_14926,N_13730,N_13340);
or U14927 (N_14927,N_13218,N_13736);
nand U14928 (N_14928,N_13686,N_13689);
or U14929 (N_14929,N_13589,N_13256);
or U14930 (N_14930,N_13724,N_13719);
nand U14931 (N_14931,N_13822,N_13478);
or U14932 (N_14932,N_13328,N_13315);
nand U14933 (N_14933,N_13208,N_13024);
and U14934 (N_14934,N_13552,N_13458);
nor U14935 (N_14935,N_13029,N_13193);
nor U14936 (N_14936,N_13081,N_13733);
or U14937 (N_14937,N_13517,N_13764);
or U14938 (N_14938,N_13688,N_13969);
nor U14939 (N_14939,N_13358,N_13565);
xnor U14940 (N_14940,N_13882,N_13954);
and U14941 (N_14941,N_13188,N_13886);
or U14942 (N_14942,N_13328,N_13176);
xor U14943 (N_14943,N_13996,N_13517);
nor U14944 (N_14944,N_13723,N_13350);
xnor U14945 (N_14945,N_13868,N_13275);
nand U14946 (N_14946,N_13052,N_13673);
and U14947 (N_14947,N_13612,N_13238);
nor U14948 (N_14948,N_13713,N_13104);
and U14949 (N_14949,N_13752,N_13935);
nor U14950 (N_14950,N_13688,N_13103);
or U14951 (N_14951,N_13191,N_13375);
and U14952 (N_14952,N_13479,N_13470);
or U14953 (N_14953,N_13455,N_13995);
or U14954 (N_14954,N_13019,N_13237);
and U14955 (N_14955,N_13223,N_13366);
nor U14956 (N_14956,N_13720,N_13965);
nor U14957 (N_14957,N_13649,N_13496);
nor U14958 (N_14958,N_13964,N_13841);
nor U14959 (N_14959,N_13242,N_13857);
nand U14960 (N_14960,N_13620,N_13326);
and U14961 (N_14961,N_13587,N_13657);
xor U14962 (N_14962,N_13193,N_13898);
nor U14963 (N_14963,N_13574,N_13316);
xnor U14964 (N_14964,N_13667,N_13139);
or U14965 (N_14965,N_13732,N_13417);
or U14966 (N_14966,N_13420,N_13967);
nor U14967 (N_14967,N_13326,N_13221);
xor U14968 (N_14968,N_13896,N_13856);
nand U14969 (N_14969,N_13996,N_13518);
nand U14970 (N_14970,N_13354,N_13041);
nand U14971 (N_14971,N_13800,N_13767);
or U14972 (N_14972,N_13487,N_13462);
or U14973 (N_14973,N_13618,N_13771);
or U14974 (N_14974,N_13280,N_13170);
nor U14975 (N_14975,N_13561,N_13111);
or U14976 (N_14976,N_13362,N_13871);
nor U14977 (N_14977,N_13416,N_13392);
xor U14978 (N_14978,N_13615,N_13599);
and U14979 (N_14979,N_13539,N_13170);
and U14980 (N_14980,N_13922,N_13577);
or U14981 (N_14981,N_13313,N_13428);
or U14982 (N_14982,N_13357,N_13717);
nor U14983 (N_14983,N_13969,N_13142);
and U14984 (N_14984,N_13996,N_13460);
and U14985 (N_14985,N_13312,N_13519);
and U14986 (N_14986,N_13861,N_13781);
nor U14987 (N_14987,N_13407,N_13461);
or U14988 (N_14988,N_13117,N_13710);
nand U14989 (N_14989,N_13357,N_13535);
and U14990 (N_14990,N_13674,N_13384);
and U14991 (N_14991,N_13996,N_13798);
nor U14992 (N_14992,N_13150,N_13577);
and U14993 (N_14993,N_13366,N_13883);
nand U14994 (N_14994,N_13229,N_13482);
nor U14995 (N_14995,N_13365,N_13873);
nand U14996 (N_14996,N_13300,N_13105);
or U14997 (N_14997,N_13751,N_13214);
nor U14998 (N_14998,N_13317,N_13990);
nor U14999 (N_14999,N_13921,N_13023);
and U15000 (N_15000,N_14985,N_14566);
and U15001 (N_15001,N_14604,N_14622);
nand U15002 (N_15002,N_14461,N_14044);
nand U15003 (N_15003,N_14617,N_14971);
or U15004 (N_15004,N_14955,N_14561);
nor U15005 (N_15005,N_14261,N_14924);
and U15006 (N_15006,N_14089,N_14518);
xor U15007 (N_15007,N_14655,N_14212);
or U15008 (N_15008,N_14587,N_14628);
or U15009 (N_15009,N_14595,N_14147);
nor U15010 (N_15010,N_14373,N_14359);
and U15011 (N_15011,N_14805,N_14228);
and U15012 (N_15012,N_14412,N_14739);
xnor U15013 (N_15013,N_14432,N_14774);
nor U15014 (N_15014,N_14603,N_14366);
nor U15015 (N_15015,N_14682,N_14067);
nor U15016 (N_15016,N_14811,N_14039);
nand U15017 (N_15017,N_14717,N_14351);
nor U15018 (N_15018,N_14681,N_14876);
and U15019 (N_15019,N_14640,N_14736);
nand U15020 (N_15020,N_14095,N_14542);
and U15021 (N_15021,N_14941,N_14426);
and U15022 (N_15022,N_14685,N_14154);
nor U15023 (N_15023,N_14288,N_14517);
nand U15024 (N_15024,N_14970,N_14792);
and U15025 (N_15025,N_14043,N_14114);
and U15026 (N_15026,N_14176,N_14397);
and U15027 (N_15027,N_14350,N_14045);
or U15028 (N_15028,N_14890,N_14661);
nand U15029 (N_15029,N_14605,N_14883);
nand U15030 (N_15030,N_14205,N_14135);
or U15031 (N_15031,N_14762,N_14945);
and U15032 (N_15032,N_14156,N_14149);
nor U15033 (N_15033,N_14014,N_14490);
nand U15034 (N_15034,N_14112,N_14384);
xor U15035 (N_15035,N_14338,N_14694);
nor U15036 (N_15036,N_14400,N_14979);
nand U15037 (N_15037,N_14069,N_14578);
nor U15038 (N_15038,N_14751,N_14616);
and U15039 (N_15039,N_14191,N_14047);
or U15040 (N_15040,N_14683,N_14544);
xnor U15041 (N_15041,N_14989,N_14269);
nor U15042 (N_15042,N_14497,N_14250);
nor U15043 (N_15043,N_14464,N_14447);
xnor U15044 (N_15044,N_14865,N_14009);
or U15045 (N_15045,N_14200,N_14433);
nand U15046 (N_15046,N_14032,N_14963);
and U15047 (N_15047,N_14019,N_14054);
nor U15048 (N_15048,N_14056,N_14732);
or U15049 (N_15049,N_14806,N_14455);
and U15050 (N_15050,N_14829,N_14998);
xor U15051 (N_15051,N_14379,N_14652);
nand U15052 (N_15052,N_14743,N_14697);
nand U15053 (N_15053,N_14253,N_14127);
and U15054 (N_15054,N_14003,N_14365);
xnor U15055 (N_15055,N_14631,N_14966);
or U15056 (N_15056,N_14050,N_14020);
nand U15057 (N_15057,N_14040,N_14929);
nor U15058 (N_15058,N_14860,N_14823);
or U15059 (N_15059,N_14656,N_14415);
or U15060 (N_15060,N_14104,N_14825);
nand U15061 (N_15061,N_14268,N_14363);
or U15062 (N_15062,N_14841,N_14568);
or U15063 (N_15063,N_14778,N_14265);
and U15064 (N_15064,N_14611,N_14010);
nand U15065 (N_15065,N_14348,N_14718);
or U15066 (N_15066,N_14651,N_14458);
nor U15067 (N_15067,N_14678,N_14887);
nand U15068 (N_15068,N_14575,N_14668);
nand U15069 (N_15069,N_14911,N_14745);
and U15070 (N_15070,N_14724,N_14788);
and U15071 (N_15071,N_14569,N_14689);
and U15072 (N_15072,N_14030,N_14466);
nand U15073 (N_15073,N_14082,N_14999);
and U15074 (N_15074,N_14336,N_14385);
xor U15075 (N_15075,N_14078,N_14192);
and U15076 (N_15076,N_14870,N_14353);
nand U15077 (N_15077,N_14435,N_14297);
and U15078 (N_15078,N_14693,N_14165);
nand U15079 (N_15079,N_14706,N_14310);
and U15080 (N_15080,N_14535,N_14854);
and U15081 (N_15081,N_14133,N_14878);
nor U15082 (N_15082,N_14645,N_14898);
and U15083 (N_15083,N_14637,N_14311);
nor U15084 (N_15084,N_14317,N_14711);
nor U15085 (N_15085,N_14855,N_14824);
and U15086 (N_15086,N_14534,N_14958);
and U15087 (N_15087,N_14072,N_14565);
and U15088 (N_15088,N_14766,N_14839);
nand U15089 (N_15089,N_14388,N_14660);
nor U15090 (N_15090,N_14287,N_14741);
xor U15091 (N_15091,N_14413,N_14822);
xor U15092 (N_15092,N_14123,N_14048);
nand U15093 (N_15093,N_14756,N_14814);
and U15094 (N_15094,N_14601,N_14174);
and U15095 (N_15095,N_14233,N_14781);
nand U15096 (N_15096,N_14041,N_14467);
and U15097 (N_15097,N_14757,N_14635);
nand U15098 (N_15098,N_14273,N_14333);
or U15099 (N_15099,N_14438,N_14213);
nor U15100 (N_15100,N_14921,N_14579);
nor U15101 (N_15101,N_14916,N_14161);
xnor U15102 (N_15102,N_14527,N_14627);
nand U15103 (N_15103,N_14471,N_14117);
nand U15104 (N_15104,N_14593,N_14832);
nand U15105 (N_15105,N_14794,N_14139);
and U15106 (N_15106,N_14239,N_14722);
or U15107 (N_15107,N_14007,N_14952);
xnor U15108 (N_15108,N_14264,N_14267);
nand U15109 (N_15109,N_14763,N_14073);
nand U15110 (N_15110,N_14087,N_14562);
or U15111 (N_15111,N_14896,N_14177);
or U15112 (N_15112,N_14111,N_14153);
nor U15113 (N_15113,N_14961,N_14529);
or U15114 (N_15114,N_14000,N_14479);
or U15115 (N_15115,N_14653,N_14609);
nor U15116 (N_15116,N_14893,N_14892);
and U15117 (N_15117,N_14954,N_14801);
and U15118 (N_15118,N_14209,N_14394);
nand U15119 (N_15119,N_14528,N_14217);
and U15120 (N_15120,N_14299,N_14767);
nor U15121 (N_15121,N_14874,N_14437);
nand U15122 (N_15122,N_14137,N_14096);
or U15123 (N_15123,N_14973,N_14950);
xor U15124 (N_15124,N_14118,N_14244);
or U15125 (N_15125,N_14122,N_14863);
or U15126 (N_15126,N_14821,N_14807);
xor U15127 (N_15127,N_14158,N_14417);
nand U15128 (N_15128,N_14439,N_14367);
or U15129 (N_15129,N_14580,N_14771);
and U15130 (N_15130,N_14939,N_14733);
nor U15131 (N_15131,N_14016,N_14493);
xor U15132 (N_15132,N_14060,N_14028);
or U15133 (N_15133,N_14869,N_14754);
and U15134 (N_15134,N_14484,N_14818);
or U15135 (N_15135,N_14589,N_14620);
nand U15136 (N_15136,N_14335,N_14401);
nand U15137 (N_15137,N_14830,N_14967);
nand U15138 (N_15138,N_14877,N_14583);
nor U15139 (N_15139,N_14769,N_14422);
nand U15140 (N_15140,N_14386,N_14431);
and U15141 (N_15141,N_14483,N_14959);
nand U15142 (N_15142,N_14256,N_14225);
nor U15143 (N_15143,N_14902,N_14926);
or U15144 (N_15144,N_14790,N_14364);
nand U15145 (N_15145,N_14782,N_14468);
xnor U15146 (N_15146,N_14899,N_14234);
nand U15147 (N_15147,N_14708,N_14163);
nand U15148 (N_15148,N_14884,N_14404);
nor U15149 (N_15149,N_14615,N_14211);
and U15150 (N_15150,N_14731,N_14251);
nand U15151 (N_15151,N_14626,N_14465);
nor U15152 (N_15152,N_14787,N_14563);
nand U15153 (N_15153,N_14880,N_14453);
or U15154 (N_15154,N_14679,N_14195);
nor U15155 (N_15155,N_14423,N_14015);
nor U15156 (N_15156,N_14285,N_14456);
or U15157 (N_15157,N_14242,N_14889);
and U15158 (N_15158,N_14026,N_14850);
xnor U15159 (N_15159,N_14927,N_14198);
nand U15160 (N_15160,N_14337,N_14314);
and U15161 (N_15161,N_14935,N_14215);
nor U15162 (N_15162,N_14813,N_14725);
xor U15163 (N_15163,N_14940,N_14917);
nand U15164 (N_15164,N_14900,N_14291);
nand U15165 (N_15165,N_14537,N_14512);
and U15166 (N_15166,N_14546,N_14738);
and U15167 (N_15167,N_14946,N_14101);
nor U15168 (N_15168,N_14735,N_14383);
nor U15169 (N_15169,N_14129,N_14862);
nor U15170 (N_15170,N_14796,N_14108);
and U15171 (N_15171,N_14474,N_14675);
and U15172 (N_15172,N_14840,N_14776);
or U15173 (N_15173,N_14765,N_14551);
xor U15174 (N_15174,N_14875,N_14584);
nand U15175 (N_15175,N_14986,N_14308);
nand U15176 (N_15176,N_14282,N_14306);
nor U15177 (N_15177,N_14925,N_14643);
or U15178 (N_15178,N_14714,N_14956);
nand U15179 (N_15179,N_14070,N_14360);
xor U15180 (N_15180,N_14328,N_14799);
nand U15181 (N_15181,N_14064,N_14614);
nand U15182 (N_15182,N_14023,N_14919);
nand U15183 (N_15183,N_14340,N_14276);
nor U15184 (N_15184,N_14298,N_14157);
and U15185 (N_15185,N_14719,N_14936);
and U15186 (N_15186,N_14079,N_14930);
nor U15187 (N_15187,N_14085,N_14221);
and U15188 (N_15188,N_14241,N_14904);
or U15189 (N_15189,N_14820,N_14457);
nand U15190 (N_15190,N_14271,N_14399);
or U15191 (N_15191,N_14463,N_14196);
xnor U15192 (N_15192,N_14076,N_14151);
or U15193 (N_15193,N_14744,N_14393);
nand U15194 (N_15194,N_14978,N_14120);
nand U15195 (N_15195,N_14031,N_14646);
or U15196 (N_15196,N_14402,N_14560);
and U15197 (N_15197,N_14644,N_14789);
and U15198 (N_15198,N_14503,N_14886);
and U15199 (N_15199,N_14380,N_14508);
xor U15200 (N_15200,N_14342,N_14664);
nand U15201 (N_15201,N_14006,N_14038);
xnor U15202 (N_15202,N_14968,N_14747);
nand U15203 (N_15203,N_14301,N_14779);
or U15204 (N_15204,N_14427,N_14696);
nor U15205 (N_15205,N_14548,N_14347);
nor U15206 (N_15206,N_14356,N_14894);
and U15207 (N_15207,N_14487,N_14680);
or U15208 (N_15208,N_14831,N_14424);
xor U15209 (N_15209,N_14057,N_14169);
nand U15210 (N_15210,N_14376,N_14444);
xor U15211 (N_15211,N_14785,N_14881);
xor U15212 (N_15212,N_14141,N_14784);
and U15213 (N_15213,N_14526,N_14252);
nor U15214 (N_15214,N_14477,N_14663);
nand U15215 (N_15215,N_14642,N_14915);
and U15216 (N_15216,N_14525,N_14473);
nor U15217 (N_15217,N_14100,N_14633);
or U15218 (N_15218,N_14327,N_14027);
and U15219 (N_15219,N_14549,N_14266);
and U15220 (N_15220,N_14770,N_14737);
nor U15221 (N_15221,N_14649,N_14772);
xor U15222 (N_15222,N_14172,N_14819);
nor U15223 (N_15223,N_14980,N_14852);
nor U15224 (N_15224,N_14879,N_14223);
nand U15225 (N_15225,N_14944,N_14080);
or U15226 (N_15226,N_14795,N_14091);
nor U15227 (N_15227,N_14075,N_14488);
or U15228 (N_15228,N_14341,N_14606);
nor U15229 (N_15229,N_14931,N_14933);
or U15230 (N_15230,N_14699,N_14222);
and U15231 (N_15231,N_14843,N_14109);
nor U15232 (N_15232,N_14318,N_14844);
xnor U15233 (N_15233,N_14816,N_14349);
and U15234 (N_15234,N_14270,N_14996);
nor U15235 (N_15235,N_14472,N_14764);
nor U15236 (N_15236,N_14184,N_14476);
nand U15237 (N_15237,N_14144,N_14160);
or U15238 (N_15238,N_14025,N_14146);
nor U15239 (N_15239,N_14389,N_14613);
and U15240 (N_15240,N_14511,N_14375);
nor U15241 (N_15241,N_14257,N_14330);
xnor U15242 (N_15242,N_14331,N_14313);
nand U15243 (N_15243,N_14136,N_14909);
or U15244 (N_15244,N_14247,N_14309);
nand U15245 (N_15245,N_14937,N_14409);
nand U15246 (N_15246,N_14168,N_14533);
or U15247 (N_15247,N_14938,N_14037);
nand U15248 (N_15248,N_14752,N_14868);
nor U15249 (N_15249,N_14162,N_14254);
nand U15250 (N_15250,N_14964,N_14066);
or U15251 (N_15251,N_14035,N_14543);
and U15252 (N_15252,N_14240,N_14284);
and U15253 (N_15253,N_14235,N_14428);
xor U15254 (N_15254,N_14536,N_14110);
nand U15255 (N_15255,N_14873,N_14758);
nor U15256 (N_15256,N_14290,N_14629);
or U15257 (N_15257,N_14849,N_14063);
nor U15258 (N_15258,N_14748,N_14498);
nand U15259 (N_15259,N_14024,N_14932);
or U15260 (N_15260,N_14173,N_14429);
nor U15261 (N_15261,N_14703,N_14071);
nor U15262 (N_15262,N_14214,N_14179);
xnor U15263 (N_15263,N_14665,N_14727);
and U15264 (N_15264,N_14740,N_14332);
nor U15265 (N_15265,N_14227,N_14126);
and U15266 (N_15266,N_14322,N_14407);
nand U15267 (N_15267,N_14815,N_14289);
nand U15268 (N_15268,N_14055,N_14210);
or U15269 (N_15269,N_14326,N_14410);
nor U15270 (N_15270,N_14155,N_14791);
nand U15271 (N_15271,N_14721,N_14051);
nor U15272 (N_15272,N_14346,N_14405);
nor U15273 (N_15273,N_14775,N_14572);
nand U15274 (N_15274,N_14278,N_14371);
xnor U15275 (N_15275,N_14293,N_14499);
or U15276 (N_15276,N_14545,N_14654);
nand U15277 (N_15277,N_14238,N_14053);
nor U15278 (N_15278,N_14159,N_14838);
nor U15279 (N_15279,N_14848,N_14442);
nor U15280 (N_15280,N_14965,N_14369);
xor U15281 (N_15281,N_14103,N_14559);
or U15282 (N_15282,N_14768,N_14279);
and U15283 (N_15283,N_14042,N_14475);
and U15284 (N_15284,N_14142,N_14555);
nand U15285 (N_15285,N_14062,N_14382);
or U15286 (N_15286,N_14530,N_14029);
and U15287 (N_15287,N_14856,N_14190);
xnor U15288 (N_15288,N_14670,N_14864);
nor U15289 (N_15289,N_14761,N_14125);
and U15290 (N_15290,N_14590,N_14505);
or U15291 (N_15291,N_14345,N_14093);
or U15292 (N_15292,N_14218,N_14907);
nand U15293 (N_15293,N_14470,N_14510);
and U15294 (N_15294,N_14962,N_14182);
or U15295 (N_15295,N_14166,N_14502);
and U15296 (N_15296,N_14321,N_14358);
nor U15297 (N_15297,N_14283,N_14418);
xor U15298 (N_15298,N_14734,N_14099);
nor U15299 (N_15299,N_14630,N_14115);
and U15300 (N_15300,N_14574,N_14325);
nor U15301 (N_15301,N_14836,N_14280);
xor U15302 (N_15302,N_14598,N_14374);
or U15303 (N_15303,N_14355,N_14391);
xor U15304 (N_15304,N_14181,N_14798);
nand U15305 (N_15305,N_14690,N_14920);
or U15306 (N_15306,N_14846,N_14012);
or U15307 (N_15307,N_14454,N_14459);
nand U15308 (N_15308,N_14199,N_14632);
nor U15309 (N_15309,N_14949,N_14094);
nor U15310 (N_15310,N_14312,N_14912);
or U15311 (N_15311,N_14914,N_14552);
nor U15312 (N_15312,N_14148,N_14713);
xor U15313 (N_15313,N_14988,N_14203);
nand U15314 (N_15314,N_14485,N_14107);
nor U15315 (N_15315,N_14004,N_14677);
nand U15316 (N_15316,N_14990,N_14084);
nand U15317 (N_15317,N_14102,N_14403);
nor U15318 (N_15318,N_14581,N_14853);
nand U15319 (N_15319,N_14249,N_14582);
or U15320 (N_15320,N_14842,N_14749);
nor U15321 (N_15321,N_14150,N_14793);
and U15322 (N_15322,N_14259,N_14550);
or U15323 (N_15323,N_14197,N_14494);
nor U15324 (N_15324,N_14729,N_14170);
xnor U15325 (N_15325,N_14092,N_14116);
nor U15326 (N_15326,N_14372,N_14204);
or U15327 (N_15327,N_14258,N_14134);
nand U15328 (N_15328,N_14515,N_14274);
and U15329 (N_15329,N_14845,N_14777);
nor U15330 (N_15330,N_14540,N_14208);
xor U15331 (N_15331,N_14378,N_14597);
nand U15332 (N_15332,N_14891,N_14726);
nor U15333 (N_15333,N_14928,N_14232);
and U15334 (N_15334,N_14976,N_14220);
xor U15335 (N_15335,N_14230,N_14621);
nor U15336 (N_15336,N_14531,N_14707);
or U15337 (N_15337,N_14065,N_14411);
and U15338 (N_15338,N_14647,N_14994);
nor U15339 (N_15339,N_14804,N_14128);
nand U15340 (N_15340,N_14387,N_14984);
or U15341 (N_15341,N_14421,N_14316);
xor U15342 (N_15342,N_14524,N_14702);
nor U15343 (N_15343,N_14482,N_14178);
and U15344 (N_15344,N_14462,N_14624);
or U15345 (N_15345,N_14648,N_14608);
nor U15346 (N_15346,N_14594,N_14339);
nor U15347 (N_15347,N_14202,N_14913);
nand U15348 (N_15348,N_14507,N_14357);
and U15349 (N_15349,N_14728,N_14618);
nor U15350 (N_15350,N_14828,N_14716);
nor U15351 (N_15351,N_14720,N_14687);
and U15352 (N_15352,N_14833,N_14918);
nand U15353 (N_15353,N_14755,N_14121);
and U15354 (N_15354,N_14957,N_14674);
xnor U15355 (N_15355,N_14760,N_14903);
or U15356 (N_15356,N_14263,N_14676);
and U15357 (N_15357,N_14558,N_14923);
or U15358 (N_15358,N_14446,N_14977);
xor U15359 (N_15359,N_14396,N_14034);
and U15360 (N_15360,N_14077,N_14292);
and U15361 (N_15361,N_14539,N_14231);
or U15362 (N_15362,N_14324,N_14882);
nor U15363 (N_15363,N_14319,N_14827);
or U15364 (N_15364,N_14478,N_14296);
or U15365 (N_15365,N_14942,N_14623);
or U15366 (N_15366,N_14599,N_14492);
or U15367 (N_15367,N_14090,N_14248);
nand U15368 (N_15368,N_14398,N_14395);
nor U15369 (N_15369,N_14885,N_14186);
xnor U15370 (N_15370,N_14783,N_14557);
nor U15371 (N_15371,N_14180,N_14119);
or U15372 (N_15372,N_14897,N_14859);
and U15373 (N_15373,N_14011,N_14858);
nor U15374 (N_15374,N_14036,N_14362);
and U15375 (N_15375,N_14381,N_14895);
nand U15376 (N_15376,N_14612,N_14753);
or U15377 (N_15377,N_14246,N_14408);
and U15378 (N_15378,N_14553,N_14260);
and U15379 (N_15379,N_14152,N_14450);
nand U15380 (N_15380,N_14504,N_14206);
nand U15381 (N_15381,N_14097,N_14997);
nand U15382 (N_15382,N_14377,N_14441);
nand U15383 (N_15383,N_14495,N_14586);
nand U15384 (N_15384,N_14835,N_14294);
or U15385 (N_15385,N_14607,N_14547);
and U15386 (N_15386,N_14662,N_14201);
and U15387 (N_15387,N_14803,N_14698);
nand U15388 (N_15388,N_14780,N_14981);
nand U15389 (N_15389,N_14255,N_14052);
nor U15390 (N_15390,N_14138,N_14513);
nand U15391 (N_15391,N_14443,N_14419);
nor U15392 (N_15392,N_14773,N_14320);
and U15393 (N_15393,N_14851,N_14817);
nand U15394 (N_15394,N_14684,N_14344);
nor U15395 (N_15395,N_14207,N_14081);
nand U15396 (N_15396,N_14295,N_14216);
or U15397 (N_15397,N_14974,N_14519);
nand U15398 (N_15398,N_14390,N_14002);
nor U15399 (N_15399,N_14183,N_14812);
or U15400 (N_15400,N_14500,N_14947);
or U15401 (N_15401,N_14641,N_14837);
nor U15402 (N_15402,N_14658,N_14602);
nand U15403 (N_15403,N_14434,N_14591);
xnor U15404 (N_15404,N_14995,N_14448);
nand U15405 (N_15405,N_14742,N_14871);
and U15406 (N_15406,N_14709,N_14808);
and U15407 (N_15407,N_14969,N_14489);
or U15408 (N_15408,N_14867,N_14866);
nor U15409 (N_15409,N_14522,N_14991);
or U15410 (N_15410,N_14625,N_14619);
and U15411 (N_15411,N_14786,N_14420);
and U15412 (N_15412,N_14700,N_14021);
nand U15413 (N_15413,N_14514,N_14068);
nor U15414 (N_15414,N_14993,N_14059);
nand U15415 (N_15415,N_14538,N_14236);
nor U15416 (N_15416,N_14826,N_14541);
and U15417 (N_15417,N_14224,N_14281);
and U15418 (N_15418,N_14074,N_14600);
nand U15419 (N_15419,N_14520,N_14272);
nor U15420 (N_15420,N_14809,N_14307);
or U15421 (N_15421,N_14746,N_14303);
nor U15422 (N_15422,N_14573,N_14008);
nand U15423 (N_15423,N_14140,N_14592);
nand U15424 (N_15424,N_14577,N_14334);
xor U15425 (N_15425,N_14960,N_14229);
nor U15426 (N_15426,N_14800,N_14667);
nand U15427 (N_15427,N_14975,N_14650);
nand U15428 (N_15428,N_14452,N_14343);
or U15429 (N_15429,N_14521,N_14953);
nand U15430 (N_15430,N_14414,N_14124);
nand U15431 (N_15431,N_14810,N_14673);
nand U15432 (N_15432,N_14275,N_14797);
and U15433 (N_15433,N_14571,N_14449);
or U15434 (N_15434,N_14083,N_14516);
or U15435 (N_15435,N_14058,N_14486);
or U15436 (N_15436,N_14130,N_14901);
nor U15437 (N_15437,N_14370,N_14657);
nor U15438 (N_15438,N_14802,N_14509);
and U15439 (N_15439,N_14132,N_14834);
and U15440 (N_15440,N_14392,N_14175);
xor U15441 (N_15441,N_14688,N_14469);
nor U15442 (N_15442,N_14910,N_14033);
or U15443 (N_15443,N_14430,N_14013);
and U15444 (N_15444,N_14145,N_14302);
nand U15445 (N_15445,N_14634,N_14329);
or U15446 (N_15446,N_14193,N_14934);
and U15447 (N_15447,N_14857,N_14368);
or U15448 (N_15448,N_14872,N_14022);
nor U15449 (N_15449,N_14323,N_14596);
or U15450 (N_15450,N_14445,N_14245);
or U15451 (N_15451,N_14481,N_14906);
or U15452 (N_15452,N_14639,N_14086);
and U15453 (N_15453,N_14691,N_14187);
nand U15454 (N_15454,N_14219,N_14304);
nand U15455 (N_15455,N_14352,N_14106);
or U15456 (N_15456,N_14046,N_14987);
nand U15457 (N_15457,N_14460,N_14567);
or U15458 (N_15458,N_14672,N_14088);
nor U15459 (N_15459,N_14948,N_14188);
nand U15460 (N_15460,N_14712,N_14436);
nand U15461 (N_15461,N_14723,N_14972);
nor U15462 (N_15462,N_14610,N_14554);
nand U15463 (N_15463,N_14710,N_14659);
and U15464 (N_15464,N_14237,N_14226);
and U15465 (N_15465,N_14440,N_14638);
and U15466 (N_15466,N_14564,N_14570);
or U15467 (N_15467,N_14262,N_14983);
and U15468 (N_15468,N_14185,N_14705);
or U15469 (N_15469,N_14686,N_14523);
nor U15470 (N_15470,N_14354,N_14704);
or U15471 (N_15471,N_14425,N_14701);
nand U15472 (N_15472,N_14113,N_14532);
and U15473 (N_15473,N_14105,N_14361);
nand U15474 (N_15474,N_14005,N_14194);
nand U15475 (N_15475,N_14189,N_14556);
nor U15476 (N_15476,N_14847,N_14300);
and U15477 (N_15477,N_14451,N_14061);
and U15478 (N_15478,N_14861,N_14001);
or U15479 (N_15479,N_14669,N_14131);
or U15480 (N_15480,N_14506,N_14908);
or U15481 (N_15481,N_14585,N_14406);
nand U15482 (N_15482,N_14171,N_14491);
nor U15483 (N_15483,N_14098,N_14695);
and U15484 (N_15484,N_14164,N_14286);
and U15485 (N_15485,N_14277,N_14049);
nand U15486 (N_15486,N_14480,N_14576);
or U15487 (N_15487,N_14315,N_14666);
nor U15488 (N_15488,N_14692,N_14167);
or U15489 (N_15489,N_14715,N_14496);
nor U15490 (N_15490,N_14588,N_14636);
or U15491 (N_15491,N_14501,N_14888);
and U15492 (N_15492,N_14922,N_14905);
nand U15493 (N_15493,N_14750,N_14759);
or U15494 (N_15494,N_14143,N_14671);
nor U15495 (N_15495,N_14017,N_14982);
and U15496 (N_15496,N_14730,N_14243);
and U15497 (N_15497,N_14943,N_14992);
or U15498 (N_15498,N_14018,N_14416);
nor U15499 (N_15499,N_14951,N_14305);
nand U15500 (N_15500,N_14133,N_14489);
and U15501 (N_15501,N_14201,N_14652);
nand U15502 (N_15502,N_14880,N_14232);
nand U15503 (N_15503,N_14179,N_14188);
and U15504 (N_15504,N_14467,N_14986);
nand U15505 (N_15505,N_14542,N_14995);
nand U15506 (N_15506,N_14529,N_14112);
or U15507 (N_15507,N_14107,N_14147);
nand U15508 (N_15508,N_14892,N_14583);
and U15509 (N_15509,N_14223,N_14091);
or U15510 (N_15510,N_14902,N_14152);
nor U15511 (N_15511,N_14492,N_14278);
and U15512 (N_15512,N_14342,N_14602);
or U15513 (N_15513,N_14243,N_14835);
xor U15514 (N_15514,N_14563,N_14449);
xor U15515 (N_15515,N_14305,N_14704);
xnor U15516 (N_15516,N_14190,N_14353);
nor U15517 (N_15517,N_14422,N_14471);
nand U15518 (N_15518,N_14347,N_14812);
or U15519 (N_15519,N_14450,N_14918);
nand U15520 (N_15520,N_14272,N_14218);
or U15521 (N_15521,N_14494,N_14928);
and U15522 (N_15522,N_14895,N_14732);
nor U15523 (N_15523,N_14654,N_14005);
nor U15524 (N_15524,N_14535,N_14818);
nor U15525 (N_15525,N_14796,N_14402);
nor U15526 (N_15526,N_14329,N_14389);
or U15527 (N_15527,N_14929,N_14437);
and U15528 (N_15528,N_14511,N_14835);
or U15529 (N_15529,N_14851,N_14401);
nor U15530 (N_15530,N_14824,N_14225);
or U15531 (N_15531,N_14095,N_14534);
and U15532 (N_15532,N_14069,N_14128);
or U15533 (N_15533,N_14655,N_14191);
or U15534 (N_15534,N_14951,N_14242);
and U15535 (N_15535,N_14339,N_14784);
nor U15536 (N_15536,N_14462,N_14369);
and U15537 (N_15537,N_14838,N_14327);
and U15538 (N_15538,N_14114,N_14812);
and U15539 (N_15539,N_14489,N_14329);
nand U15540 (N_15540,N_14395,N_14706);
nor U15541 (N_15541,N_14387,N_14162);
and U15542 (N_15542,N_14363,N_14777);
nand U15543 (N_15543,N_14001,N_14110);
or U15544 (N_15544,N_14884,N_14388);
nand U15545 (N_15545,N_14267,N_14282);
and U15546 (N_15546,N_14581,N_14325);
nor U15547 (N_15547,N_14410,N_14546);
xor U15548 (N_15548,N_14297,N_14152);
and U15549 (N_15549,N_14330,N_14047);
nor U15550 (N_15550,N_14139,N_14822);
and U15551 (N_15551,N_14101,N_14272);
nand U15552 (N_15552,N_14235,N_14919);
nand U15553 (N_15553,N_14875,N_14323);
nor U15554 (N_15554,N_14536,N_14746);
or U15555 (N_15555,N_14110,N_14951);
and U15556 (N_15556,N_14260,N_14338);
or U15557 (N_15557,N_14291,N_14697);
nor U15558 (N_15558,N_14661,N_14676);
or U15559 (N_15559,N_14267,N_14370);
or U15560 (N_15560,N_14192,N_14764);
nor U15561 (N_15561,N_14419,N_14336);
xor U15562 (N_15562,N_14765,N_14934);
and U15563 (N_15563,N_14728,N_14015);
or U15564 (N_15564,N_14948,N_14970);
xnor U15565 (N_15565,N_14657,N_14724);
nand U15566 (N_15566,N_14560,N_14140);
or U15567 (N_15567,N_14981,N_14548);
and U15568 (N_15568,N_14860,N_14921);
or U15569 (N_15569,N_14669,N_14014);
nand U15570 (N_15570,N_14427,N_14831);
nor U15571 (N_15571,N_14459,N_14089);
or U15572 (N_15572,N_14890,N_14371);
or U15573 (N_15573,N_14552,N_14908);
or U15574 (N_15574,N_14047,N_14117);
and U15575 (N_15575,N_14367,N_14519);
nand U15576 (N_15576,N_14365,N_14327);
nor U15577 (N_15577,N_14048,N_14814);
or U15578 (N_15578,N_14037,N_14935);
nor U15579 (N_15579,N_14468,N_14997);
nand U15580 (N_15580,N_14178,N_14841);
nand U15581 (N_15581,N_14717,N_14455);
nand U15582 (N_15582,N_14234,N_14678);
nand U15583 (N_15583,N_14067,N_14704);
xor U15584 (N_15584,N_14726,N_14654);
or U15585 (N_15585,N_14027,N_14783);
xnor U15586 (N_15586,N_14954,N_14895);
xor U15587 (N_15587,N_14412,N_14789);
or U15588 (N_15588,N_14092,N_14611);
xnor U15589 (N_15589,N_14145,N_14539);
nand U15590 (N_15590,N_14180,N_14545);
or U15591 (N_15591,N_14328,N_14916);
xnor U15592 (N_15592,N_14640,N_14180);
nand U15593 (N_15593,N_14407,N_14502);
and U15594 (N_15594,N_14731,N_14703);
nand U15595 (N_15595,N_14505,N_14053);
and U15596 (N_15596,N_14409,N_14987);
and U15597 (N_15597,N_14673,N_14815);
and U15598 (N_15598,N_14495,N_14964);
nand U15599 (N_15599,N_14061,N_14332);
xor U15600 (N_15600,N_14688,N_14244);
xnor U15601 (N_15601,N_14959,N_14671);
and U15602 (N_15602,N_14468,N_14118);
and U15603 (N_15603,N_14529,N_14793);
nand U15604 (N_15604,N_14433,N_14903);
nand U15605 (N_15605,N_14852,N_14540);
and U15606 (N_15606,N_14876,N_14813);
or U15607 (N_15607,N_14406,N_14774);
and U15608 (N_15608,N_14372,N_14327);
or U15609 (N_15609,N_14195,N_14585);
nor U15610 (N_15610,N_14950,N_14408);
and U15611 (N_15611,N_14984,N_14351);
and U15612 (N_15612,N_14170,N_14321);
nand U15613 (N_15613,N_14834,N_14832);
nand U15614 (N_15614,N_14417,N_14807);
nor U15615 (N_15615,N_14060,N_14952);
and U15616 (N_15616,N_14910,N_14824);
xnor U15617 (N_15617,N_14647,N_14030);
xor U15618 (N_15618,N_14801,N_14482);
and U15619 (N_15619,N_14149,N_14256);
and U15620 (N_15620,N_14840,N_14593);
or U15621 (N_15621,N_14838,N_14871);
or U15622 (N_15622,N_14068,N_14796);
nor U15623 (N_15623,N_14974,N_14766);
or U15624 (N_15624,N_14746,N_14581);
and U15625 (N_15625,N_14960,N_14627);
and U15626 (N_15626,N_14701,N_14982);
nand U15627 (N_15627,N_14063,N_14536);
nand U15628 (N_15628,N_14160,N_14536);
and U15629 (N_15629,N_14477,N_14560);
nor U15630 (N_15630,N_14573,N_14430);
nand U15631 (N_15631,N_14834,N_14397);
nand U15632 (N_15632,N_14932,N_14604);
nand U15633 (N_15633,N_14647,N_14730);
nor U15634 (N_15634,N_14324,N_14532);
nand U15635 (N_15635,N_14683,N_14353);
and U15636 (N_15636,N_14769,N_14811);
and U15637 (N_15637,N_14727,N_14614);
xor U15638 (N_15638,N_14828,N_14929);
or U15639 (N_15639,N_14574,N_14288);
xnor U15640 (N_15640,N_14195,N_14923);
and U15641 (N_15641,N_14887,N_14764);
nor U15642 (N_15642,N_14731,N_14007);
or U15643 (N_15643,N_14516,N_14520);
and U15644 (N_15644,N_14172,N_14048);
nor U15645 (N_15645,N_14412,N_14595);
nor U15646 (N_15646,N_14595,N_14688);
nor U15647 (N_15647,N_14105,N_14624);
nand U15648 (N_15648,N_14579,N_14685);
and U15649 (N_15649,N_14668,N_14631);
nor U15650 (N_15650,N_14350,N_14337);
nor U15651 (N_15651,N_14359,N_14133);
or U15652 (N_15652,N_14832,N_14926);
nand U15653 (N_15653,N_14804,N_14379);
and U15654 (N_15654,N_14947,N_14338);
nor U15655 (N_15655,N_14149,N_14893);
nor U15656 (N_15656,N_14289,N_14538);
and U15657 (N_15657,N_14693,N_14489);
and U15658 (N_15658,N_14615,N_14691);
nand U15659 (N_15659,N_14460,N_14033);
and U15660 (N_15660,N_14450,N_14933);
or U15661 (N_15661,N_14425,N_14112);
or U15662 (N_15662,N_14451,N_14644);
nand U15663 (N_15663,N_14456,N_14357);
xor U15664 (N_15664,N_14615,N_14148);
nand U15665 (N_15665,N_14614,N_14918);
nand U15666 (N_15666,N_14553,N_14529);
nand U15667 (N_15667,N_14634,N_14069);
and U15668 (N_15668,N_14885,N_14977);
nand U15669 (N_15669,N_14418,N_14185);
nand U15670 (N_15670,N_14928,N_14585);
xor U15671 (N_15671,N_14334,N_14043);
nor U15672 (N_15672,N_14756,N_14343);
and U15673 (N_15673,N_14848,N_14521);
and U15674 (N_15674,N_14567,N_14357);
xor U15675 (N_15675,N_14455,N_14983);
nand U15676 (N_15676,N_14706,N_14401);
nor U15677 (N_15677,N_14616,N_14808);
and U15678 (N_15678,N_14266,N_14489);
or U15679 (N_15679,N_14563,N_14351);
and U15680 (N_15680,N_14008,N_14236);
or U15681 (N_15681,N_14325,N_14620);
or U15682 (N_15682,N_14914,N_14963);
nor U15683 (N_15683,N_14414,N_14616);
or U15684 (N_15684,N_14921,N_14557);
nor U15685 (N_15685,N_14757,N_14284);
nor U15686 (N_15686,N_14028,N_14620);
xnor U15687 (N_15687,N_14734,N_14481);
xor U15688 (N_15688,N_14851,N_14162);
nor U15689 (N_15689,N_14577,N_14547);
and U15690 (N_15690,N_14985,N_14640);
xnor U15691 (N_15691,N_14967,N_14341);
nand U15692 (N_15692,N_14229,N_14660);
nand U15693 (N_15693,N_14311,N_14010);
and U15694 (N_15694,N_14902,N_14944);
nand U15695 (N_15695,N_14773,N_14120);
nand U15696 (N_15696,N_14484,N_14765);
and U15697 (N_15697,N_14075,N_14403);
nor U15698 (N_15698,N_14384,N_14327);
or U15699 (N_15699,N_14608,N_14664);
and U15700 (N_15700,N_14316,N_14582);
nor U15701 (N_15701,N_14612,N_14374);
nor U15702 (N_15702,N_14449,N_14846);
nor U15703 (N_15703,N_14602,N_14005);
nand U15704 (N_15704,N_14738,N_14057);
nor U15705 (N_15705,N_14022,N_14068);
or U15706 (N_15706,N_14740,N_14616);
and U15707 (N_15707,N_14171,N_14149);
nor U15708 (N_15708,N_14077,N_14369);
or U15709 (N_15709,N_14016,N_14405);
nand U15710 (N_15710,N_14879,N_14904);
nor U15711 (N_15711,N_14321,N_14428);
xor U15712 (N_15712,N_14310,N_14927);
nand U15713 (N_15713,N_14553,N_14512);
nand U15714 (N_15714,N_14447,N_14458);
or U15715 (N_15715,N_14917,N_14519);
nand U15716 (N_15716,N_14379,N_14527);
or U15717 (N_15717,N_14426,N_14335);
nand U15718 (N_15718,N_14730,N_14775);
nor U15719 (N_15719,N_14690,N_14648);
nor U15720 (N_15720,N_14816,N_14568);
and U15721 (N_15721,N_14536,N_14686);
nor U15722 (N_15722,N_14001,N_14205);
xor U15723 (N_15723,N_14124,N_14049);
nor U15724 (N_15724,N_14683,N_14711);
nand U15725 (N_15725,N_14294,N_14189);
nor U15726 (N_15726,N_14066,N_14128);
or U15727 (N_15727,N_14357,N_14101);
nor U15728 (N_15728,N_14092,N_14013);
nand U15729 (N_15729,N_14837,N_14895);
nand U15730 (N_15730,N_14593,N_14818);
nand U15731 (N_15731,N_14900,N_14864);
and U15732 (N_15732,N_14644,N_14469);
nor U15733 (N_15733,N_14097,N_14571);
or U15734 (N_15734,N_14920,N_14828);
nor U15735 (N_15735,N_14568,N_14303);
nand U15736 (N_15736,N_14698,N_14374);
and U15737 (N_15737,N_14632,N_14132);
or U15738 (N_15738,N_14331,N_14379);
and U15739 (N_15739,N_14638,N_14512);
and U15740 (N_15740,N_14113,N_14744);
or U15741 (N_15741,N_14286,N_14730);
nand U15742 (N_15742,N_14108,N_14183);
and U15743 (N_15743,N_14905,N_14030);
or U15744 (N_15744,N_14341,N_14865);
nand U15745 (N_15745,N_14199,N_14349);
nand U15746 (N_15746,N_14990,N_14532);
nand U15747 (N_15747,N_14648,N_14065);
nor U15748 (N_15748,N_14886,N_14797);
nor U15749 (N_15749,N_14207,N_14523);
nor U15750 (N_15750,N_14187,N_14734);
nand U15751 (N_15751,N_14832,N_14392);
or U15752 (N_15752,N_14849,N_14227);
or U15753 (N_15753,N_14552,N_14911);
nand U15754 (N_15754,N_14101,N_14528);
xor U15755 (N_15755,N_14895,N_14943);
and U15756 (N_15756,N_14122,N_14993);
nor U15757 (N_15757,N_14803,N_14628);
nand U15758 (N_15758,N_14379,N_14797);
or U15759 (N_15759,N_14122,N_14833);
xor U15760 (N_15760,N_14766,N_14767);
nand U15761 (N_15761,N_14732,N_14710);
nand U15762 (N_15762,N_14200,N_14429);
and U15763 (N_15763,N_14424,N_14579);
xor U15764 (N_15764,N_14032,N_14345);
or U15765 (N_15765,N_14196,N_14205);
or U15766 (N_15766,N_14003,N_14727);
and U15767 (N_15767,N_14562,N_14428);
xnor U15768 (N_15768,N_14924,N_14146);
and U15769 (N_15769,N_14936,N_14488);
or U15770 (N_15770,N_14176,N_14868);
nand U15771 (N_15771,N_14827,N_14279);
nor U15772 (N_15772,N_14143,N_14372);
or U15773 (N_15773,N_14810,N_14627);
nand U15774 (N_15774,N_14188,N_14293);
or U15775 (N_15775,N_14670,N_14853);
nand U15776 (N_15776,N_14403,N_14460);
nor U15777 (N_15777,N_14155,N_14824);
nor U15778 (N_15778,N_14067,N_14463);
nor U15779 (N_15779,N_14170,N_14934);
xor U15780 (N_15780,N_14755,N_14800);
nor U15781 (N_15781,N_14181,N_14439);
nor U15782 (N_15782,N_14418,N_14067);
nor U15783 (N_15783,N_14821,N_14590);
nand U15784 (N_15784,N_14177,N_14844);
nand U15785 (N_15785,N_14813,N_14441);
nand U15786 (N_15786,N_14864,N_14080);
xor U15787 (N_15787,N_14625,N_14374);
or U15788 (N_15788,N_14087,N_14962);
or U15789 (N_15789,N_14480,N_14737);
nor U15790 (N_15790,N_14316,N_14008);
nand U15791 (N_15791,N_14508,N_14215);
or U15792 (N_15792,N_14513,N_14002);
and U15793 (N_15793,N_14548,N_14825);
nand U15794 (N_15794,N_14255,N_14469);
and U15795 (N_15795,N_14314,N_14002);
or U15796 (N_15796,N_14912,N_14899);
or U15797 (N_15797,N_14108,N_14623);
or U15798 (N_15798,N_14028,N_14445);
and U15799 (N_15799,N_14330,N_14254);
nor U15800 (N_15800,N_14111,N_14520);
and U15801 (N_15801,N_14212,N_14805);
xor U15802 (N_15802,N_14585,N_14040);
xor U15803 (N_15803,N_14700,N_14793);
nand U15804 (N_15804,N_14533,N_14749);
or U15805 (N_15805,N_14478,N_14699);
nand U15806 (N_15806,N_14778,N_14015);
or U15807 (N_15807,N_14661,N_14850);
and U15808 (N_15808,N_14342,N_14810);
or U15809 (N_15809,N_14965,N_14719);
nor U15810 (N_15810,N_14217,N_14070);
and U15811 (N_15811,N_14737,N_14343);
nor U15812 (N_15812,N_14609,N_14121);
or U15813 (N_15813,N_14854,N_14679);
or U15814 (N_15814,N_14842,N_14744);
nand U15815 (N_15815,N_14244,N_14255);
nor U15816 (N_15816,N_14886,N_14973);
nor U15817 (N_15817,N_14815,N_14119);
or U15818 (N_15818,N_14222,N_14812);
and U15819 (N_15819,N_14021,N_14498);
nand U15820 (N_15820,N_14066,N_14651);
xor U15821 (N_15821,N_14773,N_14041);
nor U15822 (N_15822,N_14738,N_14450);
and U15823 (N_15823,N_14427,N_14981);
nand U15824 (N_15824,N_14632,N_14415);
nor U15825 (N_15825,N_14308,N_14739);
nor U15826 (N_15826,N_14930,N_14464);
nand U15827 (N_15827,N_14043,N_14144);
xor U15828 (N_15828,N_14239,N_14743);
nand U15829 (N_15829,N_14385,N_14706);
xnor U15830 (N_15830,N_14736,N_14099);
and U15831 (N_15831,N_14341,N_14529);
or U15832 (N_15832,N_14044,N_14762);
xor U15833 (N_15833,N_14895,N_14156);
or U15834 (N_15834,N_14378,N_14420);
nand U15835 (N_15835,N_14903,N_14407);
xor U15836 (N_15836,N_14912,N_14180);
nand U15837 (N_15837,N_14489,N_14837);
or U15838 (N_15838,N_14984,N_14667);
and U15839 (N_15839,N_14074,N_14586);
and U15840 (N_15840,N_14013,N_14870);
nor U15841 (N_15841,N_14034,N_14960);
nor U15842 (N_15842,N_14058,N_14767);
nor U15843 (N_15843,N_14698,N_14559);
or U15844 (N_15844,N_14498,N_14432);
or U15845 (N_15845,N_14637,N_14358);
nor U15846 (N_15846,N_14010,N_14947);
nand U15847 (N_15847,N_14102,N_14700);
nor U15848 (N_15848,N_14004,N_14285);
nand U15849 (N_15849,N_14248,N_14598);
nand U15850 (N_15850,N_14612,N_14876);
or U15851 (N_15851,N_14415,N_14732);
nor U15852 (N_15852,N_14375,N_14721);
and U15853 (N_15853,N_14597,N_14573);
nor U15854 (N_15854,N_14989,N_14096);
or U15855 (N_15855,N_14240,N_14135);
or U15856 (N_15856,N_14049,N_14242);
or U15857 (N_15857,N_14702,N_14346);
and U15858 (N_15858,N_14293,N_14677);
and U15859 (N_15859,N_14167,N_14102);
nor U15860 (N_15860,N_14750,N_14069);
nand U15861 (N_15861,N_14634,N_14899);
xnor U15862 (N_15862,N_14081,N_14765);
xor U15863 (N_15863,N_14544,N_14899);
xnor U15864 (N_15864,N_14294,N_14043);
or U15865 (N_15865,N_14654,N_14263);
and U15866 (N_15866,N_14341,N_14617);
and U15867 (N_15867,N_14717,N_14429);
or U15868 (N_15868,N_14915,N_14328);
and U15869 (N_15869,N_14361,N_14852);
and U15870 (N_15870,N_14738,N_14930);
nor U15871 (N_15871,N_14802,N_14632);
xnor U15872 (N_15872,N_14215,N_14928);
or U15873 (N_15873,N_14433,N_14673);
nand U15874 (N_15874,N_14701,N_14128);
and U15875 (N_15875,N_14886,N_14228);
xor U15876 (N_15876,N_14932,N_14082);
and U15877 (N_15877,N_14417,N_14960);
nor U15878 (N_15878,N_14749,N_14631);
nand U15879 (N_15879,N_14925,N_14258);
or U15880 (N_15880,N_14014,N_14486);
and U15881 (N_15881,N_14990,N_14005);
nor U15882 (N_15882,N_14290,N_14896);
or U15883 (N_15883,N_14934,N_14497);
nor U15884 (N_15884,N_14232,N_14904);
or U15885 (N_15885,N_14024,N_14937);
or U15886 (N_15886,N_14554,N_14742);
or U15887 (N_15887,N_14670,N_14621);
nand U15888 (N_15888,N_14619,N_14219);
or U15889 (N_15889,N_14232,N_14669);
nand U15890 (N_15890,N_14860,N_14026);
nor U15891 (N_15891,N_14137,N_14248);
or U15892 (N_15892,N_14463,N_14529);
and U15893 (N_15893,N_14480,N_14790);
or U15894 (N_15894,N_14665,N_14230);
and U15895 (N_15895,N_14461,N_14995);
and U15896 (N_15896,N_14523,N_14704);
and U15897 (N_15897,N_14486,N_14668);
nor U15898 (N_15898,N_14892,N_14670);
or U15899 (N_15899,N_14138,N_14362);
nand U15900 (N_15900,N_14033,N_14118);
or U15901 (N_15901,N_14245,N_14360);
nand U15902 (N_15902,N_14222,N_14462);
or U15903 (N_15903,N_14331,N_14834);
nor U15904 (N_15904,N_14199,N_14796);
nand U15905 (N_15905,N_14095,N_14212);
xor U15906 (N_15906,N_14878,N_14879);
or U15907 (N_15907,N_14600,N_14380);
nand U15908 (N_15908,N_14408,N_14937);
nor U15909 (N_15909,N_14989,N_14558);
or U15910 (N_15910,N_14174,N_14746);
xor U15911 (N_15911,N_14659,N_14074);
or U15912 (N_15912,N_14704,N_14436);
xnor U15913 (N_15913,N_14735,N_14312);
or U15914 (N_15914,N_14712,N_14923);
and U15915 (N_15915,N_14081,N_14486);
nor U15916 (N_15916,N_14228,N_14832);
and U15917 (N_15917,N_14354,N_14548);
and U15918 (N_15918,N_14014,N_14589);
or U15919 (N_15919,N_14684,N_14379);
nand U15920 (N_15920,N_14120,N_14778);
nand U15921 (N_15921,N_14776,N_14030);
and U15922 (N_15922,N_14851,N_14156);
and U15923 (N_15923,N_14849,N_14091);
nand U15924 (N_15924,N_14888,N_14591);
nor U15925 (N_15925,N_14105,N_14790);
and U15926 (N_15926,N_14762,N_14824);
nand U15927 (N_15927,N_14222,N_14724);
nand U15928 (N_15928,N_14320,N_14163);
or U15929 (N_15929,N_14852,N_14823);
and U15930 (N_15930,N_14562,N_14155);
or U15931 (N_15931,N_14327,N_14846);
nand U15932 (N_15932,N_14704,N_14580);
or U15933 (N_15933,N_14762,N_14947);
nand U15934 (N_15934,N_14711,N_14772);
and U15935 (N_15935,N_14227,N_14796);
nor U15936 (N_15936,N_14805,N_14913);
and U15937 (N_15937,N_14920,N_14837);
xnor U15938 (N_15938,N_14872,N_14278);
xor U15939 (N_15939,N_14479,N_14621);
nor U15940 (N_15940,N_14340,N_14275);
xnor U15941 (N_15941,N_14108,N_14412);
nand U15942 (N_15942,N_14224,N_14839);
or U15943 (N_15943,N_14878,N_14949);
and U15944 (N_15944,N_14211,N_14773);
xnor U15945 (N_15945,N_14846,N_14437);
or U15946 (N_15946,N_14015,N_14026);
xor U15947 (N_15947,N_14253,N_14353);
nand U15948 (N_15948,N_14728,N_14630);
or U15949 (N_15949,N_14856,N_14535);
and U15950 (N_15950,N_14505,N_14106);
and U15951 (N_15951,N_14153,N_14830);
nand U15952 (N_15952,N_14763,N_14523);
and U15953 (N_15953,N_14687,N_14281);
nand U15954 (N_15954,N_14296,N_14610);
or U15955 (N_15955,N_14037,N_14057);
nand U15956 (N_15956,N_14776,N_14726);
nand U15957 (N_15957,N_14609,N_14796);
or U15958 (N_15958,N_14543,N_14853);
nand U15959 (N_15959,N_14653,N_14862);
and U15960 (N_15960,N_14867,N_14808);
and U15961 (N_15961,N_14037,N_14564);
and U15962 (N_15962,N_14566,N_14990);
and U15963 (N_15963,N_14708,N_14862);
or U15964 (N_15964,N_14948,N_14036);
or U15965 (N_15965,N_14050,N_14509);
nand U15966 (N_15966,N_14484,N_14524);
or U15967 (N_15967,N_14365,N_14731);
or U15968 (N_15968,N_14846,N_14588);
or U15969 (N_15969,N_14379,N_14647);
and U15970 (N_15970,N_14433,N_14712);
or U15971 (N_15971,N_14626,N_14516);
or U15972 (N_15972,N_14671,N_14385);
and U15973 (N_15973,N_14233,N_14253);
nand U15974 (N_15974,N_14462,N_14532);
nor U15975 (N_15975,N_14509,N_14164);
xor U15976 (N_15976,N_14717,N_14650);
xnor U15977 (N_15977,N_14546,N_14299);
xnor U15978 (N_15978,N_14746,N_14650);
nand U15979 (N_15979,N_14118,N_14012);
nand U15980 (N_15980,N_14191,N_14478);
and U15981 (N_15981,N_14206,N_14301);
or U15982 (N_15982,N_14650,N_14897);
xnor U15983 (N_15983,N_14881,N_14052);
and U15984 (N_15984,N_14164,N_14128);
nor U15985 (N_15985,N_14047,N_14121);
or U15986 (N_15986,N_14026,N_14479);
and U15987 (N_15987,N_14610,N_14772);
and U15988 (N_15988,N_14575,N_14799);
nor U15989 (N_15989,N_14616,N_14952);
and U15990 (N_15990,N_14676,N_14984);
nand U15991 (N_15991,N_14398,N_14098);
nand U15992 (N_15992,N_14493,N_14466);
and U15993 (N_15993,N_14619,N_14256);
and U15994 (N_15994,N_14847,N_14157);
xnor U15995 (N_15995,N_14758,N_14553);
and U15996 (N_15996,N_14951,N_14318);
or U15997 (N_15997,N_14647,N_14446);
or U15998 (N_15998,N_14749,N_14260);
nand U15999 (N_15999,N_14089,N_14644);
nor U16000 (N_16000,N_15049,N_15722);
nand U16001 (N_16001,N_15747,N_15269);
nor U16002 (N_16002,N_15430,N_15846);
and U16003 (N_16003,N_15466,N_15808);
nor U16004 (N_16004,N_15817,N_15376);
nor U16005 (N_16005,N_15922,N_15210);
nor U16006 (N_16006,N_15490,N_15016);
or U16007 (N_16007,N_15972,N_15708);
nor U16008 (N_16008,N_15677,N_15789);
and U16009 (N_16009,N_15800,N_15758);
nand U16010 (N_16010,N_15050,N_15001);
nor U16011 (N_16011,N_15865,N_15406);
nand U16012 (N_16012,N_15870,N_15869);
and U16013 (N_16013,N_15033,N_15187);
nor U16014 (N_16014,N_15285,N_15811);
xnor U16015 (N_16015,N_15666,N_15636);
nor U16016 (N_16016,N_15436,N_15215);
or U16017 (N_16017,N_15750,N_15769);
or U16018 (N_16018,N_15943,N_15839);
and U16019 (N_16019,N_15516,N_15634);
nand U16020 (N_16020,N_15208,N_15385);
nor U16021 (N_16021,N_15093,N_15759);
nand U16022 (N_16022,N_15075,N_15774);
nand U16023 (N_16023,N_15855,N_15268);
nor U16024 (N_16024,N_15852,N_15900);
and U16025 (N_16025,N_15960,N_15624);
nand U16026 (N_16026,N_15003,N_15421);
and U16027 (N_16027,N_15939,N_15894);
nor U16028 (N_16028,N_15332,N_15567);
or U16029 (N_16029,N_15102,N_15165);
xor U16030 (N_16030,N_15270,N_15927);
or U16031 (N_16031,N_15505,N_15161);
and U16032 (N_16032,N_15889,N_15909);
nand U16033 (N_16033,N_15999,N_15314);
nand U16034 (N_16034,N_15345,N_15105);
or U16035 (N_16035,N_15162,N_15279);
nor U16036 (N_16036,N_15947,N_15657);
nor U16037 (N_16037,N_15382,N_15893);
or U16038 (N_16038,N_15521,N_15916);
or U16039 (N_16039,N_15932,N_15265);
and U16040 (N_16040,N_15837,N_15973);
nor U16041 (N_16041,N_15045,N_15663);
and U16042 (N_16042,N_15310,N_15699);
nand U16043 (N_16043,N_15561,N_15358);
or U16044 (N_16044,N_15252,N_15445);
xor U16045 (N_16045,N_15111,N_15908);
or U16046 (N_16046,N_15712,N_15654);
or U16047 (N_16047,N_15146,N_15531);
nor U16048 (N_16048,N_15099,N_15827);
and U16049 (N_16049,N_15929,N_15040);
and U16050 (N_16050,N_15910,N_15524);
nor U16051 (N_16051,N_15174,N_15984);
or U16052 (N_16052,N_15234,N_15553);
nand U16053 (N_16053,N_15764,N_15849);
and U16054 (N_16054,N_15831,N_15606);
nand U16055 (N_16055,N_15670,N_15071);
or U16056 (N_16056,N_15935,N_15925);
and U16057 (N_16057,N_15621,N_15773);
and U16058 (N_16058,N_15957,N_15956);
xor U16059 (N_16059,N_15125,N_15739);
nor U16060 (N_16060,N_15572,N_15951);
nor U16061 (N_16061,N_15807,N_15189);
nor U16062 (N_16062,N_15583,N_15812);
and U16063 (N_16063,N_15416,N_15588);
or U16064 (N_16064,N_15316,N_15224);
nand U16065 (N_16065,N_15112,N_15244);
nand U16066 (N_16066,N_15848,N_15840);
and U16067 (N_16067,N_15734,N_15410);
or U16068 (N_16068,N_15619,N_15170);
nor U16069 (N_16069,N_15482,N_15440);
or U16070 (N_16070,N_15625,N_15177);
and U16071 (N_16071,N_15976,N_15294);
or U16072 (N_16072,N_15938,N_15336);
nor U16073 (N_16073,N_15199,N_15288);
nor U16074 (N_16074,N_15213,N_15048);
or U16075 (N_16075,N_15184,N_15245);
xnor U16076 (N_16076,N_15204,N_15679);
or U16077 (N_16077,N_15323,N_15547);
and U16078 (N_16078,N_15667,N_15305);
or U16079 (N_16079,N_15608,N_15222);
nor U16080 (N_16080,N_15477,N_15727);
and U16081 (N_16081,N_15228,N_15261);
nand U16082 (N_16082,N_15958,N_15859);
and U16083 (N_16083,N_15079,N_15731);
nor U16084 (N_16084,N_15132,N_15662);
and U16085 (N_16085,N_15744,N_15481);
nand U16086 (N_16086,N_15605,N_15611);
nand U16087 (N_16087,N_15881,N_15297);
or U16088 (N_16088,N_15772,N_15328);
nor U16089 (N_16089,N_15655,N_15687);
and U16090 (N_16090,N_15373,N_15381);
and U16091 (N_16091,N_15114,N_15063);
and U16092 (N_16092,N_15777,N_15710);
xor U16093 (N_16093,N_15429,N_15835);
nor U16094 (N_16094,N_15729,N_15127);
or U16095 (N_16095,N_15562,N_15962);
or U16096 (N_16096,N_15716,N_15415);
nand U16097 (N_16097,N_15923,N_15448);
nand U16098 (N_16098,N_15100,N_15380);
or U16099 (N_16099,N_15020,N_15355);
or U16100 (N_16100,N_15728,N_15009);
nor U16101 (N_16101,N_15286,N_15472);
and U16102 (N_16102,N_15882,N_15838);
and U16103 (N_16103,N_15289,N_15593);
and U16104 (N_16104,N_15604,N_15299);
and U16105 (N_16105,N_15950,N_15640);
nand U16106 (N_16106,N_15124,N_15641);
or U16107 (N_16107,N_15778,N_15023);
xnor U16108 (N_16108,N_15362,N_15390);
nand U16109 (N_16109,N_15128,N_15301);
or U16110 (N_16110,N_15235,N_15700);
or U16111 (N_16111,N_15186,N_15665);
nor U16112 (N_16112,N_15157,N_15696);
or U16113 (N_16113,N_15961,N_15039);
and U16114 (N_16114,N_15786,N_15072);
xor U16115 (N_16115,N_15143,N_15863);
nand U16116 (N_16116,N_15044,N_15232);
or U16117 (N_16117,N_15046,N_15029);
nor U16118 (N_16118,N_15136,N_15303);
nand U16119 (N_16119,N_15431,N_15717);
nand U16120 (N_16120,N_15450,N_15584);
nor U16121 (N_16121,N_15229,N_15497);
or U16122 (N_16122,N_15272,N_15331);
nor U16123 (N_16123,N_15348,N_15338);
nor U16124 (N_16124,N_15196,N_15159);
nor U16125 (N_16125,N_15087,N_15587);
nor U16126 (N_16126,N_15674,N_15578);
or U16127 (N_16127,N_15056,N_15681);
or U16128 (N_16128,N_15220,N_15726);
and U16129 (N_16129,N_15183,N_15080);
xor U16130 (N_16130,N_15954,N_15342);
or U16131 (N_16131,N_15799,N_15260);
nor U16132 (N_16132,N_15979,N_15532);
nor U16133 (N_16133,N_15118,N_15387);
and U16134 (N_16134,N_15590,N_15560);
nor U16135 (N_16135,N_15818,N_15586);
and U16136 (N_16136,N_15070,N_15678);
or U16137 (N_16137,N_15110,N_15325);
and U16138 (N_16138,N_15293,N_15522);
or U16139 (N_16139,N_15083,N_15978);
or U16140 (N_16140,N_15755,N_15902);
and U16141 (N_16141,N_15158,N_15824);
nor U16142 (N_16142,N_15478,N_15825);
nand U16143 (N_16143,N_15403,N_15783);
nor U16144 (N_16144,N_15779,N_15433);
or U16145 (N_16145,N_15366,N_15469);
or U16146 (N_16146,N_15246,N_15513);
xor U16147 (N_16147,N_15703,N_15295);
and U16148 (N_16148,N_15405,N_15646);
or U16149 (N_16149,N_15610,N_15613);
xnor U16150 (N_16150,N_15509,N_15926);
or U16151 (N_16151,N_15462,N_15372);
or U16152 (N_16152,N_15540,N_15695);
nand U16153 (N_16153,N_15074,N_15138);
and U16154 (N_16154,N_15231,N_15378);
nor U16155 (N_16155,N_15496,N_15259);
or U16156 (N_16156,N_15797,N_15256);
nand U16157 (N_16157,N_15137,N_15868);
nand U16158 (N_16158,N_15660,N_15308);
and U16159 (N_16159,N_15313,N_15528);
and U16160 (N_16160,N_15595,N_15903);
nand U16161 (N_16161,N_15659,N_15485);
or U16162 (N_16162,N_15460,N_15077);
nor U16163 (N_16163,N_15644,N_15324);
or U16164 (N_16164,N_15698,N_15991);
nand U16165 (N_16165,N_15113,N_15467);
or U16166 (N_16166,N_15008,N_15475);
or U16167 (N_16167,N_15026,N_15834);
and U16168 (N_16168,N_15267,N_15239);
nor U16169 (N_16169,N_15997,N_15351);
or U16170 (N_16170,N_15617,N_15983);
xnor U16171 (N_16171,N_15171,N_15874);
and U16172 (N_16172,N_15768,N_15092);
nor U16173 (N_16173,N_15694,N_15918);
nand U16174 (N_16174,N_15880,N_15395);
and U16175 (N_16175,N_15898,N_15569);
nor U16176 (N_16176,N_15411,N_15980);
and U16177 (N_16177,N_15761,N_15122);
or U16178 (N_16178,N_15630,N_15451);
nand U16179 (N_16179,N_15539,N_15051);
nor U16180 (N_16180,N_15262,N_15751);
or U16181 (N_16181,N_15438,N_15527);
nor U16182 (N_16182,N_15147,N_15091);
xor U16183 (N_16183,N_15271,N_15027);
or U16184 (N_16184,N_15059,N_15317);
nand U16185 (N_16185,N_15153,N_15781);
nor U16186 (N_16186,N_15274,N_15441);
xnor U16187 (N_16187,N_15223,N_15990);
and U16188 (N_16188,N_15287,N_15830);
and U16189 (N_16189,N_15740,N_15452);
xnor U16190 (N_16190,N_15784,N_15533);
nand U16191 (N_16191,N_15886,N_15725);
or U16192 (N_16192,N_15047,N_15885);
and U16193 (N_16193,N_15707,N_15221);
nor U16194 (N_16194,N_15914,N_15375);
nand U16195 (N_16195,N_15684,N_15018);
nor U16196 (N_16196,N_15814,N_15892);
nor U16197 (N_16197,N_15141,N_15686);
or U16198 (N_16198,N_15276,N_15545);
nor U16199 (N_16199,N_15603,N_15104);
nand U16200 (N_16200,N_15335,N_15340);
nand U16201 (N_16201,N_15393,N_15930);
or U16202 (N_16202,N_15770,N_15484);
and U16203 (N_16203,N_15249,N_15844);
nand U16204 (N_16204,N_15052,N_15815);
nand U16205 (N_16205,N_15804,N_15594);
xor U16206 (N_16206,N_15422,N_15822);
nand U16207 (N_16207,N_15283,N_15017);
or U16208 (N_16208,N_15873,N_15709);
and U16209 (N_16209,N_15803,N_15793);
nand U16210 (N_16210,N_15692,N_15845);
or U16211 (N_16211,N_15273,N_15361);
or U16212 (N_16212,N_15188,N_15088);
nor U16213 (N_16213,N_15302,N_15194);
nor U16214 (N_16214,N_15058,N_15457);
xnor U16215 (N_16215,N_15209,N_15760);
nand U16216 (N_16216,N_15185,N_15697);
nand U16217 (N_16217,N_15119,N_15264);
or U16218 (N_16218,N_15250,N_15298);
and U16219 (N_16219,N_15370,N_15237);
nand U16220 (N_16220,N_15721,N_15327);
and U16221 (N_16221,N_15765,N_15771);
nor U16222 (N_16222,N_15549,N_15629);
nor U16223 (N_16223,N_15247,N_15704);
nor U16224 (N_16224,N_15541,N_15094);
nand U16225 (N_16225,N_15628,N_15488);
and U16226 (N_16226,N_15591,N_15115);
nand U16227 (N_16227,N_15551,N_15981);
nor U16228 (N_16228,N_15995,N_15656);
or U16229 (N_16229,N_15167,N_15581);
and U16230 (N_16230,N_15368,N_15166);
and U16231 (N_16231,N_15756,N_15913);
nand U16232 (N_16232,N_15139,N_15350);
or U16233 (N_16233,N_15622,N_15673);
nor U16234 (N_16234,N_15359,N_15354);
nor U16235 (N_16235,N_15263,N_15015);
nand U16236 (N_16236,N_15790,N_15470);
and U16237 (N_16237,N_15529,N_15501);
nor U16238 (N_16238,N_15919,N_15084);
and U16239 (N_16239,N_15631,N_15471);
and U16240 (N_16240,N_15861,N_15510);
nand U16241 (N_16241,N_15638,N_15206);
xor U16242 (N_16242,N_15862,N_15546);
nand U16243 (N_16243,N_15872,N_15917);
nor U16244 (N_16244,N_15579,N_15465);
or U16245 (N_16245,N_15955,N_15977);
nor U16246 (N_16246,N_15851,N_15520);
or U16247 (N_16247,N_15690,N_15409);
or U16248 (N_16248,N_15347,N_15915);
or U16249 (N_16249,N_15735,N_15805);
or U16250 (N_16250,N_15671,N_15306);
nand U16251 (N_16251,N_15435,N_15555);
nor U16252 (N_16252,N_15312,N_15321);
or U16253 (N_16253,N_15905,N_15201);
or U16254 (N_16254,N_15689,N_15538);
nor U16255 (N_16255,N_15367,N_15198);
xnor U16256 (N_16256,N_15899,N_15589);
nor U16257 (N_16257,N_15688,N_15389);
or U16258 (N_16258,N_15019,N_15633);
and U16259 (N_16259,N_15650,N_15364);
or U16260 (N_16260,N_15349,N_15180);
nand U16261 (N_16261,N_15398,N_15211);
and U16262 (N_16262,N_15878,N_15024);
nor U16263 (N_16263,N_15453,N_15014);
and U16264 (N_16264,N_15255,N_15004);
and U16265 (N_16265,N_15836,N_15192);
xor U16266 (N_16266,N_15733,N_15599);
or U16267 (N_16267,N_15007,N_15498);
or U16268 (N_16268,N_15178,N_15934);
nor U16269 (N_16269,N_15330,N_15282);
or U16270 (N_16270,N_15963,N_15858);
and U16271 (N_16271,N_15195,N_15341);
nand U16272 (N_16272,N_15000,N_15277);
or U16273 (N_16273,N_15802,N_15653);
or U16274 (N_16274,N_15495,N_15661);
xnor U16275 (N_16275,N_15503,N_15748);
nand U16276 (N_16276,N_15427,N_15944);
nor U16277 (N_16277,N_15344,N_15940);
nand U16278 (N_16278,N_15548,N_15720);
nor U16279 (N_16279,N_15291,N_15512);
and U16280 (N_16280,N_15596,N_15006);
or U16281 (N_16281,N_15565,N_15682);
or U16282 (N_16282,N_15369,N_15573);
xor U16283 (N_16283,N_15907,N_15145);
nand U16284 (N_16284,N_15447,N_15618);
nor U16285 (N_16285,N_15996,N_15197);
or U16286 (N_16286,N_15754,N_15401);
nand U16287 (N_16287,N_15975,N_15702);
nand U16288 (N_16288,N_15966,N_15993);
or U16289 (N_16289,N_15504,N_15676);
nand U16290 (N_16290,N_15906,N_15871);
or U16291 (N_16291,N_15135,N_15096);
nand U16292 (N_16292,N_15536,N_15499);
or U16293 (N_16293,N_15134,N_15508);
and U16294 (N_16294,N_15928,N_15753);
and U16295 (N_16295,N_15154,N_15637);
nor U16296 (N_16296,N_15468,N_15737);
nand U16297 (N_16297,N_15648,N_15238);
xnor U16298 (N_16298,N_15626,N_15506);
and U16299 (N_16299,N_15685,N_15543);
and U16300 (N_16300,N_15842,N_15920);
xnor U16301 (N_16301,N_15123,N_15106);
xnor U16302 (N_16302,N_15570,N_15517);
or U16303 (N_16303,N_15988,N_15149);
or U16304 (N_16304,N_15173,N_15025);
xor U16305 (N_16305,N_15742,N_15404);
or U16306 (N_16306,N_15876,N_15021);
or U16307 (N_16307,N_15172,N_15217);
nor U16308 (N_16308,N_15097,N_15998);
nand U16309 (N_16309,N_15967,N_15428);
and U16310 (N_16310,N_15275,N_15319);
nor U16311 (N_16311,N_15714,N_15826);
and U16312 (N_16312,N_15182,N_15597);
nor U16313 (N_16313,N_15365,N_15476);
and U16314 (N_16314,N_15557,N_15888);
nor U16315 (N_16315,N_15525,N_15683);
nor U16316 (N_16316,N_15492,N_15607);
nor U16317 (N_16317,N_15311,N_15121);
or U16318 (N_16318,N_15518,N_15795);
and U16319 (N_16319,N_15642,N_15566);
nand U16320 (N_16320,N_15575,N_15623);
and U16321 (N_16321,N_15813,N_15664);
and U16322 (N_16322,N_15054,N_15732);
and U16323 (N_16323,N_15242,N_15062);
nor U16324 (N_16324,N_15064,N_15425);
nor U16325 (N_16325,N_15592,N_15461);
or U16326 (N_16326,N_15443,N_15841);
nor U16327 (N_16327,N_15164,N_15969);
or U16328 (N_16328,N_15864,N_15821);
or U16329 (N_16329,N_15843,N_15374);
nand U16330 (N_16330,N_15363,N_15819);
nor U16331 (N_16331,N_15635,N_15502);
and U16332 (N_16332,N_15266,N_15647);
xor U16333 (N_16333,N_15081,N_15952);
nand U16334 (N_16334,N_15432,N_15258);
and U16335 (N_16335,N_15152,N_15455);
nand U16336 (N_16336,N_15931,N_15985);
or U16337 (N_16337,N_15176,N_15791);
nand U16338 (N_16338,N_15109,N_15407);
xnor U16339 (N_16339,N_15437,N_15911);
or U16340 (N_16340,N_15060,N_15131);
xnor U16341 (N_16341,N_15002,N_15680);
nand U16342 (N_16342,N_15828,N_15775);
and U16343 (N_16343,N_15743,N_15190);
nand U16344 (N_16344,N_15776,N_15388);
and U16345 (N_16345,N_15941,N_15163);
nand U16346 (N_16346,N_15544,N_15877);
and U16347 (N_16347,N_15419,N_15600);
nor U16348 (N_16348,N_15423,N_15946);
or U16349 (N_16349,N_15823,N_15028);
nor U16350 (N_16350,N_15140,N_15820);
nand U16351 (N_16351,N_15658,N_15537);
or U16352 (N_16352,N_15307,N_15396);
nor U16353 (N_16353,N_15493,N_15491);
nand U16354 (N_16354,N_15417,N_15292);
and U16355 (N_16355,N_15300,N_15010);
nand U16356 (N_16356,N_15090,N_15126);
or U16357 (N_16357,N_15459,N_15191);
or U16358 (N_16358,N_15035,N_15031);
nor U16359 (N_16359,N_15895,N_15489);
nor U16360 (N_16360,N_15103,N_15169);
and U16361 (N_16361,N_15724,N_15936);
nand U16362 (N_16362,N_15212,N_15523);
and U16363 (N_16363,N_15318,N_15794);
or U16364 (N_16364,N_15434,N_15278);
or U16365 (N_16365,N_15896,N_15563);
nand U16366 (N_16366,N_15480,N_15379);
nor U16367 (N_16367,N_15711,N_15078);
xnor U16368 (N_16368,N_15280,N_15701);
or U16369 (N_16369,N_15486,N_15965);
nor U16370 (N_16370,N_15494,N_15151);
and U16371 (N_16371,N_15352,N_15526);
nand U16372 (N_16372,N_15326,N_15968);
xnor U16373 (N_16373,N_15571,N_15066);
nand U16374 (N_16374,N_15749,N_15970);
nand U16375 (N_16375,N_15782,N_15402);
and U16376 (N_16376,N_15067,N_15652);
and U16377 (N_16377,N_15408,N_15251);
nor U16378 (N_16378,N_15043,N_15377);
xor U16379 (N_16379,N_15816,N_15713);
and U16380 (N_16380,N_15582,N_15474);
nor U16381 (N_16381,N_15809,N_15243);
or U16382 (N_16382,N_15576,N_15762);
nand U16383 (N_16383,N_15038,N_15933);
nor U16384 (N_16384,N_15854,N_15296);
or U16385 (N_16385,N_15086,N_15346);
and U16386 (N_16386,N_15986,N_15989);
or U16387 (N_16387,N_15011,N_15598);
nor U16388 (N_16388,N_15449,N_15949);
or U16389 (N_16389,N_15334,N_15337);
or U16390 (N_16390,N_15444,N_15420);
and U16391 (N_16391,N_15400,N_15357);
nor U16392 (N_16392,N_15577,N_15248);
nor U16393 (N_16393,N_15884,N_15953);
nand U16394 (N_16394,N_15257,N_15639);
nand U16395 (N_16395,N_15627,N_15620);
or U16396 (N_16396,N_15609,N_15005);
nand U16397 (N_16397,N_15130,N_15036);
xnor U16398 (N_16398,N_15937,N_15384);
and U16399 (N_16399,N_15193,N_15095);
or U16400 (N_16400,N_15875,N_15612);
xnor U16401 (N_16401,N_15254,N_15550);
nand U16402 (N_16402,N_15030,N_15101);
nand U16403 (N_16403,N_15343,N_15200);
nor U16404 (N_16404,N_15168,N_15643);
nand U16405 (N_16405,N_15181,N_15847);
and U16406 (N_16406,N_15867,N_15391);
and U16407 (N_16407,N_15442,N_15107);
nor U16408 (N_16408,N_15718,N_15290);
nor U16409 (N_16409,N_15780,N_15022);
nor U16410 (N_16410,N_15788,N_15240);
and U16411 (N_16411,N_15833,N_15487);
nor U16412 (N_16412,N_15155,N_15360);
xnor U16413 (N_16413,N_15315,N_15715);
or U16414 (N_16414,N_15601,N_15034);
xor U16415 (N_16415,N_15745,N_15089);
or U16416 (N_16416,N_15418,N_15339);
or U16417 (N_16417,N_15120,N_15329);
nand U16418 (N_16418,N_15236,N_15992);
and U16419 (N_16419,N_15424,N_15853);
nor U16420 (N_16420,N_15116,N_15383);
or U16421 (N_16421,N_15971,N_15479);
nor U16422 (N_16422,N_15558,N_15669);
nand U16423 (N_16423,N_15065,N_15399);
and U16424 (N_16424,N_15281,N_15556);
and U16425 (N_16425,N_15156,N_15012);
or U16426 (N_16426,N_15866,N_15741);
nor U16427 (N_16427,N_15574,N_15736);
nor U16428 (N_16428,N_15233,N_15668);
nor U16429 (N_16429,N_15304,N_15706);
or U16430 (N_16430,N_15829,N_15767);
or U16431 (N_16431,N_15483,N_15397);
xor U16432 (N_16432,N_15810,N_15041);
or U16433 (N_16433,N_15160,N_15564);
nand U16434 (N_16434,N_15032,N_15061);
and U16435 (N_16435,N_15850,N_15055);
and U16436 (N_16436,N_15148,N_15832);
nand U16437 (N_16437,N_15068,N_15921);
nor U16438 (N_16438,N_15085,N_15142);
or U16439 (N_16439,N_15353,N_15890);
nand U16440 (N_16440,N_15942,N_15394);
nor U16441 (N_16441,N_15133,N_15253);
xor U16442 (N_16442,N_15796,N_15798);
or U16443 (N_16443,N_15456,N_15801);
or U16444 (N_16444,N_15860,N_15511);
nor U16445 (N_16445,N_15230,N_15446);
nor U16446 (N_16446,N_15904,N_15585);
nor U16447 (N_16447,N_15057,N_15987);
and U16448 (N_16448,N_15473,N_15412);
and U16449 (N_16449,N_15982,N_15507);
nand U16450 (N_16450,N_15042,N_15924);
nand U16451 (N_16451,N_15719,N_15787);
nor U16452 (N_16452,N_15530,N_15333);
and U16453 (N_16453,N_15632,N_15568);
or U16454 (N_16454,N_15069,N_15535);
nand U16455 (N_16455,N_15226,N_15948);
xor U16456 (N_16456,N_15738,N_15757);
nor U16457 (N_16457,N_15693,N_15413);
and U16458 (N_16458,N_15225,N_15150);
and U16459 (N_16459,N_15013,N_15454);
and U16460 (N_16460,N_15883,N_15672);
and U16461 (N_16461,N_15108,N_15901);
and U16462 (N_16462,N_15897,N_15227);
nor U16463 (N_16463,N_15356,N_15144);
nand U16464 (N_16464,N_15098,N_15205);
xnor U16465 (N_16465,N_15320,N_15322);
xnor U16466 (N_16466,N_15792,N_15053);
nand U16467 (N_16467,N_15284,N_15414);
and U16468 (N_16468,N_15766,N_15887);
and U16469 (N_16469,N_15309,N_15763);
xnor U16470 (N_16470,N_15891,N_15559);
or U16471 (N_16471,N_15974,N_15439);
nand U16472 (N_16472,N_15785,N_15426);
or U16473 (N_16473,N_15806,N_15614);
nor U16474 (N_16474,N_15076,N_15386);
nor U16475 (N_16475,N_15534,N_15514);
nand U16476 (N_16476,N_15912,N_15515);
nand U16477 (N_16477,N_15202,N_15175);
xnor U16478 (N_16478,N_15037,N_15856);
or U16479 (N_16479,N_15705,N_15241);
nand U16480 (N_16480,N_15500,N_15464);
or U16481 (N_16481,N_15082,N_15645);
nand U16482 (N_16482,N_15675,N_15879);
and U16483 (N_16483,N_15723,N_15746);
or U16484 (N_16484,N_15214,N_15216);
nor U16485 (N_16485,N_15179,N_15554);
and U16486 (N_16486,N_15519,N_15651);
and U16487 (N_16487,N_15371,N_15219);
or U16488 (N_16488,N_15542,N_15392);
nand U16489 (N_16489,N_15463,N_15602);
nand U16490 (N_16490,N_15203,N_15117);
or U16491 (N_16491,N_15580,N_15616);
or U16492 (N_16492,N_15964,N_15959);
xor U16493 (N_16493,N_15730,N_15218);
and U16494 (N_16494,N_15691,N_15857);
and U16495 (N_16495,N_15207,N_15073);
and U16496 (N_16496,N_15129,N_15615);
and U16497 (N_16497,N_15552,N_15752);
nand U16498 (N_16498,N_15458,N_15994);
nor U16499 (N_16499,N_15945,N_15649);
nand U16500 (N_16500,N_15775,N_15767);
nand U16501 (N_16501,N_15878,N_15258);
or U16502 (N_16502,N_15393,N_15117);
and U16503 (N_16503,N_15294,N_15149);
nor U16504 (N_16504,N_15650,N_15943);
nand U16505 (N_16505,N_15519,N_15493);
or U16506 (N_16506,N_15931,N_15023);
nand U16507 (N_16507,N_15767,N_15994);
nand U16508 (N_16508,N_15377,N_15148);
and U16509 (N_16509,N_15890,N_15100);
nor U16510 (N_16510,N_15419,N_15058);
xnor U16511 (N_16511,N_15572,N_15428);
and U16512 (N_16512,N_15408,N_15110);
or U16513 (N_16513,N_15621,N_15490);
and U16514 (N_16514,N_15993,N_15095);
or U16515 (N_16515,N_15782,N_15611);
and U16516 (N_16516,N_15994,N_15581);
and U16517 (N_16517,N_15794,N_15346);
and U16518 (N_16518,N_15327,N_15578);
nand U16519 (N_16519,N_15170,N_15425);
or U16520 (N_16520,N_15570,N_15373);
or U16521 (N_16521,N_15661,N_15665);
nand U16522 (N_16522,N_15344,N_15960);
nand U16523 (N_16523,N_15380,N_15326);
or U16524 (N_16524,N_15929,N_15099);
and U16525 (N_16525,N_15935,N_15649);
nand U16526 (N_16526,N_15301,N_15306);
or U16527 (N_16527,N_15890,N_15601);
nand U16528 (N_16528,N_15110,N_15375);
or U16529 (N_16529,N_15652,N_15730);
nor U16530 (N_16530,N_15710,N_15416);
xor U16531 (N_16531,N_15187,N_15997);
nand U16532 (N_16532,N_15565,N_15780);
or U16533 (N_16533,N_15962,N_15953);
nor U16534 (N_16534,N_15370,N_15934);
nor U16535 (N_16535,N_15899,N_15176);
nand U16536 (N_16536,N_15255,N_15644);
or U16537 (N_16537,N_15366,N_15089);
nor U16538 (N_16538,N_15521,N_15586);
nor U16539 (N_16539,N_15075,N_15101);
or U16540 (N_16540,N_15682,N_15478);
and U16541 (N_16541,N_15514,N_15500);
or U16542 (N_16542,N_15311,N_15564);
and U16543 (N_16543,N_15253,N_15486);
nand U16544 (N_16544,N_15947,N_15876);
xnor U16545 (N_16545,N_15141,N_15732);
nand U16546 (N_16546,N_15436,N_15890);
and U16547 (N_16547,N_15968,N_15800);
and U16548 (N_16548,N_15238,N_15603);
or U16549 (N_16549,N_15904,N_15320);
and U16550 (N_16550,N_15918,N_15258);
xor U16551 (N_16551,N_15420,N_15402);
or U16552 (N_16552,N_15381,N_15209);
nor U16553 (N_16553,N_15453,N_15141);
xor U16554 (N_16554,N_15442,N_15877);
nor U16555 (N_16555,N_15859,N_15661);
nor U16556 (N_16556,N_15530,N_15997);
or U16557 (N_16557,N_15854,N_15398);
or U16558 (N_16558,N_15089,N_15298);
nand U16559 (N_16559,N_15801,N_15433);
nand U16560 (N_16560,N_15026,N_15919);
nor U16561 (N_16561,N_15976,N_15712);
xnor U16562 (N_16562,N_15693,N_15485);
or U16563 (N_16563,N_15696,N_15768);
and U16564 (N_16564,N_15731,N_15104);
xor U16565 (N_16565,N_15432,N_15674);
nor U16566 (N_16566,N_15966,N_15850);
nand U16567 (N_16567,N_15081,N_15492);
and U16568 (N_16568,N_15719,N_15276);
nand U16569 (N_16569,N_15735,N_15267);
and U16570 (N_16570,N_15631,N_15890);
and U16571 (N_16571,N_15748,N_15559);
and U16572 (N_16572,N_15269,N_15563);
or U16573 (N_16573,N_15990,N_15191);
nand U16574 (N_16574,N_15993,N_15032);
and U16575 (N_16575,N_15462,N_15212);
or U16576 (N_16576,N_15154,N_15088);
and U16577 (N_16577,N_15689,N_15679);
and U16578 (N_16578,N_15933,N_15793);
nor U16579 (N_16579,N_15759,N_15142);
nor U16580 (N_16580,N_15669,N_15363);
and U16581 (N_16581,N_15048,N_15025);
nor U16582 (N_16582,N_15955,N_15509);
nand U16583 (N_16583,N_15785,N_15371);
nor U16584 (N_16584,N_15269,N_15567);
and U16585 (N_16585,N_15457,N_15356);
nand U16586 (N_16586,N_15701,N_15198);
or U16587 (N_16587,N_15877,N_15995);
nand U16588 (N_16588,N_15475,N_15685);
nand U16589 (N_16589,N_15878,N_15915);
nor U16590 (N_16590,N_15494,N_15447);
nand U16591 (N_16591,N_15957,N_15543);
nand U16592 (N_16592,N_15641,N_15063);
or U16593 (N_16593,N_15511,N_15289);
and U16594 (N_16594,N_15719,N_15495);
or U16595 (N_16595,N_15089,N_15923);
or U16596 (N_16596,N_15747,N_15367);
nor U16597 (N_16597,N_15502,N_15557);
nor U16598 (N_16598,N_15274,N_15331);
nor U16599 (N_16599,N_15635,N_15746);
nand U16600 (N_16600,N_15165,N_15849);
nor U16601 (N_16601,N_15464,N_15082);
nor U16602 (N_16602,N_15689,N_15246);
or U16603 (N_16603,N_15969,N_15422);
or U16604 (N_16604,N_15741,N_15196);
or U16605 (N_16605,N_15814,N_15771);
or U16606 (N_16606,N_15390,N_15429);
nand U16607 (N_16607,N_15013,N_15816);
and U16608 (N_16608,N_15136,N_15122);
xor U16609 (N_16609,N_15357,N_15313);
and U16610 (N_16610,N_15762,N_15891);
and U16611 (N_16611,N_15511,N_15830);
or U16612 (N_16612,N_15782,N_15491);
or U16613 (N_16613,N_15922,N_15027);
nand U16614 (N_16614,N_15214,N_15236);
and U16615 (N_16615,N_15303,N_15167);
or U16616 (N_16616,N_15735,N_15965);
or U16617 (N_16617,N_15449,N_15641);
or U16618 (N_16618,N_15532,N_15023);
xnor U16619 (N_16619,N_15563,N_15676);
or U16620 (N_16620,N_15041,N_15697);
or U16621 (N_16621,N_15065,N_15374);
nand U16622 (N_16622,N_15690,N_15858);
nand U16623 (N_16623,N_15581,N_15722);
nor U16624 (N_16624,N_15982,N_15313);
nand U16625 (N_16625,N_15179,N_15770);
nand U16626 (N_16626,N_15588,N_15687);
or U16627 (N_16627,N_15316,N_15389);
or U16628 (N_16628,N_15134,N_15797);
or U16629 (N_16629,N_15223,N_15616);
nor U16630 (N_16630,N_15589,N_15525);
or U16631 (N_16631,N_15073,N_15405);
or U16632 (N_16632,N_15053,N_15611);
or U16633 (N_16633,N_15609,N_15359);
nand U16634 (N_16634,N_15569,N_15695);
and U16635 (N_16635,N_15462,N_15338);
or U16636 (N_16636,N_15380,N_15881);
and U16637 (N_16637,N_15226,N_15233);
and U16638 (N_16638,N_15837,N_15442);
nor U16639 (N_16639,N_15384,N_15443);
or U16640 (N_16640,N_15800,N_15557);
nor U16641 (N_16641,N_15635,N_15260);
or U16642 (N_16642,N_15698,N_15013);
or U16643 (N_16643,N_15021,N_15447);
xnor U16644 (N_16644,N_15252,N_15658);
nand U16645 (N_16645,N_15379,N_15569);
nor U16646 (N_16646,N_15274,N_15801);
or U16647 (N_16647,N_15098,N_15767);
nand U16648 (N_16648,N_15118,N_15265);
nor U16649 (N_16649,N_15158,N_15568);
nand U16650 (N_16650,N_15725,N_15126);
and U16651 (N_16651,N_15935,N_15170);
nand U16652 (N_16652,N_15949,N_15122);
nor U16653 (N_16653,N_15615,N_15831);
nand U16654 (N_16654,N_15465,N_15681);
or U16655 (N_16655,N_15437,N_15567);
nor U16656 (N_16656,N_15666,N_15176);
or U16657 (N_16657,N_15167,N_15059);
or U16658 (N_16658,N_15306,N_15153);
xor U16659 (N_16659,N_15918,N_15508);
or U16660 (N_16660,N_15423,N_15122);
nand U16661 (N_16661,N_15392,N_15762);
nand U16662 (N_16662,N_15945,N_15127);
or U16663 (N_16663,N_15963,N_15242);
nand U16664 (N_16664,N_15713,N_15546);
nor U16665 (N_16665,N_15244,N_15649);
and U16666 (N_16666,N_15692,N_15485);
and U16667 (N_16667,N_15396,N_15949);
nand U16668 (N_16668,N_15941,N_15705);
or U16669 (N_16669,N_15362,N_15372);
nor U16670 (N_16670,N_15703,N_15241);
or U16671 (N_16671,N_15412,N_15071);
or U16672 (N_16672,N_15753,N_15123);
nand U16673 (N_16673,N_15538,N_15365);
and U16674 (N_16674,N_15679,N_15134);
or U16675 (N_16675,N_15272,N_15723);
nor U16676 (N_16676,N_15648,N_15119);
or U16677 (N_16677,N_15429,N_15604);
or U16678 (N_16678,N_15606,N_15531);
xor U16679 (N_16679,N_15576,N_15983);
nand U16680 (N_16680,N_15551,N_15832);
or U16681 (N_16681,N_15196,N_15671);
xor U16682 (N_16682,N_15159,N_15219);
nand U16683 (N_16683,N_15214,N_15333);
xnor U16684 (N_16684,N_15468,N_15878);
or U16685 (N_16685,N_15381,N_15071);
and U16686 (N_16686,N_15112,N_15387);
nor U16687 (N_16687,N_15524,N_15891);
nor U16688 (N_16688,N_15036,N_15978);
nor U16689 (N_16689,N_15234,N_15517);
nor U16690 (N_16690,N_15144,N_15659);
and U16691 (N_16691,N_15690,N_15681);
nor U16692 (N_16692,N_15478,N_15519);
nor U16693 (N_16693,N_15753,N_15995);
xnor U16694 (N_16694,N_15686,N_15317);
and U16695 (N_16695,N_15282,N_15517);
and U16696 (N_16696,N_15861,N_15316);
nor U16697 (N_16697,N_15719,N_15875);
nand U16698 (N_16698,N_15084,N_15350);
or U16699 (N_16699,N_15756,N_15946);
nand U16700 (N_16700,N_15969,N_15281);
nand U16701 (N_16701,N_15799,N_15859);
or U16702 (N_16702,N_15285,N_15542);
or U16703 (N_16703,N_15470,N_15688);
or U16704 (N_16704,N_15649,N_15977);
and U16705 (N_16705,N_15052,N_15782);
nand U16706 (N_16706,N_15088,N_15142);
and U16707 (N_16707,N_15071,N_15151);
nor U16708 (N_16708,N_15920,N_15081);
or U16709 (N_16709,N_15111,N_15866);
nand U16710 (N_16710,N_15219,N_15199);
nor U16711 (N_16711,N_15331,N_15714);
xor U16712 (N_16712,N_15232,N_15848);
nor U16713 (N_16713,N_15006,N_15513);
nor U16714 (N_16714,N_15079,N_15865);
or U16715 (N_16715,N_15121,N_15869);
nor U16716 (N_16716,N_15711,N_15135);
and U16717 (N_16717,N_15383,N_15821);
and U16718 (N_16718,N_15205,N_15366);
nor U16719 (N_16719,N_15106,N_15286);
or U16720 (N_16720,N_15390,N_15183);
nor U16721 (N_16721,N_15513,N_15387);
and U16722 (N_16722,N_15399,N_15606);
or U16723 (N_16723,N_15796,N_15986);
or U16724 (N_16724,N_15435,N_15595);
xnor U16725 (N_16725,N_15640,N_15645);
nand U16726 (N_16726,N_15464,N_15180);
and U16727 (N_16727,N_15101,N_15692);
nor U16728 (N_16728,N_15382,N_15093);
nand U16729 (N_16729,N_15244,N_15473);
nand U16730 (N_16730,N_15112,N_15596);
and U16731 (N_16731,N_15068,N_15837);
or U16732 (N_16732,N_15848,N_15099);
nand U16733 (N_16733,N_15538,N_15634);
nor U16734 (N_16734,N_15635,N_15399);
nand U16735 (N_16735,N_15992,N_15770);
or U16736 (N_16736,N_15437,N_15703);
nor U16737 (N_16737,N_15811,N_15678);
and U16738 (N_16738,N_15715,N_15187);
and U16739 (N_16739,N_15297,N_15788);
nand U16740 (N_16740,N_15391,N_15961);
nor U16741 (N_16741,N_15316,N_15410);
nor U16742 (N_16742,N_15563,N_15636);
nor U16743 (N_16743,N_15402,N_15248);
xor U16744 (N_16744,N_15754,N_15866);
and U16745 (N_16745,N_15371,N_15035);
or U16746 (N_16746,N_15894,N_15452);
and U16747 (N_16747,N_15761,N_15208);
and U16748 (N_16748,N_15747,N_15439);
xnor U16749 (N_16749,N_15820,N_15826);
and U16750 (N_16750,N_15980,N_15198);
nor U16751 (N_16751,N_15747,N_15952);
nand U16752 (N_16752,N_15028,N_15626);
xnor U16753 (N_16753,N_15989,N_15951);
or U16754 (N_16754,N_15178,N_15278);
nand U16755 (N_16755,N_15827,N_15649);
or U16756 (N_16756,N_15696,N_15746);
nor U16757 (N_16757,N_15246,N_15023);
nor U16758 (N_16758,N_15947,N_15357);
nand U16759 (N_16759,N_15342,N_15240);
or U16760 (N_16760,N_15160,N_15830);
nand U16761 (N_16761,N_15282,N_15116);
xnor U16762 (N_16762,N_15864,N_15724);
and U16763 (N_16763,N_15684,N_15454);
or U16764 (N_16764,N_15114,N_15694);
nand U16765 (N_16765,N_15849,N_15889);
nand U16766 (N_16766,N_15442,N_15242);
or U16767 (N_16767,N_15019,N_15067);
or U16768 (N_16768,N_15655,N_15429);
xor U16769 (N_16769,N_15461,N_15872);
nand U16770 (N_16770,N_15148,N_15851);
and U16771 (N_16771,N_15172,N_15269);
nor U16772 (N_16772,N_15163,N_15802);
nand U16773 (N_16773,N_15871,N_15352);
nand U16774 (N_16774,N_15491,N_15264);
nand U16775 (N_16775,N_15867,N_15854);
nand U16776 (N_16776,N_15992,N_15249);
nor U16777 (N_16777,N_15110,N_15122);
or U16778 (N_16778,N_15664,N_15638);
nand U16779 (N_16779,N_15404,N_15175);
nand U16780 (N_16780,N_15130,N_15615);
nand U16781 (N_16781,N_15575,N_15336);
or U16782 (N_16782,N_15332,N_15487);
xor U16783 (N_16783,N_15079,N_15228);
nor U16784 (N_16784,N_15368,N_15826);
nor U16785 (N_16785,N_15854,N_15761);
and U16786 (N_16786,N_15074,N_15285);
and U16787 (N_16787,N_15714,N_15822);
or U16788 (N_16788,N_15376,N_15836);
nor U16789 (N_16789,N_15726,N_15184);
xnor U16790 (N_16790,N_15674,N_15719);
and U16791 (N_16791,N_15399,N_15128);
nor U16792 (N_16792,N_15285,N_15569);
nor U16793 (N_16793,N_15033,N_15919);
nor U16794 (N_16794,N_15758,N_15177);
nand U16795 (N_16795,N_15954,N_15606);
and U16796 (N_16796,N_15998,N_15813);
xnor U16797 (N_16797,N_15680,N_15338);
and U16798 (N_16798,N_15218,N_15921);
nand U16799 (N_16799,N_15777,N_15962);
xor U16800 (N_16800,N_15700,N_15198);
and U16801 (N_16801,N_15636,N_15373);
nor U16802 (N_16802,N_15401,N_15940);
nor U16803 (N_16803,N_15338,N_15790);
or U16804 (N_16804,N_15748,N_15441);
nor U16805 (N_16805,N_15539,N_15684);
nor U16806 (N_16806,N_15555,N_15673);
and U16807 (N_16807,N_15056,N_15662);
and U16808 (N_16808,N_15135,N_15886);
or U16809 (N_16809,N_15090,N_15834);
xnor U16810 (N_16810,N_15711,N_15770);
and U16811 (N_16811,N_15814,N_15185);
and U16812 (N_16812,N_15677,N_15587);
and U16813 (N_16813,N_15650,N_15790);
or U16814 (N_16814,N_15309,N_15157);
and U16815 (N_16815,N_15256,N_15296);
or U16816 (N_16816,N_15110,N_15872);
or U16817 (N_16817,N_15488,N_15507);
nand U16818 (N_16818,N_15130,N_15760);
xor U16819 (N_16819,N_15670,N_15635);
and U16820 (N_16820,N_15996,N_15859);
or U16821 (N_16821,N_15981,N_15328);
or U16822 (N_16822,N_15978,N_15599);
nor U16823 (N_16823,N_15118,N_15025);
and U16824 (N_16824,N_15549,N_15396);
and U16825 (N_16825,N_15269,N_15374);
xor U16826 (N_16826,N_15836,N_15255);
and U16827 (N_16827,N_15244,N_15715);
and U16828 (N_16828,N_15932,N_15054);
and U16829 (N_16829,N_15637,N_15236);
nand U16830 (N_16830,N_15351,N_15084);
nand U16831 (N_16831,N_15473,N_15196);
nand U16832 (N_16832,N_15710,N_15177);
nor U16833 (N_16833,N_15758,N_15536);
xor U16834 (N_16834,N_15413,N_15744);
nor U16835 (N_16835,N_15862,N_15172);
and U16836 (N_16836,N_15193,N_15931);
nand U16837 (N_16837,N_15432,N_15554);
or U16838 (N_16838,N_15100,N_15085);
and U16839 (N_16839,N_15499,N_15314);
or U16840 (N_16840,N_15082,N_15692);
or U16841 (N_16841,N_15528,N_15555);
and U16842 (N_16842,N_15600,N_15815);
xnor U16843 (N_16843,N_15571,N_15291);
or U16844 (N_16844,N_15552,N_15594);
xor U16845 (N_16845,N_15694,N_15529);
and U16846 (N_16846,N_15480,N_15887);
xnor U16847 (N_16847,N_15767,N_15745);
and U16848 (N_16848,N_15851,N_15505);
and U16849 (N_16849,N_15054,N_15931);
nor U16850 (N_16850,N_15796,N_15709);
xnor U16851 (N_16851,N_15157,N_15457);
nor U16852 (N_16852,N_15911,N_15789);
nand U16853 (N_16853,N_15596,N_15118);
xor U16854 (N_16854,N_15545,N_15912);
and U16855 (N_16855,N_15285,N_15237);
and U16856 (N_16856,N_15466,N_15410);
nand U16857 (N_16857,N_15830,N_15482);
nor U16858 (N_16858,N_15804,N_15236);
nand U16859 (N_16859,N_15722,N_15215);
or U16860 (N_16860,N_15378,N_15069);
or U16861 (N_16861,N_15843,N_15671);
nor U16862 (N_16862,N_15869,N_15558);
and U16863 (N_16863,N_15994,N_15812);
or U16864 (N_16864,N_15449,N_15621);
or U16865 (N_16865,N_15318,N_15012);
nor U16866 (N_16866,N_15105,N_15125);
xor U16867 (N_16867,N_15219,N_15618);
and U16868 (N_16868,N_15491,N_15611);
nor U16869 (N_16869,N_15391,N_15460);
xor U16870 (N_16870,N_15365,N_15926);
nand U16871 (N_16871,N_15100,N_15439);
and U16872 (N_16872,N_15656,N_15000);
and U16873 (N_16873,N_15826,N_15262);
and U16874 (N_16874,N_15757,N_15770);
or U16875 (N_16875,N_15356,N_15530);
or U16876 (N_16876,N_15536,N_15504);
or U16877 (N_16877,N_15488,N_15340);
xnor U16878 (N_16878,N_15489,N_15421);
or U16879 (N_16879,N_15775,N_15633);
nor U16880 (N_16880,N_15107,N_15603);
nor U16881 (N_16881,N_15622,N_15230);
and U16882 (N_16882,N_15510,N_15713);
or U16883 (N_16883,N_15402,N_15176);
nor U16884 (N_16884,N_15030,N_15276);
nand U16885 (N_16885,N_15691,N_15277);
and U16886 (N_16886,N_15104,N_15660);
and U16887 (N_16887,N_15688,N_15249);
or U16888 (N_16888,N_15331,N_15693);
and U16889 (N_16889,N_15552,N_15093);
nor U16890 (N_16890,N_15630,N_15992);
and U16891 (N_16891,N_15993,N_15026);
nor U16892 (N_16892,N_15111,N_15713);
or U16893 (N_16893,N_15955,N_15370);
and U16894 (N_16894,N_15627,N_15306);
xnor U16895 (N_16895,N_15507,N_15472);
and U16896 (N_16896,N_15305,N_15860);
nor U16897 (N_16897,N_15946,N_15471);
nand U16898 (N_16898,N_15452,N_15230);
xnor U16899 (N_16899,N_15155,N_15829);
nand U16900 (N_16900,N_15593,N_15396);
nor U16901 (N_16901,N_15905,N_15381);
nor U16902 (N_16902,N_15165,N_15455);
xor U16903 (N_16903,N_15796,N_15658);
nor U16904 (N_16904,N_15042,N_15778);
nand U16905 (N_16905,N_15345,N_15806);
and U16906 (N_16906,N_15416,N_15536);
nor U16907 (N_16907,N_15303,N_15924);
or U16908 (N_16908,N_15721,N_15595);
nor U16909 (N_16909,N_15163,N_15262);
nand U16910 (N_16910,N_15325,N_15101);
nor U16911 (N_16911,N_15639,N_15750);
or U16912 (N_16912,N_15066,N_15920);
nand U16913 (N_16913,N_15144,N_15513);
and U16914 (N_16914,N_15285,N_15658);
and U16915 (N_16915,N_15552,N_15472);
nor U16916 (N_16916,N_15114,N_15048);
nand U16917 (N_16917,N_15586,N_15177);
or U16918 (N_16918,N_15506,N_15059);
nand U16919 (N_16919,N_15889,N_15593);
nor U16920 (N_16920,N_15462,N_15825);
nand U16921 (N_16921,N_15982,N_15250);
nor U16922 (N_16922,N_15414,N_15577);
nand U16923 (N_16923,N_15698,N_15462);
nor U16924 (N_16924,N_15140,N_15106);
nand U16925 (N_16925,N_15214,N_15459);
nand U16926 (N_16926,N_15283,N_15913);
xnor U16927 (N_16927,N_15788,N_15967);
nand U16928 (N_16928,N_15253,N_15258);
nor U16929 (N_16929,N_15117,N_15376);
nand U16930 (N_16930,N_15256,N_15521);
and U16931 (N_16931,N_15555,N_15116);
and U16932 (N_16932,N_15684,N_15530);
nand U16933 (N_16933,N_15230,N_15357);
nor U16934 (N_16934,N_15630,N_15600);
nand U16935 (N_16935,N_15110,N_15594);
xor U16936 (N_16936,N_15096,N_15903);
nand U16937 (N_16937,N_15297,N_15067);
nand U16938 (N_16938,N_15876,N_15478);
nand U16939 (N_16939,N_15536,N_15376);
or U16940 (N_16940,N_15452,N_15552);
or U16941 (N_16941,N_15178,N_15241);
or U16942 (N_16942,N_15182,N_15843);
or U16943 (N_16943,N_15316,N_15621);
nor U16944 (N_16944,N_15533,N_15571);
or U16945 (N_16945,N_15434,N_15665);
xnor U16946 (N_16946,N_15596,N_15683);
or U16947 (N_16947,N_15014,N_15505);
and U16948 (N_16948,N_15142,N_15043);
or U16949 (N_16949,N_15472,N_15801);
xor U16950 (N_16950,N_15812,N_15390);
and U16951 (N_16951,N_15897,N_15253);
nand U16952 (N_16952,N_15045,N_15462);
nor U16953 (N_16953,N_15364,N_15169);
or U16954 (N_16954,N_15301,N_15714);
and U16955 (N_16955,N_15660,N_15908);
and U16956 (N_16956,N_15428,N_15717);
or U16957 (N_16957,N_15518,N_15613);
or U16958 (N_16958,N_15541,N_15527);
nor U16959 (N_16959,N_15663,N_15237);
xor U16960 (N_16960,N_15157,N_15442);
nand U16961 (N_16961,N_15215,N_15665);
nor U16962 (N_16962,N_15273,N_15889);
nand U16963 (N_16963,N_15541,N_15844);
nand U16964 (N_16964,N_15572,N_15390);
or U16965 (N_16965,N_15922,N_15347);
or U16966 (N_16966,N_15503,N_15616);
nand U16967 (N_16967,N_15716,N_15564);
xnor U16968 (N_16968,N_15739,N_15710);
or U16969 (N_16969,N_15420,N_15735);
xnor U16970 (N_16970,N_15770,N_15617);
and U16971 (N_16971,N_15886,N_15985);
and U16972 (N_16972,N_15325,N_15100);
nand U16973 (N_16973,N_15327,N_15794);
or U16974 (N_16974,N_15018,N_15782);
or U16975 (N_16975,N_15185,N_15114);
or U16976 (N_16976,N_15348,N_15150);
nor U16977 (N_16977,N_15146,N_15447);
nor U16978 (N_16978,N_15190,N_15164);
nand U16979 (N_16979,N_15949,N_15842);
or U16980 (N_16980,N_15456,N_15755);
nor U16981 (N_16981,N_15436,N_15699);
nor U16982 (N_16982,N_15471,N_15327);
or U16983 (N_16983,N_15832,N_15051);
nor U16984 (N_16984,N_15255,N_15275);
and U16985 (N_16985,N_15999,N_15725);
or U16986 (N_16986,N_15973,N_15593);
nand U16987 (N_16987,N_15736,N_15321);
nand U16988 (N_16988,N_15333,N_15461);
nand U16989 (N_16989,N_15549,N_15812);
xnor U16990 (N_16990,N_15579,N_15188);
xor U16991 (N_16991,N_15519,N_15373);
or U16992 (N_16992,N_15538,N_15265);
nand U16993 (N_16993,N_15105,N_15553);
nor U16994 (N_16994,N_15806,N_15380);
nand U16995 (N_16995,N_15426,N_15676);
and U16996 (N_16996,N_15569,N_15208);
nor U16997 (N_16997,N_15808,N_15260);
and U16998 (N_16998,N_15081,N_15302);
and U16999 (N_16999,N_15169,N_15075);
and U17000 (N_17000,N_16857,N_16154);
and U17001 (N_17001,N_16266,N_16715);
and U17002 (N_17002,N_16921,N_16671);
nand U17003 (N_17003,N_16637,N_16369);
or U17004 (N_17004,N_16994,N_16400);
and U17005 (N_17005,N_16679,N_16863);
nand U17006 (N_17006,N_16823,N_16457);
nor U17007 (N_17007,N_16646,N_16316);
or U17008 (N_17008,N_16327,N_16383);
nor U17009 (N_17009,N_16574,N_16467);
nor U17010 (N_17010,N_16880,N_16676);
nand U17011 (N_17011,N_16083,N_16523);
nor U17012 (N_17012,N_16524,N_16969);
or U17013 (N_17013,N_16270,N_16352);
and U17014 (N_17014,N_16726,N_16579);
or U17015 (N_17015,N_16746,N_16179);
nand U17016 (N_17016,N_16696,N_16714);
and U17017 (N_17017,N_16584,N_16985);
and U17018 (N_17018,N_16955,N_16599);
or U17019 (N_17019,N_16189,N_16056);
or U17020 (N_17020,N_16868,N_16058);
or U17021 (N_17021,N_16759,N_16820);
nor U17022 (N_17022,N_16354,N_16871);
and U17023 (N_17023,N_16368,N_16454);
xor U17024 (N_17024,N_16546,N_16009);
nand U17025 (N_17025,N_16918,N_16366);
xnor U17026 (N_17026,N_16935,N_16243);
nand U17027 (N_17027,N_16652,N_16982);
and U17028 (N_17028,N_16408,N_16041);
and U17029 (N_17029,N_16613,N_16735);
nor U17030 (N_17030,N_16993,N_16178);
nor U17031 (N_17031,N_16468,N_16604);
nand U17032 (N_17032,N_16013,N_16043);
or U17033 (N_17033,N_16989,N_16567);
nand U17034 (N_17034,N_16209,N_16160);
and U17035 (N_17035,N_16476,N_16502);
or U17036 (N_17036,N_16670,N_16601);
or U17037 (N_17037,N_16807,N_16732);
or U17038 (N_17038,N_16719,N_16940);
or U17039 (N_17039,N_16643,N_16277);
nand U17040 (N_17040,N_16936,N_16267);
or U17041 (N_17041,N_16626,N_16108);
and U17042 (N_17042,N_16288,N_16849);
and U17043 (N_17043,N_16365,N_16201);
and U17044 (N_17044,N_16012,N_16247);
or U17045 (N_17045,N_16183,N_16103);
nor U17046 (N_17046,N_16516,N_16278);
or U17047 (N_17047,N_16387,N_16256);
xor U17048 (N_17048,N_16177,N_16785);
xor U17049 (N_17049,N_16085,N_16490);
or U17050 (N_17050,N_16981,N_16385);
nor U17051 (N_17051,N_16057,N_16335);
nand U17052 (N_17052,N_16772,N_16202);
nand U17053 (N_17053,N_16246,N_16812);
nor U17054 (N_17054,N_16886,N_16059);
and U17055 (N_17055,N_16392,N_16691);
nand U17056 (N_17056,N_16787,N_16786);
and U17057 (N_17057,N_16867,N_16675);
or U17058 (N_17058,N_16410,N_16261);
or U17059 (N_17059,N_16141,N_16445);
or U17060 (N_17060,N_16583,N_16724);
xor U17061 (N_17061,N_16914,N_16832);
nor U17062 (N_17062,N_16110,N_16082);
nand U17063 (N_17063,N_16757,N_16139);
nand U17064 (N_17064,N_16238,N_16397);
and U17065 (N_17065,N_16663,N_16866);
nor U17066 (N_17066,N_16357,N_16314);
nand U17067 (N_17067,N_16176,N_16210);
or U17068 (N_17068,N_16928,N_16299);
and U17069 (N_17069,N_16016,N_16437);
nor U17070 (N_17070,N_16655,N_16435);
or U17071 (N_17071,N_16846,N_16121);
nor U17072 (N_17072,N_16023,N_16744);
nor U17073 (N_17073,N_16796,N_16349);
and U17074 (N_17074,N_16711,N_16231);
nor U17075 (N_17075,N_16406,N_16472);
nand U17076 (N_17076,N_16539,N_16608);
and U17077 (N_17077,N_16355,N_16263);
nor U17078 (N_17078,N_16856,N_16548);
nor U17079 (N_17079,N_16045,N_16004);
nand U17080 (N_17080,N_16708,N_16835);
nand U17081 (N_17081,N_16602,N_16011);
nand U17082 (N_17082,N_16014,N_16099);
nor U17083 (N_17083,N_16425,N_16146);
nand U17084 (N_17084,N_16345,N_16561);
and U17085 (N_17085,N_16782,N_16089);
nand U17086 (N_17086,N_16060,N_16126);
or U17087 (N_17087,N_16917,N_16883);
nand U17088 (N_17088,N_16098,N_16487);
and U17089 (N_17089,N_16875,N_16999);
nor U17090 (N_17090,N_16066,N_16162);
or U17091 (N_17091,N_16590,N_16802);
nand U17092 (N_17092,N_16976,N_16919);
nor U17093 (N_17093,N_16764,N_16658);
and U17094 (N_17094,N_16501,N_16434);
nand U17095 (N_17095,N_16455,N_16544);
or U17096 (N_17096,N_16821,N_16598);
nor U17097 (N_17097,N_16296,N_16610);
and U17098 (N_17098,N_16251,N_16444);
xnor U17099 (N_17099,N_16432,N_16331);
xor U17100 (N_17100,N_16594,N_16720);
or U17101 (N_17101,N_16614,N_16379);
nand U17102 (N_17102,N_16957,N_16493);
xor U17103 (N_17103,N_16566,N_16254);
nor U17104 (N_17104,N_16063,N_16843);
and U17105 (N_17105,N_16187,N_16079);
nand U17106 (N_17106,N_16326,N_16362);
or U17107 (N_17107,N_16104,N_16636);
or U17108 (N_17108,N_16514,N_16363);
nand U17109 (N_17109,N_16306,N_16689);
or U17110 (N_17110,N_16838,N_16713);
and U17111 (N_17111,N_16656,N_16905);
nand U17112 (N_17112,N_16239,N_16941);
and U17113 (N_17113,N_16088,N_16972);
xor U17114 (N_17114,N_16760,N_16305);
nand U17115 (N_17115,N_16390,N_16107);
or U17116 (N_17116,N_16244,N_16859);
nor U17117 (N_17117,N_16570,N_16117);
and U17118 (N_17118,N_16198,N_16519);
xor U17119 (N_17119,N_16386,N_16578);
nor U17120 (N_17120,N_16699,N_16906);
and U17121 (N_17121,N_16289,N_16394);
nand U17122 (N_17122,N_16471,N_16792);
or U17123 (N_17123,N_16228,N_16925);
xor U17124 (N_17124,N_16893,N_16865);
and U17125 (N_17125,N_16418,N_16855);
nand U17126 (N_17126,N_16414,N_16473);
nand U17127 (N_17127,N_16833,N_16252);
and U17128 (N_17128,N_16384,N_16814);
nand U17129 (N_17129,N_16460,N_16374);
nand U17130 (N_17130,N_16946,N_16742);
nor U17131 (N_17131,N_16743,N_16320);
or U17132 (N_17132,N_16236,N_16692);
nor U17133 (N_17133,N_16283,N_16970);
and U17134 (N_17134,N_16053,N_16974);
nor U17135 (N_17135,N_16144,N_16112);
xor U17136 (N_17136,N_16172,N_16947);
nor U17137 (N_17137,N_16262,N_16756);
or U17138 (N_17138,N_16419,N_16372);
nor U17139 (N_17139,N_16749,N_16297);
nor U17140 (N_17140,N_16870,N_16538);
or U17141 (N_17141,N_16540,N_16529);
xnor U17142 (N_17142,N_16453,N_16811);
xor U17143 (N_17143,N_16114,N_16517);
nor U17144 (N_17144,N_16125,N_16312);
and U17145 (N_17145,N_16790,N_16988);
nand U17146 (N_17146,N_16956,N_16775);
or U17147 (N_17147,N_16370,N_16361);
nand U17148 (N_17148,N_16442,N_16486);
nor U17149 (N_17149,N_16217,N_16282);
nor U17150 (N_17150,N_16153,N_16770);
nand U17151 (N_17151,N_16163,N_16309);
and U17152 (N_17152,N_16531,N_16255);
xor U17153 (N_17153,N_16226,N_16353);
nand U17154 (N_17154,N_16752,N_16428);
or U17155 (N_17155,N_16907,N_16642);
or U17156 (N_17156,N_16304,N_16142);
nand U17157 (N_17157,N_16470,N_16495);
and U17158 (N_17158,N_16559,N_16977);
or U17159 (N_17159,N_16723,N_16640);
or U17160 (N_17160,N_16730,N_16836);
and U17161 (N_17161,N_16431,N_16573);
nor U17162 (N_17162,N_16980,N_16618);
xor U17163 (N_17163,N_16151,N_16830);
and U17164 (N_17164,N_16841,N_16987);
nor U17165 (N_17165,N_16302,N_16284);
nand U17166 (N_17166,N_16729,N_16322);
nor U17167 (N_17167,N_16499,N_16959);
nor U17168 (N_17168,N_16482,N_16762);
or U17169 (N_17169,N_16157,N_16515);
nor U17170 (N_17170,N_16206,N_16525);
and U17171 (N_17171,N_16754,N_16170);
nand U17172 (N_17172,N_16033,N_16339);
or U17173 (N_17173,N_16116,N_16795);
nor U17174 (N_17174,N_16026,N_16155);
nor U17175 (N_17175,N_16801,N_16902);
nor U17176 (N_17176,N_16718,N_16845);
nor U17177 (N_17177,N_16556,N_16081);
xnor U17178 (N_17178,N_16965,N_16200);
nor U17179 (N_17179,N_16837,N_16076);
or U17180 (N_17180,N_16412,N_16269);
nor U17181 (N_17181,N_16565,N_16869);
and U17182 (N_17182,N_16440,N_16219);
nand U17183 (N_17183,N_16128,N_16564);
nor U17184 (N_17184,N_16595,N_16912);
nor U17185 (N_17185,N_16413,N_16364);
and U17186 (N_17186,N_16067,N_16257);
or U17187 (N_17187,N_16064,N_16568);
and U17188 (N_17188,N_16411,N_16332);
xor U17189 (N_17189,N_16481,N_16647);
xnor U17190 (N_17190,N_16650,N_16077);
nor U17191 (N_17191,N_16505,N_16586);
xnor U17192 (N_17192,N_16963,N_16951);
nand U17193 (N_17193,N_16190,N_16315);
nor U17194 (N_17194,N_16204,N_16196);
nor U17195 (N_17195,N_16851,N_16224);
or U17196 (N_17196,N_16300,N_16587);
nand U17197 (N_17197,N_16702,N_16736);
or U17198 (N_17198,N_16186,N_16904);
and U17199 (N_17199,N_16896,N_16264);
nor U17200 (N_17200,N_16070,N_16660);
nor U17201 (N_17201,N_16275,N_16235);
nor U17202 (N_17202,N_16221,N_16136);
nand U17203 (N_17203,N_16452,N_16734);
nand U17204 (N_17204,N_16265,N_16657);
xor U17205 (N_17205,N_16276,N_16769);
and U17206 (N_17206,N_16697,N_16822);
and U17207 (N_17207,N_16002,N_16684);
and U17208 (N_17208,N_16683,N_16952);
nand U17209 (N_17209,N_16616,N_16542);
and U17210 (N_17210,N_16813,N_16479);
or U17211 (N_17211,N_16403,N_16036);
nand U17212 (N_17212,N_16526,N_16380);
or U17213 (N_17213,N_16323,N_16130);
nor U17214 (N_17214,N_16872,N_16274);
xor U17215 (N_17215,N_16591,N_16712);
xnor U17216 (N_17216,N_16717,N_16527);
and U17217 (N_17217,N_16464,N_16954);
and U17218 (N_17218,N_16038,N_16042);
xor U17219 (N_17219,N_16627,N_16483);
nor U17220 (N_17220,N_16751,N_16208);
or U17221 (N_17221,N_16873,N_16168);
nand U17222 (N_17222,N_16480,N_16973);
xnor U17223 (N_17223,N_16503,N_16509);
nand U17224 (N_17224,N_16779,N_16840);
nand U17225 (N_17225,N_16436,N_16211);
or U17226 (N_17226,N_16592,N_16285);
or U17227 (N_17227,N_16609,N_16641);
nor U17228 (N_17228,N_16105,N_16260);
and U17229 (N_17229,N_16377,N_16000);
nor U17230 (N_17230,N_16337,N_16554);
nor U17231 (N_17231,N_16700,N_16273);
and U17232 (N_17232,N_16182,N_16903);
or U17233 (N_17233,N_16649,N_16205);
nor U17234 (N_17234,N_16706,N_16929);
nor U17235 (N_17235,N_16945,N_16253);
nand U17236 (N_17236,N_16203,N_16698);
and U17237 (N_17237,N_16961,N_16430);
nand U17238 (N_17238,N_16839,N_16055);
or U17239 (N_17239,N_16500,N_16924);
nor U17240 (N_17240,N_16688,N_16659);
and U17241 (N_17241,N_16890,N_16728);
and U17242 (N_17242,N_16932,N_16800);
xor U17243 (N_17243,N_16662,N_16341);
and U17244 (N_17244,N_16996,N_16010);
nor U17245 (N_17245,N_16465,N_16844);
nor U17246 (N_17246,N_16447,N_16311);
nand U17247 (N_17247,N_16100,N_16831);
nand U17248 (N_17248,N_16740,N_16789);
and U17249 (N_17249,N_16777,N_16421);
nand U17250 (N_17250,N_16901,N_16678);
nand U17251 (N_17251,N_16555,N_16143);
nor U17252 (N_17252,N_16521,N_16635);
nand U17253 (N_17253,N_16569,N_16021);
xnor U17254 (N_17254,N_16307,N_16860);
and U17255 (N_17255,N_16420,N_16218);
nor U17256 (N_17256,N_16159,N_16137);
nor U17257 (N_17257,N_16249,N_16286);
nor U17258 (N_17258,N_16737,N_16407);
nor U17259 (N_17259,N_16603,N_16047);
or U17260 (N_17260,N_16279,N_16597);
nand U17261 (N_17261,N_16984,N_16448);
or U17262 (N_17262,N_16639,N_16805);
or U17263 (N_17263,N_16313,N_16581);
nand U17264 (N_17264,N_16920,N_16328);
nand U17265 (N_17265,N_16577,N_16827);
and U17266 (N_17266,N_16998,N_16024);
nand U17267 (N_17267,N_16359,N_16788);
nor U17268 (N_17268,N_16551,N_16340);
nand U17269 (N_17269,N_16888,N_16475);
and U17270 (N_17270,N_16572,N_16072);
nand U17271 (N_17271,N_16381,N_16214);
and U17272 (N_17272,N_16496,N_16884);
and U17273 (N_17273,N_16039,N_16763);
xnor U17274 (N_17274,N_16900,N_16654);
nor U17275 (N_17275,N_16804,N_16008);
nor U17276 (N_17276,N_16979,N_16096);
nor U17277 (N_17277,N_16032,N_16748);
and U17278 (N_17278,N_16828,N_16050);
nor U17279 (N_17279,N_16768,N_16975);
nand U17280 (N_17280,N_16062,N_16001);
and U17281 (N_17281,N_16847,N_16491);
xor U17282 (N_17282,N_16817,N_16135);
or U17283 (N_17283,N_16124,N_16113);
xor U17284 (N_17284,N_16780,N_16510);
or U17285 (N_17285,N_16092,N_16793);
nand U17286 (N_17286,N_16351,N_16739);
nand U17287 (N_17287,N_16894,N_16395);
and U17288 (N_17288,N_16356,N_16575);
or U17289 (N_17289,N_16899,N_16375);
or U17290 (N_17290,N_16596,N_16223);
nand U17291 (N_17291,N_16664,N_16622);
and U17292 (N_17292,N_16798,N_16552);
nor U17293 (N_17293,N_16926,N_16477);
nand U17294 (N_17294,N_16281,N_16336);
nand U17295 (N_17295,N_16416,N_16766);
and U17296 (N_17296,N_16240,N_16382);
nor U17297 (N_17297,N_16446,N_16250);
nand U17298 (N_17298,N_16343,N_16776);
nor U17299 (N_17299,N_16630,N_16750);
nand U17300 (N_17300,N_16438,N_16019);
nor U17301 (N_17301,N_16722,N_16794);
nor U17302 (N_17302,N_16498,N_16148);
nand U17303 (N_17303,N_16119,N_16334);
nor U17304 (N_17304,N_16826,N_16194);
nand U17305 (N_17305,N_16582,N_16451);
nand U17306 (N_17306,N_16967,N_16488);
xnor U17307 (N_17307,N_16199,N_16680);
nand U17308 (N_17308,N_16753,N_16156);
or U17309 (N_17309,N_16378,N_16771);
nand U17310 (N_17310,N_16166,N_16731);
nand U17311 (N_17311,N_16129,N_16553);
nand U17312 (N_17312,N_16758,N_16034);
and U17313 (N_17313,N_16450,N_16086);
or U17314 (N_17314,N_16950,N_16549);
and U17315 (N_17315,N_16185,N_16842);
nor U17316 (N_17316,N_16733,N_16075);
or U17317 (N_17317,N_16978,N_16234);
nand U17318 (N_17318,N_16910,N_16167);
and U17319 (N_17319,N_16983,N_16628);
or U17320 (N_17320,N_16301,N_16463);
or U17321 (N_17321,N_16061,N_16535);
nor U17322 (N_17322,N_16741,N_16396);
nor U17323 (N_17323,N_16922,N_16358);
nand U17324 (N_17324,N_16485,N_16933);
nor U17325 (N_17325,N_16120,N_16459);
and U17326 (N_17326,N_16293,N_16207);
nand U17327 (N_17327,N_16492,N_16881);
nand U17328 (N_17328,N_16621,N_16931);
nor U17329 (N_17329,N_16044,N_16667);
or U17330 (N_17330,N_16291,N_16885);
nor U17331 (N_17331,N_16773,N_16709);
nand U17332 (N_17332,N_16550,N_16259);
or U17333 (N_17333,N_16938,N_16342);
xor U17334 (N_17334,N_16990,N_16220);
xnor U17335 (N_17335,N_16687,N_16571);
and U17336 (N_17336,N_16791,N_16149);
nor U17337 (N_17337,N_16816,N_16638);
nor U17338 (N_17338,N_16541,N_16031);
and U17339 (N_17339,N_16939,N_16986);
or U17340 (N_17340,N_16037,N_16703);
nand U17341 (N_17341,N_16877,N_16686);
nor U17342 (N_17342,N_16192,N_16547);
or U17343 (N_17343,N_16666,N_16625);
or U17344 (N_17344,N_16029,N_16417);
nor U17345 (N_17345,N_16545,N_16048);
nor U17346 (N_17346,N_16290,N_16393);
and U17347 (N_17347,N_16864,N_16909);
or U17348 (N_17348,N_16028,N_16188);
or U17349 (N_17349,N_16373,N_16242);
nor U17350 (N_17350,N_16858,N_16213);
nand U17351 (N_17351,N_16850,N_16399);
nor U17352 (N_17352,N_16040,N_16404);
or U17353 (N_17353,N_16593,N_16681);
and U17354 (N_17354,N_16433,N_16484);
xnor U17355 (N_17355,N_16725,N_16150);
nand U17356 (N_17356,N_16997,N_16215);
and U17357 (N_17357,N_16512,N_16180);
and U17358 (N_17358,N_16422,N_16797);
and U17359 (N_17359,N_16248,N_16809);
and U17360 (N_17360,N_16644,N_16930);
xnor U17361 (N_17361,N_16767,N_16443);
xnor U17362 (N_17362,N_16109,N_16876);
or U17363 (N_17363,N_16348,N_16949);
xnor U17364 (N_17364,N_16035,N_16562);
and U17365 (N_17365,N_16049,N_16536);
or U17366 (N_17366,N_16073,N_16147);
nand U17367 (N_17367,N_16887,N_16003);
xnor U17368 (N_17368,N_16164,N_16669);
xor U17369 (N_17369,N_16069,N_16087);
and U17370 (N_17370,N_16494,N_16175);
and U17371 (N_17371,N_16115,N_16027);
nor U17372 (N_17372,N_16580,N_16169);
nor U17373 (N_17373,N_16878,N_16915);
nor U17374 (N_17374,N_16645,N_16405);
nor U17375 (N_17375,N_16389,N_16294);
or U17376 (N_17376,N_16629,N_16449);
or U17377 (N_17377,N_16962,N_16534);
or U17378 (N_17378,N_16783,N_16233);
and U17379 (N_17379,N_16632,N_16818);
or U17380 (N_17380,N_16543,N_16462);
and U17381 (N_17381,N_16513,N_16815);
and U17382 (N_17382,N_16619,N_16272);
or U17383 (N_17383,N_16585,N_16191);
or U17384 (N_17384,N_16690,N_16781);
or U17385 (N_17385,N_16518,N_16258);
and U17386 (N_17386,N_16469,N_16889);
or U17387 (N_17387,N_16908,N_16693);
or U17388 (N_17388,N_16367,N_16091);
or U17389 (N_17389,N_16497,N_16046);
nand U17390 (N_17390,N_16966,N_16682);
nand U17391 (N_17391,N_16230,N_16897);
and U17392 (N_17392,N_16212,N_16829);
xnor U17393 (N_17393,N_16563,N_16995);
nand U17394 (N_17394,N_16017,N_16015);
or U17395 (N_17395,N_16461,N_16426);
nand U17396 (N_17396,N_16537,N_16222);
or U17397 (N_17397,N_16507,N_16799);
and U17398 (N_17398,N_16953,N_16853);
nor U17399 (N_17399,N_16329,N_16376);
or U17400 (N_17400,N_16911,N_16942);
and U17401 (N_17401,N_16106,N_16707);
and U17402 (N_17402,N_16466,N_16227);
and U17403 (N_17403,N_16268,N_16765);
nor U17404 (N_17404,N_16078,N_16441);
nor U17405 (N_17405,N_16068,N_16745);
nor U17406 (N_17406,N_16806,N_16716);
and U17407 (N_17407,N_16522,N_16232);
nor U17408 (N_17408,N_16152,N_16895);
or U17409 (N_17409,N_16344,N_16852);
nor U17410 (N_17410,N_16287,N_16080);
nand U17411 (N_17411,N_16648,N_16424);
nand U17412 (N_17412,N_16530,N_16558);
and U17413 (N_17413,N_16971,N_16427);
nand U17414 (N_17414,N_16350,N_16052);
or U17415 (N_17415,N_16118,N_16511);
xor U17416 (N_17416,N_16456,N_16409);
nor U17417 (N_17417,N_16808,N_16891);
nand U17418 (N_17418,N_16216,N_16158);
nand U17419 (N_17419,N_16668,N_16097);
nor U17420 (N_17420,N_16923,N_16774);
and U17421 (N_17421,N_16892,N_16054);
nor U17422 (N_17422,N_16007,N_16111);
and U17423 (N_17423,N_16721,N_16898);
nor U17424 (N_17424,N_16913,N_16321);
or U17425 (N_17425,N_16755,N_16308);
or U17426 (N_17426,N_16333,N_16402);
nand U17427 (N_17427,N_16489,N_16325);
xor U17428 (N_17428,N_16727,N_16295);
nand U17429 (N_17429,N_16324,N_16138);
nand U17430 (N_17430,N_16197,N_16673);
and U17431 (N_17431,N_16819,N_16653);
nand U17432 (N_17432,N_16298,N_16508);
nand U17433 (N_17433,N_16127,N_16123);
and U17434 (N_17434,N_16161,N_16589);
or U17435 (N_17435,N_16292,N_16825);
and U17436 (N_17436,N_16310,N_16834);
and U17437 (N_17437,N_16346,N_16131);
xor U17438 (N_17438,N_16705,N_16303);
xor U17439 (N_17439,N_16458,N_16319);
xnor U17440 (N_17440,N_16854,N_16824);
nor U17441 (N_17441,N_16391,N_16145);
and U17442 (N_17442,N_16195,N_16174);
or U17443 (N_17443,N_16371,N_16576);
or U17444 (N_17444,N_16937,N_16051);
nor U17445 (N_17445,N_16677,N_16784);
and U17446 (N_17446,N_16694,N_16624);
xor U17447 (N_17447,N_16992,N_16193);
or U17448 (N_17448,N_16943,N_16738);
nor U17449 (N_17449,N_16623,N_16241);
nand U17450 (N_17450,N_16101,N_16803);
xor U17451 (N_17451,N_16347,N_16588);
nor U17452 (N_17452,N_16122,N_16948);
nor U17453 (N_17453,N_16018,N_16964);
or U17454 (N_17454,N_16225,N_16605);
and U17455 (N_17455,N_16478,N_16318);
xnor U17456 (N_17456,N_16074,N_16862);
and U17457 (N_17457,N_16958,N_16006);
nor U17458 (N_17458,N_16095,N_16672);
or U17459 (N_17459,N_16474,N_16528);
nor U17460 (N_17460,N_16005,N_16022);
nor U17461 (N_17461,N_16093,N_16944);
and U17462 (N_17462,N_16600,N_16271);
nor U17463 (N_17463,N_16317,N_16848);
nand U17464 (N_17464,N_16633,N_16612);
xor U17465 (N_17465,N_16415,N_16090);
nor U17466 (N_17466,N_16171,N_16607);
or U17467 (N_17467,N_16934,N_16388);
nor U17468 (N_17468,N_16631,N_16181);
or U17469 (N_17469,N_16094,N_16991);
nand U17470 (N_17470,N_16710,N_16674);
or U17471 (N_17471,N_16184,N_16398);
and U17472 (N_17472,N_16916,N_16882);
or U17473 (N_17473,N_16701,N_16165);
and U17474 (N_17474,N_16423,N_16778);
nand U17475 (N_17475,N_16065,N_16429);
and U17476 (N_17476,N_16617,N_16695);
nor U17477 (N_17477,N_16560,N_16338);
or U17478 (N_17478,N_16132,N_16360);
xnor U17479 (N_17479,N_16133,N_16874);
nor U17480 (N_17480,N_16520,N_16140);
nor U17481 (N_17481,N_16532,N_16506);
and U17482 (N_17482,N_16173,N_16611);
xor U17483 (N_17483,N_16439,N_16134);
xnor U17484 (N_17484,N_16504,N_16665);
nand U17485 (N_17485,N_16102,N_16401);
xor U17486 (N_17486,N_16747,N_16651);
and U17487 (N_17487,N_16615,N_16533);
and U17488 (N_17488,N_16229,N_16237);
and U17489 (N_17489,N_16761,N_16025);
or U17490 (N_17490,N_16685,N_16879);
or U17491 (N_17491,N_16557,N_16661);
nor U17492 (N_17492,N_16810,N_16071);
and U17493 (N_17493,N_16861,N_16606);
and U17494 (N_17494,N_16968,N_16927);
nor U17495 (N_17495,N_16960,N_16634);
nor U17496 (N_17496,N_16245,N_16330);
xnor U17497 (N_17497,N_16020,N_16084);
nand U17498 (N_17498,N_16704,N_16030);
and U17499 (N_17499,N_16620,N_16280);
or U17500 (N_17500,N_16389,N_16137);
nand U17501 (N_17501,N_16719,N_16402);
and U17502 (N_17502,N_16327,N_16524);
or U17503 (N_17503,N_16667,N_16713);
nor U17504 (N_17504,N_16774,N_16182);
nor U17505 (N_17505,N_16127,N_16960);
or U17506 (N_17506,N_16307,N_16627);
nor U17507 (N_17507,N_16086,N_16526);
nand U17508 (N_17508,N_16344,N_16996);
nor U17509 (N_17509,N_16199,N_16957);
nand U17510 (N_17510,N_16450,N_16895);
nor U17511 (N_17511,N_16064,N_16347);
xnor U17512 (N_17512,N_16540,N_16703);
nand U17513 (N_17513,N_16994,N_16712);
nand U17514 (N_17514,N_16008,N_16361);
nor U17515 (N_17515,N_16592,N_16304);
and U17516 (N_17516,N_16855,N_16387);
and U17517 (N_17517,N_16304,N_16227);
and U17518 (N_17518,N_16754,N_16779);
and U17519 (N_17519,N_16517,N_16636);
nand U17520 (N_17520,N_16660,N_16048);
or U17521 (N_17521,N_16903,N_16992);
and U17522 (N_17522,N_16764,N_16392);
nand U17523 (N_17523,N_16021,N_16828);
nand U17524 (N_17524,N_16997,N_16347);
and U17525 (N_17525,N_16190,N_16766);
xor U17526 (N_17526,N_16208,N_16195);
nor U17527 (N_17527,N_16116,N_16947);
nand U17528 (N_17528,N_16075,N_16881);
or U17529 (N_17529,N_16469,N_16030);
or U17530 (N_17530,N_16231,N_16917);
or U17531 (N_17531,N_16381,N_16608);
nor U17532 (N_17532,N_16613,N_16270);
nor U17533 (N_17533,N_16346,N_16811);
nor U17534 (N_17534,N_16813,N_16107);
or U17535 (N_17535,N_16613,N_16573);
nand U17536 (N_17536,N_16287,N_16930);
or U17537 (N_17537,N_16295,N_16122);
nor U17538 (N_17538,N_16917,N_16970);
nor U17539 (N_17539,N_16379,N_16866);
nor U17540 (N_17540,N_16827,N_16816);
nor U17541 (N_17541,N_16225,N_16980);
or U17542 (N_17542,N_16629,N_16936);
and U17543 (N_17543,N_16203,N_16236);
and U17544 (N_17544,N_16821,N_16731);
nor U17545 (N_17545,N_16870,N_16916);
or U17546 (N_17546,N_16311,N_16060);
or U17547 (N_17547,N_16261,N_16437);
nor U17548 (N_17548,N_16253,N_16557);
xnor U17549 (N_17549,N_16013,N_16732);
and U17550 (N_17550,N_16087,N_16339);
and U17551 (N_17551,N_16418,N_16340);
or U17552 (N_17552,N_16752,N_16488);
nand U17553 (N_17553,N_16316,N_16025);
or U17554 (N_17554,N_16253,N_16724);
nor U17555 (N_17555,N_16164,N_16036);
nand U17556 (N_17556,N_16086,N_16146);
nand U17557 (N_17557,N_16418,N_16481);
nor U17558 (N_17558,N_16810,N_16193);
and U17559 (N_17559,N_16090,N_16294);
nor U17560 (N_17560,N_16374,N_16609);
nor U17561 (N_17561,N_16180,N_16120);
and U17562 (N_17562,N_16749,N_16845);
xnor U17563 (N_17563,N_16148,N_16798);
xnor U17564 (N_17564,N_16421,N_16575);
nor U17565 (N_17565,N_16378,N_16050);
and U17566 (N_17566,N_16782,N_16861);
or U17567 (N_17567,N_16197,N_16799);
and U17568 (N_17568,N_16377,N_16293);
nor U17569 (N_17569,N_16257,N_16665);
or U17570 (N_17570,N_16831,N_16687);
nand U17571 (N_17571,N_16026,N_16109);
xor U17572 (N_17572,N_16066,N_16851);
nor U17573 (N_17573,N_16962,N_16245);
nand U17574 (N_17574,N_16322,N_16987);
or U17575 (N_17575,N_16724,N_16633);
and U17576 (N_17576,N_16655,N_16204);
or U17577 (N_17577,N_16310,N_16348);
and U17578 (N_17578,N_16416,N_16546);
nor U17579 (N_17579,N_16437,N_16443);
xor U17580 (N_17580,N_16720,N_16567);
or U17581 (N_17581,N_16508,N_16819);
xnor U17582 (N_17582,N_16657,N_16517);
or U17583 (N_17583,N_16281,N_16773);
nor U17584 (N_17584,N_16565,N_16711);
and U17585 (N_17585,N_16607,N_16854);
nor U17586 (N_17586,N_16496,N_16167);
and U17587 (N_17587,N_16854,N_16073);
nor U17588 (N_17588,N_16756,N_16094);
xor U17589 (N_17589,N_16469,N_16103);
nand U17590 (N_17590,N_16883,N_16290);
nand U17591 (N_17591,N_16275,N_16151);
nor U17592 (N_17592,N_16575,N_16792);
or U17593 (N_17593,N_16053,N_16369);
nand U17594 (N_17594,N_16154,N_16004);
or U17595 (N_17595,N_16316,N_16398);
nor U17596 (N_17596,N_16054,N_16875);
nor U17597 (N_17597,N_16515,N_16706);
and U17598 (N_17598,N_16857,N_16326);
xor U17599 (N_17599,N_16258,N_16393);
and U17600 (N_17600,N_16221,N_16638);
nor U17601 (N_17601,N_16695,N_16356);
nor U17602 (N_17602,N_16788,N_16620);
and U17603 (N_17603,N_16990,N_16715);
nand U17604 (N_17604,N_16388,N_16350);
or U17605 (N_17605,N_16071,N_16025);
nor U17606 (N_17606,N_16896,N_16955);
xor U17607 (N_17607,N_16672,N_16370);
and U17608 (N_17608,N_16703,N_16010);
nand U17609 (N_17609,N_16743,N_16612);
or U17610 (N_17610,N_16952,N_16086);
or U17611 (N_17611,N_16601,N_16032);
and U17612 (N_17612,N_16206,N_16331);
or U17613 (N_17613,N_16815,N_16273);
and U17614 (N_17614,N_16552,N_16050);
nor U17615 (N_17615,N_16357,N_16352);
nand U17616 (N_17616,N_16236,N_16702);
or U17617 (N_17617,N_16982,N_16622);
nand U17618 (N_17618,N_16523,N_16526);
xnor U17619 (N_17619,N_16631,N_16834);
and U17620 (N_17620,N_16672,N_16003);
and U17621 (N_17621,N_16015,N_16342);
nor U17622 (N_17622,N_16531,N_16619);
nand U17623 (N_17623,N_16878,N_16665);
nand U17624 (N_17624,N_16351,N_16328);
nand U17625 (N_17625,N_16677,N_16783);
and U17626 (N_17626,N_16411,N_16394);
nand U17627 (N_17627,N_16244,N_16451);
or U17628 (N_17628,N_16157,N_16574);
and U17629 (N_17629,N_16561,N_16767);
and U17630 (N_17630,N_16988,N_16550);
xnor U17631 (N_17631,N_16829,N_16375);
and U17632 (N_17632,N_16108,N_16838);
and U17633 (N_17633,N_16965,N_16928);
or U17634 (N_17634,N_16360,N_16526);
nand U17635 (N_17635,N_16644,N_16297);
nand U17636 (N_17636,N_16970,N_16053);
or U17637 (N_17637,N_16647,N_16169);
or U17638 (N_17638,N_16157,N_16338);
and U17639 (N_17639,N_16348,N_16503);
nor U17640 (N_17640,N_16383,N_16483);
xnor U17641 (N_17641,N_16452,N_16051);
and U17642 (N_17642,N_16806,N_16529);
or U17643 (N_17643,N_16002,N_16236);
nand U17644 (N_17644,N_16800,N_16102);
nand U17645 (N_17645,N_16865,N_16113);
xor U17646 (N_17646,N_16155,N_16946);
and U17647 (N_17647,N_16399,N_16185);
or U17648 (N_17648,N_16197,N_16710);
nand U17649 (N_17649,N_16098,N_16754);
nor U17650 (N_17650,N_16357,N_16452);
and U17651 (N_17651,N_16213,N_16782);
nor U17652 (N_17652,N_16133,N_16007);
or U17653 (N_17653,N_16655,N_16445);
nand U17654 (N_17654,N_16890,N_16641);
nor U17655 (N_17655,N_16030,N_16309);
and U17656 (N_17656,N_16346,N_16593);
or U17657 (N_17657,N_16909,N_16602);
nor U17658 (N_17658,N_16462,N_16390);
or U17659 (N_17659,N_16047,N_16341);
or U17660 (N_17660,N_16922,N_16356);
nor U17661 (N_17661,N_16868,N_16446);
or U17662 (N_17662,N_16152,N_16317);
or U17663 (N_17663,N_16749,N_16097);
or U17664 (N_17664,N_16684,N_16532);
or U17665 (N_17665,N_16882,N_16200);
or U17666 (N_17666,N_16894,N_16624);
xor U17667 (N_17667,N_16929,N_16441);
xnor U17668 (N_17668,N_16081,N_16182);
xor U17669 (N_17669,N_16180,N_16114);
and U17670 (N_17670,N_16208,N_16000);
or U17671 (N_17671,N_16233,N_16865);
nand U17672 (N_17672,N_16780,N_16022);
xor U17673 (N_17673,N_16979,N_16187);
and U17674 (N_17674,N_16304,N_16759);
nand U17675 (N_17675,N_16403,N_16404);
or U17676 (N_17676,N_16674,N_16804);
and U17677 (N_17677,N_16295,N_16353);
nand U17678 (N_17678,N_16845,N_16449);
xor U17679 (N_17679,N_16472,N_16741);
nor U17680 (N_17680,N_16421,N_16437);
or U17681 (N_17681,N_16397,N_16910);
xnor U17682 (N_17682,N_16767,N_16424);
or U17683 (N_17683,N_16562,N_16527);
nand U17684 (N_17684,N_16987,N_16517);
or U17685 (N_17685,N_16608,N_16837);
or U17686 (N_17686,N_16010,N_16013);
xnor U17687 (N_17687,N_16995,N_16493);
xnor U17688 (N_17688,N_16523,N_16399);
and U17689 (N_17689,N_16558,N_16964);
nor U17690 (N_17690,N_16422,N_16055);
nand U17691 (N_17691,N_16618,N_16497);
xor U17692 (N_17692,N_16972,N_16425);
nor U17693 (N_17693,N_16464,N_16751);
nor U17694 (N_17694,N_16096,N_16209);
nor U17695 (N_17695,N_16572,N_16303);
nand U17696 (N_17696,N_16148,N_16376);
nand U17697 (N_17697,N_16887,N_16824);
and U17698 (N_17698,N_16282,N_16128);
or U17699 (N_17699,N_16743,N_16708);
or U17700 (N_17700,N_16794,N_16937);
nand U17701 (N_17701,N_16827,N_16930);
or U17702 (N_17702,N_16356,N_16559);
nor U17703 (N_17703,N_16616,N_16443);
or U17704 (N_17704,N_16628,N_16646);
and U17705 (N_17705,N_16631,N_16427);
nor U17706 (N_17706,N_16829,N_16099);
and U17707 (N_17707,N_16818,N_16584);
nor U17708 (N_17708,N_16583,N_16647);
and U17709 (N_17709,N_16598,N_16950);
or U17710 (N_17710,N_16318,N_16564);
and U17711 (N_17711,N_16035,N_16279);
or U17712 (N_17712,N_16961,N_16002);
nand U17713 (N_17713,N_16154,N_16329);
nand U17714 (N_17714,N_16565,N_16361);
nand U17715 (N_17715,N_16147,N_16084);
nand U17716 (N_17716,N_16889,N_16853);
and U17717 (N_17717,N_16156,N_16272);
or U17718 (N_17718,N_16134,N_16079);
nor U17719 (N_17719,N_16206,N_16145);
and U17720 (N_17720,N_16441,N_16007);
xnor U17721 (N_17721,N_16325,N_16895);
nand U17722 (N_17722,N_16779,N_16555);
xor U17723 (N_17723,N_16144,N_16541);
or U17724 (N_17724,N_16363,N_16248);
nand U17725 (N_17725,N_16603,N_16245);
nand U17726 (N_17726,N_16660,N_16077);
nand U17727 (N_17727,N_16661,N_16559);
nor U17728 (N_17728,N_16432,N_16456);
and U17729 (N_17729,N_16900,N_16496);
and U17730 (N_17730,N_16692,N_16367);
or U17731 (N_17731,N_16930,N_16705);
nand U17732 (N_17732,N_16266,N_16890);
nor U17733 (N_17733,N_16097,N_16884);
or U17734 (N_17734,N_16765,N_16414);
or U17735 (N_17735,N_16358,N_16151);
nand U17736 (N_17736,N_16421,N_16508);
nor U17737 (N_17737,N_16547,N_16207);
nor U17738 (N_17738,N_16826,N_16328);
xnor U17739 (N_17739,N_16794,N_16032);
nand U17740 (N_17740,N_16306,N_16686);
or U17741 (N_17741,N_16563,N_16886);
xnor U17742 (N_17742,N_16038,N_16248);
nor U17743 (N_17743,N_16067,N_16084);
nor U17744 (N_17744,N_16265,N_16523);
nand U17745 (N_17745,N_16686,N_16703);
nor U17746 (N_17746,N_16646,N_16171);
or U17747 (N_17747,N_16527,N_16053);
xnor U17748 (N_17748,N_16548,N_16845);
nor U17749 (N_17749,N_16820,N_16314);
nand U17750 (N_17750,N_16973,N_16751);
nand U17751 (N_17751,N_16483,N_16439);
nand U17752 (N_17752,N_16884,N_16757);
and U17753 (N_17753,N_16999,N_16476);
nor U17754 (N_17754,N_16659,N_16742);
and U17755 (N_17755,N_16253,N_16928);
nor U17756 (N_17756,N_16021,N_16534);
nor U17757 (N_17757,N_16638,N_16229);
nor U17758 (N_17758,N_16900,N_16961);
nor U17759 (N_17759,N_16363,N_16463);
and U17760 (N_17760,N_16525,N_16492);
xnor U17761 (N_17761,N_16580,N_16162);
and U17762 (N_17762,N_16348,N_16119);
and U17763 (N_17763,N_16040,N_16578);
xor U17764 (N_17764,N_16747,N_16739);
or U17765 (N_17765,N_16571,N_16827);
nand U17766 (N_17766,N_16670,N_16512);
or U17767 (N_17767,N_16955,N_16719);
nand U17768 (N_17768,N_16800,N_16229);
nand U17769 (N_17769,N_16738,N_16750);
nand U17770 (N_17770,N_16026,N_16776);
and U17771 (N_17771,N_16469,N_16156);
and U17772 (N_17772,N_16357,N_16021);
and U17773 (N_17773,N_16998,N_16815);
nand U17774 (N_17774,N_16873,N_16733);
nand U17775 (N_17775,N_16457,N_16033);
nand U17776 (N_17776,N_16750,N_16293);
nor U17777 (N_17777,N_16459,N_16342);
nand U17778 (N_17778,N_16065,N_16899);
nand U17779 (N_17779,N_16841,N_16850);
xor U17780 (N_17780,N_16614,N_16599);
nand U17781 (N_17781,N_16023,N_16942);
or U17782 (N_17782,N_16486,N_16956);
and U17783 (N_17783,N_16337,N_16539);
nand U17784 (N_17784,N_16623,N_16208);
and U17785 (N_17785,N_16436,N_16463);
or U17786 (N_17786,N_16467,N_16347);
nand U17787 (N_17787,N_16530,N_16018);
nand U17788 (N_17788,N_16585,N_16419);
nor U17789 (N_17789,N_16030,N_16579);
nor U17790 (N_17790,N_16210,N_16692);
or U17791 (N_17791,N_16627,N_16447);
or U17792 (N_17792,N_16563,N_16311);
nand U17793 (N_17793,N_16205,N_16187);
nand U17794 (N_17794,N_16182,N_16374);
nand U17795 (N_17795,N_16444,N_16506);
nor U17796 (N_17796,N_16344,N_16138);
or U17797 (N_17797,N_16054,N_16377);
and U17798 (N_17798,N_16644,N_16452);
xnor U17799 (N_17799,N_16087,N_16238);
and U17800 (N_17800,N_16753,N_16941);
and U17801 (N_17801,N_16118,N_16120);
nand U17802 (N_17802,N_16968,N_16770);
or U17803 (N_17803,N_16685,N_16352);
nor U17804 (N_17804,N_16826,N_16578);
nor U17805 (N_17805,N_16765,N_16736);
nor U17806 (N_17806,N_16726,N_16563);
nand U17807 (N_17807,N_16964,N_16839);
nand U17808 (N_17808,N_16217,N_16798);
nor U17809 (N_17809,N_16809,N_16451);
or U17810 (N_17810,N_16386,N_16446);
and U17811 (N_17811,N_16244,N_16613);
and U17812 (N_17812,N_16728,N_16674);
xnor U17813 (N_17813,N_16933,N_16012);
nor U17814 (N_17814,N_16746,N_16519);
xnor U17815 (N_17815,N_16252,N_16310);
nor U17816 (N_17816,N_16029,N_16104);
nor U17817 (N_17817,N_16585,N_16404);
nor U17818 (N_17818,N_16290,N_16841);
and U17819 (N_17819,N_16564,N_16541);
and U17820 (N_17820,N_16241,N_16110);
nor U17821 (N_17821,N_16217,N_16409);
and U17822 (N_17822,N_16247,N_16813);
nor U17823 (N_17823,N_16539,N_16817);
nor U17824 (N_17824,N_16482,N_16879);
xor U17825 (N_17825,N_16680,N_16071);
or U17826 (N_17826,N_16227,N_16970);
and U17827 (N_17827,N_16076,N_16788);
or U17828 (N_17828,N_16910,N_16819);
nand U17829 (N_17829,N_16749,N_16222);
or U17830 (N_17830,N_16059,N_16266);
nor U17831 (N_17831,N_16476,N_16947);
xor U17832 (N_17832,N_16100,N_16469);
nand U17833 (N_17833,N_16148,N_16241);
nor U17834 (N_17834,N_16156,N_16001);
nor U17835 (N_17835,N_16881,N_16796);
nor U17836 (N_17836,N_16103,N_16637);
and U17837 (N_17837,N_16859,N_16965);
nand U17838 (N_17838,N_16164,N_16192);
nand U17839 (N_17839,N_16825,N_16661);
or U17840 (N_17840,N_16980,N_16630);
xnor U17841 (N_17841,N_16836,N_16031);
nor U17842 (N_17842,N_16370,N_16151);
or U17843 (N_17843,N_16797,N_16242);
xor U17844 (N_17844,N_16725,N_16157);
nor U17845 (N_17845,N_16991,N_16847);
nand U17846 (N_17846,N_16017,N_16656);
and U17847 (N_17847,N_16127,N_16743);
or U17848 (N_17848,N_16808,N_16085);
or U17849 (N_17849,N_16254,N_16193);
xor U17850 (N_17850,N_16434,N_16918);
xnor U17851 (N_17851,N_16095,N_16036);
nand U17852 (N_17852,N_16150,N_16521);
nor U17853 (N_17853,N_16334,N_16729);
xor U17854 (N_17854,N_16776,N_16725);
or U17855 (N_17855,N_16265,N_16189);
and U17856 (N_17856,N_16509,N_16911);
xor U17857 (N_17857,N_16447,N_16448);
and U17858 (N_17858,N_16288,N_16614);
nor U17859 (N_17859,N_16866,N_16989);
nor U17860 (N_17860,N_16534,N_16935);
and U17861 (N_17861,N_16901,N_16861);
nor U17862 (N_17862,N_16349,N_16475);
and U17863 (N_17863,N_16735,N_16977);
nand U17864 (N_17864,N_16616,N_16400);
nand U17865 (N_17865,N_16840,N_16879);
or U17866 (N_17866,N_16234,N_16336);
or U17867 (N_17867,N_16056,N_16819);
and U17868 (N_17868,N_16784,N_16566);
nor U17869 (N_17869,N_16042,N_16440);
xnor U17870 (N_17870,N_16233,N_16270);
or U17871 (N_17871,N_16151,N_16109);
nand U17872 (N_17872,N_16442,N_16784);
nor U17873 (N_17873,N_16588,N_16993);
nand U17874 (N_17874,N_16827,N_16051);
and U17875 (N_17875,N_16110,N_16316);
xor U17876 (N_17876,N_16209,N_16273);
nor U17877 (N_17877,N_16274,N_16464);
or U17878 (N_17878,N_16476,N_16434);
nand U17879 (N_17879,N_16297,N_16030);
or U17880 (N_17880,N_16542,N_16623);
xor U17881 (N_17881,N_16239,N_16320);
and U17882 (N_17882,N_16293,N_16715);
or U17883 (N_17883,N_16170,N_16970);
nand U17884 (N_17884,N_16571,N_16105);
nand U17885 (N_17885,N_16591,N_16724);
nand U17886 (N_17886,N_16764,N_16245);
nand U17887 (N_17887,N_16809,N_16108);
or U17888 (N_17888,N_16376,N_16992);
nor U17889 (N_17889,N_16298,N_16082);
nor U17890 (N_17890,N_16754,N_16852);
nor U17891 (N_17891,N_16456,N_16718);
and U17892 (N_17892,N_16843,N_16497);
nand U17893 (N_17893,N_16331,N_16368);
nand U17894 (N_17894,N_16214,N_16937);
nor U17895 (N_17895,N_16597,N_16215);
xnor U17896 (N_17896,N_16410,N_16612);
nand U17897 (N_17897,N_16078,N_16294);
nor U17898 (N_17898,N_16807,N_16554);
and U17899 (N_17899,N_16701,N_16859);
nand U17900 (N_17900,N_16286,N_16470);
or U17901 (N_17901,N_16644,N_16051);
or U17902 (N_17902,N_16595,N_16869);
and U17903 (N_17903,N_16646,N_16071);
xnor U17904 (N_17904,N_16450,N_16280);
and U17905 (N_17905,N_16729,N_16345);
or U17906 (N_17906,N_16983,N_16325);
and U17907 (N_17907,N_16023,N_16296);
nor U17908 (N_17908,N_16727,N_16782);
or U17909 (N_17909,N_16126,N_16681);
nand U17910 (N_17910,N_16265,N_16249);
or U17911 (N_17911,N_16933,N_16005);
xnor U17912 (N_17912,N_16339,N_16563);
or U17913 (N_17913,N_16016,N_16702);
or U17914 (N_17914,N_16956,N_16401);
and U17915 (N_17915,N_16677,N_16723);
and U17916 (N_17916,N_16458,N_16776);
or U17917 (N_17917,N_16998,N_16868);
nor U17918 (N_17918,N_16181,N_16029);
nand U17919 (N_17919,N_16380,N_16252);
nand U17920 (N_17920,N_16708,N_16010);
nor U17921 (N_17921,N_16355,N_16390);
nand U17922 (N_17922,N_16558,N_16377);
nor U17923 (N_17923,N_16631,N_16679);
nand U17924 (N_17924,N_16697,N_16288);
or U17925 (N_17925,N_16443,N_16991);
nor U17926 (N_17926,N_16500,N_16134);
nor U17927 (N_17927,N_16622,N_16401);
nor U17928 (N_17928,N_16658,N_16898);
nor U17929 (N_17929,N_16214,N_16505);
and U17930 (N_17930,N_16255,N_16034);
xnor U17931 (N_17931,N_16340,N_16148);
nor U17932 (N_17932,N_16685,N_16599);
xor U17933 (N_17933,N_16244,N_16915);
nand U17934 (N_17934,N_16483,N_16064);
or U17935 (N_17935,N_16993,N_16882);
nor U17936 (N_17936,N_16511,N_16971);
nor U17937 (N_17937,N_16739,N_16515);
and U17938 (N_17938,N_16015,N_16800);
or U17939 (N_17939,N_16270,N_16450);
or U17940 (N_17940,N_16858,N_16458);
nor U17941 (N_17941,N_16259,N_16434);
or U17942 (N_17942,N_16823,N_16153);
nand U17943 (N_17943,N_16939,N_16278);
and U17944 (N_17944,N_16751,N_16703);
or U17945 (N_17945,N_16518,N_16338);
or U17946 (N_17946,N_16597,N_16490);
xnor U17947 (N_17947,N_16170,N_16426);
or U17948 (N_17948,N_16951,N_16415);
or U17949 (N_17949,N_16148,N_16719);
nor U17950 (N_17950,N_16713,N_16126);
nor U17951 (N_17951,N_16664,N_16420);
or U17952 (N_17952,N_16831,N_16498);
or U17953 (N_17953,N_16116,N_16995);
xnor U17954 (N_17954,N_16950,N_16863);
nand U17955 (N_17955,N_16297,N_16461);
and U17956 (N_17956,N_16446,N_16481);
nand U17957 (N_17957,N_16314,N_16039);
or U17958 (N_17958,N_16766,N_16882);
and U17959 (N_17959,N_16361,N_16591);
nand U17960 (N_17960,N_16722,N_16387);
nand U17961 (N_17961,N_16097,N_16191);
and U17962 (N_17962,N_16302,N_16674);
xor U17963 (N_17963,N_16719,N_16160);
nand U17964 (N_17964,N_16531,N_16301);
or U17965 (N_17965,N_16920,N_16311);
and U17966 (N_17966,N_16586,N_16648);
nor U17967 (N_17967,N_16299,N_16922);
xnor U17968 (N_17968,N_16535,N_16957);
nand U17969 (N_17969,N_16761,N_16035);
nand U17970 (N_17970,N_16861,N_16897);
or U17971 (N_17971,N_16140,N_16837);
nand U17972 (N_17972,N_16130,N_16977);
nor U17973 (N_17973,N_16220,N_16585);
or U17974 (N_17974,N_16914,N_16909);
nor U17975 (N_17975,N_16759,N_16806);
nor U17976 (N_17976,N_16601,N_16992);
nor U17977 (N_17977,N_16592,N_16578);
xor U17978 (N_17978,N_16924,N_16060);
nand U17979 (N_17979,N_16799,N_16376);
and U17980 (N_17980,N_16223,N_16630);
xnor U17981 (N_17981,N_16862,N_16429);
nand U17982 (N_17982,N_16636,N_16118);
nor U17983 (N_17983,N_16586,N_16470);
xor U17984 (N_17984,N_16508,N_16764);
nor U17985 (N_17985,N_16387,N_16854);
nand U17986 (N_17986,N_16759,N_16674);
nor U17987 (N_17987,N_16911,N_16785);
or U17988 (N_17988,N_16645,N_16404);
and U17989 (N_17989,N_16989,N_16708);
and U17990 (N_17990,N_16734,N_16469);
or U17991 (N_17991,N_16134,N_16081);
nor U17992 (N_17992,N_16534,N_16626);
nor U17993 (N_17993,N_16936,N_16505);
xor U17994 (N_17994,N_16845,N_16339);
xor U17995 (N_17995,N_16927,N_16503);
nor U17996 (N_17996,N_16573,N_16333);
and U17997 (N_17997,N_16761,N_16696);
nand U17998 (N_17998,N_16369,N_16964);
nor U17999 (N_17999,N_16271,N_16982);
nor U18000 (N_18000,N_17838,N_17368);
nand U18001 (N_18001,N_17090,N_17162);
and U18002 (N_18002,N_17187,N_17289);
or U18003 (N_18003,N_17207,N_17278);
or U18004 (N_18004,N_17038,N_17412);
and U18005 (N_18005,N_17859,N_17301);
or U18006 (N_18006,N_17843,N_17102);
nand U18007 (N_18007,N_17883,N_17803);
or U18008 (N_18008,N_17664,N_17758);
xor U18009 (N_18009,N_17250,N_17672);
and U18010 (N_18010,N_17435,N_17612);
and U18011 (N_18011,N_17510,N_17668);
nor U18012 (N_18012,N_17127,N_17957);
xor U18013 (N_18013,N_17943,N_17600);
nand U18014 (N_18014,N_17543,N_17697);
and U18015 (N_18015,N_17736,N_17534);
or U18016 (N_18016,N_17946,N_17969);
or U18017 (N_18017,N_17202,N_17133);
nand U18018 (N_18018,N_17780,N_17474);
xor U18019 (N_18019,N_17495,N_17635);
nor U18020 (N_18020,N_17651,N_17243);
nor U18021 (N_18021,N_17784,N_17869);
and U18022 (N_18022,N_17523,N_17363);
nand U18023 (N_18023,N_17271,N_17332);
nand U18024 (N_18024,N_17824,N_17912);
or U18025 (N_18025,N_17342,N_17813);
nor U18026 (N_18026,N_17210,N_17568);
nand U18027 (N_18027,N_17227,N_17837);
or U18028 (N_18028,N_17190,N_17654);
nor U18029 (N_18029,N_17005,N_17361);
nor U18030 (N_18030,N_17681,N_17279);
nand U18031 (N_18031,N_17918,N_17825);
nand U18032 (N_18032,N_17045,N_17414);
or U18033 (N_18033,N_17872,N_17965);
or U18034 (N_18034,N_17461,N_17839);
and U18035 (N_18035,N_17639,N_17975);
nor U18036 (N_18036,N_17625,N_17198);
nor U18037 (N_18037,N_17298,N_17076);
and U18038 (N_18038,N_17172,N_17742);
nand U18039 (N_18039,N_17015,N_17094);
and U18040 (N_18040,N_17092,N_17194);
or U18041 (N_18041,N_17911,N_17739);
nand U18042 (N_18042,N_17083,N_17772);
xnor U18043 (N_18043,N_17862,N_17307);
nor U18044 (N_18044,N_17616,N_17046);
or U18045 (N_18045,N_17677,N_17136);
nand U18046 (N_18046,N_17032,N_17470);
or U18047 (N_18047,N_17445,N_17456);
nand U18048 (N_18048,N_17857,N_17966);
nand U18049 (N_18049,N_17426,N_17258);
nor U18050 (N_18050,N_17521,N_17955);
and U18051 (N_18051,N_17561,N_17177);
nand U18052 (N_18052,N_17844,N_17188);
nand U18053 (N_18053,N_17261,N_17611);
or U18054 (N_18054,N_17774,N_17499);
nand U18055 (N_18055,N_17346,N_17787);
nor U18056 (N_18056,N_17373,N_17021);
or U18057 (N_18057,N_17782,N_17374);
xnor U18058 (N_18058,N_17558,N_17218);
nor U18059 (N_18059,N_17444,N_17476);
nand U18060 (N_18060,N_17904,N_17998);
or U18061 (N_18061,N_17204,N_17880);
nor U18062 (N_18062,N_17593,N_17648);
or U18063 (N_18063,N_17786,N_17330);
and U18064 (N_18064,N_17276,N_17728);
nand U18065 (N_18065,N_17179,N_17108);
nand U18066 (N_18066,N_17566,N_17466);
nand U18067 (N_18067,N_17981,N_17410);
and U18068 (N_18068,N_17900,N_17356);
nor U18069 (N_18069,N_17737,N_17832);
or U18070 (N_18070,N_17684,N_17638);
or U18071 (N_18071,N_17422,N_17846);
xnor U18072 (N_18072,N_17240,N_17026);
and U18073 (N_18073,N_17120,N_17686);
nor U18074 (N_18074,N_17798,N_17174);
nand U18075 (N_18075,N_17115,N_17746);
nor U18076 (N_18076,N_17365,N_17529);
nand U18077 (N_18077,N_17173,N_17425);
and U18078 (N_18078,N_17603,N_17820);
nor U18079 (N_18079,N_17488,N_17691);
nor U18080 (N_18080,N_17889,N_17449);
nand U18081 (N_18081,N_17496,N_17808);
xnor U18082 (N_18082,N_17216,N_17448);
nor U18083 (N_18083,N_17548,N_17049);
nand U18084 (N_18084,N_17637,N_17500);
nor U18085 (N_18085,N_17709,N_17554);
and U18086 (N_18086,N_17641,N_17819);
xnor U18087 (N_18087,N_17376,N_17123);
and U18088 (N_18088,N_17084,N_17321);
and U18089 (N_18089,N_17805,N_17674);
or U18090 (N_18090,N_17164,N_17489);
xnor U18091 (N_18091,N_17415,N_17753);
nor U18092 (N_18092,N_17086,N_17687);
or U18093 (N_18093,N_17947,N_17138);
or U18094 (N_18094,N_17799,N_17956);
and U18095 (N_18095,N_17621,N_17704);
nor U18096 (N_18096,N_17925,N_17852);
or U18097 (N_18097,N_17427,N_17296);
and U18098 (N_18098,N_17436,N_17926);
nor U18099 (N_18099,N_17631,N_17159);
nor U18100 (N_18100,N_17882,N_17605);
xor U18101 (N_18101,N_17696,N_17260);
nand U18102 (N_18102,N_17773,N_17310);
and U18103 (N_18103,N_17357,N_17088);
and U18104 (N_18104,N_17973,N_17506);
nor U18105 (N_18105,N_17486,N_17362);
or U18106 (N_18106,N_17682,N_17785);
and U18107 (N_18107,N_17100,N_17952);
nand U18108 (N_18108,N_17482,N_17297);
xor U18109 (N_18109,N_17281,N_17991);
nand U18110 (N_18110,N_17724,N_17581);
and U18111 (N_18111,N_17630,N_17735);
and U18112 (N_18112,N_17884,N_17740);
nor U18113 (N_18113,N_17795,N_17520);
nand U18114 (N_18114,N_17669,N_17339);
xor U18115 (N_18115,N_17041,N_17788);
nor U18116 (N_18116,N_17666,N_17033);
nand U18117 (N_18117,N_17228,N_17160);
or U18118 (N_18118,N_17155,N_17552);
xnor U18119 (N_18119,N_17077,N_17822);
and U18120 (N_18120,N_17318,N_17231);
nor U18121 (N_18121,N_17923,N_17472);
nand U18122 (N_18122,N_17781,N_17665);
or U18123 (N_18123,N_17615,N_17526);
and U18124 (N_18124,N_17917,N_17713);
nor U18125 (N_18125,N_17024,N_17014);
nor U18126 (N_18126,N_17814,N_17420);
nand U18127 (N_18127,N_17576,N_17383);
nor U18128 (N_18128,N_17986,N_17269);
nand U18129 (N_18129,N_17096,N_17934);
and U18130 (N_18130,N_17875,N_17961);
and U18131 (N_18131,N_17056,N_17176);
and U18132 (N_18132,N_17892,N_17438);
and U18133 (N_18133,N_17633,N_17890);
nand U18134 (N_18134,N_17129,N_17055);
nor U18135 (N_18135,N_17070,N_17663);
nor U18136 (N_18136,N_17878,N_17165);
xor U18137 (N_18137,N_17256,N_17707);
or U18138 (N_18138,N_17241,N_17335);
or U18139 (N_18139,N_17430,N_17185);
xnor U18140 (N_18140,N_17545,N_17519);
nor U18141 (N_18141,N_17382,N_17268);
xor U18142 (N_18142,N_17416,N_17344);
nor U18143 (N_18143,N_17058,N_17804);
or U18144 (N_18144,N_17294,N_17932);
nor U18145 (N_18145,N_17478,N_17539);
nor U18146 (N_18146,N_17743,N_17895);
and U18147 (N_18147,N_17987,N_17602);
or U18148 (N_18148,N_17467,N_17492);
nand U18149 (N_18149,N_17891,N_17594);
and U18150 (N_18150,N_17652,N_17930);
nand U18151 (N_18151,N_17775,N_17992);
or U18152 (N_18152,N_17226,N_17508);
nand U18153 (N_18153,N_17182,N_17010);
nor U18154 (N_18154,N_17967,N_17481);
nand U18155 (N_18155,N_17469,N_17450);
nor U18156 (N_18156,N_17167,N_17777);
or U18157 (N_18157,N_17013,N_17395);
nand U18158 (N_18158,N_17797,N_17715);
and U18159 (N_18159,N_17954,N_17477);
or U18160 (N_18160,N_17976,N_17065);
nor U18161 (N_18161,N_17212,N_17407);
nor U18162 (N_18162,N_17902,N_17679);
or U18163 (N_18163,N_17812,N_17836);
nor U18164 (N_18164,N_17877,N_17371);
and U18165 (N_18165,N_17575,N_17587);
nand U18166 (N_18166,N_17752,N_17741);
nor U18167 (N_18167,N_17494,N_17675);
nor U18168 (N_18168,N_17985,N_17779);
or U18169 (N_18169,N_17285,N_17604);
and U18170 (N_18170,N_17656,N_17459);
and U18171 (N_18171,N_17348,N_17103);
xnor U18172 (N_18172,N_17263,N_17315);
nand U18173 (N_18173,N_17408,N_17390);
xnor U18174 (N_18174,N_17460,N_17984);
or U18175 (N_18175,N_17340,N_17091);
xor U18176 (N_18176,N_17234,N_17017);
or U18177 (N_18177,N_17380,N_17893);
nand U18178 (N_18178,N_17721,N_17860);
nand U18179 (N_18179,N_17711,N_17725);
nor U18180 (N_18180,N_17647,N_17560);
nor U18181 (N_18181,N_17706,N_17870);
nor U18182 (N_18182,N_17006,N_17072);
nor U18183 (N_18183,N_17002,N_17039);
and U18184 (N_18184,N_17366,N_17802);
or U18185 (N_18185,N_17044,N_17433);
nand U18186 (N_18186,N_17700,N_17744);
or U18187 (N_18187,N_17886,N_17452);
nand U18188 (N_18188,N_17053,N_17154);
and U18189 (N_18189,N_17131,N_17439);
nand U18190 (N_18190,N_17671,N_17104);
xor U18191 (N_18191,N_17359,N_17057);
or U18192 (N_18192,N_17827,N_17614);
nand U18193 (N_18193,N_17591,N_17040);
nand U18194 (N_18194,N_17480,N_17977);
nor U18195 (N_18195,N_17557,N_17874);
and U18196 (N_18196,N_17485,N_17559);
nor U18197 (N_18197,N_17280,N_17314);
nor U18198 (N_18198,N_17722,N_17640);
nand U18199 (N_18199,N_17491,N_17004);
nand U18200 (N_18200,N_17405,N_17059);
nor U18201 (N_18201,N_17451,N_17750);
or U18202 (N_18202,N_17936,N_17413);
xnor U18203 (N_18203,N_17302,N_17255);
nand U18204 (N_18204,N_17311,N_17290);
or U18205 (N_18205,N_17504,N_17484);
nand U18206 (N_18206,N_17191,N_17790);
nand U18207 (N_18207,N_17454,N_17765);
nor U18208 (N_18208,N_17673,N_17815);
or U18209 (N_18209,N_17791,N_17483);
or U18210 (N_18210,N_17397,N_17994);
and U18211 (N_18211,N_17751,N_17214);
and U18212 (N_18212,N_17453,N_17577);
and U18213 (N_18213,N_17338,N_17341);
nand U18214 (N_18214,N_17418,N_17437);
or U18215 (N_18215,N_17716,N_17622);
nor U18216 (N_18216,N_17888,N_17695);
and U18217 (N_18217,N_17379,N_17586);
or U18218 (N_18218,N_17308,N_17513);
nand U18219 (N_18219,N_17432,N_17121);
or U18220 (N_18220,N_17583,N_17939);
nand U18221 (N_18221,N_17446,N_17197);
nand U18222 (N_18222,N_17398,N_17749);
nand U18223 (N_18223,N_17035,N_17370);
or U18224 (N_18224,N_17292,N_17107);
or U18225 (N_18225,N_17745,N_17730);
nand U18226 (N_18226,N_17579,N_17219);
and U18227 (N_18227,N_17493,N_17331);
or U18228 (N_18228,N_17067,N_17109);
or U18229 (N_18229,N_17458,N_17336);
nor U18230 (N_18230,N_17702,N_17989);
nor U18231 (N_18231,N_17596,N_17016);
xor U18232 (N_18232,N_17205,N_17145);
nand U18233 (N_18233,N_17333,N_17606);
and U18234 (N_18234,N_17396,N_17885);
nand U18235 (N_18235,N_17941,N_17644);
nand U18236 (N_18236,N_17968,N_17209);
nor U18237 (N_18237,N_17146,N_17937);
and U18238 (N_18238,N_17649,N_17778);
xor U18239 (N_18239,N_17610,N_17897);
nor U18240 (N_18240,N_17367,N_17229);
and U18241 (N_18241,N_17019,N_17501);
and U18242 (N_18242,N_17254,N_17050);
nor U18243 (N_18243,N_17963,N_17854);
nor U18244 (N_18244,N_17312,N_17447);
and U18245 (N_18245,N_17497,N_17157);
xor U18246 (N_18246,N_17546,N_17719);
nand U18247 (N_18247,N_17211,N_17029);
nor U18248 (N_18248,N_17001,N_17238);
nor U18249 (N_18249,N_17747,N_17252);
nor U18250 (N_18250,N_17899,N_17817);
and U18251 (N_18251,N_17277,N_17512);
and U18252 (N_18252,N_17244,N_17617);
nor U18253 (N_18253,N_17689,N_17879);
nor U18254 (N_18254,N_17392,N_17848);
or U18255 (N_18255,N_17062,N_17514);
nand U18256 (N_18256,N_17144,N_17220);
or U18257 (N_18257,N_17525,N_17826);
or U18258 (N_18258,N_17248,N_17137);
and U18259 (N_18259,N_17200,N_17538);
nor U18260 (N_18260,N_17267,N_17284);
nand U18261 (N_18261,N_17221,N_17273);
nand U18262 (N_18262,N_17286,N_17364);
nor U18263 (N_18263,N_17087,N_17699);
nand U18264 (N_18264,N_17845,N_17921);
and U18265 (N_18265,N_17562,N_17518);
nor U18266 (N_18266,N_17463,N_17794);
nor U18267 (N_18267,N_17201,N_17502);
nor U18268 (N_18268,N_17999,N_17841);
or U18269 (N_18269,N_17511,N_17051);
xor U18270 (N_18270,N_17770,N_17468);
and U18271 (N_18271,N_17731,N_17208);
nor U18272 (N_18272,N_17022,N_17855);
nor U18273 (N_18273,N_17720,N_17385);
nor U18274 (N_18274,N_17871,N_17350);
nand U18275 (N_18275,N_17517,N_17515);
nand U18276 (N_18276,N_17487,N_17224);
or U18277 (N_18277,N_17712,N_17972);
nand U18278 (N_18278,N_17189,N_17345);
and U18279 (N_18279,N_17093,N_17178);
nor U18280 (N_18280,N_17597,N_17074);
and U18281 (N_18281,N_17233,N_17595);
nor U18282 (N_18282,N_17152,N_17849);
or U18283 (N_18283,N_17828,N_17266);
and U18284 (N_18284,N_17343,N_17949);
and U18285 (N_18285,N_17896,N_17317);
nor U18286 (N_18286,N_17599,N_17717);
nand U18287 (N_18287,N_17783,N_17553);
or U18288 (N_18288,N_17993,N_17983);
nand U18289 (N_18289,N_17295,N_17935);
nor U18290 (N_18290,N_17776,N_17873);
xnor U18291 (N_18291,N_17537,N_17628);
nand U18292 (N_18292,N_17106,N_17011);
nand U18293 (N_18293,N_17023,N_17360);
or U18294 (N_18294,N_17894,N_17111);
nor U18295 (N_18295,N_17223,N_17169);
and U18296 (N_18296,N_17215,N_17105);
nor U18297 (N_18297,N_17761,N_17660);
nor U18298 (N_18298,N_17662,N_17944);
nand U18299 (N_18299,N_17061,N_17908);
nor U18300 (N_18300,N_17764,N_17095);
nor U18301 (N_18301,N_17075,N_17037);
or U18302 (N_18302,N_17796,N_17222);
and U18303 (N_18303,N_17206,N_17126);
nand U18304 (N_18304,N_17288,N_17978);
or U18305 (N_18305,N_17726,N_17763);
and U18306 (N_18306,N_17320,N_17128);
or U18307 (N_18307,N_17801,N_17283);
and U18308 (N_18308,N_17655,N_17140);
nand U18309 (N_18309,N_17970,N_17465);
or U18310 (N_18310,N_17574,N_17116);
nor U18311 (N_18311,N_17582,N_17589);
xnor U18312 (N_18312,N_17809,N_17230);
and U18313 (N_18313,N_17000,N_17818);
nand U18314 (N_18314,N_17768,N_17962);
and U18315 (N_18315,N_17913,N_17275);
xor U18316 (N_18316,N_17851,N_17110);
or U18317 (N_18317,N_17555,N_17264);
xnor U18318 (N_18318,N_17516,N_17253);
nand U18319 (N_18319,N_17953,N_17052);
nand U18320 (N_18320,N_17195,N_17097);
or U18321 (N_18321,N_17247,N_17831);
or U18322 (N_18322,N_17262,N_17861);
and U18323 (N_18323,N_17082,N_17536);
nand U18324 (N_18324,N_17400,N_17471);
xor U18325 (N_18325,N_17570,N_17565);
nand U18326 (N_18326,N_17192,N_17306);
and U18327 (N_18327,N_17375,N_17945);
nand U18328 (N_18328,N_17161,N_17964);
and U18329 (N_18329,N_17239,N_17287);
xor U18330 (N_18330,N_17569,N_17729);
nand U18331 (N_18331,N_17353,N_17907);
nor U18332 (N_18332,N_17428,N_17112);
nand U18333 (N_18333,N_17592,N_17193);
nand U18334 (N_18334,N_17007,N_17847);
and U18335 (N_18335,N_17876,N_17354);
and U18336 (N_18336,N_17394,N_17982);
and U18337 (N_18337,N_17842,N_17071);
or U18338 (N_18338,N_17646,N_17585);
nand U18339 (N_18339,N_17149,N_17117);
and U18340 (N_18340,N_17319,N_17073);
nor U18341 (N_18341,N_17670,N_17355);
nand U18342 (N_18342,N_17503,N_17509);
or U18343 (N_18343,N_17718,N_17225);
and U18344 (N_18344,N_17830,N_17829);
nand U18345 (N_18345,N_17864,N_17031);
xor U18346 (N_18346,N_17170,N_17036);
xnor U18347 (N_18347,N_17018,N_17714);
nor U18348 (N_18348,N_17678,N_17997);
nor U18349 (N_18349,N_17924,N_17657);
and U18350 (N_18350,N_17246,N_17609);
or U18351 (N_18351,N_17431,N_17661);
xor U18352 (N_18352,N_17440,N_17835);
nand U18353 (N_18353,N_17156,N_17866);
and U18354 (N_18354,N_17800,N_17951);
or U18355 (N_18355,N_17667,N_17974);
or U18356 (N_18356,N_17676,N_17066);
nand U18357 (N_18357,N_17867,N_17078);
nor U18358 (N_18358,N_17399,N_17996);
and U18359 (N_18359,N_17940,N_17429);
and U18360 (N_18360,N_17748,N_17175);
xnor U18361 (N_18361,N_17910,N_17821);
xor U18362 (N_18362,N_17423,N_17386);
or U18363 (N_18363,N_17540,N_17524);
nand U18364 (N_18364,N_17358,N_17898);
or U18365 (N_18365,N_17384,N_17150);
nor U18366 (N_18366,N_17455,N_17650);
xor U18367 (N_18367,N_17645,N_17099);
or U18368 (N_18368,N_17980,N_17168);
nand U18369 (N_18369,N_17441,N_17337);
nor U18370 (N_18370,N_17323,N_17113);
and U18371 (N_18371,N_17530,N_17909);
nor U18372 (N_18372,N_17688,N_17535);
xor U18373 (N_18373,N_17950,N_17158);
or U18374 (N_18374,N_17634,N_17334);
nor U18375 (N_18375,N_17550,N_17098);
nor U18376 (N_18376,N_17629,N_17738);
nor U18377 (N_18377,N_17624,N_17556);
or U18378 (N_18378,N_17130,N_17409);
nand U18379 (N_18379,N_17235,N_17401);
xnor U18380 (N_18380,N_17213,N_17920);
nor U18381 (N_18381,N_17028,N_17328);
and U18382 (N_18382,N_17858,N_17300);
and U18383 (N_18383,N_17387,N_17755);
or U18384 (N_18384,N_17756,N_17403);
and U18385 (N_18385,N_17727,N_17598);
and U18386 (N_18386,N_17572,N_17995);
xnor U18387 (N_18387,N_17054,N_17089);
nand U18388 (N_18388,N_17642,N_17643);
nand U18389 (N_18389,N_17916,N_17305);
and U18390 (N_18390,N_17771,N_17723);
xor U18391 (N_18391,N_17148,N_17166);
or U18392 (N_18392,N_17404,N_17291);
or U18393 (N_18393,N_17085,N_17081);
nand U18394 (N_18394,N_17402,N_17064);
xnor U18395 (N_18395,N_17101,N_17759);
or U18396 (N_18396,N_17958,N_17443);
nand U18397 (N_18397,N_17601,N_17377);
xnor U18398 (N_18398,N_17959,N_17948);
nand U18399 (N_18399,N_17856,N_17479);
or U18400 (N_18400,N_17326,N_17457);
nor U18401 (N_18401,N_17806,N_17658);
and U18402 (N_18402,N_17544,N_17003);
and U18403 (N_18403,N_17047,N_17927);
xnor U18404 (N_18404,N_17203,N_17184);
nor U18405 (N_18405,N_17270,N_17025);
and U18406 (N_18406,N_17659,N_17034);
nor U18407 (N_18407,N_17887,N_17153);
and U18408 (N_18408,N_17690,N_17299);
or U18409 (N_18409,N_17464,N_17626);
or U18410 (N_18410,N_17417,N_17960);
nand U18411 (N_18411,N_17183,N_17701);
and U18412 (N_18412,N_17282,N_17623);
nand U18413 (N_18413,N_17079,N_17251);
and U18414 (N_18414,N_17351,N_17027);
or U18415 (N_18415,N_17698,N_17531);
nand U18416 (N_18416,N_17372,N_17807);
nand U18417 (N_18417,N_17922,N_17369);
nand U18418 (N_18418,N_17265,N_17551);
and U18419 (N_18419,N_17434,N_17063);
nand U18420 (N_18420,N_17473,N_17578);
nor U18421 (N_18421,N_17125,N_17309);
or U18422 (N_18422,N_17833,N_17680);
xnor U18423 (N_18423,N_17259,N_17619);
and U18424 (N_18424,N_17132,N_17030);
xnor U18425 (N_18425,N_17505,N_17733);
and U18426 (N_18426,N_17938,N_17442);
nand U18427 (N_18427,N_17919,N_17789);
and U18428 (N_18428,N_17590,N_17792);
or U18429 (N_18429,N_17840,N_17906);
or U18430 (N_18430,N_17710,N_17527);
and U18431 (N_18431,N_17541,N_17199);
nand U18432 (N_18432,N_17549,N_17012);
or U18433 (N_18433,N_17881,N_17547);
nor U18434 (N_18434,N_17048,N_17766);
or U18435 (N_18435,N_17462,N_17732);
nor U18436 (N_18436,N_17068,N_17901);
and U18437 (N_18437,N_17313,N_17942);
nor U18438 (N_18438,N_17119,N_17683);
nand U18439 (N_18439,N_17114,N_17060);
xor U18440 (N_18440,N_17734,N_17705);
nor U18441 (N_18441,N_17563,N_17141);
nor U18442 (N_18442,N_17171,N_17588);
nand U18443 (N_18443,N_17142,N_17135);
nand U18444 (N_18444,N_17694,N_17419);
nand U18445 (N_18445,N_17865,N_17971);
or U18446 (N_18446,N_17236,N_17388);
nand U18447 (N_18447,N_17834,N_17381);
xor U18448 (N_18448,N_17163,N_17542);
or U18449 (N_18449,N_17580,N_17424);
nand U18450 (N_18450,N_17522,N_17245);
xor U18451 (N_18451,N_17811,N_17378);
nor U18452 (N_18452,N_17043,N_17237);
nand U18453 (N_18453,N_17573,N_17122);
nor U18454 (N_18454,N_17124,N_17767);
nor U18455 (N_18455,N_17528,N_17931);
or U18456 (N_18456,N_17903,N_17393);
xnor U18457 (N_18457,N_17134,N_17863);
xor U18458 (N_18458,N_17069,N_17693);
or U18459 (N_18459,N_17653,N_17352);
nor U18460 (N_18460,N_17249,N_17272);
nand U18461 (N_18461,N_17754,N_17475);
and U18462 (N_18462,N_17349,N_17928);
nand U18463 (N_18463,N_17915,N_17143);
nor U18464 (N_18464,N_17685,N_17608);
nand U18465 (N_18465,N_17257,N_17914);
nor U18466 (N_18466,N_17868,N_17151);
xnor U18467 (N_18467,N_17632,N_17933);
nand U18468 (N_18468,N_17533,N_17181);
xor U18469 (N_18469,N_17316,N_17303);
nand U18470 (N_18470,N_17708,N_17929);
nor U18471 (N_18471,N_17327,N_17990);
or U18472 (N_18472,N_17760,N_17020);
nor U18473 (N_18473,N_17325,N_17080);
and U18474 (N_18474,N_17905,N_17490);
or U18475 (N_18475,N_17180,N_17988);
nand U18476 (N_18476,N_17567,N_17322);
and U18477 (N_18477,N_17274,N_17498);
and U18478 (N_18478,N_17324,N_17584);
nor U18479 (N_18479,N_17147,N_17692);
xnor U18480 (N_18480,N_17703,N_17620);
and U18481 (N_18481,N_17816,N_17008);
and U18482 (N_18482,N_17391,N_17564);
nor U18483 (N_18483,N_17532,N_17853);
nor U18484 (N_18484,N_17823,N_17636);
nor U18485 (N_18485,N_17139,N_17406);
and U18486 (N_18486,N_17186,N_17347);
and U18487 (N_18487,N_17769,N_17232);
xnor U18488 (N_18488,N_17507,N_17762);
nand U18489 (N_18489,N_17571,N_17389);
nand U18490 (N_18490,N_17217,N_17850);
nand U18491 (N_18491,N_17118,N_17793);
nand U18492 (N_18492,N_17042,N_17618);
nor U18493 (N_18493,N_17196,N_17242);
nor U18494 (N_18494,N_17613,N_17810);
nand U18495 (N_18495,N_17627,N_17009);
nor U18496 (N_18496,N_17411,N_17329);
and U18497 (N_18497,N_17421,N_17293);
or U18498 (N_18498,N_17757,N_17304);
nand U18499 (N_18499,N_17979,N_17607);
or U18500 (N_18500,N_17126,N_17395);
or U18501 (N_18501,N_17087,N_17041);
nand U18502 (N_18502,N_17380,N_17063);
or U18503 (N_18503,N_17595,N_17009);
or U18504 (N_18504,N_17454,N_17452);
nor U18505 (N_18505,N_17446,N_17646);
and U18506 (N_18506,N_17906,N_17913);
or U18507 (N_18507,N_17911,N_17555);
and U18508 (N_18508,N_17400,N_17171);
nand U18509 (N_18509,N_17928,N_17996);
nor U18510 (N_18510,N_17449,N_17612);
nand U18511 (N_18511,N_17911,N_17458);
or U18512 (N_18512,N_17257,N_17674);
or U18513 (N_18513,N_17488,N_17739);
nor U18514 (N_18514,N_17232,N_17979);
nand U18515 (N_18515,N_17707,N_17135);
nand U18516 (N_18516,N_17471,N_17016);
xor U18517 (N_18517,N_17934,N_17297);
and U18518 (N_18518,N_17571,N_17319);
nor U18519 (N_18519,N_17406,N_17431);
or U18520 (N_18520,N_17768,N_17953);
or U18521 (N_18521,N_17591,N_17032);
nor U18522 (N_18522,N_17324,N_17634);
nor U18523 (N_18523,N_17921,N_17991);
nor U18524 (N_18524,N_17207,N_17461);
nor U18525 (N_18525,N_17551,N_17919);
or U18526 (N_18526,N_17818,N_17853);
and U18527 (N_18527,N_17991,N_17071);
nor U18528 (N_18528,N_17634,N_17392);
nand U18529 (N_18529,N_17523,N_17994);
nor U18530 (N_18530,N_17527,N_17711);
nor U18531 (N_18531,N_17257,N_17258);
or U18532 (N_18532,N_17216,N_17710);
xnor U18533 (N_18533,N_17634,N_17858);
or U18534 (N_18534,N_17213,N_17718);
and U18535 (N_18535,N_17940,N_17140);
nor U18536 (N_18536,N_17153,N_17737);
or U18537 (N_18537,N_17888,N_17095);
nand U18538 (N_18538,N_17722,N_17009);
or U18539 (N_18539,N_17218,N_17844);
xor U18540 (N_18540,N_17182,N_17193);
or U18541 (N_18541,N_17142,N_17000);
or U18542 (N_18542,N_17376,N_17481);
or U18543 (N_18543,N_17098,N_17595);
nor U18544 (N_18544,N_17680,N_17203);
nand U18545 (N_18545,N_17968,N_17874);
and U18546 (N_18546,N_17288,N_17121);
and U18547 (N_18547,N_17566,N_17775);
nor U18548 (N_18548,N_17176,N_17168);
nand U18549 (N_18549,N_17077,N_17657);
and U18550 (N_18550,N_17143,N_17670);
nor U18551 (N_18551,N_17224,N_17881);
and U18552 (N_18552,N_17385,N_17278);
xor U18553 (N_18553,N_17903,N_17368);
nor U18554 (N_18554,N_17910,N_17680);
and U18555 (N_18555,N_17193,N_17626);
or U18556 (N_18556,N_17167,N_17879);
xor U18557 (N_18557,N_17696,N_17935);
nor U18558 (N_18558,N_17990,N_17127);
and U18559 (N_18559,N_17211,N_17395);
and U18560 (N_18560,N_17114,N_17994);
nand U18561 (N_18561,N_17029,N_17010);
and U18562 (N_18562,N_17252,N_17392);
or U18563 (N_18563,N_17219,N_17164);
nand U18564 (N_18564,N_17659,N_17276);
nor U18565 (N_18565,N_17667,N_17645);
nor U18566 (N_18566,N_17821,N_17837);
xnor U18567 (N_18567,N_17554,N_17818);
nand U18568 (N_18568,N_17037,N_17083);
or U18569 (N_18569,N_17390,N_17717);
nand U18570 (N_18570,N_17534,N_17935);
and U18571 (N_18571,N_17076,N_17504);
or U18572 (N_18572,N_17646,N_17374);
or U18573 (N_18573,N_17742,N_17954);
and U18574 (N_18574,N_17823,N_17084);
nor U18575 (N_18575,N_17135,N_17658);
xnor U18576 (N_18576,N_17745,N_17621);
or U18577 (N_18577,N_17165,N_17094);
nand U18578 (N_18578,N_17272,N_17823);
or U18579 (N_18579,N_17617,N_17877);
xnor U18580 (N_18580,N_17741,N_17570);
xor U18581 (N_18581,N_17145,N_17789);
nand U18582 (N_18582,N_17182,N_17616);
nor U18583 (N_18583,N_17576,N_17088);
nor U18584 (N_18584,N_17997,N_17338);
nand U18585 (N_18585,N_17028,N_17324);
and U18586 (N_18586,N_17971,N_17868);
and U18587 (N_18587,N_17161,N_17093);
nand U18588 (N_18588,N_17124,N_17995);
and U18589 (N_18589,N_17885,N_17502);
or U18590 (N_18590,N_17259,N_17871);
and U18591 (N_18591,N_17888,N_17472);
and U18592 (N_18592,N_17519,N_17689);
and U18593 (N_18593,N_17905,N_17302);
and U18594 (N_18594,N_17012,N_17090);
or U18595 (N_18595,N_17629,N_17013);
nand U18596 (N_18596,N_17777,N_17535);
or U18597 (N_18597,N_17982,N_17790);
and U18598 (N_18598,N_17917,N_17073);
nor U18599 (N_18599,N_17048,N_17841);
xor U18600 (N_18600,N_17491,N_17496);
and U18601 (N_18601,N_17210,N_17124);
and U18602 (N_18602,N_17100,N_17622);
nor U18603 (N_18603,N_17833,N_17568);
nor U18604 (N_18604,N_17817,N_17190);
xor U18605 (N_18605,N_17393,N_17878);
and U18606 (N_18606,N_17819,N_17941);
and U18607 (N_18607,N_17220,N_17539);
nor U18608 (N_18608,N_17894,N_17681);
or U18609 (N_18609,N_17301,N_17352);
or U18610 (N_18610,N_17017,N_17888);
and U18611 (N_18611,N_17605,N_17255);
and U18612 (N_18612,N_17166,N_17854);
nor U18613 (N_18613,N_17187,N_17796);
or U18614 (N_18614,N_17450,N_17396);
nor U18615 (N_18615,N_17308,N_17447);
nand U18616 (N_18616,N_17863,N_17275);
xnor U18617 (N_18617,N_17072,N_17079);
xor U18618 (N_18618,N_17163,N_17101);
nor U18619 (N_18619,N_17351,N_17618);
nor U18620 (N_18620,N_17810,N_17937);
or U18621 (N_18621,N_17122,N_17582);
and U18622 (N_18622,N_17014,N_17789);
and U18623 (N_18623,N_17938,N_17513);
or U18624 (N_18624,N_17686,N_17902);
nor U18625 (N_18625,N_17938,N_17916);
or U18626 (N_18626,N_17659,N_17095);
or U18627 (N_18627,N_17964,N_17621);
and U18628 (N_18628,N_17399,N_17454);
or U18629 (N_18629,N_17359,N_17096);
nand U18630 (N_18630,N_17498,N_17847);
and U18631 (N_18631,N_17021,N_17840);
nand U18632 (N_18632,N_17372,N_17287);
nor U18633 (N_18633,N_17372,N_17147);
or U18634 (N_18634,N_17355,N_17247);
and U18635 (N_18635,N_17482,N_17869);
nand U18636 (N_18636,N_17398,N_17532);
or U18637 (N_18637,N_17516,N_17156);
and U18638 (N_18638,N_17357,N_17225);
or U18639 (N_18639,N_17885,N_17813);
and U18640 (N_18640,N_17359,N_17630);
nand U18641 (N_18641,N_17727,N_17773);
nand U18642 (N_18642,N_17514,N_17280);
nor U18643 (N_18643,N_17331,N_17192);
or U18644 (N_18644,N_17142,N_17261);
nor U18645 (N_18645,N_17045,N_17039);
nand U18646 (N_18646,N_17903,N_17433);
and U18647 (N_18647,N_17794,N_17438);
nor U18648 (N_18648,N_17406,N_17287);
or U18649 (N_18649,N_17109,N_17202);
nor U18650 (N_18650,N_17020,N_17735);
nor U18651 (N_18651,N_17310,N_17096);
nand U18652 (N_18652,N_17811,N_17753);
nand U18653 (N_18653,N_17601,N_17028);
and U18654 (N_18654,N_17332,N_17214);
nand U18655 (N_18655,N_17019,N_17562);
and U18656 (N_18656,N_17296,N_17035);
nand U18657 (N_18657,N_17694,N_17073);
xnor U18658 (N_18658,N_17578,N_17960);
or U18659 (N_18659,N_17279,N_17854);
or U18660 (N_18660,N_17193,N_17538);
nand U18661 (N_18661,N_17052,N_17989);
xor U18662 (N_18662,N_17156,N_17095);
and U18663 (N_18663,N_17871,N_17656);
nand U18664 (N_18664,N_17727,N_17319);
nor U18665 (N_18665,N_17513,N_17199);
nor U18666 (N_18666,N_17900,N_17146);
nor U18667 (N_18667,N_17726,N_17718);
nand U18668 (N_18668,N_17724,N_17175);
nor U18669 (N_18669,N_17640,N_17483);
or U18670 (N_18670,N_17897,N_17047);
nand U18671 (N_18671,N_17821,N_17893);
nand U18672 (N_18672,N_17054,N_17968);
nor U18673 (N_18673,N_17203,N_17884);
nor U18674 (N_18674,N_17173,N_17591);
and U18675 (N_18675,N_17286,N_17723);
nor U18676 (N_18676,N_17977,N_17426);
nand U18677 (N_18677,N_17462,N_17077);
nor U18678 (N_18678,N_17223,N_17963);
nand U18679 (N_18679,N_17232,N_17013);
or U18680 (N_18680,N_17625,N_17213);
or U18681 (N_18681,N_17987,N_17834);
nor U18682 (N_18682,N_17576,N_17434);
nand U18683 (N_18683,N_17582,N_17236);
and U18684 (N_18684,N_17117,N_17550);
or U18685 (N_18685,N_17566,N_17331);
nor U18686 (N_18686,N_17186,N_17494);
nand U18687 (N_18687,N_17436,N_17405);
and U18688 (N_18688,N_17439,N_17305);
nand U18689 (N_18689,N_17492,N_17136);
xor U18690 (N_18690,N_17212,N_17959);
and U18691 (N_18691,N_17019,N_17461);
nand U18692 (N_18692,N_17295,N_17006);
xnor U18693 (N_18693,N_17031,N_17190);
xor U18694 (N_18694,N_17798,N_17287);
and U18695 (N_18695,N_17765,N_17939);
nand U18696 (N_18696,N_17890,N_17577);
nor U18697 (N_18697,N_17098,N_17603);
and U18698 (N_18698,N_17034,N_17161);
nor U18699 (N_18699,N_17316,N_17107);
xor U18700 (N_18700,N_17242,N_17529);
nand U18701 (N_18701,N_17337,N_17393);
nor U18702 (N_18702,N_17661,N_17829);
and U18703 (N_18703,N_17374,N_17825);
and U18704 (N_18704,N_17188,N_17249);
nor U18705 (N_18705,N_17839,N_17252);
nand U18706 (N_18706,N_17556,N_17912);
and U18707 (N_18707,N_17849,N_17218);
and U18708 (N_18708,N_17892,N_17052);
nor U18709 (N_18709,N_17279,N_17668);
nor U18710 (N_18710,N_17126,N_17907);
nor U18711 (N_18711,N_17565,N_17933);
nor U18712 (N_18712,N_17722,N_17882);
nor U18713 (N_18713,N_17020,N_17181);
or U18714 (N_18714,N_17292,N_17168);
xor U18715 (N_18715,N_17360,N_17488);
nand U18716 (N_18716,N_17135,N_17387);
xnor U18717 (N_18717,N_17871,N_17433);
nand U18718 (N_18718,N_17120,N_17371);
or U18719 (N_18719,N_17706,N_17327);
and U18720 (N_18720,N_17312,N_17402);
and U18721 (N_18721,N_17750,N_17870);
xor U18722 (N_18722,N_17435,N_17775);
or U18723 (N_18723,N_17946,N_17038);
and U18724 (N_18724,N_17427,N_17318);
and U18725 (N_18725,N_17701,N_17137);
nor U18726 (N_18726,N_17161,N_17019);
xnor U18727 (N_18727,N_17914,N_17527);
nor U18728 (N_18728,N_17212,N_17285);
xnor U18729 (N_18729,N_17485,N_17306);
or U18730 (N_18730,N_17614,N_17658);
nand U18731 (N_18731,N_17833,N_17519);
nand U18732 (N_18732,N_17697,N_17744);
nor U18733 (N_18733,N_17099,N_17130);
nor U18734 (N_18734,N_17190,N_17990);
or U18735 (N_18735,N_17551,N_17134);
nor U18736 (N_18736,N_17867,N_17331);
nor U18737 (N_18737,N_17430,N_17540);
xor U18738 (N_18738,N_17473,N_17821);
nor U18739 (N_18739,N_17901,N_17830);
or U18740 (N_18740,N_17376,N_17877);
nor U18741 (N_18741,N_17048,N_17847);
nor U18742 (N_18742,N_17519,N_17524);
and U18743 (N_18743,N_17899,N_17009);
nor U18744 (N_18744,N_17498,N_17148);
nand U18745 (N_18745,N_17080,N_17104);
xnor U18746 (N_18746,N_17697,N_17387);
or U18747 (N_18747,N_17334,N_17438);
or U18748 (N_18748,N_17917,N_17351);
nand U18749 (N_18749,N_17033,N_17598);
and U18750 (N_18750,N_17713,N_17653);
or U18751 (N_18751,N_17998,N_17934);
xnor U18752 (N_18752,N_17637,N_17378);
or U18753 (N_18753,N_17512,N_17057);
nor U18754 (N_18754,N_17966,N_17457);
nand U18755 (N_18755,N_17021,N_17249);
nand U18756 (N_18756,N_17876,N_17941);
nor U18757 (N_18757,N_17563,N_17946);
nand U18758 (N_18758,N_17388,N_17263);
and U18759 (N_18759,N_17559,N_17049);
and U18760 (N_18760,N_17686,N_17708);
and U18761 (N_18761,N_17101,N_17036);
and U18762 (N_18762,N_17361,N_17508);
nor U18763 (N_18763,N_17169,N_17115);
nor U18764 (N_18764,N_17803,N_17729);
nor U18765 (N_18765,N_17414,N_17987);
nor U18766 (N_18766,N_17905,N_17716);
nand U18767 (N_18767,N_17561,N_17095);
xor U18768 (N_18768,N_17348,N_17504);
and U18769 (N_18769,N_17263,N_17981);
nor U18770 (N_18770,N_17686,N_17405);
and U18771 (N_18771,N_17737,N_17802);
nand U18772 (N_18772,N_17408,N_17000);
nor U18773 (N_18773,N_17625,N_17654);
and U18774 (N_18774,N_17227,N_17292);
nand U18775 (N_18775,N_17043,N_17345);
nor U18776 (N_18776,N_17068,N_17762);
xor U18777 (N_18777,N_17041,N_17035);
nand U18778 (N_18778,N_17155,N_17685);
and U18779 (N_18779,N_17282,N_17577);
nand U18780 (N_18780,N_17857,N_17233);
nor U18781 (N_18781,N_17256,N_17757);
or U18782 (N_18782,N_17338,N_17450);
and U18783 (N_18783,N_17720,N_17372);
nand U18784 (N_18784,N_17247,N_17281);
nand U18785 (N_18785,N_17875,N_17993);
and U18786 (N_18786,N_17534,N_17881);
nand U18787 (N_18787,N_17483,N_17002);
nor U18788 (N_18788,N_17880,N_17750);
nand U18789 (N_18789,N_17648,N_17760);
and U18790 (N_18790,N_17225,N_17801);
and U18791 (N_18791,N_17906,N_17584);
nor U18792 (N_18792,N_17408,N_17119);
or U18793 (N_18793,N_17583,N_17859);
nor U18794 (N_18794,N_17606,N_17231);
nand U18795 (N_18795,N_17202,N_17825);
nor U18796 (N_18796,N_17730,N_17226);
and U18797 (N_18797,N_17070,N_17664);
nor U18798 (N_18798,N_17540,N_17299);
nand U18799 (N_18799,N_17190,N_17531);
nor U18800 (N_18800,N_17749,N_17719);
or U18801 (N_18801,N_17416,N_17678);
and U18802 (N_18802,N_17609,N_17318);
and U18803 (N_18803,N_17318,N_17887);
nor U18804 (N_18804,N_17715,N_17871);
nor U18805 (N_18805,N_17854,N_17410);
nand U18806 (N_18806,N_17865,N_17793);
xor U18807 (N_18807,N_17575,N_17551);
nor U18808 (N_18808,N_17277,N_17879);
nand U18809 (N_18809,N_17483,N_17115);
and U18810 (N_18810,N_17204,N_17652);
nor U18811 (N_18811,N_17088,N_17514);
nand U18812 (N_18812,N_17824,N_17485);
nor U18813 (N_18813,N_17451,N_17025);
xor U18814 (N_18814,N_17310,N_17816);
and U18815 (N_18815,N_17753,N_17258);
xor U18816 (N_18816,N_17480,N_17296);
and U18817 (N_18817,N_17040,N_17569);
or U18818 (N_18818,N_17123,N_17002);
or U18819 (N_18819,N_17305,N_17172);
xnor U18820 (N_18820,N_17760,N_17174);
nor U18821 (N_18821,N_17343,N_17392);
and U18822 (N_18822,N_17609,N_17647);
nor U18823 (N_18823,N_17500,N_17093);
and U18824 (N_18824,N_17620,N_17181);
or U18825 (N_18825,N_17298,N_17131);
or U18826 (N_18826,N_17756,N_17647);
xor U18827 (N_18827,N_17802,N_17371);
xnor U18828 (N_18828,N_17468,N_17159);
or U18829 (N_18829,N_17910,N_17646);
nor U18830 (N_18830,N_17863,N_17729);
and U18831 (N_18831,N_17549,N_17478);
or U18832 (N_18832,N_17606,N_17817);
and U18833 (N_18833,N_17924,N_17881);
and U18834 (N_18834,N_17160,N_17079);
or U18835 (N_18835,N_17493,N_17439);
and U18836 (N_18836,N_17983,N_17953);
nand U18837 (N_18837,N_17685,N_17141);
or U18838 (N_18838,N_17015,N_17342);
nor U18839 (N_18839,N_17452,N_17720);
nor U18840 (N_18840,N_17612,N_17671);
nor U18841 (N_18841,N_17374,N_17387);
nor U18842 (N_18842,N_17571,N_17934);
nand U18843 (N_18843,N_17651,N_17492);
nand U18844 (N_18844,N_17580,N_17896);
nor U18845 (N_18845,N_17691,N_17983);
or U18846 (N_18846,N_17580,N_17076);
nand U18847 (N_18847,N_17350,N_17031);
and U18848 (N_18848,N_17172,N_17778);
and U18849 (N_18849,N_17601,N_17878);
nor U18850 (N_18850,N_17586,N_17290);
nor U18851 (N_18851,N_17917,N_17360);
xor U18852 (N_18852,N_17831,N_17823);
or U18853 (N_18853,N_17246,N_17120);
nor U18854 (N_18854,N_17575,N_17056);
nor U18855 (N_18855,N_17553,N_17373);
or U18856 (N_18856,N_17995,N_17415);
and U18857 (N_18857,N_17605,N_17316);
nor U18858 (N_18858,N_17690,N_17116);
and U18859 (N_18859,N_17785,N_17014);
or U18860 (N_18860,N_17863,N_17853);
nor U18861 (N_18861,N_17945,N_17468);
xor U18862 (N_18862,N_17415,N_17862);
nand U18863 (N_18863,N_17565,N_17076);
and U18864 (N_18864,N_17337,N_17182);
nand U18865 (N_18865,N_17455,N_17250);
or U18866 (N_18866,N_17840,N_17641);
or U18867 (N_18867,N_17021,N_17391);
nand U18868 (N_18868,N_17284,N_17521);
and U18869 (N_18869,N_17995,N_17380);
nand U18870 (N_18870,N_17831,N_17431);
and U18871 (N_18871,N_17639,N_17790);
nor U18872 (N_18872,N_17867,N_17241);
and U18873 (N_18873,N_17798,N_17312);
nor U18874 (N_18874,N_17530,N_17916);
nor U18875 (N_18875,N_17838,N_17601);
and U18876 (N_18876,N_17044,N_17741);
or U18877 (N_18877,N_17151,N_17703);
nand U18878 (N_18878,N_17813,N_17551);
nor U18879 (N_18879,N_17874,N_17957);
nor U18880 (N_18880,N_17813,N_17072);
nor U18881 (N_18881,N_17217,N_17139);
or U18882 (N_18882,N_17354,N_17318);
nand U18883 (N_18883,N_17715,N_17018);
and U18884 (N_18884,N_17134,N_17480);
and U18885 (N_18885,N_17621,N_17695);
nand U18886 (N_18886,N_17580,N_17510);
nand U18887 (N_18887,N_17580,N_17933);
xor U18888 (N_18888,N_17923,N_17545);
and U18889 (N_18889,N_17495,N_17704);
nand U18890 (N_18890,N_17189,N_17503);
nand U18891 (N_18891,N_17367,N_17089);
and U18892 (N_18892,N_17512,N_17638);
xor U18893 (N_18893,N_17494,N_17821);
nand U18894 (N_18894,N_17643,N_17401);
nor U18895 (N_18895,N_17309,N_17200);
nor U18896 (N_18896,N_17517,N_17957);
or U18897 (N_18897,N_17218,N_17655);
xnor U18898 (N_18898,N_17975,N_17099);
nand U18899 (N_18899,N_17749,N_17771);
nor U18900 (N_18900,N_17046,N_17818);
and U18901 (N_18901,N_17328,N_17865);
or U18902 (N_18902,N_17496,N_17660);
nor U18903 (N_18903,N_17580,N_17984);
and U18904 (N_18904,N_17040,N_17249);
and U18905 (N_18905,N_17518,N_17793);
or U18906 (N_18906,N_17400,N_17851);
nand U18907 (N_18907,N_17436,N_17365);
xor U18908 (N_18908,N_17325,N_17153);
nor U18909 (N_18909,N_17518,N_17835);
nor U18910 (N_18910,N_17233,N_17214);
and U18911 (N_18911,N_17979,N_17778);
xor U18912 (N_18912,N_17072,N_17647);
or U18913 (N_18913,N_17944,N_17329);
and U18914 (N_18914,N_17577,N_17377);
and U18915 (N_18915,N_17126,N_17555);
nor U18916 (N_18916,N_17513,N_17329);
or U18917 (N_18917,N_17207,N_17748);
nor U18918 (N_18918,N_17680,N_17219);
nand U18919 (N_18919,N_17854,N_17817);
or U18920 (N_18920,N_17693,N_17959);
nand U18921 (N_18921,N_17652,N_17535);
or U18922 (N_18922,N_17372,N_17117);
and U18923 (N_18923,N_17450,N_17918);
nor U18924 (N_18924,N_17479,N_17259);
and U18925 (N_18925,N_17408,N_17810);
and U18926 (N_18926,N_17155,N_17636);
nor U18927 (N_18927,N_17486,N_17608);
nor U18928 (N_18928,N_17269,N_17526);
and U18929 (N_18929,N_17916,N_17517);
or U18930 (N_18930,N_17411,N_17430);
and U18931 (N_18931,N_17965,N_17251);
xor U18932 (N_18932,N_17106,N_17533);
and U18933 (N_18933,N_17148,N_17595);
and U18934 (N_18934,N_17350,N_17281);
xnor U18935 (N_18935,N_17078,N_17474);
nor U18936 (N_18936,N_17083,N_17884);
nor U18937 (N_18937,N_17190,N_17775);
nor U18938 (N_18938,N_17240,N_17548);
nand U18939 (N_18939,N_17927,N_17700);
nand U18940 (N_18940,N_17562,N_17807);
or U18941 (N_18941,N_17061,N_17687);
and U18942 (N_18942,N_17249,N_17956);
or U18943 (N_18943,N_17749,N_17534);
nand U18944 (N_18944,N_17926,N_17592);
or U18945 (N_18945,N_17283,N_17110);
xnor U18946 (N_18946,N_17237,N_17020);
xnor U18947 (N_18947,N_17368,N_17870);
nor U18948 (N_18948,N_17532,N_17830);
and U18949 (N_18949,N_17261,N_17467);
and U18950 (N_18950,N_17471,N_17946);
nor U18951 (N_18951,N_17952,N_17200);
nand U18952 (N_18952,N_17416,N_17205);
and U18953 (N_18953,N_17750,N_17281);
nor U18954 (N_18954,N_17044,N_17655);
or U18955 (N_18955,N_17747,N_17424);
nand U18956 (N_18956,N_17649,N_17350);
or U18957 (N_18957,N_17566,N_17752);
or U18958 (N_18958,N_17417,N_17496);
nor U18959 (N_18959,N_17118,N_17916);
nand U18960 (N_18960,N_17115,N_17790);
nor U18961 (N_18961,N_17055,N_17248);
nand U18962 (N_18962,N_17641,N_17209);
nor U18963 (N_18963,N_17416,N_17890);
and U18964 (N_18964,N_17794,N_17741);
or U18965 (N_18965,N_17871,N_17893);
or U18966 (N_18966,N_17721,N_17551);
and U18967 (N_18967,N_17335,N_17099);
nor U18968 (N_18968,N_17565,N_17126);
nor U18969 (N_18969,N_17540,N_17813);
or U18970 (N_18970,N_17601,N_17511);
nand U18971 (N_18971,N_17456,N_17968);
nor U18972 (N_18972,N_17475,N_17848);
nand U18973 (N_18973,N_17001,N_17090);
nor U18974 (N_18974,N_17703,N_17661);
or U18975 (N_18975,N_17951,N_17288);
and U18976 (N_18976,N_17811,N_17428);
or U18977 (N_18977,N_17725,N_17389);
nand U18978 (N_18978,N_17998,N_17337);
nor U18979 (N_18979,N_17692,N_17966);
nor U18980 (N_18980,N_17108,N_17203);
nor U18981 (N_18981,N_17390,N_17454);
xnor U18982 (N_18982,N_17300,N_17184);
nand U18983 (N_18983,N_17177,N_17151);
nor U18984 (N_18984,N_17527,N_17270);
and U18985 (N_18985,N_17081,N_17405);
or U18986 (N_18986,N_17802,N_17929);
or U18987 (N_18987,N_17585,N_17745);
nor U18988 (N_18988,N_17048,N_17006);
and U18989 (N_18989,N_17283,N_17472);
nand U18990 (N_18990,N_17432,N_17904);
and U18991 (N_18991,N_17428,N_17618);
and U18992 (N_18992,N_17863,N_17897);
nor U18993 (N_18993,N_17223,N_17609);
or U18994 (N_18994,N_17606,N_17084);
nor U18995 (N_18995,N_17517,N_17272);
nor U18996 (N_18996,N_17275,N_17745);
nor U18997 (N_18997,N_17988,N_17395);
or U18998 (N_18998,N_17225,N_17912);
and U18999 (N_18999,N_17182,N_17049);
or U19000 (N_19000,N_18458,N_18248);
nor U19001 (N_19001,N_18508,N_18745);
nand U19002 (N_19002,N_18700,N_18868);
nor U19003 (N_19003,N_18333,N_18402);
nor U19004 (N_19004,N_18223,N_18672);
nor U19005 (N_19005,N_18730,N_18072);
nand U19006 (N_19006,N_18470,N_18404);
nor U19007 (N_19007,N_18279,N_18069);
and U19008 (N_19008,N_18340,N_18909);
nand U19009 (N_19009,N_18557,N_18687);
or U19010 (N_19010,N_18294,N_18516);
xnor U19011 (N_19011,N_18242,N_18477);
nand U19012 (N_19012,N_18866,N_18990);
nor U19013 (N_19013,N_18750,N_18732);
nor U19014 (N_19014,N_18257,N_18350);
nand U19015 (N_19015,N_18618,N_18442);
and U19016 (N_19016,N_18729,N_18473);
and U19017 (N_19017,N_18252,N_18722);
nor U19018 (N_19018,N_18798,N_18727);
or U19019 (N_19019,N_18754,N_18101);
xor U19020 (N_19020,N_18921,N_18204);
nor U19021 (N_19021,N_18769,N_18879);
nand U19022 (N_19022,N_18147,N_18400);
nand U19023 (N_19023,N_18980,N_18770);
xor U19024 (N_19024,N_18758,N_18264);
xnor U19025 (N_19025,N_18523,N_18630);
or U19026 (N_19026,N_18092,N_18375);
xnor U19027 (N_19027,N_18940,N_18901);
and U19028 (N_19028,N_18873,N_18551);
xnor U19029 (N_19029,N_18033,N_18341);
nand U19030 (N_19030,N_18456,N_18309);
nor U19031 (N_19031,N_18927,N_18225);
nand U19032 (N_19032,N_18002,N_18032);
nor U19033 (N_19033,N_18850,N_18144);
nand U19034 (N_19034,N_18426,N_18148);
or U19035 (N_19035,N_18747,N_18505);
nor U19036 (N_19036,N_18411,N_18718);
nand U19037 (N_19037,N_18467,N_18075);
or U19038 (N_19038,N_18638,N_18544);
xnor U19039 (N_19039,N_18414,N_18027);
and U19040 (N_19040,N_18555,N_18013);
or U19041 (N_19041,N_18418,N_18760);
or U19042 (N_19042,N_18399,N_18303);
and U19043 (N_19043,N_18851,N_18406);
nor U19044 (N_19044,N_18606,N_18542);
nor U19045 (N_19045,N_18496,N_18803);
nand U19046 (N_19046,N_18864,N_18584);
xnor U19047 (N_19047,N_18983,N_18941);
nand U19048 (N_19048,N_18054,N_18500);
and U19049 (N_19049,N_18193,N_18627);
nor U19050 (N_19050,N_18933,N_18838);
nand U19051 (N_19051,N_18553,N_18472);
nand U19052 (N_19052,N_18143,N_18845);
or U19053 (N_19053,N_18886,N_18623);
nor U19054 (N_19054,N_18967,N_18669);
nor U19055 (N_19055,N_18044,N_18869);
and U19056 (N_19056,N_18179,N_18659);
nand U19057 (N_19057,N_18448,N_18049);
nand U19058 (N_19058,N_18714,N_18017);
nor U19059 (N_19059,N_18734,N_18648);
and U19060 (N_19060,N_18527,N_18572);
and U19061 (N_19061,N_18911,N_18778);
nor U19062 (N_19062,N_18965,N_18562);
xor U19063 (N_19063,N_18432,N_18317);
or U19064 (N_19064,N_18498,N_18964);
xor U19065 (N_19065,N_18050,N_18371);
and U19066 (N_19066,N_18910,N_18843);
or U19067 (N_19067,N_18993,N_18592);
xor U19068 (N_19068,N_18665,N_18338);
and U19069 (N_19069,N_18334,N_18060);
and U19070 (N_19070,N_18305,N_18118);
xnor U19071 (N_19071,N_18945,N_18041);
nor U19072 (N_19072,N_18512,N_18914);
nor U19073 (N_19073,N_18543,N_18263);
nor U19074 (N_19074,N_18425,N_18858);
and U19075 (N_19075,N_18635,N_18634);
and U19076 (N_19076,N_18209,N_18127);
nor U19077 (N_19077,N_18501,N_18796);
nor U19078 (N_19078,N_18369,N_18749);
xor U19079 (N_19079,N_18348,N_18538);
or U19080 (N_19080,N_18042,N_18834);
nand U19081 (N_19081,N_18676,N_18091);
xnor U19082 (N_19082,N_18654,N_18434);
and U19083 (N_19083,N_18289,N_18382);
and U19084 (N_19084,N_18293,N_18691);
or U19085 (N_19085,N_18491,N_18468);
xnor U19086 (N_19086,N_18398,N_18612);
nand U19087 (N_19087,N_18882,N_18820);
nand U19088 (N_19088,N_18765,N_18358);
or U19089 (N_19089,N_18475,N_18609);
xor U19090 (N_19090,N_18019,N_18986);
and U19091 (N_19091,N_18438,N_18856);
or U19092 (N_19092,N_18578,N_18102);
nand U19093 (N_19093,N_18645,N_18234);
and U19094 (N_19094,N_18785,N_18871);
or U19095 (N_19095,N_18247,N_18662);
and U19096 (N_19096,N_18195,N_18846);
xnor U19097 (N_19097,N_18943,N_18619);
nor U19098 (N_19098,N_18168,N_18755);
xor U19099 (N_19099,N_18847,N_18217);
and U19100 (N_19100,N_18196,N_18707);
nand U19101 (N_19101,N_18620,N_18325);
or U19102 (N_19102,N_18108,N_18640);
nand U19103 (N_19103,N_18924,N_18385);
or U19104 (N_19104,N_18359,N_18644);
and U19105 (N_19105,N_18878,N_18329);
nor U19106 (N_19106,N_18416,N_18464);
nor U19107 (N_19107,N_18715,N_18484);
nor U19108 (N_19108,N_18246,N_18804);
nor U19109 (N_19109,N_18029,N_18479);
nor U19110 (N_19110,N_18877,N_18146);
nor U19111 (N_19111,N_18138,N_18950);
nand U19112 (N_19112,N_18064,N_18974);
nand U19113 (N_19113,N_18719,N_18712);
nor U19114 (N_19114,N_18692,N_18462);
nand U19115 (N_19115,N_18387,N_18984);
and U19116 (N_19116,N_18413,N_18253);
and U19117 (N_19117,N_18567,N_18867);
nor U19118 (N_19118,N_18583,N_18025);
xor U19119 (N_19119,N_18848,N_18018);
or U19120 (N_19120,N_18313,N_18614);
and U19121 (N_19121,N_18073,N_18646);
or U19122 (N_19122,N_18150,N_18517);
nor U19123 (N_19123,N_18229,N_18232);
nand U19124 (N_19124,N_18430,N_18920);
or U19125 (N_19125,N_18568,N_18628);
and U19126 (N_19126,N_18084,N_18392);
nor U19127 (N_19127,N_18968,N_18511);
nor U19128 (N_19128,N_18693,N_18801);
nand U19129 (N_19129,N_18660,N_18880);
nor U19130 (N_19130,N_18607,N_18439);
or U19131 (N_19131,N_18935,N_18162);
nand U19132 (N_19132,N_18030,N_18779);
nor U19133 (N_19133,N_18189,N_18994);
nand U19134 (N_19134,N_18753,N_18238);
nand U19135 (N_19135,N_18395,N_18736);
xor U19136 (N_19136,N_18942,N_18431);
nor U19137 (N_19137,N_18717,N_18704);
or U19138 (N_19138,N_18565,N_18047);
or U19139 (N_19139,N_18191,N_18603);
nand U19140 (N_19140,N_18186,N_18507);
nor U19141 (N_19141,N_18113,N_18087);
xor U19142 (N_19142,N_18504,N_18696);
and U19143 (N_19143,N_18109,N_18429);
xor U19144 (N_19144,N_18744,N_18589);
nor U19145 (N_19145,N_18530,N_18107);
xnor U19146 (N_19146,N_18996,N_18723);
nand U19147 (N_19147,N_18938,N_18632);
nor U19148 (N_19148,N_18036,N_18708);
nor U19149 (N_19149,N_18452,N_18997);
or U19150 (N_19150,N_18735,N_18494);
nor U19151 (N_19151,N_18214,N_18768);
nand U19152 (N_19152,N_18061,N_18254);
nor U19153 (N_19153,N_18891,N_18503);
nor U19154 (N_19154,N_18525,N_18424);
and U19155 (N_19155,N_18016,N_18902);
and U19156 (N_19156,N_18678,N_18790);
nand U19157 (N_19157,N_18080,N_18674);
and U19158 (N_19158,N_18639,N_18916);
nor U19159 (N_19159,N_18236,N_18605);
nor U19160 (N_19160,N_18541,N_18600);
nand U19161 (N_19161,N_18142,N_18417);
and U19162 (N_19162,N_18761,N_18694);
nor U19163 (N_19163,N_18836,N_18841);
and U19164 (N_19164,N_18872,N_18969);
and U19165 (N_19165,N_18522,N_18586);
nand U19166 (N_19166,N_18937,N_18782);
nor U19167 (N_19167,N_18135,N_18633);
nor U19168 (N_19168,N_18021,N_18045);
nand U19169 (N_19169,N_18183,N_18040);
or U19170 (N_19170,N_18459,N_18825);
nand U19171 (N_19171,N_18637,N_18203);
nor U19172 (N_19172,N_18130,N_18261);
xnor U19173 (N_19173,N_18463,N_18376);
nor U19174 (N_19174,N_18184,N_18808);
nor U19175 (N_19175,N_18563,N_18251);
nor U19176 (N_19176,N_18471,N_18751);
nor U19177 (N_19177,N_18043,N_18422);
or U19178 (N_19178,N_18067,N_18420);
nand U19179 (N_19179,N_18119,N_18746);
nor U19180 (N_19180,N_18310,N_18666);
and U19181 (N_19181,N_18987,N_18766);
and U19182 (N_19182,N_18705,N_18534);
nand U19183 (N_19183,N_18668,N_18653);
xor U19184 (N_19184,N_18482,N_18690);
and U19185 (N_19185,N_18152,N_18208);
or U19186 (N_19186,N_18774,N_18290);
nor U19187 (N_19187,N_18367,N_18571);
or U19188 (N_19188,N_18124,N_18335);
and U19189 (N_19189,N_18772,N_18832);
and U19190 (N_19190,N_18613,N_18963);
or U19191 (N_19191,N_18111,N_18898);
or U19192 (N_19192,N_18881,N_18908);
and U19193 (N_19193,N_18158,N_18673);
nand U19194 (N_19194,N_18437,N_18390);
nor U19195 (N_19195,N_18591,N_18647);
nand U19196 (N_19196,N_18220,N_18893);
nand U19197 (N_19197,N_18270,N_18089);
or U19198 (N_19198,N_18741,N_18161);
or U19199 (N_19199,N_18037,N_18821);
nand U19200 (N_19200,N_18272,N_18952);
and U19201 (N_19201,N_18185,N_18651);
or U19202 (N_19202,N_18837,N_18728);
or U19203 (N_19203,N_18657,N_18393);
or U19204 (N_19204,N_18213,N_18946);
or U19205 (N_19205,N_18602,N_18245);
or U19206 (N_19206,N_18275,N_18088);
or U19207 (N_19207,N_18266,N_18314);
xnor U19208 (N_19208,N_18816,N_18068);
or U19209 (N_19209,N_18912,N_18039);
and U19210 (N_19210,N_18379,N_18394);
or U19211 (N_19211,N_18026,N_18918);
nand U19212 (N_19212,N_18810,N_18355);
or U19213 (N_19213,N_18926,N_18683);
or U19214 (N_19214,N_18331,N_18174);
and U19215 (N_19215,N_18149,N_18716);
nand U19216 (N_19216,N_18917,N_18216);
and U19217 (N_19217,N_18954,N_18115);
or U19218 (N_19218,N_18664,N_18799);
and U19219 (N_19219,N_18540,N_18888);
nor U19220 (N_19220,N_18368,N_18133);
and U19221 (N_19221,N_18281,N_18206);
nor U19222 (N_19222,N_18145,N_18642);
or U19223 (N_19223,N_18853,N_18502);
nor U19224 (N_19224,N_18787,N_18132);
or U19225 (N_19225,N_18116,N_18829);
and U19226 (N_19226,N_18703,N_18256);
or U19227 (N_19227,N_18670,N_18007);
or U19228 (N_19228,N_18802,N_18518);
and U19229 (N_19229,N_18097,N_18949);
or U19230 (N_19230,N_18066,N_18733);
or U19231 (N_19231,N_18546,N_18698);
nor U19232 (N_19232,N_18330,N_18739);
or U19233 (N_19233,N_18197,N_18156);
nand U19234 (N_19234,N_18991,N_18655);
xor U19235 (N_19235,N_18260,N_18580);
and U19236 (N_19236,N_18469,N_18128);
nor U19237 (N_19237,N_18677,N_18265);
and U19238 (N_19238,N_18302,N_18001);
or U19239 (N_19239,N_18364,N_18461);
xor U19240 (N_19240,N_18055,N_18970);
nor U19241 (N_19241,N_18188,N_18221);
and U19242 (N_19242,N_18169,N_18806);
and U19243 (N_19243,N_18874,N_18053);
or U19244 (N_19244,N_18865,N_18939);
or U19245 (N_19245,N_18885,N_18318);
nand U19246 (N_19246,N_18748,N_18493);
nor U19247 (N_19247,N_18928,N_18190);
nand U19248 (N_19248,N_18056,N_18440);
and U19249 (N_19249,N_18661,N_18913);
and U19250 (N_19250,N_18370,N_18046);
and U19251 (N_19251,N_18742,N_18791);
or U19252 (N_19252,N_18324,N_18680);
or U19253 (N_19253,N_18173,N_18667);
nor U19254 (N_19254,N_18929,N_18616);
xnor U19255 (N_19255,N_18887,N_18547);
nand U19256 (N_19256,N_18786,N_18164);
nand U19257 (N_19257,N_18312,N_18320);
nor U19258 (N_19258,N_18282,N_18552);
and U19259 (N_19259,N_18163,N_18381);
or U19260 (N_19260,N_18308,N_18485);
or U19261 (N_19261,N_18497,N_18906);
nor U19262 (N_19262,N_18224,N_18611);
or U19263 (N_19263,N_18192,N_18353);
nor U19264 (N_19264,N_18818,N_18581);
nor U19265 (N_19265,N_18028,N_18894);
nor U19266 (N_19266,N_18215,N_18982);
or U19267 (N_19267,N_18105,N_18407);
or U19268 (N_19268,N_18861,N_18112);
nor U19269 (N_19269,N_18773,N_18298);
xor U19270 (N_19270,N_18824,N_18922);
and U19271 (N_19271,N_18337,N_18889);
nand U19272 (N_19272,N_18951,N_18684);
and U19273 (N_19273,N_18962,N_18476);
nand U19274 (N_19274,N_18139,N_18085);
xnor U19275 (N_19275,N_18100,N_18656);
or U19276 (N_19276,N_18811,N_18936);
nor U19277 (N_19277,N_18307,N_18481);
or U19278 (N_19278,N_18792,N_18784);
and U19279 (N_19279,N_18137,N_18815);
nor U19280 (N_19280,N_18483,N_18579);
nor U19281 (N_19281,N_18957,N_18271);
nand U19282 (N_19282,N_18608,N_18134);
nand U19283 (N_19283,N_18200,N_18288);
or U19284 (N_19284,N_18593,N_18658);
and U19285 (N_19285,N_18795,N_18240);
or U19286 (N_19286,N_18235,N_18890);
and U19287 (N_19287,N_18278,N_18365);
nor U19288 (N_19288,N_18564,N_18629);
xnor U19289 (N_19289,N_18830,N_18243);
or U19290 (N_19290,N_18737,N_18255);
or U19291 (N_19291,N_18233,N_18062);
nand U19292 (N_19292,N_18789,N_18450);
or U19293 (N_19293,N_18351,N_18297);
nand U19294 (N_19294,N_18095,N_18349);
nand U19295 (N_19295,N_18435,N_18160);
or U19296 (N_19296,N_18386,N_18433);
and U19297 (N_19297,N_18120,N_18219);
nor U19298 (N_19298,N_18362,N_18363);
nor U19299 (N_19299,N_18762,N_18875);
nor U19300 (N_19300,N_18269,N_18083);
nand U19301 (N_19301,N_18129,N_18495);
or U19302 (N_19302,N_18539,N_18126);
nor U19303 (N_19303,N_18944,N_18577);
nand U19304 (N_19304,N_18321,N_18977);
or U19305 (N_19305,N_18177,N_18180);
nand U19306 (N_19306,N_18397,N_18159);
xnor U19307 (N_19307,N_18131,N_18490);
xnor U19308 (N_19308,N_18277,N_18514);
nor U19309 (N_19309,N_18923,N_18587);
or U19310 (N_19310,N_18280,N_18304);
nor U19311 (N_19311,N_18998,N_18681);
nor U19312 (N_19312,N_18166,N_18566);
and U19313 (N_19313,N_18383,N_18899);
and U19314 (N_19314,N_18403,N_18250);
nor U19315 (N_19315,N_18332,N_18421);
nand U19316 (N_19316,N_18022,N_18823);
nor U19317 (N_19317,N_18315,N_18573);
nand U19318 (N_19318,N_18038,N_18560);
nor U19319 (N_19319,N_18812,N_18915);
xnor U19320 (N_19320,N_18339,N_18415);
nand U19321 (N_19321,N_18826,N_18720);
or U19322 (N_19322,N_18024,N_18155);
or U19323 (N_19323,N_18961,N_18117);
nor U19324 (N_19324,N_18862,N_18372);
nand U19325 (N_19325,N_18199,N_18817);
nor U19326 (N_19326,N_18299,N_18958);
and U19327 (N_19327,N_18601,N_18679);
nor U19328 (N_19328,N_18740,N_18506);
or U19329 (N_19329,N_18374,N_18771);
or U19330 (N_19330,N_18165,N_18389);
or U19331 (N_19331,N_18098,N_18897);
or U19332 (N_19332,N_18989,N_18081);
xnor U19333 (N_19333,N_18978,N_18559);
nor U19334 (N_19334,N_18524,N_18863);
and U19335 (N_19335,N_18366,N_18455);
nor U19336 (N_19336,N_18446,N_18451);
nand U19337 (N_19337,N_18813,N_18356);
or U19338 (N_19338,N_18797,N_18903);
nor U19339 (N_19339,N_18621,N_18594);
nand U19340 (N_19340,N_18172,N_18695);
xnor U19341 (N_19341,N_18034,N_18550);
and U19342 (N_19342,N_18093,N_18548);
xor U19343 (N_19343,N_18096,N_18859);
or U19344 (N_19344,N_18070,N_18059);
or U19345 (N_19345,N_18099,N_18776);
and U19346 (N_19346,N_18883,N_18336);
and U19347 (N_19347,N_18857,N_18625);
or U19348 (N_19348,N_18852,N_18842);
nor U19349 (N_19349,N_18063,N_18285);
nand U19350 (N_19350,N_18354,N_18373);
nor U19351 (N_19351,N_18110,N_18474);
nor U19352 (N_19352,N_18342,N_18763);
nor U19353 (N_19353,N_18035,N_18671);
or U19354 (N_19354,N_18685,N_18819);
nor U19355 (N_19355,N_18757,N_18925);
nor U19356 (N_19356,N_18000,N_18569);
and U19357 (N_19357,N_18210,N_18082);
or U19358 (N_19358,N_18752,N_18649);
nand U19359 (N_19359,N_18532,N_18274);
and U19360 (N_19360,N_18948,N_18876);
and U19361 (N_19361,N_18140,N_18556);
nand U19362 (N_19362,N_18839,N_18011);
xnor U19363 (N_19363,N_18006,N_18956);
or U19364 (N_19364,N_18284,N_18777);
and U19365 (N_19365,N_18136,N_18775);
and U19366 (N_19366,N_18545,N_18870);
nand U19367 (N_19367,N_18973,N_18268);
nor U19368 (N_19368,N_18622,N_18724);
nand U19369 (N_19369,N_18521,N_18999);
xnor U19370 (N_19370,N_18079,N_18835);
nor U19371 (N_19371,N_18178,N_18709);
and U19372 (N_19372,N_18104,N_18953);
or U19373 (N_19373,N_18230,N_18441);
nor U19374 (N_19374,N_18896,N_18610);
xnor U19375 (N_19375,N_18194,N_18489);
nand U19376 (N_19376,N_18057,N_18300);
or U19377 (N_19377,N_18805,N_18443);
nor U19378 (N_19378,N_18058,N_18346);
nand U19379 (N_19379,N_18380,N_18972);
and U19380 (N_19380,N_18157,N_18689);
nor U19381 (N_19381,N_18478,N_18981);
nand U19382 (N_19382,N_18377,N_18588);
or U19383 (N_19383,N_18125,N_18682);
nand U19384 (N_19384,N_18357,N_18202);
nand U19385 (N_19385,N_18151,N_18767);
nor U19386 (N_19386,N_18731,N_18012);
and U19387 (N_19387,N_18617,N_18453);
and U19388 (N_19388,N_18615,N_18900);
or U19389 (N_19389,N_18960,N_18992);
or U19390 (N_19390,N_18860,N_18531);
nand U19391 (N_19391,N_18286,N_18574);
and U19392 (N_19392,N_18004,N_18905);
nand U19393 (N_19393,N_18114,N_18959);
and U19394 (N_19394,N_18537,N_18457);
nand U19395 (N_19395,N_18449,N_18316);
nor U19396 (N_19396,N_18181,N_18241);
nand U19397 (N_19397,N_18895,N_18076);
nor U19398 (N_19398,N_18599,N_18408);
nor U19399 (N_19399,N_18650,N_18175);
or U19400 (N_19400,N_18322,N_18436);
nand U19401 (N_19401,N_18401,N_18249);
nand U19402 (N_19402,N_18971,N_18781);
xnor U19403 (N_19403,N_18283,N_18686);
nand U19404 (N_19404,N_18227,N_18345);
xor U19405 (N_19405,N_18743,N_18287);
nand U19406 (N_19406,N_18010,N_18447);
nor U19407 (N_19407,N_18576,N_18934);
or U19408 (N_19408,N_18979,N_18636);
nand U19409 (N_19409,N_18509,N_18003);
and U19410 (N_19410,N_18410,N_18176);
or U19411 (N_19411,N_18561,N_18207);
or U19412 (N_19412,N_18201,N_18725);
or U19413 (N_19413,N_18788,N_18170);
xor U19414 (N_19414,N_18244,N_18713);
and U19415 (N_19415,N_18412,N_18074);
nand U19416 (N_19416,N_18405,N_18419);
nor U19417 (N_19417,N_18077,N_18427);
and U19418 (N_19418,N_18396,N_18975);
and U19419 (N_19419,N_18182,N_18409);
nor U19420 (N_19420,N_18326,N_18466);
or U19421 (N_19421,N_18328,N_18738);
and U19422 (N_19422,N_18276,N_18226);
or U19423 (N_19423,N_18121,N_18809);
nor U19424 (N_19424,N_18460,N_18258);
or U19425 (N_19425,N_18759,N_18536);
or U19426 (N_19426,N_18702,N_18205);
nor U19427 (N_19427,N_18187,N_18465);
or U19428 (N_19428,N_18499,N_18154);
nand U19429 (N_19429,N_18123,N_18919);
or U19430 (N_19430,N_18932,N_18631);
or U19431 (N_19431,N_18849,N_18153);
or U19432 (N_19432,N_18688,N_18595);
xor U19433 (N_19433,N_18344,N_18212);
xor U19434 (N_19434,N_18259,N_18955);
or U19435 (N_19435,N_18023,N_18549);
nor U19436 (N_19436,N_18515,N_18005);
or U19437 (N_19437,N_18701,N_18697);
or U19438 (N_19438,N_18319,N_18624);
or U19439 (N_19439,N_18384,N_18807);
nor U19440 (N_19440,N_18590,N_18598);
xor U19441 (N_19441,N_18103,N_18756);
and U19442 (N_19442,N_18930,N_18855);
nand U19443 (N_19443,N_18078,N_18840);
xnor U19444 (N_19444,N_18947,N_18343);
and U19445 (N_19445,N_18711,N_18988);
and U19446 (N_19446,N_18218,N_18513);
or U19447 (N_19447,N_18726,N_18361);
and U19448 (N_19448,N_18575,N_18822);
nor U19449 (N_19449,N_18800,N_18301);
nand U19450 (N_19450,N_18273,N_18292);
and U19451 (N_19451,N_18122,N_18597);
nor U19452 (N_19452,N_18071,N_18570);
nand U19453 (N_19453,N_18663,N_18844);
nor U19454 (N_19454,N_18428,N_18764);
nand U19455 (N_19455,N_18699,N_18106);
nor U19456 (N_19456,N_18228,N_18486);
nor U19457 (N_19457,N_18052,N_18854);
xor U19458 (N_19458,N_18231,N_18492);
nand U19459 (N_19459,N_18884,N_18904);
or U19460 (N_19460,N_18675,N_18327);
or U19461 (N_19461,N_18020,N_18706);
or U19462 (N_19462,N_18323,N_18828);
nand U19463 (N_19463,N_18827,N_18582);
xor U19464 (N_19464,N_18907,N_18528);
and U19465 (N_19465,N_18222,N_18794);
and U19466 (N_19466,N_18526,N_18008);
nor U19467 (N_19467,N_18833,N_18094);
xor U19468 (N_19468,N_18931,N_18710);
or U19469 (N_19469,N_18558,N_18480);
xnor U19470 (N_19470,N_18090,N_18976);
and U19471 (N_19471,N_18520,N_18454);
nand U19472 (N_19472,N_18198,N_18783);
nand U19473 (N_19473,N_18966,N_18141);
and U19474 (N_19474,N_18015,N_18554);
or U19475 (N_19475,N_18239,N_18048);
or U19476 (N_19476,N_18211,N_18487);
and U19477 (N_19477,N_18652,N_18780);
and U19478 (N_19478,N_18388,N_18237);
and U19479 (N_19479,N_18641,N_18262);
nor U19480 (N_19480,N_18360,N_18445);
nor U19481 (N_19481,N_18585,N_18014);
and U19482 (N_19482,N_18596,N_18510);
xnor U19483 (N_19483,N_18444,N_18171);
nor U19484 (N_19484,N_18519,N_18295);
xor U19485 (N_19485,N_18291,N_18793);
nand U19486 (N_19486,N_18009,N_18267);
or U19487 (N_19487,N_18065,N_18306);
nand U19488 (N_19488,N_18311,N_18347);
or U19489 (N_19489,N_18535,N_18995);
xor U19490 (N_19490,N_18423,N_18378);
nor U19491 (N_19491,N_18892,N_18086);
nor U19492 (N_19492,N_18985,N_18721);
or U19493 (N_19493,N_18814,N_18296);
and U19494 (N_19494,N_18391,N_18488);
nand U19495 (N_19495,N_18167,N_18831);
nand U19496 (N_19496,N_18643,N_18031);
nand U19497 (N_19497,N_18626,N_18051);
or U19498 (N_19498,N_18529,N_18533);
and U19499 (N_19499,N_18604,N_18352);
or U19500 (N_19500,N_18227,N_18058);
nor U19501 (N_19501,N_18597,N_18945);
and U19502 (N_19502,N_18413,N_18857);
or U19503 (N_19503,N_18497,N_18592);
nand U19504 (N_19504,N_18568,N_18651);
xor U19505 (N_19505,N_18659,N_18752);
or U19506 (N_19506,N_18664,N_18652);
and U19507 (N_19507,N_18997,N_18999);
nor U19508 (N_19508,N_18983,N_18421);
and U19509 (N_19509,N_18238,N_18532);
xor U19510 (N_19510,N_18142,N_18759);
and U19511 (N_19511,N_18205,N_18851);
nand U19512 (N_19512,N_18468,N_18372);
or U19513 (N_19513,N_18901,N_18904);
nor U19514 (N_19514,N_18477,N_18613);
xnor U19515 (N_19515,N_18826,N_18916);
nor U19516 (N_19516,N_18911,N_18627);
and U19517 (N_19517,N_18620,N_18305);
or U19518 (N_19518,N_18377,N_18442);
nand U19519 (N_19519,N_18898,N_18385);
xnor U19520 (N_19520,N_18065,N_18452);
and U19521 (N_19521,N_18575,N_18303);
nor U19522 (N_19522,N_18893,N_18969);
nand U19523 (N_19523,N_18875,N_18081);
nor U19524 (N_19524,N_18911,N_18380);
nand U19525 (N_19525,N_18442,N_18495);
nor U19526 (N_19526,N_18994,N_18581);
or U19527 (N_19527,N_18621,N_18179);
or U19528 (N_19528,N_18501,N_18460);
or U19529 (N_19529,N_18929,N_18973);
nand U19530 (N_19530,N_18403,N_18950);
xnor U19531 (N_19531,N_18838,N_18667);
nand U19532 (N_19532,N_18381,N_18970);
or U19533 (N_19533,N_18434,N_18323);
or U19534 (N_19534,N_18044,N_18005);
nor U19535 (N_19535,N_18951,N_18284);
and U19536 (N_19536,N_18893,N_18034);
or U19537 (N_19537,N_18003,N_18005);
xor U19538 (N_19538,N_18051,N_18383);
and U19539 (N_19539,N_18310,N_18179);
and U19540 (N_19540,N_18907,N_18997);
nor U19541 (N_19541,N_18510,N_18313);
nand U19542 (N_19542,N_18545,N_18812);
xor U19543 (N_19543,N_18111,N_18175);
or U19544 (N_19544,N_18112,N_18692);
nor U19545 (N_19545,N_18175,N_18436);
nor U19546 (N_19546,N_18505,N_18166);
nand U19547 (N_19547,N_18919,N_18726);
and U19548 (N_19548,N_18518,N_18730);
or U19549 (N_19549,N_18209,N_18919);
nand U19550 (N_19550,N_18924,N_18086);
and U19551 (N_19551,N_18505,N_18775);
or U19552 (N_19552,N_18978,N_18584);
nand U19553 (N_19553,N_18697,N_18939);
nand U19554 (N_19554,N_18567,N_18093);
xor U19555 (N_19555,N_18091,N_18126);
nand U19556 (N_19556,N_18090,N_18637);
xnor U19557 (N_19557,N_18824,N_18059);
or U19558 (N_19558,N_18502,N_18205);
nor U19559 (N_19559,N_18185,N_18514);
or U19560 (N_19560,N_18500,N_18073);
nand U19561 (N_19561,N_18650,N_18624);
nand U19562 (N_19562,N_18797,N_18866);
and U19563 (N_19563,N_18087,N_18852);
or U19564 (N_19564,N_18339,N_18439);
nand U19565 (N_19565,N_18046,N_18787);
and U19566 (N_19566,N_18573,N_18072);
or U19567 (N_19567,N_18992,N_18354);
nor U19568 (N_19568,N_18684,N_18234);
nand U19569 (N_19569,N_18727,N_18211);
nor U19570 (N_19570,N_18513,N_18216);
or U19571 (N_19571,N_18259,N_18711);
and U19572 (N_19572,N_18729,N_18188);
and U19573 (N_19573,N_18583,N_18246);
xnor U19574 (N_19574,N_18116,N_18915);
or U19575 (N_19575,N_18587,N_18961);
nor U19576 (N_19576,N_18761,N_18513);
or U19577 (N_19577,N_18929,N_18808);
nand U19578 (N_19578,N_18405,N_18913);
nand U19579 (N_19579,N_18295,N_18079);
xnor U19580 (N_19580,N_18182,N_18261);
and U19581 (N_19581,N_18394,N_18263);
nor U19582 (N_19582,N_18205,N_18050);
nand U19583 (N_19583,N_18923,N_18897);
and U19584 (N_19584,N_18146,N_18354);
nor U19585 (N_19585,N_18792,N_18398);
nor U19586 (N_19586,N_18196,N_18279);
nand U19587 (N_19587,N_18280,N_18765);
nand U19588 (N_19588,N_18910,N_18326);
xnor U19589 (N_19589,N_18310,N_18732);
or U19590 (N_19590,N_18237,N_18169);
and U19591 (N_19591,N_18056,N_18219);
or U19592 (N_19592,N_18807,N_18698);
nor U19593 (N_19593,N_18799,N_18122);
nor U19594 (N_19594,N_18828,N_18893);
and U19595 (N_19595,N_18909,N_18629);
and U19596 (N_19596,N_18112,N_18049);
or U19597 (N_19597,N_18715,N_18356);
xor U19598 (N_19598,N_18321,N_18801);
and U19599 (N_19599,N_18496,N_18285);
or U19600 (N_19600,N_18514,N_18508);
nor U19601 (N_19601,N_18820,N_18085);
nand U19602 (N_19602,N_18555,N_18398);
xor U19603 (N_19603,N_18467,N_18813);
nor U19604 (N_19604,N_18945,N_18755);
and U19605 (N_19605,N_18495,N_18248);
or U19606 (N_19606,N_18042,N_18714);
and U19607 (N_19607,N_18070,N_18135);
nor U19608 (N_19608,N_18302,N_18445);
nand U19609 (N_19609,N_18634,N_18903);
or U19610 (N_19610,N_18777,N_18346);
xor U19611 (N_19611,N_18423,N_18029);
nand U19612 (N_19612,N_18291,N_18454);
or U19613 (N_19613,N_18095,N_18760);
or U19614 (N_19614,N_18865,N_18242);
or U19615 (N_19615,N_18069,N_18842);
and U19616 (N_19616,N_18030,N_18630);
nand U19617 (N_19617,N_18604,N_18984);
and U19618 (N_19618,N_18795,N_18143);
nor U19619 (N_19619,N_18159,N_18309);
nor U19620 (N_19620,N_18537,N_18376);
and U19621 (N_19621,N_18973,N_18832);
nor U19622 (N_19622,N_18274,N_18903);
xor U19623 (N_19623,N_18399,N_18032);
xor U19624 (N_19624,N_18021,N_18652);
xnor U19625 (N_19625,N_18626,N_18653);
or U19626 (N_19626,N_18285,N_18098);
nand U19627 (N_19627,N_18165,N_18551);
nor U19628 (N_19628,N_18383,N_18178);
and U19629 (N_19629,N_18269,N_18716);
or U19630 (N_19630,N_18329,N_18089);
nand U19631 (N_19631,N_18215,N_18114);
nand U19632 (N_19632,N_18424,N_18169);
xnor U19633 (N_19633,N_18693,N_18360);
nor U19634 (N_19634,N_18033,N_18775);
nor U19635 (N_19635,N_18264,N_18505);
nand U19636 (N_19636,N_18238,N_18730);
nand U19637 (N_19637,N_18210,N_18031);
and U19638 (N_19638,N_18672,N_18114);
nand U19639 (N_19639,N_18278,N_18656);
or U19640 (N_19640,N_18813,N_18593);
nand U19641 (N_19641,N_18909,N_18645);
or U19642 (N_19642,N_18830,N_18373);
nor U19643 (N_19643,N_18124,N_18016);
xor U19644 (N_19644,N_18234,N_18330);
xor U19645 (N_19645,N_18372,N_18981);
nand U19646 (N_19646,N_18362,N_18250);
nor U19647 (N_19647,N_18728,N_18680);
xnor U19648 (N_19648,N_18524,N_18311);
or U19649 (N_19649,N_18586,N_18001);
and U19650 (N_19650,N_18789,N_18237);
nand U19651 (N_19651,N_18310,N_18889);
nand U19652 (N_19652,N_18033,N_18971);
nand U19653 (N_19653,N_18189,N_18411);
nand U19654 (N_19654,N_18279,N_18387);
and U19655 (N_19655,N_18513,N_18634);
nand U19656 (N_19656,N_18582,N_18279);
nor U19657 (N_19657,N_18120,N_18027);
or U19658 (N_19658,N_18701,N_18295);
and U19659 (N_19659,N_18987,N_18223);
nor U19660 (N_19660,N_18716,N_18482);
and U19661 (N_19661,N_18318,N_18690);
nand U19662 (N_19662,N_18239,N_18433);
nand U19663 (N_19663,N_18922,N_18840);
and U19664 (N_19664,N_18857,N_18108);
or U19665 (N_19665,N_18452,N_18049);
and U19666 (N_19666,N_18681,N_18010);
or U19667 (N_19667,N_18197,N_18256);
and U19668 (N_19668,N_18894,N_18395);
or U19669 (N_19669,N_18155,N_18203);
nand U19670 (N_19670,N_18495,N_18855);
and U19671 (N_19671,N_18776,N_18020);
and U19672 (N_19672,N_18732,N_18736);
nor U19673 (N_19673,N_18781,N_18254);
or U19674 (N_19674,N_18333,N_18322);
nor U19675 (N_19675,N_18994,N_18841);
nor U19676 (N_19676,N_18520,N_18055);
or U19677 (N_19677,N_18322,N_18352);
nor U19678 (N_19678,N_18653,N_18177);
nor U19679 (N_19679,N_18684,N_18562);
and U19680 (N_19680,N_18371,N_18567);
and U19681 (N_19681,N_18813,N_18758);
xor U19682 (N_19682,N_18463,N_18337);
xor U19683 (N_19683,N_18548,N_18657);
nor U19684 (N_19684,N_18105,N_18901);
and U19685 (N_19685,N_18224,N_18729);
and U19686 (N_19686,N_18334,N_18776);
or U19687 (N_19687,N_18834,N_18754);
and U19688 (N_19688,N_18220,N_18306);
nor U19689 (N_19689,N_18644,N_18225);
and U19690 (N_19690,N_18495,N_18804);
or U19691 (N_19691,N_18437,N_18528);
nand U19692 (N_19692,N_18715,N_18160);
or U19693 (N_19693,N_18798,N_18308);
nand U19694 (N_19694,N_18603,N_18814);
nand U19695 (N_19695,N_18530,N_18263);
and U19696 (N_19696,N_18949,N_18140);
nor U19697 (N_19697,N_18699,N_18016);
and U19698 (N_19698,N_18206,N_18612);
and U19699 (N_19699,N_18708,N_18975);
nor U19700 (N_19700,N_18069,N_18714);
and U19701 (N_19701,N_18899,N_18390);
nor U19702 (N_19702,N_18136,N_18836);
nand U19703 (N_19703,N_18789,N_18340);
and U19704 (N_19704,N_18814,N_18881);
nand U19705 (N_19705,N_18858,N_18107);
or U19706 (N_19706,N_18431,N_18463);
and U19707 (N_19707,N_18717,N_18686);
nand U19708 (N_19708,N_18158,N_18619);
or U19709 (N_19709,N_18234,N_18242);
or U19710 (N_19710,N_18305,N_18161);
or U19711 (N_19711,N_18981,N_18744);
nor U19712 (N_19712,N_18482,N_18823);
and U19713 (N_19713,N_18271,N_18088);
nor U19714 (N_19714,N_18792,N_18820);
and U19715 (N_19715,N_18148,N_18637);
or U19716 (N_19716,N_18454,N_18218);
and U19717 (N_19717,N_18916,N_18499);
nand U19718 (N_19718,N_18806,N_18170);
nor U19719 (N_19719,N_18949,N_18159);
and U19720 (N_19720,N_18479,N_18363);
or U19721 (N_19721,N_18239,N_18337);
and U19722 (N_19722,N_18860,N_18116);
or U19723 (N_19723,N_18131,N_18740);
and U19724 (N_19724,N_18994,N_18350);
nor U19725 (N_19725,N_18958,N_18020);
nor U19726 (N_19726,N_18466,N_18969);
nor U19727 (N_19727,N_18392,N_18746);
nand U19728 (N_19728,N_18336,N_18309);
and U19729 (N_19729,N_18059,N_18653);
or U19730 (N_19730,N_18626,N_18851);
xnor U19731 (N_19731,N_18295,N_18052);
nand U19732 (N_19732,N_18805,N_18880);
nor U19733 (N_19733,N_18282,N_18831);
nor U19734 (N_19734,N_18375,N_18928);
or U19735 (N_19735,N_18026,N_18398);
nand U19736 (N_19736,N_18935,N_18647);
nand U19737 (N_19737,N_18489,N_18880);
or U19738 (N_19738,N_18831,N_18057);
and U19739 (N_19739,N_18623,N_18740);
and U19740 (N_19740,N_18372,N_18156);
nor U19741 (N_19741,N_18436,N_18303);
nand U19742 (N_19742,N_18624,N_18388);
and U19743 (N_19743,N_18413,N_18462);
or U19744 (N_19744,N_18988,N_18250);
or U19745 (N_19745,N_18171,N_18388);
xor U19746 (N_19746,N_18703,N_18696);
xnor U19747 (N_19747,N_18036,N_18395);
and U19748 (N_19748,N_18611,N_18594);
or U19749 (N_19749,N_18181,N_18331);
and U19750 (N_19750,N_18896,N_18366);
or U19751 (N_19751,N_18895,N_18074);
xnor U19752 (N_19752,N_18557,N_18674);
or U19753 (N_19753,N_18019,N_18752);
or U19754 (N_19754,N_18603,N_18806);
nor U19755 (N_19755,N_18564,N_18090);
nand U19756 (N_19756,N_18998,N_18296);
nor U19757 (N_19757,N_18499,N_18862);
nand U19758 (N_19758,N_18260,N_18296);
nor U19759 (N_19759,N_18238,N_18137);
nand U19760 (N_19760,N_18472,N_18807);
or U19761 (N_19761,N_18720,N_18621);
nor U19762 (N_19762,N_18009,N_18703);
and U19763 (N_19763,N_18808,N_18161);
xnor U19764 (N_19764,N_18555,N_18154);
or U19765 (N_19765,N_18247,N_18197);
nor U19766 (N_19766,N_18421,N_18904);
nor U19767 (N_19767,N_18745,N_18050);
or U19768 (N_19768,N_18254,N_18514);
and U19769 (N_19769,N_18344,N_18252);
nand U19770 (N_19770,N_18913,N_18430);
or U19771 (N_19771,N_18627,N_18328);
nand U19772 (N_19772,N_18889,N_18163);
xor U19773 (N_19773,N_18846,N_18428);
or U19774 (N_19774,N_18250,N_18377);
xor U19775 (N_19775,N_18468,N_18676);
or U19776 (N_19776,N_18714,N_18111);
nor U19777 (N_19777,N_18795,N_18956);
nand U19778 (N_19778,N_18700,N_18981);
and U19779 (N_19779,N_18725,N_18697);
and U19780 (N_19780,N_18116,N_18335);
nor U19781 (N_19781,N_18759,N_18458);
and U19782 (N_19782,N_18672,N_18906);
nand U19783 (N_19783,N_18959,N_18656);
nand U19784 (N_19784,N_18712,N_18727);
xor U19785 (N_19785,N_18965,N_18597);
or U19786 (N_19786,N_18352,N_18184);
and U19787 (N_19787,N_18717,N_18369);
and U19788 (N_19788,N_18501,N_18120);
and U19789 (N_19789,N_18291,N_18387);
or U19790 (N_19790,N_18625,N_18378);
nand U19791 (N_19791,N_18172,N_18455);
and U19792 (N_19792,N_18604,N_18709);
and U19793 (N_19793,N_18745,N_18537);
nor U19794 (N_19794,N_18939,N_18037);
nand U19795 (N_19795,N_18952,N_18569);
or U19796 (N_19796,N_18949,N_18586);
and U19797 (N_19797,N_18728,N_18627);
nor U19798 (N_19798,N_18802,N_18928);
or U19799 (N_19799,N_18372,N_18902);
xnor U19800 (N_19800,N_18720,N_18097);
and U19801 (N_19801,N_18429,N_18785);
and U19802 (N_19802,N_18453,N_18417);
nor U19803 (N_19803,N_18510,N_18522);
nand U19804 (N_19804,N_18117,N_18254);
and U19805 (N_19805,N_18551,N_18780);
or U19806 (N_19806,N_18317,N_18696);
or U19807 (N_19807,N_18962,N_18217);
nand U19808 (N_19808,N_18197,N_18614);
nand U19809 (N_19809,N_18898,N_18231);
xor U19810 (N_19810,N_18965,N_18804);
nand U19811 (N_19811,N_18666,N_18869);
nor U19812 (N_19812,N_18643,N_18516);
nor U19813 (N_19813,N_18106,N_18254);
nand U19814 (N_19814,N_18880,N_18225);
and U19815 (N_19815,N_18267,N_18418);
nand U19816 (N_19816,N_18467,N_18610);
and U19817 (N_19817,N_18074,N_18826);
nor U19818 (N_19818,N_18649,N_18403);
nor U19819 (N_19819,N_18054,N_18408);
or U19820 (N_19820,N_18776,N_18520);
nor U19821 (N_19821,N_18704,N_18252);
nand U19822 (N_19822,N_18510,N_18602);
nor U19823 (N_19823,N_18094,N_18421);
and U19824 (N_19824,N_18596,N_18501);
nor U19825 (N_19825,N_18091,N_18536);
or U19826 (N_19826,N_18921,N_18268);
xor U19827 (N_19827,N_18758,N_18534);
and U19828 (N_19828,N_18903,N_18265);
nand U19829 (N_19829,N_18335,N_18529);
or U19830 (N_19830,N_18251,N_18826);
and U19831 (N_19831,N_18033,N_18162);
nand U19832 (N_19832,N_18154,N_18105);
nand U19833 (N_19833,N_18569,N_18736);
and U19834 (N_19834,N_18732,N_18119);
nor U19835 (N_19835,N_18487,N_18277);
xor U19836 (N_19836,N_18688,N_18628);
and U19837 (N_19837,N_18645,N_18611);
nor U19838 (N_19838,N_18645,N_18163);
nor U19839 (N_19839,N_18355,N_18789);
xnor U19840 (N_19840,N_18857,N_18704);
nand U19841 (N_19841,N_18480,N_18037);
nor U19842 (N_19842,N_18660,N_18062);
and U19843 (N_19843,N_18577,N_18667);
and U19844 (N_19844,N_18573,N_18513);
and U19845 (N_19845,N_18354,N_18785);
xor U19846 (N_19846,N_18742,N_18220);
or U19847 (N_19847,N_18447,N_18164);
nor U19848 (N_19848,N_18797,N_18543);
nor U19849 (N_19849,N_18166,N_18115);
nor U19850 (N_19850,N_18505,N_18859);
nor U19851 (N_19851,N_18363,N_18972);
or U19852 (N_19852,N_18305,N_18419);
nand U19853 (N_19853,N_18790,N_18541);
or U19854 (N_19854,N_18291,N_18495);
nor U19855 (N_19855,N_18918,N_18983);
nor U19856 (N_19856,N_18525,N_18830);
and U19857 (N_19857,N_18295,N_18310);
and U19858 (N_19858,N_18614,N_18747);
nand U19859 (N_19859,N_18961,N_18454);
or U19860 (N_19860,N_18462,N_18215);
nor U19861 (N_19861,N_18228,N_18411);
nand U19862 (N_19862,N_18822,N_18215);
xor U19863 (N_19863,N_18848,N_18815);
or U19864 (N_19864,N_18811,N_18462);
or U19865 (N_19865,N_18955,N_18320);
or U19866 (N_19866,N_18898,N_18507);
nor U19867 (N_19867,N_18144,N_18373);
nand U19868 (N_19868,N_18089,N_18421);
nor U19869 (N_19869,N_18637,N_18963);
nand U19870 (N_19870,N_18661,N_18398);
xnor U19871 (N_19871,N_18591,N_18055);
nand U19872 (N_19872,N_18131,N_18012);
nor U19873 (N_19873,N_18235,N_18440);
and U19874 (N_19874,N_18287,N_18346);
nor U19875 (N_19875,N_18723,N_18069);
nand U19876 (N_19876,N_18989,N_18342);
nand U19877 (N_19877,N_18917,N_18069);
nand U19878 (N_19878,N_18850,N_18138);
and U19879 (N_19879,N_18900,N_18167);
xor U19880 (N_19880,N_18947,N_18235);
xor U19881 (N_19881,N_18391,N_18836);
nor U19882 (N_19882,N_18223,N_18996);
nand U19883 (N_19883,N_18106,N_18535);
or U19884 (N_19884,N_18921,N_18494);
and U19885 (N_19885,N_18027,N_18720);
nand U19886 (N_19886,N_18857,N_18139);
nor U19887 (N_19887,N_18667,N_18829);
and U19888 (N_19888,N_18878,N_18776);
nor U19889 (N_19889,N_18547,N_18878);
and U19890 (N_19890,N_18074,N_18234);
nor U19891 (N_19891,N_18512,N_18167);
nand U19892 (N_19892,N_18410,N_18381);
nand U19893 (N_19893,N_18375,N_18113);
and U19894 (N_19894,N_18142,N_18839);
nand U19895 (N_19895,N_18278,N_18808);
or U19896 (N_19896,N_18051,N_18816);
nand U19897 (N_19897,N_18612,N_18622);
and U19898 (N_19898,N_18125,N_18022);
or U19899 (N_19899,N_18476,N_18560);
nor U19900 (N_19900,N_18772,N_18704);
and U19901 (N_19901,N_18227,N_18480);
nor U19902 (N_19902,N_18044,N_18887);
and U19903 (N_19903,N_18991,N_18458);
and U19904 (N_19904,N_18484,N_18797);
or U19905 (N_19905,N_18633,N_18618);
or U19906 (N_19906,N_18979,N_18414);
nand U19907 (N_19907,N_18845,N_18725);
or U19908 (N_19908,N_18324,N_18107);
and U19909 (N_19909,N_18740,N_18690);
and U19910 (N_19910,N_18584,N_18963);
and U19911 (N_19911,N_18346,N_18444);
nor U19912 (N_19912,N_18283,N_18438);
nor U19913 (N_19913,N_18032,N_18352);
nand U19914 (N_19914,N_18146,N_18922);
nand U19915 (N_19915,N_18044,N_18466);
nor U19916 (N_19916,N_18286,N_18313);
nor U19917 (N_19917,N_18110,N_18497);
nor U19918 (N_19918,N_18738,N_18728);
or U19919 (N_19919,N_18548,N_18520);
and U19920 (N_19920,N_18616,N_18211);
or U19921 (N_19921,N_18086,N_18449);
nand U19922 (N_19922,N_18803,N_18106);
and U19923 (N_19923,N_18309,N_18243);
and U19924 (N_19924,N_18316,N_18642);
and U19925 (N_19925,N_18742,N_18376);
and U19926 (N_19926,N_18795,N_18851);
and U19927 (N_19927,N_18473,N_18171);
nor U19928 (N_19928,N_18766,N_18145);
xnor U19929 (N_19929,N_18270,N_18338);
and U19930 (N_19930,N_18787,N_18560);
nor U19931 (N_19931,N_18321,N_18778);
and U19932 (N_19932,N_18231,N_18028);
or U19933 (N_19933,N_18491,N_18473);
or U19934 (N_19934,N_18864,N_18006);
and U19935 (N_19935,N_18650,N_18326);
nor U19936 (N_19936,N_18670,N_18562);
nand U19937 (N_19937,N_18531,N_18468);
nand U19938 (N_19938,N_18877,N_18137);
nand U19939 (N_19939,N_18918,N_18539);
xnor U19940 (N_19940,N_18685,N_18436);
nor U19941 (N_19941,N_18619,N_18937);
nand U19942 (N_19942,N_18512,N_18840);
nor U19943 (N_19943,N_18476,N_18024);
nand U19944 (N_19944,N_18620,N_18380);
nand U19945 (N_19945,N_18785,N_18860);
and U19946 (N_19946,N_18622,N_18333);
nor U19947 (N_19947,N_18719,N_18877);
or U19948 (N_19948,N_18162,N_18222);
xor U19949 (N_19949,N_18096,N_18850);
nand U19950 (N_19950,N_18966,N_18158);
nor U19951 (N_19951,N_18898,N_18444);
nor U19952 (N_19952,N_18775,N_18923);
or U19953 (N_19953,N_18145,N_18071);
xor U19954 (N_19954,N_18511,N_18393);
or U19955 (N_19955,N_18595,N_18883);
nand U19956 (N_19956,N_18336,N_18337);
or U19957 (N_19957,N_18491,N_18395);
and U19958 (N_19958,N_18301,N_18976);
nand U19959 (N_19959,N_18613,N_18686);
nor U19960 (N_19960,N_18466,N_18421);
or U19961 (N_19961,N_18223,N_18702);
or U19962 (N_19962,N_18956,N_18774);
nand U19963 (N_19963,N_18121,N_18269);
and U19964 (N_19964,N_18756,N_18842);
xor U19965 (N_19965,N_18566,N_18278);
and U19966 (N_19966,N_18745,N_18253);
and U19967 (N_19967,N_18319,N_18487);
nand U19968 (N_19968,N_18558,N_18200);
nand U19969 (N_19969,N_18997,N_18475);
nor U19970 (N_19970,N_18776,N_18359);
nor U19971 (N_19971,N_18055,N_18330);
nand U19972 (N_19972,N_18179,N_18772);
xnor U19973 (N_19973,N_18405,N_18607);
nand U19974 (N_19974,N_18216,N_18829);
nand U19975 (N_19975,N_18664,N_18564);
or U19976 (N_19976,N_18285,N_18677);
or U19977 (N_19977,N_18308,N_18752);
nor U19978 (N_19978,N_18148,N_18998);
and U19979 (N_19979,N_18123,N_18840);
or U19980 (N_19980,N_18027,N_18034);
nor U19981 (N_19981,N_18126,N_18749);
nand U19982 (N_19982,N_18301,N_18522);
or U19983 (N_19983,N_18697,N_18884);
nand U19984 (N_19984,N_18845,N_18800);
or U19985 (N_19985,N_18206,N_18683);
or U19986 (N_19986,N_18566,N_18381);
or U19987 (N_19987,N_18769,N_18064);
nand U19988 (N_19988,N_18991,N_18133);
and U19989 (N_19989,N_18319,N_18589);
nand U19990 (N_19990,N_18088,N_18365);
nor U19991 (N_19991,N_18282,N_18114);
nand U19992 (N_19992,N_18791,N_18755);
nand U19993 (N_19993,N_18663,N_18803);
nor U19994 (N_19994,N_18973,N_18129);
and U19995 (N_19995,N_18793,N_18065);
xnor U19996 (N_19996,N_18797,N_18514);
or U19997 (N_19997,N_18293,N_18339);
or U19998 (N_19998,N_18479,N_18804);
xnor U19999 (N_19999,N_18601,N_18369);
or UO_0 (O_0,N_19466,N_19706);
xor UO_1 (O_1,N_19389,N_19935);
nor UO_2 (O_2,N_19863,N_19021);
or UO_3 (O_3,N_19836,N_19397);
nand UO_4 (O_4,N_19536,N_19552);
nor UO_5 (O_5,N_19481,N_19001);
nor UO_6 (O_6,N_19516,N_19338);
nand UO_7 (O_7,N_19562,N_19968);
nor UO_8 (O_8,N_19175,N_19460);
nor UO_9 (O_9,N_19344,N_19554);
and UO_10 (O_10,N_19928,N_19019);
or UO_11 (O_11,N_19447,N_19665);
nand UO_12 (O_12,N_19709,N_19921);
or UO_13 (O_13,N_19699,N_19680);
xnor UO_14 (O_14,N_19085,N_19559);
nor UO_15 (O_15,N_19845,N_19158);
and UO_16 (O_16,N_19905,N_19975);
and UO_17 (O_17,N_19463,N_19683);
xnor UO_18 (O_18,N_19764,N_19022);
and UO_19 (O_19,N_19452,N_19999);
xnor UO_20 (O_20,N_19118,N_19633);
or UO_21 (O_21,N_19780,N_19626);
xnor UO_22 (O_22,N_19675,N_19396);
nor UO_23 (O_23,N_19597,N_19588);
nor UO_24 (O_24,N_19926,N_19471);
or UO_25 (O_25,N_19223,N_19601);
nor UO_26 (O_26,N_19914,N_19939);
or UO_27 (O_27,N_19393,N_19087);
nor UO_28 (O_28,N_19334,N_19268);
nand UO_29 (O_29,N_19897,N_19073);
nand UO_30 (O_30,N_19607,N_19574);
nor UO_31 (O_31,N_19482,N_19029);
or UO_32 (O_32,N_19809,N_19537);
and UO_33 (O_33,N_19840,N_19095);
nand UO_34 (O_34,N_19216,N_19962);
nand UO_35 (O_35,N_19341,N_19711);
or UO_36 (O_36,N_19644,N_19464);
nor UO_37 (O_37,N_19350,N_19685);
nand UO_38 (O_38,N_19070,N_19079);
nor UO_39 (O_39,N_19708,N_19982);
and UO_40 (O_40,N_19589,N_19099);
or UO_41 (O_41,N_19187,N_19220);
or UO_42 (O_42,N_19412,N_19714);
nand UO_43 (O_43,N_19960,N_19547);
or UO_44 (O_44,N_19732,N_19953);
and UO_45 (O_45,N_19760,N_19369);
nand UO_46 (O_46,N_19852,N_19144);
nand UO_47 (O_47,N_19787,N_19814);
or UO_48 (O_48,N_19386,N_19376);
nand UO_49 (O_49,N_19240,N_19703);
nand UO_50 (O_50,N_19956,N_19077);
and UO_51 (O_51,N_19600,N_19235);
and UO_52 (O_52,N_19662,N_19151);
xor UO_53 (O_53,N_19720,N_19551);
nand UO_54 (O_54,N_19372,N_19180);
nand UO_55 (O_55,N_19194,N_19045);
nand UO_56 (O_56,N_19735,N_19571);
or UO_57 (O_57,N_19289,N_19617);
xnor UO_58 (O_58,N_19632,N_19034);
nand UO_59 (O_59,N_19147,N_19170);
and UO_60 (O_60,N_19434,N_19692);
or UO_61 (O_61,N_19278,N_19459);
nor UO_62 (O_62,N_19865,N_19731);
nor UO_63 (O_63,N_19918,N_19239);
nor UO_64 (O_64,N_19517,N_19518);
and UO_65 (O_65,N_19005,N_19741);
or UO_66 (O_66,N_19707,N_19855);
and UO_67 (O_67,N_19477,N_19440);
or UO_68 (O_68,N_19391,N_19217);
xnor UO_69 (O_69,N_19721,N_19702);
or UO_70 (O_70,N_19909,N_19371);
or UO_71 (O_71,N_19544,N_19945);
and UO_72 (O_72,N_19587,N_19647);
or UO_73 (O_73,N_19538,N_19724);
or UO_74 (O_74,N_19184,N_19990);
or UO_75 (O_75,N_19103,N_19263);
and UO_76 (O_76,N_19530,N_19322);
nand UO_77 (O_77,N_19567,N_19590);
nand UO_78 (O_78,N_19432,N_19284);
nor UO_79 (O_79,N_19039,N_19564);
or UO_80 (O_80,N_19867,N_19832);
xnor UO_81 (O_81,N_19546,N_19943);
nor UO_82 (O_82,N_19745,N_19690);
nor UO_83 (O_83,N_19718,N_19541);
nand UO_84 (O_84,N_19221,N_19660);
nand UO_85 (O_85,N_19676,N_19456);
nand UO_86 (O_86,N_19385,N_19575);
and UO_87 (O_87,N_19249,N_19468);
and UO_88 (O_88,N_19024,N_19779);
or UO_89 (O_89,N_19006,N_19861);
or UO_90 (O_90,N_19150,N_19295);
nor UO_91 (O_91,N_19382,N_19038);
and UO_92 (O_92,N_19752,N_19992);
or UO_93 (O_93,N_19238,N_19788);
nand UO_94 (O_94,N_19354,N_19258);
nor UO_95 (O_95,N_19831,N_19766);
nand UO_96 (O_96,N_19869,N_19756);
nand UO_97 (O_97,N_19816,N_19879);
nor UO_98 (O_98,N_19302,N_19612);
xnor UO_99 (O_99,N_19859,N_19112);
xor UO_100 (O_100,N_19958,N_19729);
and UO_101 (O_101,N_19271,N_19673);
or UO_102 (O_102,N_19117,N_19494);
nand UO_103 (O_103,N_19976,N_19124);
and UO_104 (O_104,N_19066,N_19230);
or UO_105 (O_105,N_19842,N_19507);
nor UO_106 (O_106,N_19234,N_19134);
or UO_107 (O_107,N_19149,N_19098);
nand UO_108 (O_108,N_19667,N_19421);
or UO_109 (O_109,N_19018,N_19654);
nor UO_110 (O_110,N_19072,N_19603);
xor UO_111 (O_111,N_19093,N_19555);
and UO_112 (O_112,N_19485,N_19512);
and UO_113 (O_113,N_19204,N_19428);
or UO_114 (O_114,N_19191,N_19920);
nor UO_115 (O_115,N_19650,N_19782);
or UO_116 (O_116,N_19496,N_19671);
nor UO_117 (O_117,N_19586,N_19986);
or UO_118 (O_118,N_19651,N_19339);
xnor UO_119 (O_119,N_19717,N_19321);
nor UO_120 (O_120,N_19435,N_19980);
nand UO_121 (O_121,N_19267,N_19137);
nand UO_122 (O_122,N_19044,N_19243);
nand UO_123 (O_123,N_19715,N_19854);
nor UO_124 (O_124,N_19798,N_19102);
or UO_125 (O_125,N_19674,N_19880);
or UO_126 (O_126,N_19526,N_19261);
nor UO_127 (O_127,N_19153,N_19778);
or UO_128 (O_128,N_19264,N_19462);
nor UO_129 (O_129,N_19876,N_19944);
nand UO_130 (O_130,N_19989,N_19241);
and UO_131 (O_131,N_19378,N_19292);
nor UO_132 (O_132,N_19535,N_19672);
and UO_133 (O_133,N_19197,N_19682);
xor UO_134 (O_134,N_19661,N_19819);
or UO_135 (O_135,N_19226,N_19057);
xnor UO_136 (O_136,N_19110,N_19067);
and UO_137 (O_137,N_19540,N_19236);
nand UO_138 (O_138,N_19668,N_19425);
xnor UO_139 (O_139,N_19196,N_19262);
xor UO_140 (O_140,N_19046,N_19490);
or UO_141 (O_141,N_19606,N_19542);
and UO_142 (O_142,N_19367,N_19154);
nor UO_143 (O_143,N_19366,N_19701);
nor UO_144 (O_144,N_19027,N_19207);
nor UO_145 (O_145,N_19188,N_19282);
nor UO_146 (O_146,N_19395,N_19993);
nand UO_147 (O_147,N_19892,N_19767);
or UO_148 (O_148,N_19037,N_19895);
and UO_149 (O_149,N_19898,N_19211);
or UO_150 (O_150,N_19251,N_19276);
xor UO_151 (O_151,N_19844,N_19529);
or UO_152 (O_152,N_19377,N_19792);
or UO_153 (O_153,N_19758,N_19763);
or UO_154 (O_154,N_19624,N_19791);
and UO_155 (O_155,N_19915,N_19585);
and UO_156 (O_156,N_19062,N_19345);
nor UO_157 (O_157,N_19418,N_19069);
nand UO_158 (O_158,N_19417,N_19550);
nor UO_159 (O_159,N_19116,N_19531);
nand UO_160 (O_160,N_19437,N_19646);
nor UO_161 (O_161,N_19265,N_19352);
or UO_162 (O_162,N_19141,N_19618);
or UO_163 (O_163,N_19470,N_19358);
or UO_164 (O_164,N_19314,N_19998);
nor UO_165 (O_165,N_19594,N_19402);
nand UO_166 (O_166,N_19736,N_19145);
or UO_167 (O_167,N_19298,N_19817);
nor UO_168 (O_168,N_19679,N_19948);
nand UO_169 (O_169,N_19598,N_19380);
and UO_170 (O_170,N_19873,N_19957);
and UO_171 (O_171,N_19076,N_19955);
xnor UO_172 (O_172,N_19625,N_19894);
or UO_173 (O_173,N_19131,N_19013);
xnor UO_174 (O_174,N_19088,N_19139);
and UO_175 (O_175,N_19521,N_19950);
and UO_176 (O_176,N_19055,N_19566);
or UO_177 (O_177,N_19363,N_19784);
or UO_178 (O_178,N_19242,N_19419);
nand UO_179 (O_179,N_19457,N_19669);
nor UO_180 (O_180,N_19113,N_19813);
nor UO_181 (O_181,N_19106,N_19010);
and UO_182 (O_182,N_19203,N_19925);
and UO_183 (O_183,N_19743,N_19441);
and UO_184 (O_184,N_19253,N_19337);
and UO_185 (O_185,N_19983,N_19476);
or UO_186 (O_186,N_19886,N_19047);
xor UO_187 (O_187,N_19907,N_19004);
or UO_188 (O_188,N_19882,N_19506);
nor UO_189 (O_189,N_19874,N_19599);
nor UO_190 (O_190,N_19696,N_19722);
nor UO_191 (O_191,N_19871,N_19532);
xnor UO_192 (O_192,N_19759,N_19580);
nand UO_193 (O_193,N_19578,N_19190);
or UO_194 (O_194,N_19681,N_19610);
nor UO_195 (O_195,N_19157,N_19308);
nor UO_196 (O_196,N_19080,N_19299);
or UO_197 (O_197,N_19237,N_19210);
and UO_198 (O_198,N_19539,N_19591);
nand UO_199 (O_199,N_19163,N_19212);
nor UO_200 (O_200,N_19218,N_19307);
nand UO_201 (O_201,N_19431,N_19052);
nand UO_202 (O_202,N_19115,N_19877);
nand UO_203 (O_203,N_19105,N_19275);
or UO_204 (O_204,N_19138,N_19866);
and UO_205 (O_205,N_19257,N_19858);
and UO_206 (O_206,N_19781,N_19405);
and UO_207 (O_207,N_19269,N_19123);
nor UO_208 (O_208,N_19177,N_19033);
and UO_209 (O_209,N_19850,N_19408);
nor UO_210 (O_210,N_19558,N_19804);
nor UO_211 (O_211,N_19728,N_19427);
nor UO_212 (O_212,N_19611,N_19572);
and UO_213 (O_213,N_19126,N_19359);
nor UO_214 (O_214,N_19186,N_19753);
nor UO_215 (O_215,N_19403,N_19515);
and UO_216 (O_216,N_19082,N_19560);
nor UO_217 (O_217,N_19061,N_19719);
and UO_218 (O_218,N_19812,N_19991);
nor UO_219 (O_219,N_19426,N_19383);
nor UO_220 (O_220,N_19347,N_19981);
nor UO_221 (O_221,N_19751,N_19056);
and UO_222 (O_222,N_19520,N_19996);
and UO_223 (O_223,N_19195,N_19014);
nand UO_224 (O_224,N_19762,N_19007);
nor UO_225 (O_225,N_19486,N_19978);
and UO_226 (O_226,N_19899,N_19750);
nand UO_227 (O_227,N_19246,N_19635);
and UO_228 (O_228,N_19274,N_19636);
nor UO_229 (O_229,N_19849,N_19379);
or UO_230 (O_230,N_19505,N_19285);
or UO_231 (O_231,N_19213,N_19342);
xor UO_232 (O_232,N_19648,N_19390);
xnor UO_233 (O_233,N_19484,N_19025);
or UO_234 (O_234,N_19255,N_19162);
nor UO_235 (O_235,N_19997,N_19492);
nor UO_236 (O_236,N_19748,N_19155);
and UO_237 (O_237,N_19630,N_19890);
nand UO_238 (O_238,N_19400,N_19670);
nor UO_239 (O_239,N_19838,N_19906);
and UO_240 (O_240,N_19091,N_19872);
and UO_241 (O_241,N_19577,N_19775);
or UO_242 (O_242,N_19266,N_19569);
xor UO_243 (O_243,N_19937,N_19399);
nor UO_244 (O_244,N_19181,N_19684);
nor UO_245 (O_245,N_19313,N_19938);
and UO_246 (O_246,N_19444,N_19465);
nand UO_247 (O_247,N_19208,N_19286);
nor UO_248 (O_248,N_19805,N_19451);
and UO_249 (O_249,N_19416,N_19710);
nor UO_250 (O_250,N_19161,N_19356);
nand UO_251 (O_251,N_19628,N_19678);
nor UO_252 (O_252,N_19726,N_19165);
or UO_253 (O_253,N_19026,N_19754);
nor UO_254 (O_254,N_19023,N_19772);
or UO_255 (O_255,N_19747,N_19398);
and UO_256 (O_256,N_19202,N_19830);
and UO_257 (O_257,N_19705,N_19988);
and UO_258 (O_258,N_19483,N_19723);
nor UO_259 (O_259,N_19443,N_19972);
nor UO_260 (O_260,N_19458,N_19868);
nor UO_261 (O_261,N_19401,N_19254);
nand UO_262 (O_262,N_19800,N_19891);
nor UO_263 (O_263,N_19064,N_19900);
or UO_264 (O_264,N_19222,N_19534);
nand UO_265 (O_265,N_19946,N_19525);
and UO_266 (O_266,N_19214,N_19329);
nor UO_267 (O_267,N_19473,N_19697);
nor UO_268 (O_268,N_19835,N_19060);
or UO_269 (O_269,N_19016,N_19498);
nor UO_270 (O_270,N_19640,N_19801);
and UO_271 (O_271,N_19545,N_19936);
nor UO_272 (O_272,N_19059,N_19063);
and UO_273 (O_273,N_19104,N_19793);
and UO_274 (O_274,N_19727,N_19040);
nor UO_275 (O_275,N_19666,N_19910);
nand UO_276 (O_276,N_19058,N_19929);
xor UO_277 (O_277,N_19325,N_19826);
and UO_278 (O_278,N_19248,N_19769);
and UO_279 (O_279,N_19164,N_19965);
nand UO_280 (O_280,N_19084,N_19689);
or UO_281 (O_281,N_19821,N_19698);
and UO_282 (O_282,N_19415,N_19078);
or UO_283 (O_283,N_19200,N_19818);
nand UO_284 (O_284,N_19663,N_19129);
or UO_285 (O_285,N_19595,N_19883);
nor UO_286 (O_286,N_19148,N_19947);
or UO_287 (O_287,N_19449,N_19009);
nand UO_288 (O_288,N_19942,N_19889);
or UO_289 (O_289,N_19771,N_19049);
or UO_290 (O_290,N_19912,N_19120);
xnor UO_291 (O_291,N_19933,N_19857);
nor UO_292 (O_292,N_19107,N_19686);
nand UO_293 (O_293,N_19357,N_19119);
and UO_294 (O_294,N_19785,N_19041);
and UO_295 (O_295,N_19613,N_19035);
or UO_296 (O_296,N_19198,N_19904);
or UO_297 (O_297,N_19343,N_19192);
or UO_298 (O_298,N_19846,N_19453);
xnor UO_299 (O_299,N_19738,N_19860);
nand UO_300 (O_300,N_19959,N_19260);
xor UO_301 (O_301,N_19627,N_19837);
or UO_302 (O_302,N_19475,N_19407);
xor UO_303 (O_303,N_19908,N_19290);
and UO_304 (O_304,N_19533,N_19584);
xor UO_305 (O_305,N_19768,N_19178);
xor UO_306 (O_306,N_19827,N_19114);
and UO_307 (O_307,N_19713,N_19469);
or UO_308 (O_308,N_19365,N_19108);
nand UO_309 (O_309,N_19851,N_19963);
xor UO_310 (O_310,N_19664,N_19461);
or UO_311 (O_311,N_19050,N_19259);
or UO_312 (O_312,N_19799,N_19310);
or UO_313 (O_313,N_19966,N_19096);
and UO_314 (O_314,N_19430,N_19183);
nand UO_315 (O_315,N_19450,N_19159);
nand UO_316 (O_316,N_19319,N_19903);
and UO_317 (O_317,N_19615,N_19878);
nor UO_318 (O_318,N_19495,N_19323);
xnor UO_319 (O_319,N_19374,N_19875);
nor UO_320 (O_320,N_19896,N_19094);
and UO_321 (O_321,N_19169,N_19219);
nand UO_322 (O_322,N_19987,N_19229);
nand UO_323 (O_323,N_19881,N_19224);
or UO_324 (O_324,N_19524,N_19362);
nor UO_325 (O_325,N_19620,N_19433);
nor UO_326 (O_326,N_19796,N_19749);
or UO_327 (O_327,N_19740,N_19283);
nand UO_328 (O_328,N_19609,N_19130);
and UO_329 (O_329,N_19328,N_19065);
nand UO_330 (O_330,N_19977,N_19913);
and UO_331 (O_331,N_19641,N_19927);
xor UO_332 (O_332,N_19100,N_19304);
nand UO_333 (O_333,N_19649,N_19316);
and UO_334 (O_334,N_19841,N_19244);
or UO_335 (O_335,N_19279,N_19333);
and UO_336 (O_336,N_19300,N_19227);
or UO_337 (O_337,N_19967,N_19193);
nand UO_338 (O_338,N_19324,N_19331);
nor UO_339 (O_339,N_19634,N_19346);
nor UO_340 (O_340,N_19971,N_19215);
nor UO_341 (O_341,N_19409,N_19504);
nand UO_342 (O_342,N_19658,N_19291);
nor UO_343 (O_343,N_19135,N_19786);
nand UO_344 (O_344,N_19730,N_19422);
xnor UO_345 (O_345,N_19795,N_19949);
nand UO_346 (O_346,N_19491,N_19637);
and UO_347 (O_347,N_19127,N_19081);
nor UO_348 (O_348,N_19783,N_19445);
xor UO_349 (O_349,N_19125,N_19514);
or UO_350 (O_350,N_19931,N_19870);
nor UO_351 (O_351,N_19653,N_19593);
nand UO_352 (O_352,N_19802,N_19036);
nand UO_353 (O_353,N_19327,N_19561);
nor UO_354 (O_354,N_19694,N_19774);
nand UO_355 (O_355,N_19487,N_19790);
nor UO_356 (O_356,N_19737,N_19543);
nand UO_357 (O_357,N_19002,N_19406);
and UO_358 (O_358,N_19152,N_19509);
or UO_359 (O_359,N_19493,N_19765);
nand UO_360 (O_360,N_19757,N_19582);
nor UO_361 (O_361,N_19773,N_19031);
xor UO_362 (O_362,N_19296,N_19761);
and UO_363 (O_363,N_19326,N_19631);
or UO_364 (O_364,N_19508,N_19312);
nor UO_365 (O_365,N_19233,N_19605);
and UO_366 (O_366,N_19133,N_19250);
nand UO_367 (O_367,N_19604,N_19053);
xnor UO_368 (O_368,N_19252,N_19008);
and UO_369 (O_369,N_19777,N_19888);
or UO_370 (O_370,N_19042,N_19810);
nor UO_371 (O_371,N_19472,N_19205);
nand UO_372 (O_372,N_19716,N_19825);
nor UO_373 (O_373,N_19951,N_19501);
nand UO_374 (O_374,N_19351,N_19166);
or UO_375 (O_375,N_19317,N_19581);
or UO_376 (O_376,N_19924,N_19528);
and UO_377 (O_377,N_19964,N_19335);
or UO_378 (O_378,N_19301,N_19413);
or UO_379 (O_379,N_19423,N_19862);
or UO_380 (O_380,N_19281,N_19442);
nand UO_381 (O_381,N_19922,N_19160);
and UO_382 (O_382,N_19712,N_19232);
nand UO_383 (O_383,N_19639,N_19392);
nor UO_384 (O_384,N_19424,N_19746);
and UO_385 (O_385,N_19287,N_19853);
and UO_386 (O_386,N_19048,N_19370);
nor UO_387 (O_387,N_19693,N_19985);
xnor UO_388 (O_388,N_19020,N_19655);
and UO_389 (O_389,N_19885,N_19622);
nor UO_390 (O_390,N_19293,N_19368);
nor UO_391 (O_391,N_19003,N_19388);
and UO_392 (O_392,N_19619,N_19438);
nor UO_393 (O_393,N_19340,N_19090);
or UO_394 (O_394,N_19256,N_19930);
nor UO_395 (O_395,N_19375,N_19101);
nand UO_396 (O_396,N_19051,N_19122);
nor UO_397 (O_397,N_19332,N_19902);
or UO_398 (O_398,N_19303,N_19974);
and UO_399 (O_399,N_19309,N_19028);
nor UO_400 (O_400,N_19995,N_19820);
nor UO_401 (O_401,N_19136,N_19206);
nor UO_402 (O_402,N_19373,N_19277);
and UO_403 (O_403,N_19823,N_19923);
or UO_404 (O_404,N_19414,N_19502);
nand UO_405 (O_405,N_19270,N_19436);
and UO_406 (O_406,N_19602,N_19563);
nand UO_407 (O_407,N_19455,N_19742);
or UO_408 (O_408,N_19807,N_19228);
nand UO_409 (O_409,N_19306,N_19527);
nand UO_410 (O_410,N_19755,N_19075);
nand UO_411 (O_411,N_19856,N_19553);
and UO_412 (O_412,N_19089,N_19608);
xor UO_413 (O_413,N_19806,N_19847);
or UO_414 (O_414,N_19803,N_19596);
or UO_415 (O_415,N_19522,N_19932);
xnor UO_416 (O_416,N_19272,N_19828);
or UO_417 (O_417,N_19348,N_19556);
or UO_418 (O_418,N_19794,N_19111);
and UO_419 (O_419,N_19349,N_19305);
or UO_420 (O_420,N_19511,N_19488);
xor UO_421 (O_421,N_19688,N_19704);
xor UO_422 (O_422,N_19245,N_19074);
xor UO_423 (O_423,N_19012,N_19086);
or UO_424 (O_424,N_19973,N_19592);
and UO_425 (O_425,N_19848,N_19174);
and UO_426 (O_426,N_19623,N_19071);
nor UO_427 (O_427,N_19404,N_19916);
nand UO_428 (O_428,N_19361,N_19815);
nor UO_429 (O_429,N_19645,N_19387);
and UO_430 (O_430,N_19568,N_19725);
or UO_431 (O_431,N_19201,N_19961);
nand UO_432 (O_432,N_19017,N_19140);
or UO_433 (O_433,N_19011,N_19969);
nand UO_434 (O_434,N_19043,N_19565);
nor UO_435 (O_435,N_19573,N_19616);
or UO_436 (O_436,N_19934,N_19231);
nor UO_437 (O_437,N_19513,N_19700);
and UO_438 (O_438,N_19739,N_19979);
xor UO_439 (O_439,N_19919,N_19384);
and UO_440 (O_440,N_19420,N_19173);
or UO_441 (O_441,N_19032,N_19311);
nand UO_442 (O_442,N_19657,N_19189);
and UO_443 (O_443,N_19887,N_19143);
or UO_444 (O_444,N_19901,N_19132);
nor UO_445 (O_445,N_19503,N_19288);
nor UO_446 (O_446,N_19811,N_19410);
or UO_447 (O_447,N_19621,N_19315);
nor UO_448 (O_448,N_19360,N_19294);
nand UO_449 (O_449,N_19652,N_19179);
nand UO_450 (O_450,N_19121,N_19446);
or UO_451 (O_451,N_19557,N_19097);
nand UO_452 (O_452,N_19954,N_19941);
xor UO_453 (O_453,N_19054,N_19583);
or UO_454 (O_454,N_19172,N_19695);
xor UO_455 (O_455,N_19834,N_19744);
and UO_456 (O_456,N_19474,N_19917);
nor UO_457 (O_457,N_19579,N_19394);
nand UO_458 (O_458,N_19970,N_19911);
nand UO_459 (O_459,N_19364,N_19994);
nor UO_460 (O_460,N_19167,N_19355);
nor UO_461 (O_461,N_19448,N_19691);
or UO_462 (O_462,N_19297,N_19952);
nand UO_463 (O_463,N_19770,N_19336);
nor UO_464 (O_464,N_19893,N_19176);
and UO_465 (O_465,N_19318,N_19185);
or UO_466 (O_466,N_19411,N_19822);
or UO_467 (O_467,N_19128,N_19109);
or UO_468 (O_468,N_19797,N_19734);
and UO_469 (O_469,N_19168,N_19500);
or UO_470 (O_470,N_19156,N_19940);
nand UO_471 (O_471,N_19642,N_19146);
xor UO_472 (O_472,N_19523,N_19677);
or UO_473 (O_473,N_19864,N_19499);
or UO_474 (O_474,N_19643,N_19068);
xor UO_475 (O_475,N_19353,N_19199);
and UO_476 (O_476,N_19629,N_19548);
nand UO_477 (O_477,N_19280,N_19776);
or UO_478 (O_478,N_19083,N_19000);
nor UO_479 (O_479,N_19171,N_19439);
nor UO_480 (O_480,N_19549,N_19570);
nand UO_481 (O_481,N_19519,N_19454);
and UO_482 (O_482,N_19142,N_19656);
or UO_483 (O_483,N_19479,N_19467);
nand UO_484 (O_484,N_19984,N_19320);
nor UO_485 (O_485,N_19478,N_19480);
nor UO_486 (O_486,N_19638,N_19687);
or UO_487 (O_487,N_19733,N_19182);
and UO_488 (O_488,N_19659,N_19833);
nor UO_489 (O_489,N_19015,N_19829);
nor UO_490 (O_490,N_19030,N_19884);
nor UO_491 (O_491,N_19576,N_19839);
nand UO_492 (O_492,N_19843,N_19510);
nor UO_493 (O_493,N_19330,N_19497);
or UO_494 (O_494,N_19614,N_19092);
and UO_495 (O_495,N_19824,N_19429);
nor UO_496 (O_496,N_19225,N_19209);
and UO_497 (O_497,N_19789,N_19808);
nor UO_498 (O_498,N_19273,N_19381);
or UO_499 (O_499,N_19489,N_19247);
nand UO_500 (O_500,N_19286,N_19235);
and UO_501 (O_501,N_19946,N_19643);
nand UO_502 (O_502,N_19094,N_19145);
or UO_503 (O_503,N_19842,N_19906);
nor UO_504 (O_504,N_19797,N_19386);
nand UO_505 (O_505,N_19497,N_19316);
nor UO_506 (O_506,N_19147,N_19723);
or UO_507 (O_507,N_19804,N_19763);
xor UO_508 (O_508,N_19174,N_19148);
nor UO_509 (O_509,N_19952,N_19919);
nand UO_510 (O_510,N_19904,N_19249);
and UO_511 (O_511,N_19994,N_19708);
xor UO_512 (O_512,N_19915,N_19924);
or UO_513 (O_513,N_19654,N_19069);
nor UO_514 (O_514,N_19322,N_19902);
or UO_515 (O_515,N_19399,N_19916);
nor UO_516 (O_516,N_19147,N_19656);
and UO_517 (O_517,N_19502,N_19059);
and UO_518 (O_518,N_19236,N_19361);
and UO_519 (O_519,N_19268,N_19584);
nor UO_520 (O_520,N_19466,N_19872);
xor UO_521 (O_521,N_19093,N_19338);
or UO_522 (O_522,N_19103,N_19210);
and UO_523 (O_523,N_19750,N_19481);
or UO_524 (O_524,N_19286,N_19787);
or UO_525 (O_525,N_19356,N_19920);
nor UO_526 (O_526,N_19885,N_19833);
or UO_527 (O_527,N_19512,N_19349);
and UO_528 (O_528,N_19665,N_19583);
nor UO_529 (O_529,N_19234,N_19915);
or UO_530 (O_530,N_19688,N_19056);
nand UO_531 (O_531,N_19840,N_19259);
or UO_532 (O_532,N_19954,N_19872);
nand UO_533 (O_533,N_19353,N_19610);
or UO_534 (O_534,N_19835,N_19716);
and UO_535 (O_535,N_19739,N_19062);
or UO_536 (O_536,N_19860,N_19757);
or UO_537 (O_537,N_19134,N_19566);
or UO_538 (O_538,N_19347,N_19784);
or UO_539 (O_539,N_19337,N_19857);
and UO_540 (O_540,N_19372,N_19833);
or UO_541 (O_541,N_19874,N_19175);
nor UO_542 (O_542,N_19559,N_19449);
xor UO_543 (O_543,N_19172,N_19876);
or UO_544 (O_544,N_19472,N_19036);
or UO_545 (O_545,N_19142,N_19186);
or UO_546 (O_546,N_19509,N_19820);
or UO_547 (O_547,N_19988,N_19210);
nand UO_548 (O_548,N_19284,N_19309);
or UO_549 (O_549,N_19194,N_19889);
and UO_550 (O_550,N_19679,N_19530);
or UO_551 (O_551,N_19942,N_19575);
xnor UO_552 (O_552,N_19973,N_19752);
or UO_553 (O_553,N_19046,N_19507);
and UO_554 (O_554,N_19516,N_19520);
and UO_555 (O_555,N_19408,N_19388);
nand UO_556 (O_556,N_19364,N_19241);
nand UO_557 (O_557,N_19348,N_19077);
nand UO_558 (O_558,N_19597,N_19494);
nand UO_559 (O_559,N_19912,N_19237);
and UO_560 (O_560,N_19339,N_19850);
or UO_561 (O_561,N_19339,N_19854);
xnor UO_562 (O_562,N_19496,N_19343);
or UO_563 (O_563,N_19605,N_19421);
and UO_564 (O_564,N_19626,N_19611);
nor UO_565 (O_565,N_19550,N_19927);
nor UO_566 (O_566,N_19651,N_19136);
and UO_567 (O_567,N_19410,N_19140);
or UO_568 (O_568,N_19511,N_19751);
and UO_569 (O_569,N_19064,N_19467);
nor UO_570 (O_570,N_19580,N_19092);
nor UO_571 (O_571,N_19287,N_19122);
and UO_572 (O_572,N_19238,N_19054);
nor UO_573 (O_573,N_19753,N_19617);
xor UO_574 (O_574,N_19286,N_19733);
nor UO_575 (O_575,N_19751,N_19789);
nor UO_576 (O_576,N_19907,N_19680);
nor UO_577 (O_577,N_19581,N_19822);
and UO_578 (O_578,N_19328,N_19165);
or UO_579 (O_579,N_19466,N_19633);
nand UO_580 (O_580,N_19941,N_19025);
nand UO_581 (O_581,N_19762,N_19312);
and UO_582 (O_582,N_19470,N_19969);
and UO_583 (O_583,N_19866,N_19790);
nor UO_584 (O_584,N_19987,N_19352);
nor UO_585 (O_585,N_19632,N_19151);
or UO_586 (O_586,N_19484,N_19886);
nand UO_587 (O_587,N_19578,N_19154);
and UO_588 (O_588,N_19023,N_19176);
nor UO_589 (O_589,N_19042,N_19460);
and UO_590 (O_590,N_19550,N_19816);
nor UO_591 (O_591,N_19799,N_19633);
nand UO_592 (O_592,N_19320,N_19756);
nand UO_593 (O_593,N_19367,N_19939);
nor UO_594 (O_594,N_19886,N_19307);
nor UO_595 (O_595,N_19889,N_19617);
nor UO_596 (O_596,N_19392,N_19753);
nor UO_597 (O_597,N_19542,N_19567);
or UO_598 (O_598,N_19312,N_19817);
nor UO_599 (O_599,N_19831,N_19787);
or UO_600 (O_600,N_19710,N_19204);
nor UO_601 (O_601,N_19292,N_19344);
nor UO_602 (O_602,N_19455,N_19143);
or UO_603 (O_603,N_19918,N_19905);
nand UO_604 (O_604,N_19414,N_19626);
nor UO_605 (O_605,N_19946,N_19806);
and UO_606 (O_606,N_19863,N_19967);
and UO_607 (O_607,N_19200,N_19151);
or UO_608 (O_608,N_19472,N_19965);
and UO_609 (O_609,N_19533,N_19936);
nand UO_610 (O_610,N_19571,N_19608);
or UO_611 (O_611,N_19105,N_19086);
nand UO_612 (O_612,N_19456,N_19284);
or UO_613 (O_613,N_19579,N_19776);
and UO_614 (O_614,N_19079,N_19010);
xor UO_615 (O_615,N_19816,N_19220);
and UO_616 (O_616,N_19021,N_19746);
and UO_617 (O_617,N_19416,N_19326);
nor UO_618 (O_618,N_19351,N_19721);
nor UO_619 (O_619,N_19909,N_19773);
or UO_620 (O_620,N_19353,N_19670);
nand UO_621 (O_621,N_19525,N_19709);
nor UO_622 (O_622,N_19070,N_19307);
nor UO_623 (O_623,N_19746,N_19677);
or UO_624 (O_624,N_19716,N_19102);
xor UO_625 (O_625,N_19274,N_19773);
nor UO_626 (O_626,N_19290,N_19916);
nor UO_627 (O_627,N_19718,N_19599);
and UO_628 (O_628,N_19702,N_19680);
and UO_629 (O_629,N_19611,N_19028);
nor UO_630 (O_630,N_19637,N_19106);
nor UO_631 (O_631,N_19264,N_19864);
xnor UO_632 (O_632,N_19125,N_19864);
or UO_633 (O_633,N_19428,N_19560);
or UO_634 (O_634,N_19994,N_19488);
nand UO_635 (O_635,N_19486,N_19887);
nor UO_636 (O_636,N_19209,N_19569);
nor UO_637 (O_637,N_19085,N_19934);
nand UO_638 (O_638,N_19479,N_19054);
and UO_639 (O_639,N_19830,N_19684);
nor UO_640 (O_640,N_19148,N_19424);
nand UO_641 (O_641,N_19439,N_19886);
nor UO_642 (O_642,N_19472,N_19428);
or UO_643 (O_643,N_19042,N_19103);
nand UO_644 (O_644,N_19306,N_19270);
nor UO_645 (O_645,N_19930,N_19054);
nor UO_646 (O_646,N_19184,N_19236);
and UO_647 (O_647,N_19307,N_19602);
or UO_648 (O_648,N_19926,N_19385);
xnor UO_649 (O_649,N_19848,N_19724);
nor UO_650 (O_650,N_19520,N_19538);
or UO_651 (O_651,N_19341,N_19139);
nor UO_652 (O_652,N_19219,N_19822);
and UO_653 (O_653,N_19187,N_19788);
and UO_654 (O_654,N_19755,N_19239);
or UO_655 (O_655,N_19345,N_19011);
nor UO_656 (O_656,N_19356,N_19777);
or UO_657 (O_657,N_19818,N_19210);
or UO_658 (O_658,N_19049,N_19556);
and UO_659 (O_659,N_19468,N_19075);
nor UO_660 (O_660,N_19795,N_19900);
nand UO_661 (O_661,N_19151,N_19207);
or UO_662 (O_662,N_19555,N_19720);
nand UO_663 (O_663,N_19465,N_19359);
and UO_664 (O_664,N_19953,N_19089);
nand UO_665 (O_665,N_19618,N_19799);
xor UO_666 (O_666,N_19056,N_19112);
nand UO_667 (O_667,N_19980,N_19601);
nor UO_668 (O_668,N_19835,N_19796);
or UO_669 (O_669,N_19124,N_19470);
or UO_670 (O_670,N_19948,N_19999);
xnor UO_671 (O_671,N_19579,N_19852);
nor UO_672 (O_672,N_19729,N_19902);
and UO_673 (O_673,N_19558,N_19864);
nand UO_674 (O_674,N_19350,N_19405);
or UO_675 (O_675,N_19317,N_19135);
or UO_676 (O_676,N_19802,N_19268);
and UO_677 (O_677,N_19465,N_19413);
or UO_678 (O_678,N_19226,N_19291);
and UO_679 (O_679,N_19616,N_19065);
or UO_680 (O_680,N_19024,N_19762);
or UO_681 (O_681,N_19515,N_19116);
xnor UO_682 (O_682,N_19666,N_19870);
xor UO_683 (O_683,N_19884,N_19275);
and UO_684 (O_684,N_19000,N_19356);
xor UO_685 (O_685,N_19641,N_19113);
nor UO_686 (O_686,N_19706,N_19977);
nor UO_687 (O_687,N_19333,N_19039);
and UO_688 (O_688,N_19274,N_19520);
nand UO_689 (O_689,N_19187,N_19015);
and UO_690 (O_690,N_19539,N_19041);
xnor UO_691 (O_691,N_19228,N_19608);
nand UO_692 (O_692,N_19502,N_19461);
nand UO_693 (O_693,N_19691,N_19225);
and UO_694 (O_694,N_19459,N_19024);
nor UO_695 (O_695,N_19772,N_19074);
nor UO_696 (O_696,N_19088,N_19746);
or UO_697 (O_697,N_19122,N_19396);
nand UO_698 (O_698,N_19288,N_19859);
nand UO_699 (O_699,N_19308,N_19553);
and UO_700 (O_700,N_19293,N_19714);
or UO_701 (O_701,N_19542,N_19422);
and UO_702 (O_702,N_19527,N_19014);
or UO_703 (O_703,N_19467,N_19699);
or UO_704 (O_704,N_19338,N_19949);
and UO_705 (O_705,N_19256,N_19828);
nor UO_706 (O_706,N_19490,N_19400);
xor UO_707 (O_707,N_19234,N_19930);
and UO_708 (O_708,N_19542,N_19628);
nor UO_709 (O_709,N_19505,N_19265);
xnor UO_710 (O_710,N_19073,N_19754);
xor UO_711 (O_711,N_19373,N_19913);
and UO_712 (O_712,N_19334,N_19799);
nand UO_713 (O_713,N_19440,N_19262);
or UO_714 (O_714,N_19691,N_19903);
nor UO_715 (O_715,N_19248,N_19200);
and UO_716 (O_716,N_19784,N_19202);
nor UO_717 (O_717,N_19714,N_19049);
nand UO_718 (O_718,N_19865,N_19321);
nand UO_719 (O_719,N_19405,N_19340);
or UO_720 (O_720,N_19814,N_19587);
nor UO_721 (O_721,N_19750,N_19654);
nor UO_722 (O_722,N_19190,N_19437);
nor UO_723 (O_723,N_19607,N_19007);
nand UO_724 (O_724,N_19937,N_19098);
nor UO_725 (O_725,N_19419,N_19399);
or UO_726 (O_726,N_19159,N_19993);
or UO_727 (O_727,N_19732,N_19280);
nand UO_728 (O_728,N_19601,N_19940);
nor UO_729 (O_729,N_19054,N_19407);
xnor UO_730 (O_730,N_19207,N_19902);
and UO_731 (O_731,N_19851,N_19179);
and UO_732 (O_732,N_19002,N_19574);
and UO_733 (O_733,N_19633,N_19789);
nor UO_734 (O_734,N_19472,N_19020);
nor UO_735 (O_735,N_19070,N_19101);
or UO_736 (O_736,N_19843,N_19207);
nor UO_737 (O_737,N_19533,N_19506);
nand UO_738 (O_738,N_19845,N_19605);
nand UO_739 (O_739,N_19222,N_19647);
nor UO_740 (O_740,N_19553,N_19270);
nand UO_741 (O_741,N_19712,N_19955);
and UO_742 (O_742,N_19137,N_19224);
nor UO_743 (O_743,N_19563,N_19316);
xor UO_744 (O_744,N_19317,N_19128);
xor UO_745 (O_745,N_19095,N_19586);
and UO_746 (O_746,N_19056,N_19457);
nor UO_747 (O_747,N_19686,N_19452);
and UO_748 (O_748,N_19973,N_19136);
or UO_749 (O_749,N_19372,N_19877);
nor UO_750 (O_750,N_19536,N_19145);
nor UO_751 (O_751,N_19139,N_19170);
or UO_752 (O_752,N_19491,N_19006);
nand UO_753 (O_753,N_19687,N_19685);
nand UO_754 (O_754,N_19503,N_19565);
or UO_755 (O_755,N_19880,N_19815);
nor UO_756 (O_756,N_19488,N_19171);
nand UO_757 (O_757,N_19570,N_19935);
nor UO_758 (O_758,N_19294,N_19966);
nor UO_759 (O_759,N_19456,N_19696);
and UO_760 (O_760,N_19595,N_19089);
xnor UO_761 (O_761,N_19995,N_19122);
or UO_762 (O_762,N_19489,N_19271);
or UO_763 (O_763,N_19179,N_19253);
and UO_764 (O_764,N_19716,N_19894);
nand UO_765 (O_765,N_19834,N_19479);
xnor UO_766 (O_766,N_19813,N_19807);
or UO_767 (O_767,N_19500,N_19646);
nand UO_768 (O_768,N_19461,N_19251);
nand UO_769 (O_769,N_19988,N_19327);
nand UO_770 (O_770,N_19139,N_19269);
and UO_771 (O_771,N_19766,N_19309);
nor UO_772 (O_772,N_19828,N_19169);
nor UO_773 (O_773,N_19564,N_19698);
nor UO_774 (O_774,N_19394,N_19165);
nand UO_775 (O_775,N_19333,N_19497);
and UO_776 (O_776,N_19978,N_19412);
xor UO_777 (O_777,N_19321,N_19104);
nor UO_778 (O_778,N_19261,N_19126);
nand UO_779 (O_779,N_19144,N_19526);
and UO_780 (O_780,N_19909,N_19960);
or UO_781 (O_781,N_19958,N_19526);
nand UO_782 (O_782,N_19994,N_19715);
and UO_783 (O_783,N_19321,N_19921);
nand UO_784 (O_784,N_19260,N_19694);
nor UO_785 (O_785,N_19841,N_19202);
nand UO_786 (O_786,N_19331,N_19900);
and UO_787 (O_787,N_19312,N_19106);
nor UO_788 (O_788,N_19108,N_19546);
and UO_789 (O_789,N_19134,N_19141);
and UO_790 (O_790,N_19874,N_19362);
or UO_791 (O_791,N_19497,N_19771);
nor UO_792 (O_792,N_19087,N_19016);
and UO_793 (O_793,N_19146,N_19034);
or UO_794 (O_794,N_19254,N_19433);
and UO_795 (O_795,N_19005,N_19106);
nor UO_796 (O_796,N_19515,N_19269);
nor UO_797 (O_797,N_19145,N_19298);
and UO_798 (O_798,N_19290,N_19003);
or UO_799 (O_799,N_19758,N_19610);
nor UO_800 (O_800,N_19947,N_19080);
nand UO_801 (O_801,N_19161,N_19850);
and UO_802 (O_802,N_19365,N_19925);
or UO_803 (O_803,N_19912,N_19161);
nor UO_804 (O_804,N_19512,N_19623);
xor UO_805 (O_805,N_19310,N_19705);
nor UO_806 (O_806,N_19975,N_19096);
nor UO_807 (O_807,N_19010,N_19971);
xnor UO_808 (O_808,N_19777,N_19919);
xnor UO_809 (O_809,N_19070,N_19707);
nor UO_810 (O_810,N_19518,N_19844);
or UO_811 (O_811,N_19351,N_19879);
or UO_812 (O_812,N_19021,N_19160);
nor UO_813 (O_813,N_19006,N_19077);
or UO_814 (O_814,N_19535,N_19439);
and UO_815 (O_815,N_19792,N_19853);
and UO_816 (O_816,N_19046,N_19323);
or UO_817 (O_817,N_19290,N_19684);
and UO_818 (O_818,N_19881,N_19664);
nor UO_819 (O_819,N_19644,N_19928);
or UO_820 (O_820,N_19605,N_19662);
nand UO_821 (O_821,N_19235,N_19559);
and UO_822 (O_822,N_19761,N_19110);
or UO_823 (O_823,N_19030,N_19520);
nand UO_824 (O_824,N_19961,N_19498);
nand UO_825 (O_825,N_19730,N_19109);
nor UO_826 (O_826,N_19733,N_19830);
and UO_827 (O_827,N_19886,N_19582);
and UO_828 (O_828,N_19707,N_19770);
or UO_829 (O_829,N_19767,N_19787);
nor UO_830 (O_830,N_19042,N_19697);
nor UO_831 (O_831,N_19495,N_19284);
xnor UO_832 (O_832,N_19441,N_19945);
nand UO_833 (O_833,N_19040,N_19332);
nand UO_834 (O_834,N_19531,N_19482);
and UO_835 (O_835,N_19993,N_19669);
nand UO_836 (O_836,N_19598,N_19516);
and UO_837 (O_837,N_19320,N_19917);
or UO_838 (O_838,N_19588,N_19547);
or UO_839 (O_839,N_19189,N_19063);
or UO_840 (O_840,N_19195,N_19585);
or UO_841 (O_841,N_19766,N_19239);
and UO_842 (O_842,N_19984,N_19893);
or UO_843 (O_843,N_19987,N_19558);
nand UO_844 (O_844,N_19163,N_19590);
nand UO_845 (O_845,N_19654,N_19012);
or UO_846 (O_846,N_19965,N_19681);
and UO_847 (O_847,N_19730,N_19738);
nand UO_848 (O_848,N_19418,N_19604);
or UO_849 (O_849,N_19566,N_19518);
xor UO_850 (O_850,N_19391,N_19644);
nand UO_851 (O_851,N_19783,N_19126);
nor UO_852 (O_852,N_19401,N_19328);
or UO_853 (O_853,N_19409,N_19517);
or UO_854 (O_854,N_19505,N_19966);
nor UO_855 (O_855,N_19249,N_19867);
nor UO_856 (O_856,N_19374,N_19725);
or UO_857 (O_857,N_19909,N_19740);
or UO_858 (O_858,N_19115,N_19387);
xnor UO_859 (O_859,N_19342,N_19682);
nand UO_860 (O_860,N_19737,N_19657);
xnor UO_861 (O_861,N_19242,N_19673);
xor UO_862 (O_862,N_19430,N_19387);
and UO_863 (O_863,N_19148,N_19143);
and UO_864 (O_864,N_19912,N_19001);
nand UO_865 (O_865,N_19981,N_19482);
nand UO_866 (O_866,N_19555,N_19670);
nand UO_867 (O_867,N_19455,N_19035);
nand UO_868 (O_868,N_19681,N_19324);
or UO_869 (O_869,N_19414,N_19009);
nor UO_870 (O_870,N_19880,N_19910);
nor UO_871 (O_871,N_19653,N_19171);
xnor UO_872 (O_872,N_19986,N_19208);
and UO_873 (O_873,N_19096,N_19604);
nor UO_874 (O_874,N_19774,N_19862);
or UO_875 (O_875,N_19778,N_19497);
and UO_876 (O_876,N_19108,N_19733);
nor UO_877 (O_877,N_19149,N_19980);
and UO_878 (O_878,N_19349,N_19513);
nor UO_879 (O_879,N_19612,N_19710);
nand UO_880 (O_880,N_19929,N_19950);
nor UO_881 (O_881,N_19155,N_19253);
nor UO_882 (O_882,N_19150,N_19642);
or UO_883 (O_883,N_19420,N_19448);
nor UO_884 (O_884,N_19493,N_19134);
and UO_885 (O_885,N_19109,N_19963);
or UO_886 (O_886,N_19942,N_19925);
or UO_887 (O_887,N_19970,N_19910);
or UO_888 (O_888,N_19147,N_19905);
xnor UO_889 (O_889,N_19795,N_19650);
nor UO_890 (O_890,N_19328,N_19666);
nand UO_891 (O_891,N_19945,N_19660);
and UO_892 (O_892,N_19673,N_19288);
nor UO_893 (O_893,N_19666,N_19056);
nor UO_894 (O_894,N_19734,N_19056);
nor UO_895 (O_895,N_19045,N_19255);
xor UO_896 (O_896,N_19230,N_19582);
and UO_897 (O_897,N_19766,N_19980);
or UO_898 (O_898,N_19763,N_19593);
and UO_899 (O_899,N_19278,N_19750);
and UO_900 (O_900,N_19041,N_19176);
nor UO_901 (O_901,N_19702,N_19628);
nand UO_902 (O_902,N_19792,N_19044);
or UO_903 (O_903,N_19768,N_19120);
nand UO_904 (O_904,N_19884,N_19907);
or UO_905 (O_905,N_19080,N_19667);
or UO_906 (O_906,N_19855,N_19328);
and UO_907 (O_907,N_19499,N_19074);
nand UO_908 (O_908,N_19769,N_19639);
or UO_909 (O_909,N_19347,N_19336);
nor UO_910 (O_910,N_19482,N_19694);
nand UO_911 (O_911,N_19208,N_19559);
and UO_912 (O_912,N_19564,N_19459);
nor UO_913 (O_913,N_19927,N_19705);
or UO_914 (O_914,N_19869,N_19495);
xnor UO_915 (O_915,N_19513,N_19224);
xor UO_916 (O_916,N_19936,N_19498);
xor UO_917 (O_917,N_19500,N_19924);
nor UO_918 (O_918,N_19059,N_19017);
and UO_919 (O_919,N_19308,N_19265);
nand UO_920 (O_920,N_19718,N_19641);
or UO_921 (O_921,N_19077,N_19969);
nor UO_922 (O_922,N_19850,N_19596);
or UO_923 (O_923,N_19052,N_19229);
and UO_924 (O_924,N_19996,N_19863);
xor UO_925 (O_925,N_19081,N_19408);
or UO_926 (O_926,N_19303,N_19338);
nor UO_927 (O_927,N_19919,N_19115);
or UO_928 (O_928,N_19399,N_19837);
and UO_929 (O_929,N_19711,N_19565);
xor UO_930 (O_930,N_19171,N_19212);
nor UO_931 (O_931,N_19442,N_19335);
nand UO_932 (O_932,N_19361,N_19907);
nand UO_933 (O_933,N_19296,N_19214);
nand UO_934 (O_934,N_19181,N_19678);
and UO_935 (O_935,N_19417,N_19469);
xor UO_936 (O_936,N_19160,N_19640);
nor UO_937 (O_937,N_19688,N_19900);
or UO_938 (O_938,N_19072,N_19705);
or UO_939 (O_939,N_19578,N_19651);
nand UO_940 (O_940,N_19168,N_19108);
and UO_941 (O_941,N_19982,N_19657);
nand UO_942 (O_942,N_19236,N_19789);
xor UO_943 (O_943,N_19922,N_19565);
nand UO_944 (O_944,N_19872,N_19254);
nand UO_945 (O_945,N_19651,N_19298);
nand UO_946 (O_946,N_19830,N_19497);
xnor UO_947 (O_947,N_19059,N_19864);
or UO_948 (O_948,N_19394,N_19049);
or UO_949 (O_949,N_19485,N_19900);
or UO_950 (O_950,N_19944,N_19872);
and UO_951 (O_951,N_19188,N_19874);
nor UO_952 (O_952,N_19944,N_19330);
or UO_953 (O_953,N_19305,N_19118);
xnor UO_954 (O_954,N_19602,N_19667);
or UO_955 (O_955,N_19269,N_19662);
nor UO_956 (O_956,N_19069,N_19650);
nand UO_957 (O_957,N_19674,N_19665);
or UO_958 (O_958,N_19438,N_19678);
xor UO_959 (O_959,N_19421,N_19462);
nor UO_960 (O_960,N_19263,N_19297);
or UO_961 (O_961,N_19509,N_19190);
and UO_962 (O_962,N_19286,N_19050);
nand UO_963 (O_963,N_19111,N_19685);
nor UO_964 (O_964,N_19062,N_19433);
or UO_965 (O_965,N_19535,N_19291);
nor UO_966 (O_966,N_19312,N_19078);
nor UO_967 (O_967,N_19368,N_19017);
and UO_968 (O_968,N_19963,N_19671);
nand UO_969 (O_969,N_19068,N_19766);
nand UO_970 (O_970,N_19616,N_19902);
nor UO_971 (O_971,N_19895,N_19155);
or UO_972 (O_972,N_19086,N_19118);
nand UO_973 (O_973,N_19279,N_19443);
nor UO_974 (O_974,N_19591,N_19234);
or UO_975 (O_975,N_19482,N_19160);
or UO_976 (O_976,N_19356,N_19849);
or UO_977 (O_977,N_19132,N_19707);
or UO_978 (O_978,N_19877,N_19440);
nor UO_979 (O_979,N_19806,N_19382);
or UO_980 (O_980,N_19109,N_19149);
or UO_981 (O_981,N_19061,N_19692);
nor UO_982 (O_982,N_19489,N_19366);
xnor UO_983 (O_983,N_19092,N_19330);
and UO_984 (O_984,N_19702,N_19886);
nor UO_985 (O_985,N_19834,N_19864);
or UO_986 (O_986,N_19326,N_19886);
nand UO_987 (O_987,N_19298,N_19896);
nand UO_988 (O_988,N_19115,N_19311);
nand UO_989 (O_989,N_19361,N_19424);
or UO_990 (O_990,N_19571,N_19440);
xnor UO_991 (O_991,N_19119,N_19953);
or UO_992 (O_992,N_19624,N_19996);
or UO_993 (O_993,N_19269,N_19285);
nand UO_994 (O_994,N_19991,N_19696);
nand UO_995 (O_995,N_19583,N_19866);
xnor UO_996 (O_996,N_19599,N_19541);
nor UO_997 (O_997,N_19815,N_19153);
xnor UO_998 (O_998,N_19375,N_19498);
nand UO_999 (O_999,N_19428,N_19363);
nand UO_1000 (O_1000,N_19266,N_19988);
nor UO_1001 (O_1001,N_19976,N_19358);
or UO_1002 (O_1002,N_19395,N_19298);
or UO_1003 (O_1003,N_19369,N_19535);
and UO_1004 (O_1004,N_19729,N_19732);
nand UO_1005 (O_1005,N_19069,N_19168);
or UO_1006 (O_1006,N_19002,N_19785);
and UO_1007 (O_1007,N_19111,N_19391);
or UO_1008 (O_1008,N_19349,N_19580);
and UO_1009 (O_1009,N_19539,N_19554);
and UO_1010 (O_1010,N_19994,N_19424);
xor UO_1011 (O_1011,N_19716,N_19107);
or UO_1012 (O_1012,N_19132,N_19269);
nand UO_1013 (O_1013,N_19981,N_19882);
or UO_1014 (O_1014,N_19839,N_19157);
and UO_1015 (O_1015,N_19945,N_19250);
nor UO_1016 (O_1016,N_19575,N_19431);
nor UO_1017 (O_1017,N_19275,N_19464);
and UO_1018 (O_1018,N_19022,N_19453);
nand UO_1019 (O_1019,N_19854,N_19851);
and UO_1020 (O_1020,N_19238,N_19888);
nand UO_1021 (O_1021,N_19172,N_19775);
and UO_1022 (O_1022,N_19070,N_19857);
and UO_1023 (O_1023,N_19693,N_19975);
nand UO_1024 (O_1024,N_19006,N_19518);
and UO_1025 (O_1025,N_19965,N_19266);
or UO_1026 (O_1026,N_19350,N_19488);
or UO_1027 (O_1027,N_19675,N_19029);
nor UO_1028 (O_1028,N_19544,N_19348);
and UO_1029 (O_1029,N_19971,N_19296);
xnor UO_1030 (O_1030,N_19828,N_19496);
xor UO_1031 (O_1031,N_19581,N_19454);
and UO_1032 (O_1032,N_19589,N_19971);
nand UO_1033 (O_1033,N_19363,N_19102);
nand UO_1034 (O_1034,N_19625,N_19263);
nor UO_1035 (O_1035,N_19829,N_19291);
nor UO_1036 (O_1036,N_19230,N_19776);
and UO_1037 (O_1037,N_19402,N_19500);
nand UO_1038 (O_1038,N_19394,N_19582);
and UO_1039 (O_1039,N_19035,N_19517);
nor UO_1040 (O_1040,N_19320,N_19829);
nor UO_1041 (O_1041,N_19355,N_19314);
or UO_1042 (O_1042,N_19386,N_19464);
nand UO_1043 (O_1043,N_19428,N_19725);
xnor UO_1044 (O_1044,N_19993,N_19825);
or UO_1045 (O_1045,N_19119,N_19290);
nand UO_1046 (O_1046,N_19632,N_19857);
or UO_1047 (O_1047,N_19674,N_19198);
nor UO_1048 (O_1048,N_19281,N_19354);
xor UO_1049 (O_1049,N_19726,N_19031);
nor UO_1050 (O_1050,N_19485,N_19646);
nand UO_1051 (O_1051,N_19340,N_19256);
nor UO_1052 (O_1052,N_19274,N_19121);
and UO_1053 (O_1053,N_19186,N_19799);
nor UO_1054 (O_1054,N_19255,N_19966);
xor UO_1055 (O_1055,N_19840,N_19485);
nor UO_1056 (O_1056,N_19337,N_19314);
or UO_1057 (O_1057,N_19507,N_19218);
and UO_1058 (O_1058,N_19301,N_19933);
and UO_1059 (O_1059,N_19329,N_19067);
xor UO_1060 (O_1060,N_19466,N_19415);
nand UO_1061 (O_1061,N_19774,N_19337);
or UO_1062 (O_1062,N_19636,N_19946);
or UO_1063 (O_1063,N_19528,N_19565);
and UO_1064 (O_1064,N_19599,N_19094);
nor UO_1065 (O_1065,N_19343,N_19777);
nor UO_1066 (O_1066,N_19642,N_19215);
and UO_1067 (O_1067,N_19305,N_19619);
and UO_1068 (O_1068,N_19077,N_19071);
and UO_1069 (O_1069,N_19458,N_19625);
or UO_1070 (O_1070,N_19937,N_19182);
nand UO_1071 (O_1071,N_19823,N_19574);
nand UO_1072 (O_1072,N_19036,N_19888);
and UO_1073 (O_1073,N_19857,N_19303);
nor UO_1074 (O_1074,N_19210,N_19736);
nand UO_1075 (O_1075,N_19612,N_19860);
or UO_1076 (O_1076,N_19975,N_19955);
nor UO_1077 (O_1077,N_19064,N_19632);
nor UO_1078 (O_1078,N_19894,N_19311);
nand UO_1079 (O_1079,N_19770,N_19877);
or UO_1080 (O_1080,N_19587,N_19863);
and UO_1081 (O_1081,N_19239,N_19512);
and UO_1082 (O_1082,N_19016,N_19023);
or UO_1083 (O_1083,N_19428,N_19919);
nor UO_1084 (O_1084,N_19441,N_19678);
or UO_1085 (O_1085,N_19773,N_19443);
or UO_1086 (O_1086,N_19006,N_19606);
nor UO_1087 (O_1087,N_19337,N_19666);
nand UO_1088 (O_1088,N_19044,N_19446);
nand UO_1089 (O_1089,N_19385,N_19229);
xnor UO_1090 (O_1090,N_19107,N_19769);
and UO_1091 (O_1091,N_19199,N_19961);
nand UO_1092 (O_1092,N_19637,N_19068);
nand UO_1093 (O_1093,N_19524,N_19788);
or UO_1094 (O_1094,N_19089,N_19684);
xor UO_1095 (O_1095,N_19672,N_19324);
nor UO_1096 (O_1096,N_19049,N_19486);
or UO_1097 (O_1097,N_19614,N_19417);
xnor UO_1098 (O_1098,N_19144,N_19487);
and UO_1099 (O_1099,N_19980,N_19881);
nor UO_1100 (O_1100,N_19197,N_19980);
nor UO_1101 (O_1101,N_19519,N_19798);
xnor UO_1102 (O_1102,N_19684,N_19620);
nand UO_1103 (O_1103,N_19557,N_19324);
or UO_1104 (O_1104,N_19238,N_19329);
and UO_1105 (O_1105,N_19864,N_19338);
nor UO_1106 (O_1106,N_19758,N_19983);
nand UO_1107 (O_1107,N_19858,N_19845);
nand UO_1108 (O_1108,N_19803,N_19675);
nor UO_1109 (O_1109,N_19433,N_19050);
nor UO_1110 (O_1110,N_19206,N_19863);
nor UO_1111 (O_1111,N_19504,N_19848);
and UO_1112 (O_1112,N_19648,N_19552);
or UO_1113 (O_1113,N_19574,N_19585);
or UO_1114 (O_1114,N_19085,N_19527);
or UO_1115 (O_1115,N_19169,N_19525);
nand UO_1116 (O_1116,N_19828,N_19744);
and UO_1117 (O_1117,N_19821,N_19797);
nand UO_1118 (O_1118,N_19911,N_19778);
nor UO_1119 (O_1119,N_19065,N_19386);
and UO_1120 (O_1120,N_19670,N_19931);
nor UO_1121 (O_1121,N_19019,N_19024);
or UO_1122 (O_1122,N_19248,N_19900);
or UO_1123 (O_1123,N_19157,N_19663);
or UO_1124 (O_1124,N_19261,N_19560);
or UO_1125 (O_1125,N_19343,N_19146);
nor UO_1126 (O_1126,N_19775,N_19728);
and UO_1127 (O_1127,N_19418,N_19796);
xor UO_1128 (O_1128,N_19494,N_19802);
and UO_1129 (O_1129,N_19369,N_19101);
nand UO_1130 (O_1130,N_19010,N_19202);
nand UO_1131 (O_1131,N_19989,N_19769);
and UO_1132 (O_1132,N_19453,N_19245);
nor UO_1133 (O_1133,N_19130,N_19618);
nor UO_1134 (O_1134,N_19695,N_19727);
nor UO_1135 (O_1135,N_19923,N_19335);
or UO_1136 (O_1136,N_19991,N_19783);
or UO_1137 (O_1137,N_19398,N_19810);
or UO_1138 (O_1138,N_19696,N_19704);
or UO_1139 (O_1139,N_19293,N_19019);
nor UO_1140 (O_1140,N_19833,N_19618);
nor UO_1141 (O_1141,N_19444,N_19169);
or UO_1142 (O_1142,N_19364,N_19584);
or UO_1143 (O_1143,N_19370,N_19682);
and UO_1144 (O_1144,N_19405,N_19285);
nor UO_1145 (O_1145,N_19433,N_19274);
and UO_1146 (O_1146,N_19659,N_19825);
and UO_1147 (O_1147,N_19104,N_19996);
nand UO_1148 (O_1148,N_19261,N_19677);
and UO_1149 (O_1149,N_19074,N_19876);
nand UO_1150 (O_1150,N_19891,N_19572);
nand UO_1151 (O_1151,N_19439,N_19287);
nor UO_1152 (O_1152,N_19367,N_19298);
or UO_1153 (O_1153,N_19548,N_19580);
or UO_1154 (O_1154,N_19307,N_19704);
nand UO_1155 (O_1155,N_19475,N_19862);
and UO_1156 (O_1156,N_19977,N_19455);
and UO_1157 (O_1157,N_19878,N_19684);
or UO_1158 (O_1158,N_19503,N_19112);
and UO_1159 (O_1159,N_19874,N_19761);
nand UO_1160 (O_1160,N_19379,N_19877);
xor UO_1161 (O_1161,N_19451,N_19336);
xnor UO_1162 (O_1162,N_19585,N_19919);
nand UO_1163 (O_1163,N_19475,N_19591);
or UO_1164 (O_1164,N_19061,N_19564);
xnor UO_1165 (O_1165,N_19047,N_19913);
xor UO_1166 (O_1166,N_19320,N_19792);
nand UO_1167 (O_1167,N_19810,N_19955);
and UO_1168 (O_1168,N_19508,N_19792);
nand UO_1169 (O_1169,N_19157,N_19253);
and UO_1170 (O_1170,N_19450,N_19239);
or UO_1171 (O_1171,N_19213,N_19946);
xnor UO_1172 (O_1172,N_19423,N_19707);
xor UO_1173 (O_1173,N_19829,N_19300);
or UO_1174 (O_1174,N_19993,N_19448);
and UO_1175 (O_1175,N_19710,N_19908);
and UO_1176 (O_1176,N_19898,N_19782);
nor UO_1177 (O_1177,N_19455,N_19362);
or UO_1178 (O_1178,N_19133,N_19539);
nand UO_1179 (O_1179,N_19892,N_19789);
or UO_1180 (O_1180,N_19109,N_19082);
nand UO_1181 (O_1181,N_19197,N_19852);
nand UO_1182 (O_1182,N_19350,N_19576);
and UO_1183 (O_1183,N_19377,N_19663);
and UO_1184 (O_1184,N_19304,N_19571);
nor UO_1185 (O_1185,N_19880,N_19289);
nand UO_1186 (O_1186,N_19850,N_19702);
nor UO_1187 (O_1187,N_19437,N_19676);
and UO_1188 (O_1188,N_19805,N_19202);
nor UO_1189 (O_1189,N_19285,N_19346);
and UO_1190 (O_1190,N_19748,N_19478);
nor UO_1191 (O_1191,N_19441,N_19634);
nor UO_1192 (O_1192,N_19707,N_19639);
nand UO_1193 (O_1193,N_19810,N_19489);
or UO_1194 (O_1194,N_19505,N_19056);
or UO_1195 (O_1195,N_19915,N_19784);
xnor UO_1196 (O_1196,N_19260,N_19573);
or UO_1197 (O_1197,N_19795,N_19750);
nand UO_1198 (O_1198,N_19967,N_19893);
or UO_1199 (O_1199,N_19508,N_19560);
or UO_1200 (O_1200,N_19458,N_19313);
nand UO_1201 (O_1201,N_19797,N_19049);
or UO_1202 (O_1202,N_19096,N_19673);
and UO_1203 (O_1203,N_19665,N_19606);
or UO_1204 (O_1204,N_19784,N_19198);
nand UO_1205 (O_1205,N_19526,N_19674);
and UO_1206 (O_1206,N_19302,N_19002);
nand UO_1207 (O_1207,N_19086,N_19496);
nand UO_1208 (O_1208,N_19018,N_19081);
nand UO_1209 (O_1209,N_19544,N_19210);
nor UO_1210 (O_1210,N_19212,N_19240);
nor UO_1211 (O_1211,N_19070,N_19527);
and UO_1212 (O_1212,N_19869,N_19138);
and UO_1213 (O_1213,N_19468,N_19181);
nand UO_1214 (O_1214,N_19711,N_19227);
nand UO_1215 (O_1215,N_19496,N_19975);
nor UO_1216 (O_1216,N_19114,N_19847);
nand UO_1217 (O_1217,N_19958,N_19535);
nand UO_1218 (O_1218,N_19758,N_19626);
nand UO_1219 (O_1219,N_19191,N_19491);
and UO_1220 (O_1220,N_19325,N_19578);
nand UO_1221 (O_1221,N_19092,N_19497);
nand UO_1222 (O_1222,N_19639,N_19371);
or UO_1223 (O_1223,N_19231,N_19852);
or UO_1224 (O_1224,N_19272,N_19972);
or UO_1225 (O_1225,N_19241,N_19782);
and UO_1226 (O_1226,N_19681,N_19034);
or UO_1227 (O_1227,N_19435,N_19519);
nand UO_1228 (O_1228,N_19417,N_19142);
nand UO_1229 (O_1229,N_19527,N_19235);
or UO_1230 (O_1230,N_19143,N_19761);
or UO_1231 (O_1231,N_19683,N_19283);
and UO_1232 (O_1232,N_19732,N_19161);
xor UO_1233 (O_1233,N_19182,N_19391);
and UO_1234 (O_1234,N_19905,N_19314);
or UO_1235 (O_1235,N_19491,N_19413);
nor UO_1236 (O_1236,N_19185,N_19341);
nor UO_1237 (O_1237,N_19525,N_19113);
or UO_1238 (O_1238,N_19428,N_19272);
nand UO_1239 (O_1239,N_19853,N_19885);
nand UO_1240 (O_1240,N_19889,N_19683);
nand UO_1241 (O_1241,N_19818,N_19562);
nor UO_1242 (O_1242,N_19689,N_19263);
xor UO_1243 (O_1243,N_19509,N_19932);
or UO_1244 (O_1244,N_19462,N_19790);
nand UO_1245 (O_1245,N_19032,N_19338);
and UO_1246 (O_1246,N_19909,N_19920);
and UO_1247 (O_1247,N_19292,N_19291);
and UO_1248 (O_1248,N_19036,N_19544);
and UO_1249 (O_1249,N_19049,N_19582);
nor UO_1250 (O_1250,N_19297,N_19492);
nor UO_1251 (O_1251,N_19604,N_19618);
nor UO_1252 (O_1252,N_19599,N_19102);
and UO_1253 (O_1253,N_19501,N_19254);
nand UO_1254 (O_1254,N_19381,N_19193);
or UO_1255 (O_1255,N_19430,N_19617);
nand UO_1256 (O_1256,N_19311,N_19477);
nor UO_1257 (O_1257,N_19985,N_19510);
nor UO_1258 (O_1258,N_19865,N_19788);
nand UO_1259 (O_1259,N_19192,N_19217);
and UO_1260 (O_1260,N_19270,N_19471);
nand UO_1261 (O_1261,N_19461,N_19911);
nor UO_1262 (O_1262,N_19780,N_19145);
and UO_1263 (O_1263,N_19797,N_19699);
nor UO_1264 (O_1264,N_19674,N_19143);
and UO_1265 (O_1265,N_19232,N_19480);
or UO_1266 (O_1266,N_19840,N_19076);
and UO_1267 (O_1267,N_19898,N_19592);
nand UO_1268 (O_1268,N_19703,N_19149);
or UO_1269 (O_1269,N_19655,N_19683);
nor UO_1270 (O_1270,N_19945,N_19161);
nor UO_1271 (O_1271,N_19946,N_19541);
nand UO_1272 (O_1272,N_19243,N_19769);
and UO_1273 (O_1273,N_19330,N_19953);
and UO_1274 (O_1274,N_19875,N_19716);
and UO_1275 (O_1275,N_19340,N_19723);
nor UO_1276 (O_1276,N_19601,N_19784);
nand UO_1277 (O_1277,N_19356,N_19083);
or UO_1278 (O_1278,N_19459,N_19763);
or UO_1279 (O_1279,N_19855,N_19083);
or UO_1280 (O_1280,N_19820,N_19826);
nand UO_1281 (O_1281,N_19762,N_19547);
nor UO_1282 (O_1282,N_19467,N_19329);
nor UO_1283 (O_1283,N_19827,N_19199);
or UO_1284 (O_1284,N_19952,N_19642);
and UO_1285 (O_1285,N_19832,N_19184);
or UO_1286 (O_1286,N_19277,N_19319);
nor UO_1287 (O_1287,N_19314,N_19739);
or UO_1288 (O_1288,N_19457,N_19934);
nor UO_1289 (O_1289,N_19721,N_19387);
or UO_1290 (O_1290,N_19730,N_19983);
and UO_1291 (O_1291,N_19962,N_19297);
and UO_1292 (O_1292,N_19035,N_19110);
and UO_1293 (O_1293,N_19049,N_19652);
and UO_1294 (O_1294,N_19506,N_19586);
and UO_1295 (O_1295,N_19593,N_19394);
or UO_1296 (O_1296,N_19880,N_19834);
nand UO_1297 (O_1297,N_19885,N_19520);
nand UO_1298 (O_1298,N_19643,N_19322);
or UO_1299 (O_1299,N_19034,N_19134);
nor UO_1300 (O_1300,N_19211,N_19839);
nor UO_1301 (O_1301,N_19569,N_19677);
nor UO_1302 (O_1302,N_19920,N_19882);
and UO_1303 (O_1303,N_19829,N_19296);
and UO_1304 (O_1304,N_19787,N_19331);
and UO_1305 (O_1305,N_19539,N_19640);
nand UO_1306 (O_1306,N_19949,N_19103);
nor UO_1307 (O_1307,N_19333,N_19562);
nand UO_1308 (O_1308,N_19858,N_19174);
or UO_1309 (O_1309,N_19560,N_19316);
and UO_1310 (O_1310,N_19146,N_19471);
or UO_1311 (O_1311,N_19018,N_19870);
nand UO_1312 (O_1312,N_19764,N_19951);
nor UO_1313 (O_1313,N_19539,N_19954);
nor UO_1314 (O_1314,N_19643,N_19187);
nor UO_1315 (O_1315,N_19290,N_19746);
or UO_1316 (O_1316,N_19210,N_19901);
or UO_1317 (O_1317,N_19147,N_19045);
nand UO_1318 (O_1318,N_19685,N_19574);
nor UO_1319 (O_1319,N_19294,N_19769);
nand UO_1320 (O_1320,N_19585,N_19140);
nand UO_1321 (O_1321,N_19321,N_19358);
xnor UO_1322 (O_1322,N_19887,N_19315);
xnor UO_1323 (O_1323,N_19282,N_19200);
xnor UO_1324 (O_1324,N_19169,N_19264);
and UO_1325 (O_1325,N_19354,N_19869);
or UO_1326 (O_1326,N_19321,N_19426);
or UO_1327 (O_1327,N_19580,N_19967);
or UO_1328 (O_1328,N_19522,N_19592);
nand UO_1329 (O_1329,N_19419,N_19107);
and UO_1330 (O_1330,N_19352,N_19115);
nor UO_1331 (O_1331,N_19644,N_19397);
or UO_1332 (O_1332,N_19480,N_19660);
or UO_1333 (O_1333,N_19894,N_19380);
or UO_1334 (O_1334,N_19598,N_19912);
or UO_1335 (O_1335,N_19384,N_19367);
xor UO_1336 (O_1336,N_19774,N_19974);
and UO_1337 (O_1337,N_19885,N_19980);
or UO_1338 (O_1338,N_19123,N_19061);
and UO_1339 (O_1339,N_19631,N_19801);
or UO_1340 (O_1340,N_19708,N_19950);
nand UO_1341 (O_1341,N_19233,N_19061);
nand UO_1342 (O_1342,N_19845,N_19133);
and UO_1343 (O_1343,N_19868,N_19649);
and UO_1344 (O_1344,N_19397,N_19857);
or UO_1345 (O_1345,N_19481,N_19421);
and UO_1346 (O_1346,N_19118,N_19882);
nor UO_1347 (O_1347,N_19490,N_19040);
nor UO_1348 (O_1348,N_19206,N_19739);
nand UO_1349 (O_1349,N_19707,N_19051);
nand UO_1350 (O_1350,N_19641,N_19179);
nand UO_1351 (O_1351,N_19502,N_19236);
nor UO_1352 (O_1352,N_19977,N_19511);
and UO_1353 (O_1353,N_19959,N_19582);
nor UO_1354 (O_1354,N_19009,N_19269);
nand UO_1355 (O_1355,N_19841,N_19111);
nand UO_1356 (O_1356,N_19862,N_19815);
nor UO_1357 (O_1357,N_19007,N_19322);
xnor UO_1358 (O_1358,N_19302,N_19809);
nand UO_1359 (O_1359,N_19722,N_19614);
or UO_1360 (O_1360,N_19035,N_19037);
nand UO_1361 (O_1361,N_19406,N_19830);
and UO_1362 (O_1362,N_19986,N_19673);
nor UO_1363 (O_1363,N_19053,N_19016);
and UO_1364 (O_1364,N_19431,N_19462);
nor UO_1365 (O_1365,N_19639,N_19882);
xor UO_1366 (O_1366,N_19828,N_19938);
and UO_1367 (O_1367,N_19074,N_19163);
nor UO_1368 (O_1368,N_19618,N_19351);
nand UO_1369 (O_1369,N_19608,N_19813);
nor UO_1370 (O_1370,N_19921,N_19736);
and UO_1371 (O_1371,N_19659,N_19265);
or UO_1372 (O_1372,N_19735,N_19158);
and UO_1373 (O_1373,N_19132,N_19006);
and UO_1374 (O_1374,N_19362,N_19968);
nor UO_1375 (O_1375,N_19809,N_19133);
nor UO_1376 (O_1376,N_19653,N_19656);
and UO_1377 (O_1377,N_19786,N_19682);
or UO_1378 (O_1378,N_19093,N_19317);
nand UO_1379 (O_1379,N_19246,N_19830);
and UO_1380 (O_1380,N_19318,N_19103);
and UO_1381 (O_1381,N_19217,N_19674);
and UO_1382 (O_1382,N_19742,N_19999);
and UO_1383 (O_1383,N_19121,N_19498);
or UO_1384 (O_1384,N_19445,N_19394);
and UO_1385 (O_1385,N_19826,N_19342);
xnor UO_1386 (O_1386,N_19606,N_19794);
nor UO_1387 (O_1387,N_19645,N_19876);
nor UO_1388 (O_1388,N_19146,N_19184);
and UO_1389 (O_1389,N_19408,N_19650);
xnor UO_1390 (O_1390,N_19333,N_19680);
or UO_1391 (O_1391,N_19153,N_19649);
nand UO_1392 (O_1392,N_19354,N_19123);
and UO_1393 (O_1393,N_19410,N_19639);
or UO_1394 (O_1394,N_19249,N_19260);
or UO_1395 (O_1395,N_19197,N_19914);
nand UO_1396 (O_1396,N_19035,N_19675);
nor UO_1397 (O_1397,N_19399,N_19141);
nor UO_1398 (O_1398,N_19831,N_19682);
and UO_1399 (O_1399,N_19735,N_19473);
nor UO_1400 (O_1400,N_19127,N_19881);
nor UO_1401 (O_1401,N_19582,N_19955);
or UO_1402 (O_1402,N_19160,N_19848);
nand UO_1403 (O_1403,N_19589,N_19949);
and UO_1404 (O_1404,N_19937,N_19480);
or UO_1405 (O_1405,N_19341,N_19115);
nor UO_1406 (O_1406,N_19288,N_19498);
and UO_1407 (O_1407,N_19747,N_19874);
nor UO_1408 (O_1408,N_19318,N_19899);
and UO_1409 (O_1409,N_19549,N_19828);
or UO_1410 (O_1410,N_19257,N_19823);
nand UO_1411 (O_1411,N_19243,N_19481);
and UO_1412 (O_1412,N_19250,N_19855);
nand UO_1413 (O_1413,N_19496,N_19246);
or UO_1414 (O_1414,N_19784,N_19785);
or UO_1415 (O_1415,N_19510,N_19806);
and UO_1416 (O_1416,N_19495,N_19442);
or UO_1417 (O_1417,N_19315,N_19081);
or UO_1418 (O_1418,N_19743,N_19095);
or UO_1419 (O_1419,N_19442,N_19959);
and UO_1420 (O_1420,N_19033,N_19190);
nor UO_1421 (O_1421,N_19809,N_19544);
nor UO_1422 (O_1422,N_19113,N_19896);
nand UO_1423 (O_1423,N_19336,N_19127);
and UO_1424 (O_1424,N_19898,N_19748);
or UO_1425 (O_1425,N_19494,N_19342);
and UO_1426 (O_1426,N_19278,N_19699);
nor UO_1427 (O_1427,N_19288,N_19437);
or UO_1428 (O_1428,N_19873,N_19543);
nand UO_1429 (O_1429,N_19048,N_19685);
or UO_1430 (O_1430,N_19965,N_19518);
nor UO_1431 (O_1431,N_19984,N_19963);
and UO_1432 (O_1432,N_19372,N_19536);
xor UO_1433 (O_1433,N_19251,N_19237);
xnor UO_1434 (O_1434,N_19276,N_19345);
nor UO_1435 (O_1435,N_19682,N_19426);
and UO_1436 (O_1436,N_19899,N_19912);
nand UO_1437 (O_1437,N_19680,N_19516);
nor UO_1438 (O_1438,N_19453,N_19064);
and UO_1439 (O_1439,N_19032,N_19826);
nand UO_1440 (O_1440,N_19463,N_19705);
and UO_1441 (O_1441,N_19557,N_19939);
or UO_1442 (O_1442,N_19524,N_19299);
nand UO_1443 (O_1443,N_19770,N_19303);
and UO_1444 (O_1444,N_19074,N_19410);
or UO_1445 (O_1445,N_19471,N_19181);
nand UO_1446 (O_1446,N_19932,N_19708);
nor UO_1447 (O_1447,N_19992,N_19399);
and UO_1448 (O_1448,N_19730,N_19243);
xnor UO_1449 (O_1449,N_19800,N_19990);
nand UO_1450 (O_1450,N_19145,N_19806);
nand UO_1451 (O_1451,N_19868,N_19755);
or UO_1452 (O_1452,N_19743,N_19187);
nand UO_1453 (O_1453,N_19171,N_19311);
and UO_1454 (O_1454,N_19411,N_19044);
and UO_1455 (O_1455,N_19495,N_19155);
nor UO_1456 (O_1456,N_19173,N_19814);
or UO_1457 (O_1457,N_19109,N_19589);
nor UO_1458 (O_1458,N_19728,N_19421);
nand UO_1459 (O_1459,N_19144,N_19986);
or UO_1460 (O_1460,N_19146,N_19783);
nand UO_1461 (O_1461,N_19485,N_19553);
nor UO_1462 (O_1462,N_19296,N_19819);
nor UO_1463 (O_1463,N_19649,N_19595);
nor UO_1464 (O_1464,N_19849,N_19352);
and UO_1465 (O_1465,N_19859,N_19488);
nand UO_1466 (O_1466,N_19845,N_19953);
or UO_1467 (O_1467,N_19340,N_19400);
or UO_1468 (O_1468,N_19498,N_19863);
and UO_1469 (O_1469,N_19470,N_19031);
or UO_1470 (O_1470,N_19701,N_19285);
nand UO_1471 (O_1471,N_19926,N_19903);
and UO_1472 (O_1472,N_19606,N_19924);
xor UO_1473 (O_1473,N_19935,N_19630);
nor UO_1474 (O_1474,N_19429,N_19292);
and UO_1475 (O_1475,N_19468,N_19325);
or UO_1476 (O_1476,N_19197,N_19645);
xnor UO_1477 (O_1477,N_19396,N_19840);
and UO_1478 (O_1478,N_19014,N_19191);
or UO_1479 (O_1479,N_19855,N_19260);
xnor UO_1480 (O_1480,N_19049,N_19297);
nor UO_1481 (O_1481,N_19821,N_19432);
xnor UO_1482 (O_1482,N_19647,N_19987);
or UO_1483 (O_1483,N_19509,N_19357);
or UO_1484 (O_1484,N_19940,N_19463);
or UO_1485 (O_1485,N_19013,N_19726);
nand UO_1486 (O_1486,N_19053,N_19726);
nand UO_1487 (O_1487,N_19220,N_19612);
nand UO_1488 (O_1488,N_19948,N_19511);
nor UO_1489 (O_1489,N_19859,N_19419);
nor UO_1490 (O_1490,N_19611,N_19124);
nand UO_1491 (O_1491,N_19365,N_19954);
and UO_1492 (O_1492,N_19478,N_19287);
nor UO_1493 (O_1493,N_19618,N_19206);
or UO_1494 (O_1494,N_19083,N_19748);
or UO_1495 (O_1495,N_19937,N_19277);
and UO_1496 (O_1496,N_19525,N_19185);
or UO_1497 (O_1497,N_19413,N_19036);
and UO_1498 (O_1498,N_19733,N_19265);
nand UO_1499 (O_1499,N_19358,N_19804);
and UO_1500 (O_1500,N_19881,N_19459);
xnor UO_1501 (O_1501,N_19518,N_19912);
nor UO_1502 (O_1502,N_19548,N_19001);
nand UO_1503 (O_1503,N_19978,N_19030);
nor UO_1504 (O_1504,N_19473,N_19114);
nand UO_1505 (O_1505,N_19027,N_19911);
nand UO_1506 (O_1506,N_19940,N_19058);
and UO_1507 (O_1507,N_19641,N_19058);
or UO_1508 (O_1508,N_19170,N_19014);
nor UO_1509 (O_1509,N_19539,N_19275);
xnor UO_1510 (O_1510,N_19715,N_19876);
nand UO_1511 (O_1511,N_19739,N_19911);
nor UO_1512 (O_1512,N_19497,N_19699);
xor UO_1513 (O_1513,N_19237,N_19460);
and UO_1514 (O_1514,N_19006,N_19971);
and UO_1515 (O_1515,N_19730,N_19687);
or UO_1516 (O_1516,N_19921,N_19871);
or UO_1517 (O_1517,N_19543,N_19173);
nor UO_1518 (O_1518,N_19180,N_19876);
or UO_1519 (O_1519,N_19780,N_19373);
nand UO_1520 (O_1520,N_19632,N_19746);
and UO_1521 (O_1521,N_19700,N_19402);
or UO_1522 (O_1522,N_19659,N_19215);
and UO_1523 (O_1523,N_19931,N_19714);
and UO_1524 (O_1524,N_19384,N_19884);
xnor UO_1525 (O_1525,N_19351,N_19184);
nand UO_1526 (O_1526,N_19265,N_19972);
and UO_1527 (O_1527,N_19742,N_19840);
nand UO_1528 (O_1528,N_19090,N_19988);
and UO_1529 (O_1529,N_19768,N_19688);
nor UO_1530 (O_1530,N_19468,N_19611);
nand UO_1531 (O_1531,N_19026,N_19163);
nand UO_1532 (O_1532,N_19921,N_19052);
nand UO_1533 (O_1533,N_19652,N_19020);
nor UO_1534 (O_1534,N_19802,N_19487);
xnor UO_1535 (O_1535,N_19193,N_19345);
nor UO_1536 (O_1536,N_19691,N_19093);
or UO_1537 (O_1537,N_19537,N_19451);
and UO_1538 (O_1538,N_19562,N_19695);
nor UO_1539 (O_1539,N_19209,N_19325);
nand UO_1540 (O_1540,N_19665,N_19150);
xnor UO_1541 (O_1541,N_19369,N_19853);
xor UO_1542 (O_1542,N_19018,N_19910);
nand UO_1543 (O_1543,N_19858,N_19457);
nor UO_1544 (O_1544,N_19721,N_19166);
or UO_1545 (O_1545,N_19848,N_19413);
xnor UO_1546 (O_1546,N_19043,N_19120);
and UO_1547 (O_1547,N_19300,N_19714);
or UO_1548 (O_1548,N_19084,N_19399);
or UO_1549 (O_1549,N_19722,N_19782);
and UO_1550 (O_1550,N_19666,N_19942);
nand UO_1551 (O_1551,N_19304,N_19352);
or UO_1552 (O_1552,N_19165,N_19632);
nor UO_1553 (O_1553,N_19130,N_19607);
xor UO_1554 (O_1554,N_19024,N_19791);
and UO_1555 (O_1555,N_19045,N_19962);
or UO_1556 (O_1556,N_19077,N_19706);
nand UO_1557 (O_1557,N_19622,N_19488);
or UO_1558 (O_1558,N_19962,N_19480);
nand UO_1559 (O_1559,N_19375,N_19694);
or UO_1560 (O_1560,N_19264,N_19496);
and UO_1561 (O_1561,N_19321,N_19949);
nor UO_1562 (O_1562,N_19718,N_19061);
nand UO_1563 (O_1563,N_19423,N_19700);
nand UO_1564 (O_1564,N_19358,N_19728);
nor UO_1565 (O_1565,N_19799,N_19703);
nand UO_1566 (O_1566,N_19016,N_19918);
nor UO_1567 (O_1567,N_19616,N_19758);
nor UO_1568 (O_1568,N_19047,N_19336);
nand UO_1569 (O_1569,N_19956,N_19218);
xor UO_1570 (O_1570,N_19100,N_19748);
and UO_1571 (O_1571,N_19324,N_19104);
xnor UO_1572 (O_1572,N_19662,N_19172);
nand UO_1573 (O_1573,N_19521,N_19085);
nand UO_1574 (O_1574,N_19318,N_19371);
nand UO_1575 (O_1575,N_19598,N_19193);
and UO_1576 (O_1576,N_19976,N_19549);
nand UO_1577 (O_1577,N_19313,N_19608);
nor UO_1578 (O_1578,N_19337,N_19051);
and UO_1579 (O_1579,N_19886,N_19150);
and UO_1580 (O_1580,N_19949,N_19486);
nand UO_1581 (O_1581,N_19811,N_19846);
and UO_1582 (O_1582,N_19361,N_19463);
and UO_1583 (O_1583,N_19958,N_19776);
nand UO_1584 (O_1584,N_19285,N_19289);
or UO_1585 (O_1585,N_19722,N_19432);
and UO_1586 (O_1586,N_19822,N_19588);
or UO_1587 (O_1587,N_19301,N_19258);
and UO_1588 (O_1588,N_19177,N_19399);
nor UO_1589 (O_1589,N_19682,N_19317);
and UO_1590 (O_1590,N_19299,N_19867);
nand UO_1591 (O_1591,N_19863,N_19266);
nand UO_1592 (O_1592,N_19948,N_19154);
nor UO_1593 (O_1593,N_19466,N_19237);
and UO_1594 (O_1594,N_19323,N_19088);
or UO_1595 (O_1595,N_19348,N_19270);
xor UO_1596 (O_1596,N_19089,N_19012);
nor UO_1597 (O_1597,N_19123,N_19008);
or UO_1598 (O_1598,N_19846,N_19572);
and UO_1599 (O_1599,N_19005,N_19583);
nor UO_1600 (O_1600,N_19731,N_19189);
nor UO_1601 (O_1601,N_19734,N_19820);
and UO_1602 (O_1602,N_19153,N_19111);
xor UO_1603 (O_1603,N_19286,N_19372);
nor UO_1604 (O_1604,N_19444,N_19837);
and UO_1605 (O_1605,N_19919,N_19145);
nand UO_1606 (O_1606,N_19103,N_19809);
or UO_1607 (O_1607,N_19482,N_19957);
nand UO_1608 (O_1608,N_19469,N_19114);
and UO_1609 (O_1609,N_19163,N_19004);
nand UO_1610 (O_1610,N_19497,N_19269);
nor UO_1611 (O_1611,N_19993,N_19404);
and UO_1612 (O_1612,N_19891,N_19723);
nand UO_1613 (O_1613,N_19860,N_19185);
nor UO_1614 (O_1614,N_19350,N_19423);
nand UO_1615 (O_1615,N_19930,N_19956);
nor UO_1616 (O_1616,N_19969,N_19096);
nor UO_1617 (O_1617,N_19635,N_19567);
nand UO_1618 (O_1618,N_19112,N_19293);
or UO_1619 (O_1619,N_19518,N_19888);
nor UO_1620 (O_1620,N_19272,N_19933);
nand UO_1621 (O_1621,N_19593,N_19148);
nand UO_1622 (O_1622,N_19379,N_19158);
xor UO_1623 (O_1623,N_19766,N_19770);
and UO_1624 (O_1624,N_19195,N_19722);
and UO_1625 (O_1625,N_19575,N_19007);
and UO_1626 (O_1626,N_19173,N_19608);
and UO_1627 (O_1627,N_19913,N_19725);
and UO_1628 (O_1628,N_19534,N_19118);
nand UO_1629 (O_1629,N_19497,N_19108);
nand UO_1630 (O_1630,N_19559,N_19856);
and UO_1631 (O_1631,N_19486,N_19796);
or UO_1632 (O_1632,N_19452,N_19921);
nor UO_1633 (O_1633,N_19816,N_19798);
nor UO_1634 (O_1634,N_19883,N_19276);
and UO_1635 (O_1635,N_19391,N_19239);
nor UO_1636 (O_1636,N_19607,N_19455);
nand UO_1637 (O_1637,N_19603,N_19728);
nor UO_1638 (O_1638,N_19278,N_19065);
nor UO_1639 (O_1639,N_19464,N_19452);
nand UO_1640 (O_1640,N_19816,N_19984);
or UO_1641 (O_1641,N_19135,N_19820);
nor UO_1642 (O_1642,N_19838,N_19341);
or UO_1643 (O_1643,N_19588,N_19615);
or UO_1644 (O_1644,N_19939,N_19833);
xor UO_1645 (O_1645,N_19362,N_19700);
nand UO_1646 (O_1646,N_19002,N_19257);
nand UO_1647 (O_1647,N_19763,N_19498);
and UO_1648 (O_1648,N_19220,N_19209);
or UO_1649 (O_1649,N_19547,N_19021);
nor UO_1650 (O_1650,N_19232,N_19118);
xnor UO_1651 (O_1651,N_19639,N_19458);
nor UO_1652 (O_1652,N_19791,N_19649);
and UO_1653 (O_1653,N_19588,N_19382);
xor UO_1654 (O_1654,N_19164,N_19250);
nor UO_1655 (O_1655,N_19409,N_19312);
nand UO_1656 (O_1656,N_19504,N_19941);
xnor UO_1657 (O_1657,N_19770,N_19254);
nand UO_1658 (O_1658,N_19728,N_19023);
nand UO_1659 (O_1659,N_19022,N_19345);
and UO_1660 (O_1660,N_19172,N_19311);
or UO_1661 (O_1661,N_19865,N_19894);
nor UO_1662 (O_1662,N_19449,N_19552);
nor UO_1663 (O_1663,N_19246,N_19862);
nor UO_1664 (O_1664,N_19251,N_19676);
nor UO_1665 (O_1665,N_19185,N_19761);
and UO_1666 (O_1666,N_19903,N_19148);
or UO_1667 (O_1667,N_19842,N_19178);
or UO_1668 (O_1668,N_19313,N_19353);
or UO_1669 (O_1669,N_19554,N_19102);
and UO_1670 (O_1670,N_19016,N_19624);
or UO_1671 (O_1671,N_19699,N_19055);
nand UO_1672 (O_1672,N_19109,N_19607);
and UO_1673 (O_1673,N_19624,N_19240);
or UO_1674 (O_1674,N_19442,N_19354);
nand UO_1675 (O_1675,N_19253,N_19630);
or UO_1676 (O_1676,N_19104,N_19778);
or UO_1677 (O_1677,N_19422,N_19304);
xor UO_1678 (O_1678,N_19934,N_19161);
or UO_1679 (O_1679,N_19863,N_19750);
nand UO_1680 (O_1680,N_19863,N_19673);
and UO_1681 (O_1681,N_19335,N_19053);
xor UO_1682 (O_1682,N_19211,N_19413);
and UO_1683 (O_1683,N_19238,N_19724);
or UO_1684 (O_1684,N_19819,N_19204);
or UO_1685 (O_1685,N_19039,N_19844);
nand UO_1686 (O_1686,N_19987,N_19549);
nor UO_1687 (O_1687,N_19645,N_19621);
nand UO_1688 (O_1688,N_19649,N_19194);
xor UO_1689 (O_1689,N_19971,N_19320);
xor UO_1690 (O_1690,N_19646,N_19623);
or UO_1691 (O_1691,N_19571,N_19132);
or UO_1692 (O_1692,N_19588,N_19869);
nand UO_1693 (O_1693,N_19790,N_19324);
or UO_1694 (O_1694,N_19175,N_19882);
nor UO_1695 (O_1695,N_19713,N_19536);
and UO_1696 (O_1696,N_19694,N_19175);
or UO_1697 (O_1697,N_19049,N_19023);
xnor UO_1698 (O_1698,N_19345,N_19393);
or UO_1699 (O_1699,N_19257,N_19248);
or UO_1700 (O_1700,N_19759,N_19656);
nor UO_1701 (O_1701,N_19565,N_19994);
or UO_1702 (O_1702,N_19798,N_19779);
nand UO_1703 (O_1703,N_19015,N_19446);
and UO_1704 (O_1704,N_19969,N_19828);
nand UO_1705 (O_1705,N_19182,N_19536);
or UO_1706 (O_1706,N_19320,N_19548);
nand UO_1707 (O_1707,N_19428,N_19285);
nor UO_1708 (O_1708,N_19825,N_19978);
or UO_1709 (O_1709,N_19087,N_19698);
or UO_1710 (O_1710,N_19198,N_19158);
and UO_1711 (O_1711,N_19232,N_19742);
nand UO_1712 (O_1712,N_19904,N_19483);
nor UO_1713 (O_1713,N_19472,N_19488);
and UO_1714 (O_1714,N_19418,N_19545);
nor UO_1715 (O_1715,N_19420,N_19772);
and UO_1716 (O_1716,N_19832,N_19885);
xor UO_1717 (O_1717,N_19295,N_19674);
or UO_1718 (O_1718,N_19452,N_19200);
nor UO_1719 (O_1719,N_19232,N_19919);
and UO_1720 (O_1720,N_19326,N_19979);
or UO_1721 (O_1721,N_19321,N_19985);
nand UO_1722 (O_1722,N_19947,N_19484);
nor UO_1723 (O_1723,N_19035,N_19983);
or UO_1724 (O_1724,N_19291,N_19273);
and UO_1725 (O_1725,N_19851,N_19039);
nor UO_1726 (O_1726,N_19745,N_19610);
xnor UO_1727 (O_1727,N_19049,N_19416);
nor UO_1728 (O_1728,N_19183,N_19359);
or UO_1729 (O_1729,N_19341,N_19736);
and UO_1730 (O_1730,N_19764,N_19715);
or UO_1731 (O_1731,N_19605,N_19871);
xnor UO_1732 (O_1732,N_19288,N_19264);
or UO_1733 (O_1733,N_19569,N_19988);
and UO_1734 (O_1734,N_19467,N_19856);
xnor UO_1735 (O_1735,N_19925,N_19994);
nand UO_1736 (O_1736,N_19015,N_19702);
or UO_1737 (O_1737,N_19530,N_19764);
nand UO_1738 (O_1738,N_19770,N_19833);
and UO_1739 (O_1739,N_19685,N_19722);
xnor UO_1740 (O_1740,N_19134,N_19848);
or UO_1741 (O_1741,N_19453,N_19906);
nor UO_1742 (O_1742,N_19213,N_19752);
and UO_1743 (O_1743,N_19840,N_19711);
and UO_1744 (O_1744,N_19338,N_19948);
and UO_1745 (O_1745,N_19144,N_19170);
nor UO_1746 (O_1746,N_19499,N_19035);
or UO_1747 (O_1747,N_19550,N_19409);
and UO_1748 (O_1748,N_19618,N_19898);
and UO_1749 (O_1749,N_19343,N_19864);
and UO_1750 (O_1750,N_19022,N_19033);
or UO_1751 (O_1751,N_19904,N_19012);
and UO_1752 (O_1752,N_19675,N_19722);
and UO_1753 (O_1753,N_19284,N_19248);
and UO_1754 (O_1754,N_19353,N_19635);
nand UO_1755 (O_1755,N_19729,N_19909);
or UO_1756 (O_1756,N_19111,N_19105);
and UO_1757 (O_1757,N_19105,N_19503);
or UO_1758 (O_1758,N_19998,N_19527);
nand UO_1759 (O_1759,N_19743,N_19670);
nand UO_1760 (O_1760,N_19146,N_19145);
xnor UO_1761 (O_1761,N_19712,N_19492);
nor UO_1762 (O_1762,N_19865,N_19166);
nand UO_1763 (O_1763,N_19687,N_19844);
and UO_1764 (O_1764,N_19649,N_19526);
xor UO_1765 (O_1765,N_19406,N_19122);
nand UO_1766 (O_1766,N_19366,N_19556);
or UO_1767 (O_1767,N_19762,N_19062);
nand UO_1768 (O_1768,N_19510,N_19479);
xnor UO_1769 (O_1769,N_19194,N_19534);
nand UO_1770 (O_1770,N_19770,N_19933);
nor UO_1771 (O_1771,N_19036,N_19411);
nand UO_1772 (O_1772,N_19077,N_19878);
nor UO_1773 (O_1773,N_19918,N_19031);
or UO_1774 (O_1774,N_19291,N_19408);
xor UO_1775 (O_1775,N_19044,N_19313);
and UO_1776 (O_1776,N_19718,N_19561);
nor UO_1777 (O_1777,N_19825,N_19110);
or UO_1778 (O_1778,N_19859,N_19579);
xor UO_1779 (O_1779,N_19291,N_19745);
nand UO_1780 (O_1780,N_19589,N_19453);
and UO_1781 (O_1781,N_19228,N_19688);
or UO_1782 (O_1782,N_19234,N_19259);
and UO_1783 (O_1783,N_19580,N_19747);
nor UO_1784 (O_1784,N_19000,N_19661);
and UO_1785 (O_1785,N_19790,N_19017);
and UO_1786 (O_1786,N_19793,N_19703);
and UO_1787 (O_1787,N_19331,N_19568);
or UO_1788 (O_1788,N_19742,N_19223);
or UO_1789 (O_1789,N_19824,N_19556);
nor UO_1790 (O_1790,N_19490,N_19910);
or UO_1791 (O_1791,N_19144,N_19096);
and UO_1792 (O_1792,N_19682,N_19442);
nor UO_1793 (O_1793,N_19627,N_19504);
xnor UO_1794 (O_1794,N_19668,N_19061);
or UO_1795 (O_1795,N_19144,N_19739);
and UO_1796 (O_1796,N_19699,N_19623);
and UO_1797 (O_1797,N_19966,N_19694);
and UO_1798 (O_1798,N_19797,N_19564);
xor UO_1799 (O_1799,N_19789,N_19943);
nor UO_1800 (O_1800,N_19533,N_19687);
nand UO_1801 (O_1801,N_19064,N_19759);
nor UO_1802 (O_1802,N_19153,N_19550);
nor UO_1803 (O_1803,N_19215,N_19247);
xor UO_1804 (O_1804,N_19304,N_19881);
or UO_1805 (O_1805,N_19805,N_19621);
xnor UO_1806 (O_1806,N_19511,N_19963);
nor UO_1807 (O_1807,N_19563,N_19732);
or UO_1808 (O_1808,N_19658,N_19728);
and UO_1809 (O_1809,N_19176,N_19376);
or UO_1810 (O_1810,N_19367,N_19190);
nor UO_1811 (O_1811,N_19890,N_19718);
xnor UO_1812 (O_1812,N_19596,N_19895);
nor UO_1813 (O_1813,N_19970,N_19430);
nor UO_1814 (O_1814,N_19795,N_19473);
nand UO_1815 (O_1815,N_19976,N_19668);
and UO_1816 (O_1816,N_19884,N_19302);
nor UO_1817 (O_1817,N_19657,N_19957);
nand UO_1818 (O_1818,N_19959,N_19608);
and UO_1819 (O_1819,N_19367,N_19400);
nand UO_1820 (O_1820,N_19172,N_19734);
nor UO_1821 (O_1821,N_19097,N_19780);
or UO_1822 (O_1822,N_19025,N_19809);
or UO_1823 (O_1823,N_19812,N_19443);
or UO_1824 (O_1824,N_19364,N_19615);
and UO_1825 (O_1825,N_19347,N_19527);
or UO_1826 (O_1826,N_19890,N_19011);
or UO_1827 (O_1827,N_19762,N_19699);
nand UO_1828 (O_1828,N_19434,N_19594);
nand UO_1829 (O_1829,N_19178,N_19874);
and UO_1830 (O_1830,N_19953,N_19502);
nand UO_1831 (O_1831,N_19044,N_19006);
and UO_1832 (O_1832,N_19739,N_19124);
and UO_1833 (O_1833,N_19770,N_19110);
xnor UO_1834 (O_1834,N_19860,N_19935);
nor UO_1835 (O_1835,N_19373,N_19942);
nand UO_1836 (O_1836,N_19069,N_19216);
xor UO_1837 (O_1837,N_19274,N_19517);
and UO_1838 (O_1838,N_19159,N_19610);
or UO_1839 (O_1839,N_19278,N_19001);
or UO_1840 (O_1840,N_19499,N_19178);
nor UO_1841 (O_1841,N_19960,N_19947);
nor UO_1842 (O_1842,N_19216,N_19235);
and UO_1843 (O_1843,N_19759,N_19641);
and UO_1844 (O_1844,N_19248,N_19137);
nand UO_1845 (O_1845,N_19723,N_19365);
and UO_1846 (O_1846,N_19147,N_19796);
and UO_1847 (O_1847,N_19591,N_19139);
and UO_1848 (O_1848,N_19741,N_19046);
nand UO_1849 (O_1849,N_19495,N_19353);
and UO_1850 (O_1850,N_19181,N_19820);
or UO_1851 (O_1851,N_19488,N_19728);
or UO_1852 (O_1852,N_19592,N_19322);
or UO_1853 (O_1853,N_19736,N_19446);
or UO_1854 (O_1854,N_19803,N_19306);
nor UO_1855 (O_1855,N_19461,N_19009);
xnor UO_1856 (O_1856,N_19764,N_19523);
and UO_1857 (O_1857,N_19255,N_19140);
nand UO_1858 (O_1858,N_19988,N_19310);
or UO_1859 (O_1859,N_19055,N_19863);
xor UO_1860 (O_1860,N_19516,N_19327);
nor UO_1861 (O_1861,N_19170,N_19612);
nand UO_1862 (O_1862,N_19491,N_19596);
and UO_1863 (O_1863,N_19385,N_19830);
and UO_1864 (O_1864,N_19164,N_19730);
nor UO_1865 (O_1865,N_19715,N_19088);
or UO_1866 (O_1866,N_19482,N_19886);
or UO_1867 (O_1867,N_19365,N_19446);
or UO_1868 (O_1868,N_19599,N_19074);
and UO_1869 (O_1869,N_19864,N_19416);
nand UO_1870 (O_1870,N_19908,N_19100);
or UO_1871 (O_1871,N_19235,N_19872);
or UO_1872 (O_1872,N_19801,N_19513);
nand UO_1873 (O_1873,N_19009,N_19801);
or UO_1874 (O_1874,N_19971,N_19235);
nand UO_1875 (O_1875,N_19367,N_19927);
and UO_1876 (O_1876,N_19295,N_19282);
nor UO_1877 (O_1877,N_19352,N_19165);
or UO_1878 (O_1878,N_19823,N_19676);
or UO_1879 (O_1879,N_19018,N_19842);
nor UO_1880 (O_1880,N_19049,N_19011);
nand UO_1881 (O_1881,N_19836,N_19002);
nand UO_1882 (O_1882,N_19171,N_19281);
and UO_1883 (O_1883,N_19386,N_19892);
nand UO_1884 (O_1884,N_19410,N_19096);
and UO_1885 (O_1885,N_19560,N_19233);
or UO_1886 (O_1886,N_19202,N_19151);
nand UO_1887 (O_1887,N_19182,N_19527);
or UO_1888 (O_1888,N_19575,N_19046);
or UO_1889 (O_1889,N_19433,N_19033);
and UO_1890 (O_1890,N_19289,N_19531);
and UO_1891 (O_1891,N_19383,N_19434);
and UO_1892 (O_1892,N_19840,N_19979);
xor UO_1893 (O_1893,N_19127,N_19292);
nor UO_1894 (O_1894,N_19624,N_19448);
and UO_1895 (O_1895,N_19955,N_19644);
and UO_1896 (O_1896,N_19963,N_19165);
or UO_1897 (O_1897,N_19330,N_19553);
xor UO_1898 (O_1898,N_19762,N_19465);
nand UO_1899 (O_1899,N_19229,N_19212);
nor UO_1900 (O_1900,N_19244,N_19286);
xor UO_1901 (O_1901,N_19594,N_19405);
nor UO_1902 (O_1902,N_19662,N_19543);
nor UO_1903 (O_1903,N_19976,N_19472);
or UO_1904 (O_1904,N_19617,N_19395);
nor UO_1905 (O_1905,N_19981,N_19579);
nor UO_1906 (O_1906,N_19292,N_19540);
nand UO_1907 (O_1907,N_19846,N_19109);
nor UO_1908 (O_1908,N_19347,N_19061);
nand UO_1909 (O_1909,N_19497,N_19116);
and UO_1910 (O_1910,N_19202,N_19964);
or UO_1911 (O_1911,N_19882,N_19260);
nor UO_1912 (O_1912,N_19545,N_19658);
and UO_1913 (O_1913,N_19540,N_19937);
or UO_1914 (O_1914,N_19837,N_19831);
xnor UO_1915 (O_1915,N_19081,N_19072);
or UO_1916 (O_1916,N_19824,N_19107);
nor UO_1917 (O_1917,N_19721,N_19281);
nor UO_1918 (O_1918,N_19609,N_19728);
nand UO_1919 (O_1919,N_19934,N_19353);
nand UO_1920 (O_1920,N_19832,N_19815);
xnor UO_1921 (O_1921,N_19283,N_19286);
or UO_1922 (O_1922,N_19920,N_19619);
nand UO_1923 (O_1923,N_19401,N_19474);
and UO_1924 (O_1924,N_19323,N_19263);
or UO_1925 (O_1925,N_19469,N_19443);
xnor UO_1926 (O_1926,N_19483,N_19616);
or UO_1927 (O_1927,N_19665,N_19807);
nand UO_1928 (O_1928,N_19870,N_19792);
nand UO_1929 (O_1929,N_19838,N_19225);
and UO_1930 (O_1930,N_19737,N_19011);
xnor UO_1931 (O_1931,N_19940,N_19838);
nor UO_1932 (O_1932,N_19574,N_19152);
or UO_1933 (O_1933,N_19450,N_19934);
or UO_1934 (O_1934,N_19733,N_19767);
xor UO_1935 (O_1935,N_19390,N_19485);
nor UO_1936 (O_1936,N_19837,N_19073);
nor UO_1937 (O_1937,N_19208,N_19383);
and UO_1938 (O_1938,N_19899,N_19988);
xnor UO_1939 (O_1939,N_19626,N_19937);
or UO_1940 (O_1940,N_19017,N_19597);
nor UO_1941 (O_1941,N_19498,N_19773);
nand UO_1942 (O_1942,N_19033,N_19858);
and UO_1943 (O_1943,N_19049,N_19649);
and UO_1944 (O_1944,N_19563,N_19295);
nor UO_1945 (O_1945,N_19478,N_19378);
nor UO_1946 (O_1946,N_19287,N_19503);
nor UO_1947 (O_1947,N_19516,N_19263);
and UO_1948 (O_1948,N_19570,N_19058);
and UO_1949 (O_1949,N_19858,N_19083);
and UO_1950 (O_1950,N_19335,N_19738);
nand UO_1951 (O_1951,N_19714,N_19923);
nor UO_1952 (O_1952,N_19860,N_19441);
or UO_1953 (O_1953,N_19953,N_19903);
or UO_1954 (O_1954,N_19432,N_19508);
nand UO_1955 (O_1955,N_19047,N_19882);
nor UO_1956 (O_1956,N_19031,N_19607);
nand UO_1957 (O_1957,N_19004,N_19703);
nor UO_1958 (O_1958,N_19445,N_19238);
and UO_1959 (O_1959,N_19740,N_19889);
nor UO_1960 (O_1960,N_19471,N_19321);
nand UO_1961 (O_1961,N_19090,N_19951);
nor UO_1962 (O_1962,N_19111,N_19980);
and UO_1963 (O_1963,N_19277,N_19915);
xor UO_1964 (O_1964,N_19051,N_19836);
and UO_1965 (O_1965,N_19303,N_19297);
or UO_1966 (O_1966,N_19458,N_19172);
nor UO_1967 (O_1967,N_19860,N_19747);
nor UO_1968 (O_1968,N_19620,N_19793);
xor UO_1969 (O_1969,N_19015,N_19632);
and UO_1970 (O_1970,N_19665,N_19899);
or UO_1971 (O_1971,N_19515,N_19528);
or UO_1972 (O_1972,N_19511,N_19353);
or UO_1973 (O_1973,N_19212,N_19333);
or UO_1974 (O_1974,N_19810,N_19666);
and UO_1975 (O_1975,N_19286,N_19689);
xor UO_1976 (O_1976,N_19074,N_19757);
and UO_1977 (O_1977,N_19647,N_19142);
nand UO_1978 (O_1978,N_19146,N_19099);
nand UO_1979 (O_1979,N_19481,N_19648);
and UO_1980 (O_1980,N_19418,N_19317);
or UO_1981 (O_1981,N_19871,N_19319);
nor UO_1982 (O_1982,N_19767,N_19453);
or UO_1983 (O_1983,N_19443,N_19944);
or UO_1984 (O_1984,N_19352,N_19385);
nor UO_1985 (O_1985,N_19804,N_19967);
or UO_1986 (O_1986,N_19556,N_19968);
nand UO_1987 (O_1987,N_19147,N_19972);
and UO_1988 (O_1988,N_19937,N_19616);
nand UO_1989 (O_1989,N_19992,N_19757);
or UO_1990 (O_1990,N_19661,N_19058);
nand UO_1991 (O_1991,N_19969,N_19294);
xnor UO_1992 (O_1992,N_19202,N_19029);
or UO_1993 (O_1993,N_19953,N_19563);
nor UO_1994 (O_1994,N_19502,N_19981);
xor UO_1995 (O_1995,N_19343,N_19600);
nor UO_1996 (O_1996,N_19076,N_19242);
nor UO_1997 (O_1997,N_19446,N_19981);
nand UO_1998 (O_1998,N_19264,N_19509);
xnor UO_1999 (O_1999,N_19149,N_19730);
and UO_2000 (O_2000,N_19982,N_19208);
or UO_2001 (O_2001,N_19180,N_19431);
and UO_2002 (O_2002,N_19226,N_19977);
xnor UO_2003 (O_2003,N_19335,N_19141);
or UO_2004 (O_2004,N_19662,N_19825);
nand UO_2005 (O_2005,N_19510,N_19080);
nor UO_2006 (O_2006,N_19966,N_19251);
and UO_2007 (O_2007,N_19137,N_19028);
nand UO_2008 (O_2008,N_19668,N_19079);
or UO_2009 (O_2009,N_19028,N_19219);
and UO_2010 (O_2010,N_19434,N_19691);
or UO_2011 (O_2011,N_19683,N_19107);
nand UO_2012 (O_2012,N_19634,N_19813);
nand UO_2013 (O_2013,N_19638,N_19112);
nand UO_2014 (O_2014,N_19204,N_19462);
and UO_2015 (O_2015,N_19531,N_19486);
xnor UO_2016 (O_2016,N_19065,N_19952);
nand UO_2017 (O_2017,N_19815,N_19716);
nand UO_2018 (O_2018,N_19598,N_19584);
and UO_2019 (O_2019,N_19071,N_19709);
or UO_2020 (O_2020,N_19414,N_19333);
or UO_2021 (O_2021,N_19788,N_19249);
or UO_2022 (O_2022,N_19041,N_19281);
or UO_2023 (O_2023,N_19646,N_19566);
xnor UO_2024 (O_2024,N_19024,N_19383);
or UO_2025 (O_2025,N_19830,N_19726);
xor UO_2026 (O_2026,N_19355,N_19423);
nor UO_2027 (O_2027,N_19614,N_19285);
nor UO_2028 (O_2028,N_19259,N_19481);
nand UO_2029 (O_2029,N_19787,N_19783);
nor UO_2030 (O_2030,N_19759,N_19145);
or UO_2031 (O_2031,N_19731,N_19679);
nand UO_2032 (O_2032,N_19423,N_19732);
nand UO_2033 (O_2033,N_19475,N_19346);
and UO_2034 (O_2034,N_19754,N_19476);
and UO_2035 (O_2035,N_19371,N_19442);
or UO_2036 (O_2036,N_19574,N_19577);
or UO_2037 (O_2037,N_19117,N_19611);
or UO_2038 (O_2038,N_19891,N_19716);
nor UO_2039 (O_2039,N_19716,N_19074);
nand UO_2040 (O_2040,N_19412,N_19005);
and UO_2041 (O_2041,N_19270,N_19490);
nand UO_2042 (O_2042,N_19557,N_19009);
nand UO_2043 (O_2043,N_19520,N_19829);
or UO_2044 (O_2044,N_19560,N_19932);
or UO_2045 (O_2045,N_19176,N_19654);
or UO_2046 (O_2046,N_19822,N_19109);
nand UO_2047 (O_2047,N_19033,N_19286);
or UO_2048 (O_2048,N_19050,N_19984);
or UO_2049 (O_2049,N_19157,N_19925);
nor UO_2050 (O_2050,N_19257,N_19987);
or UO_2051 (O_2051,N_19559,N_19772);
nor UO_2052 (O_2052,N_19087,N_19241);
xnor UO_2053 (O_2053,N_19214,N_19466);
and UO_2054 (O_2054,N_19855,N_19320);
xor UO_2055 (O_2055,N_19477,N_19587);
nand UO_2056 (O_2056,N_19764,N_19110);
and UO_2057 (O_2057,N_19751,N_19968);
nor UO_2058 (O_2058,N_19819,N_19688);
nand UO_2059 (O_2059,N_19673,N_19091);
nand UO_2060 (O_2060,N_19077,N_19449);
or UO_2061 (O_2061,N_19601,N_19283);
or UO_2062 (O_2062,N_19798,N_19696);
and UO_2063 (O_2063,N_19125,N_19304);
and UO_2064 (O_2064,N_19326,N_19463);
nand UO_2065 (O_2065,N_19915,N_19101);
or UO_2066 (O_2066,N_19489,N_19818);
or UO_2067 (O_2067,N_19444,N_19039);
or UO_2068 (O_2068,N_19721,N_19224);
and UO_2069 (O_2069,N_19615,N_19842);
nand UO_2070 (O_2070,N_19626,N_19967);
and UO_2071 (O_2071,N_19125,N_19190);
or UO_2072 (O_2072,N_19126,N_19940);
nor UO_2073 (O_2073,N_19582,N_19145);
nor UO_2074 (O_2074,N_19553,N_19304);
nand UO_2075 (O_2075,N_19790,N_19918);
nor UO_2076 (O_2076,N_19623,N_19477);
and UO_2077 (O_2077,N_19328,N_19565);
and UO_2078 (O_2078,N_19306,N_19671);
nor UO_2079 (O_2079,N_19522,N_19011);
xnor UO_2080 (O_2080,N_19559,N_19507);
or UO_2081 (O_2081,N_19157,N_19449);
nand UO_2082 (O_2082,N_19917,N_19186);
and UO_2083 (O_2083,N_19090,N_19008);
and UO_2084 (O_2084,N_19355,N_19433);
and UO_2085 (O_2085,N_19729,N_19004);
nor UO_2086 (O_2086,N_19531,N_19253);
nand UO_2087 (O_2087,N_19658,N_19676);
nand UO_2088 (O_2088,N_19439,N_19993);
nand UO_2089 (O_2089,N_19138,N_19530);
nand UO_2090 (O_2090,N_19986,N_19121);
or UO_2091 (O_2091,N_19555,N_19837);
or UO_2092 (O_2092,N_19242,N_19236);
nand UO_2093 (O_2093,N_19294,N_19786);
nand UO_2094 (O_2094,N_19959,N_19122);
xor UO_2095 (O_2095,N_19130,N_19324);
or UO_2096 (O_2096,N_19227,N_19186);
and UO_2097 (O_2097,N_19436,N_19973);
and UO_2098 (O_2098,N_19272,N_19852);
xnor UO_2099 (O_2099,N_19425,N_19885);
nor UO_2100 (O_2100,N_19911,N_19700);
or UO_2101 (O_2101,N_19341,N_19467);
nand UO_2102 (O_2102,N_19704,N_19673);
xor UO_2103 (O_2103,N_19062,N_19912);
xor UO_2104 (O_2104,N_19956,N_19728);
and UO_2105 (O_2105,N_19831,N_19852);
nand UO_2106 (O_2106,N_19405,N_19708);
or UO_2107 (O_2107,N_19369,N_19902);
and UO_2108 (O_2108,N_19097,N_19487);
nand UO_2109 (O_2109,N_19452,N_19742);
nor UO_2110 (O_2110,N_19083,N_19675);
nor UO_2111 (O_2111,N_19279,N_19913);
and UO_2112 (O_2112,N_19215,N_19462);
nand UO_2113 (O_2113,N_19588,N_19774);
and UO_2114 (O_2114,N_19630,N_19309);
and UO_2115 (O_2115,N_19696,N_19312);
and UO_2116 (O_2116,N_19406,N_19993);
nor UO_2117 (O_2117,N_19232,N_19355);
and UO_2118 (O_2118,N_19924,N_19429);
xor UO_2119 (O_2119,N_19316,N_19943);
xor UO_2120 (O_2120,N_19305,N_19484);
and UO_2121 (O_2121,N_19559,N_19043);
nor UO_2122 (O_2122,N_19042,N_19645);
nor UO_2123 (O_2123,N_19833,N_19865);
nand UO_2124 (O_2124,N_19192,N_19531);
nand UO_2125 (O_2125,N_19940,N_19507);
nand UO_2126 (O_2126,N_19566,N_19497);
and UO_2127 (O_2127,N_19403,N_19522);
or UO_2128 (O_2128,N_19208,N_19114);
or UO_2129 (O_2129,N_19054,N_19875);
xor UO_2130 (O_2130,N_19322,N_19938);
nor UO_2131 (O_2131,N_19644,N_19674);
nor UO_2132 (O_2132,N_19993,N_19713);
and UO_2133 (O_2133,N_19973,N_19664);
or UO_2134 (O_2134,N_19552,N_19486);
nand UO_2135 (O_2135,N_19947,N_19489);
nand UO_2136 (O_2136,N_19626,N_19899);
nand UO_2137 (O_2137,N_19114,N_19033);
nand UO_2138 (O_2138,N_19506,N_19619);
or UO_2139 (O_2139,N_19840,N_19178);
and UO_2140 (O_2140,N_19336,N_19667);
xnor UO_2141 (O_2141,N_19627,N_19167);
nand UO_2142 (O_2142,N_19053,N_19781);
or UO_2143 (O_2143,N_19171,N_19650);
or UO_2144 (O_2144,N_19142,N_19295);
nor UO_2145 (O_2145,N_19211,N_19149);
nand UO_2146 (O_2146,N_19123,N_19261);
or UO_2147 (O_2147,N_19996,N_19592);
or UO_2148 (O_2148,N_19141,N_19672);
and UO_2149 (O_2149,N_19057,N_19462);
nand UO_2150 (O_2150,N_19302,N_19352);
nor UO_2151 (O_2151,N_19603,N_19445);
or UO_2152 (O_2152,N_19135,N_19426);
nor UO_2153 (O_2153,N_19528,N_19964);
or UO_2154 (O_2154,N_19883,N_19187);
nor UO_2155 (O_2155,N_19092,N_19689);
or UO_2156 (O_2156,N_19970,N_19501);
nor UO_2157 (O_2157,N_19939,N_19448);
nand UO_2158 (O_2158,N_19628,N_19382);
or UO_2159 (O_2159,N_19151,N_19687);
or UO_2160 (O_2160,N_19749,N_19929);
xnor UO_2161 (O_2161,N_19201,N_19289);
or UO_2162 (O_2162,N_19777,N_19519);
nand UO_2163 (O_2163,N_19913,N_19288);
nand UO_2164 (O_2164,N_19288,N_19258);
nor UO_2165 (O_2165,N_19967,N_19585);
nor UO_2166 (O_2166,N_19980,N_19860);
xor UO_2167 (O_2167,N_19869,N_19590);
nor UO_2168 (O_2168,N_19025,N_19603);
nand UO_2169 (O_2169,N_19105,N_19644);
nand UO_2170 (O_2170,N_19559,N_19476);
or UO_2171 (O_2171,N_19884,N_19892);
and UO_2172 (O_2172,N_19331,N_19821);
nand UO_2173 (O_2173,N_19274,N_19567);
and UO_2174 (O_2174,N_19405,N_19155);
nor UO_2175 (O_2175,N_19761,N_19399);
nor UO_2176 (O_2176,N_19112,N_19765);
nor UO_2177 (O_2177,N_19075,N_19113);
nor UO_2178 (O_2178,N_19107,N_19010);
nand UO_2179 (O_2179,N_19213,N_19491);
nand UO_2180 (O_2180,N_19559,N_19598);
and UO_2181 (O_2181,N_19847,N_19448);
and UO_2182 (O_2182,N_19746,N_19119);
or UO_2183 (O_2183,N_19525,N_19199);
nor UO_2184 (O_2184,N_19112,N_19848);
xor UO_2185 (O_2185,N_19323,N_19080);
nor UO_2186 (O_2186,N_19340,N_19346);
and UO_2187 (O_2187,N_19924,N_19947);
nand UO_2188 (O_2188,N_19839,N_19060);
and UO_2189 (O_2189,N_19065,N_19955);
and UO_2190 (O_2190,N_19767,N_19355);
nor UO_2191 (O_2191,N_19350,N_19325);
nor UO_2192 (O_2192,N_19633,N_19724);
nor UO_2193 (O_2193,N_19707,N_19438);
and UO_2194 (O_2194,N_19592,N_19545);
nand UO_2195 (O_2195,N_19075,N_19820);
xor UO_2196 (O_2196,N_19041,N_19768);
nor UO_2197 (O_2197,N_19175,N_19494);
or UO_2198 (O_2198,N_19831,N_19290);
nor UO_2199 (O_2199,N_19075,N_19151);
and UO_2200 (O_2200,N_19745,N_19606);
nor UO_2201 (O_2201,N_19995,N_19872);
nand UO_2202 (O_2202,N_19845,N_19208);
xnor UO_2203 (O_2203,N_19517,N_19591);
and UO_2204 (O_2204,N_19851,N_19658);
nand UO_2205 (O_2205,N_19798,N_19377);
nor UO_2206 (O_2206,N_19852,N_19338);
or UO_2207 (O_2207,N_19795,N_19643);
nor UO_2208 (O_2208,N_19571,N_19636);
or UO_2209 (O_2209,N_19200,N_19952);
nand UO_2210 (O_2210,N_19373,N_19179);
or UO_2211 (O_2211,N_19531,N_19578);
nand UO_2212 (O_2212,N_19725,N_19334);
xnor UO_2213 (O_2213,N_19534,N_19048);
or UO_2214 (O_2214,N_19905,N_19100);
nor UO_2215 (O_2215,N_19528,N_19939);
and UO_2216 (O_2216,N_19329,N_19739);
and UO_2217 (O_2217,N_19118,N_19335);
or UO_2218 (O_2218,N_19604,N_19228);
or UO_2219 (O_2219,N_19647,N_19552);
nand UO_2220 (O_2220,N_19387,N_19375);
and UO_2221 (O_2221,N_19645,N_19793);
and UO_2222 (O_2222,N_19643,N_19682);
or UO_2223 (O_2223,N_19198,N_19304);
and UO_2224 (O_2224,N_19027,N_19456);
nor UO_2225 (O_2225,N_19350,N_19547);
or UO_2226 (O_2226,N_19974,N_19852);
or UO_2227 (O_2227,N_19397,N_19726);
and UO_2228 (O_2228,N_19252,N_19537);
nand UO_2229 (O_2229,N_19385,N_19925);
nand UO_2230 (O_2230,N_19123,N_19237);
xnor UO_2231 (O_2231,N_19449,N_19594);
and UO_2232 (O_2232,N_19151,N_19477);
and UO_2233 (O_2233,N_19437,N_19722);
nand UO_2234 (O_2234,N_19289,N_19500);
nand UO_2235 (O_2235,N_19012,N_19767);
nor UO_2236 (O_2236,N_19987,N_19800);
xor UO_2237 (O_2237,N_19736,N_19549);
nor UO_2238 (O_2238,N_19272,N_19529);
nand UO_2239 (O_2239,N_19086,N_19234);
and UO_2240 (O_2240,N_19652,N_19883);
and UO_2241 (O_2241,N_19956,N_19039);
nor UO_2242 (O_2242,N_19518,N_19962);
or UO_2243 (O_2243,N_19551,N_19385);
nand UO_2244 (O_2244,N_19911,N_19360);
nor UO_2245 (O_2245,N_19919,N_19333);
nor UO_2246 (O_2246,N_19041,N_19098);
or UO_2247 (O_2247,N_19743,N_19671);
nand UO_2248 (O_2248,N_19567,N_19877);
and UO_2249 (O_2249,N_19326,N_19032);
or UO_2250 (O_2250,N_19227,N_19245);
and UO_2251 (O_2251,N_19660,N_19688);
nor UO_2252 (O_2252,N_19739,N_19301);
or UO_2253 (O_2253,N_19117,N_19710);
nor UO_2254 (O_2254,N_19734,N_19281);
and UO_2255 (O_2255,N_19456,N_19927);
nor UO_2256 (O_2256,N_19376,N_19727);
or UO_2257 (O_2257,N_19751,N_19972);
or UO_2258 (O_2258,N_19176,N_19295);
nand UO_2259 (O_2259,N_19010,N_19577);
or UO_2260 (O_2260,N_19573,N_19425);
nand UO_2261 (O_2261,N_19128,N_19230);
or UO_2262 (O_2262,N_19226,N_19065);
or UO_2263 (O_2263,N_19369,N_19635);
or UO_2264 (O_2264,N_19342,N_19670);
nand UO_2265 (O_2265,N_19582,N_19914);
nand UO_2266 (O_2266,N_19304,N_19009);
nor UO_2267 (O_2267,N_19661,N_19577);
xnor UO_2268 (O_2268,N_19381,N_19643);
xor UO_2269 (O_2269,N_19758,N_19115);
nor UO_2270 (O_2270,N_19213,N_19951);
nor UO_2271 (O_2271,N_19715,N_19792);
nor UO_2272 (O_2272,N_19979,N_19779);
and UO_2273 (O_2273,N_19819,N_19206);
and UO_2274 (O_2274,N_19769,N_19203);
nand UO_2275 (O_2275,N_19420,N_19787);
or UO_2276 (O_2276,N_19562,N_19265);
and UO_2277 (O_2277,N_19040,N_19867);
nand UO_2278 (O_2278,N_19772,N_19334);
nand UO_2279 (O_2279,N_19403,N_19096);
nand UO_2280 (O_2280,N_19340,N_19371);
nand UO_2281 (O_2281,N_19607,N_19040);
xor UO_2282 (O_2282,N_19284,N_19904);
xnor UO_2283 (O_2283,N_19731,N_19874);
nand UO_2284 (O_2284,N_19818,N_19189);
or UO_2285 (O_2285,N_19116,N_19465);
or UO_2286 (O_2286,N_19504,N_19700);
and UO_2287 (O_2287,N_19304,N_19280);
and UO_2288 (O_2288,N_19999,N_19074);
or UO_2289 (O_2289,N_19450,N_19039);
nand UO_2290 (O_2290,N_19820,N_19709);
xnor UO_2291 (O_2291,N_19603,N_19405);
nand UO_2292 (O_2292,N_19771,N_19325);
or UO_2293 (O_2293,N_19205,N_19497);
or UO_2294 (O_2294,N_19285,N_19024);
or UO_2295 (O_2295,N_19119,N_19504);
and UO_2296 (O_2296,N_19039,N_19471);
nor UO_2297 (O_2297,N_19262,N_19264);
nand UO_2298 (O_2298,N_19979,N_19142);
nor UO_2299 (O_2299,N_19326,N_19885);
nand UO_2300 (O_2300,N_19211,N_19072);
and UO_2301 (O_2301,N_19948,N_19101);
xnor UO_2302 (O_2302,N_19555,N_19316);
and UO_2303 (O_2303,N_19705,N_19734);
or UO_2304 (O_2304,N_19911,N_19609);
or UO_2305 (O_2305,N_19870,N_19165);
and UO_2306 (O_2306,N_19609,N_19022);
nand UO_2307 (O_2307,N_19588,N_19722);
and UO_2308 (O_2308,N_19956,N_19115);
nand UO_2309 (O_2309,N_19400,N_19158);
or UO_2310 (O_2310,N_19517,N_19329);
nor UO_2311 (O_2311,N_19552,N_19720);
nor UO_2312 (O_2312,N_19455,N_19254);
or UO_2313 (O_2313,N_19396,N_19201);
and UO_2314 (O_2314,N_19366,N_19183);
nor UO_2315 (O_2315,N_19583,N_19482);
nand UO_2316 (O_2316,N_19149,N_19677);
nand UO_2317 (O_2317,N_19980,N_19726);
nor UO_2318 (O_2318,N_19285,N_19662);
and UO_2319 (O_2319,N_19153,N_19862);
or UO_2320 (O_2320,N_19378,N_19833);
and UO_2321 (O_2321,N_19285,N_19307);
nor UO_2322 (O_2322,N_19558,N_19622);
nor UO_2323 (O_2323,N_19385,N_19726);
and UO_2324 (O_2324,N_19346,N_19168);
or UO_2325 (O_2325,N_19713,N_19305);
xor UO_2326 (O_2326,N_19843,N_19745);
nand UO_2327 (O_2327,N_19385,N_19236);
or UO_2328 (O_2328,N_19951,N_19654);
xor UO_2329 (O_2329,N_19586,N_19516);
or UO_2330 (O_2330,N_19258,N_19611);
nand UO_2331 (O_2331,N_19380,N_19909);
nor UO_2332 (O_2332,N_19221,N_19523);
nor UO_2333 (O_2333,N_19884,N_19564);
nand UO_2334 (O_2334,N_19592,N_19138);
nor UO_2335 (O_2335,N_19433,N_19691);
xor UO_2336 (O_2336,N_19743,N_19238);
and UO_2337 (O_2337,N_19081,N_19840);
or UO_2338 (O_2338,N_19363,N_19801);
and UO_2339 (O_2339,N_19066,N_19489);
or UO_2340 (O_2340,N_19494,N_19908);
and UO_2341 (O_2341,N_19329,N_19798);
and UO_2342 (O_2342,N_19826,N_19480);
nor UO_2343 (O_2343,N_19510,N_19326);
xor UO_2344 (O_2344,N_19447,N_19148);
nand UO_2345 (O_2345,N_19294,N_19830);
or UO_2346 (O_2346,N_19139,N_19191);
xnor UO_2347 (O_2347,N_19493,N_19041);
or UO_2348 (O_2348,N_19545,N_19188);
or UO_2349 (O_2349,N_19401,N_19064);
or UO_2350 (O_2350,N_19995,N_19210);
or UO_2351 (O_2351,N_19674,N_19542);
nor UO_2352 (O_2352,N_19014,N_19553);
nand UO_2353 (O_2353,N_19694,N_19843);
nand UO_2354 (O_2354,N_19354,N_19326);
nand UO_2355 (O_2355,N_19406,N_19585);
nand UO_2356 (O_2356,N_19176,N_19022);
and UO_2357 (O_2357,N_19182,N_19482);
or UO_2358 (O_2358,N_19938,N_19819);
nor UO_2359 (O_2359,N_19341,N_19873);
nor UO_2360 (O_2360,N_19188,N_19547);
nand UO_2361 (O_2361,N_19159,N_19144);
nor UO_2362 (O_2362,N_19376,N_19604);
nor UO_2363 (O_2363,N_19885,N_19288);
nor UO_2364 (O_2364,N_19925,N_19754);
nand UO_2365 (O_2365,N_19433,N_19597);
and UO_2366 (O_2366,N_19164,N_19957);
and UO_2367 (O_2367,N_19615,N_19504);
or UO_2368 (O_2368,N_19962,N_19106);
or UO_2369 (O_2369,N_19826,N_19664);
xor UO_2370 (O_2370,N_19513,N_19965);
nor UO_2371 (O_2371,N_19342,N_19613);
xor UO_2372 (O_2372,N_19372,N_19862);
nand UO_2373 (O_2373,N_19270,N_19050);
nand UO_2374 (O_2374,N_19834,N_19388);
nor UO_2375 (O_2375,N_19887,N_19970);
nand UO_2376 (O_2376,N_19471,N_19996);
and UO_2377 (O_2377,N_19316,N_19587);
nand UO_2378 (O_2378,N_19545,N_19860);
or UO_2379 (O_2379,N_19099,N_19912);
nor UO_2380 (O_2380,N_19235,N_19732);
nor UO_2381 (O_2381,N_19929,N_19823);
and UO_2382 (O_2382,N_19864,N_19376);
nor UO_2383 (O_2383,N_19505,N_19877);
or UO_2384 (O_2384,N_19286,N_19223);
xnor UO_2385 (O_2385,N_19358,N_19120);
or UO_2386 (O_2386,N_19805,N_19009);
or UO_2387 (O_2387,N_19579,N_19738);
nor UO_2388 (O_2388,N_19103,N_19871);
and UO_2389 (O_2389,N_19600,N_19840);
nand UO_2390 (O_2390,N_19769,N_19086);
nor UO_2391 (O_2391,N_19455,N_19012);
and UO_2392 (O_2392,N_19415,N_19074);
nor UO_2393 (O_2393,N_19156,N_19409);
or UO_2394 (O_2394,N_19518,N_19166);
and UO_2395 (O_2395,N_19333,N_19738);
or UO_2396 (O_2396,N_19297,N_19037);
nor UO_2397 (O_2397,N_19935,N_19043);
nor UO_2398 (O_2398,N_19054,N_19490);
nor UO_2399 (O_2399,N_19562,N_19089);
nand UO_2400 (O_2400,N_19755,N_19921);
and UO_2401 (O_2401,N_19102,N_19958);
xnor UO_2402 (O_2402,N_19323,N_19154);
nor UO_2403 (O_2403,N_19830,N_19794);
nor UO_2404 (O_2404,N_19403,N_19627);
nor UO_2405 (O_2405,N_19827,N_19997);
nand UO_2406 (O_2406,N_19380,N_19073);
nor UO_2407 (O_2407,N_19977,N_19389);
xnor UO_2408 (O_2408,N_19993,N_19211);
or UO_2409 (O_2409,N_19287,N_19442);
or UO_2410 (O_2410,N_19083,N_19082);
or UO_2411 (O_2411,N_19348,N_19167);
nand UO_2412 (O_2412,N_19176,N_19409);
xor UO_2413 (O_2413,N_19503,N_19006);
or UO_2414 (O_2414,N_19081,N_19068);
nand UO_2415 (O_2415,N_19906,N_19284);
or UO_2416 (O_2416,N_19813,N_19278);
and UO_2417 (O_2417,N_19610,N_19774);
nand UO_2418 (O_2418,N_19317,N_19549);
nor UO_2419 (O_2419,N_19123,N_19615);
or UO_2420 (O_2420,N_19251,N_19319);
and UO_2421 (O_2421,N_19058,N_19648);
and UO_2422 (O_2422,N_19700,N_19532);
and UO_2423 (O_2423,N_19335,N_19555);
or UO_2424 (O_2424,N_19372,N_19830);
or UO_2425 (O_2425,N_19818,N_19517);
nor UO_2426 (O_2426,N_19100,N_19961);
nor UO_2427 (O_2427,N_19176,N_19901);
nor UO_2428 (O_2428,N_19547,N_19969);
and UO_2429 (O_2429,N_19909,N_19317);
nor UO_2430 (O_2430,N_19050,N_19630);
nor UO_2431 (O_2431,N_19994,N_19222);
and UO_2432 (O_2432,N_19219,N_19423);
nor UO_2433 (O_2433,N_19582,N_19876);
nor UO_2434 (O_2434,N_19687,N_19900);
nand UO_2435 (O_2435,N_19426,N_19591);
nor UO_2436 (O_2436,N_19155,N_19206);
nor UO_2437 (O_2437,N_19156,N_19902);
and UO_2438 (O_2438,N_19679,N_19770);
or UO_2439 (O_2439,N_19767,N_19592);
nand UO_2440 (O_2440,N_19330,N_19996);
and UO_2441 (O_2441,N_19303,N_19688);
and UO_2442 (O_2442,N_19504,N_19866);
nand UO_2443 (O_2443,N_19148,N_19274);
nor UO_2444 (O_2444,N_19836,N_19106);
nor UO_2445 (O_2445,N_19748,N_19470);
xnor UO_2446 (O_2446,N_19548,N_19047);
and UO_2447 (O_2447,N_19175,N_19974);
or UO_2448 (O_2448,N_19283,N_19041);
nand UO_2449 (O_2449,N_19036,N_19777);
and UO_2450 (O_2450,N_19162,N_19882);
or UO_2451 (O_2451,N_19821,N_19833);
or UO_2452 (O_2452,N_19516,N_19757);
and UO_2453 (O_2453,N_19334,N_19739);
and UO_2454 (O_2454,N_19084,N_19342);
or UO_2455 (O_2455,N_19671,N_19423);
nor UO_2456 (O_2456,N_19135,N_19435);
or UO_2457 (O_2457,N_19234,N_19820);
or UO_2458 (O_2458,N_19198,N_19534);
or UO_2459 (O_2459,N_19539,N_19181);
nor UO_2460 (O_2460,N_19773,N_19172);
nand UO_2461 (O_2461,N_19070,N_19817);
nand UO_2462 (O_2462,N_19780,N_19705);
xor UO_2463 (O_2463,N_19153,N_19877);
nand UO_2464 (O_2464,N_19411,N_19066);
or UO_2465 (O_2465,N_19755,N_19083);
nor UO_2466 (O_2466,N_19131,N_19878);
nor UO_2467 (O_2467,N_19036,N_19582);
nand UO_2468 (O_2468,N_19737,N_19352);
nor UO_2469 (O_2469,N_19821,N_19269);
or UO_2470 (O_2470,N_19452,N_19870);
and UO_2471 (O_2471,N_19423,N_19583);
or UO_2472 (O_2472,N_19478,N_19529);
or UO_2473 (O_2473,N_19136,N_19593);
and UO_2474 (O_2474,N_19232,N_19535);
nand UO_2475 (O_2475,N_19198,N_19804);
nor UO_2476 (O_2476,N_19602,N_19208);
nand UO_2477 (O_2477,N_19595,N_19928);
or UO_2478 (O_2478,N_19829,N_19903);
nand UO_2479 (O_2479,N_19843,N_19291);
nand UO_2480 (O_2480,N_19650,N_19360);
nand UO_2481 (O_2481,N_19839,N_19633);
xnor UO_2482 (O_2482,N_19090,N_19629);
nand UO_2483 (O_2483,N_19272,N_19653);
and UO_2484 (O_2484,N_19067,N_19546);
or UO_2485 (O_2485,N_19882,N_19642);
nor UO_2486 (O_2486,N_19151,N_19404);
nor UO_2487 (O_2487,N_19125,N_19006);
and UO_2488 (O_2488,N_19987,N_19692);
nor UO_2489 (O_2489,N_19981,N_19292);
nor UO_2490 (O_2490,N_19948,N_19259);
or UO_2491 (O_2491,N_19711,N_19280);
nor UO_2492 (O_2492,N_19288,N_19647);
and UO_2493 (O_2493,N_19203,N_19236);
nand UO_2494 (O_2494,N_19122,N_19786);
or UO_2495 (O_2495,N_19386,N_19626);
or UO_2496 (O_2496,N_19270,N_19572);
and UO_2497 (O_2497,N_19015,N_19054);
xor UO_2498 (O_2498,N_19270,N_19736);
xnor UO_2499 (O_2499,N_19937,N_19487);
endmodule