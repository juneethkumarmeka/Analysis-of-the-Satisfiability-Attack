module basic_1500_15000_2000_20_levels_10xor_9(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999;
or U0 (N_0,In_1371,In_930);
or U1 (N_1,In_824,In_610);
or U2 (N_2,In_888,In_682);
and U3 (N_3,In_492,In_306);
or U4 (N_4,In_1168,In_431);
nor U5 (N_5,In_599,In_889);
and U6 (N_6,In_1259,In_1192);
and U7 (N_7,In_1461,In_157);
and U8 (N_8,In_329,In_146);
and U9 (N_9,In_1488,In_1026);
xnor U10 (N_10,In_669,In_818);
and U11 (N_11,In_229,In_1060);
and U12 (N_12,In_35,In_1012);
and U13 (N_13,In_1317,In_558);
nor U14 (N_14,In_1092,In_23);
nor U15 (N_15,In_21,In_1122);
or U16 (N_16,In_1398,In_445);
nor U17 (N_17,In_619,In_1491);
xnor U18 (N_18,In_112,In_8);
nand U19 (N_19,In_688,In_1016);
or U20 (N_20,In_410,In_1209);
or U21 (N_21,In_426,In_1089);
and U22 (N_22,In_743,In_508);
and U23 (N_23,In_1311,In_1276);
nand U24 (N_24,In_311,In_368);
xnor U25 (N_25,In_862,In_1391);
and U26 (N_26,In_654,In_524);
xnor U27 (N_27,In_1352,In_1431);
xnor U28 (N_28,In_603,In_335);
and U29 (N_29,In_1250,In_167);
and U30 (N_30,In_886,In_559);
or U31 (N_31,In_830,In_1284);
and U32 (N_32,In_276,In_119);
or U33 (N_33,In_1437,In_580);
and U34 (N_34,In_1077,In_1109);
nor U35 (N_35,In_1331,In_20);
and U36 (N_36,In_1085,In_677);
nor U37 (N_37,In_142,In_759);
nand U38 (N_38,In_435,In_623);
or U39 (N_39,In_239,In_339);
nor U40 (N_40,In_790,In_348);
xnor U41 (N_41,In_513,In_1161);
and U42 (N_42,In_796,In_1141);
or U43 (N_43,In_1131,In_952);
xor U44 (N_44,In_547,In_185);
or U45 (N_45,In_355,In_1345);
nor U46 (N_46,In_337,In_177);
nor U47 (N_47,In_1421,In_1434);
or U48 (N_48,In_984,In_483);
nor U49 (N_49,In_75,In_200);
and U50 (N_50,In_582,In_913);
or U51 (N_51,In_1307,In_140);
and U52 (N_52,In_845,In_1022);
or U53 (N_53,In_327,In_1083);
xor U54 (N_54,In_264,In_1356);
or U55 (N_55,In_243,In_648);
xnor U56 (N_56,In_979,In_707);
nor U57 (N_57,In_434,In_39);
and U58 (N_58,In_217,In_1279);
and U59 (N_59,In_250,In_531);
xnor U60 (N_60,In_838,In_1001);
and U61 (N_61,In_1258,In_381);
nor U62 (N_62,In_1393,In_1466);
nor U63 (N_63,In_1353,In_1441);
or U64 (N_64,In_461,In_812);
nor U65 (N_65,In_1002,In_73);
nand U66 (N_66,In_620,In_1385);
xnor U67 (N_67,In_1329,In_55);
nor U68 (N_68,In_174,In_1357);
and U69 (N_69,In_338,In_1127);
nand U70 (N_70,In_937,In_615);
xor U71 (N_71,In_220,In_585);
nor U72 (N_72,In_85,In_132);
nor U73 (N_73,In_1006,In_1333);
and U74 (N_74,In_501,In_999);
nand U75 (N_75,In_1492,In_1087);
nor U76 (N_76,In_877,In_923);
and U77 (N_77,In_609,In_1283);
or U78 (N_78,In_636,In_423);
and U79 (N_79,In_1302,In_295);
nor U80 (N_80,In_725,In_716);
and U81 (N_81,In_965,In_1478);
nor U82 (N_82,In_933,In_641);
or U83 (N_83,In_265,In_1113);
xor U84 (N_84,In_1040,In_735);
xor U85 (N_85,In_367,In_454);
and U86 (N_86,In_991,In_980);
xor U87 (N_87,In_1303,In_1145);
xor U88 (N_88,In_496,In_864);
and U89 (N_89,In_439,In_542);
or U90 (N_90,In_60,In_450);
and U91 (N_91,In_831,In_1044);
nor U92 (N_92,In_419,In_386);
nor U93 (N_93,In_113,In_594);
nor U94 (N_94,In_1110,In_491);
nor U95 (N_95,In_750,In_42);
nand U96 (N_96,In_874,In_65);
or U97 (N_97,In_315,In_429);
nand U98 (N_98,In_593,In_1163);
nor U99 (N_99,In_15,In_216);
nand U100 (N_100,In_98,In_6);
nor U101 (N_101,In_1170,In_1452);
and U102 (N_102,In_689,In_36);
or U103 (N_103,In_354,In_1414);
or U104 (N_104,In_145,In_1337);
nor U105 (N_105,In_126,In_813);
xor U106 (N_106,In_1041,In_987);
nand U107 (N_107,In_94,In_983);
nand U108 (N_108,In_1201,In_1156);
nor U109 (N_109,In_1378,In_1249);
nand U110 (N_110,In_822,In_1397);
and U111 (N_111,In_189,In_127);
nand U112 (N_112,In_1342,In_883);
nor U113 (N_113,In_1082,In_639);
nor U114 (N_114,In_770,In_388);
nand U115 (N_115,In_690,In_309);
or U116 (N_116,In_463,In_1182);
or U117 (N_117,In_522,In_97);
nand U118 (N_118,In_1216,In_941);
nor U119 (N_119,In_89,In_499);
xnor U120 (N_120,In_901,In_1227);
or U121 (N_121,In_1212,In_296);
nor U122 (N_122,In_884,In_130);
xnor U123 (N_123,In_22,In_76);
xor U124 (N_124,In_717,In_184);
and U125 (N_125,In_1103,In_1467);
or U126 (N_126,In_1166,In_227);
nand U127 (N_127,In_61,In_872);
nand U128 (N_128,In_573,In_695);
nand U129 (N_129,In_1314,In_906);
xnor U130 (N_130,In_737,In_403);
nor U131 (N_131,In_789,In_665);
and U132 (N_132,In_1052,In_782);
and U133 (N_133,In_986,In_1328);
nand U134 (N_134,In_1149,In_1334);
nor U135 (N_135,In_1305,In_821);
and U136 (N_136,In_494,In_1154);
nor U137 (N_137,In_1453,In_938);
or U138 (N_138,In_588,In_1118);
and U139 (N_139,In_27,In_1176);
nor U140 (N_140,In_1230,In_1389);
or U141 (N_141,In_1396,In_597);
or U142 (N_142,In_702,In_963);
or U143 (N_143,In_175,In_135);
nor U144 (N_144,In_579,In_1386);
and U145 (N_145,In_1120,In_618);
and U146 (N_146,In_521,In_951);
and U147 (N_147,In_940,In_1003);
and U148 (N_148,In_482,In_754);
and U149 (N_149,In_826,In_659);
nand U150 (N_150,In_964,In_263);
or U151 (N_151,In_846,In_51);
nor U152 (N_152,In_260,In_1290);
or U153 (N_153,In_24,In_545);
and U154 (N_154,In_54,In_658);
and U155 (N_155,In_1320,In_1462);
or U156 (N_156,In_1394,In_170);
nor U157 (N_157,In_1099,In_1031);
nor U158 (N_158,In_1050,In_1197);
nand U159 (N_159,In_430,In_387);
nor U160 (N_160,In_141,In_1335);
and U161 (N_161,In_854,In_324);
nand U162 (N_162,In_1056,In_977);
nand U163 (N_163,In_1173,In_875);
nor U164 (N_164,In_129,In_396);
nand U165 (N_165,In_171,In_709);
nor U166 (N_166,In_108,In_481);
or U167 (N_167,In_314,In_458);
nand U168 (N_168,In_116,In_749);
nor U169 (N_169,In_1440,In_520);
or U170 (N_170,In_1098,In_93);
nor U171 (N_171,In_536,In_614);
nor U172 (N_172,In_1379,In_1436);
nand U173 (N_173,In_1446,In_1313);
xnor U174 (N_174,In_313,In_131);
xor U175 (N_175,In_1009,In_277);
or U176 (N_176,In_1175,In_1377);
and U177 (N_177,In_882,In_803);
nor U178 (N_178,In_880,In_261);
and U179 (N_179,In_456,In_1021);
or U180 (N_180,In_1341,In_621);
xnor U181 (N_181,In_1047,In_1494);
or U182 (N_182,In_1285,In_385);
xnor U183 (N_183,In_1151,In_1429);
and U184 (N_184,In_606,In_1366);
or U185 (N_185,In_612,In_776);
xnor U186 (N_186,In_172,In_19);
and U187 (N_187,In_562,In_553);
xnor U188 (N_188,In_1264,In_369);
nand U189 (N_189,In_257,In_820);
or U190 (N_190,In_1088,In_1220);
or U191 (N_191,In_1454,In_713);
or U192 (N_192,In_595,In_62);
xor U193 (N_193,In_507,In_1194);
nor U194 (N_194,In_288,In_397);
and U195 (N_195,In_225,In_7);
nor U196 (N_196,In_152,In_78);
or U197 (N_197,In_490,In_527);
xnor U198 (N_198,In_258,In_1306);
xor U199 (N_199,In_356,In_32);
xor U200 (N_200,In_1256,In_1435);
nand U201 (N_201,In_729,In_1024);
nor U202 (N_202,In_1346,In_100);
nand U203 (N_203,In_1097,In_1210);
and U204 (N_204,In_996,In_52);
or U205 (N_205,In_405,In_926);
xnor U206 (N_206,In_1057,In_1215);
nand U207 (N_207,In_896,In_625);
or U208 (N_208,In_462,In_164);
and U209 (N_209,In_498,In_742);
nand U210 (N_210,In_406,In_190);
nand U211 (N_211,In_59,In_331);
xnor U212 (N_212,In_968,In_1233);
xor U213 (N_213,In_1196,In_985);
nor U214 (N_214,In_1301,In_5);
xnor U215 (N_215,In_392,In_1028);
nand U216 (N_216,In_851,In_829);
xnor U217 (N_217,In_1254,In_1029);
xnor U218 (N_218,In_245,In_230);
xnor U219 (N_219,In_179,In_1180);
nor U220 (N_220,In_891,In_664);
nor U221 (N_221,In_566,In_109);
nand U222 (N_222,In_569,In_26);
nand U223 (N_223,In_765,In_640);
nand U224 (N_224,In_394,In_1030);
and U225 (N_225,In_1105,In_1291);
nand U226 (N_226,In_298,In_1229);
and U227 (N_227,In_767,In_1075);
nor U228 (N_228,In_262,In_1046);
or U229 (N_229,In_687,In_916);
nand U230 (N_230,In_681,In_1292);
nor U231 (N_231,In_256,In_325);
xor U232 (N_232,In_1117,In_638);
nor U233 (N_233,In_350,In_1179);
nand U234 (N_234,In_1235,In_819);
and U235 (N_235,In_1142,In_777);
or U236 (N_236,In_857,In_342);
nand U237 (N_237,In_1253,In_1493);
or U238 (N_238,In_535,In_911);
nand U239 (N_239,In_804,In_1222);
or U240 (N_240,In_756,In_1130);
xnor U241 (N_241,In_1344,In_1255);
and U242 (N_242,In_351,In_1094);
nand U243 (N_243,In_1204,In_675);
nand U244 (N_244,In_74,In_1164);
xor U245 (N_245,In_914,In_1458);
nor U246 (N_246,In_917,In_575);
nor U247 (N_247,In_1382,In_753);
xor U248 (N_248,In_652,In_1199);
nor U249 (N_249,In_1277,In_1160);
nand U250 (N_250,In_607,In_1020);
and U251 (N_251,In_115,In_193);
or U252 (N_252,In_866,In_1239);
nor U253 (N_253,In_438,In_1497);
and U254 (N_254,In_412,In_995);
xor U255 (N_255,In_1084,In_1295);
xor U256 (N_256,In_312,In_835);
or U257 (N_257,In_349,In_653);
xor U258 (N_258,In_904,In_376);
or U259 (N_259,In_1426,In_511);
nand U260 (N_260,In_1129,In_817);
nand U261 (N_261,In_541,In_495);
nand U262 (N_262,In_485,In_1079);
xnor U263 (N_263,In_981,In_876);
or U264 (N_264,In_1489,In_897);
or U265 (N_265,In_576,In_1420);
nor U266 (N_266,In_422,In_1217);
xnor U267 (N_267,In_488,In_1469);
or U268 (N_268,In_1401,In_165);
nor U269 (N_269,In_1240,In_1365);
or U270 (N_270,In_12,In_365);
xnor U271 (N_271,In_973,In_45);
nand U272 (N_272,In_1416,In_1051);
nand U273 (N_273,In_453,In_158);
nor U274 (N_274,In_1459,In_960);
and U275 (N_275,In_253,In_1043);
or U276 (N_276,In_379,In_752);
nor U277 (N_277,In_1177,In_1274);
or U278 (N_278,In_841,In_1281);
nand U279 (N_279,In_1372,In_711);
or U280 (N_280,In_87,In_117);
xor U281 (N_281,In_371,In_1315);
or U282 (N_282,In_989,In_358);
nor U283 (N_283,In_443,In_291);
xnor U284 (N_284,In_909,In_1045);
nand U285 (N_285,In_186,In_939);
and U286 (N_286,In_1450,In_228);
xnor U287 (N_287,In_1287,In_1018);
xnor U288 (N_288,In_798,In_1428);
or U289 (N_289,In_465,In_332);
nor U290 (N_290,In_1399,In_57);
xor U291 (N_291,In_255,In_1412);
nor U292 (N_292,In_1390,In_642);
or U293 (N_293,In_532,In_953);
and U294 (N_294,In_807,In_1464);
nand U295 (N_295,In_670,In_1107);
xor U296 (N_296,In_219,In_1178);
and U297 (N_297,In_1112,In_71);
and U298 (N_298,In_278,In_894);
and U299 (N_299,In_279,In_1269);
nand U300 (N_300,In_994,In_971);
xnor U301 (N_301,In_353,In_699);
and U302 (N_302,In_1247,In_70);
nand U303 (N_303,In_178,In_10);
nand U304 (N_304,In_1387,In_630);
xor U305 (N_305,In_201,In_209);
nand U306 (N_306,In_758,In_283);
or U307 (N_307,In_714,In_604);
nor U308 (N_308,In_544,In_1361);
or U309 (N_309,In_294,In_746);
xor U310 (N_310,In_757,In_802);
or U311 (N_311,In_328,In_517);
nor U312 (N_312,In_1388,In_961);
nor U313 (N_313,In_668,In_137);
and U314 (N_314,In_235,In_0);
or U315 (N_315,In_823,In_134);
and U316 (N_316,In_44,In_899);
or U317 (N_317,In_334,In_732);
xor U318 (N_318,In_210,In_469);
xor U319 (N_319,In_751,In_221);
nand U320 (N_320,In_236,In_155);
xnor U321 (N_321,In_608,In_1340);
or U322 (N_322,In_878,In_1165);
nand U323 (N_323,In_691,In_160);
and U324 (N_324,In_417,In_1147);
or U325 (N_325,In_159,In_1409);
xor U326 (N_326,In_203,In_853);
xnor U327 (N_327,In_1169,In_107);
xor U328 (N_328,In_869,In_1095);
nor U329 (N_329,In_1066,In_176);
and U330 (N_330,In_705,In_676);
xor U331 (N_331,In_449,In_370);
xor U332 (N_332,In_962,In_1309);
xor U333 (N_333,In_970,In_246);
or U334 (N_334,In_247,In_304);
nand U335 (N_335,In_1481,In_1336);
nand U336 (N_336,In_447,In_1139);
xnor U337 (N_337,In_811,In_1096);
nor U338 (N_338,In_254,In_1424);
or U339 (N_339,In_847,In_1271);
and U340 (N_340,In_1000,In_111);
nand U341 (N_341,In_459,In_58);
nor U342 (N_342,In_881,In_95);
and U343 (N_343,In_1392,In_708);
and U344 (N_344,In_663,In_323);
and U345 (N_345,In_444,In_1486);
xnor U346 (N_346,In_1368,In_46);
xnor U347 (N_347,In_634,In_448);
or U348 (N_348,In_816,In_395);
and U349 (N_349,In_1081,In_1187);
nand U350 (N_350,In_1495,In_1438);
xor U351 (N_351,In_617,In_1144);
and U352 (N_352,In_733,In_1137);
xor U353 (N_353,In_1153,In_269);
nor U354 (N_354,In_1260,In_762);
nand U355 (N_355,In_336,In_53);
xnor U356 (N_356,In_69,In_1069);
and U357 (N_357,In_1119,In_934);
nand U358 (N_358,In_105,In_515);
nand U359 (N_359,In_967,In_801);
nor U360 (N_360,In_982,In_738);
xor U361 (N_361,In_950,In_1064);
nand U362 (N_362,In_679,In_928);
and U363 (N_363,In_290,In_487);
nor U364 (N_364,In_144,In_834);
nand U365 (N_365,In_1327,In_921);
nand U366 (N_366,In_139,In_249);
nand U367 (N_367,In_800,In_516);
and U368 (N_368,In_1067,In_1432);
xor U369 (N_369,In_919,In_1423);
nand U370 (N_370,In_760,In_1411);
xnor U371 (N_371,In_404,In_1267);
nor U372 (N_372,In_1244,In_202);
or U373 (N_373,In_840,In_1415);
nand U374 (N_374,In_627,In_1054);
xor U375 (N_375,In_451,In_1148);
or U376 (N_376,In_30,In_1116);
or U377 (N_377,In_543,In_1228);
and U378 (N_378,In_268,In_1484);
xor U379 (N_379,In_1351,In_1004);
xnor U380 (N_380,In_104,In_194);
nand U381 (N_381,In_446,In_285);
nand U382 (N_382,In_442,In_468);
xor U383 (N_383,In_478,In_1332);
nor U384 (N_384,In_374,In_1155);
or U385 (N_385,In_1111,In_726);
or U386 (N_386,In_557,In_1482);
nand U387 (N_387,In_1465,In_136);
or U388 (N_388,In_1405,In_1483);
or U389 (N_389,In_18,In_1070);
or U390 (N_390,In_143,In_859);
xor U391 (N_391,In_584,In_1027);
and U392 (N_392,In_359,In_34);
nand U393 (N_393,In_616,In_1299);
xnor U394 (N_394,In_1471,In_1174);
or U395 (N_395,In_797,In_724);
nand U396 (N_396,In_121,In_1364);
and U397 (N_397,In_1451,In_280);
or U398 (N_398,In_1207,In_3);
nand U399 (N_399,In_740,In_1055);
or U400 (N_400,In_924,In_1310);
nor U401 (N_401,In_704,In_432);
and U402 (N_402,In_1190,In_972);
and U403 (N_403,In_583,In_25);
and U404 (N_404,In_1140,In_825);
or U405 (N_405,In_282,In_715);
nor U406 (N_406,In_90,In_734);
xor U407 (N_407,In_151,In_223);
xor U408 (N_408,In_993,In_1363);
nor U409 (N_409,In_848,In_1380);
or U410 (N_410,In_915,In_945);
xnor U411 (N_411,In_1203,In_769);
or U412 (N_412,In_1101,In_1049);
nor U413 (N_413,In_427,In_787);
xor U414 (N_414,In_666,In_480);
and U415 (N_415,In_600,In_86);
or U416 (N_416,In_1286,In_975);
xor U417 (N_417,In_920,In_944);
or U418 (N_418,In_1133,In_1456);
xnor U419 (N_419,In_1410,In_1433);
nand U420 (N_420,In_1039,In_1183);
or U421 (N_421,In_1078,In_457);
or U422 (N_422,In_150,In_533);
nand U423 (N_423,In_763,In_645);
nand U424 (N_424,In_123,In_1257);
nor U425 (N_425,In_384,In_50);
or U426 (N_426,In_635,In_362);
and U427 (N_427,In_1498,In_377);
nor U428 (N_428,In_156,In_1293);
nand U429 (N_429,In_1134,In_1487);
or U430 (N_430,In_844,In_651);
and U431 (N_431,In_748,In_1205);
or U432 (N_432,In_401,In_1172);
xor U433 (N_433,In_340,In_680);
nor U434 (N_434,In_1062,In_997);
and U435 (N_435,In_731,In_1395);
nand U436 (N_436,In_1350,In_101);
or U437 (N_437,In_678,In_273);
nor U438 (N_438,In_1490,In_1157);
xor U439 (N_439,In_1184,In_124);
nor U440 (N_440,In_551,In_1479);
nor U441 (N_441,In_736,In_1065);
nand U442 (N_442,In_1408,In_9);
nand U443 (N_443,In_703,In_650);
nand U444 (N_444,In_561,In_552);
or U445 (N_445,In_719,In_722);
or U446 (N_446,In_1121,In_514);
xnor U447 (N_447,In_655,In_198);
and U448 (N_448,In_577,In_13);
xnor U449 (N_449,In_81,In_942);
and U450 (N_450,In_259,In_601);
nand U451 (N_451,In_380,In_560);
or U452 (N_452,In_320,In_242);
nand U453 (N_453,In_773,In_780);
nand U454 (N_454,In_455,In_550);
xor U455 (N_455,In_281,In_38);
nor U456 (N_456,In_1093,In_460);
nor U457 (N_457,In_37,In_199);
and U458 (N_458,In_1477,In_400);
nand U459 (N_459,In_464,In_1241);
nor U460 (N_460,In_556,In_29);
nor U461 (N_461,In_927,In_205);
or U462 (N_462,In_1444,In_1347);
xnor U463 (N_463,In_1102,In_287);
nand U464 (N_464,In_697,In_477);
and U465 (N_465,In_1403,In_297);
nand U466 (N_466,In_411,In_103);
nand U467 (N_467,In_206,In_855);
or U468 (N_468,In_125,In_540);
nor U469 (N_469,In_1280,In_512);
nor U470 (N_470,In_1015,In_1213);
nor U471 (N_471,In_77,In_1198);
nor U472 (N_472,In_1242,In_1251);
xor U473 (N_473,In_389,In_549);
and U474 (N_474,In_922,In_43);
or U475 (N_475,In_1445,In_1297);
nor U476 (N_476,In_162,In_1090);
and U477 (N_477,In_852,In_504);
nor U478 (N_478,In_212,In_472);
or U479 (N_479,In_1013,In_307);
xor U480 (N_480,In_563,In_525);
or U481 (N_481,In_310,In_1289);
xnor U482 (N_482,In_879,In_433);
xor U483 (N_483,In_694,In_809);
and U484 (N_484,In_1422,In_484);
nand U485 (N_485,In_1246,In_1407);
nand U486 (N_486,In_657,In_1005);
or U487 (N_487,In_1138,In_173);
or U488 (N_488,In_63,In_2);
nand U489 (N_489,In_420,In_503);
or U490 (N_490,In_474,In_1473);
nor U491 (N_491,In_322,In_4);
xor U492 (N_492,In_302,In_318);
or U493 (N_493,In_643,In_624);
nand U494 (N_494,In_300,In_333);
nor U495 (N_495,In_1348,In_161);
and U496 (N_496,In_187,In_1243);
xor U497 (N_497,In_133,In_40);
and U498 (N_498,In_631,In_360);
and U499 (N_499,In_1191,In_873);
xnor U500 (N_500,In_1376,In_272);
nand U501 (N_501,In_436,In_241);
nor U502 (N_502,In_153,In_1496);
and U503 (N_503,In_1017,In_784);
nor U504 (N_504,In_646,In_622);
or U505 (N_505,In_120,In_476);
nand U506 (N_506,In_425,In_1343);
or U507 (N_507,In_122,In_637);
xor U508 (N_508,In_795,In_1234);
or U509 (N_509,In_572,In_856);
xnor U510 (N_510,In_1330,In_728);
and U511 (N_511,In_1036,In_828);
or U512 (N_512,In_958,In_598);
nand U513 (N_513,In_1262,In_118);
or U514 (N_514,In_1032,In_486);
and U515 (N_515,In_1126,In_1374);
nor U516 (N_516,In_1265,In_1418);
nor U517 (N_517,In_505,In_343);
and U518 (N_518,In_741,In_128);
nor U519 (N_519,In_414,In_1188);
xor U520 (N_520,In_966,In_428);
xor U521 (N_521,In_589,In_284);
xor U522 (N_522,In_893,In_378);
nand U523 (N_523,In_195,In_1442);
nand U524 (N_524,In_1007,In_1023);
nor U525 (N_525,In_799,In_571);
and U526 (N_526,In_102,In_1245);
and U527 (N_527,In_110,In_308);
xor U528 (N_528,In_1014,In_827);
nand U529 (N_529,In_632,In_1338);
xnor U530 (N_530,In_605,In_237);
nor U531 (N_531,In_1238,In_305);
nor U532 (N_532,In_602,In_900);
nand U533 (N_533,In_806,In_1288);
xnor U534 (N_534,In_863,In_587);
nand U535 (N_535,In_99,In_1323);
or U536 (N_536,In_935,In_698);
nand U537 (N_537,In_1048,In_674);
nor U538 (N_538,In_1370,In_11);
or U539 (N_539,In_1143,In_895);
or U540 (N_540,In_564,In_500);
nand U541 (N_541,In_363,In_700);
nand U542 (N_542,In_1460,In_502);
or U543 (N_543,In_79,In_1485);
xnor U544 (N_544,In_251,In_41);
nor U545 (N_545,In_1360,In_382);
or U546 (N_546,In_1214,In_792);
or U547 (N_547,In_67,In_570);
nand U548 (N_548,In_1206,In_1402);
xnor U549 (N_549,In_226,In_1275);
and U550 (N_550,In_166,In_667);
nand U551 (N_551,In_91,In_692);
xnor U552 (N_552,In_1189,In_191);
nand U553 (N_553,In_843,In_1339);
nor U554 (N_554,In_418,In_17);
and U555 (N_555,In_509,In_1034);
or U556 (N_556,In_364,In_684);
xor U557 (N_557,In_548,In_832);
and U558 (N_558,In_660,In_1304);
nand U559 (N_559,In_671,In_317);
or U560 (N_560,In_947,In_84);
nor U561 (N_561,In_1294,In_421);
nor U562 (N_562,In_1463,In_718);
nor U563 (N_563,In_788,In_1171);
or U564 (N_564,In_207,In_506);
nand U565 (N_565,In_1162,In_808);
nor U566 (N_566,In_1202,In_860);
nand U567 (N_567,In_1322,In_321);
xor U568 (N_568,In_534,In_530);
or U569 (N_569,In_1058,In_1449);
and U570 (N_570,In_1076,In_1349);
nor U571 (N_571,In_929,In_470);
or U572 (N_572,In_1367,In_1124);
nand U573 (N_573,In_772,In_1167);
nor U574 (N_574,In_274,In_849);
and U575 (N_575,In_1135,In_1221);
and U576 (N_576,In_1358,In_293);
or U577 (N_577,In_344,In_771);
nor U578 (N_578,In_932,In_286);
xor U579 (N_579,In_842,In_1159);
and U580 (N_580,In_1448,In_271);
nand U581 (N_581,In_890,In_778);
xnor U582 (N_582,In_1086,In_526);
nor U583 (N_583,In_685,In_892);
or U584 (N_584,In_64,In_466);
xor U585 (N_585,In_1186,In_147);
or U586 (N_586,In_978,In_416);
or U587 (N_587,In_188,In_390);
and U588 (N_588,In_114,In_538);
xor U589 (N_589,In_836,In_413);
nand U590 (N_590,In_775,In_931);
nand U591 (N_591,In_1455,In_837);
nand U592 (N_592,In_1404,In_907);
or U593 (N_593,In_1324,In_424);
nand U594 (N_594,In_1325,In_786);
and U595 (N_595,In_316,In_528);
and U596 (N_596,In_949,In_1224);
xnor U597 (N_597,In_1226,In_82);
and U598 (N_598,In_218,In_1261);
or U599 (N_599,In_346,In_1232);
or U600 (N_600,In_974,In_1319);
nand U601 (N_601,In_683,In_1080);
nand U602 (N_602,In_347,In_1447);
and U603 (N_603,In_1059,In_661);
nor U604 (N_604,In_903,In_224);
xnor U605 (N_605,In_180,In_647);
xnor U606 (N_606,In_222,In_696);
nor U607 (N_607,In_1270,In_399);
nand U608 (N_608,In_706,In_998);
xor U609 (N_609,In_1146,In_1300);
or U610 (N_610,In_154,In_169);
nor U611 (N_611,In_633,In_568);
and U612 (N_612,In_1298,In_266);
nand U613 (N_613,In_1033,In_192);
nor U614 (N_614,In_629,In_1430);
nand U615 (N_615,In_149,In_1425);
xnor U616 (N_616,In_1115,In_1200);
nand U617 (N_617,In_943,In_1218);
and U618 (N_618,In_745,In_1106);
or U619 (N_619,In_1132,In_275);
and U620 (N_620,In_1181,In_211);
and U621 (N_621,In_1439,In_204);
xnor U622 (N_622,In_805,In_1114);
nor U623 (N_623,In_1355,In_861);
nor U624 (N_624,In_781,In_1068);
xnor U625 (N_625,In_613,In_341);
nand U626 (N_626,In_992,In_592);
or U627 (N_627,In_1359,In_138);
and U628 (N_628,In_1208,In_31);
nor U629 (N_629,In_301,In_898);
nand U630 (N_630,In_299,In_1185);
and U631 (N_631,In_1499,In_814);
or U632 (N_632,In_1211,In_1193);
and U633 (N_633,In_833,In_1072);
xnor U634 (N_634,In_467,In_990);
xor U635 (N_635,In_398,In_649);
and U636 (N_636,In_1266,In_955);
or U637 (N_637,In_106,In_791);
nand U638 (N_638,In_1042,In_723);
nor U639 (N_639,In_49,In_83);
nor U640 (N_640,In_197,In_539);
and U641 (N_641,In_1252,In_72);
or U642 (N_642,In_815,In_1128);
or U643 (N_643,In_946,In_794);
or U644 (N_644,In_1158,In_578);
or U645 (N_645,In_885,In_1231);
nor U646 (N_646,In_783,In_744);
nand U647 (N_647,In_372,In_196);
xor U648 (N_648,In_345,In_415);
and U649 (N_649,In_1108,In_766);
and U650 (N_650,In_440,In_720);
or U651 (N_651,In_574,In_183);
nor U652 (N_652,In_68,In_1318);
xnor U653 (N_653,In_871,In_248);
nand U654 (N_654,In_567,In_1476);
nand U655 (N_655,In_391,In_1470);
xnor U656 (N_656,In_810,In_739);
or U657 (N_657,In_954,In_774);
or U658 (N_658,In_1237,In_1354);
nor U659 (N_659,In_755,In_1104);
and U660 (N_660,In_1400,In_546);
nor U661 (N_661,In_1091,In_1123);
nand U662 (N_662,In_1025,In_918);
nor U663 (N_663,In_867,In_1268);
nor U664 (N_664,In_148,In_1443);
or U665 (N_665,In_510,In_1474);
or U666 (N_666,In_1362,In_710);
nand U667 (N_667,In_1375,In_785);
xor U668 (N_668,In_489,In_1263);
nand U669 (N_669,In_88,In_1413);
nand U670 (N_670,In_870,In_352);
xnor U671 (N_671,In_1011,In_902);
and U672 (N_672,In_252,In_730);
or U673 (N_673,In_473,In_1383);
nor U674 (N_674,In_905,In_858);
or U675 (N_675,In_1321,In_581);
nand U676 (N_676,In_591,In_1417);
nand U677 (N_677,In_1272,In_92);
and U678 (N_678,In_1475,In_330);
nand U679 (N_679,In_497,In_1053);
and U680 (N_680,In_1308,In_936);
or U681 (N_681,In_839,In_1472);
nor U682 (N_682,In_383,In_1316);
or U683 (N_683,In_887,In_270);
nor U684 (N_684,In_693,In_686);
or U685 (N_685,In_292,In_673);
nand U686 (N_686,In_33,In_1);
nand U687 (N_687,In_441,In_1248);
xor U688 (N_688,In_233,In_865);
nor U689 (N_689,In_1195,In_1427);
xor U690 (N_690,In_493,In_409);
nand U691 (N_691,In_1061,In_518);
xnor U692 (N_692,In_644,In_1219);
xor U693 (N_693,In_721,In_361);
or U694 (N_694,In_611,In_244);
nor U695 (N_695,In_590,In_1278);
nand U696 (N_696,In_701,In_240);
nand U697 (N_697,In_1074,In_662);
or U698 (N_698,In_912,In_1152);
and U699 (N_699,In_1480,In_232);
xnor U700 (N_700,In_959,In_850);
nand U701 (N_701,In_214,In_764);
or U702 (N_702,In_868,In_238);
xor U703 (N_703,In_910,In_554);
or U704 (N_704,In_479,In_66);
nor U705 (N_705,In_925,In_957);
and U706 (N_706,In_1019,In_956);
nand U707 (N_707,In_1326,In_1406);
xor U708 (N_708,In_1035,In_779);
xnor U709 (N_709,In_452,In_303);
xor U710 (N_710,In_523,In_373);
nand U711 (N_711,In_1037,In_747);
and U712 (N_712,In_357,In_1236);
xnor U713 (N_713,In_1273,In_1296);
and U714 (N_714,In_366,In_326);
xnor U715 (N_715,In_1225,In_96);
xor U716 (N_716,In_319,In_1223);
or U717 (N_717,In_555,In_14);
xnor U718 (N_718,In_628,In_1100);
xor U719 (N_719,In_1373,In_672);
nand U720 (N_720,In_289,In_208);
nand U721 (N_721,In_475,In_471);
nand U722 (N_722,In_267,In_168);
nand U723 (N_723,In_181,In_626);
and U724 (N_724,In_519,In_407);
nor U725 (N_725,In_402,In_1312);
and U726 (N_726,In_16,In_1008);
nor U727 (N_727,In_28,In_213);
nor U728 (N_728,In_375,In_231);
and U729 (N_729,In_1419,In_48);
and U730 (N_730,In_215,In_565);
xor U731 (N_731,In_1384,In_56);
nor U732 (N_732,In_1125,In_529);
or U733 (N_733,In_908,In_969);
nor U734 (N_734,In_408,In_586);
or U735 (N_735,In_80,In_596);
and U736 (N_736,In_768,In_656);
or U737 (N_737,In_437,In_1071);
nor U738 (N_738,In_182,In_1457);
or U739 (N_739,In_234,In_163);
nand U740 (N_740,In_1073,In_948);
and U741 (N_741,In_1282,In_537);
nor U742 (N_742,In_1468,In_393);
or U743 (N_743,In_1369,In_1063);
and U744 (N_744,In_47,In_1381);
nand U745 (N_745,In_727,In_712);
xnor U746 (N_746,In_1038,In_1010);
nand U747 (N_747,In_761,In_976);
and U748 (N_748,In_988,In_1136);
nor U749 (N_749,In_793,In_1150);
nor U750 (N_750,N_113,N_590);
nand U751 (N_751,N_704,N_609);
xnor U752 (N_752,N_26,N_566);
xor U753 (N_753,N_347,N_735);
nand U754 (N_754,N_409,N_650);
xnor U755 (N_755,N_371,N_660);
xnor U756 (N_756,N_680,N_578);
xor U757 (N_757,N_270,N_728);
or U758 (N_758,N_212,N_730);
nand U759 (N_759,N_537,N_27);
xnor U760 (N_760,N_644,N_96);
nor U761 (N_761,N_277,N_534);
or U762 (N_762,N_60,N_373);
nand U763 (N_763,N_634,N_424);
nand U764 (N_764,N_32,N_444);
nor U765 (N_765,N_86,N_407);
nor U766 (N_766,N_346,N_269);
or U767 (N_767,N_726,N_119);
nor U768 (N_768,N_261,N_125);
xor U769 (N_769,N_29,N_8);
nor U770 (N_770,N_37,N_209);
nor U771 (N_771,N_288,N_619);
xnor U772 (N_772,N_642,N_52);
nor U773 (N_773,N_84,N_106);
xor U774 (N_774,N_232,N_14);
xnor U775 (N_775,N_28,N_602);
and U776 (N_776,N_313,N_394);
or U777 (N_777,N_653,N_46);
nor U778 (N_778,N_18,N_514);
xor U779 (N_779,N_364,N_700);
xnor U780 (N_780,N_562,N_197);
nor U781 (N_781,N_72,N_575);
xnor U782 (N_782,N_250,N_595);
or U783 (N_783,N_41,N_219);
and U784 (N_784,N_607,N_34);
xor U785 (N_785,N_260,N_116);
and U786 (N_786,N_740,N_745);
nand U787 (N_787,N_396,N_658);
xnor U788 (N_788,N_530,N_554);
and U789 (N_789,N_31,N_624);
nor U790 (N_790,N_552,N_45);
or U791 (N_791,N_716,N_92);
xnor U792 (N_792,N_676,N_525);
and U793 (N_793,N_275,N_1);
xor U794 (N_794,N_16,N_421);
or U795 (N_795,N_276,N_128);
xnor U796 (N_796,N_379,N_714);
and U797 (N_797,N_576,N_510);
xor U798 (N_798,N_675,N_312);
or U799 (N_799,N_103,N_494);
and U800 (N_800,N_733,N_83);
xnor U801 (N_801,N_6,N_742);
and U802 (N_802,N_337,N_162);
or U803 (N_803,N_392,N_140);
xor U804 (N_804,N_507,N_249);
or U805 (N_805,N_511,N_329);
nor U806 (N_806,N_647,N_90);
xnor U807 (N_807,N_121,N_251);
nand U808 (N_808,N_520,N_306);
nor U809 (N_809,N_117,N_491);
or U810 (N_810,N_478,N_414);
nor U811 (N_811,N_154,N_199);
nand U812 (N_812,N_341,N_605);
or U813 (N_813,N_406,N_493);
xor U814 (N_814,N_79,N_451);
xor U815 (N_815,N_10,N_701);
xor U816 (N_816,N_105,N_279);
or U817 (N_817,N_588,N_721);
and U818 (N_818,N_725,N_258);
and U819 (N_819,N_599,N_539);
nor U820 (N_820,N_15,N_296);
nor U821 (N_821,N_214,N_57);
nand U822 (N_822,N_354,N_632);
and U823 (N_823,N_321,N_627);
or U824 (N_824,N_230,N_338);
nor U825 (N_825,N_49,N_483);
xnor U826 (N_826,N_12,N_638);
nor U827 (N_827,N_630,N_376);
nor U828 (N_828,N_684,N_666);
nor U829 (N_829,N_692,N_107);
or U830 (N_830,N_21,N_468);
nand U831 (N_831,N_361,N_559);
nor U832 (N_832,N_369,N_355);
nor U833 (N_833,N_293,N_448);
xnor U834 (N_834,N_274,N_727);
nor U835 (N_835,N_59,N_436);
nor U836 (N_836,N_304,N_126);
or U837 (N_837,N_403,N_51);
nor U838 (N_838,N_422,N_343);
nor U839 (N_839,N_150,N_298);
nor U840 (N_840,N_268,N_423);
nor U841 (N_841,N_732,N_583);
xor U842 (N_842,N_368,N_25);
and U843 (N_843,N_487,N_153);
or U844 (N_844,N_340,N_715);
and U845 (N_845,N_694,N_365);
nand U846 (N_846,N_476,N_631);
xnor U847 (N_847,N_486,N_481);
and U848 (N_848,N_617,N_557);
xnor U849 (N_849,N_120,N_0);
nand U850 (N_850,N_538,N_669);
xnor U851 (N_851,N_519,N_523);
nor U852 (N_852,N_189,N_561);
and U853 (N_853,N_683,N_429);
xor U854 (N_854,N_264,N_223);
nor U855 (N_855,N_574,N_245);
or U856 (N_856,N_427,N_563);
or U857 (N_857,N_524,N_101);
nor U858 (N_858,N_362,N_352);
nand U859 (N_859,N_350,N_68);
nor U860 (N_860,N_143,N_235);
or U861 (N_861,N_518,N_351);
and U862 (N_862,N_592,N_673);
nor U863 (N_863,N_78,N_532);
or U864 (N_864,N_73,N_400);
and U865 (N_865,N_213,N_36);
and U866 (N_866,N_85,N_287);
or U867 (N_867,N_504,N_157);
xnor U868 (N_868,N_689,N_316);
and U869 (N_869,N_388,N_513);
nor U870 (N_870,N_332,N_540);
nor U871 (N_871,N_528,N_639);
nor U872 (N_872,N_446,N_185);
or U873 (N_873,N_97,N_109);
nor U874 (N_874,N_170,N_567);
or U875 (N_875,N_431,N_194);
nand U876 (N_876,N_458,N_207);
nor U877 (N_877,N_682,N_267);
and U878 (N_878,N_48,N_211);
nand U879 (N_879,N_734,N_512);
nor U880 (N_880,N_506,N_271);
xnor U881 (N_881,N_98,N_196);
xor U882 (N_882,N_134,N_192);
or U883 (N_883,N_702,N_294);
and U884 (N_884,N_699,N_454);
nand U885 (N_885,N_160,N_404);
and U886 (N_886,N_40,N_178);
xor U887 (N_887,N_501,N_11);
or U888 (N_888,N_174,N_475);
xor U889 (N_889,N_297,N_344);
nor U890 (N_890,N_273,N_254);
nor U891 (N_891,N_42,N_311);
nand U892 (N_892,N_408,N_378);
nand U893 (N_893,N_470,N_142);
nand U894 (N_894,N_241,N_171);
or U895 (N_895,N_257,N_253);
nor U896 (N_896,N_449,N_712);
or U897 (N_897,N_286,N_114);
xnor U898 (N_898,N_353,N_67);
or U899 (N_899,N_248,N_205);
or U900 (N_900,N_147,N_87);
xnor U901 (N_901,N_466,N_179);
and U902 (N_902,N_330,N_44);
or U903 (N_903,N_685,N_224);
or U904 (N_904,N_603,N_262);
nor U905 (N_905,N_225,N_746);
or U906 (N_906,N_442,N_367);
and U907 (N_907,N_710,N_50);
or U908 (N_908,N_22,N_169);
and U909 (N_909,N_697,N_415);
and U910 (N_910,N_227,N_381);
nor U911 (N_911,N_656,N_357);
xnor U912 (N_912,N_457,N_743);
and U913 (N_913,N_281,N_320);
and U914 (N_914,N_594,N_259);
nand U915 (N_915,N_425,N_94);
or U916 (N_916,N_202,N_322);
nor U917 (N_917,N_533,N_687);
nand U918 (N_918,N_272,N_711);
nand U919 (N_919,N_628,N_163);
xnor U920 (N_920,N_318,N_738);
xnor U921 (N_921,N_503,N_399);
and U922 (N_922,N_641,N_593);
xnor U923 (N_923,N_324,N_747);
and U924 (N_924,N_342,N_71);
nand U925 (N_925,N_587,N_488);
xor U926 (N_926,N_233,N_326);
xnor U927 (N_927,N_719,N_244);
xor U928 (N_928,N_579,N_646);
nand U929 (N_929,N_127,N_461);
nor U930 (N_930,N_151,N_645);
nand U931 (N_931,N_323,N_499);
or U932 (N_932,N_53,N_420);
xor U933 (N_933,N_387,N_585);
and U934 (N_934,N_331,N_247);
xor U935 (N_935,N_410,N_548);
xnor U936 (N_936,N_741,N_469);
xnor U937 (N_937,N_496,N_386);
or U938 (N_938,N_455,N_348);
xor U939 (N_939,N_278,N_536);
and U940 (N_940,N_200,N_531);
xor U941 (N_941,N_377,N_345);
nand U942 (N_942,N_139,N_589);
xnor U943 (N_943,N_465,N_584);
or U944 (N_944,N_543,N_623);
nand U945 (N_945,N_58,N_718);
xnor U946 (N_946,N_447,N_416);
nor U947 (N_947,N_222,N_176);
and U948 (N_948,N_191,N_419);
or U949 (N_949,N_74,N_526);
and U950 (N_950,N_598,N_542);
nand U951 (N_951,N_411,N_240);
nor U952 (N_952,N_629,N_636);
xnor U953 (N_953,N_484,N_572);
nor U954 (N_954,N_319,N_314);
nand U955 (N_955,N_678,N_705);
xnor U956 (N_956,N_615,N_545);
and U957 (N_957,N_480,N_691);
nand U958 (N_958,N_145,N_527);
or U959 (N_959,N_604,N_360);
nand U960 (N_960,N_158,N_195);
or U961 (N_961,N_129,N_382);
nor U962 (N_962,N_606,N_502);
nor U963 (N_963,N_662,N_736);
xor U964 (N_964,N_183,N_370);
xor U965 (N_965,N_77,N_359);
and U966 (N_966,N_317,N_130);
nand U967 (N_967,N_621,N_182);
and U968 (N_968,N_155,N_626);
nand U969 (N_969,N_159,N_443);
xor U970 (N_970,N_172,N_608);
and U971 (N_971,N_201,N_556);
or U972 (N_972,N_549,N_450);
nor U973 (N_973,N_460,N_307);
and U974 (N_974,N_81,N_291);
nand U975 (N_975,N_635,N_335);
xnor U976 (N_976,N_23,N_70);
xor U977 (N_977,N_435,N_17);
or U978 (N_978,N_210,N_490);
or U979 (N_979,N_111,N_301);
nand U980 (N_980,N_544,N_66);
and U981 (N_981,N_265,N_110);
xnor U982 (N_982,N_141,N_398);
and U983 (N_983,N_482,N_216);
or U984 (N_984,N_385,N_285);
nor U985 (N_985,N_333,N_280);
nand U986 (N_986,N_62,N_108);
nand U987 (N_987,N_391,N_413);
nor U988 (N_988,N_652,N_156);
nand U989 (N_989,N_664,N_610);
nor U990 (N_990,N_236,N_144);
or U991 (N_991,N_356,N_20);
xnor U992 (N_992,N_184,N_30);
and U993 (N_993,N_464,N_24);
nand U994 (N_994,N_428,N_580);
nor U995 (N_995,N_255,N_167);
and U996 (N_996,N_625,N_439);
or U997 (N_997,N_600,N_440);
or U998 (N_998,N_252,N_437);
nor U999 (N_999,N_180,N_266);
xnor U1000 (N_1000,N_325,N_75);
or U1001 (N_1001,N_495,N_243);
and U1002 (N_1002,N_418,N_591);
or U1003 (N_1003,N_551,N_445);
xnor U1004 (N_1004,N_479,N_681);
xor U1005 (N_1005,N_61,N_375);
nand U1006 (N_1006,N_693,N_80);
xor U1007 (N_1007,N_535,N_723);
or U1008 (N_1008,N_173,N_47);
nor U1009 (N_1009,N_517,N_565);
or U1010 (N_1010,N_299,N_198);
nor U1011 (N_1011,N_568,N_349);
xor U1012 (N_1012,N_614,N_88);
or U1013 (N_1013,N_472,N_115);
and U1014 (N_1014,N_19,N_166);
or U1015 (N_1015,N_165,N_620);
nand U1016 (N_1016,N_674,N_308);
and U1017 (N_1017,N_569,N_739);
nand U1018 (N_1018,N_215,N_263);
nand U1019 (N_1019,N_132,N_69);
nor U1020 (N_1020,N_99,N_521);
nor U1021 (N_1021,N_550,N_206);
nand U1022 (N_1022,N_300,N_405);
xor U1023 (N_1023,N_149,N_168);
or U1024 (N_1024,N_295,N_146);
nor U1025 (N_1025,N_327,N_509);
nand U1026 (N_1026,N_412,N_65);
xor U1027 (N_1027,N_7,N_547);
and U1028 (N_1028,N_655,N_654);
and U1029 (N_1029,N_516,N_616);
and U1030 (N_1030,N_677,N_679);
or U1031 (N_1031,N_695,N_748);
nor U1032 (N_1032,N_402,N_193);
or U1033 (N_1033,N_720,N_383);
and U1034 (N_1034,N_508,N_546);
nand U1035 (N_1035,N_637,N_434);
or U1036 (N_1036,N_438,N_239);
xnor U1037 (N_1037,N_3,N_217);
xnor U1038 (N_1038,N_577,N_133);
nand U1039 (N_1039,N_138,N_100);
nand U1040 (N_1040,N_729,N_724);
or U1041 (N_1041,N_242,N_124);
nand U1042 (N_1042,N_611,N_622);
nor U1043 (N_1043,N_393,N_473);
nand U1044 (N_1044,N_686,N_713);
or U1045 (N_1045,N_722,N_570);
and U1046 (N_1046,N_95,N_175);
nand U1047 (N_1047,N_384,N_238);
xor U1048 (N_1048,N_661,N_148);
nand U1049 (N_1049,N_571,N_82);
nand U1050 (N_1050,N_553,N_459);
xor U1051 (N_1051,N_649,N_35);
or U1052 (N_1052,N_39,N_54);
nand U1053 (N_1053,N_441,N_586);
or U1054 (N_1054,N_485,N_474);
or U1055 (N_1055,N_613,N_43);
nand U1056 (N_1056,N_717,N_374);
and U1057 (N_1057,N_208,N_9);
and U1058 (N_1058,N_703,N_582);
nor U1059 (N_1059,N_237,N_256);
xor U1060 (N_1060,N_515,N_497);
nand U1061 (N_1061,N_395,N_401);
nand U1062 (N_1062,N_112,N_56);
nor U1063 (N_1063,N_136,N_417);
or U1064 (N_1064,N_289,N_453);
xnor U1065 (N_1065,N_492,N_282);
xor U1066 (N_1066,N_33,N_177);
xor U1067 (N_1067,N_529,N_187);
and U1068 (N_1068,N_5,N_505);
xor U1069 (N_1069,N_397,N_618);
xnor U1070 (N_1070,N_389,N_696);
nor U1071 (N_1071,N_284,N_204);
nor U1072 (N_1072,N_597,N_328);
nand U1073 (N_1073,N_737,N_93);
and U1074 (N_1074,N_339,N_456);
or U1075 (N_1075,N_498,N_612);
or U1076 (N_1076,N_670,N_462);
xor U1077 (N_1077,N_663,N_731);
nor U1078 (N_1078,N_63,N_560);
xor U1079 (N_1079,N_643,N_665);
xnor U1080 (N_1080,N_380,N_471);
nand U1081 (N_1081,N_309,N_657);
and U1082 (N_1082,N_601,N_426);
or U1083 (N_1083,N_708,N_477);
xnor U1084 (N_1084,N_432,N_633);
xor U1085 (N_1085,N_188,N_433);
and U1086 (N_1086,N_709,N_659);
or U1087 (N_1087,N_671,N_246);
xnor U1088 (N_1088,N_190,N_500);
nor U1089 (N_1089,N_651,N_334);
nand U1090 (N_1090,N_707,N_231);
nand U1091 (N_1091,N_152,N_89);
xor U1092 (N_1092,N_315,N_290);
xnor U1093 (N_1093,N_161,N_467);
nand U1094 (N_1094,N_672,N_749);
nor U1095 (N_1095,N_310,N_122);
and U1096 (N_1096,N_573,N_303);
nand U1097 (N_1097,N_541,N_302);
nor U1098 (N_1098,N_186,N_688);
xnor U1099 (N_1099,N_118,N_221);
nand U1100 (N_1100,N_363,N_283);
nor U1101 (N_1101,N_104,N_596);
or U1102 (N_1102,N_226,N_430);
or U1103 (N_1103,N_55,N_4);
nand U1104 (N_1104,N_706,N_690);
nor U1105 (N_1105,N_164,N_522);
nand U1106 (N_1106,N_489,N_38);
and U1107 (N_1107,N_220,N_581);
xor U1108 (N_1108,N_76,N_667);
nand U1109 (N_1109,N_137,N_558);
and U1110 (N_1110,N_463,N_668);
xnor U1111 (N_1111,N_64,N_744);
nor U1112 (N_1112,N_131,N_372);
or U1113 (N_1113,N_2,N_390);
xnor U1114 (N_1114,N_181,N_292);
nand U1115 (N_1115,N_564,N_366);
nor U1116 (N_1116,N_640,N_228);
nor U1117 (N_1117,N_555,N_135);
xnor U1118 (N_1118,N_91,N_102);
xor U1119 (N_1119,N_234,N_336);
xor U1120 (N_1120,N_358,N_452);
xor U1121 (N_1121,N_123,N_698);
nand U1122 (N_1122,N_203,N_305);
or U1123 (N_1123,N_13,N_218);
nor U1124 (N_1124,N_648,N_229);
or U1125 (N_1125,N_646,N_693);
and U1126 (N_1126,N_383,N_248);
nand U1127 (N_1127,N_711,N_191);
or U1128 (N_1128,N_1,N_148);
and U1129 (N_1129,N_648,N_696);
nand U1130 (N_1130,N_692,N_452);
nand U1131 (N_1131,N_412,N_644);
nor U1132 (N_1132,N_49,N_213);
or U1133 (N_1133,N_305,N_748);
xnor U1134 (N_1134,N_68,N_700);
or U1135 (N_1135,N_275,N_334);
nand U1136 (N_1136,N_544,N_323);
or U1137 (N_1137,N_652,N_590);
nor U1138 (N_1138,N_180,N_449);
and U1139 (N_1139,N_383,N_567);
and U1140 (N_1140,N_593,N_510);
and U1141 (N_1141,N_627,N_142);
nor U1142 (N_1142,N_341,N_402);
nand U1143 (N_1143,N_737,N_525);
nand U1144 (N_1144,N_227,N_650);
nand U1145 (N_1145,N_649,N_26);
or U1146 (N_1146,N_305,N_632);
or U1147 (N_1147,N_322,N_740);
nor U1148 (N_1148,N_616,N_388);
xnor U1149 (N_1149,N_362,N_652);
or U1150 (N_1150,N_185,N_638);
nor U1151 (N_1151,N_509,N_217);
or U1152 (N_1152,N_640,N_637);
and U1153 (N_1153,N_649,N_246);
nor U1154 (N_1154,N_504,N_384);
xor U1155 (N_1155,N_669,N_505);
xor U1156 (N_1156,N_384,N_129);
nor U1157 (N_1157,N_400,N_331);
nor U1158 (N_1158,N_673,N_723);
or U1159 (N_1159,N_549,N_253);
xor U1160 (N_1160,N_349,N_140);
xor U1161 (N_1161,N_324,N_241);
or U1162 (N_1162,N_58,N_255);
nand U1163 (N_1163,N_666,N_197);
xor U1164 (N_1164,N_631,N_300);
or U1165 (N_1165,N_612,N_526);
xnor U1166 (N_1166,N_174,N_152);
xor U1167 (N_1167,N_455,N_388);
nor U1168 (N_1168,N_122,N_445);
nor U1169 (N_1169,N_159,N_705);
or U1170 (N_1170,N_556,N_672);
nand U1171 (N_1171,N_412,N_735);
and U1172 (N_1172,N_191,N_261);
nor U1173 (N_1173,N_717,N_190);
or U1174 (N_1174,N_118,N_667);
or U1175 (N_1175,N_631,N_353);
xor U1176 (N_1176,N_336,N_558);
and U1177 (N_1177,N_142,N_265);
and U1178 (N_1178,N_238,N_726);
xnor U1179 (N_1179,N_688,N_184);
and U1180 (N_1180,N_112,N_717);
nand U1181 (N_1181,N_397,N_131);
xnor U1182 (N_1182,N_187,N_158);
and U1183 (N_1183,N_221,N_636);
nor U1184 (N_1184,N_48,N_24);
xnor U1185 (N_1185,N_102,N_545);
nor U1186 (N_1186,N_27,N_580);
or U1187 (N_1187,N_3,N_369);
xnor U1188 (N_1188,N_406,N_69);
and U1189 (N_1189,N_120,N_495);
nand U1190 (N_1190,N_467,N_424);
or U1191 (N_1191,N_194,N_348);
and U1192 (N_1192,N_250,N_353);
nand U1193 (N_1193,N_745,N_435);
and U1194 (N_1194,N_337,N_319);
nand U1195 (N_1195,N_110,N_644);
or U1196 (N_1196,N_738,N_382);
xnor U1197 (N_1197,N_262,N_414);
nand U1198 (N_1198,N_257,N_125);
nor U1199 (N_1199,N_180,N_705);
nand U1200 (N_1200,N_200,N_87);
or U1201 (N_1201,N_694,N_661);
and U1202 (N_1202,N_83,N_320);
or U1203 (N_1203,N_534,N_571);
or U1204 (N_1204,N_713,N_485);
nand U1205 (N_1205,N_497,N_123);
nand U1206 (N_1206,N_696,N_621);
nand U1207 (N_1207,N_354,N_427);
or U1208 (N_1208,N_21,N_480);
nand U1209 (N_1209,N_556,N_13);
xor U1210 (N_1210,N_84,N_577);
and U1211 (N_1211,N_280,N_236);
nand U1212 (N_1212,N_151,N_593);
nand U1213 (N_1213,N_637,N_72);
xor U1214 (N_1214,N_489,N_304);
nand U1215 (N_1215,N_686,N_741);
nand U1216 (N_1216,N_432,N_144);
and U1217 (N_1217,N_480,N_442);
nand U1218 (N_1218,N_6,N_349);
nor U1219 (N_1219,N_175,N_29);
nor U1220 (N_1220,N_432,N_214);
or U1221 (N_1221,N_641,N_521);
xor U1222 (N_1222,N_633,N_187);
nor U1223 (N_1223,N_494,N_690);
or U1224 (N_1224,N_517,N_569);
nand U1225 (N_1225,N_737,N_255);
or U1226 (N_1226,N_17,N_442);
nor U1227 (N_1227,N_34,N_114);
nor U1228 (N_1228,N_99,N_81);
or U1229 (N_1229,N_16,N_573);
or U1230 (N_1230,N_552,N_120);
nand U1231 (N_1231,N_670,N_269);
and U1232 (N_1232,N_254,N_189);
and U1233 (N_1233,N_374,N_578);
nor U1234 (N_1234,N_553,N_206);
or U1235 (N_1235,N_449,N_668);
or U1236 (N_1236,N_601,N_124);
or U1237 (N_1237,N_618,N_143);
or U1238 (N_1238,N_641,N_714);
or U1239 (N_1239,N_229,N_347);
or U1240 (N_1240,N_253,N_306);
or U1241 (N_1241,N_681,N_91);
nor U1242 (N_1242,N_306,N_593);
xor U1243 (N_1243,N_549,N_538);
or U1244 (N_1244,N_473,N_448);
or U1245 (N_1245,N_384,N_347);
nor U1246 (N_1246,N_404,N_540);
nor U1247 (N_1247,N_138,N_223);
nor U1248 (N_1248,N_226,N_36);
nor U1249 (N_1249,N_485,N_609);
xnor U1250 (N_1250,N_664,N_324);
nand U1251 (N_1251,N_511,N_63);
and U1252 (N_1252,N_434,N_55);
nor U1253 (N_1253,N_533,N_149);
xor U1254 (N_1254,N_320,N_244);
or U1255 (N_1255,N_551,N_410);
nand U1256 (N_1256,N_161,N_97);
and U1257 (N_1257,N_221,N_206);
and U1258 (N_1258,N_109,N_127);
nand U1259 (N_1259,N_589,N_677);
or U1260 (N_1260,N_690,N_595);
or U1261 (N_1261,N_375,N_726);
xor U1262 (N_1262,N_250,N_288);
and U1263 (N_1263,N_645,N_242);
nand U1264 (N_1264,N_592,N_131);
xor U1265 (N_1265,N_571,N_384);
nand U1266 (N_1266,N_303,N_449);
nor U1267 (N_1267,N_428,N_197);
or U1268 (N_1268,N_303,N_341);
xnor U1269 (N_1269,N_126,N_35);
or U1270 (N_1270,N_635,N_271);
nor U1271 (N_1271,N_465,N_23);
nor U1272 (N_1272,N_262,N_588);
nor U1273 (N_1273,N_419,N_8);
nand U1274 (N_1274,N_677,N_278);
nand U1275 (N_1275,N_341,N_240);
xnor U1276 (N_1276,N_625,N_307);
nor U1277 (N_1277,N_339,N_51);
or U1278 (N_1278,N_379,N_48);
nand U1279 (N_1279,N_326,N_377);
xnor U1280 (N_1280,N_87,N_312);
or U1281 (N_1281,N_467,N_738);
nand U1282 (N_1282,N_558,N_624);
nand U1283 (N_1283,N_394,N_268);
or U1284 (N_1284,N_553,N_34);
or U1285 (N_1285,N_58,N_574);
and U1286 (N_1286,N_731,N_447);
or U1287 (N_1287,N_110,N_675);
nand U1288 (N_1288,N_70,N_61);
nor U1289 (N_1289,N_290,N_178);
and U1290 (N_1290,N_452,N_466);
or U1291 (N_1291,N_37,N_239);
xnor U1292 (N_1292,N_151,N_176);
and U1293 (N_1293,N_93,N_14);
or U1294 (N_1294,N_1,N_472);
nor U1295 (N_1295,N_458,N_699);
nor U1296 (N_1296,N_58,N_287);
and U1297 (N_1297,N_426,N_259);
nand U1298 (N_1298,N_572,N_474);
nor U1299 (N_1299,N_112,N_473);
or U1300 (N_1300,N_181,N_422);
nand U1301 (N_1301,N_287,N_554);
or U1302 (N_1302,N_689,N_343);
xor U1303 (N_1303,N_108,N_267);
nand U1304 (N_1304,N_103,N_738);
nor U1305 (N_1305,N_565,N_505);
and U1306 (N_1306,N_378,N_267);
and U1307 (N_1307,N_466,N_170);
xor U1308 (N_1308,N_328,N_603);
nor U1309 (N_1309,N_88,N_385);
and U1310 (N_1310,N_605,N_710);
nand U1311 (N_1311,N_652,N_592);
and U1312 (N_1312,N_232,N_258);
or U1313 (N_1313,N_438,N_638);
xnor U1314 (N_1314,N_93,N_744);
nand U1315 (N_1315,N_589,N_257);
and U1316 (N_1316,N_72,N_712);
or U1317 (N_1317,N_280,N_413);
or U1318 (N_1318,N_227,N_611);
or U1319 (N_1319,N_338,N_718);
or U1320 (N_1320,N_634,N_673);
or U1321 (N_1321,N_437,N_215);
or U1322 (N_1322,N_135,N_52);
xor U1323 (N_1323,N_728,N_69);
nand U1324 (N_1324,N_256,N_654);
nor U1325 (N_1325,N_598,N_421);
nor U1326 (N_1326,N_181,N_110);
or U1327 (N_1327,N_560,N_228);
nand U1328 (N_1328,N_734,N_201);
and U1329 (N_1329,N_209,N_355);
xnor U1330 (N_1330,N_415,N_5);
or U1331 (N_1331,N_352,N_439);
xnor U1332 (N_1332,N_272,N_155);
or U1333 (N_1333,N_295,N_422);
nor U1334 (N_1334,N_451,N_37);
nor U1335 (N_1335,N_416,N_576);
or U1336 (N_1336,N_143,N_328);
and U1337 (N_1337,N_587,N_27);
nand U1338 (N_1338,N_159,N_445);
and U1339 (N_1339,N_105,N_648);
and U1340 (N_1340,N_642,N_472);
nand U1341 (N_1341,N_144,N_194);
and U1342 (N_1342,N_508,N_513);
xor U1343 (N_1343,N_515,N_401);
xnor U1344 (N_1344,N_236,N_499);
and U1345 (N_1345,N_236,N_304);
nor U1346 (N_1346,N_627,N_312);
or U1347 (N_1347,N_648,N_405);
xor U1348 (N_1348,N_151,N_350);
xor U1349 (N_1349,N_738,N_705);
or U1350 (N_1350,N_263,N_267);
xor U1351 (N_1351,N_485,N_653);
xnor U1352 (N_1352,N_731,N_295);
and U1353 (N_1353,N_257,N_399);
xnor U1354 (N_1354,N_458,N_288);
nand U1355 (N_1355,N_613,N_362);
and U1356 (N_1356,N_265,N_427);
xor U1357 (N_1357,N_173,N_604);
and U1358 (N_1358,N_477,N_384);
and U1359 (N_1359,N_363,N_163);
or U1360 (N_1360,N_676,N_276);
xor U1361 (N_1361,N_97,N_349);
nor U1362 (N_1362,N_557,N_225);
and U1363 (N_1363,N_652,N_70);
or U1364 (N_1364,N_719,N_251);
or U1365 (N_1365,N_286,N_186);
xor U1366 (N_1366,N_706,N_155);
or U1367 (N_1367,N_283,N_532);
nand U1368 (N_1368,N_708,N_441);
nand U1369 (N_1369,N_176,N_312);
nor U1370 (N_1370,N_684,N_621);
xnor U1371 (N_1371,N_486,N_238);
xnor U1372 (N_1372,N_222,N_266);
and U1373 (N_1373,N_397,N_320);
or U1374 (N_1374,N_702,N_550);
or U1375 (N_1375,N_554,N_458);
nor U1376 (N_1376,N_110,N_585);
and U1377 (N_1377,N_329,N_242);
nor U1378 (N_1378,N_746,N_715);
xor U1379 (N_1379,N_434,N_213);
and U1380 (N_1380,N_226,N_623);
xor U1381 (N_1381,N_554,N_228);
and U1382 (N_1382,N_723,N_7);
or U1383 (N_1383,N_597,N_292);
xor U1384 (N_1384,N_655,N_62);
xnor U1385 (N_1385,N_711,N_484);
nor U1386 (N_1386,N_740,N_439);
xnor U1387 (N_1387,N_472,N_244);
xnor U1388 (N_1388,N_365,N_378);
xnor U1389 (N_1389,N_497,N_114);
or U1390 (N_1390,N_745,N_181);
and U1391 (N_1391,N_707,N_367);
or U1392 (N_1392,N_458,N_747);
nor U1393 (N_1393,N_552,N_376);
nand U1394 (N_1394,N_231,N_641);
nor U1395 (N_1395,N_309,N_564);
and U1396 (N_1396,N_183,N_19);
xnor U1397 (N_1397,N_322,N_308);
and U1398 (N_1398,N_432,N_101);
xnor U1399 (N_1399,N_682,N_467);
and U1400 (N_1400,N_544,N_435);
nor U1401 (N_1401,N_329,N_266);
and U1402 (N_1402,N_242,N_649);
and U1403 (N_1403,N_41,N_332);
xnor U1404 (N_1404,N_430,N_360);
or U1405 (N_1405,N_745,N_615);
nor U1406 (N_1406,N_400,N_490);
nor U1407 (N_1407,N_656,N_578);
and U1408 (N_1408,N_464,N_634);
and U1409 (N_1409,N_636,N_100);
and U1410 (N_1410,N_379,N_112);
and U1411 (N_1411,N_647,N_322);
or U1412 (N_1412,N_607,N_731);
nand U1413 (N_1413,N_141,N_139);
nor U1414 (N_1414,N_137,N_304);
xnor U1415 (N_1415,N_201,N_218);
nor U1416 (N_1416,N_719,N_635);
nand U1417 (N_1417,N_566,N_5);
and U1418 (N_1418,N_151,N_669);
xnor U1419 (N_1419,N_237,N_542);
xnor U1420 (N_1420,N_544,N_135);
nor U1421 (N_1421,N_679,N_725);
nand U1422 (N_1422,N_448,N_736);
and U1423 (N_1423,N_100,N_363);
nand U1424 (N_1424,N_695,N_28);
nor U1425 (N_1425,N_57,N_63);
and U1426 (N_1426,N_458,N_731);
nand U1427 (N_1427,N_170,N_456);
nor U1428 (N_1428,N_411,N_219);
nand U1429 (N_1429,N_692,N_38);
and U1430 (N_1430,N_635,N_31);
nor U1431 (N_1431,N_14,N_701);
xor U1432 (N_1432,N_540,N_164);
nor U1433 (N_1433,N_685,N_657);
xnor U1434 (N_1434,N_546,N_674);
nor U1435 (N_1435,N_73,N_176);
nand U1436 (N_1436,N_270,N_457);
nand U1437 (N_1437,N_105,N_8);
xnor U1438 (N_1438,N_43,N_563);
nor U1439 (N_1439,N_62,N_385);
nand U1440 (N_1440,N_83,N_297);
and U1441 (N_1441,N_604,N_543);
and U1442 (N_1442,N_36,N_388);
and U1443 (N_1443,N_422,N_374);
nand U1444 (N_1444,N_210,N_336);
xnor U1445 (N_1445,N_526,N_402);
nor U1446 (N_1446,N_277,N_72);
and U1447 (N_1447,N_508,N_138);
xnor U1448 (N_1448,N_323,N_193);
or U1449 (N_1449,N_648,N_208);
or U1450 (N_1450,N_274,N_347);
xnor U1451 (N_1451,N_729,N_593);
nor U1452 (N_1452,N_268,N_166);
nor U1453 (N_1453,N_212,N_50);
xnor U1454 (N_1454,N_499,N_85);
nor U1455 (N_1455,N_231,N_101);
nor U1456 (N_1456,N_471,N_285);
and U1457 (N_1457,N_266,N_403);
nand U1458 (N_1458,N_16,N_682);
xor U1459 (N_1459,N_239,N_737);
nor U1460 (N_1460,N_1,N_594);
nand U1461 (N_1461,N_669,N_643);
nand U1462 (N_1462,N_421,N_212);
xnor U1463 (N_1463,N_232,N_683);
nor U1464 (N_1464,N_167,N_444);
nand U1465 (N_1465,N_282,N_516);
and U1466 (N_1466,N_561,N_183);
or U1467 (N_1467,N_435,N_122);
nor U1468 (N_1468,N_649,N_34);
and U1469 (N_1469,N_15,N_619);
and U1470 (N_1470,N_105,N_555);
nand U1471 (N_1471,N_465,N_495);
nand U1472 (N_1472,N_432,N_412);
nand U1473 (N_1473,N_666,N_269);
nand U1474 (N_1474,N_516,N_479);
and U1475 (N_1475,N_143,N_583);
and U1476 (N_1476,N_113,N_186);
or U1477 (N_1477,N_18,N_214);
nor U1478 (N_1478,N_447,N_463);
xor U1479 (N_1479,N_569,N_701);
nor U1480 (N_1480,N_3,N_470);
nand U1481 (N_1481,N_391,N_184);
or U1482 (N_1482,N_33,N_735);
xnor U1483 (N_1483,N_114,N_352);
nand U1484 (N_1484,N_554,N_30);
xnor U1485 (N_1485,N_666,N_446);
nand U1486 (N_1486,N_695,N_328);
xor U1487 (N_1487,N_620,N_164);
and U1488 (N_1488,N_45,N_202);
nor U1489 (N_1489,N_507,N_50);
xor U1490 (N_1490,N_125,N_415);
nand U1491 (N_1491,N_616,N_23);
or U1492 (N_1492,N_410,N_235);
and U1493 (N_1493,N_370,N_632);
nor U1494 (N_1494,N_317,N_315);
nand U1495 (N_1495,N_588,N_305);
nor U1496 (N_1496,N_427,N_370);
nand U1497 (N_1497,N_4,N_623);
nand U1498 (N_1498,N_354,N_96);
nor U1499 (N_1499,N_195,N_700);
xor U1500 (N_1500,N_1270,N_880);
nor U1501 (N_1501,N_1352,N_831);
or U1502 (N_1502,N_1374,N_1087);
nand U1503 (N_1503,N_1021,N_1291);
xor U1504 (N_1504,N_1071,N_861);
or U1505 (N_1505,N_890,N_1310);
and U1506 (N_1506,N_1471,N_1223);
nor U1507 (N_1507,N_827,N_878);
nor U1508 (N_1508,N_1314,N_998);
nand U1509 (N_1509,N_1331,N_1033);
nor U1510 (N_1510,N_1007,N_1118);
xnor U1511 (N_1511,N_982,N_1212);
or U1512 (N_1512,N_1416,N_965);
and U1513 (N_1513,N_1181,N_884);
nand U1514 (N_1514,N_1442,N_960);
and U1515 (N_1515,N_1487,N_1348);
nand U1516 (N_1516,N_825,N_1450);
nand U1517 (N_1517,N_1174,N_1128);
and U1518 (N_1518,N_1182,N_828);
nand U1519 (N_1519,N_1138,N_1232);
and U1520 (N_1520,N_1214,N_1124);
nor U1521 (N_1521,N_1447,N_1378);
nor U1522 (N_1522,N_986,N_1261);
nand U1523 (N_1523,N_868,N_1465);
nor U1524 (N_1524,N_1405,N_1122);
or U1525 (N_1525,N_783,N_894);
nor U1526 (N_1526,N_1220,N_967);
nand U1527 (N_1527,N_1211,N_830);
nand U1528 (N_1528,N_1404,N_1161);
and U1529 (N_1529,N_871,N_1157);
xor U1530 (N_1530,N_1362,N_1417);
and U1531 (N_1531,N_1130,N_835);
and U1532 (N_1532,N_882,N_1105);
xnor U1533 (N_1533,N_762,N_1386);
and U1534 (N_1534,N_1113,N_1280);
xor U1535 (N_1535,N_1200,N_1461);
xnor U1536 (N_1536,N_1025,N_1454);
and U1537 (N_1537,N_1491,N_1483);
nand U1538 (N_1538,N_1463,N_834);
and U1539 (N_1539,N_1170,N_1457);
and U1540 (N_1540,N_1060,N_909);
nor U1541 (N_1541,N_1150,N_1394);
and U1542 (N_1542,N_1375,N_1363);
nand U1543 (N_1543,N_901,N_1083);
nand U1544 (N_1544,N_812,N_942);
nand U1545 (N_1545,N_1089,N_771);
and U1546 (N_1546,N_885,N_1193);
nand U1547 (N_1547,N_1354,N_1458);
and U1548 (N_1548,N_1215,N_1349);
xor U1549 (N_1549,N_1149,N_794);
or U1550 (N_1550,N_1322,N_1210);
nor U1551 (N_1551,N_1476,N_972);
or U1552 (N_1552,N_898,N_1344);
or U1553 (N_1553,N_1142,N_1330);
nand U1554 (N_1554,N_1289,N_1018);
or U1555 (N_1555,N_1302,N_1222);
or U1556 (N_1556,N_1068,N_1075);
or U1557 (N_1557,N_1045,N_1109);
or U1558 (N_1558,N_1057,N_1047);
nor U1559 (N_1559,N_1077,N_1178);
or U1560 (N_1560,N_1058,N_968);
xnor U1561 (N_1561,N_1350,N_849);
or U1562 (N_1562,N_1472,N_1159);
and U1563 (N_1563,N_1162,N_1345);
nand U1564 (N_1564,N_1301,N_946);
xor U1565 (N_1565,N_1316,N_1441);
xnor U1566 (N_1566,N_799,N_1426);
and U1567 (N_1567,N_1470,N_1423);
nand U1568 (N_1568,N_1088,N_852);
and U1569 (N_1569,N_1144,N_977);
xor U1570 (N_1570,N_1251,N_1041);
nor U1571 (N_1571,N_1327,N_931);
nand U1572 (N_1572,N_1154,N_1246);
nand U1573 (N_1573,N_949,N_1117);
xnor U1574 (N_1574,N_999,N_786);
nand U1575 (N_1575,N_1437,N_805);
or U1576 (N_1576,N_1422,N_1034);
or U1577 (N_1577,N_1104,N_1067);
nor U1578 (N_1578,N_1095,N_1413);
xor U1579 (N_1579,N_1420,N_761);
and U1580 (N_1580,N_774,N_932);
or U1581 (N_1581,N_1133,N_1321);
nor U1582 (N_1582,N_975,N_873);
nand U1583 (N_1583,N_1368,N_906);
nor U1584 (N_1584,N_1244,N_800);
and U1585 (N_1585,N_869,N_1462);
nor U1586 (N_1586,N_821,N_897);
and U1587 (N_1587,N_1421,N_976);
nor U1588 (N_1588,N_1481,N_1286);
nand U1589 (N_1589,N_987,N_1184);
or U1590 (N_1590,N_1172,N_922);
xor U1591 (N_1591,N_1010,N_1397);
or U1592 (N_1592,N_940,N_1234);
nor U1593 (N_1593,N_1097,N_838);
and U1594 (N_1594,N_1230,N_781);
nand U1595 (N_1595,N_1414,N_1311);
and U1596 (N_1596,N_1282,N_1433);
nor U1597 (N_1597,N_1427,N_1380);
nand U1598 (N_1598,N_1005,N_1435);
nand U1599 (N_1599,N_864,N_1474);
and U1600 (N_1600,N_1262,N_1229);
xor U1601 (N_1601,N_1176,N_1365);
and U1602 (N_1602,N_1451,N_1361);
and U1603 (N_1603,N_757,N_1046);
xnor U1604 (N_1604,N_796,N_1179);
and U1605 (N_1605,N_903,N_853);
xor U1606 (N_1606,N_1020,N_1241);
nor U1607 (N_1607,N_1489,N_951);
and U1608 (N_1608,N_1001,N_1279);
nor U1609 (N_1609,N_914,N_916);
xnor U1610 (N_1610,N_1078,N_939);
xnor U1611 (N_1611,N_839,N_814);
nor U1612 (N_1612,N_1392,N_921);
nor U1613 (N_1613,N_1439,N_1052);
nor U1614 (N_1614,N_1120,N_1115);
and U1615 (N_1615,N_981,N_883);
or U1616 (N_1616,N_845,N_979);
nand U1617 (N_1617,N_778,N_983);
xor U1618 (N_1618,N_1479,N_764);
nor U1619 (N_1619,N_801,N_1191);
nor U1620 (N_1620,N_1111,N_1475);
xor U1621 (N_1621,N_911,N_1165);
or U1622 (N_1622,N_1247,N_1141);
and U1623 (N_1623,N_1208,N_1236);
nand U1624 (N_1624,N_1499,N_959);
nand U1625 (N_1625,N_855,N_1090);
xnor U1626 (N_1626,N_1248,N_1391);
or U1627 (N_1627,N_854,N_1225);
nand U1628 (N_1628,N_1091,N_1164);
or U1629 (N_1629,N_1203,N_1094);
or U1630 (N_1630,N_1081,N_1228);
nor U1631 (N_1631,N_813,N_1055);
nand U1632 (N_1632,N_1395,N_1218);
nor U1633 (N_1633,N_1026,N_1367);
nand U1634 (N_1634,N_1424,N_1412);
nor U1635 (N_1635,N_1002,N_1024);
or U1636 (N_1636,N_1073,N_1132);
xnor U1637 (N_1637,N_877,N_1408);
nand U1638 (N_1638,N_888,N_963);
or U1639 (N_1639,N_973,N_941);
xnor U1640 (N_1640,N_978,N_810);
nand U1641 (N_1641,N_820,N_1080);
nor U1642 (N_1642,N_1456,N_1035);
nand U1643 (N_1643,N_1264,N_867);
nand U1644 (N_1644,N_777,N_1177);
nor U1645 (N_1645,N_770,N_950);
nand U1646 (N_1646,N_957,N_1309);
nor U1647 (N_1647,N_900,N_1379);
or U1648 (N_1648,N_1351,N_1151);
nor U1649 (N_1649,N_1432,N_1296);
nand U1650 (N_1650,N_847,N_1155);
nor U1651 (N_1651,N_1146,N_1290);
xor U1652 (N_1652,N_784,N_776);
and U1653 (N_1653,N_1359,N_912);
nand U1654 (N_1654,N_974,N_1064);
and U1655 (N_1655,N_944,N_1429);
or U1656 (N_1656,N_804,N_1213);
xor U1657 (N_1657,N_1342,N_823);
or U1658 (N_1658,N_1103,N_948);
xnor U1659 (N_1659,N_1242,N_809);
and U1660 (N_1660,N_829,N_1259);
nand U1661 (N_1661,N_1431,N_874);
or U1662 (N_1662,N_1082,N_1326);
xor U1663 (N_1663,N_1096,N_1198);
xor U1664 (N_1664,N_840,N_1468);
nand U1665 (N_1665,N_1283,N_819);
nand U1666 (N_1666,N_1168,N_1364);
xor U1667 (N_1667,N_970,N_893);
xor U1668 (N_1668,N_1147,N_848);
or U1669 (N_1669,N_1267,N_1340);
and U1670 (N_1670,N_991,N_1235);
xor U1671 (N_1671,N_1255,N_907);
or U1672 (N_1672,N_896,N_1346);
or U1673 (N_1673,N_1304,N_943);
and U1674 (N_1674,N_889,N_1336);
nand U1675 (N_1675,N_1143,N_775);
or U1676 (N_1676,N_1153,N_1139);
or U1677 (N_1677,N_1086,N_1305);
and U1678 (N_1678,N_995,N_1003);
and U1679 (N_1679,N_961,N_844);
and U1680 (N_1680,N_899,N_857);
and U1681 (N_1681,N_1163,N_971);
nand U1682 (N_1682,N_1389,N_1185);
nand U1683 (N_1683,N_887,N_1418);
and U1684 (N_1684,N_858,N_841);
nand U1685 (N_1685,N_1328,N_1313);
and U1686 (N_1686,N_779,N_1042);
nand U1687 (N_1687,N_1206,N_1455);
nor U1688 (N_1688,N_808,N_1353);
nand U1689 (N_1689,N_876,N_923);
and U1690 (N_1690,N_1308,N_1406);
and U1691 (N_1691,N_1129,N_1148);
xnor U1692 (N_1692,N_792,N_1099);
and U1693 (N_1693,N_1272,N_765);
nor U1694 (N_1694,N_1050,N_1123);
nor U1695 (N_1695,N_863,N_1016);
nand U1696 (N_1696,N_1383,N_1183);
and U1697 (N_1697,N_1278,N_1469);
and U1698 (N_1698,N_1108,N_1004);
or U1699 (N_1699,N_1085,N_1171);
xnor U1700 (N_1700,N_1051,N_1287);
nand U1701 (N_1701,N_836,N_1201);
xor U1702 (N_1702,N_1195,N_1127);
nand U1703 (N_1703,N_935,N_1023);
and U1704 (N_1704,N_994,N_1102);
nor U1705 (N_1705,N_958,N_795);
and U1706 (N_1706,N_1271,N_1258);
and U1707 (N_1707,N_879,N_1188);
nand U1708 (N_1708,N_1011,N_1219);
xnor U1709 (N_1709,N_1022,N_1482);
nor U1710 (N_1710,N_1371,N_1428);
nor U1711 (N_1711,N_1445,N_750);
nor U1712 (N_1712,N_1131,N_803);
or U1713 (N_1713,N_811,N_773);
nor U1714 (N_1714,N_1173,N_1485);
xor U1715 (N_1715,N_856,N_1459);
and U1716 (N_1716,N_1300,N_1297);
and U1717 (N_1717,N_1460,N_752);
nor U1718 (N_1718,N_1125,N_798);
xnor U1719 (N_1719,N_1032,N_988);
xnor U1720 (N_1720,N_1093,N_1156);
xnor U1721 (N_1721,N_769,N_1260);
and U1722 (N_1722,N_1399,N_891);
nor U1723 (N_1723,N_1373,N_1061);
xor U1724 (N_1724,N_1409,N_1288);
and U1725 (N_1725,N_1369,N_850);
xor U1726 (N_1726,N_1382,N_1398);
or U1727 (N_1727,N_1062,N_1112);
and U1728 (N_1728,N_1044,N_993);
xnor U1729 (N_1729,N_1338,N_859);
nor U1730 (N_1730,N_1252,N_833);
xor U1731 (N_1731,N_1495,N_1190);
nor U1732 (N_1732,N_791,N_1434);
xnor U1733 (N_1733,N_1038,N_1204);
or U1734 (N_1734,N_1037,N_1245);
nor U1735 (N_1735,N_1084,N_1407);
and U1736 (N_1736,N_1430,N_1175);
or U1737 (N_1737,N_1325,N_789);
nand U1738 (N_1738,N_851,N_1292);
nand U1739 (N_1739,N_843,N_1226);
or U1740 (N_1740,N_1333,N_996);
and U1741 (N_1741,N_1145,N_1039);
or U1742 (N_1742,N_1306,N_1192);
xor U1743 (N_1743,N_1334,N_1317);
xnor U1744 (N_1744,N_1347,N_1400);
nor U1745 (N_1745,N_1000,N_1323);
nor U1746 (N_1746,N_1028,N_1199);
or U1747 (N_1747,N_1269,N_1043);
and U1748 (N_1748,N_1009,N_1186);
xnor U1749 (N_1749,N_815,N_1339);
nand U1750 (N_1750,N_1356,N_758);
xor U1751 (N_1751,N_925,N_927);
xnor U1752 (N_1752,N_766,N_1227);
or U1753 (N_1753,N_895,N_1017);
and U1754 (N_1754,N_832,N_1238);
xnor U1755 (N_1755,N_1372,N_1197);
and U1756 (N_1756,N_930,N_937);
nand U1757 (N_1757,N_1014,N_772);
nor U1758 (N_1758,N_1180,N_1167);
or U1759 (N_1759,N_1040,N_1209);
nand U1760 (N_1760,N_1393,N_1320);
or U1761 (N_1761,N_1008,N_1303);
nand U1762 (N_1762,N_1135,N_929);
or U1763 (N_1763,N_908,N_1049);
and U1764 (N_1764,N_1275,N_790);
or U1765 (N_1765,N_1137,N_862);
and U1766 (N_1766,N_997,N_1263);
nor U1767 (N_1767,N_1256,N_1063);
nand U1768 (N_1768,N_1335,N_1384);
nor U1769 (N_1769,N_837,N_1307);
nor U1770 (N_1770,N_1467,N_1250);
xnor U1771 (N_1771,N_1376,N_1464);
nand U1772 (N_1772,N_952,N_1152);
or U1773 (N_1773,N_1066,N_1295);
nand U1774 (N_1774,N_1285,N_754);
and U1775 (N_1775,N_902,N_1187);
or U1776 (N_1776,N_1189,N_1121);
nand U1777 (N_1777,N_989,N_1031);
nand U1778 (N_1778,N_926,N_1140);
nand U1779 (N_1779,N_818,N_865);
xnor U1780 (N_1780,N_938,N_1484);
nor U1781 (N_1781,N_870,N_1449);
nand U1782 (N_1782,N_817,N_962);
xor U1783 (N_1783,N_910,N_788);
or U1784 (N_1784,N_1134,N_787);
nor U1785 (N_1785,N_1415,N_1355);
or U1786 (N_1786,N_1013,N_1443);
nor U1787 (N_1787,N_956,N_1106);
nor U1788 (N_1788,N_866,N_1056);
nand U1789 (N_1789,N_1169,N_782);
and U1790 (N_1790,N_802,N_1160);
and U1791 (N_1791,N_1217,N_1494);
nand U1792 (N_1792,N_1281,N_1315);
or U1793 (N_1793,N_1438,N_1284);
and U1794 (N_1794,N_767,N_1254);
or U1795 (N_1795,N_1194,N_1401);
and U1796 (N_1796,N_1268,N_954);
or U1797 (N_1797,N_822,N_1015);
or U1798 (N_1798,N_1233,N_1480);
nand U1799 (N_1799,N_990,N_1419);
nor U1800 (N_1800,N_1496,N_933);
nor U1801 (N_1801,N_760,N_985);
and U1802 (N_1802,N_905,N_1403);
xnor U1803 (N_1803,N_1243,N_1337);
or U1804 (N_1804,N_1332,N_1059);
nand U1805 (N_1805,N_1012,N_1265);
nand U1806 (N_1806,N_955,N_1231);
nand U1807 (N_1807,N_1054,N_1473);
nand U1808 (N_1808,N_1490,N_1107);
or U1809 (N_1809,N_1266,N_915);
xor U1810 (N_1810,N_1274,N_1019);
and U1811 (N_1811,N_1253,N_1497);
nor U1812 (N_1812,N_768,N_1377);
and U1813 (N_1813,N_920,N_969);
xnor U1814 (N_1814,N_1410,N_1119);
or U1815 (N_1815,N_1100,N_807);
nand U1816 (N_1816,N_1101,N_1411);
or U1817 (N_1817,N_924,N_1249);
nand U1818 (N_1818,N_1452,N_953);
or U1819 (N_1819,N_1070,N_966);
or U1820 (N_1820,N_1358,N_1486);
and U1821 (N_1821,N_756,N_1453);
or U1822 (N_1822,N_1076,N_1224);
nor U1823 (N_1823,N_846,N_1216);
or U1824 (N_1824,N_881,N_945);
and U1825 (N_1825,N_1273,N_1136);
nor U1826 (N_1826,N_886,N_806);
xnor U1827 (N_1827,N_1488,N_1360);
nand U1828 (N_1828,N_1477,N_913);
and U1829 (N_1829,N_1402,N_1116);
xnor U1830 (N_1830,N_1074,N_1072);
nor U1831 (N_1831,N_826,N_1048);
xor U1832 (N_1832,N_1030,N_1202);
nor U1833 (N_1833,N_1440,N_793);
or U1834 (N_1834,N_984,N_1396);
nand U1835 (N_1835,N_875,N_860);
or U1836 (N_1836,N_1257,N_1357);
or U1837 (N_1837,N_1385,N_1079);
and U1838 (N_1838,N_980,N_1341);
or U1839 (N_1839,N_1381,N_1370);
and U1840 (N_1840,N_917,N_785);
nor U1841 (N_1841,N_1294,N_1065);
nand U1842 (N_1842,N_1390,N_1318);
nand U1843 (N_1843,N_1237,N_1098);
nor U1844 (N_1844,N_1069,N_1126);
nor U1845 (N_1845,N_1293,N_1027);
nor U1846 (N_1846,N_1366,N_919);
xor U1847 (N_1847,N_872,N_1446);
xnor U1848 (N_1848,N_1444,N_1425);
xnor U1849 (N_1849,N_1036,N_1319);
nor U1850 (N_1850,N_1196,N_904);
nand U1851 (N_1851,N_928,N_759);
or U1852 (N_1852,N_1492,N_751);
or U1853 (N_1853,N_1312,N_1110);
and U1854 (N_1854,N_842,N_753);
or U1855 (N_1855,N_992,N_1299);
xnor U1856 (N_1856,N_1298,N_936);
or U1857 (N_1857,N_1493,N_1436);
and U1858 (N_1858,N_1114,N_1478);
or U1859 (N_1859,N_1029,N_964);
or U1860 (N_1860,N_1277,N_918);
xnor U1861 (N_1861,N_1329,N_1221);
nand U1862 (N_1862,N_947,N_1276);
and U1863 (N_1863,N_797,N_755);
and U1864 (N_1864,N_1006,N_1466);
and U1865 (N_1865,N_1343,N_1053);
or U1866 (N_1866,N_824,N_1092);
nor U1867 (N_1867,N_1205,N_1387);
or U1868 (N_1868,N_816,N_1324);
xnor U1869 (N_1869,N_1158,N_1498);
nor U1870 (N_1870,N_934,N_892);
and U1871 (N_1871,N_1388,N_1240);
or U1872 (N_1872,N_1239,N_763);
and U1873 (N_1873,N_1166,N_780);
nor U1874 (N_1874,N_1448,N_1207);
and U1875 (N_1875,N_991,N_985);
nand U1876 (N_1876,N_970,N_781);
or U1877 (N_1877,N_773,N_1411);
xor U1878 (N_1878,N_788,N_1035);
nand U1879 (N_1879,N_758,N_1411);
and U1880 (N_1880,N_1147,N_1303);
nand U1881 (N_1881,N_950,N_979);
xor U1882 (N_1882,N_822,N_880);
nand U1883 (N_1883,N_1345,N_1074);
nor U1884 (N_1884,N_1220,N_1465);
nor U1885 (N_1885,N_846,N_771);
xnor U1886 (N_1886,N_1170,N_1109);
and U1887 (N_1887,N_1131,N_915);
and U1888 (N_1888,N_947,N_1265);
nand U1889 (N_1889,N_903,N_1493);
and U1890 (N_1890,N_1106,N_1066);
or U1891 (N_1891,N_1284,N_1417);
xnor U1892 (N_1892,N_1189,N_846);
nor U1893 (N_1893,N_1265,N_1307);
nand U1894 (N_1894,N_1188,N_823);
or U1895 (N_1895,N_1458,N_1211);
or U1896 (N_1896,N_1297,N_1184);
or U1897 (N_1897,N_1329,N_910);
nor U1898 (N_1898,N_1318,N_1286);
nor U1899 (N_1899,N_1088,N_1124);
nor U1900 (N_1900,N_1170,N_1233);
xnor U1901 (N_1901,N_834,N_1147);
xor U1902 (N_1902,N_1280,N_1017);
or U1903 (N_1903,N_863,N_1496);
nor U1904 (N_1904,N_1412,N_1344);
nor U1905 (N_1905,N_1313,N_773);
nor U1906 (N_1906,N_1190,N_1470);
or U1907 (N_1907,N_855,N_992);
or U1908 (N_1908,N_951,N_1322);
or U1909 (N_1909,N_1101,N_1405);
nor U1910 (N_1910,N_819,N_772);
nand U1911 (N_1911,N_1069,N_947);
nor U1912 (N_1912,N_1180,N_803);
and U1913 (N_1913,N_1166,N_1175);
nand U1914 (N_1914,N_899,N_1322);
nor U1915 (N_1915,N_1095,N_1447);
xor U1916 (N_1916,N_1066,N_1192);
and U1917 (N_1917,N_1127,N_1048);
or U1918 (N_1918,N_998,N_862);
nor U1919 (N_1919,N_1131,N_1112);
or U1920 (N_1920,N_1034,N_826);
and U1921 (N_1921,N_1071,N_1415);
or U1922 (N_1922,N_858,N_1461);
nor U1923 (N_1923,N_1027,N_1436);
nor U1924 (N_1924,N_1432,N_1406);
and U1925 (N_1925,N_1243,N_934);
nand U1926 (N_1926,N_1067,N_1256);
nor U1927 (N_1927,N_1379,N_994);
and U1928 (N_1928,N_1120,N_1384);
xnor U1929 (N_1929,N_1319,N_943);
nand U1930 (N_1930,N_811,N_1141);
or U1931 (N_1931,N_1475,N_1412);
or U1932 (N_1932,N_1371,N_1101);
xor U1933 (N_1933,N_1097,N_1378);
nand U1934 (N_1934,N_1243,N_1461);
and U1935 (N_1935,N_906,N_940);
nand U1936 (N_1936,N_916,N_1397);
nor U1937 (N_1937,N_1039,N_1131);
xor U1938 (N_1938,N_1132,N_1017);
or U1939 (N_1939,N_956,N_1451);
xnor U1940 (N_1940,N_1400,N_918);
or U1941 (N_1941,N_1273,N_1222);
nand U1942 (N_1942,N_990,N_993);
nor U1943 (N_1943,N_854,N_830);
or U1944 (N_1944,N_1196,N_950);
nor U1945 (N_1945,N_1286,N_1220);
or U1946 (N_1946,N_1041,N_1334);
nor U1947 (N_1947,N_1444,N_1253);
or U1948 (N_1948,N_765,N_800);
and U1949 (N_1949,N_888,N_1332);
and U1950 (N_1950,N_1306,N_1257);
nand U1951 (N_1951,N_963,N_1237);
nand U1952 (N_1952,N_933,N_1171);
and U1953 (N_1953,N_1413,N_1398);
nand U1954 (N_1954,N_1157,N_1245);
and U1955 (N_1955,N_1068,N_1053);
nand U1956 (N_1956,N_1270,N_913);
and U1957 (N_1957,N_1214,N_914);
nand U1958 (N_1958,N_986,N_1455);
nor U1959 (N_1959,N_842,N_1028);
nand U1960 (N_1960,N_1455,N_1449);
nor U1961 (N_1961,N_913,N_752);
nor U1962 (N_1962,N_942,N_1142);
and U1963 (N_1963,N_1081,N_1019);
nor U1964 (N_1964,N_1239,N_1214);
or U1965 (N_1965,N_856,N_1151);
xor U1966 (N_1966,N_821,N_1473);
and U1967 (N_1967,N_857,N_810);
nand U1968 (N_1968,N_839,N_1228);
or U1969 (N_1969,N_783,N_991);
or U1970 (N_1970,N_995,N_1273);
or U1971 (N_1971,N_1353,N_1124);
nor U1972 (N_1972,N_849,N_1422);
and U1973 (N_1973,N_1421,N_1374);
or U1974 (N_1974,N_1314,N_1044);
and U1975 (N_1975,N_848,N_851);
nor U1976 (N_1976,N_824,N_1098);
nand U1977 (N_1977,N_1282,N_1204);
nand U1978 (N_1978,N_1143,N_1481);
nor U1979 (N_1979,N_1007,N_1264);
nor U1980 (N_1980,N_1410,N_894);
xor U1981 (N_1981,N_1440,N_754);
nor U1982 (N_1982,N_1029,N_1449);
nor U1983 (N_1983,N_1377,N_839);
nand U1984 (N_1984,N_861,N_1115);
or U1985 (N_1985,N_923,N_1184);
or U1986 (N_1986,N_1291,N_1270);
and U1987 (N_1987,N_1294,N_1345);
xnor U1988 (N_1988,N_1440,N_1443);
xnor U1989 (N_1989,N_1314,N_1345);
nand U1990 (N_1990,N_910,N_933);
nand U1991 (N_1991,N_1216,N_835);
nor U1992 (N_1992,N_1001,N_855);
nand U1993 (N_1993,N_1394,N_839);
nand U1994 (N_1994,N_1434,N_1451);
and U1995 (N_1995,N_1420,N_1147);
nor U1996 (N_1996,N_1169,N_990);
nand U1997 (N_1997,N_834,N_1239);
and U1998 (N_1998,N_1412,N_1338);
xnor U1999 (N_1999,N_1438,N_1434);
nand U2000 (N_2000,N_1043,N_1166);
or U2001 (N_2001,N_1168,N_1209);
or U2002 (N_2002,N_1473,N_1170);
xnor U2003 (N_2003,N_1223,N_1008);
xor U2004 (N_2004,N_1189,N_795);
nand U2005 (N_2005,N_1124,N_1387);
nor U2006 (N_2006,N_1174,N_1352);
and U2007 (N_2007,N_1036,N_1488);
nor U2008 (N_2008,N_1239,N_1310);
nor U2009 (N_2009,N_1005,N_1371);
nor U2010 (N_2010,N_1248,N_1349);
nor U2011 (N_2011,N_922,N_1065);
or U2012 (N_2012,N_764,N_815);
nor U2013 (N_2013,N_803,N_1409);
nor U2014 (N_2014,N_1355,N_1460);
or U2015 (N_2015,N_1435,N_922);
or U2016 (N_2016,N_1291,N_856);
xnor U2017 (N_2017,N_857,N_1280);
xnor U2018 (N_2018,N_1362,N_776);
xnor U2019 (N_2019,N_934,N_1019);
nor U2020 (N_2020,N_859,N_1118);
nand U2021 (N_2021,N_1382,N_1351);
nor U2022 (N_2022,N_1131,N_1225);
nand U2023 (N_2023,N_1127,N_1371);
xor U2024 (N_2024,N_943,N_1429);
xnor U2025 (N_2025,N_1311,N_1267);
or U2026 (N_2026,N_1450,N_1337);
nor U2027 (N_2027,N_1457,N_1200);
or U2028 (N_2028,N_1158,N_1283);
or U2029 (N_2029,N_897,N_1455);
or U2030 (N_2030,N_1113,N_1082);
or U2031 (N_2031,N_1240,N_1195);
or U2032 (N_2032,N_1298,N_895);
or U2033 (N_2033,N_981,N_1319);
nand U2034 (N_2034,N_903,N_925);
or U2035 (N_2035,N_1495,N_860);
xor U2036 (N_2036,N_761,N_1415);
and U2037 (N_2037,N_1360,N_1448);
nor U2038 (N_2038,N_920,N_843);
xor U2039 (N_2039,N_1333,N_836);
xor U2040 (N_2040,N_789,N_785);
or U2041 (N_2041,N_984,N_1437);
nor U2042 (N_2042,N_1456,N_1237);
xor U2043 (N_2043,N_881,N_1454);
nor U2044 (N_2044,N_936,N_1485);
nand U2045 (N_2045,N_870,N_965);
nor U2046 (N_2046,N_1290,N_1015);
xnor U2047 (N_2047,N_1380,N_1107);
and U2048 (N_2048,N_851,N_1217);
and U2049 (N_2049,N_934,N_1480);
nand U2050 (N_2050,N_1043,N_1000);
or U2051 (N_2051,N_1193,N_1032);
xor U2052 (N_2052,N_971,N_1338);
xnor U2053 (N_2053,N_1190,N_780);
nor U2054 (N_2054,N_905,N_931);
xnor U2055 (N_2055,N_1032,N_1177);
nand U2056 (N_2056,N_798,N_1212);
nor U2057 (N_2057,N_1106,N_889);
or U2058 (N_2058,N_759,N_1296);
and U2059 (N_2059,N_1009,N_1385);
and U2060 (N_2060,N_951,N_803);
xor U2061 (N_2061,N_771,N_1072);
xnor U2062 (N_2062,N_912,N_1310);
or U2063 (N_2063,N_906,N_1158);
and U2064 (N_2064,N_1303,N_1062);
nand U2065 (N_2065,N_1119,N_1088);
or U2066 (N_2066,N_1266,N_883);
or U2067 (N_2067,N_1302,N_932);
or U2068 (N_2068,N_1120,N_790);
xor U2069 (N_2069,N_901,N_946);
and U2070 (N_2070,N_792,N_819);
xor U2071 (N_2071,N_760,N_1486);
or U2072 (N_2072,N_1414,N_1364);
and U2073 (N_2073,N_1392,N_1190);
and U2074 (N_2074,N_977,N_1437);
and U2075 (N_2075,N_1260,N_1044);
or U2076 (N_2076,N_1455,N_827);
nand U2077 (N_2077,N_805,N_1049);
xor U2078 (N_2078,N_1338,N_922);
nand U2079 (N_2079,N_1430,N_841);
and U2080 (N_2080,N_811,N_1284);
and U2081 (N_2081,N_869,N_1260);
xnor U2082 (N_2082,N_1322,N_1243);
and U2083 (N_2083,N_1208,N_1375);
nand U2084 (N_2084,N_1356,N_1349);
nor U2085 (N_2085,N_906,N_1060);
nor U2086 (N_2086,N_997,N_1042);
or U2087 (N_2087,N_1094,N_1052);
nor U2088 (N_2088,N_1213,N_1029);
xnor U2089 (N_2089,N_1265,N_951);
xnor U2090 (N_2090,N_1100,N_1493);
xnor U2091 (N_2091,N_942,N_804);
and U2092 (N_2092,N_1005,N_943);
and U2093 (N_2093,N_1469,N_1119);
nor U2094 (N_2094,N_766,N_849);
xnor U2095 (N_2095,N_803,N_1072);
nor U2096 (N_2096,N_979,N_1389);
nor U2097 (N_2097,N_823,N_1409);
xnor U2098 (N_2098,N_1189,N_1449);
xnor U2099 (N_2099,N_808,N_1000);
xnor U2100 (N_2100,N_894,N_977);
and U2101 (N_2101,N_1052,N_876);
and U2102 (N_2102,N_1233,N_1496);
or U2103 (N_2103,N_758,N_1155);
nand U2104 (N_2104,N_1446,N_788);
nor U2105 (N_2105,N_1184,N_921);
xor U2106 (N_2106,N_969,N_1243);
nor U2107 (N_2107,N_1021,N_863);
and U2108 (N_2108,N_1270,N_1408);
or U2109 (N_2109,N_980,N_997);
and U2110 (N_2110,N_985,N_1184);
and U2111 (N_2111,N_1203,N_909);
and U2112 (N_2112,N_1028,N_797);
xor U2113 (N_2113,N_1385,N_1083);
and U2114 (N_2114,N_1134,N_1280);
and U2115 (N_2115,N_1099,N_1330);
and U2116 (N_2116,N_1106,N_1224);
nor U2117 (N_2117,N_1217,N_1445);
and U2118 (N_2118,N_1019,N_1461);
and U2119 (N_2119,N_1073,N_1357);
nand U2120 (N_2120,N_1401,N_1053);
nand U2121 (N_2121,N_1088,N_1234);
or U2122 (N_2122,N_1132,N_1264);
nand U2123 (N_2123,N_1421,N_1487);
or U2124 (N_2124,N_1409,N_1296);
xnor U2125 (N_2125,N_1474,N_951);
nand U2126 (N_2126,N_875,N_1052);
and U2127 (N_2127,N_1138,N_1282);
nor U2128 (N_2128,N_953,N_1430);
nor U2129 (N_2129,N_998,N_1261);
or U2130 (N_2130,N_763,N_1244);
and U2131 (N_2131,N_766,N_1359);
or U2132 (N_2132,N_1018,N_1168);
nor U2133 (N_2133,N_1261,N_928);
nor U2134 (N_2134,N_1106,N_1450);
and U2135 (N_2135,N_1439,N_1275);
nand U2136 (N_2136,N_1087,N_1008);
and U2137 (N_2137,N_1243,N_767);
nand U2138 (N_2138,N_1219,N_1356);
nand U2139 (N_2139,N_1220,N_1056);
or U2140 (N_2140,N_1018,N_777);
xor U2141 (N_2141,N_1271,N_902);
nor U2142 (N_2142,N_1077,N_1455);
or U2143 (N_2143,N_1272,N_1255);
and U2144 (N_2144,N_1050,N_1166);
or U2145 (N_2145,N_752,N_1411);
nor U2146 (N_2146,N_879,N_1360);
and U2147 (N_2147,N_1470,N_1008);
nor U2148 (N_2148,N_1144,N_1492);
and U2149 (N_2149,N_1000,N_1029);
and U2150 (N_2150,N_1083,N_955);
or U2151 (N_2151,N_935,N_999);
xnor U2152 (N_2152,N_883,N_760);
nor U2153 (N_2153,N_1080,N_978);
nand U2154 (N_2154,N_795,N_983);
and U2155 (N_2155,N_1435,N_1057);
xnor U2156 (N_2156,N_813,N_864);
xor U2157 (N_2157,N_1103,N_828);
or U2158 (N_2158,N_1351,N_1360);
or U2159 (N_2159,N_1191,N_897);
nand U2160 (N_2160,N_1419,N_866);
xnor U2161 (N_2161,N_1197,N_1220);
and U2162 (N_2162,N_1421,N_1424);
nand U2163 (N_2163,N_1121,N_969);
nand U2164 (N_2164,N_818,N_1121);
xnor U2165 (N_2165,N_1233,N_798);
nor U2166 (N_2166,N_1261,N_1157);
nor U2167 (N_2167,N_1052,N_1202);
and U2168 (N_2168,N_869,N_1157);
nor U2169 (N_2169,N_1375,N_937);
or U2170 (N_2170,N_1163,N_1044);
or U2171 (N_2171,N_841,N_1150);
xor U2172 (N_2172,N_1287,N_1296);
and U2173 (N_2173,N_971,N_1351);
or U2174 (N_2174,N_1283,N_917);
nand U2175 (N_2175,N_802,N_1220);
or U2176 (N_2176,N_1484,N_1353);
xnor U2177 (N_2177,N_827,N_1462);
xnor U2178 (N_2178,N_1303,N_1198);
nor U2179 (N_2179,N_1215,N_1158);
nor U2180 (N_2180,N_1331,N_759);
xor U2181 (N_2181,N_1324,N_791);
xor U2182 (N_2182,N_1093,N_1393);
and U2183 (N_2183,N_1027,N_947);
xnor U2184 (N_2184,N_774,N_970);
xnor U2185 (N_2185,N_1154,N_1369);
nor U2186 (N_2186,N_817,N_1358);
xnor U2187 (N_2187,N_825,N_904);
and U2188 (N_2188,N_1230,N_1194);
or U2189 (N_2189,N_856,N_1001);
nor U2190 (N_2190,N_1197,N_1274);
or U2191 (N_2191,N_1166,N_1473);
nor U2192 (N_2192,N_1184,N_758);
nand U2193 (N_2193,N_1196,N_845);
or U2194 (N_2194,N_953,N_1080);
or U2195 (N_2195,N_1240,N_1164);
xor U2196 (N_2196,N_936,N_1157);
nand U2197 (N_2197,N_1121,N_831);
xnor U2198 (N_2198,N_1167,N_1301);
or U2199 (N_2199,N_886,N_1457);
nand U2200 (N_2200,N_1143,N_823);
xor U2201 (N_2201,N_873,N_1103);
nor U2202 (N_2202,N_1252,N_1434);
nand U2203 (N_2203,N_1478,N_875);
nor U2204 (N_2204,N_1393,N_754);
nand U2205 (N_2205,N_1418,N_836);
xnor U2206 (N_2206,N_1480,N_798);
xor U2207 (N_2207,N_1328,N_1188);
nor U2208 (N_2208,N_1274,N_1498);
nor U2209 (N_2209,N_1467,N_1052);
nand U2210 (N_2210,N_1457,N_1494);
xnor U2211 (N_2211,N_1018,N_1486);
or U2212 (N_2212,N_1446,N_1441);
and U2213 (N_2213,N_1439,N_1244);
xnor U2214 (N_2214,N_883,N_1312);
nor U2215 (N_2215,N_1052,N_975);
or U2216 (N_2216,N_1413,N_1290);
or U2217 (N_2217,N_1191,N_1383);
nand U2218 (N_2218,N_784,N_1406);
nand U2219 (N_2219,N_959,N_1019);
nor U2220 (N_2220,N_1152,N_1214);
xnor U2221 (N_2221,N_1405,N_1356);
nand U2222 (N_2222,N_1376,N_908);
nand U2223 (N_2223,N_1464,N_1003);
or U2224 (N_2224,N_1109,N_1039);
xor U2225 (N_2225,N_935,N_994);
nand U2226 (N_2226,N_799,N_926);
nor U2227 (N_2227,N_926,N_1437);
and U2228 (N_2228,N_800,N_1041);
xnor U2229 (N_2229,N_1433,N_1107);
xnor U2230 (N_2230,N_1386,N_1065);
xor U2231 (N_2231,N_1055,N_1304);
xnor U2232 (N_2232,N_821,N_1492);
or U2233 (N_2233,N_942,N_1075);
xnor U2234 (N_2234,N_1084,N_1398);
and U2235 (N_2235,N_851,N_1324);
xor U2236 (N_2236,N_778,N_1126);
xor U2237 (N_2237,N_1167,N_1352);
xnor U2238 (N_2238,N_840,N_1004);
or U2239 (N_2239,N_972,N_1097);
and U2240 (N_2240,N_981,N_1291);
nand U2241 (N_2241,N_784,N_1305);
xor U2242 (N_2242,N_1118,N_1266);
nor U2243 (N_2243,N_897,N_960);
xor U2244 (N_2244,N_1182,N_1389);
nand U2245 (N_2245,N_1123,N_846);
or U2246 (N_2246,N_755,N_1420);
nand U2247 (N_2247,N_1114,N_885);
and U2248 (N_2248,N_822,N_1194);
or U2249 (N_2249,N_843,N_1368);
nand U2250 (N_2250,N_2077,N_2195);
nand U2251 (N_2251,N_1512,N_2170);
xor U2252 (N_2252,N_1572,N_1626);
and U2253 (N_2253,N_1841,N_2097);
xor U2254 (N_2254,N_1828,N_2171);
and U2255 (N_2255,N_1967,N_2124);
and U2256 (N_2256,N_1526,N_1984);
xor U2257 (N_2257,N_2237,N_1994);
or U2258 (N_2258,N_1800,N_2096);
or U2259 (N_2259,N_1642,N_2193);
nor U2260 (N_2260,N_1951,N_1565);
and U2261 (N_2261,N_1613,N_2030);
nor U2262 (N_2262,N_1627,N_1639);
nand U2263 (N_2263,N_1679,N_2115);
or U2264 (N_2264,N_1655,N_1759);
and U2265 (N_2265,N_1935,N_1570);
nand U2266 (N_2266,N_1713,N_2128);
xor U2267 (N_2267,N_1564,N_2024);
xor U2268 (N_2268,N_2015,N_2009);
nor U2269 (N_2269,N_1827,N_2153);
nor U2270 (N_2270,N_1976,N_1578);
and U2271 (N_2271,N_2241,N_1813);
xnor U2272 (N_2272,N_2040,N_2181);
and U2273 (N_2273,N_1647,N_1753);
and U2274 (N_2274,N_1840,N_1523);
and U2275 (N_2275,N_1518,N_2150);
and U2276 (N_2276,N_2178,N_1847);
and U2277 (N_2277,N_1592,N_1785);
and U2278 (N_2278,N_1911,N_1640);
xnor U2279 (N_2279,N_2071,N_2199);
nand U2280 (N_2280,N_2005,N_2172);
xnor U2281 (N_2281,N_2225,N_1772);
or U2282 (N_2282,N_1693,N_2032);
and U2283 (N_2283,N_1632,N_1850);
nor U2284 (N_2284,N_2160,N_1543);
xor U2285 (N_2285,N_2017,N_1694);
nand U2286 (N_2286,N_2034,N_1608);
xor U2287 (N_2287,N_1648,N_1576);
xor U2288 (N_2288,N_1587,N_1882);
or U2289 (N_2289,N_2223,N_1701);
or U2290 (N_2290,N_1584,N_1870);
or U2291 (N_2291,N_1541,N_1652);
xnor U2292 (N_2292,N_2156,N_1844);
or U2293 (N_2293,N_1599,N_1688);
xnor U2294 (N_2294,N_1696,N_1992);
nor U2295 (N_2295,N_1861,N_1862);
and U2296 (N_2296,N_2233,N_1952);
nand U2297 (N_2297,N_2014,N_2122);
or U2298 (N_2298,N_1638,N_1798);
xor U2299 (N_2299,N_1858,N_1932);
nor U2300 (N_2300,N_1818,N_1871);
or U2301 (N_2301,N_1692,N_2143);
xor U2302 (N_2302,N_1734,N_1604);
nor U2303 (N_2303,N_2242,N_1631);
xnor U2304 (N_2304,N_1622,N_1706);
and U2305 (N_2305,N_2104,N_2146);
or U2306 (N_2306,N_1915,N_1566);
nand U2307 (N_2307,N_2101,N_2126);
nor U2308 (N_2308,N_2113,N_1756);
nand U2309 (N_2309,N_1936,N_1943);
and U2310 (N_2310,N_1575,N_1516);
or U2311 (N_2311,N_2068,N_1620);
and U2312 (N_2312,N_1600,N_2121);
and U2313 (N_2313,N_2159,N_2038);
nor U2314 (N_2314,N_2012,N_1560);
or U2315 (N_2315,N_1624,N_1883);
nor U2316 (N_2316,N_1928,N_2207);
and U2317 (N_2317,N_1938,N_1629);
and U2318 (N_2318,N_1905,N_1663);
nor U2319 (N_2319,N_2025,N_1633);
and U2320 (N_2320,N_1845,N_1559);
or U2321 (N_2321,N_1860,N_1670);
or U2322 (N_2322,N_1906,N_1875);
nand U2323 (N_2323,N_1815,N_2063);
or U2324 (N_2324,N_2119,N_2167);
and U2325 (N_2325,N_1553,N_1520);
nand U2326 (N_2326,N_1762,N_2080);
nor U2327 (N_2327,N_2131,N_2190);
nand U2328 (N_2328,N_1719,N_2092);
and U2329 (N_2329,N_1654,N_1881);
nor U2330 (N_2330,N_1986,N_1773);
xnor U2331 (N_2331,N_2175,N_1509);
or U2332 (N_2332,N_1635,N_1894);
and U2333 (N_2333,N_1605,N_2042);
or U2334 (N_2334,N_1649,N_1980);
nor U2335 (N_2335,N_1996,N_1700);
or U2336 (N_2336,N_1767,N_1909);
xnor U2337 (N_2337,N_1950,N_1751);
or U2338 (N_2338,N_1920,N_1784);
nand U2339 (N_2339,N_1904,N_1973);
and U2340 (N_2340,N_1926,N_1825);
nor U2341 (N_2341,N_1889,N_2154);
nor U2342 (N_2342,N_1671,N_2102);
xnor U2343 (N_2343,N_2161,N_1876);
and U2344 (N_2344,N_1832,N_1852);
nand U2345 (N_2345,N_1568,N_1893);
or U2346 (N_2346,N_1855,N_1569);
xor U2347 (N_2347,N_1697,N_2201);
or U2348 (N_2348,N_2236,N_1710);
and U2349 (N_2349,N_1979,N_1801);
and U2350 (N_2350,N_1517,N_1752);
and U2351 (N_2351,N_1704,N_1787);
or U2352 (N_2352,N_1805,N_2185);
or U2353 (N_2353,N_1758,N_1991);
xor U2354 (N_2354,N_1764,N_1792);
or U2355 (N_2355,N_1609,N_1908);
nor U2356 (N_2356,N_1808,N_1879);
xnor U2357 (N_2357,N_1834,N_1830);
nor U2358 (N_2358,N_2016,N_1807);
and U2359 (N_2359,N_1941,N_1867);
nor U2360 (N_2360,N_2238,N_1571);
nor U2361 (N_2361,N_1506,N_2050);
xor U2362 (N_2362,N_2021,N_1746);
xor U2363 (N_2363,N_1975,N_1525);
xor U2364 (N_2364,N_2070,N_1775);
and U2365 (N_2365,N_2189,N_1720);
and U2366 (N_2366,N_1816,N_1750);
or U2367 (N_2367,N_1786,N_2197);
nand U2368 (N_2368,N_2202,N_1736);
nand U2369 (N_2369,N_2106,N_1680);
or U2370 (N_2370,N_1757,N_2123);
xnor U2371 (N_2371,N_1795,N_2148);
and U2372 (N_2372,N_2033,N_2100);
or U2373 (N_2373,N_2191,N_2120);
xnor U2374 (N_2374,N_1983,N_2053);
and U2375 (N_2375,N_1567,N_2039);
xor U2376 (N_2376,N_1903,N_1511);
or U2377 (N_2377,N_2088,N_1755);
nor U2378 (N_2378,N_1799,N_1831);
and U2379 (N_2379,N_1645,N_2125);
nor U2380 (N_2380,N_2176,N_1958);
and U2381 (N_2381,N_2114,N_1957);
nand U2382 (N_2382,N_1942,N_1666);
nand U2383 (N_2383,N_2147,N_1948);
and U2384 (N_2384,N_1944,N_1745);
nand U2385 (N_2385,N_1698,N_1997);
nor U2386 (N_2386,N_1930,N_1820);
nor U2387 (N_2387,N_1641,N_2108);
nor U2388 (N_2388,N_2116,N_2142);
nand U2389 (N_2389,N_1536,N_1835);
xor U2390 (N_2390,N_1874,N_2151);
nor U2391 (N_2391,N_2169,N_2222);
or U2392 (N_2392,N_2111,N_1732);
nor U2393 (N_2393,N_1502,N_1548);
or U2394 (N_2394,N_2246,N_2245);
and U2395 (N_2395,N_1657,N_1669);
nor U2396 (N_2396,N_2078,N_1527);
xor U2397 (N_2397,N_1849,N_2180);
nand U2398 (N_2398,N_2132,N_1708);
xor U2399 (N_2399,N_1999,N_2234);
nand U2400 (N_2400,N_1658,N_1607);
nor U2401 (N_2401,N_1829,N_2130);
and U2402 (N_2402,N_1782,N_1561);
nand U2403 (N_2403,N_1718,N_2065);
or U2404 (N_2404,N_1691,N_1937);
or U2405 (N_2405,N_1922,N_1885);
xnor U2406 (N_2406,N_1797,N_2211);
nand U2407 (N_2407,N_1978,N_2019);
nand U2408 (N_2408,N_1896,N_1966);
and U2409 (N_2409,N_2057,N_2001);
nand U2410 (N_2410,N_1778,N_2184);
nand U2411 (N_2411,N_1848,N_1927);
nand U2412 (N_2412,N_2164,N_2141);
or U2413 (N_2413,N_1577,N_1637);
or U2414 (N_2414,N_1838,N_1779);
and U2415 (N_2415,N_1636,N_2004);
and U2416 (N_2416,N_1743,N_1674);
nand U2417 (N_2417,N_1596,N_1695);
nor U2418 (N_2418,N_1611,N_1895);
xnor U2419 (N_2419,N_1595,N_1741);
nor U2420 (N_2420,N_1659,N_2018);
nor U2421 (N_2421,N_1890,N_1985);
or U2422 (N_2422,N_2129,N_2035);
nand U2423 (N_2423,N_1551,N_1836);
nor U2424 (N_2424,N_2069,N_2109);
nor U2425 (N_2425,N_2056,N_1628);
nor U2426 (N_2426,N_1601,N_1528);
and U2427 (N_2427,N_1998,N_1910);
xnor U2428 (N_2428,N_1880,N_1583);
nor U2429 (N_2429,N_2067,N_1522);
and U2430 (N_2430,N_1916,N_2074);
nand U2431 (N_2431,N_1803,N_1651);
and U2432 (N_2432,N_2247,N_2200);
nand U2433 (N_2433,N_1661,N_1727);
or U2434 (N_2434,N_2192,N_2023);
or U2435 (N_2435,N_2118,N_1644);
nor U2436 (N_2436,N_2219,N_1804);
xor U2437 (N_2437,N_1678,N_1665);
nand U2438 (N_2438,N_1982,N_1731);
and U2439 (N_2439,N_1555,N_2230);
nor U2440 (N_2440,N_1900,N_2182);
nand U2441 (N_2441,N_1714,N_2044);
xnor U2442 (N_2442,N_1970,N_1810);
and U2443 (N_2443,N_1721,N_2052);
nand U2444 (N_2444,N_1793,N_1537);
or U2445 (N_2445,N_2226,N_1524);
nand U2446 (N_2446,N_1542,N_2135);
xnor U2447 (N_2447,N_1846,N_2105);
nor U2448 (N_2448,N_1783,N_1519);
and U2449 (N_2449,N_2045,N_1707);
and U2450 (N_2450,N_2240,N_1869);
and U2451 (N_2451,N_1796,N_2007);
nand U2452 (N_2452,N_1619,N_1535);
nor U2453 (N_2453,N_2006,N_1739);
nand U2454 (N_2454,N_2196,N_1851);
or U2455 (N_2455,N_1933,N_1558);
nand U2456 (N_2456,N_2049,N_1790);
or U2457 (N_2457,N_2000,N_2008);
nand U2458 (N_2458,N_1740,N_2058);
or U2459 (N_2459,N_1562,N_1949);
and U2460 (N_2460,N_1589,N_1833);
and U2461 (N_2461,N_2086,N_2215);
xor U2462 (N_2462,N_1888,N_2037);
nor U2463 (N_2463,N_1768,N_2158);
or U2464 (N_2464,N_2212,N_1914);
nor U2465 (N_2465,N_2162,N_2082);
nor U2466 (N_2466,N_1988,N_2140);
xnor U2467 (N_2467,N_2031,N_1917);
and U2468 (N_2468,N_1514,N_1769);
nand U2469 (N_2469,N_2177,N_2217);
nand U2470 (N_2470,N_1770,N_1856);
nor U2471 (N_2471,N_1532,N_1995);
xnor U2472 (N_2472,N_1971,N_1515);
or U2473 (N_2473,N_2249,N_1923);
nand U2474 (N_2474,N_2026,N_1912);
xor U2475 (N_2475,N_1748,N_1974);
or U2476 (N_2476,N_2188,N_2205);
xnor U2477 (N_2477,N_1684,N_2220);
nor U2478 (N_2478,N_1668,N_1588);
nand U2479 (N_2479,N_2165,N_2036);
or U2480 (N_2480,N_2059,N_1709);
nor U2481 (N_2481,N_2235,N_1919);
nand U2482 (N_2482,N_1591,N_1962);
nor U2483 (N_2483,N_2022,N_1580);
nand U2484 (N_2484,N_1539,N_1872);
nand U2485 (N_2485,N_2221,N_1653);
nand U2486 (N_2486,N_1728,N_1886);
nor U2487 (N_2487,N_2076,N_1618);
xnor U2488 (N_2488,N_1842,N_1533);
or U2489 (N_2489,N_2204,N_1868);
or U2490 (N_2490,N_2085,N_1981);
nor U2491 (N_2491,N_1689,N_2210);
nand U2492 (N_2492,N_1602,N_2127);
and U2493 (N_2493,N_1538,N_1664);
or U2494 (N_2494,N_1687,N_1606);
or U2495 (N_2495,N_1573,N_2244);
xnor U2496 (N_2496,N_1615,N_1504);
or U2497 (N_2497,N_2138,N_2183);
nand U2498 (N_2498,N_1898,N_1929);
nor U2499 (N_2499,N_1878,N_1550);
nor U2500 (N_2500,N_2061,N_1545);
nand U2501 (N_2501,N_1507,N_2232);
and U2502 (N_2502,N_1843,N_2099);
or U2503 (N_2503,N_1530,N_1946);
xnor U2504 (N_2504,N_2157,N_1940);
nand U2505 (N_2505,N_1683,N_2048);
and U2506 (N_2506,N_2213,N_1837);
and U2507 (N_2507,N_1907,N_2194);
or U2508 (N_2508,N_2072,N_2243);
nand U2509 (N_2509,N_2152,N_1857);
xor U2510 (N_2510,N_1625,N_2228);
nor U2511 (N_2511,N_1598,N_1702);
nor U2512 (N_2512,N_2010,N_1774);
xnor U2513 (N_2513,N_1662,N_1956);
xor U2514 (N_2514,N_1723,N_1989);
nor U2515 (N_2515,N_1968,N_1924);
nand U2516 (N_2516,N_2090,N_1722);
or U2517 (N_2517,N_2139,N_1546);
and U2518 (N_2518,N_2218,N_1594);
or U2519 (N_2519,N_1617,N_1913);
and U2520 (N_2520,N_2041,N_2149);
nand U2521 (N_2521,N_2187,N_1776);
or U2522 (N_2522,N_2229,N_1819);
or U2523 (N_2523,N_1682,N_2231);
nand U2524 (N_2524,N_1972,N_1969);
and U2525 (N_2525,N_1513,N_1547);
nor U2526 (N_2526,N_2144,N_2073);
or U2527 (N_2527,N_2110,N_1939);
xor U2528 (N_2528,N_2224,N_1771);
xnor U2529 (N_2529,N_2089,N_2083);
and U2530 (N_2530,N_1500,N_2079);
nand U2531 (N_2531,N_1703,N_1540);
or U2532 (N_2532,N_1579,N_2003);
nand U2533 (N_2533,N_2013,N_1733);
and U2534 (N_2534,N_1593,N_1791);
nor U2535 (N_2535,N_2084,N_2062);
xnor U2536 (N_2536,N_2112,N_1965);
or U2537 (N_2537,N_1521,N_2064);
nor U2538 (N_2538,N_1960,N_1959);
or U2539 (N_2539,N_1877,N_1646);
xor U2540 (N_2540,N_2054,N_1725);
xor U2541 (N_2541,N_1554,N_1884);
xor U2542 (N_2542,N_2208,N_1676);
and U2543 (N_2543,N_1574,N_2103);
nor U2544 (N_2544,N_1614,N_1508);
or U2545 (N_2545,N_1824,N_2216);
nand U2546 (N_2546,N_2203,N_1760);
nand U2547 (N_2547,N_1616,N_2055);
and U2548 (N_2548,N_2136,N_2093);
nand U2549 (N_2549,N_1823,N_1749);
xor U2550 (N_2550,N_1961,N_1544);
nor U2551 (N_2551,N_1623,N_1863);
xor U2552 (N_2552,N_1963,N_1918);
or U2553 (N_2553,N_1826,N_1634);
or U2554 (N_2554,N_1667,N_2186);
nand U2555 (N_2555,N_1892,N_1735);
xor U2556 (N_2556,N_1754,N_1947);
or U2557 (N_2557,N_1814,N_1556);
nand U2558 (N_2558,N_2107,N_1742);
or U2559 (N_2559,N_1789,N_1766);
or U2560 (N_2560,N_1812,N_2166);
nand U2561 (N_2561,N_1738,N_2011);
or U2562 (N_2562,N_1597,N_1586);
or U2563 (N_2563,N_2134,N_2046);
xor U2564 (N_2564,N_1681,N_1853);
xnor U2565 (N_2565,N_2002,N_1529);
xnor U2566 (N_2566,N_1777,N_2117);
xor U2567 (N_2567,N_2155,N_1859);
or U2568 (N_2568,N_1964,N_1672);
or U2569 (N_2569,N_1953,N_2081);
nor U2570 (N_2570,N_1934,N_1582);
and U2571 (N_2571,N_1610,N_1549);
or U2572 (N_2572,N_2095,N_1690);
nand U2573 (N_2573,N_2091,N_2027);
xnor U2574 (N_2574,N_1630,N_1899);
xor U2575 (N_2575,N_2206,N_1557);
nand U2576 (N_2576,N_2020,N_1590);
and U2577 (N_2577,N_1794,N_2066);
or U2578 (N_2578,N_1761,N_1854);
or U2579 (N_2579,N_1724,N_1821);
nor U2580 (N_2580,N_1685,N_1726);
and U2581 (N_2581,N_1505,N_2043);
nor U2582 (N_2582,N_1612,N_2168);
nand U2583 (N_2583,N_1954,N_1717);
and U2584 (N_2584,N_1677,N_2029);
nor U2585 (N_2585,N_2174,N_1699);
xor U2586 (N_2586,N_1806,N_2145);
xor U2587 (N_2587,N_1747,N_2087);
xnor U2588 (N_2588,N_1763,N_1673);
or U2589 (N_2589,N_1552,N_1921);
or U2590 (N_2590,N_1650,N_2075);
or U2591 (N_2591,N_2028,N_1531);
nor U2592 (N_2592,N_1987,N_2051);
nor U2593 (N_2593,N_1715,N_2173);
or U2594 (N_2594,N_1866,N_2094);
xnor U2595 (N_2595,N_1729,N_1809);
xnor U2596 (N_2596,N_1817,N_1945);
nand U2597 (N_2597,N_2098,N_1931);
xnor U2598 (N_2598,N_1712,N_1744);
and U2599 (N_2599,N_2214,N_2198);
xor U2600 (N_2600,N_1643,N_1802);
or U2601 (N_2601,N_1503,N_2047);
nand U2602 (N_2602,N_1788,N_1534);
nor U2603 (N_2603,N_1864,N_1510);
nor U2604 (N_2604,N_1656,N_1711);
xnor U2605 (N_2605,N_2179,N_1675);
and U2606 (N_2606,N_2163,N_2248);
and U2607 (N_2607,N_1822,N_1902);
xor U2608 (N_2608,N_1730,N_1716);
nor U2609 (N_2609,N_2133,N_1621);
nor U2610 (N_2610,N_1897,N_1781);
nor U2611 (N_2611,N_1865,N_2137);
nand U2612 (N_2612,N_2060,N_1891);
nand U2613 (N_2613,N_1993,N_1603);
nand U2614 (N_2614,N_1887,N_1811);
and U2615 (N_2615,N_1977,N_1925);
or U2616 (N_2616,N_1737,N_2209);
and U2617 (N_2617,N_1501,N_1990);
xor U2618 (N_2618,N_1581,N_1705);
xor U2619 (N_2619,N_1839,N_1955);
nor U2620 (N_2620,N_1686,N_1660);
nand U2621 (N_2621,N_1901,N_2239);
and U2622 (N_2622,N_1765,N_1585);
nand U2623 (N_2623,N_1780,N_1563);
or U2624 (N_2624,N_1873,N_2227);
xnor U2625 (N_2625,N_1851,N_2005);
and U2626 (N_2626,N_1949,N_1752);
xor U2627 (N_2627,N_1762,N_2158);
or U2628 (N_2628,N_1842,N_1580);
nand U2629 (N_2629,N_2163,N_2195);
xnor U2630 (N_2630,N_1873,N_2044);
nor U2631 (N_2631,N_1896,N_1851);
or U2632 (N_2632,N_1591,N_1662);
nor U2633 (N_2633,N_1959,N_1529);
nor U2634 (N_2634,N_1634,N_1971);
or U2635 (N_2635,N_1891,N_2103);
or U2636 (N_2636,N_1817,N_2019);
or U2637 (N_2637,N_1713,N_1512);
or U2638 (N_2638,N_1787,N_1832);
xor U2639 (N_2639,N_1583,N_2155);
and U2640 (N_2640,N_2136,N_2022);
nor U2641 (N_2641,N_1755,N_1888);
nor U2642 (N_2642,N_2074,N_1844);
xor U2643 (N_2643,N_2148,N_2105);
nand U2644 (N_2644,N_2156,N_1842);
nor U2645 (N_2645,N_2007,N_1858);
nor U2646 (N_2646,N_1673,N_2052);
xnor U2647 (N_2647,N_2043,N_2080);
and U2648 (N_2648,N_2219,N_1796);
nor U2649 (N_2649,N_1992,N_1990);
or U2650 (N_2650,N_1575,N_1805);
nor U2651 (N_2651,N_1788,N_1643);
and U2652 (N_2652,N_2107,N_1524);
xnor U2653 (N_2653,N_2101,N_1742);
nor U2654 (N_2654,N_2074,N_1851);
and U2655 (N_2655,N_1908,N_1905);
nand U2656 (N_2656,N_1597,N_1706);
nor U2657 (N_2657,N_1586,N_1805);
nand U2658 (N_2658,N_2088,N_2206);
and U2659 (N_2659,N_1696,N_1685);
or U2660 (N_2660,N_2229,N_1547);
or U2661 (N_2661,N_1982,N_1604);
and U2662 (N_2662,N_2165,N_1542);
or U2663 (N_2663,N_2175,N_2067);
or U2664 (N_2664,N_1886,N_2013);
or U2665 (N_2665,N_1922,N_1785);
or U2666 (N_2666,N_1669,N_1694);
or U2667 (N_2667,N_2060,N_2129);
nand U2668 (N_2668,N_2200,N_2124);
nor U2669 (N_2669,N_2015,N_2153);
xnor U2670 (N_2670,N_1694,N_2177);
or U2671 (N_2671,N_2167,N_2228);
nand U2672 (N_2672,N_2173,N_2155);
or U2673 (N_2673,N_1989,N_1572);
nor U2674 (N_2674,N_1850,N_1924);
nor U2675 (N_2675,N_1603,N_1761);
and U2676 (N_2676,N_1805,N_1639);
or U2677 (N_2677,N_2000,N_1862);
or U2678 (N_2678,N_1605,N_1556);
or U2679 (N_2679,N_1965,N_1760);
or U2680 (N_2680,N_1884,N_2100);
and U2681 (N_2681,N_1780,N_1601);
nor U2682 (N_2682,N_1560,N_1527);
nand U2683 (N_2683,N_1975,N_1574);
or U2684 (N_2684,N_2098,N_1985);
or U2685 (N_2685,N_1685,N_1660);
and U2686 (N_2686,N_1837,N_2042);
and U2687 (N_2687,N_2236,N_2017);
nor U2688 (N_2688,N_1839,N_1539);
nor U2689 (N_2689,N_2180,N_1584);
or U2690 (N_2690,N_1941,N_1926);
xnor U2691 (N_2691,N_2154,N_2035);
and U2692 (N_2692,N_1798,N_2079);
xnor U2693 (N_2693,N_1536,N_2007);
and U2694 (N_2694,N_1701,N_2133);
or U2695 (N_2695,N_1752,N_1682);
nor U2696 (N_2696,N_1927,N_1986);
nor U2697 (N_2697,N_1651,N_2209);
nor U2698 (N_2698,N_1913,N_1869);
nand U2699 (N_2699,N_1785,N_1595);
xnor U2700 (N_2700,N_1959,N_1790);
nor U2701 (N_2701,N_2006,N_1688);
xor U2702 (N_2702,N_2032,N_1706);
nor U2703 (N_2703,N_1957,N_1505);
xor U2704 (N_2704,N_1805,N_2090);
xor U2705 (N_2705,N_2028,N_1749);
or U2706 (N_2706,N_1880,N_2029);
nand U2707 (N_2707,N_1771,N_2160);
xnor U2708 (N_2708,N_2157,N_2021);
or U2709 (N_2709,N_2072,N_1778);
nand U2710 (N_2710,N_2067,N_2212);
and U2711 (N_2711,N_1586,N_2006);
nand U2712 (N_2712,N_1925,N_1847);
or U2713 (N_2713,N_1822,N_2021);
and U2714 (N_2714,N_1966,N_2120);
xor U2715 (N_2715,N_1702,N_2165);
or U2716 (N_2716,N_1918,N_2028);
and U2717 (N_2717,N_2135,N_1889);
nor U2718 (N_2718,N_1604,N_1736);
nor U2719 (N_2719,N_1806,N_1946);
nor U2720 (N_2720,N_1963,N_1786);
or U2721 (N_2721,N_1596,N_2142);
and U2722 (N_2722,N_1679,N_1841);
nor U2723 (N_2723,N_2217,N_1515);
or U2724 (N_2724,N_2170,N_1666);
nor U2725 (N_2725,N_1800,N_1632);
nor U2726 (N_2726,N_1801,N_1655);
nor U2727 (N_2727,N_2108,N_1689);
and U2728 (N_2728,N_1843,N_2166);
or U2729 (N_2729,N_2120,N_2075);
nand U2730 (N_2730,N_1520,N_1721);
xnor U2731 (N_2731,N_1788,N_2187);
or U2732 (N_2732,N_1872,N_1725);
or U2733 (N_2733,N_2222,N_1702);
or U2734 (N_2734,N_1683,N_2123);
or U2735 (N_2735,N_1622,N_2035);
xnor U2736 (N_2736,N_1754,N_2190);
xor U2737 (N_2737,N_2150,N_2247);
nor U2738 (N_2738,N_1805,N_2196);
nor U2739 (N_2739,N_2159,N_2138);
or U2740 (N_2740,N_2127,N_2097);
or U2741 (N_2741,N_1632,N_2002);
or U2742 (N_2742,N_1809,N_1698);
or U2743 (N_2743,N_1722,N_1554);
xor U2744 (N_2744,N_1699,N_1973);
nand U2745 (N_2745,N_1694,N_1681);
or U2746 (N_2746,N_1823,N_2145);
or U2747 (N_2747,N_1683,N_2152);
or U2748 (N_2748,N_1760,N_2240);
or U2749 (N_2749,N_1879,N_1551);
or U2750 (N_2750,N_1846,N_2011);
xnor U2751 (N_2751,N_1602,N_1906);
xnor U2752 (N_2752,N_2064,N_1624);
xnor U2753 (N_2753,N_1502,N_1647);
or U2754 (N_2754,N_1561,N_2113);
or U2755 (N_2755,N_1773,N_1607);
and U2756 (N_2756,N_1508,N_2161);
xnor U2757 (N_2757,N_1727,N_2148);
nor U2758 (N_2758,N_1964,N_2208);
and U2759 (N_2759,N_1749,N_1777);
or U2760 (N_2760,N_1632,N_1514);
nor U2761 (N_2761,N_1790,N_1506);
nand U2762 (N_2762,N_2151,N_1861);
or U2763 (N_2763,N_1737,N_1571);
xnor U2764 (N_2764,N_1512,N_1898);
and U2765 (N_2765,N_2181,N_2236);
xor U2766 (N_2766,N_1676,N_1505);
nor U2767 (N_2767,N_1601,N_1914);
nor U2768 (N_2768,N_2032,N_1594);
or U2769 (N_2769,N_2162,N_2059);
or U2770 (N_2770,N_1664,N_1818);
and U2771 (N_2771,N_2208,N_1879);
xnor U2772 (N_2772,N_1921,N_2115);
nand U2773 (N_2773,N_2212,N_1750);
nor U2774 (N_2774,N_1582,N_1510);
or U2775 (N_2775,N_2033,N_2123);
or U2776 (N_2776,N_2161,N_1541);
nand U2777 (N_2777,N_1528,N_2091);
or U2778 (N_2778,N_1998,N_1548);
xnor U2779 (N_2779,N_1533,N_1761);
xor U2780 (N_2780,N_1651,N_1886);
xor U2781 (N_2781,N_1733,N_1557);
nand U2782 (N_2782,N_1747,N_1945);
nand U2783 (N_2783,N_2058,N_1994);
nand U2784 (N_2784,N_2245,N_1730);
or U2785 (N_2785,N_1600,N_1958);
or U2786 (N_2786,N_2239,N_1565);
xnor U2787 (N_2787,N_2057,N_2190);
xnor U2788 (N_2788,N_2152,N_1848);
or U2789 (N_2789,N_1869,N_1630);
and U2790 (N_2790,N_1798,N_1906);
nor U2791 (N_2791,N_1829,N_2057);
nor U2792 (N_2792,N_1792,N_1824);
xor U2793 (N_2793,N_1919,N_1766);
and U2794 (N_2794,N_1770,N_1829);
or U2795 (N_2795,N_1590,N_2230);
nor U2796 (N_2796,N_1695,N_2101);
or U2797 (N_2797,N_1799,N_2004);
or U2798 (N_2798,N_1595,N_1836);
nand U2799 (N_2799,N_2049,N_1532);
xnor U2800 (N_2800,N_1928,N_1777);
nand U2801 (N_2801,N_2029,N_1526);
or U2802 (N_2802,N_1929,N_2030);
and U2803 (N_2803,N_1884,N_1662);
nand U2804 (N_2804,N_1821,N_2101);
and U2805 (N_2805,N_1828,N_1942);
and U2806 (N_2806,N_1536,N_1898);
and U2807 (N_2807,N_2127,N_2130);
nand U2808 (N_2808,N_1623,N_1702);
and U2809 (N_2809,N_2108,N_1832);
and U2810 (N_2810,N_2218,N_1571);
xnor U2811 (N_2811,N_1842,N_1986);
nand U2812 (N_2812,N_1647,N_1682);
xor U2813 (N_2813,N_2158,N_2175);
nor U2814 (N_2814,N_1576,N_1829);
nor U2815 (N_2815,N_1986,N_1566);
nor U2816 (N_2816,N_1699,N_1786);
nand U2817 (N_2817,N_2143,N_1705);
nand U2818 (N_2818,N_1919,N_2085);
xnor U2819 (N_2819,N_1856,N_2036);
nand U2820 (N_2820,N_1966,N_2119);
or U2821 (N_2821,N_1658,N_2127);
or U2822 (N_2822,N_1951,N_1776);
xor U2823 (N_2823,N_1802,N_1583);
nor U2824 (N_2824,N_2128,N_1846);
xnor U2825 (N_2825,N_1526,N_1746);
and U2826 (N_2826,N_1978,N_1697);
nand U2827 (N_2827,N_1509,N_1713);
nor U2828 (N_2828,N_1699,N_2203);
nand U2829 (N_2829,N_1552,N_1624);
or U2830 (N_2830,N_1821,N_1880);
xor U2831 (N_2831,N_2235,N_2013);
and U2832 (N_2832,N_1883,N_1654);
and U2833 (N_2833,N_1938,N_1841);
or U2834 (N_2834,N_2029,N_1641);
or U2835 (N_2835,N_2186,N_1728);
nand U2836 (N_2836,N_1707,N_1900);
or U2837 (N_2837,N_1919,N_1508);
or U2838 (N_2838,N_1628,N_2058);
or U2839 (N_2839,N_2108,N_2164);
nand U2840 (N_2840,N_2206,N_2025);
or U2841 (N_2841,N_2063,N_1610);
xor U2842 (N_2842,N_2045,N_2104);
nand U2843 (N_2843,N_1762,N_1835);
nand U2844 (N_2844,N_1665,N_1608);
nor U2845 (N_2845,N_1983,N_1771);
or U2846 (N_2846,N_1623,N_1681);
or U2847 (N_2847,N_1585,N_2229);
nor U2848 (N_2848,N_1771,N_1765);
nand U2849 (N_2849,N_1559,N_1508);
nand U2850 (N_2850,N_2070,N_1977);
nand U2851 (N_2851,N_2163,N_1998);
or U2852 (N_2852,N_1563,N_1925);
xnor U2853 (N_2853,N_1565,N_2132);
or U2854 (N_2854,N_2178,N_2222);
or U2855 (N_2855,N_1717,N_1773);
xor U2856 (N_2856,N_1906,N_2210);
or U2857 (N_2857,N_1632,N_1760);
xnor U2858 (N_2858,N_1819,N_2138);
nor U2859 (N_2859,N_2165,N_2047);
xnor U2860 (N_2860,N_1995,N_1688);
nor U2861 (N_2861,N_2039,N_1822);
xnor U2862 (N_2862,N_1776,N_1904);
xnor U2863 (N_2863,N_2079,N_1594);
or U2864 (N_2864,N_1750,N_1716);
nand U2865 (N_2865,N_2243,N_1859);
xor U2866 (N_2866,N_1974,N_2069);
or U2867 (N_2867,N_2227,N_2086);
or U2868 (N_2868,N_1620,N_1982);
nand U2869 (N_2869,N_2127,N_2208);
nor U2870 (N_2870,N_2223,N_1901);
xor U2871 (N_2871,N_2173,N_1931);
or U2872 (N_2872,N_1654,N_1905);
nor U2873 (N_2873,N_1590,N_1699);
and U2874 (N_2874,N_1567,N_1559);
nor U2875 (N_2875,N_1729,N_2130);
xnor U2876 (N_2876,N_1872,N_2215);
or U2877 (N_2877,N_2019,N_2136);
nor U2878 (N_2878,N_1587,N_1911);
and U2879 (N_2879,N_1921,N_1562);
nor U2880 (N_2880,N_1561,N_2201);
nor U2881 (N_2881,N_2141,N_1775);
nor U2882 (N_2882,N_2008,N_1872);
or U2883 (N_2883,N_2036,N_2233);
or U2884 (N_2884,N_1882,N_1506);
nand U2885 (N_2885,N_1517,N_1585);
and U2886 (N_2886,N_1748,N_1571);
and U2887 (N_2887,N_1941,N_1542);
or U2888 (N_2888,N_1864,N_2061);
xnor U2889 (N_2889,N_1583,N_1670);
nor U2890 (N_2890,N_1959,N_1547);
nor U2891 (N_2891,N_2165,N_1772);
nand U2892 (N_2892,N_1735,N_1848);
nand U2893 (N_2893,N_1935,N_2164);
or U2894 (N_2894,N_1800,N_1525);
nor U2895 (N_2895,N_1667,N_2234);
nor U2896 (N_2896,N_1812,N_1535);
or U2897 (N_2897,N_1832,N_2160);
nor U2898 (N_2898,N_2063,N_1830);
or U2899 (N_2899,N_1900,N_1669);
nand U2900 (N_2900,N_1785,N_2211);
xor U2901 (N_2901,N_2219,N_1637);
or U2902 (N_2902,N_2053,N_1930);
nand U2903 (N_2903,N_1990,N_1636);
and U2904 (N_2904,N_1673,N_1753);
xnor U2905 (N_2905,N_1509,N_2201);
or U2906 (N_2906,N_1731,N_1797);
nor U2907 (N_2907,N_1956,N_2164);
nand U2908 (N_2908,N_1946,N_1800);
and U2909 (N_2909,N_1783,N_1743);
or U2910 (N_2910,N_1827,N_1539);
or U2911 (N_2911,N_1747,N_1595);
or U2912 (N_2912,N_2114,N_2045);
and U2913 (N_2913,N_1784,N_1682);
and U2914 (N_2914,N_1697,N_1949);
and U2915 (N_2915,N_1661,N_1597);
nand U2916 (N_2916,N_1806,N_1599);
or U2917 (N_2917,N_1688,N_1657);
nand U2918 (N_2918,N_2149,N_1984);
xnor U2919 (N_2919,N_1555,N_2198);
xor U2920 (N_2920,N_1677,N_1525);
xnor U2921 (N_2921,N_1755,N_1930);
and U2922 (N_2922,N_2198,N_1576);
and U2923 (N_2923,N_2013,N_1684);
and U2924 (N_2924,N_1640,N_1657);
nor U2925 (N_2925,N_1748,N_2051);
nor U2926 (N_2926,N_1582,N_2130);
or U2927 (N_2927,N_2179,N_1791);
nor U2928 (N_2928,N_2081,N_2172);
nand U2929 (N_2929,N_1836,N_2212);
nor U2930 (N_2930,N_1818,N_1858);
nand U2931 (N_2931,N_1622,N_1838);
xor U2932 (N_2932,N_1880,N_1561);
nand U2933 (N_2933,N_1811,N_2058);
xor U2934 (N_2934,N_2212,N_1692);
nand U2935 (N_2935,N_1929,N_1594);
nor U2936 (N_2936,N_1959,N_1889);
xnor U2937 (N_2937,N_1947,N_1872);
or U2938 (N_2938,N_1829,N_1730);
nor U2939 (N_2939,N_1926,N_1771);
nand U2940 (N_2940,N_2206,N_2086);
and U2941 (N_2941,N_1872,N_2135);
nand U2942 (N_2942,N_1553,N_2033);
nand U2943 (N_2943,N_1892,N_1899);
nor U2944 (N_2944,N_2068,N_1552);
or U2945 (N_2945,N_2151,N_1863);
and U2946 (N_2946,N_1805,N_1537);
or U2947 (N_2947,N_1533,N_1824);
nor U2948 (N_2948,N_1714,N_1646);
xnor U2949 (N_2949,N_1519,N_2221);
nand U2950 (N_2950,N_2155,N_1786);
xnor U2951 (N_2951,N_1987,N_1835);
xnor U2952 (N_2952,N_1842,N_2112);
and U2953 (N_2953,N_2071,N_1797);
or U2954 (N_2954,N_2117,N_1704);
nand U2955 (N_2955,N_1681,N_1550);
xnor U2956 (N_2956,N_1781,N_1663);
or U2957 (N_2957,N_1559,N_1896);
nor U2958 (N_2958,N_1527,N_2086);
xor U2959 (N_2959,N_1563,N_1604);
nand U2960 (N_2960,N_2119,N_1988);
nor U2961 (N_2961,N_1665,N_1951);
xnor U2962 (N_2962,N_1751,N_1519);
xor U2963 (N_2963,N_1657,N_1836);
and U2964 (N_2964,N_1831,N_1956);
nor U2965 (N_2965,N_1942,N_1774);
nand U2966 (N_2966,N_2083,N_1980);
nor U2967 (N_2967,N_1624,N_1978);
or U2968 (N_2968,N_2198,N_1767);
and U2969 (N_2969,N_1583,N_1853);
nand U2970 (N_2970,N_1738,N_1960);
xor U2971 (N_2971,N_1673,N_1640);
or U2972 (N_2972,N_1870,N_2150);
xnor U2973 (N_2973,N_2017,N_2181);
and U2974 (N_2974,N_1718,N_1845);
or U2975 (N_2975,N_1772,N_1715);
or U2976 (N_2976,N_2217,N_2224);
nand U2977 (N_2977,N_2168,N_1500);
nand U2978 (N_2978,N_1586,N_1504);
and U2979 (N_2979,N_2063,N_2219);
nor U2980 (N_2980,N_1652,N_2021);
xor U2981 (N_2981,N_1681,N_1854);
and U2982 (N_2982,N_1881,N_1714);
nor U2983 (N_2983,N_1805,N_1890);
and U2984 (N_2984,N_1820,N_2230);
and U2985 (N_2985,N_1987,N_1653);
nor U2986 (N_2986,N_1674,N_1705);
nand U2987 (N_2987,N_1546,N_1564);
xnor U2988 (N_2988,N_1725,N_1638);
xor U2989 (N_2989,N_1815,N_1584);
nand U2990 (N_2990,N_1847,N_1610);
and U2991 (N_2991,N_1994,N_2166);
xnor U2992 (N_2992,N_2119,N_2187);
and U2993 (N_2993,N_1967,N_1875);
nor U2994 (N_2994,N_1717,N_2183);
nand U2995 (N_2995,N_1991,N_1646);
or U2996 (N_2996,N_1554,N_1911);
nand U2997 (N_2997,N_1983,N_1765);
and U2998 (N_2998,N_2172,N_1818);
nand U2999 (N_2999,N_1543,N_1752);
and U3000 (N_3000,N_2721,N_2419);
xor U3001 (N_3001,N_2988,N_2778);
and U3002 (N_3002,N_2411,N_2975);
nor U3003 (N_3003,N_2924,N_2341);
nand U3004 (N_3004,N_2511,N_2675);
xnor U3005 (N_3005,N_2829,N_2409);
and U3006 (N_3006,N_2361,N_2725);
nor U3007 (N_3007,N_2870,N_2743);
xor U3008 (N_3008,N_2479,N_2817);
xor U3009 (N_3009,N_2523,N_2971);
xnor U3010 (N_3010,N_2764,N_2640);
xor U3011 (N_3011,N_2755,N_2633);
or U3012 (N_3012,N_2335,N_2612);
and U3013 (N_3013,N_2587,N_2493);
nand U3014 (N_3014,N_2626,N_2739);
nor U3015 (N_3015,N_2550,N_2489);
xor U3016 (N_3016,N_2426,N_2660);
nand U3017 (N_3017,N_2785,N_2397);
or U3018 (N_3018,N_2720,N_2392);
or U3019 (N_3019,N_2637,N_2698);
or U3020 (N_3020,N_2256,N_2322);
nand U3021 (N_3021,N_2429,N_2983);
nand U3022 (N_3022,N_2485,N_2621);
xnor U3023 (N_3023,N_2330,N_2490);
xor U3024 (N_3024,N_2541,N_2772);
nand U3025 (N_3025,N_2576,N_2307);
xor U3026 (N_3026,N_2629,N_2994);
nor U3027 (N_3027,N_2303,N_2468);
nor U3028 (N_3028,N_2816,N_2950);
nand U3029 (N_3029,N_2966,N_2747);
nor U3030 (N_3030,N_2538,N_2446);
or U3031 (N_3031,N_2367,N_2590);
nand U3032 (N_3032,N_2393,N_2893);
xnor U3033 (N_3033,N_2390,N_2345);
nand U3034 (N_3034,N_2374,N_2564);
nand U3035 (N_3035,N_2664,N_2578);
and U3036 (N_3036,N_2993,N_2687);
or U3037 (N_3037,N_2467,N_2686);
nor U3038 (N_3038,N_2604,N_2445);
xor U3039 (N_3039,N_2466,N_2992);
and U3040 (N_3040,N_2391,N_2413);
or U3041 (N_3041,N_2921,N_2892);
or U3042 (N_3042,N_2338,N_2843);
and U3043 (N_3043,N_2292,N_2317);
nor U3044 (N_3044,N_2585,N_2706);
nor U3045 (N_3045,N_2423,N_2812);
nor U3046 (N_3046,N_2460,N_2737);
or U3047 (N_3047,N_2279,N_2566);
nand U3048 (N_3048,N_2630,N_2922);
or U3049 (N_3049,N_2535,N_2436);
or U3050 (N_3050,N_2592,N_2857);
or U3051 (N_3051,N_2376,N_2299);
and U3052 (N_3052,N_2635,N_2884);
or U3053 (N_3053,N_2568,N_2499);
xor U3054 (N_3054,N_2465,N_2839);
xor U3055 (N_3055,N_2744,N_2919);
and U3056 (N_3056,N_2909,N_2571);
nand U3057 (N_3057,N_2400,N_2799);
nor U3058 (N_3058,N_2756,N_2622);
nand U3059 (N_3059,N_2565,N_2741);
xnor U3060 (N_3060,N_2555,N_2252);
or U3061 (N_3061,N_2320,N_2728);
or U3062 (N_3062,N_2806,N_2949);
nand U3063 (N_3063,N_2980,N_2701);
or U3064 (N_3064,N_2934,N_2682);
xnor U3065 (N_3065,N_2900,N_2653);
nor U3066 (N_3066,N_2517,N_2608);
nor U3067 (N_3067,N_2733,N_2286);
or U3068 (N_3068,N_2654,N_2936);
nand U3069 (N_3069,N_2570,N_2960);
nor U3070 (N_3070,N_2582,N_2483);
and U3071 (N_3071,N_2697,N_2757);
xor U3072 (N_3072,N_2255,N_2674);
or U3073 (N_3073,N_2476,N_2923);
and U3074 (N_3074,N_2718,N_2288);
xnor U3075 (N_3075,N_2495,N_2984);
xor U3076 (N_3076,N_2845,N_2362);
nand U3077 (N_3077,N_2646,N_2328);
nand U3078 (N_3078,N_2827,N_2280);
nor U3079 (N_3079,N_2888,N_2681);
or U3080 (N_3080,N_2868,N_2965);
and U3081 (N_3081,N_2515,N_2628);
nor U3082 (N_3082,N_2978,N_2405);
and U3083 (N_3083,N_2650,N_2352);
and U3084 (N_3084,N_2902,N_2589);
and U3085 (N_3085,N_2441,N_2959);
or U3086 (N_3086,N_2266,N_2324);
nand U3087 (N_3087,N_2901,N_2793);
xnor U3088 (N_3088,N_2879,N_2569);
nand U3089 (N_3089,N_2583,N_2645);
or U3090 (N_3090,N_2309,N_2259);
and U3091 (N_3091,N_2351,N_2418);
or U3092 (N_3092,N_2285,N_2678);
nand U3093 (N_3093,N_2903,N_2688);
or U3094 (N_3094,N_2683,N_2987);
or U3095 (N_3095,N_2602,N_2463);
nand U3096 (N_3096,N_2863,N_2321);
xnor U3097 (N_3097,N_2616,N_2337);
nand U3098 (N_3098,N_2549,N_2703);
nor U3099 (N_3099,N_2663,N_2794);
or U3100 (N_3100,N_2492,N_2265);
xnor U3101 (N_3101,N_2841,N_2356);
xor U3102 (N_3102,N_2729,N_2671);
or U3103 (N_3103,N_2509,N_2679);
nand U3104 (N_3104,N_2780,N_2540);
or U3105 (N_3105,N_2908,N_2355);
or U3106 (N_3106,N_2749,N_2779);
and U3107 (N_3107,N_2810,N_2264);
and U3108 (N_3108,N_2271,N_2849);
nor U3109 (N_3109,N_2563,N_2472);
nor U3110 (N_3110,N_2431,N_2847);
nand U3111 (N_3111,N_2942,N_2991);
or U3112 (N_3112,N_2935,N_2680);
xnor U3113 (N_3113,N_2599,N_2801);
nand U3114 (N_3114,N_2883,N_2761);
nor U3115 (N_3115,N_2972,N_2954);
nor U3116 (N_3116,N_2709,N_2634);
and U3117 (N_3117,N_2753,N_2933);
and U3118 (N_3118,N_2605,N_2543);
nand U3119 (N_3119,N_2363,N_2291);
and U3120 (N_3120,N_2889,N_2742);
xor U3121 (N_3121,N_2389,N_2802);
nor U3122 (N_3122,N_2620,N_2677);
nor U3123 (N_3123,N_2267,N_2943);
xnor U3124 (N_3124,N_2846,N_2912);
nand U3125 (N_3125,N_2357,N_2876);
nor U3126 (N_3126,N_2504,N_2910);
and U3127 (N_3127,N_2560,N_2736);
nand U3128 (N_3128,N_2808,N_2537);
xor U3129 (N_3129,N_2520,N_2977);
or U3130 (N_3130,N_2974,N_2258);
and U3131 (N_3131,N_2457,N_2758);
xor U3132 (N_3132,N_2918,N_2371);
nor U3133 (N_3133,N_2294,N_2773);
xor U3134 (N_3134,N_2643,N_2907);
or U3135 (N_3135,N_2751,N_2562);
xor U3136 (N_3136,N_2430,N_2416);
nand U3137 (N_3137,N_2450,N_2850);
nand U3138 (N_3138,N_2407,N_2383);
nand U3139 (N_3139,N_2726,N_2348);
xor U3140 (N_3140,N_2716,N_2349);
nor U3141 (N_3141,N_2260,N_2314);
xor U3142 (N_3142,N_2359,N_2886);
or U3143 (N_3143,N_2864,N_2783);
or U3144 (N_3144,N_2860,N_2296);
xor U3145 (N_3145,N_2916,N_2617);
or U3146 (N_3146,N_2342,N_2834);
and U3147 (N_3147,N_2763,N_2710);
or U3148 (N_3148,N_2579,N_2519);
xor U3149 (N_3149,N_2533,N_2573);
or U3150 (N_3150,N_2944,N_2305);
nand U3151 (N_3151,N_2951,N_2319);
xnor U3152 (N_3152,N_2649,N_2306);
and U3153 (N_3153,N_2891,N_2415);
and U3154 (N_3154,N_2861,N_2735);
xnor U3155 (N_3155,N_2696,N_2414);
xor U3156 (N_3156,N_2480,N_2295);
nor U3157 (N_3157,N_2865,N_2998);
or U3158 (N_3158,N_2553,N_2945);
or U3159 (N_3159,N_2484,N_2557);
xor U3160 (N_3160,N_2437,N_2505);
xnor U3161 (N_3161,N_2536,N_2373);
or U3162 (N_3162,N_2826,N_2792);
nor U3163 (N_3163,N_2913,N_2364);
nand U3164 (N_3164,N_2597,N_2986);
and U3165 (N_3165,N_2399,N_2731);
or U3166 (N_3166,N_2911,N_2896);
or U3167 (N_3167,N_2524,N_2326);
or U3168 (N_3168,N_2332,N_2968);
nand U3169 (N_3169,N_2853,N_2377);
and U3170 (N_3170,N_2387,N_2594);
and U3171 (N_3171,N_2527,N_2670);
or U3172 (N_3172,N_2263,N_2408);
nand U3173 (N_3173,N_2636,N_2925);
or U3174 (N_3174,N_2516,N_2354);
or U3175 (N_3175,N_2786,N_2961);
nand U3176 (N_3176,N_2528,N_2331);
xnor U3177 (N_3177,N_2386,N_2948);
and U3178 (N_3178,N_2727,N_2370);
xnor U3179 (N_3179,N_2651,N_2932);
xor U3180 (N_3180,N_2931,N_2340);
xor U3181 (N_3181,N_2639,N_2790);
nor U3182 (N_3182,N_2880,N_2750);
xor U3183 (N_3183,N_2462,N_2448);
nor U3184 (N_3184,N_2800,N_2546);
and U3185 (N_3185,N_2828,N_2496);
nor U3186 (N_3186,N_2353,N_2837);
nand U3187 (N_3187,N_2667,N_2262);
or U3188 (N_3188,N_2378,N_2619);
or U3189 (N_3189,N_2762,N_2442);
nor U3190 (N_3190,N_2881,N_2752);
or U3191 (N_3191,N_2532,N_2930);
and U3192 (N_3192,N_2659,N_2506);
xor U3193 (N_3193,N_2281,N_2693);
nor U3194 (N_3194,N_2957,N_2473);
nand U3195 (N_3195,N_2877,N_2967);
and U3196 (N_3196,N_2607,N_2304);
or U3197 (N_3197,N_2385,N_2421);
and U3198 (N_3198,N_2920,N_2862);
xnor U3199 (N_3199,N_2491,N_2656);
nand U3200 (N_3200,N_2420,N_2526);
xnor U3201 (N_3201,N_2765,N_2798);
nor U3202 (N_3202,N_2695,N_2333);
and U3203 (N_3203,N_2795,N_2575);
nor U3204 (N_3204,N_2398,N_2647);
xor U3205 (N_3205,N_2394,N_2899);
xnor U3206 (N_3206,N_2601,N_2885);
nor U3207 (N_3207,N_2350,N_2668);
nor U3208 (N_3208,N_2301,N_2444);
or U3209 (N_3209,N_2269,N_2796);
and U3210 (N_3210,N_2732,N_2676);
and U3211 (N_3211,N_2641,N_2611);
nand U3212 (N_3212,N_2823,N_2588);
or U3213 (N_3213,N_2848,N_2477);
and U3214 (N_3214,N_2625,N_2938);
nor U3215 (N_3215,N_2251,N_2614);
xor U3216 (N_3216,N_2822,N_2872);
nor U3217 (N_3217,N_2905,N_2410);
nor U3218 (N_3218,N_2854,N_2388);
nor U3219 (N_3219,N_2325,N_2381);
nor U3220 (N_3220,N_2469,N_2874);
nor U3221 (N_3221,N_2927,N_2914);
or U3222 (N_3222,N_2719,N_2558);
and U3223 (N_3223,N_2784,N_2478);
xnor U3224 (N_3224,N_2981,N_2344);
nand U3225 (N_3225,N_2438,N_2852);
or U3226 (N_3226,N_2831,N_2851);
nor U3227 (N_3227,N_2422,N_2443);
nor U3228 (N_3228,N_2990,N_2253);
nand U3229 (N_3229,N_2453,N_2906);
or U3230 (N_3230,N_2298,N_2844);
and U3231 (N_3231,N_2503,N_2775);
or U3232 (N_3232,N_2684,N_2624);
and U3233 (N_3233,N_2963,N_2379);
or U3234 (N_3234,N_2329,N_2815);
nand U3235 (N_3235,N_2665,N_2451);
nor U3236 (N_3236,N_2833,N_2531);
xor U3237 (N_3237,N_2577,N_2278);
xnor U3238 (N_3238,N_2929,N_2372);
xnor U3239 (N_3239,N_2552,N_2487);
xnor U3240 (N_3240,N_2459,N_2427);
and U3241 (N_3241,N_2970,N_2979);
and U3242 (N_3242,N_2461,N_2894);
nand U3243 (N_3243,N_2666,N_2433);
nor U3244 (N_3244,N_2488,N_2652);
or U3245 (N_3245,N_2707,N_2768);
nor U3246 (N_3246,N_2813,N_2406);
or U3247 (N_3247,N_2382,N_2366);
or U3248 (N_3248,N_2717,N_2835);
or U3249 (N_3249,N_2791,N_2454);
nand U3250 (N_3250,N_2347,N_2284);
xnor U3251 (N_3251,N_2838,N_2606);
xor U3252 (N_3252,N_2976,N_2456);
nand U3253 (N_3253,N_2702,N_2926);
nor U3254 (N_3254,N_2730,N_2542);
xnor U3255 (N_3255,N_2644,N_2890);
xnor U3256 (N_3256,N_2738,N_2917);
nand U3257 (N_3257,N_2962,N_2691);
and U3258 (N_3258,N_2952,N_2632);
nor U3259 (N_3259,N_2513,N_2878);
xnor U3260 (N_3260,N_2904,N_2518);
nor U3261 (N_3261,N_2336,N_2989);
and U3262 (N_3262,N_2323,N_2673);
nor U3263 (N_3263,N_2770,N_2481);
and U3264 (N_3264,N_2609,N_2302);
and U3265 (N_3265,N_2871,N_2276);
nand U3266 (N_3266,N_2711,N_2435);
and U3267 (N_3267,N_2521,N_2508);
nand U3268 (N_3268,N_2417,N_2724);
nand U3269 (N_3269,N_2734,N_2940);
or U3270 (N_3270,N_2428,N_2759);
and U3271 (N_3271,N_2842,N_2598);
and U3272 (N_3272,N_2574,N_2672);
or U3273 (N_3273,N_2474,N_2627);
nand U3274 (N_3274,N_2403,N_2593);
nor U3275 (N_3275,N_2529,N_2458);
and U3276 (N_3276,N_2283,N_2887);
or U3277 (N_3277,N_2956,N_2494);
and U3278 (N_3278,N_2360,N_2722);
xnor U3279 (N_3279,N_2642,N_2507);
nor U3280 (N_3280,N_2969,N_2595);
and U3281 (N_3281,N_2638,N_2824);
or U3282 (N_3282,N_2273,N_2825);
nand U3283 (N_3283,N_2657,N_2475);
or U3284 (N_3284,N_2805,N_2782);
and U3285 (N_3285,N_2447,N_2610);
nand U3286 (N_3286,N_2803,N_2832);
and U3287 (N_3287,N_2715,N_2375);
xor U3288 (N_3288,N_2275,N_2996);
xnor U3289 (N_3289,N_2365,N_2600);
or U3290 (N_3290,N_2497,N_2502);
or U3291 (N_3291,N_2708,N_2434);
or U3292 (N_3292,N_2512,N_2766);
xnor U3293 (N_3293,N_2748,N_2522);
xor U3294 (N_3294,N_2631,N_2820);
or U3295 (N_3295,N_2316,N_2997);
nor U3296 (N_3296,N_2787,N_2973);
or U3297 (N_3297,N_2586,N_2402);
and U3298 (N_3298,N_2358,N_2580);
nor U3299 (N_3299,N_2939,N_2958);
nor U3300 (N_3300,N_2424,N_2858);
and U3301 (N_3301,N_2544,N_2836);
xnor U3302 (N_3302,N_2648,N_2486);
or U3303 (N_3303,N_2547,N_2346);
nand U3304 (N_3304,N_2714,N_2623);
xnor U3305 (N_3305,N_2819,N_2797);
nand U3306 (N_3306,N_2746,N_2500);
xor U3307 (N_3307,N_2412,N_2776);
nor U3308 (N_3308,N_2814,N_2287);
nor U3309 (N_3309,N_2498,N_2999);
and U3310 (N_3310,N_2268,N_2534);
or U3311 (N_3311,N_2425,N_2274);
or U3312 (N_3312,N_2856,N_2482);
nor U3313 (N_3313,N_2297,N_2440);
and U3314 (N_3314,N_2818,N_2545);
xnor U3315 (N_3315,N_2661,N_2689);
nand U3316 (N_3316,N_2895,N_2882);
xnor U3317 (N_3317,N_2439,N_2669);
or U3318 (N_3318,N_2897,N_2327);
nor U3319 (N_3319,N_2261,N_2811);
and U3320 (N_3320,N_2615,N_2781);
or U3321 (N_3321,N_2525,N_2723);
nor U3322 (N_3322,N_2339,N_2821);
nor U3323 (N_3323,N_2395,N_2310);
and U3324 (N_3324,N_2690,N_2318);
nand U3325 (N_3325,N_2985,N_2662);
xnor U3326 (N_3326,N_2995,N_2915);
or U3327 (N_3327,N_2539,N_2554);
and U3328 (N_3328,N_2250,N_2277);
or U3329 (N_3329,N_2947,N_2567);
nor U3330 (N_3330,N_2300,N_2771);
nor U3331 (N_3331,N_2898,N_2937);
and U3332 (N_3332,N_2455,N_2312);
and U3333 (N_3333,N_2694,N_2830);
or U3334 (N_3334,N_2343,N_2699);
and U3335 (N_3335,N_2867,N_2873);
xnor U3336 (N_3336,N_2452,N_2510);
nand U3337 (N_3337,N_2789,N_2559);
nor U3338 (N_3338,N_2270,N_2712);
xnor U3339 (N_3339,N_2953,N_2655);
and U3340 (N_3340,N_2807,N_2866);
or U3341 (N_3341,N_2293,N_2584);
nand U3342 (N_3342,N_2941,N_2308);
nand U3343 (N_3343,N_2613,N_2928);
nor U3344 (N_3344,N_2530,N_2596);
and U3345 (N_3345,N_2658,N_2946);
nand U3346 (N_3346,N_2432,N_2561);
nand U3347 (N_3347,N_2368,N_2760);
and U3348 (N_3348,N_2754,N_2548);
xnor U3349 (N_3349,N_2272,N_2591);
or U3350 (N_3350,N_2501,N_2769);
and U3351 (N_3351,N_2869,N_2685);
or U3352 (N_3352,N_2471,N_2745);
xnor U3353 (N_3353,N_2704,N_2369);
and U3354 (N_3354,N_2282,N_2401);
nor U3355 (N_3355,N_2384,N_2692);
and U3356 (N_3356,N_2313,N_2964);
nor U3357 (N_3357,N_2311,N_2572);
nor U3358 (N_3358,N_2464,N_2315);
xor U3359 (N_3359,N_2777,N_2840);
and U3360 (N_3360,N_2254,N_2514);
nor U3361 (N_3361,N_2788,N_2855);
nor U3362 (N_3362,N_2804,N_2380);
and U3363 (N_3363,N_2449,N_2404);
or U3364 (N_3364,N_2700,N_2859);
nor U3365 (N_3365,N_2290,N_2705);
or U3366 (N_3366,N_2470,N_2982);
or U3367 (N_3367,N_2955,N_2556);
nand U3368 (N_3368,N_2774,N_2767);
nand U3369 (N_3369,N_2740,N_2551);
nor U3370 (N_3370,N_2618,N_2289);
and U3371 (N_3371,N_2396,N_2334);
xnor U3372 (N_3372,N_2713,N_2809);
or U3373 (N_3373,N_2581,N_2603);
xnor U3374 (N_3374,N_2257,N_2875);
or U3375 (N_3375,N_2378,N_2638);
or U3376 (N_3376,N_2560,N_2528);
and U3377 (N_3377,N_2853,N_2485);
nand U3378 (N_3378,N_2779,N_2661);
xnor U3379 (N_3379,N_2796,N_2475);
or U3380 (N_3380,N_2922,N_2936);
and U3381 (N_3381,N_2771,N_2673);
xnor U3382 (N_3382,N_2361,N_2558);
nand U3383 (N_3383,N_2416,N_2341);
nor U3384 (N_3384,N_2815,N_2891);
or U3385 (N_3385,N_2903,N_2264);
nor U3386 (N_3386,N_2966,N_2382);
nand U3387 (N_3387,N_2496,N_2996);
and U3388 (N_3388,N_2939,N_2486);
nand U3389 (N_3389,N_2612,N_2955);
nor U3390 (N_3390,N_2819,N_2959);
nor U3391 (N_3391,N_2398,N_2910);
and U3392 (N_3392,N_2686,N_2457);
xnor U3393 (N_3393,N_2328,N_2978);
nor U3394 (N_3394,N_2947,N_2974);
and U3395 (N_3395,N_2667,N_2757);
or U3396 (N_3396,N_2399,N_2752);
and U3397 (N_3397,N_2464,N_2952);
and U3398 (N_3398,N_2577,N_2906);
and U3399 (N_3399,N_2543,N_2821);
nand U3400 (N_3400,N_2718,N_2392);
nand U3401 (N_3401,N_2417,N_2503);
xnor U3402 (N_3402,N_2540,N_2883);
or U3403 (N_3403,N_2473,N_2426);
nand U3404 (N_3404,N_2435,N_2350);
xnor U3405 (N_3405,N_2386,N_2849);
and U3406 (N_3406,N_2510,N_2976);
nor U3407 (N_3407,N_2396,N_2583);
nor U3408 (N_3408,N_2736,N_2495);
nand U3409 (N_3409,N_2417,N_2693);
nor U3410 (N_3410,N_2972,N_2688);
nor U3411 (N_3411,N_2492,N_2450);
nand U3412 (N_3412,N_2815,N_2965);
nand U3413 (N_3413,N_2575,N_2955);
nor U3414 (N_3414,N_2518,N_2690);
xnor U3415 (N_3415,N_2685,N_2495);
xor U3416 (N_3416,N_2970,N_2623);
and U3417 (N_3417,N_2885,N_2358);
or U3418 (N_3418,N_2322,N_2991);
nor U3419 (N_3419,N_2320,N_2820);
nand U3420 (N_3420,N_2640,N_2361);
or U3421 (N_3421,N_2999,N_2851);
nand U3422 (N_3422,N_2702,N_2255);
nor U3423 (N_3423,N_2837,N_2736);
xnor U3424 (N_3424,N_2333,N_2753);
or U3425 (N_3425,N_2677,N_2678);
xor U3426 (N_3426,N_2648,N_2332);
xnor U3427 (N_3427,N_2264,N_2390);
nand U3428 (N_3428,N_2647,N_2822);
and U3429 (N_3429,N_2874,N_2994);
and U3430 (N_3430,N_2978,N_2579);
and U3431 (N_3431,N_2492,N_2628);
nand U3432 (N_3432,N_2912,N_2527);
nand U3433 (N_3433,N_2574,N_2505);
nand U3434 (N_3434,N_2381,N_2985);
nand U3435 (N_3435,N_2922,N_2346);
xor U3436 (N_3436,N_2258,N_2553);
xor U3437 (N_3437,N_2947,N_2451);
or U3438 (N_3438,N_2540,N_2890);
nor U3439 (N_3439,N_2921,N_2267);
nand U3440 (N_3440,N_2740,N_2450);
and U3441 (N_3441,N_2255,N_2647);
or U3442 (N_3442,N_2334,N_2613);
xor U3443 (N_3443,N_2677,N_2338);
nand U3444 (N_3444,N_2447,N_2560);
xor U3445 (N_3445,N_2937,N_2457);
xnor U3446 (N_3446,N_2462,N_2626);
and U3447 (N_3447,N_2882,N_2284);
nor U3448 (N_3448,N_2825,N_2795);
and U3449 (N_3449,N_2486,N_2385);
nand U3450 (N_3450,N_2294,N_2517);
nand U3451 (N_3451,N_2921,N_2735);
or U3452 (N_3452,N_2592,N_2529);
and U3453 (N_3453,N_2955,N_2718);
xnor U3454 (N_3454,N_2843,N_2453);
nor U3455 (N_3455,N_2597,N_2785);
nand U3456 (N_3456,N_2846,N_2636);
nand U3457 (N_3457,N_2270,N_2797);
or U3458 (N_3458,N_2962,N_2568);
nand U3459 (N_3459,N_2315,N_2588);
or U3460 (N_3460,N_2802,N_2923);
and U3461 (N_3461,N_2459,N_2520);
or U3462 (N_3462,N_2377,N_2367);
and U3463 (N_3463,N_2957,N_2894);
and U3464 (N_3464,N_2687,N_2667);
nor U3465 (N_3465,N_2751,N_2724);
and U3466 (N_3466,N_2735,N_2972);
and U3467 (N_3467,N_2915,N_2536);
nor U3468 (N_3468,N_2964,N_2477);
nor U3469 (N_3469,N_2341,N_2769);
nand U3470 (N_3470,N_2443,N_2947);
nor U3471 (N_3471,N_2802,N_2349);
and U3472 (N_3472,N_2653,N_2959);
nand U3473 (N_3473,N_2332,N_2616);
and U3474 (N_3474,N_2657,N_2406);
and U3475 (N_3475,N_2336,N_2631);
nor U3476 (N_3476,N_2971,N_2985);
nor U3477 (N_3477,N_2329,N_2289);
nand U3478 (N_3478,N_2650,N_2555);
nand U3479 (N_3479,N_2891,N_2325);
xnor U3480 (N_3480,N_2860,N_2659);
xor U3481 (N_3481,N_2688,N_2927);
and U3482 (N_3482,N_2380,N_2717);
and U3483 (N_3483,N_2983,N_2855);
nand U3484 (N_3484,N_2928,N_2333);
or U3485 (N_3485,N_2917,N_2711);
and U3486 (N_3486,N_2724,N_2611);
nor U3487 (N_3487,N_2491,N_2611);
nor U3488 (N_3488,N_2639,N_2316);
nor U3489 (N_3489,N_2803,N_2497);
and U3490 (N_3490,N_2488,N_2741);
nor U3491 (N_3491,N_2984,N_2682);
nor U3492 (N_3492,N_2261,N_2981);
xor U3493 (N_3493,N_2832,N_2427);
nand U3494 (N_3494,N_2396,N_2451);
nor U3495 (N_3495,N_2577,N_2809);
and U3496 (N_3496,N_2474,N_2272);
nand U3497 (N_3497,N_2733,N_2584);
and U3498 (N_3498,N_2767,N_2606);
xnor U3499 (N_3499,N_2420,N_2974);
xnor U3500 (N_3500,N_2513,N_2891);
nand U3501 (N_3501,N_2474,N_2808);
or U3502 (N_3502,N_2568,N_2702);
and U3503 (N_3503,N_2627,N_2775);
xor U3504 (N_3504,N_2466,N_2833);
nand U3505 (N_3505,N_2474,N_2390);
nor U3506 (N_3506,N_2441,N_2588);
nor U3507 (N_3507,N_2339,N_2363);
nor U3508 (N_3508,N_2383,N_2518);
or U3509 (N_3509,N_2273,N_2549);
xor U3510 (N_3510,N_2945,N_2848);
nor U3511 (N_3511,N_2656,N_2717);
nor U3512 (N_3512,N_2801,N_2290);
nor U3513 (N_3513,N_2635,N_2493);
nand U3514 (N_3514,N_2482,N_2853);
xnor U3515 (N_3515,N_2492,N_2899);
xnor U3516 (N_3516,N_2980,N_2367);
and U3517 (N_3517,N_2467,N_2348);
xor U3518 (N_3518,N_2973,N_2455);
and U3519 (N_3519,N_2280,N_2911);
xnor U3520 (N_3520,N_2611,N_2806);
or U3521 (N_3521,N_2332,N_2821);
xor U3522 (N_3522,N_2274,N_2353);
xnor U3523 (N_3523,N_2836,N_2488);
and U3524 (N_3524,N_2964,N_2390);
xnor U3525 (N_3525,N_2957,N_2497);
and U3526 (N_3526,N_2681,N_2411);
nand U3527 (N_3527,N_2686,N_2805);
nor U3528 (N_3528,N_2421,N_2558);
xnor U3529 (N_3529,N_2731,N_2586);
nand U3530 (N_3530,N_2847,N_2645);
nand U3531 (N_3531,N_2258,N_2252);
and U3532 (N_3532,N_2641,N_2557);
and U3533 (N_3533,N_2374,N_2313);
and U3534 (N_3534,N_2649,N_2322);
and U3535 (N_3535,N_2552,N_2877);
or U3536 (N_3536,N_2774,N_2388);
nor U3537 (N_3537,N_2845,N_2318);
nand U3538 (N_3538,N_2448,N_2771);
xnor U3539 (N_3539,N_2918,N_2621);
or U3540 (N_3540,N_2301,N_2393);
nor U3541 (N_3541,N_2802,N_2707);
nand U3542 (N_3542,N_2316,N_2269);
or U3543 (N_3543,N_2544,N_2944);
xor U3544 (N_3544,N_2870,N_2399);
and U3545 (N_3545,N_2490,N_2395);
nor U3546 (N_3546,N_2632,N_2902);
nand U3547 (N_3547,N_2567,N_2440);
nand U3548 (N_3548,N_2529,N_2853);
and U3549 (N_3549,N_2658,N_2538);
and U3550 (N_3550,N_2311,N_2394);
and U3551 (N_3551,N_2271,N_2270);
nand U3552 (N_3552,N_2419,N_2961);
or U3553 (N_3553,N_2688,N_2595);
or U3554 (N_3554,N_2974,N_2364);
nand U3555 (N_3555,N_2921,N_2606);
xnor U3556 (N_3556,N_2844,N_2451);
nor U3557 (N_3557,N_2994,N_2955);
xor U3558 (N_3558,N_2810,N_2695);
or U3559 (N_3559,N_2700,N_2784);
nand U3560 (N_3560,N_2532,N_2553);
and U3561 (N_3561,N_2320,N_2800);
nor U3562 (N_3562,N_2667,N_2473);
nand U3563 (N_3563,N_2823,N_2261);
and U3564 (N_3564,N_2718,N_2847);
xor U3565 (N_3565,N_2542,N_2922);
or U3566 (N_3566,N_2837,N_2317);
and U3567 (N_3567,N_2373,N_2364);
nor U3568 (N_3568,N_2274,N_2900);
nor U3569 (N_3569,N_2541,N_2257);
or U3570 (N_3570,N_2806,N_2311);
xor U3571 (N_3571,N_2876,N_2860);
xnor U3572 (N_3572,N_2907,N_2628);
nand U3573 (N_3573,N_2921,N_2996);
or U3574 (N_3574,N_2491,N_2989);
or U3575 (N_3575,N_2652,N_2268);
xnor U3576 (N_3576,N_2358,N_2318);
and U3577 (N_3577,N_2559,N_2854);
nand U3578 (N_3578,N_2595,N_2827);
xnor U3579 (N_3579,N_2420,N_2580);
nand U3580 (N_3580,N_2845,N_2951);
nand U3581 (N_3581,N_2719,N_2572);
nor U3582 (N_3582,N_2789,N_2409);
xnor U3583 (N_3583,N_2318,N_2755);
xor U3584 (N_3584,N_2454,N_2719);
nor U3585 (N_3585,N_2846,N_2506);
or U3586 (N_3586,N_2723,N_2788);
or U3587 (N_3587,N_2348,N_2668);
or U3588 (N_3588,N_2390,N_2552);
nor U3589 (N_3589,N_2784,N_2680);
or U3590 (N_3590,N_2449,N_2975);
nand U3591 (N_3591,N_2496,N_2978);
nor U3592 (N_3592,N_2935,N_2587);
nor U3593 (N_3593,N_2356,N_2990);
or U3594 (N_3594,N_2910,N_2708);
xor U3595 (N_3595,N_2658,N_2847);
and U3596 (N_3596,N_2371,N_2367);
nand U3597 (N_3597,N_2439,N_2591);
or U3598 (N_3598,N_2849,N_2702);
nor U3599 (N_3599,N_2652,N_2346);
nand U3600 (N_3600,N_2335,N_2516);
nand U3601 (N_3601,N_2635,N_2945);
and U3602 (N_3602,N_2250,N_2649);
xnor U3603 (N_3603,N_2632,N_2844);
nor U3604 (N_3604,N_2507,N_2589);
and U3605 (N_3605,N_2671,N_2992);
nand U3606 (N_3606,N_2989,N_2579);
and U3607 (N_3607,N_2515,N_2405);
nand U3608 (N_3608,N_2750,N_2863);
and U3609 (N_3609,N_2708,N_2510);
or U3610 (N_3610,N_2611,N_2686);
and U3611 (N_3611,N_2579,N_2369);
xnor U3612 (N_3612,N_2758,N_2928);
nand U3613 (N_3613,N_2496,N_2809);
nand U3614 (N_3614,N_2874,N_2997);
xnor U3615 (N_3615,N_2439,N_2837);
xor U3616 (N_3616,N_2785,N_2598);
nand U3617 (N_3617,N_2989,N_2828);
nand U3618 (N_3618,N_2691,N_2772);
nor U3619 (N_3619,N_2902,N_2336);
xor U3620 (N_3620,N_2429,N_2265);
and U3621 (N_3621,N_2904,N_2507);
xor U3622 (N_3622,N_2920,N_2457);
or U3623 (N_3623,N_2375,N_2654);
nand U3624 (N_3624,N_2366,N_2643);
or U3625 (N_3625,N_2606,N_2871);
nand U3626 (N_3626,N_2394,N_2637);
xnor U3627 (N_3627,N_2403,N_2352);
or U3628 (N_3628,N_2589,N_2906);
and U3629 (N_3629,N_2554,N_2846);
and U3630 (N_3630,N_2952,N_2440);
and U3631 (N_3631,N_2446,N_2447);
nand U3632 (N_3632,N_2998,N_2508);
or U3633 (N_3633,N_2536,N_2749);
nand U3634 (N_3634,N_2965,N_2707);
or U3635 (N_3635,N_2257,N_2727);
nor U3636 (N_3636,N_2344,N_2875);
or U3637 (N_3637,N_2437,N_2837);
or U3638 (N_3638,N_2388,N_2968);
or U3639 (N_3639,N_2493,N_2597);
xnor U3640 (N_3640,N_2703,N_2952);
nor U3641 (N_3641,N_2393,N_2650);
nor U3642 (N_3642,N_2423,N_2946);
nand U3643 (N_3643,N_2804,N_2399);
xor U3644 (N_3644,N_2545,N_2341);
xnor U3645 (N_3645,N_2541,N_2816);
and U3646 (N_3646,N_2863,N_2646);
xor U3647 (N_3647,N_2805,N_2842);
xnor U3648 (N_3648,N_2421,N_2440);
xor U3649 (N_3649,N_2283,N_2960);
and U3650 (N_3650,N_2884,N_2832);
nand U3651 (N_3651,N_2884,N_2703);
or U3652 (N_3652,N_2508,N_2600);
or U3653 (N_3653,N_2807,N_2382);
xnor U3654 (N_3654,N_2804,N_2805);
or U3655 (N_3655,N_2868,N_2577);
and U3656 (N_3656,N_2285,N_2821);
nand U3657 (N_3657,N_2766,N_2787);
and U3658 (N_3658,N_2771,N_2919);
and U3659 (N_3659,N_2828,N_2252);
or U3660 (N_3660,N_2498,N_2379);
or U3661 (N_3661,N_2304,N_2700);
and U3662 (N_3662,N_2732,N_2914);
nand U3663 (N_3663,N_2480,N_2894);
nand U3664 (N_3664,N_2798,N_2502);
or U3665 (N_3665,N_2901,N_2348);
or U3666 (N_3666,N_2583,N_2371);
nand U3667 (N_3667,N_2369,N_2446);
or U3668 (N_3668,N_2597,N_2480);
and U3669 (N_3669,N_2432,N_2406);
or U3670 (N_3670,N_2585,N_2370);
xor U3671 (N_3671,N_2615,N_2538);
nand U3672 (N_3672,N_2384,N_2424);
xor U3673 (N_3673,N_2339,N_2593);
or U3674 (N_3674,N_2987,N_2420);
xnor U3675 (N_3675,N_2377,N_2978);
nor U3676 (N_3676,N_2499,N_2956);
and U3677 (N_3677,N_2402,N_2763);
or U3678 (N_3678,N_2741,N_2552);
and U3679 (N_3679,N_2815,N_2334);
nand U3680 (N_3680,N_2739,N_2501);
or U3681 (N_3681,N_2822,N_2755);
nor U3682 (N_3682,N_2873,N_2868);
nor U3683 (N_3683,N_2259,N_2957);
nand U3684 (N_3684,N_2979,N_2738);
or U3685 (N_3685,N_2588,N_2569);
nand U3686 (N_3686,N_2953,N_2418);
and U3687 (N_3687,N_2833,N_2870);
and U3688 (N_3688,N_2591,N_2385);
nand U3689 (N_3689,N_2471,N_2526);
and U3690 (N_3690,N_2924,N_2768);
xnor U3691 (N_3691,N_2700,N_2984);
xor U3692 (N_3692,N_2275,N_2844);
xnor U3693 (N_3693,N_2735,N_2483);
xor U3694 (N_3694,N_2624,N_2746);
or U3695 (N_3695,N_2616,N_2451);
nand U3696 (N_3696,N_2956,N_2798);
or U3697 (N_3697,N_2698,N_2609);
xnor U3698 (N_3698,N_2749,N_2903);
xor U3699 (N_3699,N_2293,N_2316);
or U3700 (N_3700,N_2708,N_2884);
and U3701 (N_3701,N_2969,N_2327);
or U3702 (N_3702,N_2452,N_2301);
and U3703 (N_3703,N_2469,N_2388);
nor U3704 (N_3704,N_2334,N_2579);
or U3705 (N_3705,N_2316,N_2511);
and U3706 (N_3706,N_2971,N_2327);
nor U3707 (N_3707,N_2717,N_2497);
xnor U3708 (N_3708,N_2704,N_2761);
or U3709 (N_3709,N_2917,N_2670);
nor U3710 (N_3710,N_2344,N_2596);
xor U3711 (N_3711,N_2810,N_2702);
xnor U3712 (N_3712,N_2525,N_2427);
nand U3713 (N_3713,N_2885,N_2329);
nor U3714 (N_3714,N_2428,N_2332);
nand U3715 (N_3715,N_2768,N_2939);
xor U3716 (N_3716,N_2401,N_2637);
nand U3717 (N_3717,N_2268,N_2455);
xnor U3718 (N_3718,N_2266,N_2838);
or U3719 (N_3719,N_2777,N_2985);
nand U3720 (N_3720,N_2887,N_2273);
nor U3721 (N_3721,N_2950,N_2665);
nand U3722 (N_3722,N_2880,N_2416);
or U3723 (N_3723,N_2648,N_2527);
nor U3724 (N_3724,N_2926,N_2285);
or U3725 (N_3725,N_2321,N_2456);
nand U3726 (N_3726,N_2744,N_2490);
nor U3727 (N_3727,N_2605,N_2584);
nor U3728 (N_3728,N_2962,N_2339);
nand U3729 (N_3729,N_2987,N_2876);
nor U3730 (N_3730,N_2438,N_2405);
nor U3731 (N_3731,N_2455,N_2866);
and U3732 (N_3732,N_2586,N_2758);
nand U3733 (N_3733,N_2454,N_2865);
and U3734 (N_3734,N_2398,N_2620);
nand U3735 (N_3735,N_2802,N_2326);
or U3736 (N_3736,N_2846,N_2610);
nor U3737 (N_3737,N_2803,N_2805);
nand U3738 (N_3738,N_2492,N_2300);
nor U3739 (N_3739,N_2811,N_2292);
and U3740 (N_3740,N_2439,N_2551);
or U3741 (N_3741,N_2389,N_2542);
and U3742 (N_3742,N_2944,N_2334);
xor U3743 (N_3743,N_2411,N_2806);
xnor U3744 (N_3744,N_2444,N_2422);
or U3745 (N_3745,N_2861,N_2516);
nor U3746 (N_3746,N_2866,N_2662);
nor U3747 (N_3747,N_2425,N_2633);
nand U3748 (N_3748,N_2951,N_2978);
nor U3749 (N_3749,N_2764,N_2739);
or U3750 (N_3750,N_3447,N_3280);
nand U3751 (N_3751,N_3133,N_3442);
nor U3752 (N_3752,N_3388,N_3046);
and U3753 (N_3753,N_3591,N_3015);
or U3754 (N_3754,N_3535,N_3078);
nand U3755 (N_3755,N_3251,N_3739);
or U3756 (N_3756,N_3153,N_3742);
nor U3757 (N_3757,N_3741,N_3166);
nor U3758 (N_3758,N_3463,N_3571);
nor U3759 (N_3759,N_3714,N_3381);
xor U3760 (N_3760,N_3365,N_3728);
or U3761 (N_3761,N_3171,N_3000);
and U3762 (N_3762,N_3725,N_3623);
or U3763 (N_3763,N_3149,N_3680);
or U3764 (N_3764,N_3111,N_3290);
and U3765 (N_3765,N_3504,N_3256);
or U3766 (N_3766,N_3513,N_3259);
nor U3767 (N_3767,N_3386,N_3407);
or U3768 (N_3768,N_3083,N_3658);
xor U3769 (N_3769,N_3131,N_3268);
or U3770 (N_3770,N_3743,N_3610);
xor U3771 (N_3771,N_3126,N_3669);
nor U3772 (N_3772,N_3690,N_3635);
xnor U3773 (N_3773,N_3347,N_3211);
nor U3774 (N_3774,N_3248,N_3484);
or U3775 (N_3775,N_3552,N_3210);
nand U3776 (N_3776,N_3238,N_3048);
or U3777 (N_3777,N_3029,N_3032);
nor U3778 (N_3778,N_3637,N_3607);
nor U3779 (N_3779,N_3409,N_3295);
and U3780 (N_3780,N_3345,N_3119);
xor U3781 (N_3781,N_3713,N_3632);
or U3782 (N_3782,N_3720,N_3021);
or U3783 (N_3783,N_3639,N_3622);
and U3784 (N_3784,N_3410,N_3529);
and U3785 (N_3785,N_3218,N_3660);
and U3786 (N_3786,N_3574,N_3336);
and U3787 (N_3787,N_3170,N_3246);
or U3788 (N_3788,N_3547,N_3693);
nor U3789 (N_3789,N_3045,N_3228);
nand U3790 (N_3790,N_3040,N_3652);
nand U3791 (N_3791,N_3321,N_3364);
nor U3792 (N_3792,N_3105,N_3575);
nand U3793 (N_3793,N_3314,N_3152);
xnor U3794 (N_3794,N_3282,N_3479);
or U3795 (N_3795,N_3310,N_3666);
and U3796 (N_3796,N_3617,N_3727);
nor U3797 (N_3797,N_3262,N_3281);
nand U3798 (N_3798,N_3272,N_3536);
xnor U3799 (N_3799,N_3223,N_3208);
nand U3800 (N_3800,N_3236,N_3107);
and U3801 (N_3801,N_3049,N_3512);
and U3802 (N_3802,N_3118,N_3435);
nor U3803 (N_3803,N_3627,N_3446);
nor U3804 (N_3804,N_3288,N_3201);
or U3805 (N_3805,N_3071,N_3539);
or U3806 (N_3806,N_3052,N_3556);
nor U3807 (N_3807,N_3304,N_3412);
or U3808 (N_3808,N_3294,N_3163);
nor U3809 (N_3809,N_3235,N_3222);
nor U3810 (N_3810,N_3239,N_3139);
nor U3811 (N_3811,N_3475,N_3459);
xor U3812 (N_3812,N_3359,N_3630);
xor U3813 (N_3813,N_3101,N_3028);
xor U3814 (N_3814,N_3698,N_3317);
xor U3815 (N_3815,N_3613,N_3424);
or U3816 (N_3816,N_3538,N_3415);
nor U3817 (N_3817,N_3073,N_3093);
nor U3818 (N_3818,N_3564,N_3716);
nor U3819 (N_3819,N_3241,N_3494);
xor U3820 (N_3820,N_3379,N_3668);
nor U3821 (N_3821,N_3136,N_3501);
and U3822 (N_3822,N_3144,N_3180);
nand U3823 (N_3823,N_3206,N_3108);
nand U3824 (N_3824,N_3450,N_3335);
xnor U3825 (N_3825,N_3638,N_3156);
xor U3826 (N_3826,N_3188,N_3159);
xor U3827 (N_3827,N_3700,N_3319);
or U3828 (N_3828,N_3011,N_3005);
nor U3829 (N_3829,N_3151,N_3220);
nor U3830 (N_3830,N_3506,N_3115);
and U3831 (N_3831,N_3723,N_3296);
nor U3832 (N_3832,N_3326,N_3567);
nand U3833 (N_3833,N_3470,N_3129);
and U3834 (N_3834,N_3654,N_3064);
nand U3835 (N_3835,N_3313,N_3746);
xnor U3836 (N_3836,N_3192,N_3438);
nor U3837 (N_3837,N_3219,N_3275);
nand U3838 (N_3838,N_3573,N_3657);
xor U3839 (N_3839,N_3089,N_3642);
or U3840 (N_3840,N_3342,N_3453);
nor U3841 (N_3841,N_3305,N_3621);
and U3842 (N_3842,N_3525,N_3189);
xor U3843 (N_3843,N_3341,N_3097);
nor U3844 (N_3844,N_3261,N_3351);
and U3845 (N_3845,N_3298,N_3245);
nor U3846 (N_3846,N_3508,N_3662);
and U3847 (N_3847,N_3320,N_3123);
nand U3848 (N_3848,N_3300,N_3618);
nand U3849 (N_3849,N_3626,N_3534);
nor U3850 (N_3850,N_3628,N_3130);
nor U3851 (N_3851,N_3356,N_3437);
or U3852 (N_3852,N_3191,N_3541);
nor U3853 (N_3853,N_3376,N_3323);
nor U3854 (N_3854,N_3114,N_3570);
nand U3855 (N_3855,N_3041,N_3517);
nand U3856 (N_3856,N_3127,N_3457);
or U3857 (N_3857,N_3650,N_3629);
nand U3858 (N_3858,N_3455,N_3599);
nor U3859 (N_3859,N_3577,N_3566);
and U3860 (N_3860,N_3675,N_3553);
xor U3861 (N_3861,N_3014,N_3242);
nor U3862 (N_3862,N_3497,N_3588);
nor U3863 (N_3863,N_3197,N_3380);
xor U3864 (N_3864,N_3518,N_3393);
and U3865 (N_3865,N_3193,N_3467);
nand U3866 (N_3866,N_3584,N_3592);
nand U3867 (N_3867,N_3024,N_3499);
or U3868 (N_3868,N_3250,N_3276);
nand U3869 (N_3869,N_3677,N_3413);
nand U3870 (N_3870,N_3003,N_3138);
xnor U3871 (N_3871,N_3075,N_3441);
nand U3872 (N_3872,N_3154,N_3181);
or U3873 (N_3873,N_3002,N_3354);
or U3874 (N_3874,N_3090,N_3587);
xnor U3875 (N_3875,N_3018,N_3312);
and U3876 (N_3876,N_3582,N_3614);
and U3877 (N_3877,N_3511,N_3664);
xnor U3878 (N_3878,N_3440,N_3589);
or U3879 (N_3879,N_3085,N_3478);
xnor U3880 (N_3880,N_3094,N_3301);
xnor U3881 (N_3881,N_3401,N_3168);
and U3882 (N_3882,N_3087,N_3733);
or U3883 (N_3883,N_3065,N_3325);
nor U3884 (N_3884,N_3340,N_3661);
nor U3885 (N_3885,N_3578,N_3480);
nand U3886 (N_3886,N_3327,N_3583);
and U3887 (N_3887,N_3425,N_3404);
nor U3888 (N_3888,N_3350,N_3397);
and U3889 (N_3889,N_3708,N_3370);
or U3890 (N_3890,N_3289,N_3432);
nor U3891 (N_3891,N_3489,N_3605);
or U3892 (N_3892,N_3234,N_3520);
nand U3893 (N_3893,N_3165,N_3526);
nor U3894 (N_3894,N_3546,N_3155);
and U3895 (N_3895,N_3540,N_3731);
xor U3896 (N_3896,N_3456,N_3515);
nand U3897 (N_3897,N_3744,N_3704);
nand U3898 (N_3898,N_3549,N_3291);
nor U3899 (N_3899,N_3496,N_3625);
xor U3900 (N_3900,N_3600,N_3034);
and U3901 (N_3901,N_3724,N_3711);
nor U3902 (N_3902,N_3244,N_3017);
nor U3903 (N_3903,N_3134,N_3231);
xor U3904 (N_3904,N_3299,N_3648);
nor U3905 (N_3905,N_3263,N_3581);
nor U3906 (N_3906,N_3178,N_3361);
nand U3907 (N_3907,N_3172,N_3167);
xnor U3908 (N_3908,N_3430,N_3682);
nor U3909 (N_3909,N_3287,N_3240);
nor U3910 (N_3910,N_3150,N_3400);
xor U3911 (N_3911,N_3633,N_3173);
xor U3912 (N_3912,N_3037,N_3355);
xor U3913 (N_3913,N_3729,N_3548);
or U3914 (N_3914,N_3604,N_3116);
nand U3915 (N_3915,N_3394,N_3174);
xnor U3916 (N_3916,N_3311,N_3203);
nand U3917 (N_3917,N_3684,N_3563);
and U3918 (N_3918,N_3196,N_3039);
nor U3919 (N_3919,N_3543,N_3025);
nor U3920 (N_3920,N_3302,N_3182);
xnor U3921 (N_3921,N_3745,N_3081);
nand U3922 (N_3922,N_3697,N_3416);
and U3923 (N_3923,N_3348,N_3187);
xor U3924 (N_3924,N_3466,N_3378);
and U3925 (N_3925,N_3473,N_3051);
nand U3926 (N_3926,N_3086,N_3308);
nand U3927 (N_3927,N_3636,N_3247);
or U3928 (N_3928,N_3500,N_3550);
or U3929 (N_3929,N_3195,N_3176);
nand U3930 (N_3930,N_3339,N_3158);
and U3931 (N_3931,N_3042,N_3503);
and U3932 (N_3932,N_3352,N_3418);
and U3933 (N_3933,N_3061,N_3420);
or U3934 (N_3934,N_3070,N_3221);
nand U3935 (N_3935,N_3277,N_3460);
and U3936 (N_3936,N_3224,N_3471);
xnor U3937 (N_3937,N_3316,N_3624);
nor U3938 (N_3938,N_3428,N_3530);
nor U3939 (N_3939,N_3569,N_3315);
nor U3940 (N_3940,N_3488,N_3260);
nor U3941 (N_3941,N_3738,N_3434);
nor U3942 (N_3942,N_3140,N_3072);
xor U3943 (N_3943,N_3491,N_3059);
nand U3944 (N_3944,N_3215,N_3016);
and U3945 (N_3945,N_3035,N_3383);
or U3946 (N_3946,N_3113,N_3252);
xor U3947 (N_3947,N_3372,N_3007);
nor U3948 (N_3948,N_3279,N_3461);
nor U3949 (N_3949,N_3405,N_3514);
nor U3950 (N_3950,N_3726,N_3641);
nor U3951 (N_3951,N_3121,N_3391);
nand U3952 (N_3952,N_3721,N_3102);
and U3953 (N_3953,N_3199,N_3143);
nor U3954 (N_3954,N_3177,N_3691);
or U3955 (N_3955,N_3560,N_3226);
or U3956 (N_3956,N_3586,N_3715);
and U3957 (N_3957,N_3399,N_3330);
and U3958 (N_3958,N_3482,N_3110);
xnor U3959 (N_3959,N_3572,N_3670);
nand U3960 (N_3960,N_3160,N_3426);
nand U3961 (N_3961,N_3735,N_3419);
or U3962 (N_3962,N_3483,N_3487);
or U3963 (N_3963,N_3640,N_3609);
and U3964 (N_3964,N_3598,N_3104);
and U3965 (N_3965,N_3036,N_3063);
or U3966 (N_3966,N_3516,N_3095);
nor U3967 (N_3967,N_3490,N_3008);
or U3968 (N_3968,N_3023,N_3285);
or U3969 (N_3969,N_3096,N_3375);
xor U3970 (N_3970,N_3264,N_3695);
or U3971 (N_3971,N_3498,N_3109);
xor U3972 (N_3972,N_3679,N_3474);
or U3973 (N_3973,N_3385,N_3099);
nor U3974 (N_3974,N_3439,N_3286);
nand U3975 (N_3975,N_3145,N_3671);
nand U3976 (N_3976,N_3414,N_3053);
and U3977 (N_3977,N_3031,N_3616);
nand U3978 (N_3978,N_3528,N_3593);
nand U3979 (N_3979,N_3374,N_3472);
and U3980 (N_3980,N_3523,N_3186);
nand U3981 (N_3981,N_3674,N_3519);
and U3982 (N_3982,N_3486,N_3309);
and U3983 (N_3983,N_3324,N_3421);
xnor U3984 (N_3984,N_3360,N_3451);
xor U3985 (N_3985,N_3561,N_3137);
nand U3986 (N_3986,N_3462,N_3436);
nand U3987 (N_3987,N_3390,N_3659);
or U3988 (N_3988,N_3692,N_3062);
nor U3989 (N_3989,N_3568,N_3615);
nand U3990 (N_3990,N_3333,N_3124);
or U3991 (N_3991,N_3100,N_3185);
or U3992 (N_3992,N_3377,N_3606);
xnor U3993 (N_3993,N_3408,N_3141);
or U3994 (N_3994,N_3125,N_3284);
nor U3995 (N_3995,N_3103,N_3686);
xnor U3996 (N_3996,N_3537,N_3292);
and U3997 (N_3997,N_3334,N_3038);
xor U3998 (N_3998,N_3429,N_3595);
or U3999 (N_3999,N_3601,N_3554);
or U4000 (N_4000,N_3521,N_3502);
nand U4001 (N_4001,N_3734,N_3740);
or U4002 (N_4002,N_3343,N_3507);
and U4003 (N_4003,N_3672,N_3427);
nand U4004 (N_4004,N_3265,N_3253);
or U4005 (N_4005,N_3346,N_3655);
xnor U4006 (N_4006,N_3576,N_3392);
nor U4007 (N_4007,N_3706,N_3643);
or U4008 (N_4008,N_3273,N_3198);
or U4009 (N_4009,N_3673,N_3403);
nand U4010 (N_4010,N_3558,N_3509);
xnor U4011 (N_4011,N_3719,N_3147);
nor U4012 (N_4012,N_3357,N_3411);
nand U4013 (N_4013,N_3009,N_3631);
nor U4014 (N_4014,N_3112,N_3646);
nor U4015 (N_4015,N_3422,N_3477);
nand U4016 (N_4016,N_3495,N_3033);
xnor U4017 (N_4017,N_3194,N_3396);
nor U4018 (N_4018,N_3332,N_3243);
nand U4019 (N_4019,N_3255,N_3216);
nor U4020 (N_4020,N_3132,N_3452);
nand U4021 (N_4021,N_3656,N_3120);
or U4022 (N_4022,N_3585,N_3353);
nand U4023 (N_4023,N_3020,N_3580);
nor U4024 (N_4024,N_3233,N_3258);
nor U4025 (N_4025,N_3278,N_3492);
nor U4026 (N_4026,N_3373,N_3066);
xor U4027 (N_4027,N_3293,N_3047);
or U4028 (N_4028,N_3709,N_3322);
or U4029 (N_4029,N_3001,N_3678);
xor U4030 (N_4030,N_3209,N_3468);
nor U4031 (N_4031,N_3229,N_3645);
xor U4032 (N_4032,N_3344,N_3612);
and U4033 (N_4033,N_3212,N_3128);
or U4034 (N_4034,N_3433,N_3179);
nand U4035 (N_4035,N_3545,N_3190);
xor U4036 (N_4036,N_3481,N_3445);
nor U4037 (N_4037,N_3454,N_3161);
nand U4038 (N_4038,N_3012,N_3026);
xor U4039 (N_4039,N_3562,N_3705);
or U4040 (N_4040,N_3076,N_3270);
or U4041 (N_4041,N_3142,N_3214);
or U4042 (N_4042,N_3683,N_3079);
and U4043 (N_4043,N_3531,N_3449);
and U4044 (N_4044,N_3608,N_3069);
and U4045 (N_4045,N_3068,N_3565);
and U4046 (N_4046,N_3077,N_3307);
and U4047 (N_4047,N_3458,N_3225);
nor U4048 (N_4048,N_3694,N_3175);
nor U4049 (N_4049,N_3230,N_3329);
xnor U4050 (N_4050,N_3687,N_3712);
xnor U4051 (N_4051,N_3122,N_3559);
xnor U4052 (N_4052,N_3747,N_3485);
xnor U4053 (N_4053,N_3431,N_3649);
or U4054 (N_4054,N_3732,N_3717);
nand U4055 (N_4055,N_3469,N_3702);
nor U4056 (N_4056,N_3384,N_3510);
xnor U4057 (N_4057,N_3257,N_3685);
or U4058 (N_4058,N_3213,N_3146);
and U4059 (N_4059,N_3665,N_3611);
nand U4060 (N_4060,N_3088,N_3542);
nor U4061 (N_4061,N_3696,N_3597);
nand U4062 (N_4062,N_3013,N_3594);
nand U4063 (N_4063,N_3337,N_3368);
xor U4064 (N_4064,N_3369,N_3358);
or U4065 (N_4065,N_3688,N_3054);
nor U4066 (N_4066,N_3043,N_3067);
nor U4067 (N_4067,N_3663,N_3676);
or U4068 (N_4068,N_3402,N_3338);
xor U4069 (N_4069,N_3366,N_3620);
or U4070 (N_4070,N_3157,N_3331);
or U4071 (N_4071,N_3060,N_3464);
nor U4072 (N_4072,N_3237,N_3532);
xnor U4073 (N_4073,N_3699,N_3184);
nor U4074 (N_4074,N_3030,N_3080);
and U4075 (N_4075,N_3091,N_3707);
and U4076 (N_4076,N_3205,N_3135);
or U4077 (N_4077,N_3227,N_3204);
or U4078 (N_4078,N_3044,N_3667);
or U4079 (N_4079,N_3169,N_3701);
nor U4080 (N_4080,N_3603,N_3106);
nand U4081 (N_4081,N_3328,N_3349);
nor U4082 (N_4082,N_3730,N_3544);
xor U4083 (N_4083,N_3619,N_3162);
or U4084 (N_4084,N_3749,N_3303);
nor U4085 (N_4085,N_3019,N_3057);
xnor U4086 (N_4086,N_3602,N_3737);
or U4087 (N_4087,N_3232,N_3006);
and U4088 (N_4088,N_3703,N_3406);
or U4089 (N_4089,N_3202,N_3551);
or U4090 (N_4090,N_3050,N_3004);
nor U4091 (N_4091,N_3590,N_3363);
nor U4092 (N_4092,N_3058,N_3465);
nor U4093 (N_4093,N_3082,N_3010);
or U4094 (N_4094,N_3117,N_3267);
xor U4095 (N_4095,N_3634,N_3098);
xor U4096 (N_4096,N_3522,N_3266);
xor U4097 (N_4097,N_3183,N_3557);
xnor U4098 (N_4098,N_3249,N_3084);
or U4099 (N_4099,N_3476,N_3524);
or U4100 (N_4100,N_3207,N_3681);
or U4101 (N_4101,N_3644,N_3493);
nand U4102 (N_4102,N_3367,N_3217);
nor U4103 (N_4103,N_3722,N_3443);
nand U4104 (N_4104,N_3748,N_3164);
xor U4105 (N_4105,N_3444,N_3398);
and U4106 (N_4106,N_3382,N_3362);
xor U4107 (N_4107,N_3271,N_3318);
nor U4108 (N_4108,N_3074,N_3647);
nand U4109 (N_4109,N_3653,N_3306);
nor U4110 (N_4110,N_3027,N_3710);
xnor U4111 (N_4111,N_3417,N_3371);
xor U4112 (N_4112,N_3148,N_3596);
xnor U4113 (N_4113,N_3022,N_3092);
xnor U4114 (N_4114,N_3579,N_3423);
nand U4115 (N_4115,N_3389,N_3254);
and U4116 (N_4116,N_3056,N_3200);
and U4117 (N_4117,N_3736,N_3055);
nand U4118 (N_4118,N_3269,N_3505);
nor U4119 (N_4119,N_3533,N_3395);
nand U4120 (N_4120,N_3387,N_3527);
nand U4121 (N_4121,N_3448,N_3283);
nand U4122 (N_4122,N_3651,N_3555);
nor U4123 (N_4123,N_3718,N_3274);
nand U4124 (N_4124,N_3689,N_3297);
xnor U4125 (N_4125,N_3295,N_3230);
nand U4126 (N_4126,N_3323,N_3540);
xor U4127 (N_4127,N_3515,N_3662);
and U4128 (N_4128,N_3020,N_3200);
xor U4129 (N_4129,N_3395,N_3013);
and U4130 (N_4130,N_3286,N_3590);
and U4131 (N_4131,N_3553,N_3379);
xnor U4132 (N_4132,N_3265,N_3672);
nor U4133 (N_4133,N_3436,N_3404);
nand U4134 (N_4134,N_3115,N_3604);
nand U4135 (N_4135,N_3222,N_3649);
nand U4136 (N_4136,N_3565,N_3468);
and U4137 (N_4137,N_3261,N_3066);
or U4138 (N_4138,N_3249,N_3389);
and U4139 (N_4139,N_3562,N_3686);
or U4140 (N_4140,N_3719,N_3492);
nor U4141 (N_4141,N_3471,N_3025);
or U4142 (N_4142,N_3648,N_3573);
or U4143 (N_4143,N_3295,N_3209);
nor U4144 (N_4144,N_3513,N_3626);
xor U4145 (N_4145,N_3474,N_3211);
nand U4146 (N_4146,N_3464,N_3318);
or U4147 (N_4147,N_3286,N_3278);
and U4148 (N_4148,N_3490,N_3034);
nand U4149 (N_4149,N_3603,N_3271);
xnor U4150 (N_4150,N_3071,N_3449);
nand U4151 (N_4151,N_3385,N_3558);
nand U4152 (N_4152,N_3092,N_3233);
nor U4153 (N_4153,N_3664,N_3710);
nand U4154 (N_4154,N_3587,N_3042);
and U4155 (N_4155,N_3380,N_3184);
xor U4156 (N_4156,N_3741,N_3017);
xor U4157 (N_4157,N_3387,N_3425);
xnor U4158 (N_4158,N_3356,N_3732);
xnor U4159 (N_4159,N_3337,N_3424);
or U4160 (N_4160,N_3138,N_3322);
xnor U4161 (N_4161,N_3342,N_3363);
xnor U4162 (N_4162,N_3573,N_3520);
nor U4163 (N_4163,N_3011,N_3331);
or U4164 (N_4164,N_3550,N_3486);
nor U4165 (N_4165,N_3555,N_3625);
nand U4166 (N_4166,N_3458,N_3262);
xnor U4167 (N_4167,N_3536,N_3295);
or U4168 (N_4168,N_3241,N_3657);
xnor U4169 (N_4169,N_3032,N_3416);
xor U4170 (N_4170,N_3044,N_3520);
and U4171 (N_4171,N_3108,N_3505);
nand U4172 (N_4172,N_3674,N_3029);
nor U4173 (N_4173,N_3609,N_3255);
or U4174 (N_4174,N_3028,N_3066);
or U4175 (N_4175,N_3390,N_3429);
nor U4176 (N_4176,N_3306,N_3576);
xnor U4177 (N_4177,N_3143,N_3689);
or U4178 (N_4178,N_3164,N_3421);
or U4179 (N_4179,N_3029,N_3708);
xnor U4180 (N_4180,N_3097,N_3131);
xor U4181 (N_4181,N_3228,N_3649);
nand U4182 (N_4182,N_3592,N_3524);
xnor U4183 (N_4183,N_3456,N_3264);
and U4184 (N_4184,N_3024,N_3071);
or U4185 (N_4185,N_3341,N_3585);
and U4186 (N_4186,N_3541,N_3649);
nor U4187 (N_4187,N_3052,N_3291);
nand U4188 (N_4188,N_3459,N_3710);
nand U4189 (N_4189,N_3039,N_3598);
xor U4190 (N_4190,N_3463,N_3485);
nand U4191 (N_4191,N_3124,N_3488);
or U4192 (N_4192,N_3575,N_3036);
or U4193 (N_4193,N_3374,N_3144);
xnor U4194 (N_4194,N_3331,N_3737);
nor U4195 (N_4195,N_3270,N_3255);
nand U4196 (N_4196,N_3632,N_3133);
and U4197 (N_4197,N_3451,N_3075);
and U4198 (N_4198,N_3339,N_3538);
or U4199 (N_4199,N_3472,N_3556);
and U4200 (N_4200,N_3620,N_3491);
or U4201 (N_4201,N_3690,N_3161);
nand U4202 (N_4202,N_3020,N_3594);
xor U4203 (N_4203,N_3644,N_3295);
nor U4204 (N_4204,N_3382,N_3196);
nand U4205 (N_4205,N_3629,N_3724);
nand U4206 (N_4206,N_3346,N_3123);
nor U4207 (N_4207,N_3667,N_3448);
nand U4208 (N_4208,N_3326,N_3329);
or U4209 (N_4209,N_3513,N_3193);
and U4210 (N_4210,N_3553,N_3507);
and U4211 (N_4211,N_3213,N_3628);
nand U4212 (N_4212,N_3569,N_3363);
and U4213 (N_4213,N_3464,N_3553);
or U4214 (N_4214,N_3410,N_3537);
nand U4215 (N_4215,N_3572,N_3553);
or U4216 (N_4216,N_3101,N_3237);
and U4217 (N_4217,N_3249,N_3330);
or U4218 (N_4218,N_3314,N_3700);
nand U4219 (N_4219,N_3421,N_3724);
xor U4220 (N_4220,N_3253,N_3362);
nor U4221 (N_4221,N_3018,N_3653);
and U4222 (N_4222,N_3100,N_3176);
nor U4223 (N_4223,N_3125,N_3415);
or U4224 (N_4224,N_3600,N_3423);
or U4225 (N_4225,N_3256,N_3234);
nor U4226 (N_4226,N_3277,N_3651);
nand U4227 (N_4227,N_3139,N_3597);
nor U4228 (N_4228,N_3112,N_3539);
xnor U4229 (N_4229,N_3251,N_3663);
and U4230 (N_4230,N_3301,N_3460);
xnor U4231 (N_4231,N_3520,N_3665);
and U4232 (N_4232,N_3012,N_3469);
and U4233 (N_4233,N_3264,N_3302);
and U4234 (N_4234,N_3239,N_3426);
or U4235 (N_4235,N_3425,N_3173);
nand U4236 (N_4236,N_3485,N_3236);
and U4237 (N_4237,N_3606,N_3689);
nor U4238 (N_4238,N_3269,N_3043);
and U4239 (N_4239,N_3641,N_3186);
xnor U4240 (N_4240,N_3297,N_3719);
nor U4241 (N_4241,N_3144,N_3050);
nand U4242 (N_4242,N_3615,N_3194);
nor U4243 (N_4243,N_3478,N_3176);
xnor U4244 (N_4244,N_3247,N_3551);
and U4245 (N_4245,N_3519,N_3566);
xor U4246 (N_4246,N_3508,N_3064);
or U4247 (N_4247,N_3011,N_3568);
or U4248 (N_4248,N_3737,N_3395);
and U4249 (N_4249,N_3539,N_3592);
nor U4250 (N_4250,N_3262,N_3304);
nand U4251 (N_4251,N_3662,N_3029);
xor U4252 (N_4252,N_3253,N_3483);
nor U4253 (N_4253,N_3641,N_3662);
nand U4254 (N_4254,N_3196,N_3623);
xnor U4255 (N_4255,N_3001,N_3331);
and U4256 (N_4256,N_3598,N_3493);
xor U4257 (N_4257,N_3431,N_3097);
and U4258 (N_4258,N_3195,N_3360);
or U4259 (N_4259,N_3535,N_3140);
or U4260 (N_4260,N_3718,N_3416);
or U4261 (N_4261,N_3351,N_3387);
nand U4262 (N_4262,N_3231,N_3667);
nand U4263 (N_4263,N_3749,N_3558);
or U4264 (N_4264,N_3461,N_3660);
xnor U4265 (N_4265,N_3255,N_3452);
nor U4266 (N_4266,N_3358,N_3477);
nor U4267 (N_4267,N_3455,N_3387);
xor U4268 (N_4268,N_3015,N_3244);
and U4269 (N_4269,N_3260,N_3702);
or U4270 (N_4270,N_3323,N_3560);
or U4271 (N_4271,N_3482,N_3296);
or U4272 (N_4272,N_3157,N_3565);
or U4273 (N_4273,N_3292,N_3660);
and U4274 (N_4274,N_3621,N_3001);
and U4275 (N_4275,N_3730,N_3643);
nor U4276 (N_4276,N_3170,N_3540);
nand U4277 (N_4277,N_3115,N_3102);
xnor U4278 (N_4278,N_3045,N_3281);
nor U4279 (N_4279,N_3095,N_3044);
or U4280 (N_4280,N_3492,N_3238);
xnor U4281 (N_4281,N_3478,N_3722);
or U4282 (N_4282,N_3431,N_3492);
nor U4283 (N_4283,N_3111,N_3039);
xor U4284 (N_4284,N_3225,N_3702);
nand U4285 (N_4285,N_3639,N_3110);
and U4286 (N_4286,N_3731,N_3232);
nand U4287 (N_4287,N_3363,N_3255);
xor U4288 (N_4288,N_3037,N_3262);
nand U4289 (N_4289,N_3454,N_3494);
xnor U4290 (N_4290,N_3610,N_3154);
nand U4291 (N_4291,N_3321,N_3615);
or U4292 (N_4292,N_3514,N_3324);
and U4293 (N_4293,N_3510,N_3645);
and U4294 (N_4294,N_3356,N_3410);
xnor U4295 (N_4295,N_3632,N_3205);
nand U4296 (N_4296,N_3668,N_3623);
nor U4297 (N_4297,N_3126,N_3221);
nor U4298 (N_4298,N_3056,N_3226);
xor U4299 (N_4299,N_3560,N_3137);
xor U4300 (N_4300,N_3576,N_3557);
or U4301 (N_4301,N_3510,N_3570);
or U4302 (N_4302,N_3318,N_3529);
xnor U4303 (N_4303,N_3690,N_3712);
and U4304 (N_4304,N_3357,N_3030);
xor U4305 (N_4305,N_3047,N_3467);
xor U4306 (N_4306,N_3162,N_3142);
xnor U4307 (N_4307,N_3541,N_3493);
or U4308 (N_4308,N_3542,N_3707);
nor U4309 (N_4309,N_3076,N_3330);
and U4310 (N_4310,N_3607,N_3658);
xnor U4311 (N_4311,N_3600,N_3147);
or U4312 (N_4312,N_3725,N_3675);
or U4313 (N_4313,N_3095,N_3444);
xor U4314 (N_4314,N_3064,N_3447);
or U4315 (N_4315,N_3143,N_3625);
or U4316 (N_4316,N_3347,N_3416);
nand U4317 (N_4317,N_3352,N_3490);
nor U4318 (N_4318,N_3014,N_3548);
nand U4319 (N_4319,N_3505,N_3667);
or U4320 (N_4320,N_3271,N_3166);
nand U4321 (N_4321,N_3032,N_3730);
and U4322 (N_4322,N_3543,N_3322);
nand U4323 (N_4323,N_3276,N_3032);
nand U4324 (N_4324,N_3225,N_3735);
nand U4325 (N_4325,N_3737,N_3099);
nand U4326 (N_4326,N_3260,N_3360);
and U4327 (N_4327,N_3513,N_3223);
nor U4328 (N_4328,N_3092,N_3226);
xor U4329 (N_4329,N_3084,N_3345);
xnor U4330 (N_4330,N_3132,N_3312);
or U4331 (N_4331,N_3245,N_3178);
xnor U4332 (N_4332,N_3180,N_3145);
nor U4333 (N_4333,N_3640,N_3124);
nor U4334 (N_4334,N_3077,N_3576);
nand U4335 (N_4335,N_3014,N_3202);
nand U4336 (N_4336,N_3595,N_3300);
and U4337 (N_4337,N_3135,N_3442);
xor U4338 (N_4338,N_3587,N_3041);
nand U4339 (N_4339,N_3304,N_3368);
xor U4340 (N_4340,N_3393,N_3180);
or U4341 (N_4341,N_3159,N_3348);
nor U4342 (N_4342,N_3451,N_3156);
or U4343 (N_4343,N_3212,N_3614);
xnor U4344 (N_4344,N_3107,N_3292);
and U4345 (N_4345,N_3418,N_3745);
xnor U4346 (N_4346,N_3243,N_3637);
xnor U4347 (N_4347,N_3480,N_3604);
and U4348 (N_4348,N_3008,N_3317);
and U4349 (N_4349,N_3327,N_3632);
nand U4350 (N_4350,N_3386,N_3432);
xor U4351 (N_4351,N_3154,N_3496);
xnor U4352 (N_4352,N_3669,N_3435);
or U4353 (N_4353,N_3233,N_3281);
or U4354 (N_4354,N_3639,N_3035);
nand U4355 (N_4355,N_3393,N_3023);
nor U4356 (N_4356,N_3526,N_3243);
xnor U4357 (N_4357,N_3367,N_3417);
nor U4358 (N_4358,N_3274,N_3561);
and U4359 (N_4359,N_3350,N_3255);
and U4360 (N_4360,N_3263,N_3652);
and U4361 (N_4361,N_3053,N_3216);
or U4362 (N_4362,N_3215,N_3366);
nor U4363 (N_4363,N_3347,N_3129);
or U4364 (N_4364,N_3201,N_3129);
or U4365 (N_4365,N_3186,N_3070);
and U4366 (N_4366,N_3131,N_3288);
or U4367 (N_4367,N_3039,N_3678);
xnor U4368 (N_4368,N_3129,N_3311);
nor U4369 (N_4369,N_3338,N_3066);
nand U4370 (N_4370,N_3670,N_3531);
nor U4371 (N_4371,N_3103,N_3044);
xor U4372 (N_4372,N_3068,N_3252);
and U4373 (N_4373,N_3683,N_3595);
nand U4374 (N_4374,N_3259,N_3227);
xnor U4375 (N_4375,N_3427,N_3030);
nand U4376 (N_4376,N_3502,N_3479);
and U4377 (N_4377,N_3648,N_3088);
or U4378 (N_4378,N_3348,N_3535);
and U4379 (N_4379,N_3271,N_3002);
nand U4380 (N_4380,N_3475,N_3132);
and U4381 (N_4381,N_3733,N_3742);
nor U4382 (N_4382,N_3556,N_3433);
and U4383 (N_4383,N_3636,N_3395);
or U4384 (N_4384,N_3278,N_3219);
nand U4385 (N_4385,N_3720,N_3586);
nor U4386 (N_4386,N_3307,N_3473);
or U4387 (N_4387,N_3515,N_3443);
and U4388 (N_4388,N_3004,N_3243);
or U4389 (N_4389,N_3610,N_3328);
or U4390 (N_4390,N_3489,N_3385);
or U4391 (N_4391,N_3584,N_3479);
nor U4392 (N_4392,N_3290,N_3417);
nor U4393 (N_4393,N_3398,N_3505);
and U4394 (N_4394,N_3007,N_3022);
nor U4395 (N_4395,N_3167,N_3569);
or U4396 (N_4396,N_3320,N_3422);
nor U4397 (N_4397,N_3584,N_3384);
nand U4398 (N_4398,N_3079,N_3443);
xor U4399 (N_4399,N_3297,N_3613);
nand U4400 (N_4400,N_3023,N_3163);
xor U4401 (N_4401,N_3746,N_3455);
nor U4402 (N_4402,N_3432,N_3632);
nand U4403 (N_4403,N_3722,N_3388);
and U4404 (N_4404,N_3280,N_3338);
and U4405 (N_4405,N_3555,N_3259);
nand U4406 (N_4406,N_3495,N_3417);
and U4407 (N_4407,N_3182,N_3426);
nor U4408 (N_4408,N_3676,N_3543);
and U4409 (N_4409,N_3296,N_3565);
xor U4410 (N_4410,N_3370,N_3254);
nand U4411 (N_4411,N_3690,N_3307);
nand U4412 (N_4412,N_3398,N_3286);
nor U4413 (N_4413,N_3163,N_3042);
nor U4414 (N_4414,N_3372,N_3090);
xnor U4415 (N_4415,N_3211,N_3309);
nor U4416 (N_4416,N_3311,N_3629);
or U4417 (N_4417,N_3568,N_3455);
xnor U4418 (N_4418,N_3141,N_3478);
and U4419 (N_4419,N_3605,N_3528);
or U4420 (N_4420,N_3271,N_3484);
nor U4421 (N_4421,N_3010,N_3295);
and U4422 (N_4422,N_3509,N_3423);
nand U4423 (N_4423,N_3436,N_3431);
nor U4424 (N_4424,N_3664,N_3363);
and U4425 (N_4425,N_3483,N_3697);
nand U4426 (N_4426,N_3526,N_3239);
or U4427 (N_4427,N_3680,N_3602);
or U4428 (N_4428,N_3569,N_3547);
xnor U4429 (N_4429,N_3152,N_3074);
nand U4430 (N_4430,N_3554,N_3664);
xor U4431 (N_4431,N_3638,N_3483);
or U4432 (N_4432,N_3456,N_3288);
nand U4433 (N_4433,N_3533,N_3698);
and U4434 (N_4434,N_3535,N_3507);
or U4435 (N_4435,N_3003,N_3201);
xor U4436 (N_4436,N_3239,N_3623);
or U4437 (N_4437,N_3406,N_3162);
xor U4438 (N_4438,N_3232,N_3545);
or U4439 (N_4439,N_3112,N_3052);
nand U4440 (N_4440,N_3324,N_3164);
and U4441 (N_4441,N_3632,N_3039);
xnor U4442 (N_4442,N_3342,N_3591);
nor U4443 (N_4443,N_3519,N_3286);
xor U4444 (N_4444,N_3281,N_3358);
or U4445 (N_4445,N_3137,N_3415);
and U4446 (N_4446,N_3580,N_3333);
nor U4447 (N_4447,N_3062,N_3451);
nand U4448 (N_4448,N_3615,N_3414);
and U4449 (N_4449,N_3638,N_3366);
nand U4450 (N_4450,N_3353,N_3607);
and U4451 (N_4451,N_3279,N_3365);
or U4452 (N_4452,N_3642,N_3568);
and U4453 (N_4453,N_3723,N_3645);
and U4454 (N_4454,N_3723,N_3492);
and U4455 (N_4455,N_3574,N_3162);
nor U4456 (N_4456,N_3039,N_3540);
or U4457 (N_4457,N_3448,N_3079);
or U4458 (N_4458,N_3464,N_3195);
nand U4459 (N_4459,N_3167,N_3654);
nor U4460 (N_4460,N_3557,N_3582);
nand U4461 (N_4461,N_3662,N_3041);
and U4462 (N_4462,N_3688,N_3323);
nor U4463 (N_4463,N_3488,N_3383);
and U4464 (N_4464,N_3440,N_3624);
nand U4465 (N_4465,N_3152,N_3723);
or U4466 (N_4466,N_3327,N_3433);
and U4467 (N_4467,N_3638,N_3257);
xor U4468 (N_4468,N_3665,N_3161);
nand U4469 (N_4469,N_3117,N_3127);
nand U4470 (N_4470,N_3723,N_3198);
xnor U4471 (N_4471,N_3527,N_3021);
or U4472 (N_4472,N_3648,N_3326);
and U4473 (N_4473,N_3116,N_3230);
and U4474 (N_4474,N_3100,N_3288);
or U4475 (N_4475,N_3039,N_3098);
or U4476 (N_4476,N_3012,N_3062);
or U4477 (N_4477,N_3674,N_3685);
nor U4478 (N_4478,N_3739,N_3081);
xnor U4479 (N_4479,N_3066,N_3224);
nor U4480 (N_4480,N_3246,N_3176);
xor U4481 (N_4481,N_3331,N_3372);
and U4482 (N_4482,N_3734,N_3110);
xor U4483 (N_4483,N_3000,N_3726);
nor U4484 (N_4484,N_3315,N_3742);
xnor U4485 (N_4485,N_3567,N_3336);
and U4486 (N_4486,N_3273,N_3365);
nor U4487 (N_4487,N_3328,N_3053);
nand U4488 (N_4488,N_3572,N_3242);
xnor U4489 (N_4489,N_3043,N_3685);
or U4490 (N_4490,N_3192,N_3748);
or U4491 (N_4491,N_3143,N_3696);
or U4492 (N_4492,N_3402,N_3050);
and U4493 (N_4493,N_3128,N_3294);
nand U4494 (N_4494,N_3286,N_3007);
nand U4495 (N_4495,N_3173,N_3232);
xnor U4496 (N_4496,N_3554,N_3743);
and U4497 (N_4497,N_3170,N_3519);
or U4498 (N_4498,N_3535,N_3735);
nor U4499 (N_4499,N_3449,N_3619);
or U4500 (N_4500,N_4001,N_3783);
or U4501 (N_4501,N_4244,N_4461);
xnor U4502 (N_4502,N_4494,N_4190);
or U4503 (N_4503,N_4481,N_4052);
nor U4504 (N_4504,N_4442,N_4392);
nor U4505 (N_4505,N_3907,N_4249);
and U4506 (N_4506,N_3928,N_4310);
xnor U4507 (N_4507,N_4100,N_4431);
xnor U4508 (N_4508,N_4437,N_4388);
and U4509 (N_4509,N_3792,N_4069);
xor U4510 (N_4510,N_4467,N_4404);
or U4511 (N_4511,N_3857,N_4332);
and U4512 (N_4512,N_4355,N_4314);
nor U4513 (N_4513,N_4391,N_3956);
nand U4514 (N_4514,N_4080,N_4041);
nand U4515 (N_4515,N_4232,N_4495);
and U4516 (N_4516,N_3833,N_4172);
or U4517 (N_4517,N_3766,N_4082);
nor U4518 (N_4518,N_4476,N_4434);
and U4519 (N_4519,N_4270,N_4105);
nor U4520 (N_4520,N_3870,N_3859);
or U4521 (N_4521,N_4078,N_4179);
and U4522 (N_4522,N_4366,N_3824);
nand U4523 (N_4523,N_4073,N_4400);
nor U4524 (N_4524,N_3986,N_3891);
or U4525 (N_4525,N_3784,N_3980);
nand U4526 (N_4526,N_3968,N_4148);
and U4527 (N_4527,N_4091,N_4125);
and U4528 (N_4528,N_4225,N_4349);
and U4529 (N_4529,N_4102,N_4212);
nand U4530 (N_4530,N_4305,N_4061);
and U4531 (N_4531,N_4139,N_4129);
and U4532 (N_4532,N_4140,N_4242);
nor U4533 (N_4533,N_4356,N_4432);
nand U4534 (N_4534,N_4004,N_3781);
xor U4535 (N_4535,N_4060,N_4479);
xnor U4536 (N_4536,N_3881,N_4186);
and U4537 (N_4537,N_3752,N_4448);
nand U4538 (N_4538,N_4096,N_4047);
and U4539 (N_4539,N_3973,N_3964);
nor U4540 (N_4540,N_4385,N_3890);
or U4541 (N_4541,N_4439,N_3768);
xor U4542 (N_4542,N_4414,N_4455);
and U4543 (N_4543,N_3778,N_3946);
nor U4544 (N_4544,N_4138,N_4048);
nand U4545 (N_4545,N_4281,N_3905);
and U4546 (N_4546,N_4260,N_4440);
nor U4547 (N_4547,N_4173,N_3971);
xor U4548 (N_4548,N_3895,N_3985);
or U4549 (N_4549,N_4311,N_4303);
nor U4550 (N_4550,N_4031,N_3995);
nor U4551 (N_4551,N_3811,N_4044);
xnor U4552 (N_4552,N_4022,N_3931);
nor U4553 (N_4553,N_4407,N_4178);
or U4554 (N_4554,N_3771,N_4288);
or U4555 (N_4555,N_4452,N_3983);
nand U4556 (N_4556,N_4338,N_4177);
nor U4557 (N_4557,N_4197,N_3809);
nand U4558 (N_4558,N_3885,N_3765);
or U4559 (N_4559,N_3860,N_4194);
nor U4560 (N_4560,N_4321,N_4387);
and U4561 (N_4561,N_4368,N_4315);
or U4562 (N_4562,N_4327,N_3994);
nor U4563 (N_4563,N_3844,N_3990);
nor U4564 (N_4564,N_3865,N_4235);
xor U4565 (N_4565,N_4224,N_3921);
xnor U4566 (N_4566,N_4214,N_3789);
nand U4567 (N_4567,N_3972,N_3967);
xnor U4568 (N_4568,N_4317,N_4243);
nor U4569 (N_4569,N_4333,N_4341);
and U4570 (N_4570,N_3919,N_4456);
nor U4571 (N_4571,N_3853,N_4464);
and U4572 (N_4572,N_4119,N_3805);
and U4573 (N_4573,N_4283,N_4189);
and U4574 (N_4574,N_3879,N_4067);
or U4575 (N_4575,N_4297,N_3812);
or U4576 (N_4576,N_3757,N_3910);
and U4577 (N_4577,N_4241,N_3904);
or U4578 (N_4578,N_4154,N_4115);
xor U4579 (N_4579,N_4493,N_4365);
nor U4580 (N_4580,N_3818,N_4423);
and U4581 (N_4581,N_4227,N_3796);
xnor U4582 (N_4582,N_3991,N_4081);
and U4583 (N_4583,N_3875,N_4231);
or U4584 (N_4584,N_4378,N_4421);
nor U4585 (N_4585,N_3843,N_4162);
nand U4586 (N_4586,N_4482,N_3832);
and U4587 (N_4587,N_4131,N_4422);
nand U4588 (N_4588,N_4083,N_4465);
or U4589 (N_4589,N_4344,N_4253);
xnor U4590 (N_4590,N_3961,N_3909);
nor U4591 (N_4591,N_4438,N_4003);
and U4592 (N_4592,N_3958,N_3878);
and U4593 (N_4593,N_4141,N_4259);
nor U4594 (N_4594,N_4352,N_4059);
nand U4595 (N_4595,N_4245,N_4451);
xnor U4596 (N_4596,N_3976,N_4294);
xnor U4597 (N_4597,N_4436,N_3925);
or U4598 (N_4598,N_4399,N_4118);
xor U4599 (N_4599,N_4166,N_4357);
nand U4600 (N_4600,N_3918,N_3851);
or U4601 (N_4601,N_4114,N_4071);
nor U4602 (N_4602,N_4364,N_3916);
nor U4603 (N_4603,N_4217,N_4329);
and U4604 (N_4604,N_3948,N_4203);
and U4605 (N_4605,N_4200,N_3868);
nand U4606 (N_4606,N_3975,N_3863);
xnor U4607 (N_4607,N_4425,N_4405);
nor U4608 (N_4608,N_4480,N_4340);
and U4609 (N_4609,N_4057,N_4374);
or U4610 (N_4610,N_3871,N_4184);
and U4611 (N_4611,N_3869,N_4412);
nor U4612 (N_4612,N_4324,N_3800);
nand U4613 (N_4613,N_3930,N_3835);
xor U4614 (N_4614,N_4144,N_4360);
xor U4615 (N_4615,N_3799,N_3953);
xnor U4616 (N_4616,N_4074,N_4209);
and U4617 (N_4617,N_4109,N_4345);
nand U4618 (N_4618,N_4199,N_4343);
or U4619 (N_4619,N_4488,N_3940);
xnor U4620 (N_4620,N_3906,N_4301);
and U4621 (N_4621,N_3831,N_4441);
nor U4622 (N_4622,N_4175,N_3810);
xor U4623 (N_4623,N_3883,N_4282);
nand U4624 (N_4624,N_4049,N_3756);
nor U4625 (N_4625,N_3937,N_3776);
nor U4626 (N_4626,N_3962,N_4444);
nand U4627 (N_4627,N_4429,N_3880);
nand U4628 (N_4628,N_4468,N_4191);
xor U4629 (N_4629,N_4383,N_4171);
or U4630 (N_4630,N_3917,N_4272);
xor U4631 (N_4631,N_4009,N_4239);
and U4632 (N_4632,N_4185,N_4134);
and U4633 (N_4633,N_4336,N_4123);
nand U4634 (N_4634,N_4070,N_4371);
or U4635 (N_4635,N_4393,N_4274);
xor U4636 (N_4636,N_3888,N_3775);
nand U4637 (N_4637,N_3753,N_4248);
nand U4638 (N_4638,N_4228,N_4149);
xnor U4639 (N_4639,N_4062,N_4229);
or U4640 (N_4640,N_4150,N_3816);
or U4641 (N_4641,N_3938,N_4168);
nor U4642 (N_4642,N_4300,N_4453);
nand U4643 (N_4643,N_4251,N_3866);
nor U4644 (N_4644,N_4051,N_3798);
or U4645 (N_4645,N_4319,N_3855);
nor U4646 (N_4646,N_4183,N_4326);
xnor U4647 (N_4647,N_4126,N_3852);
and U4648 (N_4648,N_4361,N_4406);
nor U4649 (N_4649,N_4142,N_4408);
and U4650 (N_4650,N_4426,N_4111);
and U4651 (N_4651,N_3797,N_4450);
or U4652 (N_4652,N_4273,N_4198);
nor U4653 (N_4653,N_4396,N_4117);
nand U4654 (N_4654,N_4005,N_4193);
xor U4655 (N_4655,N_3817,N_3900);
xor U4656 (N_4656,N_3893,N_4316);
and U4657 (N_4657,N_4017,N_4181);
or U4658 (N_4658,N_4309,N_4269);
or U4659 (N_4659,N_3882,N_4018);
nand U4660 (N_4660,N_4328,N_3989);
or U4661 (N_4661,N_3970,N_4484);
nor U4662 (N_4662,N_3767,N_4325);
or U4663 (N_4663,N_3899,N_4420);
nor U4664 (N_4664,N_3872,N_4158);
nor U4665 (N_4665,N_3785,N_4084);
nor U4666 (N_4666,N_4362,N_3849);
xor U4667 (N_4667,N_4469,N_3957);
nor U4668 (N_4668,N_3820,N_4076);
nor U4669 (N_4669,N_4295,N_4237);
or U4670 (N_4670,N_4443,N_4471);
nor U4671 (N_4671,N_4014,N_4331);
and U4672 (N_4672,N_3760,N_4233);
xor U4673 (N_4673,N_4223,N_3836);
nand U4674 (N_4674,N_4077,N_3790);
nor U4675 (N_4675,N_3819,N_4053);
nor U4676 (N_4676,N_3960,N_3802);
or U4677 (N_4677,N_3952,N_4358);
and U4678 (N_4678,N_3988,N_4120);
or U4679 (N_4679,N_3955,N_3806);
nor U4680 (N_4680,N_4458,N_4353);
or U4681 (N_4681,N_4473,N_4024);
nand U4682 (N_4682,N_3898,N_3821);
nor U4683 (N_4683,N_4152,N_4276);
and U4684 (N_4684,N_4000,N_4234);
xor U4685 (N_4685,N_4137,N_4020);
nor U4686 (N_4686,N_3770,N_3787);
or U4687 (N_4687,N_3793,N_4055);
xnor U4688 (N_4688,N_4428,N_4106);
xnor U4689 (N_4689,N_3932,N_4130);
or U4690 (N_4690,N_4278,N_4065);
and U4691 (N_4691,N_4155,N_4033);
and U4692 (N_4692,N_4008,N_3999);
nand U4693 (N_4693,N_4221,N_3902);
and U4694 (N_4694,N_4409,N_4112);
and U4695 (N_4695,N_4489,N_4342);
nand U4696 (N_4696,N_3992,N_4038);
and U4697 (N_4697,N_4402,N_4339);
nor U4698 (N_4698,N_4165,N_4466);
xor U4699 (N_4699,N_3929,N_4007);
and U4700 (N_4700,N_4167,N_3837);
nand U4701 (N_4701,N_4085,N_4416);
xnor U4702 (N_4702,N_3842,N_4367);
xor U4703 (N_4703,N_3764,N_4287);
nand U4704 (N_4704,N_3772,N_4029);
nand U4705 (N_4705,N_4021,N_3815);
or U4706 (N_4706,N_3795,N_4213);
or U4707 (N_4707,N_3779,N_4246);
xnor U4708 (N_4708,N_4472,N_4204);
nand U4709 (N_4709,N_4323,N_3887);
nand U4710 (N_4710,N_3982,N_3808);
and U4711 (N_4711,N_3981,N_3920);
xnor U4712 (N_4712,N_4263,N_4187);
xor U4713 (N_4713,N_4320,N_4359);
and U4714 (N_4714,N_3965,N_3969);
and U4715 (N_4715,N_4116,N_4267);
nand U4716 (N_4716,N_4289,N_3814);
xor U4717 (N_4717,N_4348,N_4026);
xnor U4718 (N_4718,N_4153,N_4335);
xnor U4719 (N_4719,N_4036,N_4277);
or U4720 (N_4720,N_4216,N_3864);
nand U4721 (N_4721,N_3834,N_4394);
nor U4722 (N_4722,N_4054,N_4397);
nand U4723 (N_4723,N_4170,N_4296);
nand U4724 (N_4724,N_4491,N_4043);
nand U4725 (N_4725,N_3892,N_4334);
nand U4726 (N_4726,N_4121,N_4133);
nand U4727 (N_4727,N_4252,N_4284);
nand U4728 (N_4728,N_3762,N_3913);
or U4729 (N_4729,N_4499,N_4337);
nor U4730 (N_4730,N_3949,N_4487);
nand U4731 (N_4731,N_4090,N_4159);
nand U4732 (N_4732,N_3897,N_4164);
or U4733 (N_4733,N_4032,N_4146);
nand U4734 (N_4734,N_4382,N_4386);
xor U4735 (N_4735,N_3966,N_4035);
nor U4736 (N_4736,N_4478,N_4098);
nor U4737 (N_4737,N_3894,N_4110);
nand U4738 (N_4738,N_3791,N_4483);
xnor U4739 (N_4739,N_4463,N_3873);
nand U4740 (N_4740,N_4046,N_4006);
and U4741 (N_4741,N_4218,N_3828);
or U4742 (N_4742,N_4210,N_4066);
xor U4743 (N_4743,N_4390,N_3854);
xor U4744 (N_4744,N_4424,N_4169);
or U4745 (N_4745,N_4285,N_4013);
nand U4746 (N_4746,N_3933,N_4097);
or U4747 (N_4747,N_4298,N_4195);
or U4748 (N_4748,N_3987,N_4028);
xnor U4749 (N_4749,N_3825,N_3856);
nor U4750 (N_4750,N_4226,N_3794);
xor U4751 (N_4751,N_4485,N_3786);
xor U4752 (N_4752,N_4304,N_4180);
xnor U4753 (N_4753,N_4019,N_4446);
xor U4754 (N_4754,N_3773,N_3977);
nand U4755 (N_4755,N_4215,N_4135);
xor U4756 (N_4756,N_3823,N_4430);
nand U4757 (N_4757,N_3841,N_4376);
nor U4758 (N_4758,N_4264,N_4445);
or U4759 (N_4759,N_4350,N_4163);
and U4760 (N_4760,N_4088,N_4275);
xor U4761 (N_4761,N_4064,N_4079);
xnor U4762 (N_4762,N_3993,N_4381);
nand U4763 (N_4763,N_4373,N_3780);
and U4764 (N_4764,N_4011,N_4056);
xor U4765 (N_4765,N_4346,N_4262);
xnor U4766 (N_4766,N_4312,N_4271);
nand U4767 (N_4767,N_4354,N_4384);
nor U4768 (N_4768,N_4104,N_4286);
xnor U4769 (N_4769,N_3826,N_4261);
and U4770 (N_4770,N_3846,N_4145);
nor U4771 (N_4771,N_4208,N_3774);
nor U4772 (N_4772,N_4247,N_4042);
and U4773 (N_4773,N_4092,N_4403);
and U4774 (N_4774,N_4415,N_4457);
xor U4775 (N_4775,N_3963,N_3912);
nor U4776 (N_4776,N_3862,N_4240);
xnor U4777 (N_4777,N_3889,N_3751);
or U4778 (N_4778,N_4174,N_4498);
xnor U4779 (N_4779,N_3761,N_4474);
xnor U4780 (N_4780,N_3755,N_3908);
nand U4781 (N_4781,N_3804,N_3759);
xor U4782 (N_4782,N_3934,N_4413);
and U4783 (N_4783,N_4023,N_4419);
or U4784 (N_4784,N_4016,N_4477);
or U4785 (N_4785,N_4040,N_4127);
nor U4786 (N_4786,N_4351,N_3763);
xor U4787 (N_4787,N_4108,N_4087);
nor U4788 (N_4788,N_4449,N_3943);
and U4789 (N_4789,N_4002,N_4265);
xor U4790 (N_4790,N_4492,N_4279);
nand U4791 (N_4791,N_3822,N_4072);
xor U4792 (N_4792,N_4188,N_3874);
nand U4793 (N_4793,N_3959,N_4380);
xnor U4794 (N_4794,N_4280,N_4201);
nor U4795 (N_4795,N_4490,N_4496);
and U4796 (N_4796,N_4307,N_4068);
or U4797 (N_4797,N_4132,N_4401);
nor U4798 (N_4798,N_4250,N_3979);
or U4799 (N_4799,N_3861,N_4462);
nand U4800 (N_4800,N_3884,N_4375);
and U4801 (N_4801,N_3901,N_3840);
nand U4802 (N_4802,N_4369,N_3876);
or U4803 (N_4803,N_3922,N_4030);
or U4804 (N_4804,N_3927,N_4094);
nor U4805 (N_4805,N_4395,N_4025);
xnor U4806 (N_4806,N_4037,N_4257);
xnor U4807 (N_4807,N_4095,N_3924);
xor U4808 (N_4808,N_3950,N_3984);
nor U4809 (N_4809,N_4086,N_4459);
nand U4810 (N_4810,N_4027,N_3997);
xor U4811 (N_4811,N_3829,N_4302);
nor U4812 (N_4812,N_4230,N_4290);
and U4813 (N_4813,N_3978,N_3801);
xnor U4814 (N_4814,N_4255,N_4313);
nor U4815 (N_4815,N_3926,N_4370);
nand U4816 (N_4816,N_4211,N_3914);
nand U4817 (N_4817,N_4147,N_4010);
and U4818 (N_4818,N_4093,N_4220);
nand U4819 (N_4819,N_4156,N_3839);
xor U4820 (N_4820,N_4058,N_4258);
xnor U4821 (N_4821,N_4015,N_4306);
and U4822 (N_4822,N_4050,N_4266);
xnor U4823 (N_4823,N_3936,N_4039);
nand U4824 (N_4824,N_3944,N_3954);
and U4825 (N_4825,N_4293,N_4411);
and U4826 (N_4826,N_3777,N_4122);
nor U4827 (N_4827,N_4460,N_4207);
and U4828 (N_4828,N_4206,N_4238);
nor U4829 (N_4829,N_3945,N_4161);
xor U4830 (N_4830,N_4363,N_3996);
nand U4831 (N_4831,N_3788,N_4254);
xor U4832 (N_4832,N_4486,N_4418);
xnor U4833 (N_4833,N_4107,N_3911);
xor U4834 (N_4834,N_4435,N_4113);
or U4835 (N_4835,N_3769,N_3935);
nor U4836 (N_4836,N_4219,N_4236);
nor U4837 (N_4837,N_4136,N_3886);
xnor U4838 (N_4838,N_4417,N_4470);
nand U4839 (N_4839,N_3915,N_3903);
nor U4840 (N_4840,N_4075,N_4379);
nor U4841 (N_4841,N_3848,N_4398);
nor U4842 (N_4842,N_3877,N_3942);
nor U4843 (N_4843,N_4182,N_4045);
nand U4844 (N_4844,N_3758,N_4497);
nor U4845 (N_4845,N_4410,N_4433);
nand U4846 (N_4846,N_3896,N_3782);
xnor U4847 (N_4847,N_4427,N_4196);
xnor U4848 (N_4848,N_3850,N_4101);
or U4849 (N_4849,N_4012,N_4222);
xnor U4850 (N_4850,N_3947,N_4299);
nand U4851 (N_4851,N_3858,N_4157);
or U4852 (N_4852,N_4143,N_4256);
xor U4853 (N_4853,N_3847,N_4099);
and U4854 (N_4854,N_4475,N_3827);
xnor U4855 (N_4855,N_4160,N_4063);
xnor U4856 (N_4856,N_3867,N_3951);
nor U4857 (N_4857,N_3830,N_4103);
nor U4858 (N_4858,N_4308,N_4268);
or U4859 (N_4859,N_4377,N_4124);
nor U4860 (N_4860,N_3998,N_4205);
or U4861 (N_4861,N_4151,N_4292);
and U4862 (N_4862,N_3807,N_4454);
and U4863 (N_4863,N_4372,N_4330);
xor U4864 (N_4864,N_3941,N_4322);
xor U4865 (N_4865,N_3803,N_4291);
nand U4866 (N_4866,N_3923,N_3754);
or U4867 (N_4867,N_3750,N_4089);
nor U4868 (N_4868,N_4176,N_4128);
nor U4869 (N_4869,N_4447,N_4034);
nor U4870 (N_4870,N_3813,N_4347);
nor U4871 (N_4871,N_3974,N_4318);
xnor U4872 (N_4872,N_4389,N_3838);
nand U4873 (N_4873,N_3845,N_4192);
and U4874 (N_4874,N_3939,N_4202);
xor U4875 (N_4875,N_4138,N_4154);
xor U4876 (N_4876,N_3834,N_3899);
nor U4877 (N_4877,N_4433,N_3999);
nor U4878 (N_4878,N_4101,N_4488);
and U4879 (N_4879,N_4147,N_3987);
nor U4880 (N_4880,N_4203,N_3980);
nor U4881 (N_4881,N_4363,N_4364);
and U4882 (N_4882,N_4055,N_4481);
or U4883 (N_4883,N_4099,N_4410);
or U4884 (N_4884,N_4070,N_4425);
and U4885 (N_4885,N_4371,N_3849);
nor U4886 (N_4886,N_3985,N_3870);
or U4887 (N_4887,N_4289,N_3942);
xnor U4888 (N_4888,N_4063,N_3843);
xnor U4889 (N_4889,N_3976,N_4137);
nand U4890 (N_4890,N_4385,N_3900);
nor U4891 (N_4891,N_3838,N_4138);
or U4892 (N_4892,N_3753,N_4452);
nor U4893 (N_4893,N_4267,N_4172);
or U4894 (N_4894,N_4394,N_4286);
or U4895 (N_4895,N_4370,N_4231);
or U4896 (N_4896,N_4022,N_4016);
nor U4897 (N_4897,N_4354,N_4171);
xnor U4898 (N_4898,N_4033,N_3807);
or U4899 (N_4899,N_3897,N_4309);
nand U4900 (N_4900,N_4462,N_3966);
and U4901 (N_4901,N_3913,N_4352);
nor U4902 (N_4902,N_3994,N_4027);
xnor U4903 (N_4903,N_3926,N_4339);
or U4904 (N_4904,N_3878,N_3945);
xnor U4905 (N_4905,N_4337,N_4019);
and U4906 (N_4906,N_4230,N_4436);
and U4907 (N_4907,N_4302,N_4466);
nor U4908 (N_4908,N_3953,N_3919);
and U4909 (N_4909,N_4161,N_4068);
nand U4910 (N_4910,N_3949,N_4009);
nand U4911 (N_4911,N_3902,N_3900);
or U4912 (N_4912,N_4232,N_4102);
or U4913 (N_4913,N_4467,N_3944);
or U4914 (N_4914,N_4268,N_4203);
nand U4915 (N_4915,N_4371,N_4103);
nand U4916 (N_4916,N_4229,N_4236);
nand U4917 (N_4917,N_4266,N_4238);
nor U4918 (N_4918,N_4191,N_3884);
nand U4919 (N_4919,N_4196,N_4086);
and U4920 (N_4920,N_4080,N_3990);
and U4921 (N_4921,N_4134,N_4428);
xnor U4922 (N_4922,N_4421,N_4036);
and U4923 (N_4923,N_4198,N_3810);
xor U4924 (N_4924,N_3998,N_4432);
nand U4925 (N_4925,N_4484,N_3765);
and U4926 (N_4926,N_4013,N_3866);
and U4927 (N_4927,N_3895,N_4183);
and U4928 (N_4928,N_3961,N_4383);
xor U4929 (N_4929,N_3781,N_4069);
nand U4930 (N_4930,N_4433,N_4191);
or U4931 (N_4931,N_4019,N_4399);
xor U4932 (N_4932,N_4271,N_4058);
nor U4933 (N_4933,N_4143,N_4369);
and U4934 (N_4934,N_4121,N_3949);
xnor U4935 (N_4935,N_3969,N_4096);
nor U4936 (N_4936,N_4048,N_4425);
or U4937 (N_4937,N_3889,N_3935);
and U4938 (N_4938,N_3817,N_4072);
and U4939 (N_4939,N_4498,N_4110);
or U4940 (N_4940,N_3946,N_4220);
nand U4941 (N_4941,N_4424,N_3968);
xor U4942 (N_4942,N_3843,N_4088);
and U4943 (N_4943,N_3861,N_4363);
xnor U4944 (N_4944,N_4283,N_4417);
or U4945 (N_4945,N_4386,N_4323);
nor U4946 (N_4946,N_4196,N_4402);
or U4947 (N_4947,N_3912,N_4332);
nor U4948 (N_4948,N_4054,N_4250);
nand U4949 (N_4949,N_4279,N_4397);
nor U4950 (N_4950,N_4349,N_3849);
nand U4951 (N_4951,N_4170,N_4366);
nand U4952 (N_4952,N_3820,N_4079);
xnor U4953 (N_4953,N_3856,N_4413);
xor U4954 (N_4954,N_4092,N_4432);
nand U4955 (N_4955,N_4014,N_3775);
xor U4956 (N_4956,N_4291,N_4442);
nor U4957 (N_4957,N_3971,N_4448);
nand U4958 (N_4958,N_4393,N_4429);
xnor U4959 (N_4959,N_4411,N_3830);
nand U4960 (N_4960,N_4408,N_4373);
or U4961 (N_4961,N_4049,N_4360);
and U4962 (N_4962,N_4066,N_3860);
and U4963 (N_4963,N_4010,N_4494);
xor U4964 (N_4964,N_4404,N_3795);
xnor U4965 (N_4965,N_3820,N_4269);
nand U4966 (N_4966,N_3789,N_3886);
nor U4967 (N_4967,N_3800,N_4423);
or U4968 (N_4968,N_4092,N_4293);
and U4969 (N_4969,N_3997,N_4292);
and U4970 (N_4970,N_4020,N_3818);
xnor U4971 (N_4971,N_4391,N_4086);
xnor U4972 (N_4972,N_4468,N_4311);
or U4973 (N_4973,N_3916,N_3857);
and U4974 (N_4974,N_4248,N_3830);
or U4975 (N_4975,N_4153,N_4060);
nand U4976 (N_4976,N_4028,N_4483);
nor U4977 (N_4977,N_3820,N_3981);
xnor U4978 (N_4978,N_4259,N_3784);
and U4979 (N_4979,N_4212,N_4018);
and U4980 (N_4980,N_3819,N_4497);
nor U4981 (N_4981,N_3875,N_4088);
nor U4982 (N_4982,N_4393,N_4074);
or U4983 (N_4983,N_4252,N_4460);
or U4984 (N_4984,N_4338,N_4112);
and U4985 (N_4985,N_4360,N_3816);
xnor U4986 (N_4986,N_3995,N_4282);
and U4987 (N_4987,N_4020,N_4402);
and U4988 (N_4988,N_4042,N_3782);
nand U4989 (N_4989,N_3904,N_4107);
xor U4990 (N_4990,N_4153,N_3912);
nand U4991 (N_4991,N_4122,N_3832);
nand U4992 (N_4992,N_4075,N_4314);
nor U4993 (N_4993,N_4467,N_4023);
xnor U4994 (N_4994,N_3886,N_4288);
and U4995 (N_4995,N_4405,N_3992);
and U4996 (N_4996,N_4089,N_4484);
or U4997 (N_4997,N_4218,N_3827);
and U4998 (N_4998,N_3880,N_4145);
and U4999 (N_4999,N_4396,N_4498);
nor U5000 (N_5000,N_4378,N_3987);
nor U5001 (N_5001,N_4071,N_3787);
or U5002 (N_5002,N_3861,N_4453);
or U5003 (N_5003,N_4488,N_4448);
nor U5004 (N_5004,N_3902,N_4164);
xor U5005 (N_5005,N_4399,N_4468);
xor U5006 (N_5006,N_4153,N_4431);
xnor U5007 (N_5007,N_3976,N_3903);
xnor U5008 (N_5008,N_4070,N_3958);
and U5009 (N_5009,N_3882,N_3788);
and U5010 (N_5010,N_4132,N_4133);
nor U5011 (N_5011,N_4237,N_3767);
nor U5012 (N_5012,N_4080,N_3975);
nand U5013 (N_5013,N_3930,N_4241);
nor U5014 (N_5014,N_4371,N_3936);
and U5015 (N_5015,N_4184,N_4413);
xor U5016 (N_5016,N_4116,N_4243);
xor U5017 (N_5017,N_3923,N_4151);
nand U5018 (N_5018,N_3987,N_4486);
or U5019 (N_5019,N_4401,N_3833);
and U5020 (N_5020,N_4244,N_3767);
and U5021 (N_5021,N_3878,N_4336);
xor U5022 (N_5022,N_3769,N_4396);
or U5023 (N_5023,N_4159,N_4016);
or U5024 (N_5024,N_4019,N_4464);
or U5025 (N_5025,N_4214,N_3858);
xor U5026 (N_5026,N_4070,N_4228);
or U5027 (N_5027,N_4057,N_4343);
and U5028 (N_5028,N_3963,N_3995);
or U5029 (N_5029,N_4398,N_4279);
nand U5030 (N_5030,N_4056,N_4070);
xnor U5031 (N_5031,N_4127,N_4486);
and U5032 (N_5032,N_3780,N_4077);
nor U5033 (N_5033,N_4307,N_4283);
nand U5034 (N_5034,N_4027,N_3766);
nand U5035 (N_5035,N_3810,N_3930);
or U5036 (N_5036,N_4491,N_4071);
or U5037 (N_5037,N_4091,N_4037);
and U5038 (N_5038,N_4149,N_4418);
nor U5039 (N_5039,N_3785,N_3838);
nor U5040 (N_5040,N_4254,N_4066);
and U5041 (N_5041,N_3979,N_3778);
and U5042 (N_5042,N_4055,N_4253);
or U5043 (N_5043,N_4121,N_4253);
and U5044 (N_5044,N_4322,N_4013);
nor U5045 (N_5045,N_4002,N_4407);
and U5046 (N_5046,N_4334,N_4222);
or U5047 (N_5047,N_3975,N_3891);
nor U5048 (N_5048,N_4201,N_3985);
xor U5049 (N_5049,N_3893,N_4238);
and U5050 (N_5050,N_3979,N_4042);
nand U5051 (N_5051,N_3959,N_4225);
or U5052 (N_5052,N_4434,N_3814);
xnor U5053 (N_5053,N_4192,N_3863);
and U5054 (N_5054,N_3898,N_4261);
or U5055 (N_5055,N_4225,N_3901);
nand U5056 (N_5056,N_4217,N_4208);
xnor U5057 (N_5057,N_4133,N_4233);
nor U5058 (N_5058,N_4366,N_4125);
nand U5059 (N_5059,N_3778,N_4324);
nand U5060 (N_5060,N_4420,N_4230);
or U5061 (N_5061,N_4198,N_4463);
or U5062 (N_5062,N_4370,N_4298);
nor U5063 (N_5063,N_4204,N_3950);
nor U5064 (N_5064,N_4081,N_3999);
nor U5065 (N_5065,N_4232,N_4313);
nor U5066 (N_5066,N_3947,N_3974);
xnor U5067 (N_5067,N_4167,N_4479);
nand U5068 (N_5068,N_4450,N_3783);
and U5069 (N_5069,N_4051,N_4207);
nor U5070 (N_5070,N_4414,N_4225);
or U5071 (N_5071,N_4349,N_4299);
xnor U5072 (N_5072,N_4218,N_3871);
xor U5073 (N_5073,N_3799,N_4443);
xnor U5074 (N_5074,N_4047,N_3788);
xnor U5075 (N_5075,N_4239,N_4104);
and U5076 (N_5076,N_4253,N_4496);
or U5077 (N_5077,N_4492,N_4052);
or U5078 (N_5078,N_4438,N_4148);
xor U5079 (N_5079,N_4284,N_4067);
nor U5080 (N_5080,N_4312,N_4129);
or U5081 (N_5081,N_3961,N_3758);
or U5082 (N_5082,N_3757,N_3968);
and U5083 (N_5083,N_4236,N_4053);
nand U5084 (N_5084,N_3909,N_4115);
xnor U5085 (N_5085,N_4044,N_4329);
and U5086 (N_5086,N_4380,N_4401);
xnor U5087 (N_5087,N_4332,N_4102);
nand U5088 (N_5088,N_3880,N_3983);
xor U5089 (N_5089,N_3789,N_4466);
or U5090 (N_5090,N_3819,N_4241);
and U5091 (N_5091,N_4159,N_4173);
nor U5092 (N_5092,N_4103,N_4076);
nor U5093 (N_5093,N_4118,N_3941);
and U5094 (N_5094,N_4378,N_3992);
xnor U5095 (N_5095,N_4142,N_3854);
nor U5096 (N_5096,N_4105,N_4344);
nor U5097 (N_5097,N_3789,N_4094);
nand U5098 (N_5098,N_4223,N_4332);
xnor U5099 (N_5099,N_3883,N_4296);
or U5100 (N_5100,N_4429,N_4121);
nor U5101 (N_5101,N_4130,N_4317);
nor U5102 (N_5102,N_3868,N_4351);
and U5103 (N_5103,N_3825,N_4150);
or U5104 (N_5104,N_4416,N_3858);
xnor U5105 (N_5105,N_3755,N_3775);
xnor U5106 (N_5106,N_4097,N_4018);
xnor U5107 (N_5107,N_3838,N_4467);
and U5108 (N_5108,N_4356,N_4136);
nor U5109 (N_5109,N_4421,N_3899);
xnor U5110 (N_5110,N_4118,N_4176);
xor U5111 (N_5111,N_3956,N_4209);
and U5112 (N_5112,N_3853,N_4140);
nor U5113 (N_5113,N_4288,N_4467);
xnor U5114 (N_5114,N_3962,N_4392);
nor U5115 (N_5115,N_4136,N_4405);
nor U5116 (N_5116,N_3824,N_4493);
or U5117 (N_5117,N_4160,N_4096);
nand U5118 (N_5118,N_4021,N_3878);
nor U5119 (N_5119,N_3953,N_3853);
or U5120 (N_5120,N_3769,N_4224);
xor U5121 (N_5121,N_4478,N_4375);
nor U5122 (N_5122,N_4111,N_4190);
xor U5123 (N_5123,N_4468,N_3887);
nand U5124 (N_5124,N_4178,N_4254);
or U5125 (N_5125,N_3776,N_4218);
and U5126 (N_5126,N_4367,N_3852);
nand U5127 (N_5127,N_4377,N_4497);
nor U5128 (N_5128,N_4130,N_4410);
nor U5129 (N_5129,N_4291,N_3956);
xor U5130 (N_5130,N_4306,N_4307);
and U5131 (N_5131,N_3789,N_4398);
nand U5132 (N_5132,N_4429,N_4480);
nand U5133 (N_5133,N_3785,N_3946);
nand U5134 (N_5134,N_3751,N_4498);
nand U5135 (N_5135,N_4198,N_3837);
and U5136 (N_5136,N_4188,N_4057);
nand U5137 (N_5137,N_3868,N_4269);
and U5138 (N_5138,N_4111,N_3802);
and U5139 (N_5139,N_4048,N_4321);
xnor U5140 (N_5140,N_4271,N_3937);
nand U5141 (N_5141,N_4039,N_3817);
xor U5142 (N_5142,N_4395,N_4440);
and U5143 (N_5143,N_4043,N_4241);
nor U5144 (N_5144,N_3894,N_3797);
nand U5145 (N_5145,N_4033,N_4389);
and U5146 (N_5146,N_4179,N_4186);
xnor U5147 (N_5147,N_3872,N_3796);
xnor U5148 (N_5148,N_4088,N_3750);
nand U5149 (N_5149,N_4027,N_4089);
nand U5150 (N_5150,N_3829,N_4022);
xnor U5151 (N_5151,N_3796,N_4377);
xnor U5152 (N_5152,N_3983,N_4257);
xnor U5153 (N_5153,N_4290,N_3847);
nand U5154 (N_5154,N_3996,N_4125);
and U5155 (N_5155,N_4353,N_4473);
nand U5156 (N_5156,N_3920,N_4363);
and U5157 (N_5157,N_4243,N_4479);
or U5158 (N_5158,N_4133,N_3976);
nand U5159 (N_5159,N_4465,N_3987);
nand U5160 (N_5160,N_4253,N_4441);
nor U5161 (N_5161,N_4033,N_4489);
or U5162 (N_5162,N_3966,N_4206);
xnor U5163 (N_5163,N_3788,N_4352);
nor U5164 (N_5164,N_4159,N_4116);
nor U5165 (N_5165,N_4079,N_3795);
nor U5166 (N_5166,N_4106,N_3794);
and U5167 (N_5167,N_4418,N_4440);
nor U5168 (N_5168,N_4454,N_4374);
nor U5169 (N_5169,N_3969,N_4117);
nor U5170 (N_5170,N_3883,N_3878);
xnor U5171 (N_5171,N_4481,N_4053);
nor U5172 (N_5172,N_3840,N_4261);
or U5173 (N_5173,N_3902,N_3828);
nor U5174 (N_5174,N_3957,N_3797);
xor U5175 (N_5175,N_4104,N_3979);
and U5176 (N_5176,N_4215,N_4033);
nor U5177 (N_5177,N_4302,N_3936);
xor U5178 (N_5178,N_3956,N_3815);
or U5179 (N_5179,N_4084,N_3787);
and U5180 (N_5180,N_4096,N_4036);
and U5181 (N_5181,N_4419,N_4055);
nand U5182 (N_5182,N_4094,N_4335);
or U5183 (N_5183,N_3932,N_4301);
nor U5184 (N_5184,N_4391,N_4084);
or U5185 (N_5185,N_3791,N_3886);
nor U5186 (N_5186,N_4360,N_3876);
and U5187 (N_5187,N_3775,N_4330);
xor U5188 (N_5188,N_3929,N_4296);
or U5189 (N_5189,N_4082,N_4392);
nor U5190 (N_5190,N_3832,N_4368);
nand U5191 (N_5191,N_4052,N_4361);
xnor U5192 (N_5192,N_4050,N_3816);
and U5193 (N_5193,N_4165,N_4494);
or U5194 (N_5194,N_3768,N_4093);
or U5195 (N_5195,N_4456,N_4485);
and U5196 (N_5196,N_4495,N_3861);
xor U5197 (N_5197,N_4268,N_4470);
nand U5198 (N_5198,N_4432,N_4376);
xor U5199 (N_5199,N_4457,N_4282);
nor U5200 (N_5200,N_3967,N_4185);
nand U5201 (N_5201,N_3770,N_4266);
nor U5202 (N_5202,N_3973,N_4058);
xor U5203 (N_5203,N_4401,N_4156);
or U5204 (N_5204,N_4416,N_4410);
nor U5205 (N_5205,N_3799,N_4492);
or U5206 (N_5206,N_4104,N_4309);
or U5207 (N_5207,N_4127,N_4340);
or U5208 (N_5208,N_4058,N_3955);
and U5209 (N_5209,N_4197,N_3833);
nand U5210 (N_5210,N_4441,N_4186);
nand U5211 (N_5211,N_3895,N_4488);
xor U5212 (N_5212,N_4029,N_4348);
xnor U5213 (N_5213,N_3771,N_4065);
nor U5214 (N_5214,N_3774,N_4158);
and U5215 (N_5215,N_4499,N_3913);
nand U5216 (N_5216,N_4480,N_4392);
or U5217 (N_5217,N_4152,N_3896);
xnor U5218 (N_5218,N_4444,N_3776);
nor U5219 (N_5219,N_4200,N_4299);
nor U5220 (N_5220,N_4005,N_4398);
and U5221 (N_5221,N_4070,N_4232);
and U5222 (N_5222,N_4256,N_4254);
and U5223 (N_5223,N_4175,N_3871);
or U5224 (N_5224,N_4280,N_3955);
nand U5225 (N_5225,N_4088,N_4447);
and U5226 (N_5226,N_3952,N_4012);
and U5227 (N_5227,N_4421,N_4129);
and U5228 (N_5228,N_3903,N_4289);
nor U5229 (N_5229,N_3818,N_4067);
nor U5230 (N_5230,N_4233,N_4209);
nor U5231 (N_5231,N_4039,N_4221);
or U5232 (N_5232,N_4141,N_3975);
and U5233 (N_5233,N_3896,N_4257);
nor U5234 (N_5234,N_3838,N_4448);
and U5235 (N_5235,N_4465,N_3835);
nor U5236 (N_5236,N_3847,N_4080);
nand U5237 (N_5237,N_4212,N_3991);
or U5238 (N_5238,N_3816,N_4237);
nor U5239 (N_5239,N_4426,N_4165);
or U5240 (N_5240,N_4048,N_3818);
and U5241 (N_5241,N_4240,N_3932);
and U5242 (N_5242,N_4489,N_3909);
nand U5243 (N_5243,N_3984,N_4126);
and U5244 (N_5244,N_4396,N_4370);
xor U5245 (N_5245,N_4482,N_4031);
nand U5246 (N_5246,N_3996,N_4231);
or U5247 (N_5247,N_4286,N_4154);
and U5248 (N_5248,N_4049,N_4096);
nand U5249 (N_5249,N_4338,N_3780);
nand U5250 (N_5250,N_4705,N_4567);
nand U5251 (N_5251,N_4847,N_5126);
xor U5252 (N_5252,N_4791,N_4700);
and U5253 (N_5253,N_5020,N_4608);
xor U5254 (N_5254,N_4856,N_5242);
nor U5255 (N_5255,N_5140,N_4910);
xor U5256 (N_5256,N_4882,N_4514);
or U5257 (N_5257,N_4649,N_4616);
nand U5258 (N_5258,N_4613,N_5154);
xor U5259 (N_5259,N_4899,N_4891);
xnor U5260 (N_5260,N_4667,N_5151);
or U5261 (N_5261,N_4530,N_4892);
and U5262 (N_5262,N_5162,N_5106);
or U5263 (N_5263,N_5194,N_5215);
nand U5264 (N_5264,N_4963,N_4872);
or U5265 (N_5265,N_5229,N_5023);
nor U5266 (N_5266,N_5089,N_5227);
nor U5267 (N_5267,N_4636,N_5116);
and U5268 (N_5268,N_5193,N_4935);
xor U5269 (N_5269,N_4796,N_5067);
nor U5270 (N_5270,N_5238,N_4846);
and U5271 (N_5271,N_5223,N_5021);
xnor U5272 (N_5272,N_5121,N_4993);
nor U5273 (N_5273,N_4744,N_5143);
or U5274 (N_5274,N_5006,N_4527);
nand U5275 (N_5275,N_4546,N_5038);
or U5276 (N_5276,N_4715,N_4591);
or U5277 (N_5277,N_5137,N_4536);
and U5278 (N_5278,N_4507,N_5178);
nor U5279 (N_5279,N_4956,N_5214);
nor U5280 (N_5280,N_5171,N_4834);
or U5281 (N_5281,N_4721,N_4586);
nand U5282 (N_5282,N_4980,N_4720);
xor U5283 (N_5283,N_4742,N_4875);
and U5284 (N_5284,N_4917,N_4642);
and U5285 (N_5285,N_5108,N_4535);
nor U5286 (N_5286,N_4688,N_5192);
xor U5287 (N_5287,N_4881,N_5002);
and U5288 (N_5288,N_4752,N_5198);
xnor U5289 (N_5289,N_5147,N_4533);
xor U5290 (N_5290,N_4756,N_5197);
nand U5291 (N_5291,N_4785,N_4502);
nand U5292 (N_5292,N_4585,N_4578);
or U5293 (N_5293,N_4548,N_4988);
nor U5294 (N_5294,N_4515,N_5012);
xnor U5295 (N_5295,N_5186,N_4840);
xnor U5296 (N_5296,N_4692,N_4580);
nand U5297 (N_5297,N_4866,N_5034);
nor U5298 (N_5298,N_4898,N_4685);
nor U5299 (N_5299,N_4985,N_4628);
nor U5300 (N_5300,N_5201,N_5245);
and U5301 (N_5301,N_5249,N_4900);
xor U5302 (N_5302,N_5015,N_4661);
xor U5303 (N_5303,N_4851,N_4664);
and U5304 (N_5304,N_4886,N_4594);
nand U5305 (N_5305,N_4629,N_4707);
xor U5306 (N_5306,N_5248,N_4979);
and U5307 (N_5307,N_4562,N_5246);
or U5308 (N_5308,N_4965,N_5000);
or U5309 (N_5309,N_4815,N_4506);
nand U5310 (N_5310,N_4560,N_4644);
xnor U5311 (N_5311,N_5217,N_4942);
and U5312 (N_5312,N_4767,N_5155);
and U5313 (N_5313,N_5085,N_5101);
xor U5314 (N_5314,N_4769,N_4532);
xnor U5315 (N_5315,N_5014,N_5185);
nor U5316 (N_5316,N_5232,N_4758);
nand U5317 (N_5317,N_4571,N_5141);
nand U5318 (N_5318,N_4699,N_5160);
or U5319 (N_5319,N_4920,N_4686);
nor U5320 (N_5320,N_4836,N_4939);
xor U5321 (N_5321,N_5093,N_4736);
xor U5322 (N_5322,N_5063,N_5124);
xor U5323 (N_5323,N_4682,N_5043);
or U5324 (N_5324,N_4782,N_4668);
or U5325 (N_5325,N_4503,N_5174);
xnor U5326 (N_5326,N_5061,N_4788);
nor U5327 (N_5327,N_4549,N_4734);
or U5328 (N_5328,N_4967,N_5173);
nand U5329 (N_5329,N_5059,N_5090);
nand U5330 (N_5330,N_4635,N_4870);
and U5331 (N_5331,N_4849,N_4820);
xnor U5332 (N_5332,N_5247,N_5142);
nand U5333 (N_5333,N_4839,N_4755);
xnor U5334 (N_5334,N_5071,N_4821);
or U5335 (N_5335,N_4648,N_4805);
or U5336 (N_5336,N_4990,N_4584);
nor U5337 (N_5337,N_4991,N_4934);
and U5338 (N_5338,N_4932,N_4867);
nor U5339 (N_5339,N_4669,N_4841);
and U5340 (N_5340,N_5184,N_4904);
and U5341 (N_5341,N_4772,N_4714);
and U5342 (N_5342,N_4780,N_5136);
nor U5343 (N_5343,N_4727,N_4654);
or U5344 (N_5344,N_4986,N_4610);
xnor U5345 (N_5345,N_5019,N_4812);
or U5346 (N_5346,N_5138,N_4869);
nor U5347 (N_5347,N_5207,N_4638);
nand U5348 (N_5348,N_5199,N_5026);
xnor U5349 (N_5349,N_4749,N_4798);
or U5350 (N_5350,N_4764,N_4831);
nand U5351 (N_5351,N_5001,N_4880);
and U5352 (N_5352,N_4529,N_4592);
nand U5353 (N_5353,N_4808,N_5112);
xnor U5354 (N_5354,N_5008,N_5131);
and U5355 (N_5355,N_5128,N_4574);
nand U5356 (N_5356,N_4510,N_4770);
xnor U5357 (N_5357,N_4746,N_4633);
xor U5358 (N_5358,N_4912,N_4662);
or U5359 (N_5359,N_5132,N_4916);
and U5360 (N_5360,N_5177,N_5045);
xor U5361 (N_5361,N_4542,N_5092);
xor U5362 (N_5362,N_4620,N_4861);
nor U5363 (N_5363,N_4864,N_5161);
nand U5364 (N_5364,N_4826,N_5225);
nor U5365 (N_5365,N_4651,N_5159);
nand U5366 (N_5366,N_4817,N_4745);
and U5367 (N_5367,N_4717,N_4862);
and U5368 (N_5368,N_4829,N_4564);
nor U5369 (N_5369,N_4550,N_4858);
xnor U5370 (N_5370,N_5097,N_4865);
or U5371 (N_5371,N_4948,N_4823);
or U5372 (N_5372,N_4725,N_5125);
or U5373 (N_5373,N_4885,N_4773);
and U5374 (N_5374,N_4655,N_4809);
or U5375 (N_5375,N_5163,N_4924);
nand U5376 (N_5376,N_4587,N_4652);
xnor U5377 (N_5377,N_4978,N_4959);
xor U5378 (N_5378,N_4630,N_4656);
and U5379 (N_5379,N_4697,N_4719);
and U5380 (N_5380,N_4539,N_4940);
nand U5381 (N_5381,N_4905,N_5230);
or U5382 (N_5382,N_5050,N_4771);
xnor U5383 (N_5383,N_5057,N_5176);
nor U5384 (N_5384,N_4973,N_5032);
nand U5385 (N_5385,N_5172,N_4810);
or U5386 (N_5386,N_4952,N_5072);
nor U5387 (N_5387,N_4807,N_4625);
nand U5388 (N_5388,N_4671,N_4643);
xnor U5389 (N_5389,N_4997,N_5139);
nor U5390 (N_5390,N_4602,N_4653);
xnor U5391 (N_5391,N_5118,N_4879);
or U5392 (N_5392,N_5129,N_4680);
xnor U5393 (N_5393,N_5127,N_4888);
nand U5394 (N_5394,N_4894,N_4619);
nand U5395 (N_5395,N_5190,N_4624);
xor U5396 (N_5396,N_5158,N_4518);
xnor U5397 (N_5397,N_4737,N_5111);
nand U5398 (N_5398,N_4657,N_4766);
nand U5399 (N_5399,N_4974,N_4803);
nor U5400 (N_5400,N_5028,N_5119);
and U5401 (N_5401,N_5224,N_4738);
and U5402 (N_5402,N_4728,N_4789);
nand U5403 (N_5403,N_5054,N_4541);
xor U5404 (N_5404,N_4603,N_4696);
or U5405 (N_5405,N_4976,N_4666);
and U5406 (N_5406,N_4525,N_5003);
or U5407 (N_5407,N_4576,N_4612);
nor U5408 (N_5408,N_4845,N_4750);
nand U5409 (N_5409,N_4936,N_4950);
nand U5410 (N_5410,N_4555,N_4762);
and U5411 (N_5411,N_4921,N_4601);
nand U5412 (N_5412,N_5146,N_4693);
or U5413 (N_5413,N_4957,N_5035);
or U5414 (N_5414,N_4724,N_4855);
nand U5415 (N_5415,N_4683,N_4768);
nand U5416 (N_5416,N_5135,N_4739);
nand U5417 (N_5417,N_5243,N_4922);
or U5418 (N_5418,N_4645,N_4961);
xor U5419 (N_5419,N_4844,N_5188);
xor U5420 (N_5420,N_4689,N_4994);
and U5421 (N_5421,N_4835,N_5213);
xnor U5422 (N_5422,N_5216,N_4828);
nor U5423 (N_5423,N_4672,N_4595);
xnor U5424 (N_5424,N_4557,N_4981);
and U5425 (N_5425,N_4568,N_5182);
and U5426 (N_5426,N_4675,N_5080);
nand U5427 (N_5427,N_4837,N_4678);
and U5428 (N_5428,N_4614,N_4799);
nor U5429 (N_5429,N_4729,N_4704);
nor U5430 (N_5430,N_4786,N_5009);
or U5431 (N_5431,N_4964,N_5181);
and U5432 (N_5432,N_5191,N_4713);
nand U5433 (N_5433,N_4969,N_4760);
nand U5434 (N_5434,N_4824,N_5123);
or U5435 (N_5435,N_4565,N_4853);
or U5436 (N_5436,N_5025,N_4813);
nand U5437 (N_5437,N_4923,N_4926);
nand U5438 (N_5438,N_4660,N_4908);
or U5439 (N_5439,N_4524,N_4972);
and U5440 (N_5440,N_4761,N_5168);
and U5441 (N_5441,N_5235,N_4871);
and U5442 (N_5442,N_4694,N_4901);
xnor U5443 (N_5443,N_4522,N_5088);
xnor U5444 (N_5444,N_5079,N_4622);
or U5445 (N_5445,N_4984,N_4534);
or U5446 (N_5446,N_4702,N_4606);
xor U5447 (N_5447,N_4779,N_5029);
xor U5448 (N_5448,N_5078,N_5204);
xnor U5449 (N_5449,N_4735,N_4795);
and U5450 (N_5450,N_4511,N_5148);
nand U5451 (N_5451,N_5244,N_4609);
nand U5452 (N_5452,N_5104,N_4968);
or U5453 (N_5453,N_4520,N_4623);
nor U5454 (N_5454,N_4695,N_4552);
or U5455 (N_5455,N_5237,N_4516);
xnor U5456 (N_5456,N_4822,N_4763);
nand U5457 (N_5457,N_5145,N_5031);
nand U5458 (N_5458,N_4505,N_4572);
or U5459 (N_5459,N_5157,N_4777);
nor U5460 (N_5460,N_5110,N_4998);
nor U5461 (N_5461,N_4816,N_4982);
xnor U5462 (N_5462,N_5099,N_4521);
xnor U5463 (N_5463,N_5165,N_5241);
or U5464 (N_5464,N_5070,N_4741);
nand U5465 (N_5465,N_5222,N_4600);
xnor U5466 (N_5466,N_4759,N_4679);
and U5467 (N_5467,N_4597,N_5076);
nor U5468 (N_5468,N_4605,N_5010);
and U5469 (N_5469,N_5109,N_5098);
nand U5470 (N_5470,N_4819,N_5056);
nand U5471 (N_5471,N_4793,N_5047);
and U5472 (N_5472,N_4588,N_4911);
and U5473 (N_5473,N_4556,N_4599);
xnor U5474 (N_5474,N_4850,N_4748);
nor U5475 (N_5475,N_4537,N_4566);
nor U5476 (N_5476,N_4709,N_4838);
xor U5477 (N_5477,N_4690,N_4723);
nor U5478 (N_5478,N_5037,N_4833);
or U5479 (N_5479,N_5024,N_4797);
nor U5480 (N_5480,N_4698,N_5081);
nor U5481 (N_5481,N_4999,N_5183);
and U5482 (N_5482,N_4787,N_4681);
nand U5483 (N_5483,N_4913,N_4887);
nor U5484 (N_5484,N_5042,N_4611);
or U5485 (N_5485,N_4958,N_4531);
or U5486 (N_5486,N_5120,N_4800);
nor U5487 (N_5487,N_4801,N_4674);
and U5488 (N_5488,N_5226,N_4883);
and U5489 (N_5489,N_4776,N_4977);
nand U5490 (N_5490,N_4765,N_4554);
nand U5491 (N_5491,N_5004,N_5196);
xor U5492 (N_5492,N_4670,N_4955);
nand U5493 (N_5493,N_4874,N_5169);
nor U5494 (N_5494,N_4589,N_4684);
and U5495 (N_5495,N_4931,N_4832);
and U5496 (N_5496,N_5134,N_5150);
nand U5497 (N_5497,N_4551,N_5086);
nor U5498 (N_5498,N_4778,N_4747);
and U5499 (N_5499,N_4711,N_5077);
nand U5500 (N_5500,N_5044,N_4579);
or U5501 (N_5501,N_4582,N_4914);
or U5502 (N_5502,N_4848,N_4553);
and U5503 (N_5503,N_4621,N_5187);
xor U5504 (N_5504,N_5144,N_5007);
nor U5505 (N_5505,N_4631,N_4583);
nor U5506 (N_5506,N_4509,N_4540);
nor U5507 (N_5507,N_4634,N_5113);
nand U5508 (N_5508,N_4665,N_4966);
and U5509 (N_5509,N_4953,N_5164);
nor U5510 (N_5510,N_4938,N_4941);
xor U5511 (N_5511,N_5107,N_5049);
or U5512 (N_5512,N_5065,N_4962);
and U5513 (N_5513,N_4889,N_4607);
or U5514 (N_5514,N_4730,N_5209);
nand U5515 (N_5515,N_5195,N_4732);
nor U5516 (N_5516,N_4944,N_4712);
or U5517 (N_5517,N_4868,N_5091);
nand U5518 (N_5518,N_4946,N_4854);
nor U5519 (N_5519,N_4995,N_5220);
or U5520 (N_5520,N_5064,N_4740);
xor U5521 (N_5521,N_4877,N_5022);
nand U5522 (N_5522,N_4701,N_4570);
and U5523 (N_5523,N_5100,N_5211);
and U5524 (N_5524,N_4508,N_4577);
nand U5525 (N_5525,N_5152,N_4909);
or U5526 (N_5526,N_5203,N_4641);
nand U5527 (N_5527,N_5221,N_5005);
or U5528 (N_5528,N_4863,N_5033);
xor U5529 (N_5529,N_5218,N_4890);
and U5530 (N_5530,N_5102,N_5036);
and U5531 (N_5531,N_5200,N_4703);
xnor U5532 (N_5532,N_4663,N_4673);
nor U5533 (N_5533,N_5219,N_4647);
and U5534 (N_5534,N_4658,N_5170);
and U5535 (N_5535,N_5069,N_4627);
nor U5536 (N_5536,N_4757,N_4519);
nand U5537 (N_5537,N_4830,N_4859);
or U5538 (N_5538,N_5094,N_4708);
nand U5539 (N_5539,N_5017,N_4929);
xnor U5540 (N_5540,N_5130,N_5013);
nor U5541 (N_5541,N_4784,N_4987);
or U5542 (N_5542,N_5096,N_4563);
and U5543 (N_5543,N_4639,N_4646);
and U5544 (N_5544,N_5060,N_4852);
and U5545 (N_5545,N_5048,N_5040);
xnor U5546 (N_5546,N_4512,N_5073);
xor U5547 (N_5547,N_4706,N_4632);
xor U5548 (N_5548,N_5156,N_4504);
nor U5549 (N_5549,N_4794,N_4650);
xnor U5550 (N_5550,N_4501,N_5153);
xnor U5551 (N_5551,N_4975,N_5122);
nand U5552 (N_5552,N_4945,N_4878);
and U5553 (N_5553,N_4558,N_4710);
xor U5554 (N_5554,N_5114,N_4500);
nand U5555 (N_5555,N_4513,N_4754);
and U5556 (N_5556,N_5117,N_5205);
xnor U5557 (N_5557,N_4543,N_4691);
or U5558 (N_5558,N_5208,N_5236);
xor U5559 (N_5559,N_4726,N_5231);
and U5560 (N_5560,N_5175,N_4718);
xor U5561 (N_5561,N_4893,N_4598);
nor U5562 (N_5562,N_5083,N_4743);
nor U5563 (N_5563,N_4617,N_4903);
xnor U5564 (N_5564,N_4559,N_5068);
nand U5565 (N_5565,N_5212,N_4811);
and U5566 (N_5566,N_4989,N_5041);
nor U5567 (N_5567,N_5051,N_4676);
nor U5568 (N_5568,N_5053,N_4753);
and U5569 (N_5569,N_5055,N_4896);
nand U5570 (N_5570,N_4925,N_4781);
and U5571 (N_5571,N_4604,N_5052);
and U5572 (N_5572,N_4971,N_5084);
and U5573 (N_5573,N_4895,N_4884);
and U5574 (N_5574,N_4774,N_5234);
and U5575 (N_5575,N_4951,N_4722);
xnor U5576 (N_5576,N_5228,N_5239);
and U5577 (N_5577,N_4783,N_5103);
or U5578 (N_5578,N_4937,N_4927);
or U5579 (N_5579,N_4915,N_4897);
or U5580 (N_5580,N_5074,N_5027);
nand U5581 (N_5581,N_4873,N_5189);
nor U5582 (N_5582,N_4640,N_4569);
nor U5583 (N_5583,N_4545,N_5240);
nand U5584 (N_5584,N_4677,N_4590);
or U5585 (N_5585,N_4907,N_5058);
and U5586 (N_5586,N_4528,N_4538);
or U5587 (N_5587,N_4790,N_5167);
xor U5588 (N_5588,N_4818,N_4954);
or U5589 (N_5589,N_4996,N_4731);
xor U5590 (N_5590,N_4857,N_4775);
and U5591 (N_5591,N_5018,N_4561);
or U5592 (N_5592,N_4983,N_4716);
or U5593 (N_5593,N_4970,N_5066);
nand U5594 (N_5594,N_4593,N_5039);
or U5595 (N_5595,N_4906,N_5115);
nor U5596 (N_5596,N_5133,N_4876);
nand U5597 (N_5597,N_4947,N_5075);
or U5598 (N_5598,N_4544,N_4827);
xor U5599 (N_5599,N_4547,N_4596);
nand U5600 (N_5600,N_5087,N_4992);
and U5601 (N_5601,N_5210,N_4842);
and U5602 (N_5602,N_4792,N_4618);
nor U5603 (N_5603,N_4751,N_5233);
nor U5604 (N_5604,N_4733,N_4930);
xnor U5605 (N_5605,N_4626,N_5206);
xor U5606 (N_5606,N_4523,N_5030);
xor U5607 (N_5607,N_5166,N_4802);
nand U5608 (N_5608,N_4933,N_4928);
nand U5609 (N_5609,N_5046,N_4615);
or U5610 (N_5610,N_4843,N_4659);
or U5611 (N_5611,N_5062,N_4581);
or U5612 (N_5612,N_4919,N_5202);
nor U5613 (N_5613,N_5180,N_4575);
or U5614 (N_5614,N_4573,N_4943);
xnor U5615 (N_5615,N_4902,N_4526);
nor U5616 (N_5616,N_5105,N_5149);
or U5617 (N_5617,N_4806,N_4804);
and U5618 (N_5618,N_4860,N_5179);
nand U5619 (N_5619,N_5082,N_5016);
xor U5620 (N_5620,N_5095,N_4814);
nor U5621 (N_5621,N_4949,N_4825);
or U5622 (N_5622,N_4918,N_5011);
nor U5623 (N_5623,N_4960,N_4687);
xor U5624 (N_5624,N_4637,N_4517);
xor U5625 (N_5625,N_4898,N_4756);
and U5626 (N_5626,N_4647,N_4753);
or U5627 (N_5627,N_5160,N_4965);
nand U5628 (N_5628,N_4596,N_4810);
or U5629 (N_5629,N_4736,N_4747);
xor U5630 (N_5630,N_5005,N_4846);
and U5631 (N_5631,N_4544,N_4953);
and U5632 (N_5632,N_4812,N_5002);
or U5633 (N_5633,N_4716,N_4808);
and U5634 (N_5634,N_5051,N_4516);
nand U5635 (N_5635,N_4666,N_4871);
nor U5636 (N_5636,N_4990,N_5112);
or U5637 (N_5637,N_4808,N_4885);
and U5638 (N_5638,N_4619,N_4860);
nor U5639 (N_5639,N_4873,N_5203);
and U5640 (N_5640,N_5183,N_5159);
and U5641 (N_5641,N_5217,N_4816);
or U5642 (N_5642,N_5039,N_5046);
nor U5643 (N_5643,N_5152,N_5247);
nor U5644 (N_5644,N_5075,N_4906);
or U5645 (N_5645,N_4527,N_5066);
nor U5646 (N_5646,N_4785,N_4671);
nand U5647 (N_5647,N_5190,N_4803);
and U5648 (N_5648,N_5211,N_5079);
xor U5649 (N_5649,N_4553,N_5229);
xnor U5650 (N_5650,N_5226,N_4970);
and U5651 (N_5651,N_4505,N_5197);
nor U5652 (N_5652,N_5067,N_5174);
or U5653 (N_5653,N_4623,N_5111);
nor U5654 (N_5654,N_5161,N_4598);
or U5655 (N_5655,N_4669,N_4907);
xnor U5656 (N_5656,N_5225,N_4843);
nand U5657 (N_5657,N_5095,N_4818);
xor U5658 (N_5658,N_5193,N_5184);
xnor U5659 (N_5659,N_4770,N_4728);
nor U5660 (N_5660,N_5010,N_5176);
nand U5661 (N_5661,N_4658,N_4953);
nand U5662 (N_5662,N_4853,N_4524);
nor U5663 (N_5663,N_4716,N_5107);
and U5664 (N_5664,N_5131,N_4933);
nor U5665 (N_5665,N_4816,N_5005);
and U5666 (N_5666,N_4608,N_4831);
xnor U5667 (N_5667,N_5184,N_4656);
nor U5668 (N_5668,N_4568,N_4795);
and U5669 (N_5669,N_5168,N_5047);
nand U5670 (N_5670,N_4779,N_4754);
and U5671 (N_5671,N_4556,N_4659);
nand U5672 (N_5672,N_5193,N_4852);
and U5673 (N_5673,N_5006,N_4665);
or U5674 (N_5674,N_5029,N_4696);
xnor U5675 (N_5675,N_4847,N_4930);
nand U5676 (N_5676,N_5173,N_4932);
or U5677 (N_5677,N_4549,N_4766);
nand U5678 (N_5678,N_4921,N_4741);
xnor U5679 (N_5679,N_4615,N_5154);
and U5680 (N_5680,N_4516,N_5227);
nor U5681 (N_5681,N_4820,N_4917);
or U5682 (N_5682,N_5098,N_4860);
xnor U5683 (N_5683,N_5214,N_4616);
nand U5684 (N_5684,N_5160,N_5229);
or U5685 (N_5685,N_4637,N_5092);
and U5686 (N_5686,N_5211,N_5145);
xor U5687 (N_5687,N_5034,N_5175);
nand U5688 (N_5688,N_4669,N_4959);
nor U5689 (N_5689,N_4703,N_4938);
or U5690 (N_5690,N_5147,N_4586);
nand U5691 (N_5691,N_4703,N_5098);
nand U5692 (N_5692,N_4677,N_5163);
nand U5693 (N_5693,N_4508,N_5036);
nor U5694 (N_5694,N_4899,N_4975);
xor U5695 (N_5695,N_4557,N_4521);
and U5696 (N_5696,N_5148,N_4892);
and U5697 (N_5697,N_4750,N_4829);
nor U5698 (N_5698,N_4556,N_5119);
nand U5699 (N_5699,N_5190,N_4527);
and U5700 (N_5700,N_4664,N_5083);
and U5701 (N_5701,N_4679,N_5119);
xor U5702 (N_5702,N_5214,N_4660);
and U5703 (N_5703,N_5229,N_4923);
or U5704 (N_5704,N_4936,N_4858);
nor U5705 (N_5705,N_4724,N_4969);
xor U5706 (N_5706,N_4787,N_5223);
or U5707 (N_5707,N_5245,N_5006);
and U5708 (N_5708,N_4678,N_5027);
or U5709 (N_5709,N_5229,N_4734);
or U5710 (N_5710,N_4758,N_4642);
nand U5711 (N_5711,N_4515,N_4502);
nand U5712 (N_5712,N_4839,N_5155);
xnor U5713 (N_5713,N_4870,N_4921);
nand U5714 (N_5714,N_5015,N_5139);
xnor U5715 (N_5715,N_4887,N_4674);
and U5716 (N_5716,N_4686,N_4598);
and U5717 (N_5717,N_4973,N_4532);
xor U5718 (N_5718,N_5072,N_4883);
nor U5719 (N_5719,N_4768,N_4539);
or U5720 (N_5720,N_4724,N_4999);
nand U5721 (N_5721,N_5093,N_4907);
and U5722 (N_5722,N_4983,N_5142);
nor U5723 (N_5723,N_5081,N_5072);
and U5724 (N_5724,N_4854,N_5109);
xnor U5725 (N_5725,N_4789,N_4619);
or U5726 (N_5726,N_4549,N_4695);
and U5727 (N_5727,N_5154,N_4990);
xnor U5728 (N_5728,N_5057,N_4729);
or U5729 (N_5729,N_5124,N_4936);
or U5730 (N_5730,N_5069,N_4559);
and U5731 (N_5731,N_4981,N_4747);
and U5732 (N_5732,N_4626,N_4596);
nor U5733 (N_5733,N_5118,N_5248);
or U5734 (N_5734,N_5131,N_5232);
xnor U5735 (N_5735,N_4815,N_4832);
nand U5736 (N_5736,N_5077,N_4631);
nand U5737 (N_5737,N_4837,N_5085);
nor U5738 (N_5738,N_4622,N_5156);
nand U5739 (N_5739,N_4740,N_4876);
and U5740 (N_5740,N_4833,N_4966);
or U5741 (N_5741,N_5163,N_4737);
and U5742 (N_5742,N_4808,N_4521);
xor U5743 (N_5743,N_4530,N_4924);
or U5744 (N_5744,N_4928,N_4956);
nor U5745 (N_5745,N_4797,N_4874);
and U5746 (N_5746,N_5211,N_4942);
nand U5747 (N_5747,N_4614,N_4991);
nand U5748 (N_5748,N_4788,N_4603);
and U5749 (N_5749,N_4525,N_4590);
or U5750 (N_5750,N_4714,N_5087);
or U5751 (N_5751,N_4829,N_5059);
or U5752 (N_5752,N_4841,N_4868);
xnor U5753 (N_5753,N_4975,N_4830);
and U5754 (N_5754,N_4928,N_5035);
nand U5755 (N_5755,N_4955,N_4803);
or U5756 (N_5756,N_4609,N_4680);
or U5757 (N_5757,N_4580,N_4962);
nand U5758 (N_5758,N_4695,N_5006);
xor U5759 (N_5759,N_5042,N_4666);
nand U5760 (N_5760,N_4714,N_5225);
and U5761 (N_5761,N_5119,N_4752);
nor U5762 (N_5762,N_4949,N_5052);
and U5763 (N_5763,N_5174,N_4872);
and U5764 (N_5764,N_4833,N_4869);
or U5765 (N_5765,N_4570,N_4698);
xnor U5766 (N_5766,N_4797,N_4562);
or U5767 (N_5767,N_4590,N_4615);
nor U5768 (N_5768,N_4529,N_4582);
and U5769 (N_5769,N_4810,N_5044);
nor U5770 (N_5770,N_5009,N_4959);
and U5771 (N_5771,N_5086,N_4710);
xnor U5772 (N_5772,N_5040,N_4737);
nor U5773 (N_5773,N_4638,N_5218);
xnor U5774 (N_5774,N_4673,N_5188);
nand U5775 (N_5775,N_4775,N_4508);
nor U5776 (N_5776,N_4734,N_5086);
nand U5777 (N_5777,N_4554,N_4501);
nand U5778 (N_5778,N_4868,N_5155);
nand U5779 (N_5779,N_5231,N_4991);
xnor U5780 (N_5780,N_5043,N_4882);
nor U5781 (N_5781,N_4739,N_4946);
xnor U5782 (N_5782,N_4779,N_4737);
xor U5783 (N_5783,N_4508,N_5098);
nand U5784 (N_5784,N_5208,N_4796);
or U5785 (N_5785,N_4784,N_4942);
or U5786 (N_5786,N_5113,N_5242);
xor U5787 (N_5787,N_4648,N_5002);
and U5788 (N_5788,N_4845,N_4897);
or U5789 (N_5789,N_4520,N_5071);
or U5790 (N_5790,N_4629,N_4897);
and U5791 (N_5791,N_4967,N_4776);
nor U5792 (N_5792,N_5057,N_4529);
xnor U5793 (N_5793,N_5103,N_4974);
and U5794 (N_5794,N_4767,N_4886);
or U5795 (N_5795,N_4638,N_4635);
or U5796 (N_5796,N_5199,N_4814);
and U5797 (N_5797,N_5194,N_5136);
nand U5798 (N_5798,N_4939,N_5214);
or U5799 (N_5799,N_5227,N_5109);
xor U5800 (N_5800,N_5126,N_4709);
xnor U5801 (N_5801,N_4535,N_4511);
and U5802 (N_5802,N_5228,N_5130);
xnor U5803 (N_5803,N_4561,N_4951);
or U5804 (N_5804,N_5033,N_4518);
and U5805 (N_5805,N_4580,N_4691);
and U5806 (N_5806,N_4888,N_5198);
xnor U5807 (N_5807,N_4891,N_4518);
or U5808 (N_5808,N_4517,N_5148);
nor U5809 (N_5809,N_4813,N_5188);
nor U5810 (N_5810,N_5227,N_5033);
and U5811 (N_5811,N_4846,N_5050);
and U5812 (N_5812,N_4584,N_4901);
xnor U5813 (N_5813,N_4788,N_4683);
nor U5814 (N_5814,N_5044,N_4785);
or U5815 (N_5815,N_5225,N_4950);
nor U5816 (N_5816,N_4723,N_5131);
and U5817 (N_5817,N_4873,N_5178);
and U5818 (N_5818,N_4779,N_4871);
and U5819 (N_5819,N_4927,N_4760);
xor U5820 (N_5820,N_4766,N_5131);
nand U5821 (N_5821,N_5177,N_4898);
nand U5822 (N_5822,N_4661,N_4907);
and U5823 (N_5823,N_4756,N_4608);
nand U5824 (N_5824,N_4546,N_5155);
nor U5825 (N_5825,N_4755,N_4561);
and U5826 (N_5826,N_4769,N_5223);
nor U5827 (N_5827,N_4902,N_5201);
xor U5828 (N_5828,N_4759,N_4937);
or U5829 (N_5829,N_4944,N_4889);
nor U5830 (N_5830,N_4702,N_5046);
or U5831 (N_5831,N_4752,N_4706);
nand U5832 (N_5832,N_4635,N_4825);
nand U5833 (N_5833,N_4839,N_5088);
and U5834 (N_5834,N_5128,N_4671);
nor U5835 (N_5835,N_5162,N_4996);
nor U5836 (N_5836,N_4841,N_5222);
and U5837 (N_5837,N_4892,N_4924);
and U5838 (N_5838,N_4657,N_4557);
or U5839 (N_5839,N_4632,N_4980);
xor U5840 (N_5840,N_4636,N_5125);
nor U5841 (N_5841,N_5197,N_4513);
xnor U5842 (N_5842,N_4861,N_5029);
nand U5843 (N_5843,N_5138,N_4519);
nor U5844 (N_5844,N_5108,N_5205);
xnor U5845 (N_5845,N_4788,N_4939);
nor U5846 (N_5846,N_5071,N_5173);
xnor U5847 (N_5847,N_5235,N_5154);
or U5848 (N_5848,N_4981,N_4917);
or U5849 (N_5849,N_4872,N_4637);
or U5850 (N_5850,N_4782,N_5244);
and U5851 (N_5851,N_4998,N_5150);
and U5852 (N_5852,N_4719,N_5079);
nor U5853 (N_5853,N_5146,N_4854);
and U5854 (N_5854,N_4903,N_4699);
and U5855 (N_5855,N_5226,N_4625);
or U5856 (N_5856,N_4936,N_4669);
xor U5857 (N_5857,N_4562,N_4618);
nor U5858 (N_5858,N_4897,N_4929);
nor U5859 (N_5859,N_4706,N_4653);
nor U5860 (N_5860,N_4657,N_4800);
nand U5861 (N_5861,N_4939,N_5108);
nor U5862 (N_5862,N_4999,N_4632);
and U5863 (N_5863,N_4875,N_5078);
and U5864 (N_5864,N_4966,N_4592);
nand U5865 (N_5865,N_4562,N_5138);
and U5866 (N_5866,N_4793,N_4775);
or U5867 (N_5867,N_4619,N_4859);
or U5868 (N_5868,N_4656,N_4875);
nor U5869 (N_5869,N_4909,N_5080);
nor U5870 (N_5870,N_4659,N_4747);
nand U5871 (N_5871,N_4804,N_4768);
and U5872 (N_5872,N_5082,N_5101);
xor U5873 (N_5873,N_4591,N_5058);
nand U5874 (N_5874,N_4595,N_4778);
nand U5875 (N_5875,N_4782,N_4934);
xor U5876 (N_5876,N_4909,N_5121);
nand U5877 (N_5877,N_4521,N_4632);
nand U5878 (N_5878,N_5216,N_5193);
xor U5879 (N_5879,N_4586,N_4898);
and U5880 (N_5880,N_4602,N_4952);
xnor U5881 (N_5881,N_5073,N_4513);
and U5882 (N_5882,N_4823,N_5145);
xor U5883 (N_5883,N_5187,N_5100);
xnor U5884 (N_5884,N_4572,N_4639);
xnor U5885 (N_5885,N_4896,N_4889);
or U5886 (N_5886,N_4734,N_4641);
xnor U5887 (N_5887,N_4805,N_4963);
or U5888 (N_5888,N_4819,N_4974);
xor U5889 (N_5889,N_4618,N_4714);
nand U5890 (N_5890,N_4635,N_4845);
nor U5891 (N_5891,N_4519,N_4973);
nand U5892 (N_5892,N_4602,N_4852);
and U5893 (N_5893,N_4578,N_4948);
nor U5894 (N_5894,N_4722,N_4560);
or U5895 (N_5895,N_4959,N_5051);
or U5896 (N_5896,N_4525,N_5045);
nand U5897 (N_5897,N_4519,N_4713);
nor U5898 (N_5898,N_5215,N_5021);
nor U5899 (N_5899,N_4944,N_4906);
or U5900 (N_5900,N_5187,N_4508);
nor U5901 (N_5901,N_4960,N_5009);
xor U5902 (N_5902,N_4673,N_5120);
nand U5903 (N_5903,N_4631,N_5098);
nor U5904 (N_5904,N_4777,N_5022);
or U5905 (N_5905,N_5166,N_4815);
xor U5906 (N_5906,N_4760,N_4753);
xnor U5907 (N_5907,N_4902,N_5080);
or U5908 (N_5908,N_4540,N_4983);
nor U5909 (N_5909,N_4668,N_4865);
xnor U5910 (N_5910,N_5069,N_4788);
or U5911 (N_5911,N_4729,N_4615);
or U5912 (N_5912,N_5066,N_4729);
nand U5913 (N_5913,N_4997,N_5070);
xnor U5914 (N_5914,N_4949,N_4931);
nor U5915 (N_5915,N_5034,N_5056);
xnor U5916 (N_5916,N_4902,N_5249);
nand U5917 (N_5917,N_5091,N_4948);
or U5918 (N_5918,N_4522,N_4505);
xnor U5919 (N_5919,N_5094,N_4941);
and U5920 (N_5920,N_4561,N_4734);
nor U5921 (N_5921,N_5102,N_4984);
and U5922 (N_5922,N_5116,N_4513);
nand U5923 (N_5923,N_4545,N_5101);
nand U5924 (N_5924,N_4719,N_5160);
or U5925 (N_5925,N_4686,N_5242);
nor U5926 (N_5926,N_5074,N_4542);
and U5927 (N_5927,N_5130,N_5213);
nor U5928 (N_5928,N_5176,N_4912);
nor U5929 (N_5929,N_4876,N_5008);
or U5930 (N_5930,N_5129,N_4912);
and U5931 (N_5931,N_4918,N_5241);
and U5932 (N_5932,N_4884,N_4942);
xor U5933 (N_5933,N_5246,N_4896);
xor U5934 (N_5934,N_4699,N_4669);
xnor U5935 (N_5935,N_4777,N_4523);
and U5936 (N_5936,N_4693,N_5087);
nand U5937 (N_5937,N_5156,N_5023);
nand U5938 (N_5938,N_4562,N_4707);
nand U5939 (N_5939,N_4685,N_5239);
xnor U5940 (N_5940,N_5103,N_4569);
and U5941 (N_5941,N_4879,N_4938);
nor U5942 (N_5942,N_5170,N_5068);
and U5943 (N_5943,N_4929,N_5149);
nor U5944 (N_5944,N_4637,N_4910);
xor U5945 (N_5945,N_4619,N_5056);
nor U5946 (N_5946,N_4754,N_4841);
and U5947 (N_5947,N_5224,N_4995);
or U5948 (N_5948,N_5205,N_5110);
nor U5949 (N_5949,N_4608,N_4802);
nor U5950 (N_5950,N_4675,N_4644);
or U5951 (N_5951,N_5190,N_4747);
nand U5952 (N_5952,N_5227,N_5171);
nor U5953 (N_5953,N_4565,N_5240);
or U5954 (N_5954,N_4991,N_4710);
and U5955 (N_5955,N_5090,N_5041);
xor U5956 (N_5956,N_4760,N_4507);
or U5957 (N_5957,N_5217,N_4676);
nand U5958 (N_5958,N_5057,N_5119);
and U5959 (N_5959,N_5068,N_4821);
nor U5960 (N_5960,N_5213,N_4794);
nor U5961 (N_5961,N_4566,N_4747);
and U5962 (N_5962,N_4582,N_4648);
or U5963 (N_5963,N_4510,N_5171);
xnor U5964 (N_5964,N_4840,N_5182);
nand U5965 (N_5965,N_5079,N_5099);
xor U5966 (N_5966,N_4688,N_4618);
nor U5967 (N_5967,N_4748,N_5067);
and U5968 (N_5968,N_4595,N_5227);
or U5969 (N_5969,N_4922,N_4556);
xor U5970 (N_5970,N_4845,N_5225);
nand U5971 (N_5971,N_5163,N_4524);
or U5972 (N_5972,N_4718,N_5122);
nor U5973 (N_5973,N_4841,N_4527);
and U5974 (N_5974,N_4628,N_4808);
nor U5975 (N_5975,N_5056,N_4789);
or U5976 (N_5976,N_4767,N_4749);
and U5977 (N_5977,N_4631,N_5196);
nand U5978 (N_5978,N_4881,N_4599);
or U5979 (N_5979,N_5160,N_5190);
nor U5980 (N_5980,N_4510,N_4893);
and U5981 (N_5981,N_4892,N_5166);
or U5982 (N_5982,N_4991,N_5024);
xnor U5983 (N_5983,N_5051,N_5010);
xnor U5984 (N_5984,N_5134,N_5058);
xor U5985 (N_5985,N_5168,N_5003);
xnor U5986 (N_5986,N_5175,N_4995);
or U5987 (N_5987,N_4527,N_4778);
and U5988 (N_5988,N_4622,N_4845);
or U5989 (N_5989,N_4758,N_4736);
nor U5990 (N_5990,N_4935,N_4997);
nor U5991 (N_5991,N_4681,N_4847);
and U5992 (N_5992,N_4965,N_4708);
nor U5993 (N_5993,N_4976,N_4585);
nand U5994 (N_5994,N_4690,N_4653);
xor U5995 (N_5995,N_5220,N_4854);
and U5996 (N_5996,N_4733,N_5084);
nor U5997 (N_5997,N_4893,N_4562);
xnor U5998 (N_5998,N_4920,N_4837);
xnor U5999 (N_5999,N_4914,N_4913);
xor U6000 (N_6000,N_5914,N_5567);
xor U6001 (N_6001,N_5357,N_5749);
or U6002 (N_6002,N_5921,N_5602);
nand U6003 (N_6003,N_5833,N_5638);
and U6004 (N_6004,N_5999,N_5812);
or U6005 (N_6005,N_5796,N_5472);
nor U6006 (N_6006,N_5960,N_5656);
nand U6007 (N_6007,N_5565,N_5969);
nand U6008 (N_6008,N_5977,N_5498);
and U6009 (N_6009,N_5381,N_5781);
xor U6010 (N_6010,N_5671,N_5732);
nor U6011 (N_6011,N_5628,N_5494);
or U6012 (N_6012,N_5410,N_5646);
or U6013 (N_6013,N_5500,N_5490);
nor U6014 (N_6014,N_5353,N_5540);
and U6015 (N_6015,N_5316,N_5582);
nor U6016 (N_6016,N_5735,N_5295);
nand U6017 (N_6017,N_5529,N_5454);
and U6018 (N_6018,N_5259,N_5407);
nand U6019 (N_6019,N_5280,N_5619);
nor U6020 (N_6020,N_5533,N_5400);
or U6021 (N_6021,N_5416,N_5726);
nor U6022 (N_6022,N_5463,N_5904);
xnor U6023 (N_6023,N_5830,N_5840);
nor U6024 (N_6024,N_5466,N_5285);
nor U6025 (N_6025,N_5720,N_5837);
or U6026 (N_6026,N_5544,N_5818);
nor U6027 (N_6027,N_5508,N_5542);
nand U6028 (N_6028,N_5651,N_5346);
or U6029 (N_6029,N_5419,N_5701);
or U6030 (N_6030,N_5725,N_5491);
or U6031 (N_6031,N_5906,N_5978);
xnor U6032 (N_6032,N_5807,N_5449);
nor U6033 (N_6033,N_5378,N_5415);
nor U6034 (N_6034,N_5344,N_5517);
xor U6035 (N_6035,N_5547,N_5771);
nor U6036 (N_6036,N_5355,N_5505);
nand U6037 (N_6037,N_5459,N_5342);
nand U6038 (N_6038,N_5982,N_5924);
nand U6039 (N_6039,N_5279,N_5974);
nand U6040 (N_6040,N_5988,N_5553);
and U6041 (N_6041,N_5629,N_5739);
xor U6042 (N_6042,N_5976,N_5816);
nand U6043 (N_6043,N_5603,N_5691);
or U6044 (N_6044,N_5343,N_5823);
xor U6045 (N_6045,N_5736,N_5380);
and U6046 (N_6046,N_5849,N_5668);
nand U6047 (N_6047,N_5723,N_5728);
nor U6048 (N_6048,N_5263,N_5789);
or U6049 (N_6049,N_5809,N_5584);
or U6050 (N_6050,N_5918,N_5697);
nand U6051 (N_6051,N_5273,N_5624);
xor U6052 (N_6052,N_5276,N_5888);
xnor U6053 (N_6053,N_5990,N_5942);
and U6054 (N_6054,N_5297,N_5984);
nor U6055 (N_6055,N_5401,N_5250);
xnor U6056 (N_6056,N_5580,N_5957);
or U6057 (N_6057,N_5635,N_5323);
and U6058 (N_6058,N_5927,N_5703);
nor U6059 (N_6059,N_5559,N_5757);
nand U6060 (N_6060,N_5575,N_5621);
xor U6061 (N_6061,N_5506,N_5896);
nor U6062 (N_6062,N_5855,N_5555);
or U6063 (N_6063,N_5499,N_5753);
nor U6064 (N_6064,N_5819,N_5956);
nand U6065 (N_6065,N_5875,N_5802);
or U6066 (N_6066,N_5300,N_5948);
or U6067 (N_6067,N_5398,N_5901);
nor U6068 (N_6068,N_5859,N_5457);
nor U6069 (N_6069,N_5886,N_5554);
or U6070 (N_6070,N_5793,N_5681);
and U6071 (N_6071,N_5714,N_5480);
and U6072 (N_6072,N_5980,N_5907);
xnor U6073 (N_6073,N_5366,N_5528);
xnor U6074 (N_6074,N_5922,N_5332);
and U6075 (N_6075,N_5813,N_5939);
nand U6076 (N_6076,N_5595,N_5665);
and U6077 (N_6077,N_5836,N_5876);
nand U6078 (N_6078,N_5287,N_5255);
or U6079 (N_6079,N_5623,N_5814);
nor U6080 (N_6080,N_5427,N_5985);
or U6081 (N_6081,N_5829,N_5429);
and U6082 (N_6082,N_5981,N_5851);
xor U6083 (N_6083,N_5549,N_5538);
nand U6084 (N_6084,N_5804,N_5663);
xnor U6085 (N_6085,N_5800,N_5871);
xnor U6086 (N_6086,N_5405,N_5271);
nor U6087 (N_6087,N_5435,N_5510);
or U6088 (N_6088,N_5509,N_5399);
or U6089 (N_6089,N_5596,N_5729);
or U6090 (N_6090,N_5717,N_5310);
nand U6091 (N_6091,N_5899,N_5666);
and U6092 (N_6092,N_5778,N_5917);
nor U6093 (N_6093,N_5493,N_5867);
or U6094 (N_6094,N_5556,N_5507);
xor U6095 (N_6095,N_5546,N_5471);
nand U6096 (N_6096,N_5261,N_5425);
nor U6097 (N_6097,N_5303,N_5698);
and U6098 (N_6098,N_5590,N_5811);
or U6099 (N_6099,N_5947,N_5946);
nor U6100 (N_6100,N_5335,N_5474);
or U6101 (N_6101,N_5721,N_5755);
xor U6102 (N_6102,N_5945,N_5423);
nand U6103 (N_6103,N_5368,N_5451);
nand U6104 (N_6104,N_5933,N_5305);
or U6105 (N_6105,N_5842,N_5880);
and U6106 (N_6106,N_5317,N_5857);
or U6107 (N_6107,N_5847,N_5543);
and U6108 (N_6108,N_5846,N_5356);
or U6109 (N_6109,N_5358,N_5684);
xor U6110 (N_6110,N_5839,N_5785);
nor U6111 (N_6111,N_5563,N_5722);
or U6112 (N_6112,N_5277,N_5518);
nand U6113 (N_6113,N_5444,N_5627);
or U6114 (N_6114,N_5388,N_5607);
xor U6115 (N_6115,N_5864,N_5395);
nand U6116 (N_6116,N_5309,N_5325);
nor U6117 (N_6117,N_5620,N_5754);
nand U6118 (N_6118,N_5994,N_5660);
nand U6119 (N_6119,N_5558,N_5975);
or U6120 (N_6120,N_5586,N_5339);
xnor U6121 (N_6121,N_5570,N_5869);
nand U6122 (N_6122,N_5955,N_5311);
nand U6123 (N_6123,N_5943,N_5485);
xnor U6124 (N_6124,N_5252,N_5387);
nor U6125 (N_6125,N_5411,N_5461);
nor U6126 (N_6126,N_5970,N_5272);
or U6127 (N_6127,N_5340,N_5386);
nor U6128 (N_6128,N_5827,N_5940);
or U6129 (N_6129,N_5908,N_5515);
xnor U6130 (N_6130,N_5696,N_5568);
nor U6131 (N_6131,N_5376,N_5751);
or U6132 (N_6132,N_5594,N_5597);
and U6133 (N_6133,N_5712,N_5455);
or U6134 (N_6134,N_5326,N_5963);
xor U6135 (N_6135,N_5430,N_5931);
or U6136 (N_6136,N_5662,N_5614);
xor U6137 (N_6137,N_5686,N_5706);
nand U6138 (N_6138,N_5936,N_5286);
nor U6139 (N_6139,N_5495,N_5450);
or U6140 (N_6140,N_5699,N_5532);
nor U6141 (N_6141,N_5889,N_5959);
xnor U6142 (N_6142,N_5448,N_5986);
and U6143 (N_6143,N_5612,N_5761);
xor U6144 (N_6144,N_5296,N_5693);
xor U6145 (N_6145,N_5862,N_5653);
xnor U6146 (N_6146,N_5473,N_5692);
or U6147 (N_6147,N_5962,N_5727);
nand U6148 (N_6148,N_5639,N_5593);
and U6149 (N_6149,N_5605,N_5803);
nor U6150 (N_6150,N_5884,N_5991);
nor U6151 (N_6151,N_5930,N_5831);
nor U6152 (N_6152,N_5441,N_5989);
xnor U6153 (N_6153,N_5501,N_5756);
and U6154 (N_6154,N_5371,N_5784);
nand U6155 (N_6155,N_5282,N_5935);
nand U6156 (N_6156,N_5731,N_5676);
or U6157 (N_6157,N_5810,N_5791);
xor U6158 (N_6158,N_5768,N_5661);
and U6159 (N_6159,N_5502,N_5903);
nand U6160 (N_6160,N_5369,N_5324);
xor U6161 (N_6161,N_5961,N_5445);
and U6162 (N_6162,N_5302,N_5608);
nor U6163 (N_6163,N_5929,N_5587);
nor U6164 (N_6164,N_5599,N_5633);
and U6165 (N_6165,N_5630,N_5290);
nor U6166 (N_6166,N_5695,N_5583);
or U6167 (N_6167,N_5737,N_5359);
nand U6168 (N_6168,N_5777,N_5534);
or U6169 (N_6169,N_5709,N_5477);
nand U6170 (N_6170,N_5571,N_5915);
or U6171 (N_6171,N_5611,N_5557);
and U6172 (N_6172,N_5648,N_5911);
xnor U6173 (N_6173,N_5622,N_5504);
or U6174 (N_6174,N_5598,N_5805);
or U6175 (N_6175,N_5394,N_5436);
nor U6176 (N_6176,N_5600,N_5458);
nand U6177 (N_6177,N_5774,N_5541);
nand U6178 (N_6178,N_5251,N_5408);
or U6179 (N_6179,N_5421,N_5431);
or U6180 (N_6180,N_5674,N_5307);
or U6181 (N_6181,N_5375,N_5437);
and U6182 (N_6182,N_5258,N_5841);
or U6183 (N_6183,N_5492,N_5481);
nand U6184 (N_6184,N_5535,N_5617);
and U6185 (N_6185,N_5820,N_5397);
and U6186 (N_6186,N_5779,N_5858);
xor U6187 (N_6187,N_5524,N_5987);
or U6188 (N_6188,N_5897,N_5744);
nand U6189 (N_6189,N_5298,N_5996);
nand U6190 (N_6190,N_5320,N_5578);
nand U6191 (N_6191,N_5522,N_5641);
nor U6192 (N_6192,N_5952,N_5657);
and U6193 (N_6193,N_5604,N_5377);
or U6194 (N_6194,N_5764,N_5844);
or U6195 (N_6195,N_5750,N_5256);
nand U6196 (N_6196,N_5592,N_5782);
nor U6197 (N_6197,N_5951,N_5446);
xnor U6198 (N_6198,N_5885,N_5306);
nand U6199 (N_6199,N_5792,N_5352);
nor U6200 (N_6200,N_5759,N_5579);
nand U6201 (N_6201,N_5349,N_5367);
or U6202 (N_6202,N_5995,N_5314);
or U6203 (N_6203,N_5746,N_5776);
nand U6204 (N_6204,N_5937,N_5870);
or U6205 (N_6205,N_5513,N_5610);
and U6206 (N_6206,N_5413,N_5724);
nor U6207 (N_6207,N_5853,N_5385);
nand U6208 (N_6208,N_5467,N_5716);
or U6209 (N_6209,N_5438,N_5488);
or U6210 (N_6210,N_5404,N_5525);
or U6211 (N_6211,N_5968,N_5364);
or U6212 (N_6212,N_5516,N_5333);
xor U6213 (N_6213,N_5420,N_5391);
nor U6214 (N_6214,N_5760,N_5403);
or U6215 (N_6215,N_5512,N_5257);
and U6216 (N_6216,N_5758,N_5912);
and U6217 (N_6217,N_5878,N_5389);
nand U6218 (N_6218,N_5925,N_5905);
nand U6219 (N_6219,N_5655,N_5672);
and U6220 (N_6220,N_5428,N_5414);
and U6221 (N_6221,N_5384,N_5944);
xnor U6222 (N_6222,N_5669,N_5322);
or U6223 (N_6223,N_5898,N_5609);
xor U6224 (N_6224,N_5890,N_5283);
and U6225 (N_6225,N_5848,N_5365);
xnor U6226 (N_6226,N_5521,N_5954);
nor U6227 (N_6227,N_5462,N_5312);
or U6228 (N_6228,N_5328,N_5762);
nand U6229 (N_6229,N_5275,N_5742);
nand U6230 (N_6230,N_5783,N_5442);
nand U6231 (N_6231,N_5845,N_5993);
nor U6232 (N_6232,N_5478,N_5456);
and U6233 (N_6233,N_5550,N_5329);
nor U6234 (N_6234,N_5647,N_5564);
nand U6235 (N_6235,N_5468,N_5688);
xor U6236 (N_6236,N_5308,N_5267);
nor U6237 (N_6237,N_5766,N_5797);
nand U6238 (N_6238,N_5643,N_5971);
and U6239 (N_6239,N_5799,N_5392);
nand U6240 (N_6240,N_5511,N_5664);
nor U6241 (N_6241,N_5426,N_5531);
nand U6242 (N_6242,N_5626,N_5319);
xnor U6243 (N_6243,N_5795,N_5520);
xor U6244 (N_6244,N_5920,N_5383);
and U6245 (N_6245,N_5879,N_5685);
nor U6246 (N_6246,N_5483,N_5958);
or U6247 (N_6247,N_5824,N_5825);
nand U6248 (N_6248,N_5689,N_5748);
nor U6249 (N_6249,N_5964,N_5850);
nand U6250 (N_6250,N_5747,N_5497);
xor U6251 (N_6251,N_5682,N_5552);
nor U6252 (N_6252,N_5266,N_5265);
nor U6253 (N_6253,N_5852,N_5569);
or U6254 (N_6254,N_5496,N_5432);
nor U6255 (N_6255,N_5424,N_5433);
or U6256 (N_6256,N_5828,N_5928);
xor U6257 (N_6257,N_5469,N_5337);
or U6258 (N_6258,N_5362,N_5363);
nor U6259 (N_6259,N_5268,N_5965);
xor U6260 (N_6260,N_5270,N_5560);
xnor U6261 (N_6261,N_5562,N_5973);
xor U6262 (N_6262,N_5484,N_5801);
xnor U6263 (N_6263,N_5293,N_5460);
and U6264 (N_6264,N_5406,N_5821);
and U6265 (N_6265,N_5330,N_5770);
nand U6266 (N_6266,N_5327,N_5345);
and U6267 (N_6267,N_5637,N_5966);
nor U6268 (N_6268,N_5677,N_5338);
xor U6269 (N_6269,N_5412,N_5798);
nor U6270 (N_6270,N_5861,N_5618);
or U6271 (N_6271,N_5577,N_5763);
nor U6272 (N_6272,N_5659,N_5418);
or U6273 (N_6273,N_5895,N_5486);
xor U6274 (N_6274,N_5949,N_5872);
xnor U6275 (N_6275,N_5923,N_5834);
xor U6276 (N_6276,N_5794,N_5601);
or U6277 (N_6277,N_5576,N_5396);
and U6278 (N_6278,N_5390,N_5336);
nor U6279 (N_6279,N_5658,N_5892);
xnor U6280 (N_6280,N_5941,N_5274);
nand U6281 (N_6281,N_5281,N_5765);
and U6282 (N_6282,N_5854,N_5767);
nor U6283 (N_6283,N_5983,N_5606);
xnor U6284 (N_6284,N_5713,N_5860);
nor U6285 (N_6285,N_5642,N_5482);
nor U6286 (N_6286,N_5883,N_5979);
or U6287 (N_6287,N_5919,N_5434);
nand U6288 (N_6288,N_5301,N_5572);
nor U6289 (N_6289,N_5680,N_5289);
and U6290 (N_6290,N_5704,N_5304);
nand U6291 (N_6291,N_5745,N_5780);
and U6292 (N_6292,N_5718,N_5932);
nand U6293 (N_6293,N_5514,N_5909);
and U6294 (N_6294,N_5351,N_5788);
nor U6295 (N_6295,N_5675,N_5856);
nand U6296 (N_6296,N_5588,N_5667);
nor U6297 (N_6297,N_5752,N_5687);
nand U6298 (N_6298,N_5715,N_5616);
or U6299 (N_6299,N_5530,N_5551);
nand U6300 (N_6300,N_5694,N_5331);
nand U6301 (N_6301,N_5710,N_5683);
or U6302 (N_6302,N_5719,N_5992);
and U6303 (N_6303,N_5998,N_5519);
and U6304 (N_6304,N_5278,N_5341);
or U6305 (N_6305,N_5806,N_5645);
nand U6306 (N_6306,N_5422,N_5370);
nand U6307 (N_6307,N_5741,N_5372);
and U6308 (N_6308,N_5615,N_5972);
and U6309 (N_6309,N_5773,N_5262);
nor U6310 (N_6310,N_5347,N_5253);
xnor U6311 (N_6311,N_5393,N_5877);
nor U6312 (N_6312,N_5934,N_5561);
xor U6313 (N_6313,N_5900,N_5650);
nor U6314 (N_6314,N_5409,N_5536);
and U6315 (N_6315,N_5874,N_5470);
nand U6316 (N_6316,N_5269,N_5866);
nor U6317 (N_6317,N_5926,N_5613);
or U6318 (N_6318,N_5835,N_5464);
or U6319 (N_6319,N_5882,N_5772);
xor U6320 (N_6320,N_5284,N_5887);
nor U6321 (N_6321,N_5868,N_5953);
nand U6322 (N_6322,N_5902,N_5631);
xor U6323 (N_6323,N_5581,N_5702);
nor U6324 (N_6324,N_5260,N_5670);
nand U6325 (N_6325,N_5916,N_5863);
or U6326 (N_6326,N_5738,N_5808);
nand U6327 (N_6327,N_5527,N_5440);
or U6328 (N_6328,N_5787,N_5997);
xnor U6329 (N_6329,N_5374,N_5734);
nor U6330 (N_6330,N_5475,N_5707);
nand U6331 (N_6331,N_5967,N_5443);
and U6332 (N_6332,N_5822,N_5361);
and U6333 (N_6333,N_5817,N_5313);
and U6334 (N_6334,N_5894,N_5865);
and U6335 (N_6335,N_5354,N_5315);
or U6336 (N_6336,N_5299,N_5453);
nand U6337 (N_6337,N_5775,N_5740);
nand U6338 (N_6338,N_5649,N_5573);
nor U6339 (N_6339,N_5690,N_5881);
nand U6340 (N_6340,N_5733,N_5891);
nor U6341 (N_6341,N_5264,N_5708);
or U6342 (N_6342,N_5288,N_5838);
nand U6343 (N_6343,N_5938,N_5815);
nand U6344 (N_6344,N_5523,N_5910);
xor U6345 (N_6345,N_5644,N_5730);
or U6346 (N_6346,N_5526,N_5585);
and U6347 (N_6347,N_5636,N_5539);
nand U6348 (N_6348,N_5350,N_5487);
or U6349 (N_6349,N_5634,N_5673);
and U6350 (N_6350,N_5379,N_5640);
or U6351 (N_6351,N_5348,N_5632);
and U6352 (N_6352,N_5382,N_5743);
and U6353 (N_6353,N_5893,N_5503);
or U6354 (N_6354,N_5465,N_5545);
and U6355 (N_6355,N_5913,N_5360);
nor U6356 (N_6356,N_5318,N_5294);
xnor U6357 (N_6357,N_5950,N_5334);
and U6358 (N_6358,N_5548,N_5566);
nand U6359 (N_6359,N_5705,N_5843);
or U6360 (N_6360,N_5291,N_5652);
nand U6361 (N_6361,N_5479,N_5678);
or U6362 (N_6362,N_5476,N_5711);
xor U6363 (N_6363,N_5790,N_5786);
and U6364 (N_6364,N_5254,N_5402);
and U6365 (N_6365,N_5489,N_5873);
or U6366 (N_6366,N_5625,N_5589);
xnor U6367 (N_6367,N_5452,N_5679);
nand U6368 (N_6368,N_5832,N_5769);
xor U6369 (N_6369,N_5321,N_5447);
xnor U6370 (N_6370,N_5654,N_5292);
nor U6371 (N_6371,N_5826,N_5373);
or U6372 (N_6372,N_5537,N_5700);
xor U6373 (N_6373,N_5417,N_5574);
and U6374 (N_6374,N_5439,N_5591);
nor U6375 (N_6375,N_5529,N_5505);
nand U6376 (N_6376,N_5384,N_5443);
nand U6377 (N_6377,N_5673,N_5250);
or U6378 (N_6378,N_5449,N_5949);
nand U6379 (N_6379,N_5813,N_5560);
and U6380 (N_6380,N_5331,N_5314);
nor U6381 (N_6381,N_5829,N_5477);
and U6382 (N_6382,N_5855,N_5289);
or U6383 (N_6383,N_5333,N_5501);
xor U6384 (N_6384,N_5798,N_5771);
nor U6385 (N_6385,N_5929,N_5540);
nor U6386 (N_6386,N_5320,N_5331);
xor U6387 (N_6387,N_5255,N_5752);
xnor U6388 (N_6388,N_5959,N_5679);
or U6389 (N_6389,N_5363,N_5971);
and U6390 (N_6390,N_5722,N_5895);
or U6391 (N_6391,N_5763,N_5776);
xor U6392 (N_6392,N_5535,N_5689);
xnor U6393 (N_6393,N_5270,N_5294);
nand U6394 (N_6394,N_5644,N_5451);
and U6395 (N_6395,N_5954,N_5767);
xor U6396 (N_6396,N_5936,N_5642);
nand U6397 (N_6397,N_5622,N_5873);
or U6398 (N_6398,N_5963,N_5589);
or U6399 (N_6399,N_5393,N_5542);
nand U6400 (N_6400,N_5760,N_5461);
nand U6401 (N_6401,N_5679,N_5308);
xnor U6402 (N_6402,N_5517,N_5827);
xnor U6403 (N_6403,N_5557,N_5368);
and U6404 (N_6404,N_5450,N_5404);
nor U6405 (N_6405,N_5267,N_5469);
and U6406 (N_6406,N_5950,N_5464);
or U6407 (N_6407,N_5989,N_5827);
and U6408 (N_6408,N_5712,N_5846);
nand U6409 (N_6409,N_5644,N_5826);
nand U6410 (N_6410,N_5382,N_5496);
nor U6411 (N_6411,N_5963,N_5779);
nand U6412 (N_6412,N_5483,N_5469);
or U6413 (N_6413,N_5674,N_5282);
nand U6414 (N_6414,N_5439,N_5377);
or U6415 (N_6415,N_5960,N_5309);
xnor U6416 (N_6416,N_5397,N_5620);
xor U6417 (N_6417,N_5594,N_5605);
or U6418 (N_6418,N_5463,N_5811);
nand U6419 (N_6419,N_5668,N_5295);
and U6420 (N_6420,N_5831,N_5354);
and U6421 (N_6421,N_5595,N_5847);
or U6422 (N_6422,N_5648,N_5337);
nand U6423 (N_6423,N_5601,N_5427);
or U6424 (N_6424,N_5565,N_5639);
nand U6425 (N_6425,N_5481,N_5435);
nand U6426 (N_6426,N_5926,N_5780);
nor U6427 (N_6427,N_5830,N_5833);
or U6428 (N_6428,N_5502,N_5425);
or U6429 (N_6429,N_5706,N_5592);
xor U6430 (N_6430,N_5982,N_5349);
nor U6431 (N_6431,N_5260,N_5273);
nor U6432 (N_6432,N_5394,N_5608);
nand U6433 (N_6433,N_5372,N_5501);
xor U6434 (N_6434,N_5620,N_5322);
and U6435 (N_6435,N_5961,N_5513);
and U6436 (N_6436,N_5351,N_5416);
or U6437 (N_6437,N_5378,N_5448);
nand U6438 (N_6438,N_5453,N_5870);
or U6439 (N_6439,N_5267,N_5454);
xor U6440 (N_6440,N_5381,N_5941);
nor U6441 (N_6441,N_5581,N_5763);
and U6442 (N_6442,N_5704,N_5777);
nand U6443 (N_6443,N_5561,N_5794);
nand U6444 (N_6444,N_5260,N_5804);
nor U6445 (N_6445,N_5799,N_5849);
or U6446 (N_6446,N_5540,N_5446);
or U6447 (N_6447,N_5601,N_5436);
and U6448 (N_6448,N_5450,N_5862);
xnor U6449 (N_6449,N_5301,N_5531);
or U6450 (N_6450,N_5946,N_5443);
xor U6451 (N_6451,N_5874,N_5862);
nand U6452 (N_6452,N_5452,N_5911);
or U6453 (N_6453,N_5312,N_5482);
or U6454 (N_6454,N_5289,N_5904);
nand U6455 (N_6455,N_5720,N_5262);
or U6456 (N_6456,N_5426,N_5623);
and U6457 (N_6457,N_5774,N_5625);
and U6458 (N_6458,N_5266,N_5403);
xor U6459 (N_6459,N_5314,N_5383);
nand U6460 (N_6460,N_5423,N_5415);
or U6461 (N_6461,N_5836,N_5565);
xor U6462 (N_6462,N_5342,N_5554);
and U6463 (N_6463,N_5829,N_5288);
and U6464 (N_6464,N_5379,N_5606);
and U6465 (N_6465,N_5934,N_5659);
xnor U6466 (N_6466,N_5966,N_5539);
or U6467 (N_6467,N_5856,N_5427);
xnor U6468 (N_6468,N_5403,N_5525);
nand U6469 (N_6469,N_5539,N_5900);
and U6470 (N_6470,N_5687,N_5859);
nand U6471 (N_6471,N_5806,N_5651);
nand U6472 (N_6472,N_5635,N_5584);
xnor U6473 (N_6473,N_5637,N_5898);
xor U6474 (N_6474,N_5277,N_5363);
or U6475 (N_6475,N_5441,N_5464);
or U6476 (N_6476,N_5376,N_5424);
nor U6477 (N_6477,N_5291,N_5898);
nor U6478 (N_6478,N_5620,N_5316);
nand U6479 (N_6479,N_5506,N_5959);
xor U6480 (N_6480,N_5313,N_5541);
nor U6481 (N_6481,N_5999,N_5693);
nor U6482 (N_6482,N_5726,N_5326);
nand U6483 (N_6483,N_5460,N_5994);
xor U6484 (N_6484,N_5293,N_5772);
or U6485 (N_6485,N_5628,N_5811);
and U6486 (N_6486,N_5915,N_5481);
xor U6487 (N_6487,N_5317,N_5800);
nand U6488 (N_6488,N_5542,N_5484);
nor U6489 (N_6489,N_5476,N_5713);
or U6490 (N_6490,N_5540,N_5271);
or U6491 (N_6491,N_5440,N_5964);
and U6492 (N_6492,N_5698,N_5361);
or U6493 (N_6493,N_5407,N_5649);
and U6494 (N_6494,N_5288,N_5257);
nand U6495 (N_6495,N_5617,N_5321);
xnor U6496 (N_6496,N_5613,N_5533);
nand U6497 (N_6497,N_5459,N_5284);
nand U6498 (N_6498,N_5517,N_5551);
nand U6499 (N_6499,N_5398,N_5316);
nor U6500 (N_6500,N_5940,N_5624);
or U6501 (N_6501,N_5816,N_5809);
or U6502 (N_6502,N_5405,N_5946);
xor U6503 (N_6503,N_5607,N_5356);
nor U6504 (N_6504,N_5747,N_5414);
nor U6505 (N_6505,N_5716,N_5664);
and U6506 (N_6506,N_5589,N_5363);
and U6507 (N_6507,N_5866,N_5828);
and U6508 (N_6508,N_5396,N_5440);
xor U6509 (N_6509,N_5285,N_5267);
nand U6510 (N_6510,N_5991,N_5547);
or U6511 (N_6511,N_5542,N_5336);
nor U6512 (N_6512,N_5468,N_5386);
or U6513 (N_6513,N_5933,N_5755);
nor U6514 (N_6514,N_5799,N_5655);
or U6515 (N_6515,N_5746,N_5875);
or U6516 (N_6516,N_5994,N_5999);
nor U6517 (N_6517,N_5316,N_5958);
nand U6518 (N_6518,N_5251,N_5799);
xor U6519 (N_6519,N_5579,N_5696);
nor U6520 (N_6520,N_5326,N_5487);
and U6521 (N_6521,N_5382,N_5337);
nand U6522 (N_6522,N_5379,N_5436);
nor U6523 (N_6523,N_5605,N_5978);
and U6524 (N_6524,N_5671,N_5696);
or U6525 (N_6525,N_5618,N_5834);
xor U6526 (N_6526,N_5563,N_5317);
or U6527 (N_6527,N_5872,N_5427);
nor U6528 (N_6528,N_5964,N_5255);
xor U6529 (N_6529,N_5285,N_5740);
xnor U6530 (N_6530,N_5944,N_5267);
and U6531 (N_6531,N_5782,N_5626);
xnor U6532 (N_6532,N_5790,N_5920);
xor U6533 (N_6533,N_5533,N_5508);
and U6534 (N_6534,N_5692,N_5961);
or U6535 (N_6535,N_5550,N_5782);
nor U6536 (N_6536,N_5416,N_5709);
and U6537 (N_6537,N_5772,N_5542);
and U6538 (N_6538,N_5404,N_5393);
nor U6539 (N_6539,N_5307,N_5303);
and U6540 (N_6540,N_5537,N_5324);
nor U6541 (N_6541,N_5266,N_5510);
and U6542 (N_6542,N_5880,N_5475);
nor U6543 (N_6543,N_5694,N_5749);
xnor U6544 (N_6544,N_5856,N_5546);
nor U6545 (N_6545,N_5535,N_5954);
nor U6546 (N_6546,N_5542,N_5358);
or U6547 (N_6547,N_5285,N_5603);
nand U6548 (N_6548,N_5428,N_5965);
nand U6549 (N_6549,N_5864,N_5737);
nand U6550 (N_6550,N_5319,N_5992);
or U6551 (N_6551,N_5287,N_5312);
and U6552 (N_6552,N_5952,N_5345);
nand U6553 (N_6553,N_5681,N_5718);
nand U6554 (N_6554,N_5253,N_5914);
and U6555 (N_6555,N_5404,N_5989);
or U6556 (N_6556,N_5856,N_5867);
or U6557 (N_6557,N_5619,N_5792);
xor U6558 (N_6558,N_5363,N_5901);
nor U6559 (N_6559,N_5255,N_5376);
nor U6560 (N_6560,N_5450,N_5967);
nand U6561 (N_6561,N_5439,N_5782);
xor U6562 (N_6562,N_5687,N_5264);
nor U6563 (N_6563,N_5620,N_5698);
and U6564 (N_6564,N_5975,N_5658);
nand U6565 (N_6565,N_5382,N_5289);
xnor U6566 (N_6566,N_5356,N_5719);
and U6567 (N_6567,N_5714,N_5934);
and U6568 (N_6568,N_5666,N_5517);
nor U6569 (N_6569,N_5852,N_5696);
nand U6570 (N_6570,N_5425,N_5290);
or U6571 (N_6571,N_5438,N_5695);
nor U6572 (N_6572,N_5964,N_5896);
and U6573 (N_6573,N_5416,N_5623);
nand U6574 (N_6574,N_5682,N_5257);
and U6575 (N_6575,N_5467,N_5395);
xor U6576 (N_6576,N_5852,N_5534);
xnor U6577 (N_6577,N_5944,N_5428);
or U6578 (N_6578,N_5683,N_5300);
and U6579 (N_6579,N_5258,N_5752);
nand U6580 (N_6580,N_5996,N_5290);
xnor U6581 (N_6581,N_5936,N_5273);
and U6582 (N_6582,N_5986,N_5322);
nor U6583 (N_6583,N_5452,N_5529);
nand U6584 (N_6584,N_5414,N_5896);
and U6585 (N_6585,N_5804,N_5456);
nor U6586 (N_6586,N_5278,N_5257);
or U6587 (N_6587,N_5925,N_5487);
and U6588 (N_6588,N_5894,N_5918);
and U6589 (N_6589,N_5688,N_5264);
nand U6590 (N_6590,N_5826,N_5708);
xor U6591 (N_6591,N_5395,N_5260);
or U6592 (N_6592,N_5686,N_5371);
nor U6593 (N_6593,N_5769,N_5678);
nor U6594 (N_6594,N_5782,N_5768);
nor U6595 (N_6595,N_5265,N_5366);
nand U6596 (N_6596,N_5819,N_5301);
xor U6597 (N_6597,N_5846,N_5479);
nand U6598 (N_6598,N_5629,N_5995);
or U6599 (N_6599,N_5265,N_5705);
nor U6600 (N_6600,N_5806,N_5604);
and U6601 (N_6601,N_5973,N_5470);
and U6602 (N_6602,N_5718,N_5575);
xor U6603 (N_6603,N_5709,N_5598);
and U6604 (N_6604,N_5347,N_5474);
xor U6605 (N_6605,N_5442,N_5775);
nand U6606 (N_6606,N_5271,N_5823);
nor U6607 (N_6607,N_5250,N_5626);
nand U6608 (N_6608,N_5843,N_5453);
nor U6609 (N_6609,N_5491,N_5647);
nand U6610 (N_6610,N_5960,N_5852);
or U6611 (N_6611,N_5380,N_5539);
xor U6612 (N_6612,N_5676,N_5719);
or U6613 (N_6613,N_5382,N_5523);
or U6614 (N_6614,N_5931,N_5593);
nand U6615 (N_6615,N_5826,N_5565);
or U6616 (N_6616,N_5730,N_5392);
and U6617 (N_6617,N_5597,N_5679);
nor U6618 (N_6618,N_5659,N_5354);
nor U6619 (N_6619,N_5610,N_5884);
nand U6620 (N_6620,N_5291,N_5856);
nor U6621 (N_6621,N_5743,N_5799);
nand U6622 (N_6622,N_5660,N_5790);
xnor U6623 (N_6623,N_5630,N_5367);
or U6624 (N_6624,N_5916,N_5290);
or U6625 (N_6625,N_5936,N_5321);
and U6626 (N_6626,N_5902,N_5479);
nand U6627 (N_6627,N_5420,N_5399);
or U6628 (N_6628,N_5617,N_5925);
xor U6629 (N_6629,N_5966,N_5750);
xnor U6630 (N_6630,N_5428,N_5455);
nor U6631 (N_6631,N_5334,N_5710);
xor U6632 (N_6632,N_5959,N_5511);
nor U6633 (N_6633,N_5719,N_5839);
nor U6634 (N_6634,N_5924,N_5701);
and U6635 (N_6635,N_5668,N_5277);
nor U6636 (N_6636,N_5821,N_5931);
nor U6637 (N_6637,N_5922,N_5471);
nor U6638 (N_6638,N_5339,N_5927);
and U6639 (N_6639,N_5267,N_5754);
and U6640 (N_6640,N_5675,N_5858);
nand U6641 (N_6641,N_5835,N_5845);
xnor U6642 (N_6642,N_5306,N_5901);
nand U6643 (N_6643,N_5256,N_5396);
or U6644 (N_6644,N_5899,N_5645);
and U6645 (N_6645,N_5598,N_5795);
and U6646 (N_6646,N_5477,N_5828);
nand U6647 (N_6647,N_5530,N_5818);
and U6648 (N_6648,N_5799,N_5628);
or U6649 (N_6649,N_5937,N_5747);
nand U6650 (N_6650,N_5635,N_5756);
and U6651 (N_6651,N_5756,N_5344);
nor U6652 (N_6652,N_5977,N_5968);
nor U6653 (N_6653,N_5604,N_5968);
nand U6654 (N_6654,N_5430,N_5580);
nor U6655 (N_6655,N_5978,N_5299);
and U6656 (N_6656,N_5526,N_5514);
xnor U6657 (N_6657,N_5354,N_5258);
or U6658 (N_6658,N_5597,N_5644);
and U6659 (N_6659,N_5925,N_5401);
or U6660 (N_6660,N_5845,N_5334);
xor U6661 (N_6661,N_5856,N_5432);
and U6662 (N_6662,N_5756,N_5594);
and U6663 (N_6663,N_5366,N_5404);
and U6664 (N_6664,N_5811,N_5352);
and U6665 (N_6665,N_5787,N_5262);
and U6666 (N_6666,N_5399,N_5854);
nor U6667 (N_6667,N_5402,N_5424);
or U6668 (N_6668,N_5808,N_5783);
nand U6669 (N_6669,N_5895,N_5829);
and U6670 (N_6670,N_5617,N_5361);
xnor U6671 (N_6671,N_5252,N_5967);
nand U6672 (N_6672,N_5739,N_5703);
nor U6673 (N_6673,N_5887,N_5704);
or U6674 (N_6674,N_5920,N_5323);
xor U6675 (N_6675,N_5578,N_5860);
and U6676 (N_6676,N_5989,N_5461);
or U6677 (N_6677,N_5827,N_5825);
nor U6678 (N_6678,N_5795,N_5596);
nor U6679 (N_6679,N_5586,N_5936);
or U6680 (N_6680,N_5810,N_5831);
nor U6681 (N_6681,N_5592,N_5805);
nor U6682 (N_6682,N_5340,N_5758);
nand U6683 (N_6683,N_5713,N_5750);
xnor U6684 (N_6684,N_5943,N_5428);
or U6685 (N_6685,N_5325,N_5320);
or U6686 (N_6686,N_5482,N_5938);
or U6687 (N_6687,N_5658,N_5458);
nand U6688 (N_6688,N_5514,N_5749);
xnor U6689 (N_6689,N_5366,N_5401);
or U6690 (N_6690,N_5359,N_5944);
xor U6691 (N_6691,N_5394,N_5775);
xnor U6692 (N_6692,N_5300,N_5609);
and U6693 (N_6693,N_5332,N_5471);
or U6694 (N_6694,N_5526,N_5759);
xnor U6695 (N_6695,N_5800,N_5719);
or U6696 (N_6696,N_5946,N_5762);
and U6697 (N_6697,N_5679,N_5351);
nor U6698 (N_6698,N_5847,N_5589);
nand U6699 (N_6699,N_5452,N_5543);
xnor U6700 (N_6700,N_5931,N_5505);
nor U6701 (N_6701,N_5838,N_5397);
and U6702 (N_6702,N_5789,N_5806);
xor U6703 (N_6703,N_5337,N_5455);
xnor U6704 (N_6704,N_5659,N_5780);
nand U6705 (N_6705,N_5902,N_5577);
and U6706 (N_6706,N_5507,N_5397);
xnor U6707 (N_6707,N_5252,N_5853);
and U6708 (N_6708,N_5402,N_5706);
or U6709 (N_6709,N_5264,N_5343);
nor U6710 (N_6710,N_5985,N_5570);
nand U6711 (N_6711,N_5401,N_5785);
nand U6712 (N_6712,N_5345,N_5548);
or U6713 (N_6713,N_5736,N_5258);
xnor U6714 (N_6714,N_5944,N_5704);
xor U6715 (N_6715,N_5409,N_5814);
nor U6716 (N_6716,N_5761,N_5883);
nor U6717 (N_6717,N_5443,N_5670);
and U6718 (N_6718,N_5669,N_5420);
and U6719 (N_6719,N_5624,N_5352);
nand U6720 (N_6720,N_5995,N_5904);
nand U6721 (N_6721,N_5823,N_5874);
and U6722 (N_6722,N_5589,N_5831);
xnor U6723 (N_6723,N_5430,N_5776);
and U6724 (N_6724,N_5516,N_5265);
nor U6725 (N_6725,N_5741,N_5302);
or U6726 (N_6726,N_5959,N_5382);
nand U6727 (N_6727,N_5986,N_5696);
xor U6728 (N_6728,N_5518,N_5336);
nor U6729 (N_6729,N_5275,N_5527);
nand U6730 (N_6730,N_5483,N_5837);
nor U6731 (N_6731,N_5363,N_5291);
or U6732 (N_6732,N_5780,N_5955);
nand U6733 (N_6733,N_5350,N_5847);
xor U6734 (N_6734,N_5530,N_5278);
and U6735 (N_6735,N_5876,N_5529);
nor U6736 (N_6736,N_5262,N_5571);
or U6737 (N_6737,N_5266,N_5840);
nand U6738 (N_6738,N_5529,N_5335);
or U6739 (N_6739,N_5454,N_5906);
or U6740 (N_6740,N_5267,N_5556);
and U6741 (N_6741,N_5584,N_5877);
and U6742 (N_6742,N_5727,N_5831);
nand U6743 (N_6743,N_5764,N_5757);
nor U6744 (N_6744,N_5457,N_5419);
or U6745 (N_6745,N_5661,N_5470);
nor U6746 (N_6746,N_5709,N_5261);
or U6747 (N_6747,N_5856,N_5839);
and U6748 (N_6748,N_5375,N_5494);
nand U6749 (N_6749,N_5394,N_5849);
or U6750 (N_6750,N_6419,N_6118);
xor U6751 (N_6751,N_6328,N_6332);
xor U6752 (N_6752,N_6434,N_6081);
xnor U6753 (N_6753,N_6686,N_6177);
or U6754 (N_6754,N_6107,N_6567);
nand U6755 (N_6755,N_6404,N_6164);
xnor U6756 (N_6756,N_6439,N_6651);
nand U6757 (N_6757,N_6741,N_6226);
xnor U6758 (N_6758,N_6090,N_6306);
and U6759 (N_6759,N_6634,N_6004);
nand U6760 (N_6760,N_6505,N_6155);
nand U6761 (N_6761,N_6274,N_6114);
or U6762 (N_6762,N_6513,N_6256);
or U6763 (N_6763,N_6504,N_6447);
and U6764 (N_6764,N_6574,N_6391);
xnor U6765 (N_6765,N_6215,N_6649);
nor U6766 (N_6766,N_6141,N_6636);
nor U6767 (N_6767,N_6465,N_6063);
and U6768 (N_6768,N_6161,N_6748);
and U6769 (N_6769,N_6749,N_6554);
xor U6770 (N_6770,N_6279,N_6502);
xor U6771 (N_6771,N_6607,N_6553);
xor U6772 (N_6772,N_6194,N_6217);
xor U6773 (N_6773,N_6363,N_6096);
or U6774 (N_6774,N_6029,N_6005);
nand U6775 (N_6775,N_6045,N_6015);
and U6776 (N_6776,N_6721,N_6514);
and U6777 (N_6777,N_6714,N_6443);
and U6778 (N_6778,N_6621,N_6684);
nor U6779 (N_6779,N_6136,N_6583);
and U6780 (N_6780,N_6251,N_6094);
xor U6781 (N_6781,N_6303,N_6196);
xor U6782 (N_6782,N_6182,N_6287);
nor U6783 (N_6783,N_6253,N_6658);
or U6784 (N_6784,N_6258,N_6396);
nor U6785 (N_6785,N_6405,N_6695);
nor U6786 (N_6786,N_6219,N_6578);
xor U6787 (N_6787,N_6490,N_6524);
nor U6788 (N_6788,N_6425,N_6101);
xor U6789 (N_6789,N_6086,N_6656);
xor U6790 (N_6790,N_6003,N_6377);
nor U6791 (N_6791,N_6066,N_6216);
nor U6792 (N_6792,N_6507,N_6739);
xor U6793 (N_6793,N_6384,N_6555);
nor U6794 (N_6794,N_6406,N_6175);
and U6795 (N_6795,N_6519,N_6603);
or U6796 (N_6796,N_6282,N_6509);
nor U6797 (N_6797,N_6059,N_6228);
nand U6798 (N_6798,N_6454,N_6461);
nor U6799 (N_6799,N_6460,N_6452);
and U6800 (N_6800,N_6517,N_6707);
xor U6801 (N_6801,N_6338,N_6103);
nor U6802 (N_6802,N_6489,N_6401);
nand U6803 (N_6803,N_6740,N_6624);
nor U6804 (N_6804,N_6685,N_6629);
nand U6805 (N_6805,N_6157,N_6133);
xnor U6806 (N_6806,N_6247,N_6618);
xnor U6807 (N_6807,N_6212,N_6218);
and U6808 (N_6808,N_6412,N_6350);
nor U6809 (N_6809,N_6298,N_6520);
nand U6810 (N_6810,N_6723,N_6604);
or U6811 (N_6811,N_6704,N_6158);
nand U6812 (N_6812,N_6682,N_6010);
or U6813 (N_6813,N_6331,N_6088);
and U6814 (N_6814,N_6676,N_6522);
nor U6815 (N_6815,N_6137,N_6605);
nor U6816 (N_6816,N_6060,N_6263);
xor U6817 (N_6817,N_6462,N_6450);
nand U6818 (N_6818,N_6055,N_6568);
nor U6819 (N_6819,N_6189,N_6213);
and U6820 (N_6820,N_6195,N_6523);
and U6821 (N_6821,N_6357,N_6261);
nor U6822 (N_6822,N_6458,N_6291);
and U6823 (N_6823,N_6360,N_6020);
nor U6824 (N_6824,N_6224,N_6613);
or U6825 (N_6825,N_6599,N_6722);
and U6826 (N_6826,N_6397,N_6386);
or U6827 (N_6827,N_6433,N_6210);
nor U6828 (N_6828,N_6645,N_6209);
or U6829 (N_6829,N_6423,N_6389);
nor U6830 (N_6830,N_6596,N_6488);
nor U6831 (N_6831,N_6250,N_6672);
or U6832 (N_6832,N_6470,N_6036);
nor U6833 (N_6833,N_6097,N_6302);
nand U6834 (N_6834,N_6173,N_6466);
nand U6835 (N_6835,N_6569,N_6487);
nand U6836 (N_6836,N_6072,N_6301);
or U6837 (N_6837,N_6065,N_6403);
nor U6838 (N_6838,N_6670,N_6491);
xnor U6839 (N_6839,N_6694,N_6731);
and U6840 (N_6840,N_6556,N_6659);
and U6841 (N_6841,N_6534,N_6483);
nor U6842 (N_6842,N_6371,N_6028);
nor U6843 (N_6843,N_6409,N_6482);
or U6844 (N_6844,N_6640,N_6130);
nand U6845 (N_6845,N_6273,N_6703);
nand U6846 (N_6846,N_6231,N_6283);
or U6847 (N_6847,N_6050,N_6011);
nor U6848 (N_6848,N_6495,N_6364);
and U6849 (N_6849,N_6293,N_6529);
and U6850 (N_6850,N_6733,N_6078);
nor U6851 (N_6851,N_6597,N_6627);
nor U6852 (N_6852,N_6361,N_6587);
xnor U6853 (N_6853,N_6288,N_6187);
nand U6854 (N_6854,N_6588,N_6132);
or U6855 (N_6855,N_6162,N_6134);
or U6856 (N_6856,N_6095,N_6615);
nor U6857 (N_6857,N_6149,N_6208);
and U6858 (N_6858,N_6308,N_6211);
nor U6859 (N_6859,N_6260,N_6563);
and U6860 (N_6860,N_6420,N_6252);
or U6861 (N_6861,N_6411,N_6329);
nand U6862 (N_6862,N_6738,N_6438);
nor U6863 (N_6863,N_6558,N_6675);
and U6864 (N_6864,N_6057,N_6085);
or U6865 (N_6865,N_6160,N_6430);
nand U6866 (N_6866,N_6052,N_6435);
xnor U6867 (N_6867,N_6700,N_6170);
or U6868 (N_6868,N_6117,N_6294);
xor U6869 (N_6869,N_6580,N_6742);
xnor U6870 (N_6870,N_6521,N_6018);
nor U6871 (N_6871,N_6617,N_6321);
xor U6872 (N_6872,N_6665,N_6269);
or U6873 (N_6873,N_6343,N_6115);
and U6874 (N_6874,N_6146,N_6471);
or U6875 (N_6875,N_6091,N_6056);
or U6876 (N_6876,N_6300,N_6584);
xnor U6877 (N_6877,N_6608,N_6598);
nor U6878 (N_6878,N_6637,N_6051);
or U6879 (N_6879,N_6375,N_6385);
or U6880 (N_6880,N_6436,N_6027);
and U6881 (N_6881,N_6666,N_6100);
or U6882 (N_6882,N_6729,N_6606);
nor U6883 (N_6883,N_6381,N_6105);
and U6884 (N_6884,N_6227,N_6625);
or U6885 (N_6885,N_6345,N_6198);
or U6886 (N_6886,N_6657,N_6688);
nand U6887 (N_6887,N_6418,N_6113);
or U6888 (N_6888,N_6082,N_6647);
xnor U6889 (N_6889,N_6501,N_6075);
nor U6890 (N_6890,N_6664,N_6248);
nor U6891 (N_6891,N_6234,N_6271);
nor U6892 (N_6892,N_6153,N_6706);
nor U6893 (N_6893,N_6653,N_6545);
nor U6894 (N_6894,N_6408,N_6573);
or U6895 (N_6895,N_6201,N_6203);
nor U6896 (N_6896,N_6498,N_6687);
or U6897 (N_6897,N_6549,N_6354);
xnor U6898 (N_6898,N_6204,N_6089);
or U6899 (N_6899,N_6214,N_6362);
and U6900 (N_6900,N_6309,N_6619);
xnor U6901 (N_6901,N_6631,N_6349);
and U6902 (N_6902,N_6046,N_6414);
xor U6903 (N_6903,N_6728,N_6266);
and U6904 (N_6904,N_6286,N_6221);
and U6905 (N_6905,N_6424,N_6372);
nor U6906 (N_6906,N_6323,N_6339);
nor U6907 (N_6907,N_6064,N_6415);
xor U6908 (N_6908,N_6727,N_6123);
xnor U6909 (N_6909,N_6241,N_6152);
xor U6910 (N_6910,N_6746,N_6382);
nand U6911 (N_6911,N_6453,N_6678);
nor U6912 (N_6912,N_6237,N_6244);
nand U6913 (N_6913,N_6650,N_6594);
nand U6914 (N_6914,N_6547,N_6040);
and U6915 (N_6915,N_6632,N_6126);
nand U6916 (N_6916,N_6190,N_6643);
xnor U6917 (N_6917,N_6074,N_6239);
xnor U6918 (N_6918,N_6245,N_6142);
nand U6919 (N_6919,N_6031,N_6092);
or U6920 (N_6920,N_6037,N_6225);
nor U6921 (N_6921,N_6191,N_6510);
or U6922 (N_6922,N_6312,N_6112);
or U6923 (N_6923,N_6159,N_6131);
nand U6924 (N_6924,N_6681,N_6008);
xnor U6925 (N_6925,N_6006,N_6536);
or U6926 (N_6926,N_6525,N_6013);
nand U6927 (N_6927,N_6593,N_6426);
nor U6928 (N_6928,N_6725,N_6067);
nand U6929 (N_6929,N_6379,N_6135);
and U6930 (N_6930,N_6701,N_6730);
xor U6931 (N_6931,N_6200,N_6546);
nand U6932 (N_6932,N_6330,N_6630);
xor U6933 (N_6933,N_6232,N_6326);
and U6934 (N_6934,N_6535,N_6122);
or U6935 (N_6935,N_6500,N_6577);
and U6936 (N_6936,N_6359,N_6188);
and U6937 (N_6937,N_6511,N_6374);
or U6938 (N_6938,N_6745,N_6394);
nand U6939 (N_6939,N_6304,N_6445);
and U6940 (N_6940,N_6390,N_6641);
and U6941 (N_6941,N_6265,N_6167);
nor U6942 (N_6942,N_6320,N_6527);
xnor U6943 (N_6943,N_6340,N_6116);
nand U6944 (N_6944,N_6365,N_6468);
nand U6945 (N_6945,N_6220,N_6278);
xor U6946 (N_6946,N_6734,N_6174);
and U6947 (N_6947,N_6683,N_6099);
or U6948 (N_6948,N_6236,N_6571);
and U6949 (N_6949,N_6561,N_6348);
and U6950 (N_6950,N_6233,N_6043);
xnor U6951 (N_6951,N_6257,N_6033);
and U6952 (N_6952,N_6550,N_6373);
and U6953 (N_6953,N_6197,N_6121);
nand U6954 (N_6954,N_6459,N_6457);
xnor U6955 (N_6955,N_6367,N_6614);
nor U6956 (N_6956,N_6098,N_6575);
or U6957 (N_6957,N_6054,N_6591);
and U6958 (N_6958,N_6486,N_6717);
xor U6959 (N_6959,N_6680,N_6639);
and U6960 (N_6960,N_6551,N_6186);
xor U6961 (N_6961,N_6564,N_6319);
or U6962 (N_6962,N_6352,N_6368);
and U6963 (N_6963,N_6638,N_6652);
nor U6964 (N_6964,N_6572,N_6254);
xor U6965 (N_6965,N_6139,N_6289);
and U6966 (N_6966,N_6002,N_6327);
or U6967 (N_6967,N_6712,N_6048);
nand U6968 (N_6968,N_6726,N_6129);
or U6969 (N_6969,N_6421,N_6380);
xor U6970 (N_6970,N_6402,N_6691);
and U6971 (N_6971,N_6168,N_6281);
and U6972 (N_6972,N_6718,N_6276);
xor U6973 (N_6973,N_6277,N_6353);
nand U6974 (N_6974,N_6444,N_6313);
xor U6975 (N_6975,N_6310,N_6463);
xor U6976 (N_6976,N_6528,N_6275);
nor U6977 (N_6977,N_6422,N_6559);
nor U6978 (N_6978,N_6295,N_6047);
nand U6979 (N_6979,N_6472,N_6720);
or U6980 (N_6980,N_6125,N_6620);
or U6981 (N_6981,N_6093,N_6042);
nand U6982 (N_6982,N_6735,N_6150);
and U6983 (N_6983,N_6058,N_6635);
nand U6984 (N_6984,N_6140,N_6669);
nand U6985 (N_6985,N_6347,N_6660);
nor U6986 (N_6986,N_6284,N_6106);
xor U6987 (N_6987,N_6541,N_6689);
nor U6988 (N_6988,N_6019,N_6479);
nand U6989 (N_6989,N_6230,N_6451);
and U6990 (N_6990,N_6440,N_6202);
nand U6991 (N_6991,N_6183,N_6334);
nand U6992 (N_6992,N_6035,N_6316);
nor U6993 (N_6993,N_6655,N_6533);
nand U6994 (N_6994,N_6590,N_6026);
nor U6995 (N_6995,N_6508,N_6539);
xor U6996 (N_6996,N_6711,N_6668);
nand U6997 (N_6997,N_6407,N_6238);
or U6998 (N_6998,N_6644,N_6166);
and U6999 (N_6999,N_6469,N_6623);
nor U7000 (N_7000,N_6318,N_6083);
and U7001 (N_7001,N_6724,N_6206);
xnor U7002 (N_7002,N_6021,N_6000);
xnor U7003 (N_7003,N_6628,N_6366);
xnor U7004 (N_7004,N_6456,N_6499);
xnor U7005 (N_7005,N_6448,N_6070);
nor U7006 (N_7006,N_6181,N_6128);
or U7007 (N_7007,N_6071,N_6337);
xnor U7008 (N_7008,N_6205,N_6179);
or U7009 (N_7009,N_6586,N_6038);
xor U7010 (N_7010,N_6395,N_6172);
nor U7011 (N_7011,N_6516,N_6496);
nand U7012 (N_7012,N_6356,N_6124);
xor U7013 (N_7013,N_6292,N_6570);
xnor U7014 (N_7014,N_6165,N_6626);
and U7015 (N_7015,N_6314,N_6518);
and U7016 (N_7016,N_6007,N_6207);
and U7017 (N_7017,N_6016,N_6297);
xor U7018 (N_7018,N_6679,N_6148);
nor U7019 (N_7019,N_6009,N_6538);
or U7020 (N_7020,N_6716,N_6476);
nor U7021 (N_7021,N_6145,N_6062);
nand U7022 (N_7022,N_6151,N_6023);
and U7023 (N_7023,N_6267,N_6180);
and U7024 (N_7024,N_6437,N_6497);
or U7025 (N_7025,N_6025,N_6259);
nor U7026 (N_7026,N_6480,N_6077);
or U7027 (N_7027,N_6163,N_6467);
and U7028 (N_7028,N_6526,N_6335);
xnor U7029 (N_7029,N_6736,N_6715);
xor U7030 (N_7030,N_6531,N_6376);
and U7031 (N_7031,N_6732,N_6014);
xor U7032 (N_7032,N_6110,N_6324);
xor U7033 (N_7033,N_6378,N_6030);
nand U7034 (N_7034,N_6084,N_6264);
nand U7035 (N_7035,N_6041,N_6478);
nand U7036 (N_7036,N_6719,N_6358);
and U7037 (N_7037,N_6713,N_6565);
and U7038 (N_7038,N_6280,N_6355);
and U7039 (N_7039,N_6699,N_6240);
or U7040 (N_7040,N_6285,N_6698);
xnor U7041 (N_7041,N_6229,N_6076);
nand U7042 (N_7042,N_6481,N_6661);
xnor U7043 (N_7043,N_6512,N_6544);
or U7044 (N_7044,N_6223,N_6079);
nor U7045 (N_7045,N_6299,N_6671);
xnor U7046 (N_7046,N_6119,N_6708);
xor U7047 (N_7047,N_6441,N_6255);
and U7048 (N_7048,N_6246,N_6446);
and U7049 (N_7049,N_6032,N_6737);
or U7050 (N_7050,N_6595,N_6392);
xnor U7051 (N_7051,N_6184,N_6393);
nand U7052 (N_7052,N_6111,N_6344);
nand U7053 (N_7053,N_6455,N_6192);
nor U7054 (N_7054,N_6176,N_6169);
nand U7055 (N_7055,N_6589,N_6579);
or U7056 (N_7056,N_6642,N_6193);
and U7057 (N_7057,N_6325,N_6611);
or U7058 (N_7058,N_6185,N_6315);
and U7059 (N_7059,N_6039,N_6017);
nor U7060 (N_7060,N_6416,N_6080);
nor U7061 (N_7061,N_6609,N_6464);
or U7062 (N_7062,N_6592,N_6388);
nor U7063 (N_7063,N_6475,N_6235);
nor U7064 (N_7064,N_6581,N_6557);
xor U7065 (N_7065,N_6662,N_6370);
or U7066 (N_7066,N_6432,N_6061);
nand U7067 (N_7067,N_6410,N_6667);
nor U7068 (N_7068,N_6633,N_6108);
xnor U7069 (N_7069,N_6431,N_6317);
or U7070 (N_7070,N_6417,N_6601);
and U7071 (N_7071,N_6001,N_6109);
xnor U7072 (N_7072,N_6242,N_6542);
nor U7073 (N_7073,N_6600,N_6147);
or U7074 (N_7074,N_6034,N_6053);
nand U7075 (N_7075,N_6387,N_6616);
nor U7076 (N_7076,N_6369,N_6560);
nand U7077 (N_7077,N_6296,N_6305);
nor U7078 (N_7078,N_6747,N_6646);
nor U7079 (N_7079,N_6744,N_6663);
nor U7080 (N_7080,N_6506,N_6648);
and U7081 (N_7081,N_6024,N_6249);
nor U7082 (N_7082,N_6311,N_6351);
and U7083 (N_7083,N_6336,N_6322);
nand U7084 (N_7084,N_6612,N_6474);
nand U7085 (N_7085,N_6743,N_6674);
nor U7086 (N_7086,N_6272,N_6262);
nor U7087 (N_7087,N_6710,N_6127);
nand U7088 (N_7088,N_6429,N_6138);
xnor U7089 (N_7089,N_6199,N_6692);
and U7090 (N_7090,N_6398,N_6442);
or U7091 (N_7091,N_6400,N_6144);
nand U7092 (N_7092,N_6044,N_6610);
nand U7093 (N_7093,N_6243,N_6154);
xor U7094 (N_7094,N_6022,N_6484);
or U7095 (N_7095,N_6702,N_6576);
xnor U7096 (N_7096,N_6120,N_6696);
and U7097 (N_7097,N_6552,N_6515);
or U7098 (N_7098,N_6069,N_6537);
xor U7099 (N_7099,N_6270,N_6341);
and U7100 (N_7100,N_6473,N_6548);
or U7101 (N_7101,N_6503,N_6532);
nand U7102 (N_7102,N_6068,N_6530);
or U7103 (N_7103,N_6307,N_6494);
or U7104 (N_7104,N_6582,N_6049);
xnor U7105 (N_7105,N_6562,N_6585);
nand U7106 (N_7106,N_6222,N_6705);
and U7107 (N_7107,N_6073,N_6654);
or U7108 (N_7108,N_6493,N_6602);
xor U7109 (N_7109,N_6449,N_6156);
and U7110 (N_7110,N_6428,N_6673);
xnor U7111 (N_7111,N_6543,N_6622);
nor U7112 (N_7112,N_6171,N_6087);
nand U7113 (N_7113,N_6346,N_6178);
xnor U7114 (N_7114,N_6677,N_6709);
nand U7115 (N_7115,N_6485,N_6566);
and U7116 (N_7116,N_6477,N_6492);
nand U7117 (N_7117,N_6104,N_6413);
or U7118 (N_7118,N_6690,N_6102);
or U7119 (N_7119,N_6697,N_6143);
nor U7120 (N_7120,N_6290,N_6268);
nand U7121 (N_7121,N_6427,N_6383);
or U7122 (N_7122,N_6540,N_6399);
or U7123 (N_7123,N_6693,N_6342);
and U7124 (N_7124,N_6012,N_6333);
and U7125 (N_7125,N_6324,N_6354);
and U7126 (N_7126,N_6672,N_6383);
nor U7127 (N_7127,N_6385,N_6330);
nor U7128 (N_7128,N_6107,N_6726);
nand U7129 (N_7129,N_6601,N_6220);
nand U7130 (N_7130,N_6421,N_6726);
nand U7131 (N_7131,N_6409,N_6325);
or U7132 (N_7132,N_6233,N_6610);
or U7133 (N_7133,N_6053,N_6278);
nor U7134 (N_7134,N_6391,N_6394);
and U7135 (N_7135,N_6454,N_6436);
nor U7136 (N_7136,N_6217,N_6289);
and U7137 (N_7137,N_6160,N_6632);
or U7138 (N_7138,N_6557,N_6477);
or U7139 (N_7139,N_6671,N_6393);
nand U7140 (N_7140,N_6322,N_6618);
xnor U7141 (N_7141,N_6723,N_6277);
nor U7142 (N_7142,N_6463,N_6625);
or U7143 (N_7143,N_6355,N_6171);
xor U7144 (N_7144,N_6370,N_6499);
xnor U7145 (N_7145,N_6045,N_6192);
and U7146 (N_7146,N_6440,N_6589);
nand U7147 (N_7147,N_6510,N_6397);
nand U7148 (N_7148,N_6389,N_6551);
nor U7149 (N_7149,N_6063,N_6571);
and U7150 (N_7150,N_6663,N_6081);
and U7151 (N_7151,N_6200,N_6227);
or U7152 (N_7152,N_6344,N_6123);
nand U7153 (N_7153,N_6615,N_6186);
and U7154 (N_7154,N_6438,N_6052);
nor U7155 (N_7155,N_6101,N_6367);
nand U7156 (N_7156,N_6397,N_6591);
or U7157 (N_7157,N_6065,N_6195);
or U7158 (N_7158,N_6261,N_6694);
nor U7159 (N_7159,N_6632,N_6012);
and U7160 (N_7160,N_6673,N_6422);
xor U7161 (N_7161,N_6314,N_6009);
nor U7162 (N_7162,N_6380,N_6702);
and U7163 (N_7163,N_6712,N_6083);
and U7164 (N_7164,N_6398,N_6412);
and U7165 (N_7165,N_6723,N_6462);
xnor U7166 (N_7166,N_6379,N_6657);
nand U7167 (N_7167,N_6069,N_6039);
nor U7168 (N_7168,N_6702,N_6364);
xor U7169 (N_7169,N_6062,N_6343);
nor U7170 (N_7170,N_6397,N_6449);
nand U7171 (N_7171,N_6182,N_6094);
and U7172 (N_7172,N_6241,N_6103);
nand U7173 (N_7173,N_6160,N_6059);
or U7174 (N_7174,N_6382,N_6668);
or U7175 (N_7175,N_6274,N_6361);
nand U7176 (N_7176,N_6562,N_6364);
and U7177 (N_7177,N_6641,N_6161);
nor U7178 (N_7178,N_6219,N_6262);
or U7179 (N_7179,N_6344,N_6503);
xor U7180 (N_7180,N_6571,N_6727);
nand U7181 (N_7181,N_6311,N_6608);
and U7182 (N_7182,N_6633,N_6180);
or U7183 (N_7183,N_6261,N_6276);
or U7184 (N_7184,N_6550,N_6182);
or U7185 (N_7185,N_6736,N_6372);
xnor U7186 (N_7186,N_6347,N_6747);
and U7187 (N_7187,N_6489,N_6038);
or U7188 (N_7188,N_6014,N_6119);
xnor U7189 (N_7189,N_6176,N_6600);
xnor U7190 (N_7190,N_6334,N_6156);
nor U7191 (N_7191,N_6000,N_6709);
nand U7192 (N_7192,N_6654,N_6441);
nand U7193 (N_7193,N_6602,N_6296);
and U7194 (N_7194,N_6722,N_6357);
nand U7195 (N_7195,N_6240,N_6533);
nand U7196 (N_7196,N_6074,N_6183);
xor U7197 (N_7197,N_6635,N_6717);
xnor U7198 (N_7198,N_6325,N_6695);
nand U7199 (N_7199,N_6675,N_6149);
or U7200 (N_7200,N_6380,N_6169);
nand U7201 (N_7201,N_6576,N_6380);
nor U7202 (N_7202,N_6709,N_6445);
xnor U7203 (N_7203,N_6391,N_6132);
nand U7204 (N_7204,N_6014,N_6451);
and U7205 (N_7205,N_6056,N_6088);
xnor U7206 (N_7206,N_6096,N_6321);
nor U7207 (N_7207,N_6517,N_6605);
xnor U7208 (N_7208,N_6456,N_6028);
nor U7209 (N_7209,N_6541,N_6635);
nand U7210 (N_7210,N_6299,N_6148);
nand U7211 (N_7211,N_6521,N_6379);
nor U7212 (N_7212,N_6106,N_6483);
nor U7213 (N_7213,N_6195,N_6618);
nor U7214 (N_7214,N_6282,N_6472);
and U7215 (N_7215,N_6378,N_6570);
nand U7216 (N_7216,N_6647,N_6346);
nor U7217 (N_7217,N_6594,N_6663);
xor U7218 (N_7218,N_6591,N_6595);
xnor U7219 (N_7219,N_6209,N_6348);
nand U7220 (N_7220,N_6448,N_6238);
and U7221 (N_7221,N_6652,N_6347);
and U7222 (N_7222,N_6158,N_6131);
and U7223 (N_7223,N_6205,N_6294);
xnor U7224 (N_7224,N_6734,N_6071);
and U7225 (N_7225,N_6644,N_6048);
nor U7226 (N_7226,N_6713,N_6365);
nand U7227 (N_7227,N_6261,N_6389);
xnor U7228 (N_7228,N_6586,N_6292);
nand U7229 (N_7229,N_6002,N_6685);
nand U7230 (N_7230,N_6635,N_6658);
nand U7231 (N_7231,N_6593,N_6532);
and U7232 (N_7232,N_6182,N_6232);
nand U7233 (N_7233,N_6729,N_6474);
nand U7234 (N_7234,N_6447,N_6577);
or U7235 (N_7235,N_6065,N_6563);
nand U7236 (N_7236,N_6003,N_6434);
nor U7237 (N_7237,N_6156,N_6602);
or U7238 (N_7238,N_6671,N_6375);
nor U7239 (N_7239,N_6118,N_6734);
nand U7240 (N_7240,N_6144,N_6022);
or U7241 (N_7241,N_6535,N_6152);
nand U7242 (N_7242,N_6156,N_6680);
nor U7243 (N_7243,N_6075,N_6016);
or U7244 (N_7244,N_6646,N_6598);
and U7245 (N_7245,N_6402,N_6151);
and U7246 (N_7246,N_6566,N_6021);
nor U7247 (N_7247,N_6632,N_6046);
xor U7248 (N_7248,N_6395,N_6600);
and U7249 (N_7249,N_6417,N_6443);
nand U7250 (N_7250,N_6464,N_6060);
and U7251 (N_7251,N_6288,N_6108);
and U7252 (N_7252,N_6268,N_6343);
nand U7253 (N_7253,N_6447,N_6710);
nand U7254 (N_7254,N_6007,N_6371);
nor U7255 (N_7255,N_6233,N_6382);
and U7256 (N_7256,N_6262,N_6713);
xor U7257 (N_7257,N_6616,N_6106);
nor U7258 (N_7258,N_6270,N_6642);
xor U7259 (N_7259,N_6235,N_6001);
xor U7260 (N_7260,N_6423,N_6596);
and U7261 (N_7261,N_6180,N_6677);
xnor U7262 (N_7262,N_6103,N_6190);
or U7263 (N_7263,N_6346,N_6010);
nor U7264 (N_7264,N_6283,N_6170);
nor U7265 (N_7265,N_6489,N_6632);
nor U7266 (N_7266,N_6217,N_6578);
and U7267 (N_7267,N_6177,N_6345);
and U7268 (N_7268,N_6634,N_6464);
nor U7269 (N_7269,N_6581,N_6234);
and U7270 (N_7270,N_6380,N_6101);
xnor U7271 (N_7271,N_6482,N_6016);
or U7272 (N_7272,N_6116,N_6671);
nor U7273 (N_7273,N_6561,N_6603);
or U7274 (N_7274,N_6634,N_6298);
and U7275 (N_7275,N_6514,N_6054);
or U7276 (N_7276,N_6504,N_6342);
and U7277 (N_7277,N_6180,N_6229);
xnor U7278 (N_7278,N_6053,N_6535);
nand U7279 (N_7279,N_6284,N_6680);
or U7280 (N_7280,N_6275,N_6378);
xnor U7281 (N_7281,N_6018,N_6211);
and U7282 (N_7282,N_6025,N_6573);
nand U7283 (N_7283,N_6270,N_6715);
and U7284 (N_7284,N_6177,N_6741);
nand U7285 (N_7285,N_6633,N_6185);
nor U7286 (N_7286,N_6087,N_6485);
nand U7287 (N_7287,N_6070,N_6152);
or U7288 (N_7288,N_6030,N_6045);
nor U7289 (N_7289,N_6018,N_6366);
or U7290 (N_7290,N_6180,N_6659);
xnor U7291 (N_7291,N_6235,N_6162);
xor U7292 (N_7292,N_6330,N_6357);
xor U7293 (N_7293,N_6451,N_6437);
xor U7294 (N_7294,N_6650,N_6717);
nor U7295 (N_7295,N_6306,N_6441);
nand U7296 (N_7296,N_6135,N_6400);
nand U7297 (N_7297,N_6437,N_6384);
and U7298 (N_7298,N_6469,N_6725);
xnor U7299 (N_7299,N_6524,N_6416);
nand U7300 (N_7300,N_6270,N_6395);
nand U7301 (N_7301,N_6673,N_6278);
xnor U7302 (N_7302,N_6661,N_6402);
xor U7303 (N_7303,N_6717,N_6391);
or U7304 (N_7304,N_6119,N_6085);
or U7305 (N_7305,N_6505,N_6658);
or U7306 (N_7306,N_6239,N_6629);
and U7307 (N_7307,N_6207,N_6077);
or U7308 (N_7308,N_6117,N_6326);
xnor U7309 (N_7309,N_6699,N_6270);
nand U7310 (N_7310,N_6621,N_6217);
and U7311 (N_7311,N_6473,N_6064);
xnor U7312 (N_7312,N_6460,N_6511);
nand U7313 (N_7313,N_6689,N_6354);
xor U7314 (N_7314,N_6702,N_6625);
and U7315 (N_7315,N_6735,N_6251);
nand U7316 (N_7316,N_6011,N_6222);
nand U7317 (N_7317,N_6222,N_6436);
nor U7318 (N_7318,N_6305,N_6557);
nand U7319 (N_7319,N_6364,N_6194);
nor U7320 (N_7320,N_6244,N_6574);
xnor U7321 (N_7321,N_6196,N_6564);
xnor U7322 (N_7322,N_6536,N_6396);
and U7323 (N_7323,N_6221,N_6071);
and U7324 (N_7324,N_6323,N_6214);
or U7325 (N_7325,N_6046,N_6549);
xnor U7326 (N_7326,N_6264,N_6303);
xor U7327 (N_7327,N_6732,N_6292);
and U7328 (N_7328,N_6557,N_6128);
xnor U7329 (N_7329,N_6692,N_6368);
xnor U7330 (N_7330,N_6572,N_6566);
nand U7331 (N_7331,N_6631,N_6649);
or U7332 (N_7332,N_6694,N_6590);
and U7333 (N_7333,N_6081,N_6000);
or U7334 (N_7334,N_6397,N_6189);
nand U7335 (N_7335,N_6695,N_6501);
nand U7336 (N_7336,N_6060,N_6698);
xor U7337 (N_7337,N_6302,N_6570);
xor U7338 (N_7338,N_6038,N_6661);
xnor U7339 (N_7339,N_6265,N_6615);
nand U7340 (N_7340,N_6105,N_6319);
xor U7341 (N_7341,N_6222,N_6696);
or U7342 (N_7342,N_6640,N_6742);
or U7343 (N_7343,N_6340,N_6690);
nand U7344 (N_7344,N_6002,N_6694);
xor U7345 (N_7345,N_6198,N_6387);
nor U7346 (N_7346,N_6404,N_6619);
xor U7347 (N_7347,N_6398,N_6532);
nand U7348 (N_7348,N_6124,N_6418);
xnor U7349 (N_7349,N_6617,N_6644);
or U7350 (N_7350,N_6577,N_6717);
nor U7351 (N_7351,N_6137,N_6306);
and U7352 (N_7352,N_6644,N_6005);
and U7353 (N_7353,N_6335,N_6164);
and U7354 (N_7354,N_6137,N_6512);
or U7355 (N_7355,N_6128,N_6320);
nand U7356 (N_7356,N_6234,N_6651);
or U7357 (N_7357,N_6513,N_6393);
nor U7358 (N_7358,N_6090,N_6171);
xor U7359 (N_7359,N_6313,N_6493);
nand U7360 (N_7360,N_6611,N_6149);
nand U7361 (N_7361,N_6314,N_6512);
xnor U7362 (N_7362,N_6024,N_6600);
and U7363 (N_7363,N_6207,N_6292);
and U7364 (N_7364,N_6681,N_6725);
nand U7365 (N_7365,N_6325,N_6163);
nand U7366 (N_7366,N_6183,N_6739);
and U7367 (N_7367,N_6594,N_6279);
xor U7368 (N_7368,N_6646,N_6611);
nor U7369 (N_7369,N_6353,N_6288);
nand U7370 (N_7370,N_6490,N_6420);
xor U7371 (N_7371,N_6392,N_6643);
or U7372 (N_7372,N_6090,N_6395);
and U7373 (N_7373,N_6606,N_6300);
and U7374 (N_7374,N_6120,N_6504);
xnor U7375 (N_7375,N_6696,N_6244);
xor U7376 (N_7376,N_6730,N_6189);
and U7377 (N_7377,N_6666,N_6367);
nand U7378 (N_7378,N_6452,N_6203);
nor U7379 (N_7379,N_6056,N_6725);
xor U7380 (N_7380,N_6454,N_6399);
or U7381 (N_7381,N_6023,N_6439);
and U7382 (N_7382,N_6484,N_6443);
nor U7383 (N_7383,N_6212,N_6668);
xnor U7384 (N_7384,N_6736,N_6527);
and U7385 (N_7385,N_6078,N_6423);
xor U7386 (N_7386,N_6251,N_6178);
nand U7387 (N_7387,N_6338,N_6241);
xnor U7388 (N_7388,N_6345,N_6222);
and U7389 (N_7389,N_6527,N_6223);
or U7390 (N_7390,N_6694,N_6193);
xor U7391 (N_7391,N_6677,N_6321);
and U7392 (N_7392,N_6080,N_6352);
and U7393 (N_7393,N_6289,N_6384);
xor U7394 (N_7394,N_6705,N_6171);
nor U7395 (N_7395,N_6330,N_6125);
nand U7396 (N_7396,N_6613,N_6493);
nor U7397 (N_7397,N_6588,N_6458);
or U7398 (N_7398,N_6666,N_6580);
and U7399 (N_7399,N_6253,N_6236);
nor U7400 (N_7400,N_6645,N_6368);
and U7401 (N_7401,N_6226,N_6569);
or U7402 (N_7402,N_6728,N_6518);
xor U7403 (N_7403,N_6317,N_6542);
nor U7404 (N_7404,N_6427,N_6440);
nand U7405 (N_7405,N_6391,N_6435);
or U7406 (N_7406,N_6432,N_6480);
nand U7407 (N_7407,N_6352,N_6578);
nand U7408 (N_7408,N_6673,N_6060);
xor U7409 (N_7409,N_6412,N_6061);
nand U7410 (N_7410,N_6561,N_6291);
nand U7411 (N_7411,N_6429,N_6533);
and U7412 (N_7412,N_6498,N_6678);
and U7413 (N_7413,N_6451,N_6365);
and U7414 (N_7414,N_6713,N_6273);
xor U7415 (N_7415,N_6532,N_6534);
or U7416 (N_7416,N_6746,N_6421);
xor U7417 (N_7417,N_6549,N_6162);
and U7418 (N_7418,N_6498,N_6392);
nand U7419 (N_7419,N_6265,N_6580);
and U7420 (N_7420,N_6368,N_6216);
or U7421 (N_7421,N_6219,N_6519);
and U7422 (N_7422,N_6332,N_6052);
xnor U7423 (N_7423,N_6206,N_6214);
xnor U7424 (N_7424,N_6530,N_6329);
and U7425 (N_7425,N_6697,N_6212);
nor U7426 (N_7426,N_6713,N_6655);
or U7427 (N_7427,N_6159,N_6199);
nor U7428 (N_7428,N_6347,N_6592);
xnor U7429 (N_7429,N_6349,N_6408);
xor U7430 (N_7430,N_6247,N_6701);
xnor U7431 (N_7431,N_6567,N_6317);
and U7432 (N_7432,N_6201,N_6455);
xor U7433 (N_7433,N_6555,N_6317);
nor U7434 (N_7434,N_6724,N_6470);
xnor U7435 (N_7435,N_6033,N_6469);
or U7436 (N_7436,N_6587,N_6416);
xor U7437 (N_7437,N_6274,N_6696);
xor U7438 (N_7438,N_6636,N_6743);
or U7439 (N_7439,N_6551,N_6313);
and U7440 (N_7440,N_6587,N_6401);
nor U7441 (N_7441,N_6648,N_6680);
and U7442 (N_7442,N_6239,N_6538);
nor U7443 (N_7443,N_6206,N_6475);
xnor U7444 (N_7444,N_6400,N_6072);
and U7445 (N_7445,N_6193,N_6026);
nor U7446 (N_7446,N_6447,N_6022);
nand U7447 (N_7447,N_6321,N_6521);
or U7448 (N_7448,N_6295,N_6331);
or U7449 (N_7449,N_6742,N_6138);
and U7450 (N_7450,N_6346,N_6576);
and U7451 (N_7451,N_6408,N_6448);
nand U7452 (N_7452,N_6665,N_6249);
or U7453 (N_7453,N_6727,N_6275);
xor U7454 (N_7454,N_6363,N_6277);
xor U7455 (N_7455,N_6679,N_6009);
and U7456 (N_7456,N_6240,N_6722);
or U7457 (N_7457,N_6471,N_6443);
xor U7458 (N_7458,N_6356,N_6204);
and U7459 (N_7459,N_6140,N_6229);
or U7460 (N_7460,N_6548,N_6091);
and U7461 (N_7461,N_6129,N_6109);
and U7462 (N_7462,N_6439,N_6252);
nand U7463 (N_7463,N_6025,N_6515);
nand U7464 (N_7464,N_6314,N_6017);
or U7465 (N_7465,N_6114,N_6510);
or U7466 (N_7466,N_6277,N_6283);
nand U7467 (N_7467,N_6037,N_6095);
and U7468 (N_7468,N_6558,N_6345);
and U7469 (N_7469,N_6348,N_6468);
or U7470 (N_7470,N_6743,N_6370);
nor U7471 (N_7471,N_6591,N_6727);
nand U7472 (N_7472,N_6537,N_6507);
nor U7473 (N_7473,N_6135,N_6720);
nand U7474 (N_7474,N_6398,N_6178);
nand U7475 (N_7475,N_6123,N_6587);
or U7476 (N_7476,N_6449,N_6000);
nand U7477 (N_7477,N_6530,N_6693);
nand U7478 (N_7478,N_6085,N_6488);
xnor U7479 (N_7479,N_6735,N_6359);
nand U7480 (N_7480,N_6251,N_6443);
and U7481 (N_7481,N_6206,N_6703);
and U7482 (N_7482,N_6597,N_6407);
nand U7483 (N_7483,N_6081,N_6336);
and U7484 (N_7484,N_6306,N_6271);
and U7485 (N_7485,N_6077,N_6436);
and U7486 (N_7486,N_6141,N_6607);
or U7487 (N_7487,N_6675,N_6089);
xor U7488 (N_7488,N_6052,N_6547);
nor U7489 (N_7489,N_6081,N_6591);
nand U7490 (N_7490,N_6628,N_6571);
nor U7491 (N_7491,N_6703,N_6077);
and U7492 (N_7492,N_6645,N_6746);
or U7493 (N_7493,N_6083,N_6139);
or U7494 (N_7494,N_6104,N_6195);
or U7495 (N_7495,N_6386,N_6493);
and U7496 (N_7496,N_6525,N_6741);
nand U7497 (N_7497,N_6676,N_6703);
and U7498 (N_7498,N_6134,N_6208);
xor U7499 (N_7499,N_6370,N_6633);
nor U7500 (N_7500,N_6881,N_7061);
and U7501 (N_7501,N_7087,N_7469);
nand U7502 (N_7502,N_7324,N_7113);
and U7503 (N_7503,N_7107,N_7382);
nand U7504 (N_7504,N_7139,N_7017);
and U7505 (N_7505,N_7037,N_7339);
and U7506 (N_7506,N_7237,N_7003);
xnor U7507 (N_7507,N_7493,N_6926);
and U7508 (N_7508,N_6823,N_6831);
nor U7509 (N_7509,N_7497,N_7335);
nand U7510 (N_7510,N_6768,N_6947);
and U7511 (N_7511,N_7246,N_6878);
or U7512 (N_7512,N_6877,N_7453);
or U7513 (N_7513,N_7386,N_7196);
nor U7514 (N_7514,N_7072,N_6794);
nor U7515 (N_7515,N_7083,N_6764);
or U7516 (N_7516,N_6851,N_6889);
nor U7517 (N_7517,N_6817,N_7004);
and U7518 (N_7518,N_6999,N_7308);
xor U7519 (N_7519,N_6939,N_7240);
and U7520 (N_7520,N_7202,N_7250);
or U7521 (N_7521,N_7403,N_7415);
nand U7522 (N_7522,N_6954,N_7350);
or U7523 (N_7523,N_7440,N_7082);
or U7524 (N_7524,N_7394,N_7180);
and U7525 (N_7525,N_7219,N_7454);
xor U7526 (N_7526,N_6995,N_6998);
nand U7527 (N_7527,N_6990,N_6825);
and U7528 (N_7528,N_7269,N_6952);
nor U7529 (N_7529,N_6989,N_7381);
xor U7530 (N_7530,N_6997,N_7281);
nand U7531 (N_7531,N_7424,N_6812);
and U7532 (N_7532,N_7292,N_6972);
xnor U7533 (N_7533,N_6946,N_6876);
or U7534 (N_7534,N_7295,N_7023);
xor U7535 (N_7535,N_7106,N_7307);
and U7536 (N_7536,N_7168,N_6949);
xnor U7537 (N_7537,N_7176,N_7442);
and U7538 (N_7538,N_7228,N_7336);
and U7539 (N_7539,N_6922,N_7383);
or U7540 (N_7540,N_6879,N_6897);
nor U7541 (N_7541,N_6777,N_7195);
nor U7542 (N_7542,N_6916,N_7310);
nand U7543 (N_7543,N_6907,N_7096);
nor U7544 (N_7544,N_7368,N_7192);
nor U7545 (N_7545,N_6892,N_7416);
nor U7546 (N_7546,N_7319,N_7490);
xor U7547 (N_7547,N_7052,N_7256);
xnor U7548 (N_7548,N_7038,N_6928);
and U7549 (N_7549,N_7094,N_7133);
xnor U7550 (N_7550,N_7156,N_7387);
and U7551 (N_7551,N_6938,N_7108);
and U7552 (N_7552,N_6918,N_6941);
nand U7553 (N_7553,N_6903,N_7182);
nand U7554 (N_7554,N_7422,N_7337);
nor U7555 (N_7555,N_7464,N_6940);
xor U7556 (N_7556,N_7402,N_7364);
or U7557 (N_7557,N_7400,N_6860);
xor U7558 (N_7558,N_7258,N_6959);
or U7559 (N_7559,N_7011,N_7363);
or U7560 (N_7560,N_7448,N_6987);
or U7561 (N_7561,N_7486,N_6834);
nand U7562 (N_7562,N_7432,N_7272);
nand U7563 (N_7563,N_7078,N_6791);
or U7564 (N_7564,N_7474,N_7296);
nor U7565 (N_7565,N_7122,N_6833);
and U7566 (N_7566,N_7489,N_6988);
and U7567 (N_7567,N_6932,N_7342);
and U7568 (N_7568,N_7009,N_7357);
nand U7569 (N_7569,N_7012,N_6762);
or U7570 (N_7570,N_7391,N_7210);
and U7571 (N_7571,N_7217,N_7457);
nand U7572 (N_7572,N_7375,N_6857);
or U7573 (N_7573,N_6865,N_7356);
nand U7574 (N_7574,N_7254,N_6775);
nor U7575 (N_7575,N_7251,N_6870);
or U7576 (N_7576,N_6930,N_6837);
and U7577 (N_7577,N_6969,N_6757);
nand U7578 (N_7578,N_7073,N_6809);
nand U7579 (N_7579,N_6773,N_7185);
xnor U7580 (N_7580,N_7317,N_7321);
and U7581 (N_7581,N_7232,N_6974);
and U7582 (N_7582,N_6891,N_7160);
nor U7583 (N_7583,N_7441,N_6818);
xnor U7584 (N_7584,N_6758,N_6951);
nor U7585 (N_7585,N_6943,N_7499);
and U7586 (N_7586,N_7456,N_7111);
and U7587 (N_7587,N_7066,N_7397);
or U7588 (N_7588,N_6867,N_6802);
or U7589 (N_7589,N_6761,N_7124);
nor U7590 (N_7590,N_7380,N_7206);
or U7591 (N_7591,N_6886,N_7230);
xnor U7592 (N_7592,N_7148,N_7408);
nor U7593 (N_7593,N_7042,N_6968);
and U7594 (N_7594,N_7188,N_7374);
or U7595 (N_7595,N_6981,N_6856);
nor U7596 (N_7596,N_6958,N_6953);
nand U7597 (N_7597,N_7496,N_7393);
and U7598 (N_7598,N_6829,N_7145);
or U7599 (N_7599,N_6986,N_7290);
xnor U7600 (N_7600,N_7134,N_7132);
xor U7601 (N_7601,N_7159,N_7277);
xor U7602 (N_7602,N_7425,N_7092);
or U7603 (N_7603,N_7103,N_6979);
nand U7604 (N_7604,N_6788,N_7262);
or U7605 (N_7605,N_6843,N_7158);
nor U7606 (N_7606,N_6854,N_6924);
xor U7607 (N_7607,N_6832,N_6795);
or U7608 (N_7608,N_7478,N_7190);
and U7609 (N_7609,N_7430,N_7049);
xor U7610 (N_7610,N_7329,N_6950);
and U7611 (N_7611,N_7167,N_7117);
and U7612 (N_7612,N_6824,N_7181);
nor U7613 (N_7613,N_7164,N_6753);
xnor U7614 (N_7614,N_7309,N_6971);
nand U7615 (N_7615,N_7326,N_6967);
or U7616 (N_7616,N_7385,N_6973);
nand U7617 (N_7617,N_6965,N_7431);
nand U7618 (N_7618,N_7153,N_7455);
nand U7619 (N_7619,N_7179,N_6931);
and U7620 (N_7620,N_7089,N_7332);
nor U7621 (N_7621,N_7389,N_7349);
and U7622 (N_7622,N_7227,N_7119);
xor U7623 (N_7623,N_7125,N_6769);
or U7624 (N_7624,N_7421,N_6970);
nor U7625 (N_7625,N_7071,N_6806);
and U7626 (N_7626,N_7068,N_6838);
or U7627 (N_7627,N_7032,N_7294);
nand U7628 (N_7628,N_7014,N_7175);
and U7629 (N_7629,N_7404,N_6982);
or U7630 (N_7630,N_6944,N_7299);
nor U7631 (N_7631,N_7039,N_7316);
or U7632 (N_7632,N_7472,N_6895);
nand U7633 (N_7633,N_7361,N_6814);
or U7634 (N_7634,N_6792,N_7495);
xnor U7635 (N_7635,N_7418,N_7468);
nor U7636 (N_7636,N_7165,N_7412);
xor U7637 (N_7637,N_6925,N_7247);
nand U7638 (N_7638,N_7451,N_6799);
nand U7639 (N_7639,N_6759,N_7002);
or U7640 (N_7640,N_7305,N_7216);
nand U7641 (N_7641,N_7150,N_7201);
nor U7642 (N_7642,N_7477,N_6934);
nand U7643 (N_7643,N_7476,N_6885);
nor U7644 (N_7644,N_7444,N_7110);
xnor U7645 (N_7645,N_7370,N_7064);
or U7646 (N_7646,N_6836,N_7013);
xnor U7647 (N_7647,N_7452,N_7030);
nor U7648 (N_7648,N_7234,N_7088);
nand U7649 (N_7649,N_7396,N_7019);
nand U7650 (N_7650,N_7183,N_7118);
xnor U7651 (N_7651,N_7483,N_7213);
xor U7652 (N_7652,N_6905,N_6816);
and U7653 (N_7653,N_7470,N_7366);
or U7654 (N_7654,N_6868,N_6779);
nand U7655 (N_7655,N_7369,N_7434);
or U7656 (N_7656,N_7304,N_7267);
or U7657 (N_7657,N_7214,N_7320);
xor U7658 (N_7658,N_7266,N_7065);
or U7659 (N_7659,N_7263,N_7419);
xor U7660 (N_7660,N_7261,N_7498);
and U7661 (N_7661,N_6790,N_7312);
nand U7662 (N_7662,N_6765,N_7407);
nand U7663 (N_7663,N_7149,N_7458);
and U7664 (N_7664,N_7016,N_6751);
nand U7665 (N_7665,N_7428,N_7031);
nor U7666 (N_7666,N_6923,N_7325);
nor U7667 (N_7667,N_7084,N_7270);
and U7668 (N_7668,N_7318,N_7252);
nand U7669 (N_7669,N_7053,N_6778);
xnor U7670 (N_7670,N_6936,N_7447);
nand U7671 (N_7671,N_7438,N_6977);
xor U7672 (N_7672,N_6789,N_7093);
and U7673 (N_7673,N_7095,N_7466);
nand U7674 (N_7674,N_7146,N_7467);
nor U7675 (N_7675,N_7220,N_7022);
nand U7676 (N_7676,N_7492,N_7398);
or U7677 (N_7677,N_7200,N_7315);
nor U7678 (N_7678,N_7359,N_6909);
and U7679 (N_7679,N_7186,N_7427);
nor U7680 (N_7680,N_7482,N_7257);
nor U7681 (N_7681,N_7208,N_7475);
or U7682 (N_7682,N_7353,N_7395);
and U7683 (N_7683,N_7047,N_7136);
nor U7684 (N_7684,N_6828,N_6913);
nand U7685 (N_7685,N_6811,N_7311);
xnor U7686 (N_7686,N_6798,N_6820);
nand U7687 (N_7687,N_7449,N_7226);
and U7688 (N_7688,N_7172,N_7401);
and U7689 (N_7689,N_7115,N_7046);
xnor U7690 (N_7690,N_7334,N_7100);
nor U7691 (N_7691,N_6850,N_6840);
xnor U7692 (N_7692,N_7399,N_7333);
nand U7693 (N_7693,N_7191,N_7301);
nand U7694 (N_7694,N_7450,N_7021);
nor U7695 (N_7695,N_7135,N_7097);
nor U7696 (N_7696,N_6776,N_7354);
and U7697 (N_7697,N_7352,N_6869);
xor U7698 (N_7698,N_7373,N_6933);
and U7699 (N_7699,N_7035,N_7140);
nand U7700 (N_7700,N_6872,N_6772);
nand U7701 (N_7701,N_7062,N_6962);
xnor U7702 (N_7702,N_7233,N_6849);
nor U7703 (N_7703,N_6894,N_7367);
and U7704 (N_7704,N_6937,N_6774);
and U7705 (N_7705,N_7417,N_7372);
or U7706 (N_7706,N_7152,N_7236);
and U7707 (N_7707,N_7487,N_6844);
or U7708 (N_7708,N_7081,N_7379);
nand U7709 (N_7709,N_7147,N_7051);
and U7710 (N_7710,N_7341,N_7287);
xnor U7711 (N_7711,N_7224,N_6893);
and U7712 (N_7712,N_6985,N_7443);
nand U7713 (N_7713,N_6861,N_6984);
xor U7714 (N_7714,N_7043,N_7048);
nand U7715 (N_7715,N_6917,N_7184);
nor U7716 (N_7716,N_7435,N_6935);
nand U7717 (N_7717,N_7209,N_7197);
or U7718 (N_7718,N_7239,N_7223);
and U7719 (N_7719,N_7086,N_6900);
or U7720 (N_7720,N_7291,N_6871);
nand U7721 (N_7721,N_7346,N_6752);
nor U7722 (N_7722,N_7436,N_6908);
nor U7723 (N_7723,N_6796,N_7285);
nor U7724 (N_7724,N_6848,N_7446);
xor U7725 (N_7725,N_6980,N_7300);
xnor U7726 (N_7726,N_6859,N_7059);
nor U7727 (N_7727,N_6785,N_7297);
or U7728 (N_7728,N_7406,N_6927);
nand U7729 (N_7729,N_7138,N_7055);
or U7730 (N_7730,N_7099,N_7008);
xnor U7731 (N_7731,N_7330,N_7365);
xor U7732 (N_7732,N_7314,N_6813);
nor U7733 (N_7733,N_6766,N_7041);
nand U7734 (N_7734,N_6873,N_6793);
nor U7735 (N_7735,N_7123,N_6942);
nand U7736 (N_7736,N_6992,N_6975);
or U7737 (N_7737,N_6781,N_6921);
xnor U7738 (N_7738,N_7222,N_7024);
xor U7739 (N_7739,N_6976,N_7491);
xnor U7740 (N_7740,N_6887,N_6963);
and U7741 (N_7741,N_7343,N_7127);
nor U7742 (N_7742,N_7289,N_7242);
nand U7743 (N_7743,N_7445,N_6884);
xnor U7744 (N_7744,N_6920,N_7433);
nand U7745 (N_7745,N_6902,N_7409);
nand U7746 (N_7746,N_7238,N_7479);
or U7747 (N_7747,N_7169,N_7144);
and U7748 (N_7748,N_7481,N_7225);
nor U7749 (N_7749,N_6906,N_7392);
xnor U7750 (N_7750,N_6945,N_6803);
nor U7751 (N_7751,N_7284,N_7276);
nor U7752 (N_7752,N_7141,N_7076);
nand U7753 (N_7753,N_7303,N_7207);
nand U7754 (N_7754,N_6929,N_7293);
nor U7755 (N_7755,N_6863,N_7338);
nor U7756 (N_7756,N_7171,N_7371);
nand U7757 (N_7757,N_7271,N_6862);
xor U7758 (N_7758,N_6842,N_7120);
xnor U7759 (N_7759,N_7126,N_7355);
nand U7760 (N_7760,N_6957,N_7007);
and U7761 (N_7761,N_6787,N_7488);
and U7762 (N_7762,N_6948,N_7040);
and U7763 (N_7763,N_7034,N_7077);
xnor U7764 (N_7764,N_6901,N_6955);
and U7765 (N_7765,N_7026,N_7029);
and U7766 (N_7766,N_7005,N_7215);
and U7767 (N_7767,N_6960,N_7460);
or U7768 (N_7768,N_7288,N_6910);
nand U7769 (N_7769,N_7161,N_7060);
and U7770 (N_7770,N_7025,N_7205);
or U7771 (N_7771,N_7426,N_6888);
or U7772 (N_7772,N_7260,N_7057);
nor U7773 (N_7773,N_7420,N_7033);
nand U7774 (N_7774,N_7116,N_7278);
and U7775 (N_7775,N_7104,N_6771);
or U7776 (N_7776,N_6750,N_6804);
xor U7777 (N_7777,N_7001,N_7105);
nand U7778 (N_7778,N_6835,N_6800);
or U7779 (N_7779,N_7485,N_7328);
nand U7780 (N_7780,N_7101,N_7235);
nand U7781 (N_7781,N_6864,N_7264);
nor U7782 (N_7782,N_7121,N_6801);
and U7783 (N_7783,N_6911,N_6883);
or U7784 (N_7784,N_7286,N_6808);
or U7785 (N_7785,N_7114,N_7274);
nor U7786 (N_7786,N_7162,N_6845);
nand U7787 (N_7787,N_7229,N_7198);
nor U7788 (N_7788,N_7348,N_7283);
and U7789 (N_7789,N_6770,N_7137);
and U7790 (N_7790,N_7098,N_7473);
or U7791 (N_7791,N_7465,N_6805);
nand U7792 (N_7792,N_7170,N_6853);
nand U7793 (N_7793,N_6882,N_7045);
or U7794 (N_7794,N_7471,N_7211);
or U7795 (N_7795,N_7282,N_7020);
or U7796 (N_7796,N_7405,N_7070);
or U7797 (N_7797,N_7362,N_7313);
nand U7798 (N_7798,N_7221,N_6797);
nand U7799 (N_7799,N_7218,N_7027);
nand U7800 (N_7800,N_7413,N_7378);
or U7801 (N_7801,N_7323,N_7010);
and U7802 (N_7802,N_7275,N_6756);
or U7803 (N_7803,N_6760,N_6755);
nor U7804 (N_7804,N_7463,N_7253);
or U7805 (N_7805,N_6890,N_7155);
nor U7806 (N_7806,N_6964,N_7298);
xnor U7807 (N_7807,N_7423,N_6846);
and U7808 (N_7808,N_6966,N_7331);
and U7809 (N_7809,N_6807,N_6912);
xor U7810 (N_7810,N_7265,N_7130);
nand U7811 (N_7811,N_7075,N_6898);
nor U7812 (N_7812,N_6810,N_7044);
xnor U7813 (N_7813,N_6780,N_6899);
and U7814 (N_7814,N_7128,N_7204);
nand U7815 (N_7815,N_7050,N_6914);
or U7816 (N_7816,N_7494,N_7036);
xor U7817 (N_7817,N_7280,N_7163);
nor U7818 (N_7818,N_7174,N_7484);
nor U7819 (N_7819,N_7273,N_6983);
and U7820 (N_7820,N_6821,N_6754);
nand U7821 (N_7821,N_6783,N_7249);
or U7822 (N_7822,N_6827,N_7203);
xnor U7823 (N_7823,N_6763,N_7112);
or U7824 (N_7824,N_7166,N_7245);
nand U7825 (N_7825,N_7410,N_6822);
and U7826 (N_7826,N_7255,N_6784);
nand U7827 (N_7827,N_7154,N_6782);
nor U7828 (N_7828,N_6978,N_6991);
xnor U7829 (N_7829,N_7344,N_7129);
or U7830 (N_7830,N_7079,N_7377);
or U7831 (N_7831,N_7178,N_7067);
xnor U7832 (N_7832,N_7390,N_7189);
nand U7833 (N_7833,N_7360,N_7259);
nor U7834 (N_7834,N_6994,N_7243);
and U7835 (N_7835,N_7461,N_7102);
and U7836 (N_7836,N_7091,N_7439);
or U7837 (N_7837,N_6915,N_6956);
xnor U7838 (N_7838,N_7028,N_6874);
nor U7839 (N_7839,N_7340,N_7358);
nand U7840 (N_7840,N_7327,N_7279);
nand U7841 (N_7841,N_7151,N_7462);
xnor U7842 (N_7842,N_6767,N_7376);
and U7843 (N_7843,N_7131,N_6880);
or U7844 (N_7844,N_7212,N_7069);
nand U7845 (N_7845,N_7015,N_7063);
nor U7846 (N_7846,N_7157,N_7437);
and U7847 (N_7847,N_7000,N_7018);
nand U7848 (N_7848,N_6815,N_7414);
and U7849 (N_7849,N_7177,N_7080);
xnor U7850 (N_7850,N_7345,N_6830);
and U7851 (N_7851,N_6858,N_7006);
nor U7852 (N_7852,N_7347,N_6839);
nor U7853 (N_7853,N_7187,N_6919);
nor U7854 (N_7854,N_7085,N_7411);
and U7855 (N_7855,N_6896,N_6875);
xor U7856 (N_7856,N_6904,N_7194);
xnor U7857 (N_7857,N_7074,N_7090);
nand U7858 (N_7858,N_6855,N_7268);
or U7859 (N_7859,N_7054,N_7193);
xor U7860 (N_7860,N_7322,N_7142);
and U7861 (N_7861,N_6866,N_7459);
nand U7862 (N_7862,N_7143,N_7248);
xor U7863 (N_7863,N_7480,N_6961);
xnor U7864 (N_7864,N_7429,N_7058);
xor U7865 (N_7865,N_6847,N_6852);
xnor U7866 (N_7866,N_6786,N_7231);
or U7867 (N_7867,N_7306,N_7056);
or U7868 (N_7868,N_7302,N_6841);
nor U7869 (N_7869,N_7199,N_6826);
nor U7870 (N_7870,N_7384,N_7388);
or U7871 (N_7871,N_7109,N_6996);
nand U7872 (N_7872,N_7351,N_6819);
xnor U7873 (N_7873,N_7173,N_6993);
nor U7874 (N_7874,N_7244,N_7241);
or U7875 (N_7875,N_6931,N_6935);
or U7876 (N_7876,N_6862,N_7337);
and U7877 (N_7877,N_7456,N_7039);
and U7878 (N_7878,N_7412,N_6779);
xnor U7879 (N_7879,N_7338,N_7255);
xnor U7880 (N_7880,N_7266,N_7252);
nor U7881 (N_7881,N_7158,N_6938);
nand U7882 (N_7882,N_7048,N_7231);
xor U7883 (N_7883,N_7104,N_6975);
xnor U7884 (N_7884,N_7061,N_7045);
xor U7885 (N_7885,N_7036,N_7462);
xor U7886 (N_7886,N_7094,N_7113);
and U7887 (N_7887,N_6883,N_6850);
or U7888 (N_7888,N_6770,N_6815);
and U7889 (N_7889,N_6991,N_6967);
xnor U7890 (N_7890,N_7153,N_7305);
xnor U7891 (N_7891,N_6866,N_6907);
and U7892 (N_7892,N_6942,N_7212);
xor U7893 (N_7893,N_6954,N_7106);
and U7894 (N_7894,N_7435,N_6989);
xnor U7895 (N_7895,N_7425,N_7417);
nand U7896 (N_7896,N_7337,N_7072);
and U7897 (N_7897,N_7041,N_6841);
nand U7898 (N_7898,N_7369,N_7278);
and U7899 (N_7899,N_6772,N_7403);
nand U7900 (N_7900,N_6951,N_7201);
and U7901 (N_7901,N_7119,N_7189);
nand U7902 (N_7902,N_7482,N_7304);
and U7903 (N_7903,N_7072,N_7429);
or U7904 (N_7904,N_6781,N_7119);
or U7905 (N_7905,N_7048,N_7461);
xor U7906 (N_7906,N_7238,N_7190);
xor U7907 (N_7907,N_7180,N_6951);
nor U7908 (N_7908,N_7462,N_6797);
xor U7909 (N_7909,N_7483,N_7153);
or U7910 (N_7910,N_7285,N_7312);
xnor U7911 (N_7911,N_7171,N_6788);
nand U7912 (N_7912,N_6892,N_6822);
or U7913 (N_7913,N_7420,N_7330);
nand U7914 (N_7914,N_7444,N_7494);
xor U7915 (N_7915,N_7318,N_7116);
nor U7916 (N_7916,N_7092,N_6900);
xor U7917 (N_7917,N_7016,N_7004);
nor U7918 (N_7918,N_7255,N_7479);
and U7919 (N_7919,N_7477,N_6804);
nand U7920 (N_7920,N_7497,N_6981);
nand U7921 (N_7921,N_7318,N_7398);
and U7922 (N_7922,N_7440,N_7413);
or U7923 (N_7923,N_7229,N_6991);
xnor U7924 (N_7924,N_7186,N_7359);
or U7925 (N_7925,N_6814,N_7313);
and U7926 (N_7926,N_6815,N_7461);
xor U7927 (N_7927,N_7427,N_6895);
nor U7928 (N_7928,N_6823,N_7251);
or U7929 (N_7929,N_7128,N_7165);
or U7930 (N_7930,N_7037,N_7077);
nor U7931 (N_7931,N_6793,N_6922);
and U7932 (N_7932,N_7418,N_7481);
nor U7933 (N_7933,N_7081,N_7071);
xor U7934 (N_7934,N_6782,N_7235);
nor U7935 (N_7935,N_6943,N_6989);
nor U7936 (N_7936,N_7379,N_6961);
nor U7937 (N_7937,N_7090,N_7475);
nor U7938 (N_7938,N_7203,N_7387);
nand U7939 (N_7939,N_6906,N_6806);
xnor U7940 (N_7940,N_7242,N_7390);
nand U7941 (N_7941,N_6869,N_6916);
xnor U7942 (N_7942,N_7465,N_7163);
or U7943 (N_7943,N_7246,N_7208);
or U7944 (N_7944,N_7491,N_7060);
or U7945 (N_7945,N_6865,N_7428);
or U7946 (N_7946,N_6763,N_7214);
xor U7947 (N_7947,N_7350,N_7362);
xnor U7948 (N_7948,N_6953,N_7253);
nand U7949 (N_7949,N_7223,N_7013);
or U7950 (N_7950,N_6995,N_6875);
xor U7951 (N_7951,N_7188,N_7419);
or U7952 (N_7952,N_7212,N_6967);
xnor U7953 (N_7953,N_7029,N_7254);
nand U7954 (N_7954,N_6845,N_6978);
nand U7955 (N_7955,N_7061,N_6832);
and U7956 (N_7956,N_7156,N_6819);
and U7957 (N_7957,N_7032,N_7491);
nand U7958 (N_7958,N_7201,N_7211);
and U7959 (N_7959,N_6863,N_7087);
nor U7960 (N_7960,N_7479,N_7394);
xnor U7961 (N_7961,N_7420,N_7276);
nand U7962 (N_7962,N_7302,N_7348);
nor U7963 (N_7963,N_7333,N_6891);
xnor U7964 (N_7964,N_6991,N_7460);
nand U7965 (N_7965,N_6832,N_7424);
or U7966 (N_7966,N_6757,N_7064);
nor U7967 (N_7967,N_6837,N_7365);
and U7968 (N_7968,N_7047,N_7057);
or U7969 (N_7969,N_7470,N_7096);
and U7970 (N_7970,N_7109,N_6802);
nor U7971 (N_7971,N_7407,N_7061);
nor U7972 (N_7972,N_7202,N_7085);
or U7973 (N_7973,N_7020,N_6795);
nor U7974 (N_7974,N_6936,N_7147);
and U7975 (N_7975,N_7297,N_6968);
nor U7976 (N_7976,N_7195,N_7146);
nand U7977 (N_7977,N_7110,N_7355);
or U7978 (N_7978,N_6840,N_7254);
and U7979 (N_7979,N_6849,N_6771);
nor U7980 (N_7980,N_7387,N_7064);
nand U7981 (N_7981,N_7152,N_6930);
xor U7982 (N_7982,N_7234,N_7482);
nand U7983 (N_7983,N_6778,N_6817);
or U7984 (N_7984,N_7441,N_7407);
nor U7985 (N_7985,N_7144,N_6818);
or U7986 (N_7986,N_6872,N_6943);
nand U7987 (N_7987,N_7045,N_7302);
or U7988 (N_7988,N_7159,N_6751);
nand U7989 (N_7989,N_6805,N_6980);
or U7990 (N_7990,N_7351,N_7147);
nor U7991 (N_7991,N_7450,N_7283);
or U7992 (N_7992,N_7094,N_7262);
and U7993 (N_7993,N_6790,N_7364);
or U7994 (N_7994,N_7190,N_7016);
xnor U7995 (N_7995,N_6999,N_7186);
and U7996 (N_7996,N_7404,N_6938);
xor U7997 (N_7997,N_6777,N_6943);
or U7998 (N_7998,N_7470,N_7431);
nand U7999 (N_7999,N_7189,N_7204);
xor U8000 (N_8000,N_6943,N_7121);
xnor U8001 (N_8001,N_7129,N_7154);
xnor U8002 (N_8002,N_7183,N_7144);
and U8003 (N_8003,N_7449,N_6901);
nor U8004 (N_8004,N_7358,N_7328);
xor U8005 (N_8005,N_7126,N_6835);
nand U8006 (N_8006,N_7253,N_7149);
xnor U8007 (N_8007,N_7330,N_6969);
nor U8008 (N_8008,N_6869,N_7350);
xnor U8009 (N_8009,N_7331,N_6956);
or U8010 (N_8010,N_7098,N_6944);
and U8011 (N_8011,N_7044,N_6849);
or U8012 (N_8012,N_6825,N_7270);
nor U8013 (N_8013,N_7446,N_6987);
xor U8014 (N_8014,N_6865,N_7197);
or U8015 (N_8015,N_7177,N_6915);
xor U8016 (N_8016,N_7102,N_6841);
nor U8017 (N_8017,N_7072,N_6812);
or U8018 (N_8018,N_7292,N_6893);
and U8019 (N_8019,N_6839,N_7024);
nor U8020 (N_8020,N_7404,N_7010);
or U8021 (N_8021,N_7339,N_7474);
nor U8022 (N_8022,N_7132,N_7200);
or U8023 (N_8023,N_7066,N_6877);
or U8024 (N_8024,N_7454,N_7214);
nand U8025 (N_8025,N_6839,N_7253);
xor U8026 (N_8026,N_6886,N_6850);
or U8027 (N_8027,N_7107,N_6931);
xor U8028 (N_8028,N_7059,N_6776);
or U8029 (N_8029,N_7206,N_7298);
and U8030 (N_8030,N_7053,N_7336);
nor U8031 (N_8031,N_6986,N_6779);
or U8032 (N_8032,N_6840,N_6891);
nand U8033 (N_8033,N_7485,N_6928);
nor U8034 (N_8034,N_6960,N_6976);
and U8035 (N_8035,N_7321,N_7244);
nor U8036 (N_8036,N_7046,N_6920);
and U8037 (N_8037,N_7062,N_7214);
xor U8038 (N_8038,N_6923,N_7407);
xnor U8039 (N_8039,N_7294,N_6780);
nor U8040 (N_8040,N_7164,N_6979);
xnor U8041 (N_8041,N_6910,N_7115);
or U8042 (N_8042,N_6758,N_7122);
or U8043 (N_8043,N_6869,N_7057);
nand U8044 (N_8044,N_7069,N_7235);
and U8045 (N_8045,N_6967,N_7043);
nand U8046 (N_8046,N_7343,N_7298);
xor U8047 (N_8047,N_7231,N_7316);
nor U8048 (N_8048,N_7483,N_7288);
nand U8049 (N_8049,N_7088,N_6929);
and U8050 (N_8050,N_7291,N_7143);
xnor U8051 (N_8051,N_7151,N_6789);
or U8052 (N_8052,N_6842,N_7296);
and U8053 (N_8053,N_7328,N_6974);
nor U8054 (N_8054,N_7251,N_7313);
nor U8055 (N_8055,N_6914,N_6984);
nor U8056 (N_8056,N_6863,N_6997);
xor U8057 (N_8057,N_6959,N_7390);
xor U8058 (N_8058,N_7200,N_7345);
nand U8059 (N_8059,N_6750,N_7092);
nand U8060 (N_8060,N_7066,N_6975);
xnor U8061 (N_8061,N_7242,N_7282);
nand U8062 (N_8062,N_7457,N_7495);
nand U8063 (N_8063,N_7444,N_6903);
nand U8064 (N_8064,N_6987,N_6896);
or U8065 (N_8065,N_7194,N_7466);
nor U8066 (N_8066,N_7338,N_7429);
and U8067 (N_8067,N_7138,N_7283);
xor U8068 (N_8068,N_7182,N_7427);
or U8069 (N_8069,N_6818,N_6935);
nor U8070 (N_8070,N_7308,N_6881);
nand U8071 (N_8071,N_7336,N_7233);
and U8072 (N_8072,N_7203,N_7072);
and U8073 (N_8073,N_6952,N_6931);
nand U8074 (N_8074,N_6913,N_6989);
or U8075 (N_8075,N_7254,N_6970);
or U8076 (N_8076,N_6777,N_6798);
nand U8077 (N_8077,N_7349,N_7145);
and U8078 (N_8078,N_7253,N_7226);
xor U8079 (N_8079,N_7020,N_7455);
nand U8080 (N_8080,N_6882,N_7182);
nor U8081 (N_8081,N_6888,N_7485);
xor U8082 (N_8082,N_7363,N_7019);
nand U8083 (N_8083,N_6825,N_7298);
or U8084 (N_8084,N_7428,N_7451);
or U8085 (N_8085,N_7250,N_6975);
and U8086 (N_8086,N_6797,N_6777);
or U8087 (N_8087,N_7322,N_7438);
or U8088 (N_8088,N_7441,N_7366);
and U8089 (N_8089,N_7025,N_6826);
xor U8090 (N_8090,N_6993,N_7241);
and U8091 (N_8091,N_6835,N_7273);
and U8092 (N_8092,N_7111,N_6942);
or U8093 (N_8093,N_7138,N_7091);
xor U8094 (N_8094,N_6879,N_7252);
nor U8095 (N_8095,N_6880,N_7183);
nand U8096 (N_8096,N_7339,N_7025);
xor U8097 (N_8097,N_7499,N_7260);
xor U8098 (N_8098,N_7389,N_7330);
nor U8099 (N_8099,N_7096,N_7116);
nand U8100 (N_8100,N_6827,N_6920);
nand U8101 (N_8101,N_7491,N_6899);
nand U8102 (N_8102,N_7494,N_6892);
nand U8103 (N_8103,N_7300,N_6766);
nand U8104 (N_8104,N_7442,N_7077);
nand U8105 (N_8105,N_7158,N_7311);
and U8106 (N_8106,N_7160,N_7419);
or U8107 (N_8107,N_7287,N_7363);
and U8108 (N_8108,N_7342,N_7220);
xnor U8109 (N_8109,N_6830,N_6998);
and U8110 (N_8110,N_7131,N_6984);
nor U8111 (N_8111,N_7235,N_6903);
xnor U8112 (N_8112,N_7292,N_7429);
xor U8113 (N_8113,N_7086,N_7206);
or U8114 (N_8114,N_7436,N_7213);
or U8115 (N_8115,N_7204,N_6940);
xnor U8116 (N_8116,N_6898,N_6792);
xnor U8117 (N_8117,N_7143,N_7140);
xnor U8118 (N_8118,N_7226,N_7365);
nor U8119 (N_8119,N_7385,N_7461);
nor U8120 (N_8120,N_7364,N_7092);
nand U8121 (N_8121,N_7115,N_7456);
nor U8122 (N_8122,N_7282,N_7259);
or U8123 (N_8123,N_7383,N_7199);
nand U8124 (N_8124,N_7027,N_6885);
nand U8125 (N_8125,N_7217,N_6947);
and U8126 (N_8126,N_7418,N_7432);
nor U8127 (N_8127,N_6768,N_6825);
nor U8128 (N_8128,N_7335,N_7483);
nand U8129 (N_8129,N_6980,N_7264);
nor U8130 (N_8130,N_7052,N_7218);
xnor U8131 (N_8131,N_6950,N_7109);
and U8132 (N_8132,N_6953,N_7476);
and U8133 (N_8133,N_7310,N_7089);
xor U8134 (N_8134,N_7053,N_7477);
nor U8135 (N_8135,N_7266,N_7309);
nand U8136 (N_8136,N_7433,N_6841);
nor U8137 (N_8137,N_7279,N_6940);
nand U8138 (N_8138,N_7296,N_6878);
nand U8139 (N_8139,N_7374,N_7084);
nor U8140 (N_8140,N_7189,N_6983);
or U8141 (N_8141,N_7204,N_7495);
xor U8142 (N_8142,N_7417,N_7286);
nor U8143 (N_8143,N_6894,N_7218);
xnor U8144 (N_8144,N_6769,N_6817);
and U8145 (N_8145,N_7031,N_7341);
nand U8146 (N_8146,N_7341,N_7114);
nor U8147 (N_8147,N_6930,N_7111);
nand U8148 (N_8148,N_7460,N_7091);
and U8149 (N_8149,N_7147,N_7458);
nor U8150 (N_8150,N_7330,N_6753);
nand U8151 (N_8151,N_7113,N_7352);
or U8152 (N_8152,N_7053,N_7315);
nand U8153 (N_8153,N_7489,N_7349);
xor U8154 (N_8154,N_7388,N_7477);
nand U8155 (N_8155,N_7322,N_6890);
nor U8156 (N_8156,N_6810,N_6896);
nor U8157 (N_8157,N_7467,N_7197);
and U8158 (N_8158,N_7114,N_7142);
nor U8159 (N_8159,N_7496,N_7354);
and U8160 (N_8160,N_7307,N_7389);
xnor U8161 (N_8161,N_7357,N_7206);
nand U8162 (N_8162,N_6971,N_7284);
xor U8163 (N_8163,N_6819,N_7092);
nand U8164 (N_8164,N_6932,N_6928);
nor U8165 (N_8165,N_7128,N_6850);
nor U8166 (N_8166,N_7063,N_7059);
nor U8167 (N_8167,N_6954,N_7261);
nor U8168 (N_8168,N_7410,N_7013);
nor U8169 (N_8169,N_7109,N_7176);
and U8170 (N_8170,N_7454,N_6804);
nand U8171 (N_8171,N_6989,N_7131);
nor U8172 (N_8172,N_7395,N_6938);
nor U8173 (N_8173,N_6855,N_7115);
nand U8174 (N_8174,N_7210,N_7284);
or U8175 (N_8175,N_7028,N_7337);
or U8176 (N_8176,N_6935,N_7397);
nor U8177 (N_8177,N_7146,N_7390);
nand U8178 (N_8178,N_7080,N_7083);
or U8179 (N_8179,N_7039,N_7240);
and U8180 (N_8180,N_6976,N_7440);
xnor U8181 (N_8181,N_6833,N_6831);
and U8182 (N_8182,N_7336,N_7135);
xor U8183 (N_8183,N_7334,N_6790);
nand U8184 (N_8184,N_7485,N_7256);
xnor U8185 (N_8185,N_6797,N_7166);
or U8186 (N_8186,N_7442,N_6904);
nand U8187 (N_8187,N_6760,N_6989);
nor U8188 (N_8188,N_6841,N_7457);
or U8189 (N_8189,N_7324,N_6857);
or U8190 (N_8190,N_7086,N_7154);
nor U8191 (N_8191,N_6817,N_7274);
nand U8192 (N_8192,N_7428,N_7098);
nand U8193 (N_8193,N_6752,N_6757);
nand U8194 (N_8194,N_7003,N_7431);
xnor U8195 (N_8195,N_7351,N_7207);
xor U8196 (N_8196,N_6772,N_7160);
xor U8197 (N_8197,N_7158,N_7119);
and U8198 (N_8198,N_6804,N_6948);
and U8199 (N_8199,N_6983,N_7464);
nand U8200 (N_8200,N_7412,N_6907);
nand U8201 (N_8201,N_7347,N_6977);
nor U8202 (N_8202,N_6790,N_6854);
nand U8203 (N_8203,N_7273,N_7287);
nand U8204 (N_8204,N_7402,N_6943);
and U8205 (N_8205,N_7422,N_7038);
nor U8206 (N_8206,N_7407,N_7169);
or U8207 (N_8207,N_6957,N_7086);
nand U8208 (N_8208,N_6981,N_6974);
nand U8209 (N_8209,N_7162,N_6758);
and U8210 (N_8210,N_7142,N_7471);
nor U8211 (N_8211,N_7281,N_6807);
xor U8212 (N_8212,N_7174,N_7479);
or U8213 (N_8213,N_7111,N_7457);
xor U8214 (N_8214,N_7081,N_6971);
nand U8215 (N_8215,N_6762,N_6761);
nand U8216 (N_8216,N_7498,N_6968);
and U8217 (N_8217,N_6969,N_6956);
nor U8218 (N_8218,N_7012,N_6751);
xor U8219 (N_8219,N_6915,N_7279);
xor U8220 (N_8220,N_7137,N_7363);
or U8221 (N_8221,N_7297,N_7134);
and U8222 (N_8222,N_7366,N_7141);
and U8223 (N_8223,N_6805,N_7371);
and U8224 (N_8224,N_7397,N_6801);
nand U8225 (N_8225,N_7498,N_7381);
or U8226 (N_8226,N_7051,N_7475);
or U8227 (N_8227,N_6827,N_6971);
or U8228 (N_8228,N_7144,N_7462);
nor U8229 (N_8229,N_7013,N_6838);
nor U8230 (N_8230,N_7400,N_6862);
and U8231 (N_8231,N_7336,N_7461);
or U8232 (N_8232,N_6872,N_7465);
and U8233 (N_8233,N_7444,N_6915);
or U8234 (N_8234,N_7083,N_7182);
nor U8235 (N_8235,N_6822,N_7118);
xor U8236 (N_8236,N_7326,N_7405);
nand U8237 (N_8237,N_7352,N_6968);
and U8238 (N_8238,N_7296,N_7259);
xor U8239 (N_8239,N_7174,N_7341);
xnor U8240 (N_8240,N_7122,N_7124);
nand U8241 (N_8241,N_7122,N_6919);
or U8242 (N_8242,N_7487,N_7410);
xor U8243 (N_8243,N_6865,N_7271);
nor U8244 (N_8244,N_6849,N_6956);
nor U8245 (N_8245,N_7027,N_6863);
nand U8246 (N_8246,N_6821,N_7371);
nor U8247 (N_8247,N_6766,N_6892);
or U8248 (N_8248,N_7000,N_6784);
nand U8249 (N_8249,N_6856,N_7262);
xor U8250 (N_8250,N_8221,N_8072);
nor U8251 (N_8251,N_7951,N_7700);
nor U8252 (N_8252,N_7737,N_7738);
xor U8253 (N_8253,N_8152,N_7808);
and U8254 (N_8254,N_7598,N_7705);
or U8255 (N_8255,N_7566,N_8076);
nand U8256 (N_8256,N_8048,N_8079);
and U8257 (N_8257,N_8228,N_7628);
nand U8258 (N_8258,N_7899,N_7665);
nand U8259 (N_8259,N_7658,N_7526);
nor U8260 (N_8260,N_7975,N_8239);
or U8261 (N_8261,N_8195,N_7950);
nand U8262 (N_8262,N_8174,N_7998);
and U8263 (N_8263,N_8211,N_7543);
or U8264 (N_8264,N_7720,N_8208);
nor U8265 (N_8265,N_7818,N_8102);
and U8266 (N_8266,N_7525,N_7617);
xnor U8267 (N_8267,N_8109,N_7519);
nand U8268 (N_8268,N_7907,N_7994);
and U8269 (N_8269,N_7866,N_7666);
nand U8270 (N_8270,N_8094,N_7645);
xnor U8271 (N_8271,N_7925,N_7743);
xnor U8272 (N_8272,N_7933,N_7817);
nand U8273 (N_8273,N_7623,N_8248);
nand U8274 (N_8274,N_8240,N_7547);
nor U8275 (N_8275,N_7684,N_7978);
nor U8276 (N_8276,N_7501,N_8210);
and U8277 (N_8277,N_7806,N_7513);
xor U8278 (N_8278,N_7770,N_7548);
or U8279 (N_8279,N_7740,N_7870);
or U8280 (N_8280,N_7964,N_7886);
or U8281 (N_8281,N_7857,N_7853);
nand U8282 (N_8282,N_7932,N_8212);
nor U8283 (N_8283,N_7568,N_7643);
xor U8284 (N_8284,N_8047,N_8086);
nor U8285 (N_8285,N_8145,N_7747);
and U8286 (N_8286,N_8184,N_8038);
xnor U8287 (N_8287,N_7930,N_7939);
or U8288 (N_8288,N_7997,N_7592);
and U8289 (N_8289,N_7799,N_7839);
or U8290 (N_8290,N_7947,N_7502);
xnor U8291 (N_8291,N_8179,N_7772);
and U8292 (N_8292,N_7967,N_7744);
nand U8293 (N_8293,N_7938,N_7545);
nor U8294 (N_8294,N_7791,N_8181);
or U8295 (N_8295,N_8198,N_7797);
nand U8296 (N_8296,N_7745,N_7830);
nor U8297 (N_8297,N_7825,N_8139);
nor U8298 (N_8298,N_7692,N_7773);
nor U8299 (N_8299,N_7953,N_7582);
nor U8300 (N_8300,N_8200,N_8036);
and U8301 (N_8301,N_8037,N_7775);
nor U8302 (N_8302,N_7713,N_7602);
nor U8303 (N_8303,N_7794,N_7832);
or U8304 (N_8304,N_7533,N_8144);
and U8305 (N_8305,N_8103,N_8024);
xor U8306 (N_8306,N_8026,N_8077);
nand U8307 (N_8307,N_7649,N_7538);
nand U8308 (N_8308,N_7663,N_7911);
nor U8309 (N_8309,N_8030,N_8029);
and U8310 (N_8310,N_7673,N_8162);
xnor U8311 (N_8311,N_7650,N_7826);
nand U8312 (N_8312,N_7683,N_7622);
and U8313 (N_8313,N_8117,N_7725);
nor U8314 (N_8314,N_7562,N_7708);
xor U8315 (N_8315,N_7636,N_7807);
nand U8316 (N_8316,N_8163,N_7721);
xnor U8317 (N_8317,N_7942,N_7996);
nor U8318 (N_8318,N_7715,N_7779);
nand U8319 (N_8319,N_8236,N_7621);
and U8320 (N_8320,N_7914,N_8180);
nand U8321 (N_8321,N_7771,N_7668);
and U8322 (N_8322,N_7632,N_7667);
xor U8323 (N_8323,N_8055,N_7517);
and U8324 (N_8324,N_8101,N_8022);
and U8325 (N_8325,N_7641,N_7879);
and U8326 (N_8326,N_7966,N_7719);
and U8327 (N_8327,N_7736,N_7676);
nor U8328 (N_8328,N_7889,N_7885);
nand U8329 (N_8329,N_7924,N_7686);
nand U8330 (N_8330,N_7813,N_7837);
or U8331 (N_8331,N_8078,N_7928);
nor U8332 (N_8332,N_7861,N_7755);
and U8333 (N_8333,N_8087,N_7822);
and U8334 (N_8334,N_7695,N_8110);
and U8335 (N_8335,N_7634,N_7840);
nor U8336 (N_8336,N_8104,N_7710);
or U8337 (N_8337,N_7844,N_8189);
or U8338 (N_8338,N_7601,N_7988);
or U8339 (N_8339,N_7546,N_8057);
or U8340 (N_8340,N_8105,N_7577);
nor U8341 (N_8341,N_7786,N_7821);
xnor U8342 (N_8342,N_8068,N_7528);
or U8343 (N_8343,N_8246,N_8081);
xnor U8344 (N_8344,N_8066,N_7619);
xor U8345 (N_8345,N_7846,N_8091);
nor U8346 (N_8346,N_8218,N_8112);
nor U8347 (N_8347,N_7594,N_8199);
xnor U8348 (N_8348,N_7597,N_7854);
nand U8349 (N_8349,N_8075,N_7532);
or U8350 (N_8350,N_8201,N_7927);
nor U8351 (N_8351,N_8217,N_7958);
and U8352 (N_8352,N_8203,N_7915);
xnor U8353 (N_8353,N_8143,N_8222);
nor U8354 (N_8354,N_8099,N_7903);
and U8355 (N_8355,N_8182,N_8187);
and U8356 (N_8356,N_8125,N_8205);
nor U8357 (N_8357,N_7882,N_7963);
nor U8358 (N_8358,N_8209,N_7523);
nor U8359 (N_8359,N_7691,N_7812);
xor U8360 (N_8360,N_7760,N_8107);
and U8361 (N_8361,N_7909,N_8185);
nor U8362 (N_8362,N_8193,N_7509);
or U8363 (N_8363,N_7678,N_8007);
or U8364 (N_8364,N_7892,N_7787);
and U8365 (N_8365,N_7674,N_8067);
nor U8366 (N_8366,N_7888,N_7557);
xor U8367 (N_8367,N_8041,N_7985);
nand U8368 (N_8368,N_8229,N_7919);
xnor U8369 (N_8369,N_7835,N_7754);
nand U8370 (N_8370,N_7904,N_8090);
nand U8371 (N_8371,N_8120,N_7626);
xor U8372 (N_8372,N_7810,N_8188);
xnor U8373 (N_8373,N_7588,N_8062);
nand U8374 (N_8374,N_7918,N_8158);
xnor U8375 (N_8375,N_8082,N_7615);
nand U8376 (N_8376,N_7661,N_7908);
or U8377 (N_8377,N_8031,N_7876);
nor U8378 (N_8378,N_7605,N_7877);
xnor U8379 (N_8379,N_7793,N_8225);
and U8380 (N_8380,N_8159,N_8045);
nor U8381 (N_8381,N_7635,N_8175);
or U8382 (N_8382,N_7989,N_7644);
nand U8383 (N_8383,N_7596,N_7504);
xor U8384 (N_8384,N_8033,N_7934);
or U8385 (N_8385,N_7534,N_8183);
nor U8386 (N_8386,N_8194,N_7974);
nand U8387 (N_8387,N_7627,N_8249);
xor U8388 (N_8388,N_7630,N_7757);
nand U8389 (N_8389,N_7677,N_8234);
or U8390 (N_8390,N_7707,N_7767);
nand U8391 (N_8391,N_7979,N_8237);
nand U8392 (N_8392,N_8227,N_8032);
nand U8393 (N_8393,N_8059,N_7874);
xor U8394 (N_8394,N_7777,N_8088);
nor U8395 (N_8395,N_7539,N_7809);
and U8396 (N_8396,N_7884,N_7961);
nor U8397 (N_8397,N_7573,N_7941);
and U8398 (N_8398,N_7579,N_7672);
and U8399 (N_8399,N_7873,N_8186);
and U8400 (N_8400,N_8017,N_7995);
xor U8401 (N_8401,N_7800,N_8085);
or U8402 (N_8402,N_7954,N_7609);
xnor U8403 (N_8403,N_7593,N_7552);
xor U8404 (N_8404,N_7508,N_7860);
or U8405 (N_8405,N_7560,N_7926);
nand U8406 (N_8406,N_7828,N_8010);
or U8407 (N_8407,N_7976,N_8111);
or U8408 (N_8408,N_7701,N_7993);
nand U8409 (N_8409,N_7906,N_7783);
and U8410 (N_8410,N_7983,N_7990);
nor U8411 (N_8411,N_8106,N_7699);
and U8412 (N_8412,N_8113,N_8160);
nand U8413 (N_8413,N_7781,N_7893);
nor U8414 (N_8414,N_7518,N_7780);
xnor U8415 (N_8415,N_8133,N_8027);
and U8416 (N_8416,N_8054,N_7910);
or U8417 (N_8417,N_8148,N_7524);
and U8418 (N_8418,N_7848,N_8006);
nand U8419 (N_8419,N_8053,N_7732);
and U8420 (N_8420,N_7669,N_7803);
and U8421 (N_8421,N_8164,N_7751);
nor U8422 (N_8422,N_7714,N_8245);
nand U8423 (N_8423,N_7585,N_7805);
or U8424 (N_8424,N_7625,N_8231);
nor U8425 (N_8425,N_7992,N_7559);
and U8426 (N_8426,N_7694,N_7633);
xor U8427 (N_8427,N_7776,N_7811);
or U8428 (N_8428,N_7646,N_7733);
and U8429 (N_8429,N_7916,N_7880);
xor U8430 (N_8430,N_7782,N_7764);
and U8431 (N_8431,N_8130,N_8084);
nor U8432 (N_8432,N_7977,N_8238);
nand U8433 (N_8433,N_7662,N_7937);
nor U8434 (N_8434,N_7824,N_7789);
nand U8435 (N_8435,N_7685,N_7550);
nand U8436 (N_8436,N_7836,N_8170);
or U8437 (N_8437,N_7956,N_7957);
xnor U8438 (N_8438,N_7792,N_7746);
xor U8439 (N_8439,N_7614,N_7640);
or U8440 (N_8440,N_7895,N_8008);
and U8441 (N_8441,N_7570,N_7618);
nor U8442 (N_8442,N_7554,N_7887);
nand U8443 (N_8443,N_8242,N_7819);
nor U8444 (N_8444,N_7687,N_7834);
xnor U8445 (N_8445,N_8005,N_7717);
nand U8446 (N_8446,N_7693,N_8177);
nor U8447 (N_8447,N_7600,N_8049);
xnor U8448 (N_8448,N_8216,N_7960);
nor U8449 (N_8449,N_8131,N_7535);
nand U8450 (N_8450,N_8050,N_7574);
and U8451 (N_8451,N_7761,N_8043);
or U8452 (N_8452,N_8235,N_8165);
xor U8453 (N_8453,N_7541,N_7704);
nor U8454 (N_8454,N_8020,N_7587);
nor U8455 (N_8455,N_7702,N_8243);
xnor U8456 (N_8456,N_7580,N_7897);
nand U8457 (N_8457,N_7553,N_8069);
nor U8458 (N_8458,N_7682,N_7766);
nand U8459 (N_8459,N_8040,N_8074);
and U8460 (N_8460,N_8171,N_7616);
nand U8461 (N_8461,N_8042,N_7748);
xnor U8462 (N_8462,N_7894,N_7675);
and U8463 (N_8463,N_7639,N_7867);
and U8464 (N_8464,N_7599,N_7816);
nor U8465 (N_8465,N_7968,N_7851);
or U8466 (N_8466,N_7689,N_7631);
nor U8467 (N_8467,N_7542,N_8003);
xnor U8468 (N_8468,N_7608,N_7982);
xor U8469 (N_8469,N_7657,N_8015);
xor U8470 (N_8470,N_8060,N_7734);
and U8471 (N_8471,N_8147,N_7679);
nand U8472 (N_8472,N_7530,N_8115);
or U8473 (N_8473,N_7750,N_7804);
nor U8474 (N_8474,N_7891,N_7921);
nor U8475 (N_8475,N_7863,N_8202);
xor U8476 (N_8476,N_7936,N_7831);
or U8477 (N_8477,N_7759,N_8039);
or U8478 (N_8478,N_8097,N_7698);
nor U8479 (N_8479,N_7505,N_7955);
or U8480 (N_8480,N_7847,N_7820);
or U8481 (N_8481,N_7741,N_7637);
nand U8482 (N_8482,N_8192,N_7913);
nand U8483 (N_8483,N_7709,N_8044);
and U8484 (N_8484,N_7900,N_7540);
nor U8485 (N_8485,N_7872,N_7516);
nand U8486 (N_8486,N_7984,N_7859);
and U8487 (N_8487,N_8219,N_7972);
nand U8488 (N_8488,N_7629,N_7986);
nor U8489 (N_8489,N_7688,N_7731);
xnor U8490 (N_8490,N_7729,N_7522);
xor U8491 (N_8491,N_7917,N_8134);
nor U8492 (N_8492,N_8197,N_8046);
or U8493 (N_8493,N_7712,N_7778);
xor U8494 (N_8494,N_8070,N_8034);
xnor U8495 (N_8495,N_8220,N_7935);
nand U8496 (N_8496,N_7620,N_7814);
xor U8497 (N_8497,N_7556,N_8206);
nor U8498 (N_8498,N_7711,N_7584);
nand U8499 (N_8499,N_8065,N_7656);
xor U8500 (N_8500,N_7946,N_8244);
xor U8501 (N_8501,N_8114,N_7537);
or U8502 (N_8502,N_7652,N_7671);
and U8503 (N_8503,N_8178,N_8025);
nor U8504 (N_8504,N_8014,N_7659);
xnor U8505 (N_8505,N_8051,N_7503);
or U8506 (N_8506,N_7841,N_8156);
nand U8507 (N_8507,N_8129,N_7795);
or U8508 (N_8508,N_8128,N_8064);
or U8509 (N_8509,N_7544,N_8141);
nor U8510 (N_8510,N_8126,N_7681);
xnor U8511 (N_8511,N_7581,N_7823);
nand U8512 (N_8512,N_7739,N_8142);
nor U8513 (N_8513,N_8123,N_8155);
or U8514 (N_8514,N_8119,N_8035);
nor U8515 (N_8515,N_7647,N_7576);
nor U8516 (N_8516,N_7965,N_7752);
and U8517 (N_8517,N_8149,N_8098);
and U8518 (N_8518,N_7833,N_7604);
nand U8519 (N_8519,N_7788,N_8093);
xnor U8520 (N_8520,N_7849,N_8019);
and U8521 (N_8521,N_7558,N_7890);
nand U8522 (N_8522,N_7871,N_8167);
nor U8523 (N_8523,N_7653,N_7651);
nor U8524 (N_8524,N_8154,N_7607);
nor U8525 (N_8525,N_7586,N_7536);
and U8526 (N_8526,N_7549,N_7730);
xor U8527 (N_8527,N_7664,N_7970);
nand U8528 (N_8528,N_7922,N_8232);
and U8529 (N_8529,N_7727,N_8071);
or U8530 (N_8530,N_8204,N_7912);
xor U8531 (N_8531,N_7507,N_7852);
nand U8532 (N_8532,N_8021,N_8223);
xor U8533 (N_8533,N_7697,N_8230);
or U8534 (N_8534,N_7753,N_7829);
and U8535 (N_8535,N_7572,N_8132);
nor U8536 (N_8536,N_7898,N_8095);
nor U8537 (N_8537,N_7878,N_7929);
or U8538 (N_8538,N_7510,N_7856);
nand U8539 (N_8539,N_7749,N_7722);
nor U8540 (N_8540,N_7902,N_7583);
and U8541 (N_8541,N_7578,N_8100);
or U8542 (N_8542,N_7931,N_7512);
nand U8543 (N_8543,N_8168,N_7991);
and U8544 (N_8544,N_7500,N_7703);
xor U8545 (N_8545,N_7940,N_8214);
nand U8546 (N_8546,N_7802,N_8004);
and U8547 (N_8547,N_8196,N_7726);
or U8548 (N_8548,N_7855,N_7716);
nand U8549 (N_8549,N_7680,N_7648);
xnor U8550 (N_8550,N_7762,N_7881);
or U8551 (N_8551,N_7696,N_7529);
or U8552 (N_8552,N_8176,N_7969);
nor U8553 (N_8553,N_8224,N_8011);
or U8554 (N_8554,N_8092,N_8080);
nor U8555 (N_8555,N_7724,N_8016);
xnor U8556 (N_8556,N_7949,N_8052);
xnor U8557 (N_8557,N_7563,N_8013);
and U8558 (N_8558,N_7742,N_8135);
or U8559 (N_8559,N_7591,N_7948);
nand U8560 (N_8560,N_7561,N_8207);
and U8561 (N_8561,N_8108,N_8213);
xnor U8562 (N_8562,N_8173,N_7862);
nor U8563 (N_8563,N_7511,N_8058);
nor U8564 (N_8564,N_8012,N_7531);
and U8565 (N_8565,N_7521,N_8233);
and U8566 (N_8566,N_8140,N_8215);
or U8567 (N_8567,N_7624,N_7527);
xor U8568 (N_8568,N_7515,N_7506);
and U8569 (N_8569,N_7723,N_8001);
or U8570 (N_8570,N_7551,N_8190);
and U8571 (N_8571,N_8096,N_7590);
nor U8572 (N_8572,N_8118,N_7981);
and U8573 (N_8573,N_8002,N_7864);
and U8574 (N_8574,N_7896,N_8137);
xor U8575 (N_8575,N_7611,N_7959);
nand U8576 (N_8576,N_7868,N_7758);
nand U8577 (N_8577,N_7850,N_8161);
and U8578 (N_8578,N_7613,N_7514);
or U8579 (N_8579,N_7905,N_7763);
nand U8580 (N_8580,N_7845,N_7706);
or U8581 (N_8581,N_7796,N_7571);
or U8582 (N_8582,N_7655,N_8146);
xnor U8583 (N_8583,N_8138,N_8127);
and U8584 (N_8584,N_7567,N_7944);
and U8585 (N_8585,N_7569,N_8150);
nand U8586 (N_8586,N_7923,N_8191);
or U8587 (N_8587,N_8172,N_7565);
nor U8588 (N_8588,N_8023,N_8166);
or U8589 (N_8589,N_7612,N_8157);
xor U8590 (N_8590,N_7827,N_7575);
xnor U8591 (N_8591,N_7564,N_8151);
xnor U8592 (N_8592,N_8083,N_7842);
nand U8593 (N_8593,N_7603,N_7815);
nor U8594 (N_8594,N_7869,N_7801);
and U8595 (N_8595,N_7875,N_8226);
nand U8596 (N_8596,N_8009,N_8136);
and U8597 (N_8597,N_8028,N_7718);
xnor U8598 (N_8598,N_8169,N_8116);
nor U8599 (N_8599,N_8247,N_7901);
or U8600 (N_8600,N_7999,N_8089);
xnor U8601 (N_8601,N_7769,N_7555);
or U8602 (N_8602,N_7843,N_7971);
or U8603 (N_8603,N_8241,N_7735);
nor U8604 (N_8604,N_7728,N_7654);
xor U8605 (N_8605,N_7943,N_8124);
xnor U8606 (N_8606,N_7765,N_7790);
and U8607 (N_8607,N_8063,N_7920);
xnor U8608 (N_8608,N_7589,N_7690);
nand U8609 (N_8609,N_7973,N_8073);
nor U8610 (N_8610,N_7595,N_7768);
xnor U8611 (N_8611,N_7660,N_8122);
nor U8612 (N_8612,N_7606,N_8056);
xnor U8613 (N_8613,N_7785,N_7642);
xnor U8614 (N_8614,N_8121,N_7798);
nor U8615 (N_8615,N_7838,N_7962);
xor U8616 (N_8616,N_7865,N_7952);
xnor U8617 (N_8617,N_7987,N_7638);
and U8618 (N_8618,N_7883,N_7784);
nand U8619 (N_8619,N_8018,N_7945);
nand U8620 (N_8620,N_7858,N_7610);
and U8621 (N_8621,N_7756,N_8000);
or U8622 (N_8622,N_7520,N_7980);
and U8623 (N_8623,N_8061,N_8153);
xor U8624 (N_8624,N_7774,N_7670);
xor U8625 (N_8625,N_7692,N_8051);
and U8626 (N_8626,N_8211,N_7588);
xnor U8627 (N_8627,N_8024,N_7846);
or U8628 (N_8628,N_7796,N_7833);
or U8629 (N_8629,N_7541,N_8025);
nor U8630 (N_8630,N_7810,N_7775);
and U8631 (N_8631,N_8201,N_7614);
xnor U8632 (N_8632,N_7672,N_7607);
or U8633 (N_8633,N_8099,N_7537);
xnor U8634 (N_8634,N_8105,N_7863);
and U8635 (N_8635,N_7838,N_7688);
and U8636 (N_8636,N_7708,N_8105);
xnor U8637 (N_8637,N_7792,N_8050);
nand U8638 (N_8638,N_7931,N_7816);
or U8639 (N_8639,N_8063,N_7566);
xnor U8640 (N_8640,N_7851,N_7921);
nand U8641 (N_8641,N_7936,N_7777);
xor U8642 (N_8642,N_7960,N_8000);
nand U8643 (N_8643,N_7761,N_7766);
and U8644 (N_8644,N_7899,N_8241);
and U8645 (N_8645,N_7648,N_7720);
xor U8646 (N_8646,N_7518,N_8002);
nand U8647 (N_8647,N_7703,N_7918);
nor U8648 (N_8648,N_7588,N_7633);
and U8649 (N_8649,N_7593,N_8014);
or U8650 (N_8650,N_7538,N_7775);
or U8651 (N_8651,N_8245,N_7517);
xnor U8652 (N_8652,N_7826,N_8195);
nor U8653 (N_8653,N_8209,N_7656);
nor U8654 (N_8654,N_7899,N_7661);
nand U8655 (N_8655,N_7526,N_7521);
or U8656 (N_8656,N_7578,N_7594);
or U8657 (N_8657,N_7855,N_7863);
nor U8658 (N_8658,N_8076,N_7758);
nand U8659 (N_8659,N_7630,N_7946);
and U8660 (N_8660,N_7979,N_8143);
and U8661 (N_8661,N_8174,N_7818);
xnor U8662 (N_8662,N_7690,N_7772);
nor U8663 (N_8663,N_7600,N_8053);
nand U8664 (N_8664,N_7866,N_7611);
nor U8665 (N_8665,N_7815,N_8174);
nand U8666 (N_8666,N_7570,N_8223);
and U8667 (N_8667,N_7937,N_7988);
and U8668 (N_8668,N_7678,N_7642);
or U8669 (N_8669,N_7802,N_7591);
xor U8670 (N_8670,N_7931,N_8224);
nor U8671 (N_8671,N_7939,N_7991);
and U8672 (N_8672,N_7897,N_7574);
or U8673 (N_8673,N_7909,N_8159);
nand U8674 (N_8674,N_8157,N_7709);
nor U8675 (N_8675,N_7807,N_7919);
nand U8676 (N_8676,N_7675,N_7561);
nor U8677 (N_8677,N_7765,N_7999);
xor U8678 (N_8678,N_8056,N_7501);
nand U8679 (N_8679,N_8078,N_8185);
and U8680 (N_8680,N_7839,N_8206);
xnor U8681 (N_8681,N_8074,N_7969);
and U8682 (N_8682,N_7615,N_7640);
nand U8683 (N_8683,N_7520,N_7585);
and U8684 (N_8684,N_7874,N_7977);
or U8685 (N_8685,N_7943,N_8170);
or U8686 (N_8686,N_8051,N_8200);
nor U8687 (N_8687,N_7683,N_7810);
nand U8688 (N_8688,N_7943,N_7879);
or U8689 (N_8689,N_7867,N_7654);
nor U8690 (N_8690,N_7983,N_7514);
nor U8691 (N_8691,N_7938,N_7630);
xor U8692 (N_8692,N_7958,N_8190);
and U8693 (N_8693,N_8116,N_7849);
and U8694 (N_8694,N_7798,N_8066);
nand U8695 (N_8695,N_8090,N_7854);
xor U8696 (N_8696,N_7783,N_8099);
nor U8697 (N_8697,N_7951,N_7796);
nand U8698 (N_8698,N_7986,N_8103);
nor U8699 (N_8699,N_8106,N_8239);
nor U8700 (N_8700,N_7713,N_8197);
or U8701 (N_8701,N_7877,N_7622);
nor U8702 (N_8702,N_8077,N_7836);
nand U8703 (N_8703,N_7677,N_7648);
xnor U8704 (N_8704,N_7964,N_8093);
nand U8705 (N_8705,N_8202,N_7913);
nor U8706 (N_8706,N_7847,N_8229);
xor U8707 (N_8707,N_7977,N_7765);
nand U8708 (N_8708,N_8218,N_7580);
nor U8709 (N_8709,N_7641,N_7843);
nor U8710 (N_8710,N_8043,N_7628);
xor U8711 (N_8711,N_7740,N_7741);
or U8712 (N_8712,N_7873,N_8034);
xor U8713 (N_8713,N_7830,N_7906);
and U8714 (N_8714,N_8126,N_7628);
xnor U8715 (N_8715,N_7787,N_7652);
nor U8716 (N_8716,N_7783,N_8206);
nor U8717 (N_8717,N_7635,N_7779);
and U8718 (N_8718,N_7897,N_8082);
xnor U8719 (N_8719,N_7838,N_8091);
nand U8720 (N_8720,N_7962,N_7809);
and U8721 (N_8721,N_8176,N_8112);
xor U8722 (N_8722,N_8182,N_7647);
and U8723 (N_8723,N_7635,N_8070);
and U8724 (N_8724,N_8130,N_8033);
nand U8725 (N_8725,N_7633,N_7792);
and U8726 (N_8726,N_8183,N_7574);
and U8727 (N_8727,N_7695,N_7810);
and U8728 (N_8728,N_8184,N_8185);
or U8729 (N_8729,N_7943,N_8191);
and U8730 (N_8730,N_8152,N_7815);
nand U8731 (N_8731,N_7562,N_8114);
and U8732 (N_8732,N_7627,N_7749);
or U8733 (N_8733,N_8242,N_7696);
nand U8734 (N_8734,N_7501,N_8090);
nor U8735 (N_8735,N_8156,N_7575);
or U8736 (N_8736,N_8209,N_8002);
or U8737 (N_8737,N_7582,N_8154);
nand U8738 (N_8738,N_8012,N_7546);
xor U8739 (N_8739,N_7973,N_8162);
nand U8740 (N_8740,N_7896,N_7935);
and U8741 (N_8741,N_7875,N_7979);
or U8742 (N_8742,N_7939,N_7801);
xor U8743 (N_8743,N_8236,N_8057);
and U8744 (N_8744,N_8143,N_8180);
nor U8745 (N_8745,N_7933,N_7502);
or U8746 (N_8746,N_7833,N_7648);
xor U8747 (N_8747,N_7724,N_7864);
and U8748 (N_8748,N_7800,N_7557);
and U8749 (N_8749,N_8128,N_7892);
nor U8750 (N_8750,N_8227,N_8097);
nor U8751 (N_8751,N_7926,N_7572);
xnor U8752 (N_8752,N_7760,N_7666);
nand U8753 (N_8753,N_7978,N_7969);
and U8754 (N_8754,N_8137,N_7876);
nor U8755 (N_8755,N_7999,N_7694);
nand U8756 (N_8756,N_7625,N_7674);
xnor U8757 (N_8757,N_8023,N_7520);
nor U8758 (N_8758,N_7870,N_7729);
nand U8759 (N_8759,N_7780,N_7935);
nor U8760 (N_8760,N_7906,N_8103);
xor U8761 (N_8761,N_7900,N_7706);
nand U8762 (N_8762,N_7554,N_8057);
or U8763 (N_8763,N_7892,N_7933);
and U8764 (N_8764,N_8155,N_8235);
or U8765 (N_8765,N_7800,N_7631);
xor U8766 (N_8766,N_7631,N_7878);
nor U8767 (N_8767,N_8068,N_7749);
nor U8768 (N_8768,N_7966,N_7994);
or U8769 (N_8769,N_7752,N_7667);
or U8770 (N_8770,N_8015,N_7553);
or U8771 (N_8771,N_7891,N_7590);
xor U8772 (N_8772,N_7672,N_8018);
and U8773 (N_8773,N_8033,N_7890);
and U8774 (N_8774,N_7548,N_8038);
nor U8775 (N_8775,N_7911,N_8085);
or U8776 (N_8776,N_7790,N_7899);
xor U8777 (N_8777,N_7965,N_7764);
and U8778 (N_8778,N_7618,N_7881);
or U8779 (N_8779,N_8038,N_8138);
nand U8780 (N_8780,N_7742,N_7984);
nand U8781 (N_8781,N_8155,N_8107);
xor U8782 (N_8782,N_8135,N_7694);
and U8783 (N_8783,N_7749,N_7977);
nand U8784 (N_8784,N_7620,N_8012);
nand U8785 (N_8785,N_8001,N_7735);
xnor U8786 (N_8786,N_7875,N_7789);
nand U8787 (N_8787,N_7874,N_7984);
nor U8788 (N_8788,N_7775,N_8057);
and U8789 (N_8789,N_7684,N_7883);
nor U8790 (N_8790,N_8072,N_8093);
and U8791 (N_8791,N_7714,N_7890);
nor U8792 (N_8792,N_7798,N_7972);
and U8793 (N_8793,N_7750,N_7876);
and U8794 (N_8794,N_8046,N_8062);
nand U8795 (N_8795,N_7613,N_7972);
xor U8796 (N_8796,N_7948,N_7851);
or U8797 (N_8797,N_7728,N_7714);
nor U8798 (N_8798,N_8084,N_7611);
nand U8799 (N_8799,N_8239,N_7865);
nand U8800 (N_8800,N_7780,N_7870);
nand U8801 (N_8801,N_7721,N_8220);
and U8802 (N_8802,N_7989,N_7666);
and U8803 (N_8803,N_7808,N_7650);
or U8804 (N_8804,N_7586,N_7545);
nand U8805 (N_8805,N_8110,N_7966);
xnor U8806 (N_8806,N_7728,N_8015);
xor U8807 (N_8807,N_8224,N_8026);
or U8808 (N_8808,N_7677,N_7837);
or U8809 (N_8809,N_8214,N_7894);
nand U8810 (N_8810,N_7563,N_8239);
nand U8811 (N_8811,N_7949,N_7538);
and U8812 (N_8812,N_8187,N_7777);
xnor U8813 (N_8813,N_8184,N_8112);
and U8814 (N_8814,N_8186,N_8203);
nand U8815 (N_8815,N_7758,N_8175);
xnor U8816 (N_8816,N_7797,N_7917);
nand U8817 (N_8817,N_8017,N_7881);
and U8818 (N_8818,N_7896,N_7629);
and U8819 (N_8819,N_8169,N_7532);
nand U8820 (N_8820,N_7763,N_8226);
nand U8821 (N_8821,N_7644,N_8049);
nor U8822 (N_8822,N_7671,N_8022);
nand U8823 (N_8823,N_7965,N_7712);
or U8824 (N_8824,N_7854,N_7898);
and U8825 (N_8825,N_8188,N_7943);
or U8826 (N_8826,N_8057,N_7561);
and U8827 (N_8827,N_7517,N_8092);
nor U8828 (N_8828,N_8238,N_8004);
xor U8829 (N_8829,N_7893,N_7796);
xor U8830 (N_8830,N_7696,N_7820);
xor U8831 (N_8831,N_7757,N_7992);
xor U8832 (N_8832,N_7577,N_8154);
and U8833 (N_8833,N_8042,N_7652);
or U8834 (N_8834,N_7903,N_7553);
nor U8835 (N_8835,N_7538,N_7628);
or U8836 (N_8836,N_7837,N_7622);
and U8837 (N_8837,N_7780,N_8072);
and U8838 (N_8838,N_7692,N_8026);
nand U8839 (N_8839,N_7829,N_8043);
and U8840 (N_8840,N_7567,N_8230);
or U8841 (N_8841,N_8019,N_8030);
nor U8842 (N_8842,N_7918,N_8106);
nor U8843 (N_8843,N_7692,N_7927);
and U8844 (N_8844,N_7843,N_7584);
xnor U8845 (N_8845,N_7971,N_7582);
nor U8846 (N_8846,N_7655,N_8228);
nand U8847 (N_8847,N_8239,N_7817);
xnor U8848 (N_8848,N_7645,N_7704);
or U8849 (N_8849,N_8246,N_7816);
xnor U8850 (N_8850,N_8160,N_7861);
or U8851 (N_8851,N_8235,N_8214);
nor U8852 (N_8852,N_7832,N_7788);
xor U8853 (N_8853,N_7775,N_7945);
xor U8854 (N_8854,N_7910,N_8079);
nor U8855 (N_8855,N_8135,N_7862);
or U8856 (N_8856,N_7696,N_7606);
nor U8857 (N_8857,N_7692,N_8204);
nand U8858 (N_8858,N_8047,N_7529);
xor U8859 (N_8859,N_7720,N_8017);
xnor U8860 (N_8860,N_7570,N_7588);
and U8861 (N_8861,N_7939,N_8064);
or U8862 (N_8862,N_7787,N_8210);
and U8863 (N_8863,N_7516,N_8031);
nor U8864 (N_8864,N_7903,N_7771);
or U8865 (N_8865,N_7791,N_7865);
xnor U8866 (N_8866,N_7575,N_8111);
xnor U8867 (N_8867,N_7626,N_7613);
xor U8868 (N_8868,N_8226,N_7701);
xor U8869 (N_8869,N_7813,N_8019);
xnor U8870 (N_8870,N_7804,N_7595);
nor U8871 (N_8871,N_7585,N_7897);
nor U8872 (N_8872,N_8064,N_8198);
nand U8873 (N_8873,N_8168,N_7647);
and U8874 (N_8874,N_7833,N_8107);
nor U8875 (N_8875,N_7988,N_8051);
or U8876 (N_8876,N_8137,N_8120);
xnor U8877 (N_8877,N_7901,N_7617);
or U8878 (N_8878,N_7517,N_7642);
nor U8879 (N_8879,N_7615,N_8148);
nor U8880 (N_8880,N_7835,N_8177);
or U8881 (N_8881,N_7699,N_8175);
nor U8882 (N_8882,N_7608,N_7713);
and U8883 (N_8883,N_8134,N_7895);
or U8884 (N_8884,N_8129,N_7791);
nor U8885 (N_8885,N_7642,N_8011);
nand U8886 (N_8886,N_7652,N_7582);
nand U8887 (N_8887,N_7655,N_8066);
nand U8888 (N_8888,N_7998,N_8016);
nor U8889 (N_8889,N_7997,N_8200);
and U8890 (N_8890,N_7595,N_7927);
xor U8891 (N_8891,N_7657,N_8165);
and U8892 (N_8892,N_7704,N_7683);
nand U8893 (N_8893,N_8000,N_7942);
nor U8894 (N_8894,N_7745,N_7870);
or U8895 (N_8895,N_7553,N_8172);
or U8896 (N_8896,N_7824,N_8095);
and U8897 (N_8897,N_7719,N_8212);
nor U8898 (N_8898,N_8142,N_8048);
nand U8899 (N_8899,N_7865,N_7870);
nand U8900 (N_8900,N_8102,N_7803);
xor U8901 (N_8901,N_7801,N_7679);
nor U8902 (N_8902,N_7822,N_8173);
nor U8903 (N_8903,N_8087,N_7849);
xnor U8904 (N_8904,N_8136,N_7542);
nand U8905 (N_8905,N_7601,N_8035);
or U8906 (N_8906,N_8181,N_7980);
nand U8907 (N_8907,N_8244,N_7897);
or U8908 (N_8908,N_7892,N_7539);
or U8909 (N_8909,N_8198,N_7901);
or U8910 (N_8910,N_7761,N_8113);
nor U8911 (N_8911,N_7571,N_7533);
or U8912 (N_8912,N_7656,N_8174);
nand U8913 (N_8913,N_7581,N_8238);
nand U8914 (N_8914,N_7978,N_7754);
nor U8915 (N_8915,N_7677,N_8068);
or U8916 (N_8916,N_7788,N_7605);
or U8917 (N_8917,N_7581,N_7623);
xor U8918 (N_8918,N_7699,N_8030);
xnor U8919 (N_8919,N_7840,N_7606);
or U8920 (N_8920,N_7886,N_7803);
or U8921 (N_8921,N_7744,N_7881);
or U8922 (N_8922,N_8073,N_7549);
xor U8923 (N_8923,N_8070,N_8060);
xor U8924 (N_8924,N_8142,N_7679);
nor U8925 (N_8925,N_7837,N_7568);
and U8926 (N_8926,N_8103,N_7728);
and U8927 (N_8927,N_7951,N_8230);
or U8928 (N_8928,N_7796,N_8239);
nand U8929 (N_8929,N_7889,N_8042);
nor U8930 (N_8930,N_7771,N_7954);
nor U8931 (N_8931,N_8155,N_7798);
nand U8932 (N_8932,N_7762,N_8188);
nand U8933 (N_8933,N_7991,N_7914);
nand U8934 (N_8934,N_7845,N_8216);
nor U8935 (N_8935,N_7551,N_7935);
or U8936 (N_8936,N_8051,N_7881);
xor U8937 (N_8937,N_8232,N_7634);
or U8938 (N_8938,N_8165,N_7908);
or U8939 (N_8939,N_7957,N_7658);
or U8940 (N_8940,N_7672,N_7979);
nor U8941 (N_8941,N_7802,N_8114);
or U8942 (N_8942,N_8067,N_8176);
nor U8943 (N_8943,N_7811,N_8016);
nand U8944 (N_8944,N_7532,N_7509);
or U8945 (N_8945,N_7785,N_7601);
or U8946 (N_8946,N_7866,N_8047);
nand U8947 (N_8947,N_7693,N_7959);
xor U8948 (N_8948,N_7859,N_7780);
nand U8949 (N_8949,N_7978,N_7711);
or U8950 (N_8950,N_7991,N_7621);
xor U8951 (N_8951,N_8222,N_7620);
xor U8952 (N_8952,N_8206,N_8142);
or U8953 (N_8953,N_7946,N_8120);
xor U8954 (N_8954,N_7798,N_7524);
and U8955 (N_8955,N_8140,N_8121);
and U8956 (N_8956,N_7751,N_8116);
and U8957 (N_8957,N_8164,N_7653);
and U8958 (N_8958,N_7853,N_7827);
and U8959 (N_8959,N_7516,N_7980);
nor U8960 (N_8960,N_8063,N_7919);
xnor U8961 (N_8961,N_7943,N_8133);
nand U8962 (N_8962,N_7554,N_8139);
or U8963 (N_8963,N_8050,N_7650);
nand U8964 (N_8964,N_7674,N_7997);
xnor U8965 (N_8965,N_8121,N_7853);
nor U8966 (N_8966,N_7514,N_8118);
and U8967 (N_8967,N_7786,N_7520);
or U8968 (N_8968,N_7907,N_8018);
nand U8969 (N_8969,N_7718,N_7739);
nand U8970 (N_8970,N_8026,N_8249);
nor U8971 (N_8971,N_8058,N_7774);
xor U8972 (N_8972,N_8164,N_7986);
xor U8973 (N_8973,N_8188,N_7674);
and U8974 (N_8974,N_7694,N_8151);
nand U8975 (N_8975,N_7548,N_7944);
and U8976 (N_8976,N_8147,N_7600);
xor U8977 (N_8977,N_7661,N_8195);
nand U8978 (N_8978,N_7863,N_7821);
nor U8979 (N_8979,N_8008,N_7504);
or U8980 (N_8980,N_8240,N_7622);
or U8981 (N_8981,N_7975,N_7560);
nand U8982 (N_8982,N_7772,N_8160);
and U8983 (N_8983,N_7960,N_8217);
nand U8984 (N_8984,N_7660,N_7605);
xor U8985 (N_8985,N_8001,N_8172);
xor U8986 (N_8986,N_7949,N_8080);
and U8987 (N_8987,N_7586,N_7763);
xor U8988 (N_8988,N_8142,N_8231);
nor U8989 (N_8989,N_8087,N_7565);
nor U8990 (N_8990,N_8074,N_7847);
or U8991 (N_8991,N_8202,N_8236);
xnor U8992 (N_8992,N_7756,N_8191);
or U8993 (N_8993,N_7820,N_7844);
nor U8994 (N_8994,N_7667,N_7527);
xor U8995 (N_8995,N_7905,N_7592);
nor U8996 (N_8996,N_7528,N_8016);
nand U8997 (N_8997,N_8003,N_8247);
and U8998 (N_8998,N_8122,N_8193);
nand U8999 (N_8999,N_8090,N_7794);
nand U9000 (N_9000,N_8469,N_8654);
and U9001 (N_9001,N_8544,N_8804);
or U9002 (N_9002,N_8782,N_8607);
or U9003 (N_9003,N_8823,N_8472);
or U9004 (N_9004,N_8785,N_8969);
or U9005 (N_9005,N_8966,N_8458);
xnor U9006 (N_9006,N_8563,N_8872);
and U9007 (N_9007,N_8842,N_8790);
nand U9008 (N_9008,N_8453,N_8889);
xor U9009 (N_9009,N_8890,N_8681);
xnor U9010 (N_9010,N_8667,N_8502);
or U9011 (N_9011,N_8620,N_8911);
nor U9012 (N_9012,N_8746,N_8597);
and U9013 (N_9013,N_8987,N_8284);
nor U9014 (N_9014,N_8559,N_8673);
nor U9015 (N_9015,N_8579,N_8335);
and U9016 (N_9016,N_8765,N_8642);
nand U9017 (N_9017,N_8680,N_8379);
nor U9018 (N_9018,N_8767,N_8501);
xnor U9019 (N_9019,N_8250,N_8650);
or U9020 (N_9020,N_8271,N_8991);
nand U9021 (N_9021,N_8256,N_8383);
nor U9022 (N_9022,N_8945,N_8639);
or U9023 (N_9023,N_8314,N_8904);
xor U9024 (N_9024,N_8662,N_8440);
xor U9025 (N_9025,N_8778,N_8404);
nor U9026 (N_9026,N_8677,N_8499);
and U9027 (N_9027,N_8565,N_8611);
or U9028 (N_9028,N_8822,N_8422);
nand U9029 (N_9029,N_8954,N_8818);
nor U9030 (N_9030,N_8533,N_8830);
nand U9031 (N_9031,N_8627,N_8829);
or U9032 (N_9032,N_8512,N_8864);
nand U9033 (N_9033,N_8848,N_8323);
nor U9034 (N_9034,N_8302,N_8994);
nand U9035 (N_9035,N_8752,N_8541);
nor U9036 (N_9036,N_8744,N_8959);
or U9037 (N_9037,N_8919,N_8548);
xor U9038 (N_9038,N_8745,N_8711);
and U9039 (N_9039,N_8814,N_8968);
and U9040 (N_9040,N_8463,N_8508);
or U9041 (N_9041,N_8849,N_8769);
nand U9042 (N_9042,N_8325,N_8255);
or U9043 (N_9043,N_8496,N_8674);
and U9044 (N_9044,N_8443,N_8466);
nand U9045 (N_9045,N_8950,N_8742);
nand U9046 (N_9046,N_8771,N_8598);
xnor U9047 (N_9047,N_8590,N_8976);
nor U9048 (N_9048,N_8798,N_8529);
or U9049 (N_9049,N_8328,N_8303);
xor U9050 (N_9050,N_8339,N_8319);
nor U9051 (N_9051,N_8500,N_8407);
and U9052 (N_9052,N_8977,N_8568);
or U9053 (N_9053,N_8406,N_8887);
nor U9054 (N_9054,N_8329,N_8471);
nor U9055 (N_9055,N_8949,N_8707);
and U9056 (N_9056,N_8573,N_8476);
nand U9057 (N_9057,N_8749,N_8983);
xnor U9058 (N_9058,N_8929,N_8411);
and U9059 (N_9059,N_8768,N_8743);
nand U9060 (N_9060,N_8948,N_8613);
xor U9061 (N_9061,N_8774,N_8831);
nand U9062 (N_9062,N_8535,N_8812);
xnor U9063 (N_9063,N_8253,N_8567);
xnor U9064 (N_9064,N_8886,N_8536);
or U9065 (N_9065,N_8876,N_8805);
or U9066 (N_9066,N_8970,N_8675);
or U9067 (N_9067,N_8432,N_8923);
nor U9068 (N_9068,N_8318,N_8296);
xnor U9069 (N_9069,N_8951,N_8299);
nor U9070 (N_9070,N_8465,N_8275);
and U9071 (N_9071,N_8811,N_8420);
or U9072 (N_9072,N_8352,N_8456);
nand U9073 (N_9073,N_8350,N_8439);
and U9074 (N_9074,N_8288,N_8304);
nand U9075 (N_9075,N_8430,N_8741);
nor U9076 (N_9076,N_8716,N_8461);
xnor U9077 (N_9077,N_8753,N_8897);
and U9078 (N_9078,N_8989,N_8258);
xnor U9079 (N_9079,N_8617,N_8572);
nor U9080 (N_9080,N_8699,N_8434);
nor U9081 (N_9081,N_8298,N_8342);
or U9082 (N_9082,N_8348,N_8761);
or U9083 (N_9083,N_8960,N_8931);
and U9084 (N_9084,N_8610,N_8832);
or U9085 (N_9085,N_8580,N_8901);
nor U9086 (N_9086,N_8491,N_8845);
nor U9087 (N_9087,N_8262,N_8656);
nor U9088 (N_9088,N_8436,N_8295);
and U9089 (N_9089,N_8369,N_8583);
or U9090 (N_9090,N_8837,N_8574);
or U9091 (N_9091,N_8530,N_8622);
nor U9092 (N_9092,N_8554,N_8449);
nand U9093 (N_9093,N_8935,N_8297);
nor U9094 (N_9094,N_8992,N_8273);
or U9095 (N_9095,N_8788,N_8435);
xor U9096 (N_9096,N_8955,N_8702);
and U9097 (N_9097,N_8939,N_8584);
or U9098 (N_9098,N_8921,N_8657);
nor U9099 (N_9099,N_8853,N_8942);
nand U9100 (N_9100,N_8446,N_8514);
and U9101 (N_9101,N_8313,N_8557);
nor U9102 (N_9102,N_8286,N_8370);
xnor U9103 (N_9103,N_8448,N_8967);
and U9104 (N_9104,N_8807,N_8364);
or U9105 (N_9105,N_8760,N_8569);
and U9106 (N_9106,N_8551,N_8894);
xor U9107 (N_9107,N_8927,N_8683);
and U9108 (N_9108,N_8511,N_8386);
nand U9109 (N_9109,N_8531,N_8577);
xor U9110 (N_9110,N_8281,N_8758);
and U9111 (N_9111,N_8308,N_8547);
nand U9112 (N_9112,N_8263,N_8885);
xor U9113 (N_9113,N_8810,N_8267);
or U9114 (N_9114,N_8292,N_8558);
or U9115 (N_9115,N_8578,N_8697);
xnor U9116 (N_9116,N_8854,N_8852);
xor U9117 (N_9117,N_8777,N_8254);
and U9118 (N_9118,N_8869,N_8477);
nand U9119 (N_9119,N_8623,N_8715);
or U9120 (N_9120,N_8803,N_8631);
and U9121 (N_9121,N_8340,N_8384);
xor U9122 (N_9122,N_8635,N_8616);
or U9123 (N_9123,N_8827,N_8698);
and U9124 (N_9124,N_8513,N_8806);
or U9125 (N_9125,N_8817,N_8884);
nor U9126 (N_9126,N_8293,N_8920);
or U9127 (N_9127,N_8892,N_8349);
xor U9128 (N_9128,N_8858,N_8628);
xor U9129 (N_9129,N_8320,N_8772);
nand U9130 (N_9130,N_8265,N_8995);
nor U9131 (N_9131,N_8612,N_8757);
nor U9132 (N_9132,N_8542,N_8965);
or U9133 (N_9133,N_8478,N_8695);
xnor U9134 (N_9134,N_8280,N_8980);
nand U9135 (N_9135,N_8799,N_8570);
nor U9136 (N_9136,N_8736,N_8787);
xor U9137 (N_9137,N_8507,N_8734);
or U9138 (N_9138,N_8474,N_8641);
xor U9139 (N_9139,N_8368,N_8487);
nand U9140 (N_9140,N_8305,N_8726);
or U9141 (N_9141,N_8691,N_8483);
or U9142 (N_9142,N_8730,N_8464);
xnor U9143 (N_9143,N_8984,N_8510);
and U9144 (N_9144,N_8614,N_8390);
nor U9145 (N_9145,N_8581,N_8851);
xor U9146 (N_9146,N_8345,N_8525);
nand U9147 (N_9147,N_8721,N_8910);
or U9148 (N_9148,N_8428,N_8523);
nor U9149 (N_9149,N_8728,N_8337);
nor U9150 (N_9150,N_8532,N_8534);
nor U9151 (N_9151,N_8791,N_8421);
xor U9152 (N_9152,N_8676,N_8264);
nor U9153 (N_9153,N_8938,N_8330);
xor U9154 (N_9154,N_8317,N_8725);
xor U9155 (N_9155,N_8395,N_8649);
and U9156 (N_9156,N_8326,N_8809);
or U9157 (N_9157,N_8835,N_8587);
and U9158 (N_9158,N_8378,N_8855);
nor U9159 (N_9159,N_8593,N_8515);
and U9160 (N_9160,N_8908,N_8795);
nand U9161 (N_9161,N_8594,N_8444);
nor U9162 (N_9162,N_8333,N_8652);
xor U9163 (N_9163,N_8450,N_8779);
and U9164 (N_9164,N_8737,N_8724);
or U9165 (N_9165,N_8618,N_8455);
xor U9166 (N_9166,N_8926,N_8978);
nand U9167 (N_9167,N_8874,N_8429);
and U9168 (N_9168,N_8401,N_8306);
xor U9169 (N_9169,N_8696,N_8415);
or U9170 (N_9170,N_8601,N_8895);
xnor U9171 (N_9171,N_8905,N_8585);
nand U9172 (N_9172,N_8596,N_8821);
or U9173 (N_9173,N_8688,N_8426);
or U9174 (N_9174,N_8403,N_8924);
and U9175 (N_9175,N_8841,N_8608);
or U9176 (N_9176,N_8468,N_8883);
xnor U9177 (N_9177,N_8640,N_8538);
xor U9178 (N_9178,N_8492,N_8670);
and U9179 (N_9179,N_8621,N_8868);
or U9180 (N_9180,N_8906,N_8915);
xor U9181 (N_9181,N_8747,N_8371);
and U9182 (N_9182,N_8647,N_8494);
or U9183 (N_9183,N_8900,N_8679);
xnor U9184 (N_9184,N_8381,N_8843);
nand U9185 (N_9185,N_8710,N_8706);
xnor U9186 (N_9186,N_8417,N_8375);
or U9187 (N_9187,N_8940,N_8366);
and U9188 (N_9188,N_8775,N_8509);
and U9189 (N_9189,N_8916,N_8773);
xor U9190 (N_9190,N_8988,N_8682);
or U9191 (N_9191,N_8961,N_8668);
nand U9192 (N_9192,N_8985,N_8633);
and U9193 (N_9193,N_8755,N_8871);
nand U9194 (N_9194,N_8850,N_8460);
and U9195 (N_9195,N_8840,N_8527);
or U9196 (N_9196,N_8703,N_8555);
or U9197 (N_9197,N_8438,N_8713);
nor U9198 (N_9198,N_8424,N_8686);
and U9199 (N_9199,N_8972,N_8933);
nand U9200 (N_9200,N_8309,N_8341);
xnor U9201 (N_9201,N_8784,N_8624);
xnor U9202 (N_9202,N_8545,N_8833);
and U9203 (N_9203,N_8964,N_8692);
nor U9204 (N_9204,N_8467,N_8609);
nor U9205 (N_9205,N_8591,N_8537);
nor U9206 (N_9206,N_8934,N_8781);
nor U9207 (N_9207,N_8367,N_8459);
nor U9208 (N_9208,N_8655,N_8452);
or U9209 (N_9209,N_8283,N_8431);
and U9210 (N_9210,N_8793,N_8376);
xor U9211 (N_9211,N_8353,N_8651);
or U9212 (N_9212,N_8820,N_8861);
nor U9213 (N_9213,N_8776,N_8457);
and U9214 (N_9214,N_8740,N_8504);
or U9215 (N_9215,N_8522,N_8786);
nor U9216 (N_9216,N_8997,N_8602);
and U9217 (N_9217,N_8981,N_8354);
nand U9218 (N_9218,N_8719,N_8361);
xnor U9219 (N_9219,N_8846,N_8416);
nand U9220 (N_9220,N_8277,N_8907);
xor U9221 (N_9221,N_8355,N_8727);
nor U9222 (N_9222,N_8881,N_8660);
and U9223 (N_9223,N_8363,N_8630);
or U9224 (N_9224,N_8338,N_8556);
xor U9225 (N_9225,N_8517,N_8310);
nand U9226 (N_9226,N_8944,N_8252);
or U9227 (N_9227,N_8859,N_8482);
nor U9228 (N_9228,N_8257,N_8402);
and U9229 (N_9229,N_8604,N_8528);
nor U9230 (N_9230,N_8344,N_8372);
xor U9231 (N_9231,N_8836,N_8373);
nor U9232 (N_9232,N_8327,N_8414);
nor U9233 (N_9233,N_8731,N_8956);
and U9234 (N_9234,N_8285,N_8629);
nor U9235 (N_9235,N_8689,N_8526);
or U9236 (N_9236,N_8615,N_8825);
nor U9237 (N_9237,N_8802,N_8705);
xnor U9238 (N_9238,N_8913,N_8433);
nand U9239 (N_9239,N_8879,N_8392);
and U9240 (N_9240,N_8334,N_8918);
nor U9241 (N_9241,N_8909,N_8717);
nor U9242 (N_9242,N_8419,N_8770);
nor U9243 (N_9243,N_8437,N_8272);
and U9244 (N_9244,N_8606,N_8925);
and U9245 (N_9245,N_8947,N_8684);
or U9246 (N_9246,N_8358,N_8266);
nor U9247 (N_9247,N_8762,N_8418);
and U9248 (N_9248,N_8550,N_8505);
nor U9249 (N_9249,N_8953,N_8539);
nand U9250 (N_9250,N_8860,N_8882);
nand U9251 (N_9251,N_8503,N_8946);
nor U9252 (N_9252,N_8644,N_8495);
or U9253 (N_9253,N_8932,N_8723);
or U9254 (N_9254,N_8636,N_8553);
nor U9255 (N_9255,N_8490,N_8963);
nor U9256 (N_9256,N_8643,N_8400);
nor U9257 (N_9257,N_8754,N_8261);
nor U9258 (N_9258,N_8626,N_8739);
and U9259 (N_9259,N_8473,N_8700);
nor U9260 (N_9260,N_8405,N_8996);
or U9261 (N_9261,N_8891,N_8764);
nand U9262 (N_9262,N_8289,N_8941);
nand U9263 (N_9263,N_8866,N_8425);
xnor U9264 (N_9264,N_8479,N_8387);
nand U9265 (N_9265,N_8564,N_8797);
xor U9266 (N_9266,N_8592,N_8709);
and U9267 (N_9267,N_8546,N_8856);
nor U9268 (N_9268,N_8357,N_8315);
nor U9269 (N_9269,N_8780,N_8658);
and U9270 (N_9270,N_8666,N_8552);
nor U9271 (N_9271,N_8332,N_8862);
nor U9272 (N_9272,N_8763,N_8394);
nand U9273 (N_9273,N_8493,N_8993);
or U9274 (N_9274,N_8454,N_8637);
and U9275 (N_9275,N_8973,N_8582);
nor U9276 (N_9276,N_8575,N_8990);
xor U9277 (N_9277,N_8671,N_8413);
xor U9278 (N_9278,N_8398,N_8952);
or U9279 (N_9279,N_8322,N_8520);
xor U9280 (N_9280,N_8914,N_8307);
and U9281 (N_9281,N_8516,N_8819);
and U9282 (N_9282,N_8447,N_8377);
nor U9283 (N_9283,N_8279,N_8690);
and U9284 (N_9284,N_8873,N_8979);
xnor U9285 (N_9285,N_8408,N_8792);
nor U9286 (N_9286,N_8708,N_8576);
nand U9287 (N_9287,N_8571,N_8380);
nor U9288 (N_9288,N_8276,N_8665);
or U9289 (N_9289,N_8646,N_8259);
and U9290 (N_9290,N_8365,N_8748);
nand U9291 (N_9291,N_8423,N_8750);
nand U9292 (N_9292,N_8290,N_8957);
nor U9293 (N_9293,N_8999,N_8485);
nand U9294 (N_9294,N_8603,N_8470);
or U9295 (N_9295,N_8974,N_8374);
nor U9296 (N_9296,N_8687,N_8701);
and U9297 (N_9297,N_8789,N_8385);
or U9298 (N_9298,N_8847,N_8560);
nor U9299 (N_9299,N_8412,N_8347);
nand U9300 (N_9300,N_8712,N_8922);
nor U9301 (N_9301,N_8704,N_8489);
xor U9302 (N_9302,N_8917,N_8834);
and U9303 (N_9303,N_8351,N_8393);
nor U9304 (N_9304,N_8540,N_8462);
nand U9305 (N_9305,N_8270,N_8632);
and U9306 (N_9306,N_8783,N_8903);
nand U9307 (N_9307,N_8998,N_8751);
nor U9308 (N_9308,N_8720,N_8824);
nand U9309 (N_9309,N_8863,N_8937);
nand U9310 (N_9310,N_8898,N_8796);
or U9311 (N_9311,N_8388,N_8870);
nand U9312 (N_9312,N_8356,N_8800);
xor U9313 (N_9313,N_8659,N_8902);
and U9314 (N_9314,N_8678,N_8880);
nand U9315 (N_9315,N_8480,N_8312);
nor U9316 (N_9316,N_8738,N_8694);
and U9317 (N_9317,N_8878,N_8484);
and U9318 (N_9318,N_8519,N_8664);
xnor U9319 (N_9319,N_8943,N_8794);
nand U9320 (N_9320,N_8888,N_8278);
nor U9321 (N_9321,N_8648,N_8638);
or U9322 (N_9322,N_8549,N_8441);
or U9323 (N_9323,N_8653,N_8324);
or U9324 (N_9324,N_8685,N_8475);
xor U9325 (N_9325,N_8282,N_8971);
nand U9326 (N_9326,N_8486,N_8801);
nor U9327 (N_9327,N_8766,N_8294);
nand U9328 (N_9328,N_8359,N_8321);
or U9329 (N_9329,N_8300,N_8928);
xor U9330 (N_9330,N_8481,N_8409);
and U9331 (N_9331,N_8815,N_8930);
nor U9332 (N_9332,N_8269,N_8669);
or U9333 (N_9333,N_8877,N_8586);
or U9334 (N_9334,N_8729,N_8506);
or U9335 (N_9335,N_8498,N_8975);
or U9336 (N_9336,N_8396,N_8693);
nor U9337 (N_9337,N_8936,N_8756);
xor U9338 (N_9338,N_8518,N_8759);
nor U9339 (N_9339,N_8912,N_8331);
nor U9340 (N_9340,N_8808,N_8291);
nand U9341 (N_9341,N_8982,N_8251);
nor U9342 (N_9342,N_8661,N_8733);
nor U9343 (N_9343,N_8488,N_8867);
nand U9344 (N_9344,N_8360,N_8718);
nor U9345 (N_9345,N_8524,N_8311);
nor U9346 (N_9346,N_8497,N_8857);
and U9347 (N_9347,N_8287,N_8816);
xor U9348 (N_9348,N_8893,N_8427);
nand U9349 (N_9349,N_8599,N_8838);
or U9350 (N_9350,N_8619,N_8839);
xor U9351 (N_9351,N_8600,N_8826);
xnor U9352 (N_9352,N_8986,N_8589);
nor U9353 (N_9353,N_8813,N_8346);
nand U9354 (N_9354,N_8451,N_8588);
nand U9355 (N_9355,N_8260,N_8828);
nand U9356 (N_9356,N_8735,N_8382);
nand U9357 (N_9357,N_8896,N_8714);
nand U9358 (N_9358,N_8566,N_8442);
nor U9359 (N_9359,N_8645,N_8634);
and U9360 (N_9360,N_8625,N_8521);
nand U9361 (N_9361,N_8672,N_8336);
or U9362 (N_9362,N_8543,N_8958);
nor U9363 (N_9363,N_8391,N_8962);
nand U9364 (N_9364,N_8316,N_8663);
nor U9365 (N_9365,N_8274,N_8397);
or U9366 (N_9366,N_8268,N_8605);
nand U9367 (N_9367,N_8722,N_8562);
and U9368 (N_9368,N_8399,N_8844);
nor U9369 (N_9369,N_8410,N_8561);
nor U9370 (N_9370,N_8875,N_8732);
xnor U9371 (N_9371,N_8595,N_8389);
or U9372 (N_9372,N_8899,N_8362);
and U9373 (N_9373,N_8445,N_8865);
xor U9374 (N_9374,N_8343,N_8301);
nand U9375 (N_9375,N_8367,N_8352);
xnor U9376 (N_9376,N_8656,N_8889);
xnor U9377 (N_9377,N_8459,N_8780);
or U9378 (N_9378,N_8382,N_8983);
nor U9379 (N_9379,N_8283,N_8888);
nand U9380 (N_9380,N_8308,N_8601);
nand U9381 (N_9381,N_8264,N_8933);
nor U9382 (N_9382,N_8835,N_8912);
nor U9383 (N_9383,N_8665,N_8823);
nor U9384 (N_9384,N_8895,N_8633);
nand U9385 (N_9385,N_8427,N_8830);
nand U9386 (N_9386,N_8671,N_8861);
nand U9387 (N_9387,N_8683,N_8830);
nand U9388 (N_9388,N_8678,N_8562);
nand U9389 (N_9389,N_8571,N_8366);
and U9390 (N_9390,N_8332,N_8361);
nor U9391 (N_9391,N_8694,N_8709);
nor U9392 (N_9392,N_8691,N_8341);
and U9393 (N_9393,N_8888,N_8970);
nand U9394 (N_9394,N_8485,N_8305);
or U9395 (N_9395,N_8609,N_8417);
nand U9396 (N_9396,N_8851,N_8822);
or U9397 (N_9397,N_8698,N_8634);
or U9398 (N_9398,N_8344,N_8619);
xnor U9399 (N_9399,N_8366,N_8663);
and U9400 (N_9400,N_8945,N_8640);
xnor U9401 (N_9401,N_8737,N_8789);
or U9402 (N_9402,N_8871,N_8931);
xor U9403 (N_9403,N_8409,N_8254);
or U9404 (N_9404,N_8976,N_8356);
nand U9405 (N_9405,N_8755,N_8502);
nor U9406 (N_9406,N_8585,N_8367);
xnor U9407 (N_9407,N_8810,N_8910);
nor U9408 (N_9408,N_8783,N_8712);
or U9409 (N_9409,N_8663,N_8736);
and U9410 (N_9410,N_8592,N_8880);
xnor U9411 (N_9411,N_8498,N_8358);
and U9412 (N_9412,N_8964,N_8481);
nand U9413 (N_9413,N_8907,N_8955);
or U9414 (N_9414,N_8958,N_8352);
nor U9415 (N_9415,N_8753,N_8275);
xnor U9416 (N_9416,N_8947,N_8332);
xnor U9417 (N_9417,N_8616,N_8325);
xnor U9418 (N_9418,N_8494,N_8476);
nor U9419 (N_9419,N_8913,N_8589);
and U9420 (N_9420,N_8661,N_8410);
nand U9421 (N_9421,N_8431,N_8279);
or U9422 (N_9422,N_8751,N_8544);
nand U9423 (N_9423,N_8493,N_8712);
and U9424 (N_9424,N_8981,N_8992);
xnor U9425 (N_9425,N_8907,N_8333);
and U9426 (N_9426,N_8456,N_8964);
or U9427 (N_9427,N_8785,N_8510);
xor U9428 (N_9428,N_8876,N_8999);
and U9429 (N_9429,N_8655,N_8540);
xor U9430 (N_9430,N_8874,N_8965);
nand U9431 (N_9431,N_8866,N_8466);
nand U9432 (N_9432,N_8498,N_8303);
xnor U9433 (N_9433,N_8668,N_8933);
nor U9434 (N_9434,N_8628,N_8982);
xor U9435 (N_9435,N_8742,N_8887);
or U9436 (N_9436,N_8635,N_8483);
nor U9437 (N_9437,N_8683,N_8337);
nor U9438 (N_9438,N_8837,N_8735);
xor U9439 (N_9439,N_8713,N_8866);
or U9440 (N_9440,N_8839,N_8354);
nand U9441 (N_9441,N_8484,N_8542);
xor U9442 (N_9442,N_8767,N_8762);
xnor U9443 (N_9443,N_8537,N_8800);
nand U9444 (N_9444,N_8563,N_8989);
nand U9445 (N_9445,N_8302,N_8821);
or U9446 (N_9446,N_8796,N_8811);
nor U9447 (N_9447,N_8427,N_8768);
nand U9448 (N_9448,N_8486,N_8277);
or U9449 (N_9449,N_8270,N_8408);
nand U9450 (N_9450,N_8529,N_8431);
nand U9451 (N_9451,N_8732,N_8673);
or U9452 (N_9452,N_8727,N_8300);
and U9453 (N_9453,N_8513,N_8366);
nor U9454 (N_9454,N_8606,N_8778);
or U9455 (N_9455,N_8482,N_8739);
xnor U9456 (N_9456,N_8792,N_8332);
or U9457 (N_9457,N_8250,N_8767);
xor U9458 (N_9458,N_8432,N_8545);
or U9459 (N_9459,N_8674,N_8886);
and U9460 (N_9460,N_8927,N_8573);
nand U9461 (N_9461,N_8770,N_8890);
and U9462 (N_9462,N_8871,N_8312);
nor U9463 (N_9463,N_8446,N_8301);
and U9464 (N_9464,N_8749,N_8268);
xnor U9465 (N_9465,N_8397,N_8995);
and U9466 (N_9466,N_8974,N_8317);
nand U9467 (N_9467,N_8997,N_8735);
nand U9468 (N_9468,N_8925,N_8755);
or U9469 (N_9469,N_8466,N_8320);
or U9470 (N_9470,N_8797,N_8713);
nand U9471 (N_9471,N_8502,N_8703);
xor U9472 (N_9472,N_8908,N_8574);
xnor U9473 (N_9473,N_8821,N_8871);
nor U9474 (N_9474,N_8400,N_8926);
xor U9475 (N_9475,N_8493,N_8899);
nand U9476 (N_9476,N_8324,N_8756);
xor U9477 (N_9477,N_8838,N_8736);
and U9478 (N_9478,N_8552,N_8877);
xnor U9479 (N_9479,N_8656,N_8457);
nor U9480 (N_9480,N_8777,N_8544);
and U9481 (N_9481,N_8522,N_8918);
nor U9482 (N_9482,N_8363,N_8788);
and U9483 (N_9483,N_8766,N_8486);
or U9484 (N_9484,N_8376,N_8959);
xor U9485 (N_9485,N_8639,N_8392);
nor U9486 (N_9486,N_8656,N_8953);
nand U9487 (N_9487,N_8561,N_8611);
or U9488 (N_9488,N_8350,N_8956);
nand U9489 (N_9489,N_8454,N_8874);
nor U9490 (N_9490,N_8514,N_8451);
or U9491 (N_9491,N_8543,N_8259);
nor U9492 (N_9492,N_8460,N_8977);
nor U9493 (N_9493,N_8776,N_8432);
xor U9494 (N_9494,N_8866,N_8921);
and U9495 (N_9495,N_8899,N_8762);
xor U9496 (N_9496,N_8990,N_8925);
or U9497 (N_9497,N_8634,N_8429);
or U9498 (N_9498,N_8446,N_8305);
or U9499 (N_9499,N_8917,N_8443);
nor U9500 (N_9500,N_8590,N_8588);
xor U9501 (N_9501,N_8704,N_8897);
nand U9502 (N_9502,N_8300,N_8776);
and U9503 (N_9503,N_8916,N_8308);
nor U9504 (N_9504,N_8808,N_8474);
and U9505 (N_9505,N_8833,N_8746);
nand U9506 (N_9506,N_8699,N_8437);
and U9507 (N_9507,N_8868,N_8498);
nor U9508 (N_9508,N_8622,N_8995);
nand U9509 (N_9509,N_8769,N_8374);
nand U9510 (N_9510,N_8583,N_8469);
xor U9511 (N_9511,N_8273,N_8965);
and U9512 (N_9512,N_8410,N_8464);
and U9513 (N_9513,N_8973,N_8500);
xor U9514 (N_9514,N_8692,N_8552);
nor U9515 (N_9515,N_8694,N_8609);
or U9516 (N_9516,N_8891,N_8710);
xnor U9517 (N_9517,N_8907,N_8415);
or U9518 (N_9518,N_8415,N_8760);
nand U9519 (N_9519,N_8550,N_8405);
and U9520 (N_9520,N_8551,N_8258);
nand U9521 (N_9521,N_8574,N_8761);
or U9522 (N_9522,N_8355,N_8981);
and U9523 (N_9523,N_8451,N_8557);
nor U9524 (N_9524,N_8987,N_8846);
and U9525 (N_9525,N_8893,N_8338);
xnor U9526 (N_9526,N_8628,N_8713);
xor U9527 (N_9527,N_8478,N_8825);
and U9528 (N_9528,N_8728,N_8475);
nor U9529 (N_9529,N_8917,N_8612);
and U9530 (N_9530,N_8333,N_8341);
nor U9531 (N_9531,N_8632,N_8337);
nor U9532 (N_9532,N_8648,N_8787);
and U9533 (N_9533,N_8681,N_8976);
nor U9534 (N_9534,N_8678,N_8623);
nand U9535 (N_9535,N_8299,N_8592);
nand U9536 (N_9536,N_8939,N_8856);
xnor U9537 (N_9537,N_8940,N_8947);
xnor U9538 (N_9538,N_8922,N_8703);
and U9539 (N_9539,N_8946,N_8534);
and U9540 (N_9540,N_8576,N_8671);
xor U9541 (N_9541,N_8904,N_8542);
and U9542 (N_9542,N_8957,N_8386);
or U9543 (N_9543,N_8592,N_8359);
nor U9544 (N_9544,N_8271,N_8671);
nor U9545 (N_9545,N_8282,N_8563);
xnor U9546 (N_9546,N_8836,N_8290);
xnor U9547 (N_9547,N_8629,N_8775);
nor U9548 (N_9548,N_8980,N_8319);
or U9549 (N_9549,N_8594,N_8535);
xnor U9550 (N_9550,N_8467,N_8297);
xor U9551 (N_9551,N_8623,N_8304);
and U9552 (N_9552,N_8982,N_8558);
nand U9553 (N_9553,N_8510,N_8579);
or U9554 (N_9554,N_8490,N_8313);
nor U9555 (N_9555,N_8948,N_8843);
nor U9556 (N_9556,N_8327,N_8549);
nor U9557 (N_9557,N_8982,N_8589);
or U9558 (N_9558,N_8919,N_8729);
and U9559 (N_9559,N_8435,N_8370);
or U9560 (N_9560,N_8710,N_8341);
or U9561 (N_9561,N_8388,N_8780);
xnor U9562 (N_9562,N_8798,N_8434);
xnor U9563 (N_9563,N_8423,N_8898);
or U9564 (N_9564,N_8266,N_8947);
nand U9565 (N_9565,N_8604,N_8332);
or U9566 (N_9566,N_8292,N_8843);
xnor U9567 (N_9567,N_8925,N_8270);
nand U9568 (N_9568,N_8562,N_8649);
nor U9569 (N_9569,N_8857,N_8776);
xor U9570 (N_9570,N_8357,N_8538);
or U9571 (N_9571,N_8947,N_8386);
nor U9572 (N_9572,N_8775,N_8797);
and U9573 (N_9573,N_8872,N_8674);
nand U9574 (N_9574,N_8600,N_8520);
or U9575 (N_9575,N_8369,N_8256);
nor U9576 (N_9576,N_8315,N_8811);
nor U9577 (N_9577,N_8694,N_8942);
xor U9578 (N_9578,N_8795,N_8480);
nand U9579 (N_9579,N_8816,N_8807);
nor U9580 (N_9580,N_8293,N_8814);
nand U9581 (N_9581,N_8818,N_8323);
nand U9582 (N_9582,N_8980,N_8591);
nor U9583 (N_9583,N_8488,N_8505);
xnor U9584 (N_9584,N_8794,N_8802);
or U9585 (N_9585,N_8616,N_8757);
nand U9586 (N_9586,N_8893,N_8754);
and U9587 (N_9587,N_8736,N_8859);
nand U9588 (N_9588,N_8661,N_8607);
xnor U9589 (N_9589,N_8521,N_8939);
and U9590 (N_9590,N_8527,N_8429);
xor U9591 (N_9591,N_8644,N_8306);
xnor U9592 (N_9592,N_8593,N_8815);
and U9593 (N_9593,N_8985,N_8974);
or U9594 (N_9594,N_8904,N_8613);
nand U9595 (N_9595,N_8444,N_8767);
nand U9596 (N_9596,N_8752,N_8986);
or U9597 (N_9597,N_8746,N_8469);
or U9598 (N_9598,N_8777,N_8984);
nor U9599 (N_9599,N_8855,N_8418);
or U9600 (N_9600,N_8902,N_8666);
and U9601 (N_9601,N_8823,N_8288);
and U9602 (N_9602,N_8719,N_8274);
nand U9603 (N_9603,N_8821,N_8462);
and U9604 (N_9604,N_8417,N_8401);
and U9605 (N_9605,N_8372,N_8686);
xor U9606 (N_9606,N_8795,N_8345);
or U9607 (N_9607,N_8539,N_8744);
xnor U9608 (N_9608,N_8881,N_8651);
nand U9609 (N_9609,N_8990,N_8733);
xnor U9610 (N_9610,N_8789,N_8452);
nor U9611 (N_9611,N_8569,N_8395);
nand U9612 (N_9612,N_8886,N_8809);
or U9613 (N_9613,N_8368,N_8895);
or U9614 (N_9614,N_8635,N_8632);
xor U9615 (N_9615,N_8594,N_8917);
xnor U9616 (N_9616,N_8319,N_8779);
nand U9617 (N_9617,N_8621,N_8462);
nand U9618 (N_9618,N_8333,N_8261);
xor U9619 (N_9619,N_8883,N_8902);
nand U9620 (N_9620,N_8485,N_8347);
and U9621 (N_9621,N_8304,N_8994);
nand U9622 (N_9622,N_8381,N_8650);
or U9623 (N_9623,N_8353,N_8675);
or U9624 (N_9624,N_8876,N_8573);
xnor U9625 (N_9625,N_8875,N_8521);
or U9626 (N_9626,N_8627,N_8896);
nor U9627 (N_9627,N_8445,N_8834);
and U9628 (N_9628,N_8714,N_8971);
xor U9629 (N_9629,N_8351,N_8557);
or U9630 (N_9630,N_8631,N_8738);
nor U9631 (N_9631,N_8686,N_8944);
or U9632 (N_9632,N_8565,N_8751);
nor U9633 (N_9633,N_8317,N_8307);
xnor U9634 (N_9634,N_8747,N_8565);
and U9635 (N_9635,N_8467,N_8929);
and U9636 (N_9636,N_8917,N_8585);
nor U9637 (N_9637,N_8928,N_8351);
xor U9638 (N_9638,N_8421,N_8447);
xor U9639 (N_9639,N_8420,N_8770);
nor U9640 (N_9640,N_8593,N_8633);
xor U9641 (N_9641,N_8779,N_8296);
xnor U9642 (N_9642,N_8750,N_8986);
and U9643 (N_9643,N_8966,N_8790);
nand U9644 (N_9644,N_8572,N_8635);
or U9645 (N_9645,N_8324,N_8336);
nand U9646 (N_9646,N_8540,N_8812);
nor U9647 (N_9647,N_8844,N_8684);
xnor U9648 (N_9648,N_8493,N_8875);
and U9649 (N_9649,N_8661,N_8763);
and U9650 (N_9650,N_8879,N_8277);
xnor U9651 (N_9651,N_8758,N_8355);
and U9652 (N_9652,N_8645,N_8331);
or U9653 (N_9653,N_8935,N_8516);
and U9654 (N_9654,N_8400,N_8555);
and U9655 (N_9655,N_8978,N_8975);
xor U9656 (N_9656,N_8874,N_8942);
nand U9657 (N_9657,N_8475,N_8401);
nor U9658 (N_9658,N_8971,N_8631);
nand U9659 (N_9659,N_8702,N_8733);
nand U9660 (N_9660,N_8926,N_8314);
nor U9661 (N_9661,N_8960,N_8335);
or U9662 (N_9662,N_8506,N_8774);
or U9663 (N_9663,N_8387,N_8274);
and U9664 (N_9664,N_8446,N_8919);
xnor U9665 (N_9665,N_8904,N_8688);
nand U9666 (N_9666,N_8548,N_8683);
nor U9667 (N_9667,N_8813,N_8307);
xor U9668 (N_9668,N_8346,N_8945);
and U9669 (N_9669,N_8626,N_8408);
nand U9670 (N_9670,N_8719,N_8818);
nand U9671 (N_9671,N_8419,N_8842);
xor U9672 (N_9672,N_8255,N_8643);
or U9673 (N_9673,N_8397,N_8475);
nor U9674 (N_9674,N_8967,N_8537);
and U9675 (N_9675,N_8635,N_8320);
and U9676 (N_9676,N_8451,N_8258);
nor U9677 (N_9677,N_8513,N_8830);
xor U9678 (N_9678,N_8752,N_8951);
nand U9679 (N_9679,N_8540,N_8915);
and U9680 (N_9680,N_8948,N_8806);
nand U9681 (N_9681,N_8257,N_8330);
or U9682 (N_9682,N_8864,N_8842);
xor U9683 (N_9683,N_8422,N_8549);
xnor U9684 (N_9684,N_8441,N_8344);
or U9685 (N_9685,N_8346,N_8405);
nand U9686 (N_9686,N_8954,N_8940);
and U9687 (N_9687,N_8395,N_8427);
xnor U9688 (N_9688,N_8785,N_8609);
nor U9689 (N_9689,N_8865,N_8827);
nand U9690 (N_9690,N_8602,N_8632);
nor U9691 (N_9691,N_8607,N_8944);
xor U9692 (N_9692,N_8492,N_8514);
nor U9693 (N_9693,N_8381,N_8871);
xnor U9694 (N_9694,N_8599,N_8883);
or U9695 (N_9695,N_8604,N_8792);
nand U9696 (N_9696,N_8775,N_8947);
and U9697 (N_9697,N_8316,N_8597);
and U9698 (N_9698,N_8541,N_8876);
xnor U9699 (N_9699,N_8815,N_8457);
or U9700 (N_9700,N_8430,N_8306);
or U9701 (N_9701,N_8514,N_8612);
nor U9702 (N_9702,N_8811,N_8997);
xor U9703 (N_9703,N_8490,N_8924);
nor U9704 (N_9704,N_8711,N_8365);
xnor U9705 (N_9705,N_8877,N_8412);
or U9706 (N_9706,N_8937,N_8684);
xnor U9707 (N_9707,N_8770,N_8617);
and U9708 (N_9708,N_8884,N_8334);
and U9709 (N_9709,N_8471,N_8376);
or U9710 (N_9710,N_8545,N_8647);
xnor U9711 (N_9711,N_8642,N_8795);
nand U9712 (N_9712,N_8596,N_8612);
and U9713 (N_9713,N_8320,N_8564);
xor U9714 (N_9714,N_8729,N_8780);
nand U9715 (N_9715,N_8771,N_8632);
nand U9716 (N_9716,N_8590,N_8949);
xor U9717 (N_9717,N_8926,N_8567);
nor U9718 (N_9718,N_8896,N_8638);
xor U9719 (N_9719,N_8736,N_8772);
and U9720 (N_9720,N_8759,N_8325);
xnor U9721 (N_9721,N_8757,N_8830);
nor U9722 (N_9722,N_8861,N_8605);
nand U9723 (N_9723,N_8879,N_8544);
nor U9724 (N_9724,N_8421,N_8958);
or U9725 (N_9725,N_8926,N_8797);
xor U9726 (N_9726,N_8629,N_8881);
or U9727 (N_9727,N_8644,N_8634);
xnor U9728 (N_9728,N_8364,N_8967);
nor U9729 (N_9729,N_8341,N_8274);
nand U9730 (N_9730,N_8996,N_8795);
nand U9731 (N_9731,N_8754,N_8289);
nor U9732 (N_9732,N_8983,N_8850);
and U9733 (N_9733,N_8748,N_8413);
and U9734 (N_9734,N_8904,N_8380);
nand U9735 (N_9735,N_8290,N_8367);
or U9736 (N_9736,N_8441,N_8939);
nor U9737 (N_9737,N_8629,N_8454);
nand U9738 (N_9738,N_8259,N_8392);
nor U9739 (N_9739,N_8481,N_8492);
nand U9740 (N_9740,N_8635,N_8407);
nor U9741 (N_9741,N_8286,N_8620);
xnor U9742 (N_9742,N_8895,N_8901);
xnor U9743 (N_9743,N_8693,N_8808);
xor U9744 (N_9744,N_8940,N_8382);
nor U9745 (N_9745,N_8978,N_8746);
nand U9746 (N_9746,N_8380,N_8689);
nor U9747 (N_9747,N_8475,N_8698);
xor U9748 (N_9748,N_8846,N_8570);
nor U9749 (N_9749,N_8330,N_8822);
nand U9750 (N_9750,N_9170,N_9366);
and U9751 (N_9751,N_9495,N_9109);
xnor U9752 (N_9752,N_9613,N_9636);
and U9753 (N_9753,N_9196,N_9245);
nor U9754 (N_9754,N_9461,N_9138);
or U9755 (N_9755,N_9358,N_9313);
or U9756 (N_9756,N_9670,N_9431);
nand U9757 (N_9757,N_9097,N_9561);
or U9758 (N_9758,N_9375,N_9088);
and U9759 (N_9759,N_9304,N_9585);
or U9760 (N_9760,N_9091,N_9362);
xnor U9761 (N_9761,N_9122,N_9051);
or U9762 (N_9762,N_9294,N_9714);
nor U9763 (N_9763,N_9319,N_9413);
nor U9764 (N_9764,N_9127,N_9536);
and U9765 (N_9765,N_9404,N_9655);
xor U9766 (N_9766,N_9494,N_9333);
xnor U9767 (N_9767,N_9509,N_9022);
xnor U9768 (N_9768,N_9074,N_9142);
and U9769 (N_9769,N_9441,N_9554);
or U9770 (N_9770,N_9443,N_9310);
or U9771 (N_9771,N_9639,N_9629);
nand U9772 (N_9772,N_9457,N_9155);
xnor U9773 (N_9773,N_9606,N_9566);
xor U9774 (N_9774,N_9403,N_9252);
xor U9775 (N_9775,N_9490,N_9104);
xor U9776 (N_9776,N_9481,N_9545);
nor U9777 (N_9777,N_9343,N_9349);
nor U9778 (N_9778,N_9688,N_9623);
or U9779 (N_9779,N_9191,N_9054);
and U9780 (N_9780,N_9295,N_9312);
and U9781 (N_9781,N_9421,N_9085);
or U9782 (N_9782,N_9550,N_9448);
and U9783 (N_9783,N_9584,N_9329);
or U9784 (N_9784,N_9086,N_9041);
and U9785 (N_9785,N_9423,N_9200);
xnor U9786 (N_9786,N_9451,N_9173);
nor U9787 (N_9787,N_9466,N_9327);
and U9788 (N_9788,N_9209,N_9567);
and U9789 (N_9789,N_9478,N_9298);
or U9790 (N_9790,N_9174,N_9205);
nand U9791 (N_9791,N_9570,N_9005);
nand U9792 (N_9792,N_9438,N_9605);
and U9793 (N_9793,N_9045,N_9016);
or U9794 (N_9794,N_9720,N_9111);
or U9795 (N_9795,N_9161,N_9020);
nor U9796 (N_9796,N_9287,N_9202);
and U9797 (N_9797,N_9227,N_9105);
or U9798 (N_9798,N_9695,N_9263);
nand U9799 (N_9799,N_9530,N_9164);
or U9800 (N_9800,N_9301,N_9386);
or U9801 (N_9801,N_9163,N_9709);
nor U9802 (N_9802,N_9145,N_9344);
xor U9803 (N_9803,N_9741,N_9744);
xor U9804 (N_9804,N_9634,N_9619);
or U9805 (N_9805,N_9141,N_9216);
xor U9806 (N_9806,N_9406,N_9158);
nor U9807 (N_9807,N_9618,N_9408);
nand U9808 (N_9808,N_9282,N_9560);
or U9809 (N_9809,N_9600,N_9034);
xor U9810 (N_9810,N_9474,N_9497);
xor U9811 (N_9811,N_9070,N_9153);
nor U9812 (N_9812,N_9026,N_9711);
or U9813 (N_9813,N_9160,N_9731);
nand U9814 (N_9814,N_9713,N_9625);
and U9815 (N_9815,N_9444,N_9491);
or U9816 (N_9816,N_9674,N_9452);
xnor U9817 (N_9817,N_9283,N_9612);
nor U9818 (N_9818,N_9407,N_9427);
nor U9819 (N_9819,N_9396,N_9660);
xor U9820 (N_9820,N_9302,N_9255);
nor U9821 (N_9821,N_9399,N_9522);
nor U9822 (N_9822,N_9663,N_9390);
nand U9823 (N_9823,N_9019,N_9628);
and U9824 (N_9824,N_9220,N_9653);
and U9825 (N_9825,N_9035,N_9704);
xor U9826 (N_9826,N_9519,N_9288);
and U9827 (N_9827,N_9229,N_9735);
nand U9828 (N_9828,N_9006,N_9369);
nor U9829 (N_9829,N_9151,N_9102);
and U9830 (N_9830,N_9575,N_9120);
xnor U9831 (N_9831,N_9052,N_9487);
or U9832 (N_9832,N_9595,N_9549);
and U9833 (N_9833,N_9314,N_9637);
or U9834 (N_9834,N_9449,N_9539);
or U9835 (N_9835,N_9579,N_9620);
nand U9836 (N_9836,N_9694,N_9360);
or U9837 (N_9837,N_9658,N_9087);
nor U9838 (N_9838,N_9385,N_9568);
and U9839 (N_9839,N_9503,N_9032);
xor U9840 (N_9840,N_9395,N_9079);
nand U9841 (N_9841,N_9511,N_9011);
or U9842 (N_9842,N_9296,N_9398);
or U9843 (N_9843,N_9518,N_9093);
nand U9844 (N_9844,N_9024,N_9632);
nand U9845 (N_9845,N_9101,N_9044);
nand U9846 (N_9846,N_9543,N_9745);
or U9847 (N_9847,N_9557,N_9372);
xor U9848 (N_9848,N_9129,N_9236);
nor U9849 (N_9849,N_9544,N_9669);
and U9850 (N_9850,N_9462,N_9603);
nor U9851 (N_9851,N_9426,N_9534);
xnor U9852 (N_9852,N_9000,N_9180);
xnor U9853 (N_9853,N_9477,N_9003);
nor U9854 (N_9854,N_9089,N_9152);
xnor U9855 (N_9855,N_9128,N_9340);
nand U9856 (N_9856,N_9662,N_9521);
xor U9857 (N_9857,N_9197,N_9416);
nor U9858 (N_9858,N_9496,N_9747);
or U9859 (N_9859,N_9276,N_9702);
and U9860 (N_9860,N_9433,N_9555);
nand U9861 (N_9861,N_9265,N_9370);
and U9862 (N_9862,N_9631,N_9068);
nor U9863 (N_9863,N_9722,N_9194);
and U9864 (N_9864,N_9649,N_9640);
or U9865 (N_9865,N_9073,N_9053);
or U9866 (N_9866,N_9381,N_9090);
or U9867 (N_9867,N_9667,N_9589);
nor U9868 (N_9868,N_9689,N_9238);
or U9869 (N_9869,N_9065,N_9150);
nand U9870 (N_9870,N_9592,N_9393);
nand U9871 (N_9871,N_9267,N_9237);
nand U9872 (N_9872,N_9107,N_9001);
xor U9873 (N_9873,N_9315,N_9351);
nand U9874 (N_9874,N_9368,N_9257);
xor U9875 (N_9875,N_9707,N_9683);
and U9876 (N_9876,N_9311,N_9414);
nor U9877 (N_9877,N_9275,N_9323);
nor U9878 (N_9878,N_9643,N_9703);
xnor U9879 (N_9879,N_9384,N_9055);
xnor U9880 (N_9880,N_9739,N_9213);
xnor U9881 (N_9881,N_9099,N_9551);
xor U9882 (N_9882,N_9064,N_9293);
nor U9883 (N_9883,N_9217,N_9590);
nand U9884 (N_9884,N_9383,N_9533);
xor U9885 (N_9885,N_9428,N_9565);
nand U9886 (N_9886,N_9553,N_9712);
xnor U9887 (N_9887,N_9463,N_9030);
or U9888 (N_9888,N_9182,N_9388);
xnor U9889 (N_9889,N_9455,N_9014);
nand U9890 (N_9890,N_9526,N_9292);
nor U9891 (N_9891,N_9131,N_9425);
and U9892 (N_9892,N_9733,N_9728);
nor U9893 (N_9893,N_9624,N_9710);
and U9894 (N_9894,N_9280,N_9028);
and U9895 (N_9895,N_9246,N_9685);
nand U9896 (N_9896,N_9169,N_9743);
or U9897 (N_9897,N_9515,N_9008);
nand U9898 (N_9898,N_9661,N_9725);
and U9899 (N_9899,N_9571,N_9442);
or U9900 (N_9900,N_9548,N_9337);
nor U9901 (N_9901,N_9686,N_9488);
xor U9902 (N_9902,N_9270,N_9472);
xor U9903 (N_9903,N_9690,N_9583);
or U9904 (N_9904,N_9144,N_9110);
xnor U9905 (N_9905,N_9601,N_9475);
and U9906 (N_9906,N_9412,N_9483);
and U9907 (N_9907,N_9240,N_9531);
or U9908 (N_9908,N_9096,N_9687);
xnor U9909 (N_9909,N_9436,N_9214);
and U9910 (N_9910,N_9338,N_9588);
xor U9911 (N_9911,N_9010,N_9042);
or U9912 (N_9912,N_9582,N_9123);
xnor U9913 (N_9913,N_9742,N_9154);
nor U9914 (N_9914,N_9080,N_9394);
and U9915 (N_9915,N_9546,N_9616);
or U9916 (N_9916,N_9207,N_9211);
nor U9917 (N_9917,N_9479,N_9635);
nor U9918 (N_9918,N_9527,N_9535);
or U9919 (N_9919,N_9577,N_9289);
nor U9920 (N_9920,N_9192,N_9274);
xnor U9921 (N_9921,N_9389,N_9591);
xnor U9922 (N_9922,N_9437,N_9133);
nor U9923 (N_9923,N_9482,N_9215);
and U9924 (N_9924,N_9524,N_9597);
and U9925 (N_9925,N_9380,N_9130);
nor U9926 (N_9926,N_9541,N_9061);
nand U9927 (N_9927,N_9094,N_9617);
or U9928 (N_9928,N_9031,N_9226);
nand U9929 (N_9929,N_9325,N_9645);
or U9930 (N_9930,N_9221,N_9199);
and U9931 (N_9931,N_9058,N_9506);
or U9932 (N_9932,N_9179,N_9513);
xor U9933 (N_9933,N_9602,N_9740);
and U9934 (N_9934,N_9611,N_9063);
nor U9935 (N_9935,N_9738,N_9050);
and U9936 (N_9936,N_9195,N_9168);
nand U9937 (N_9937,N_9523,N_9185);
nor U9938 (N_9938,N_9346,N_9505);
nor U9939 (N_9939,N_9470,N_9454);
and U9940 (N_9940,N_9594,N_9260);
xnor U9941 (N_9941,N_9556,N_9664);
xnor U9942 (N_9942,N_9043,N_9009);
nor U9943 (N_9943,N_9212,N_9458);
or U9944 (N_9944,N_9581,N_9447);
xnor U9945 (N_9945,N_9023,N_9259);
nand U9946 (N_9946,N_9574,N_9071);
or U9947 (N_9947,N_9290,N_9156);
and U9948 (N_9948,N_9748,N_9465);
or U9949 (N_9949,N_9262,N_9029);
and U9950 (N_9950,N_9604,N_9228);
nor U9951 (N_9951,N_9004,N_9459);
xnor U9952 (N_9952,N_9230,N_9648);
and U9953 (N_9953,N_9036,N_9598);
nand U9954 (N_9954,N_9573,N_9593);
or U9955 (N_9955,N_9432,N_9335);
or U9956 (N_9956,N_9729,N_9317);
and U9957 (N_9957,N_9272,N_9308);
nand U9958 (N_9958,N_9322,N_9668);
or U9959 (N_9959,N_9307,N_9500);
nand U9960 (N_9960,N_9445,N_9424);
nand U9961 (N_9961,N_9318,N_9439);
nor U9962 (N_9962,N_9507,N_9134);
and U9963 (N_9963,N_9177,N_9092);
xor U9964 (N_9964,N_9514,N_9193);
xor U9965 (N_9965,N_9392,N_9320);
xor U9966 (N_9966,N_9328,N_9365);
xor U9967 (N_9967,N_9297,N_9723);
nor U9968 (N_9968,N_9253,N_9136);
nor U9969 (N_9969,N_9264,N_9721);
nand U9970 (N_9970,N_9489,N_9699);
nand U9971 (N_9971,N_9015,N_9309);
xnor U9972 (N_9972,N_9510,N_9037);
xor U9973 (N_9973,N_9642,N_9244);
and U9974 (N_9974,N_9430,N_9103);
xor U9975 (N_9975,N_9547,N_9204);
or U9976 (N_9976,N_9453,N_9420);
and U9977 (N_9977,N_9501,N_9114);
nand U9978 (N_9978,N_9017,N_9724);
or U9979 (N_9979,N_9646,N_9609);
nand U9980 (N_9980,N_9040,N_9401);
nor U9981 (N_9981,N_9355,N_9165);
nor U9982 (N_9982,N_9749,N_9665);
nand U9983 (N_9983,N_9188,N_9266);
nand U9984 (N_9984,N_9210,N_9615);
and U9985 (N_9985,N_9224,N_9486);
nor U9986 (N_9986,N_9671,N_9159);
nor U9987 (N_9987,N_9715,N_9657);
nor U9988 (N_9988,N_9502,N_9157);
nor U9989 (N_9989,N_9206,N_9135);
or U9990 (N_9990,N_9147,N_9529);
or U9991 (N_9991,N_9341,N_9285);
and U9992 (N_9992,N_9726,N_9537);
nand U9993 (N_9993,N_9559,N_9231);
and U9994 (N_9994,N_9176,N_9261);
or U9995 (N_9995,N_9198,N_9700);
nand U9996 (N_9996,N_9100,N_9512);
xor U9997 (N_9997,N_9587,N_9673);
xor U9998 (N_9998,N_9576,N_9409);
or U9999 (N_9999,N_9562,N_9627);
nand U10000 (N_10000,N_9464,N_9077);
nand U10001 (N_10001,N_9356,N_9540);
or U10002 (N_10002,N_9116,N_9132);
or U10003 (N_10003,N_9701,N_9115);
and U10004 (N_10004,N_9361,N_9354);
nand U10005 (N_10005,N_9644,N_9415);
or U10006 (N_10006,N_9347,N_9278);
nor U10007 (N_10007,N_9139,N_9038);
nor U10008 (N_10008,N_9059,N_9048);
and U10009 (N_10009,N_9607,N_9638);
nor U10010 (N_10010,N_9084,N_9018);
nor U10011 (N_10011,N_9303,N_9332);
nand U10012 (N_10012,N_9680,N_9599);
nor U10013 (N_10013,N_9652,N_9124);
or U10014 (N_10014,N_9251,N_9666);
or U10015 (N_10015,N_9316,N_9647);
nor U10016 (N_10016,N_9078,N_9350);
nor U10017 (N_10017,N_9708,N_9499);
xnor U10018 (N_10018,N_9580,N_9650);
nor U10019 (N_10019,N_9352,N_9357);
and U10020 (N_10020,N_9277,N_9268);
and U10021 (N_10021,N_9299,N_9419);
or U10022 (N_10022,N_9239,N_9256);
xnor U10023 (N_10023,N_9732,N_9007);
xnor U10024 (N_10024,N_9378,N_9201);
xor U10025 (N_10025,N_9046,N_9440);
nand U10026 (N_10026,N_9002,N_9162);
xnor U10027 (N_10027,N_9586,N_9121);
xor U10028 (N_10028,N_9626,N_9183);
and U10029 (N_10029,N_9564,N_9450);
nand U10030 (N_10030,N_9681,N_9072);
nand U10031 (N_10031,N_9025,N_9118);
xor U10032 (N_10032,N_9339,N_9076);
nand U10033 (N_10033,N_9727,N_9208);
nor U10034 (N_10034,N_9693,N_9359);
xnor U10035 (N_10035,N_9656,N_9149);
and U10036 (N_10036,N_9528,N_9374);
xor U10037 (N_10037,N_9717,N_9167);
nor U10038 (N_10038,N_9181,N_9678);
and U10039 (N_10039,N_9734,N_9258);
nor U10040 (N_10040,N_9140,N_9641);
nand U10041 (N_10041,N_9186,N_9532);
xor U10042 (N_10042,N_9387,N_9273);
xor U10043 (N_10043,N_9391,N_9047);
nor U10044 (N_10044,N_9364,N_9682);
nand U10045 (N_10045,N_9232,N_9698);
nand U10046 (N_10046,N_9166,N_9730);
nor U10047 (N_10047,N_9021,N_9286);
or U10048 (N_10048,N_9517,N_9271);
or U10049 (N_10049,N_9614,N_9108);
xor U10050 (N_10050,N_9233,N_9027);
nand U10051 (N_10051,N_9069,N_9516);
nand U10052 (N_10052,N_9371,N_9379);
and U10053 (N_10053,N_9471,N_9190);
nand U10054 (N_10054,N_9235,N_9241);
and U10055 (N_10055,N_9429,N_9219);
or U10056 (N_10056,N_9676,N_9305);
or U10057 (N_10057,N_9692,N_9525);
nor U10058 (N_10058,N_9119,N_9654);
or U10059 (N_10059,N_9608,N_9106);
and U10060 (N_10060,N_9400,N_9446);
nor U10061 (N_10061,N_9095,N_9178);
nand U10062 (N_10062,N_9485,N_9057);
or U10063 (N_10063,N_9675,N_9218);
nor U10064 (N_10064,N_9397,N_9367);
xor U10065 (N_10065,N_9081,N_9254);
nand U10066 (N_10066,N_9622,N_9659);
xor U10067 (N_10067,N_9706,N_9066);
nand U10068 (N_10068,N_9321,N_9075);
nand U10069 (N_10069,N_9405,N_9435);
and U10070 (N_10070,N_9098,N_9171);
and U10071 (N_10071,N_9249,N_9284);
and U10072 (N_10072,N_9460,N_9334);
or U10073 (N_10073,N_9113,N_9247);
xor U10074 (N_10074,N_9248,N_9596);
nor U10075 (N_10075,N_9691,N_9376);
or U10076 (N_10076,N_9697,N_9326);
nand U10077 (N_10077,N_9033,N_9039);
or U10078 (N_10078,N_9473,N_9300);
nor U10079 (N_10079,N_9672,N_9480);
xor U10080 (N_10080,N_9696,N_9558);
or U10081 (N_10081,N_9677,N_9633);
or U10082 (N_10082,N_9552,N_9651);
xnor U10083 (N_10083,N_9469,N_9336);
nor U10084 (N_10084,N_9049,N_9225);
or U10085 (N_10085,N_9508,N_9067);
xnor U10086 (N_10086,N_9012,N_9083);
and U10087 (N_10087,N_9013,N_9062);
nand U10088 (N_10088,N_9250,N_9610);
xnor U10089 (N_10089,N_9146,N_9578);
and U10090 (N_10090,N_9082,N_9520);
xor U10091 (N_10091,N_9056,N_9422);
and U10092 (N_10092,N_9324,N_9137);
nand U10093 (N_10093,N_9281,N_9117);
nand U10094 (N_10094,N_9331,N_9719);
xor U10095 (N_10095,N_9373,N_9184);
nor U10096 (N_10096,N_9736,N_9172);
xnor U10097 (N_10097,N_9353,N_9223);
or U10098 (N_10098,N_9679,N_9538);
nand U10099 (N_10099,N_9269,N_9718);
or U10100 (N_10100,N_9621,N_9493);
xnor U10101 (N_10101,N_9498,N_9382);
or U10102 (N_10102,N_9630,N_9203);
xnor U10103 (N_10103,N_9705,N_9125);
and U10104 (N_10104,N_9434,N_9126);
nand U10105 (N_10105,N_9468,N_9418);
xor U10106 (N_10106,N_9492,N_9342);
and U10107 (N_10107,N_9060,N_9148);
or U10108 (N_10108,N_9410,N_9542);
or U10109 (N_10109,N_9306,N_9569);
nor U10110 (N_10110,N_9234,N_9175);
xor U10111 (N_10111,N_9242,N_9737);
or U10112 (N_10112,N_9504,N_9467);
or U10113 (N_10113,N_9222,N_9279);
or U10114 (N_10114,N_9684,N_9563);
and U10115 (N_10115,N_9345,N_9476);
nor U10116 (N_10116,N_9572,N_9348);
nand U10117 (N_10117,N_9243,N_9484);
and U10118 (N_10118,N_9456,N_9363);
nand U10119 (N_10119,N_9746,N_9291);
and U10120 (N_10120,N_9112,N_9411);
nand U10121 (N_10121,N_9716,N_9330);
nand U10122 (N_10122,N_9189,N_9417);
nor U10123 (N_10123,N_9187,N_9402);
and U10124 (N_10124,N_9377,N_9143);
xor U10125 (N_10125,N_9046,N_9024);
nand U10126 (N_10126,N_9140,N_9285);
and U10127 (N_10127,N_9728,N_9042);
nand U10128 (N_10128,N_9573,N_9516);
and U10129 (N_10129,N_9267,N_9600);
xnor U10130 (N_10130,N_9111,N_9733);
nor U10131 (N_10131,N_9029,N_9313);
or U10132 (N_10132,N_9675,N_9672);
or U10133 (N_10133,N_9727,N_9486);
and U10134 (N_10134,N_9473,N_9578);
or U10135 (N_10135,N_9354,N_9526);
and U10136 (N_10136,N_9299,N_9669);
and U10137 (N_10137,N_9029,N_9669);
nor U10138 (N_10138,N_9630,N_9034);
or U10139 (N_10139,N_9177,N_9627);
nor U10140 (N_10140,N_9082,N_9154);
nor U10141 (N_10141,N_9679,N_9029);
nor U10142 (N_10142,N_9567,N_9428);
and U10143 (N_10143,N_9233,N_9077);
nor U10144 (N_10144,N_9723,N_9703);
and U10145 (N_10145,N_9599,N_9708);
nor U10146 (N_10146,N_9625,N_9633);
nor U10147 (N_10147,N_9008,N_9463);
nand U10148 (N_10148,N_9196,N_9061);
xor U10149 (N_10149,N_9497,N_9317);
nand U10150 (N_10150,N_9057,N_9051);
nor U10151 (N_10151,N_9480,N_9225);
or U10152 (N_10152,N_9079,N_9320);
nor U10153 (N_10153,N_9132,N_9626);
xnor U10154 (N_10154,N_9459,N_9472);
and U10155 (N_10155,N_9064,N_9421);
nand U10156 (N_10156,N_9550,N_9144);
nand U10157 (N_10157,N_9631,N_9495);
and U10158 (N_10158,N_9741,N_9715);
or U10159 (N_10159,N_9130,N_9630);
nand U10160 (N_10160,N_9730,N_9281);
or U10161 (N_10161,N_9308,N_9021);
nor U10162 (N_10162,N_9338,N_9555);
xor U10163 (N_10163,N_9121,N_9349);
nand U10164 (N_10164,N_9706,N_9698);
and U10165 (N_10165,N_9021,N_9064);
xnor U10166 (N_10166,N_9104,N_9716);
nor U10167 (N_10167,N_9189,N_9149);
xnor U10168 (N_10168,N_9261,N_9318);
nand U10169 (N_10169,N_9347,N_9025);
xnor U10170 (N_10170,N_9364,N_9125);
nand U10171 (N_10171,N_9658,N_9609);
nand U10172 (N_10172,N_9422,N_9523);
and U10173 (N_10173,N_9704,N_9265);
nor U10174 (N_10174,N_9243,N_9137);
nor U10175 (N_10175,N_9166,N_9408);
and U10176 (N_10176,N_9423,N_9746);
nor U10177 (N_10177,N_9411,N_9156);
or U10178 (N_10178,N_9442,N_9597);
nor U10179 (N_10179,N_9140,N_9357);
or U10180 (N_10180,N_9224,N_9228);
or U10181 (N_10181,N_9088,N_9475);
nor U10182 (N_10182,N_9251,N_9288);
xnor U10183 (N_10183,N_9017,N_9700);
nand U10184 (N_10184,N_9498,N_9108);
or U10185 (N_10185,N_9115,N_9246);
and U10186 (N_10186,N_9302,N_9361);
nand U10187 (N_10187,N_9187,N_9596);
nor U10188 (N_10188,N_9303,N_9312);
nand U10189 (N_10189,N_9214,N_9112);
nor U10190 (N_10190,N_9365,N_9563);
nor U10191 (N_10191,N_9131,N_9580);
and U10192 (N_10192,N_9679,N_9484);
or U10193 (N_10193,N_9604,N_9101);
nor U10194 (N_10194,N_9609,N_9589);
and U10195 (N_10195,N_9149,N_9507);
nand U10196 (N_10196,N_9067,N_9367);
and U10197 (N_10197,N_9556,N_9715);
and U10198 (N_10198,N_9081,N_9130);
or U10199 (N_10199,N_9408,N_9470);
nor U10200 (N_10200,N_9453,N_9486);
xnor U10201 (N_10201,N_9109,N_9666);
xnor U10202 (N_10202,N_9523,N_9087);
xor U10203 (N_10203,N_9633,N_9216);
nand U10204 (N_10204,N_9279,N_9401);
xnor U10205 (N_10205,N_9340,N_9687);
xnor U10206 (N_10206,N_9552,N_9362);
or U10207 (N_10207,N_9251,N_9726);
nand U10208 (N_10208,N_9698,N_9440);
and U10209 (N_10209,N_9237,N_9611);
nand U10210 (N_10210,N_9546,N_9558);
nor U10211 (N_10211,N_9151,N_9043);
or U10212 (N_10212,N_9582,N_9663);
nand U10213 (N_10213,N_9478,N_9251);
nor U10214 (N_10214,N_9044,N_9627);
and U10215 (N_10215,N_9008,N_9095);
nand U10216 (N_10216,N_9334,N_9277);
xor U10217 (N_10217,N_9212,N_9711);
xnor U10218 (N_10218,N_9110,N_9515);
or U10219 (N_10219,N_9413,N_9472);
nor U10220 (N_10220,N_9143,N_9057);
xnor U10221 (N_10221,N_9526,N_9325);
nor U10222 (N_10222,N_9191,N_9405);
xor U10223 (N_10223,N_9227,N_9526);
or U10224 (N_10224,N_9238,N_9472);
xnor U10225 (N_10225,N_9336,N_9086);
and U10226 (N_10226,N_9711,N_9110);
or U10227 (N_10227,N_9276,N_9486);
nand U10228 (N_10228,N_9500,N_9744);
nor U10229 (N_10229,N_9493,N_9012);
nor U10230 (N_10230,N_9060,N_9297);
nor U10231 (N_10231,N_9319,N_9555);
nand U10232 (N_10232,N_9497,N_9529);
and U10233 (N_10233,N_9732,N_9039);
or U10234 (N_10234,N_9343,N_9711);
nand U10235 (N_10235,N_9319,N_9158);
nor U10236 (N_10236,N_9268,N_9341);
or U10237 (N_10237,N_9301,N_9747);
or U10238 (N_10238,N_9296,N_9525);
or U10239 (N_10239,N_9679,N_9537);
and U10240 (N_10240,N_9224,N_9672);
xor U10241 (N_10241,N_9502,N_9161);
or U10242 (N_10242,N_9225,N_9327);
or U10243 (N_10243,N_9663,N_9350);
and U10244 (N_10244,N_9480,N_9275);
and U10245 (N_10245,N_9251,N_9682);
xnor U10246 (N_10246,N_9358,N_9588);
and U10247 (N_10247,N_9146,N_9496);
or U10248 (N_10248,N_9087,N_9540);
or U10249 (N_10249,N_9407,N_9585);
nor U10250 (N_10250,N_9324,N_9655);
and U10251 (N_10251,N_9732,N_9415);
nor U10252 (N_10252,N_9148,N_9033);
nor U10253 (N_10253,N_9637,N_9316);
and U10254 (N_10254,N_9440,N_9696);
xor U10255 (N_10255,N_9713,N_9497);
nor U10256 (N_10256,N_9393,N_9524);
and U10257 (N_10257,N_9695,N_9499);
xor U10258 (N_10258,N_9372,N_9348);
xor U10259 (N_10259,N_9558,N_9384);
xnor U10260 (N_10260,N_9175,N_9210);
xnor U10261 (N_10261,N_9564,N_9380);
nor U10262 (N_10262,N_9703,N_9043);
nor U10263 (N_10263,N_9114,N_9161);
xor U10264 (N_10264,N_9619,N_9512);
nand U10265 (N_10265,N_9144,N_9497);
xor U10266 (N_10266,N_9035,N_9229);
xnor U10267 (N_10267,N_9158,N_9053);
nand U10268 (N_10268,N_9033,N_9098);
or U10269 (N_10269,N_9594,N_9524);
or U10270 (N_10270,N_9231,N_9672);
nor U10271 (N_10271,N_9407,N_9403);
xor U10272 (N_10272,N_9053,N_9023);
nor U10273 (N_10273,N_9594,N_9230);
or U10274 (N_10274,N_9413,N_9303);
xor U10275 (N_10275,N_9210,N_9478);
nand U10276 (N_10276,N_9270,N_9436);
xnor U10277 (N_10277,N_9166,N_9679);
and U10278 (N_10278,N_9101,N_9411);
xnor U10279 (N_10279,N_9520,N_9068);
nand U10280 (N_10280,N_9594,N_9652);
nor U10281 (N_10281,N_9121,N_9078);
xnor U10282 (N_10282,N_9320,N_9032);
or U10283 (N_10283,N_9234,N_9273);
and U10284 (N_10284,N_9414,N_9253);
and U10285 (N_10285,N_9685,N_9095);
or U10286 (N_10286,N_9627,N_9422);
or U10287 (N_10287,N_9140,N_9043);
xnor U10288 (N_10288,N_9321,N_9329);
and U10289 (N_10289,N_9584,N_9245);
nor U10290 (N_10290,N_9588,N_9126);
nor U10291 (N_10291,N_9434,N_9436);
and U10292 (N_10292,N_9682,N_9456);
xnor U10293 (N_10293,N_9431,N_9232);
xnor U10294 (N_10294,N_9147,N_9131);
and U10295 (N_10295,N_9204,N_9202);
xor U10296 (N_10296,N_9199,N_9361);
nand U10297 (N_10297,N_9564,N_9086);
and U10298 (N_10298,N_9515,N_9508);
and U10299 (N_10299,N_9266,N_9504);
or U10300 (N_10300,N_9096,N_9092);
and U10301 (N_10301,N_9671,N_9584);
xor U10302 (N_10302,N_9204,N_9646);
xor U10303 (N_10303,N_9066,N_9639);
or U10304 (N_10304,N_9664,N_9617);
nor U10305 (N_10305,N_9113,N_9117);
or U10306 (N_10306,N_9200,N_9637);
nand U10307 (N_10307,N_9130,N_9133);
and U10308 (N_10308,N_9712,N_9455);
and U10309 (N_10309,N_9456,N_9182);
or U10310 (N_10310,N_9368,N_9469);
nand U10311 (N_10311,N_9671,N_9536);
nand U10312 (N_10312,N_9329,N_9341);
xor U10313 (N_10313,N_9337,N_9411);
or U10314 (N_10314,N_9499,N_9429);
nand U10315 (N_10315,N_9037,N_9079);
or U10316 (N_10316,N_9109,N_9472);
nand U10317 (N_10317,N_9623,N_9092);
or U10318 (N_10318,N_9307,N_9567);
or U10319 (N_10319,N_9493,N_9031);
nor U10320 (N_10320,N_9474,N_9399);
nor U10321 (N_10321,N_9537,N_9227);
and U10322 (N_10322,N_9514,N_9410);
and U10323 (N_10323,N_9510,N_9105);
or U10324 (N_10324,N_9270,N_9144);
or U10325 (N_10325,N_9661,N_9501);
xor U10326 (N_10326,N_9643,N_9613);
or U10327 (N_10327,N_9683,N_9454);
or U10328 (N_10328,N_9104,N_9130);
nand U10329 (N_10329,N_9353,N_9522);
or U10330 (N_10330,N_9428,N_9448);
and U10331 (N_10331,N_9397,N_9004);
xnor U10332 (N_10332,N_9527,N_9208);
nor U10333 (N_10333,N_9094,N_9076);
and U10334 (N_10334,N_9644,N_9066);
or U10335 (N_10335,N_9664,N_9279);
nor U10336 (N_10336,N_9354,N_9535);
and U10337 (N_10337,N_9451,N_9312);
or U10338 (N_10338,N_9277,N_9165);
and U10339 (N_10339,N_9225,N_9160);
or U10340 (N_10340,N_9018,N_9349);
or U10341 (N_10341,N_9324,N_9014);
xor U10342 (N_10342,N_9466,N_9233);
xnor U10343 (N_10343,N_9486,N_9650);
or U10344 (N_10344,N_9223,N_9007);
and U10345 (N_10345,N_9476,N_9115);
xor U10346 (N_10346,N_9617,N_9546);
and U10347 (N_10347,N_9332,N_9360);
and U10348 (N_10348,N_9004,N_9503);
or U10349 (N_10349,N_9626,N_9275);
or U10350 (N_10350,N_9316,N_9282);
nor U10351 (N_10351,N_9359,N_9026);
nand U10352 (N_10352,N_9567,N_9694);
or U10353 (N_10353,N_9105,N_9260);
and U10354 (N_10354,N_9718,N_9722);
nor U10355 (N_10355,N_9725,N_9208);
xnor U10356 (N_10356,N_9557,N_9639);
nor U10357 (N_10357,N_9178,N_9021);
or U10358 (N_10358,N_9677,N_9074);
and U10359 (N_10359,N_9510,N_9202);
nor U10360 (N_10360,N_9265,N_9063);
or U10361 (N_10361,N_9433,N_9441);
xnor U10362 (N_10362,N_9678,N_9564);
nand U10363 (N_10363,N_9717,N_9725);
and U10364 (N_10364,N_9307,N_9209);
and U10365 (N_10365,N_9375,N_9741);
nor U10366 (N_10366,N_9104,N_9354);
and U10367 (N_10367,N_9615,N_9520);
and U10368 (N_10368,N_9456,N_9641);
nor U10369 (N_10369,N_9089,N_9738);
nor U10370 (N_10370,N_9161,N_9432);
nand U10371 (N_10371,N_9525,N_9362);
and U10372 (N_10372,N_9416,N_9188);
xnor U10373 (N_10373,N_9679,N_9009);
nand U10374 (N_10374,N_9650,N_9318);
nand U10375 (N_10375,N_9310,N_9626);
or U10376 (N_10376,N_9671,N_9618);
nor U10377 (N_10377,N_9408,N_9205);
nand U10378 (N_10378,N_9708,N_9735);
xor U10379 (N_10379,N_9659,N_9278);
or U10380 (N_10380,N_9015,N_9729);
nand U10381 (N_10381,N_9491,N_9239);
nand U10382 (N_10382,N_9385,N_9311);
or U10383 (N_10383,N_9323,N_9260);
nand U10384 (N_10384,N_9440,N_9727);
or U10385 (N_10385,N_9471,N_9010);
xor U10386 (N_10386,N_9458,N_9629);
and U10387 (N_10387,N_9127,N_9360);
and U10388 (N_10388,N_9623,N_9536);
nand U10389 (N_10389,N_9281,N_9516);
nand U10390 (N_10390,N_9370,N_9500);
nor U10391 (N_10391,N_9164,N_9437);
nand U10392 (N_10392,N_9229,N_9005);
xor U10393 (N_10393,N_9444,N_9725);
and U10394 (N_10394,N_9250,N_9725);
and U10395 (N_10395,N_9033,N_9261);
and U10396 (N_10396,N_9330,N_9023);
and U10397 (N_10397,N_9009,N_9693);
nand U10398 (N_10398,N_9296,N_9736);
nand U10399 (N_10399,N_9166,N_9420);
nor U10400 (N_10400,N_9043,N_9164);
or U10401 (N_10401,N_9092,N_9525);
nor U10402 (N_10402,N_9177,N_9664);
or U10403 (N_10403,N_9498,N_9039);
or U10404 (N_10404,N_9704,N_9639);
or U10405 (N_10405,N_9036,N_9498);
nor U10406 (N_10406,N_9620,N_9105);
nand U10407 (N_10407,N_9344,N_9690);
and U10408 (N_10408,N_9557,N_9554);
nand U10409 (N_10409,N_9609,N_9109);
or U10410 (N_10410,N_9616,N_9271);
and U10411 (N_10411,N_9520,N_9203);
and U10412 (N_10412,N_9210,N_9574);
or U10413 (N_10413,N_9043,N_9144);
nand U10414 (N_10414,N_9347,N_9236);
nor U10415 (N_10415,N_9337,N_9154);
or U10416 (N_10416,N_9227,N_9304);
and U10417 (N_10417,N_9015,N_9143);
xnor U10418 (N_10418,N_9129,N_9217);
xnor U10419 (N_10419,N_9359,N_9031);
nand U10420 (N_10420,N_9625,N_9482);
xnor U10421 (N_10421,N_9386,N_9495);
xnor U10422 (N_10422,N_9546,N_9119);
xnor U10423 (N_10423,N_9090,N_9748);
nor U10424 (N_10424,N_9279,N_9189);
or U10425 (N_10425,N_9679,N_9032);
and U10426 (N_10426,N_9256,N_9090);
nor U10427 (N_10427,N_9480,N_9562);
nand U10428 (N_10428,N_9548,N_9274);
nand U10429 (N_10429,N_9330,N_9697);
xnor U10430 (N_10430,N_9707,N_9445);
xor U10431 (N_10431,N_9096,N_9154);
or U10432 (N_10432,N_9147,N_9019);
nand U10433 (N_10433,N_9546,N_9556);
nand U10434 (N_10434,N_9701,N_9251);
nor U10435 (N_10435,N_9504,N_9005);
and U10436 (N_10436,N_9258,N_9030);
or U10437 (N_10437,N_9042,N_9691);
xor U10438 (N_10438,N_9262,N_9422);
and U10439 (N_10439,N_9464,N_9250);
nor U10440 (N_10440,N_9476,N_9468);
nand U10441 (N_10441,N_9342,N_9023);
nand U10442 (N_10442,N_9196,N_9314);
xnor U10443 (N_10443,N_9162,N_9748);
nor U10444 (N_10444,N_9373,N_9257);
and U10445 (N_10445,N_9141,N_9569);
nand U10446 (N_10446,N_9045,N_9308);
nand U10447 (N_10447,N_9561,N_9363);
xor U10448 (N_10448,N_9431,N_9255);
xnor U10449 (N_10449,N_9271,N_9501);
nor U10450 (N_10450,N_9019,N_9429);
xnor U10451 (N_10451,N_9594,N_9100);
or U10452 (N_10452,N_9547,N_9323);
or U10453 (N_10453,N_9691,N_9723);
xor U10454 (N_10454,N_9379,N_9450);
xor U10455 (N_10455,N_9120,N_9101);
or U10456 (N_10456,N_9410,N_9043);
nand U10457 (N_10457,N_9320,N_9039);
nor U10458 (N_10458,N_9690,N_9743);
or U10459 (N_10459,N_9349,N_9088);
nand U10460 (N_10460,N_9572,N_9413);
nor U10461 (N_10461,N_9284,N_9236);
or U10462 (N_10462,N_9426,N_9455);
nand U10463 (N_10463,N_9481,N_9203);
xor U10464 (N_10464,N_9170,N_9516);
nand U10465 (N_10465,N_9498,N_9208);
nor U10466 (N_10466,N_9015,N_9254);
or U10467 (N_10467,N_9533,N_9252);
or U10468 (N_10468,N_9008,N_9637);
or U10469 (N_10469,N_9707,N_9262);
nand U10470 (N_10470,N_9214,N_9212);
nand U10471 (N_10471,N_9242,N_9647);
or U10472 (N_10472,N_9011,N_9568);
nand U10473 (N_10473,N_9729,N_9699);
nor U10474 (N_10474,N_9042,N_9666);
and U10475 (N_10475,N_9540,N_9253);
nor U10476 (N_10476,N_9217,N_9176);
xnor U10477 (N_10477,N_9442,N_9120);
nor U10478 (N_10478,N_9457,N_9551);
and U10479 (N_10479,N_9550,N_9411);
nand U10480 (N_10480,N_9036,N_9631);
xor U10481 (N_10481,N_9365,N_9437);
and U10482 (N_10482,N_9002,N_9355);
xor U10483 (N_10483,N_9266,N_9032);
or U10484 (N_10484,N_9269,N_9588);
and U10485 (N_10485,N_9636,N_9157);
and U10486 (N_10486,N_9684,N_9186);
nor U10487 (N_10487,N_9558,N_9189);
nor U10488 (N_10488,N_9633,N_9061);
or U10489 (N_10489,N_9635,N_9053);
xor U10490 (N_10490,N_9690,N_9174);
nand U10491 (N_10491,N_9006,N_9478);
and U10492 (N_10492,N_9212,N_9194);
xor U10493 (N_10493,N_9749,N_9569);
nand U10494 (N_10494,N_9300,N_9507);
nor U10495 (N_10495,N_9492,N_9083);
xnor U10496 (N_10496,N_9297,N_9693);
and U10497 (N_10497,N_9582,N_9246);
xor U10498 (N_10498,N_9129,N_9598);
and U10499 (N_10499,N_9568,N_9544);
or U10500 (N_10500,N_10125,N_9847);
xor U10501 (N_10501,N_9974,N_10015);
and U10502 (N_10502,N_10151,N_9989);
or U10503 (N_10503,N_10312,N_9961);
or U10504 (N_10504,N_10367,N_10260);
xor U10505 (N_10505,N_10388,N_10213);
nand U10506 (N_10506,N_10341,N_10129);
nor U10507 (N_10507,N_10355,N_10262);
or U10508 (N_10508,N_10362,N_10130);
xor U10509 (N_10509,N_10373,N_9971);
and U10510 (N_10510,N_10054,N_10405);
xor U10511 (N_10511,N_10127,N_10164);
and U10512 (N_10512,N_9871,N_9824);
or U10513 (N_10513,N_9957,N_9808);
nand U10514 (N_10514,N_10263,N_10398);
and U10515 (N_10515,N_9900,N_10295);
nand U10516 (N_10516,N_9897,N_10050);
nand U10517 (N_10517,N_10119,N_10197);
nand U10518 (N_10518,N_10422,N_9868);
and U10519 (N_10519,N_10493,N_10496);
or U10520 (N_10520,N_10318,N_9785);
nor U10521 (N_10521,N_10358,N_10048);
nand U10522 (N_10522,N_10236,N_10225);
nand U10523 (N_10523,N_9857,N_10448);
nand U10524 (N_10524,N_9763,N_10472);
nor U10525 (N_10525,N_10096,N_9906);
or U10526 (N_10526,N_10321,N_10399);
xor U10527 (N_10527,N_9915,N_9817);
nor U10528 (N_10528,N_9784,N_10267);
or U10529 (N_10529,N_10171,N_9921);
or U10530 (N_10530,N_10175,N_10099);
xnor U10531 (N_10531,N_10156,N_10401);
nand U10532 (N_10532,N_9835,N_10316);
xnor U10533 (N_10533,N_10177,N_10394);
xnor U10534 (N_10534,N_10188,N_10149);
or U10535 (N_10535,N_10081,N_10074);
nor U10536 (N_10536,N_10483,N_10368);
nand U10537 (N_10537,N_10466,N_9805);
or U10538 (N_10538,N_10469,N_10354);
or U10539 (N_10539,N_10176,N_10402);
or U10540 (N_10540,N_9902,N_9872);
xor U10541 (N_10541,N_9759,N_10202);
and U10542 (N_10542,N_10086,N_10345);
or U10543 (N_10543,N_10449,N_10323);
xor U10544 (N_10544,N_9799,N_9774);
and U10545 (N_10545,N_10238,N_9832);
nor U10546 (N_10546,N_9765,N_10397);
and U10547 (N_10547,N_10100,N_10311);
xor U10548 (N_10548,N_9886,N_10499);
xnor U10549 (N_10549,N_10205,N_10073);
nor U10550 (N_10550,N_10045,N_9852);
nand U10551 (N_10551,N_10049,N_10001);
and U10552 (N_10552,N_9853,N_10384);
and U10553 (N_10553,N_10350,N_10196);
nor U10554 (N_10554,N_9814,N_10221);
and U10555 (N_10555,N_10155,N_9908);
xnor U10556 (N_10556,N_10270,N_9864);
and U10557 (N_10557,N_9925,N_10140);
nor U10558 (N_10558,N_9792,N_10037);
xor U10559 (N_10559,N_9786,N_10143);
xnor U10560 (N_10560,N_10110,N_9954);
nor U10561 (N_10561,N_9809,N_10056);
xor U10562 (N_10562,N_10277,N_9770);
or U10563 (N_10563,N_10233,N_10219);
nor U10564 (N_10564,N_9926,N_9843);
nand U10565 (N_10565,N_10080,N_10315);
nor U10566 (N_10566,N_9938,N_10082);
nand U10567 (N_10567,N_9757,N_10439);
xor U10568 (N_10568,N_9875,N_10363);
nand U10569 (N_10569,N_10133,N_9800);
and U10570 (N_10570,N_10306,N_9993);
xor U10571 (N_10571,N_10297,N_10328);
nor U10572 (N_10572,N_10419,N_10455);
nor U10573 (N_10573,N_10454,N_9910);
nor U10574 (N_10574,N_10378,N_10136);
nand U10575 (N_10575,N_9963,N_10246);
nor U10576 (N_10576,N_10087,N_9771);
and U10577 (N_10577,N_10288,N_9881);
xnor U10578 (N_10578,N_9994,N_10434);
nor U10579 (N_10579,N_10215,N_9801);
nor U10580 (N_10580,N_9812,N_9945);
xor U10581 (N_10581,N_9816,N_10486);
and U10582 (N_10582,N_10017,N_10112);
nand U10583 (N_10583,N_10418,N_9761);
and U10584 (N_10584,N_10174,N_10124);
nand U10585 (N_10585,N_10141,N_9919);
or U10586 (N_10586,N_10359,N_9754);
nand U10587 (N_10587,N_10072,N_9888);
nand U10588 (N_10588,N_9956,N_9909);
nor U10589 (N_10589,N_10022,N_10189);
or U10590 (N_10590,N_10020,N_10413);
xnor U10591 (N_10591,N_10069,N_10239);
and U10592 (N_10592,N_10446,N_10490);
and U10593 (N_10593,N_9968,N_10153);
xor U10594 (N_10594,N_10222,N_10217);
nand U10595 (N_10595,N_10374,N_10353);
xnor U10596 (N_10596,N_10357,N_10249);
nand U10597 (N_10597,N_10223,N_9969);
or U10598 (N_10598,N_10029,N_10303);
xnor U10599 (N_10599,N_10317,N_10013);
and U10600 (N_10600,N_9756,N_10060);
nand U10601 (N_10601,N_10123,N_9924);
nor U10602 (N_10602,N_10296,N_10093);
nor U10603 (N_10603,N_10337,N_9985);
and U10604 (N_10604,N_10292,N_9939);
xor U10605 (N_10605,N_10021,N_10254);
xnor U10606 (N_10606,N_9911,N_9892);
or U10607 (N_10607,N_10309,N_10108);
xor U10608 (N_10608,N_9917,N_10115);
nor U10609 (N_10609,N_10407,N_10279);
or U10610 (N_10610,N_9987,N_10476);
or U10611 (N_10611,N_9949,N_10495);
xor U10612 (N_10612,N_9865,N_10244);
nor U10613 (N_10613,N_10160,N_9807);
nor U10614 (N_10614,N_10227,N_9947);
and U10615 (N_10615,N_10165,N_10332);
nand U10616 (N_10616,N_9793,N_10370);
nand U10617 (N_10617,N_9980,N_9791);
nor U10618 (N_10618,N_10342,N_10425);
nand U10619 (N_10619,N_10033,N_9982);
or U10620 (N_10620,N_10085,N_9838);
and U10621 (N_10621,N_9927,N_9788);
xor U10622 (N_10622,N_9849,N_10247);
or U10623 (N_10623,N_9923,N_10163);
or U10624 (N_10624,N_9894,N_10391);
nor U10625 (N_10625,N_10387,N_9929);
and U10626 (N_10626,N_10343,N_9967);
or U10627 (N_10627,N_10030,N_10237);
and U10628 (N_10628,N_9932,N_9890);
nand U10629 (N_10629,N_10137,N_10242);
or U10630 (N_10630,N_10273,N_9946);
nand U10631 (N_10631,N_9914,N_10159);
nand U10632 (N_10632,N_10404,N_9753);
or U10633 (N_10633,N_10078,N_9804);
xor U10634 (N_10634,N_9896,N_10479);
or U10635 (N_10635,N_10305,N_10198);
and U10636 (N_10636,N_10464,N_10106);
nand U10637 (N_10637,N_10026,N_10480);
and U10638 (N_10638,N_9950,N_9995);
nor U10639 (N_10639,N_9782,N_9955);
xnor U10640 (N_10640,N_9827,N_10134);
nor U10641 (N_10641,N_10429,N_10460);
xnor U10642 (N_10642,N_9972,N_10104);
or U10643 (N_10643,N_9882,N_10066);
nand U10644 (N_10644,N_10302,N_10044);
xor U10645 (N_10645,N_10204,N_10284);
or U10646 (N_10646,N_9930,N_10349);
and U10647 (N_10647,N_10392,N_9964);
xor U10648 (N_10648,N_10310,N_10301);
nor U10649 (N_10649,N_9918,N_10276);
or U10650 (N_10650,N_10436,N_10327);
nand U10651 (N_10651,N_9883,N_10408);
or U10652 (N_10652,N_10032,N_10307);
and U10653 (N_10653,N_10481,N_9889);
nand U10654 (N_10654,N_10006,N_10152);
nor U10655 (N_10655,N_10102,N_10036);
nand U10656 (N_10656,N_9867,N_9895);
xnor U10657 (N_10657,N_10409,N_10132);
nand U10658 (N_10658,N_9796,N_10338);
nor U10659 (N_10659,N_10325,N_10077);
or U10660 (N_10660,N_10142,N_9940);
or U10661 (N_10661,N_9811,N_9880);
nor U10662 (N_10662,N_10488,N_10287);
nand U10663 (N_10663,N_10116,N_9819);
nand U10664 (N_10664,N_9777,N_9821);
and U10665 (N_10665,N_9986,N_10052);
or U10666 (N_10666,N_10235,N_10471);
xnor U10667 (N_10667,N_9776,N_9787);
and U10668 (N_10668,N_10041,N_10440);
xor U10669 (N_10669,N_10111,N_10462);
nor U10670 (N_10670,N_10477,N_9877);
xor U10671 (N_10671,N_10344,N_9988);
and U10672 (N_10672,N_10326,N_10194);
nor U10673 (N_10673,N_10426,N_9977);
nor U10674 (N_10674,N_10169,N_10181);
nor U10675 (N_10675,N_10375,N_9795);
nor U10676 (N_10676,N_10322,N_10084);
and U10677 (N_10677,N_9869,N_10308);
and U10678 (N_10678,N_10118,N_9903);
xor U10679 (N_10679,N_10324,N_10280);
and U10680 (N_10680,N_10062,N_10393);
nand U10681 (N_10681,N_9934,N_10039);
and U10682 (N_10682,N_10201,N_9758);
nor U10683 (N_10683,N_10079,N_9851);
nor U10684 (N_10684,N_9899,N_9887);
and U10685 (N_10685,N_10271,N_10070);
nor U10686 (N_10686,N_10269,N_10256);
nand U10687 (N_10687,N_9822,N_9813);
nor U10688 (N_10688,N_10055,N_10445);
nand U10689 (N_10689,N_9965,N_10382);
nor U10690 (N_10690,N_10335,N_9780);
or U10691 (N_10691,N_10458,N_9959);
nor U10692 (N_10692,N_10200,N_10154);
and U10693 (N_10693,N_10061,N_9992);
nor U10694 (N_10694,N_10461,N_9845);
and U10695 (N_10695,N_10494,N_10360);
nand U10696 (N_10696,N_10386,N_9933);
and U10697 (N_10697,N_9815,N_10218);
or U10698 (N_10698,N_10264,N_10441);
xnor U10699 (N_10699,N_10012,N_10379);
or U10700 (N_10700,N_10075,N_10424);
or U10701 (N_10701,N_10145,N_10047);
nor U10702 (N_10702,N_9767,N_9844);
nand U10703 (N_10703,N_9751,N_10234);
and U10704 (N_10704,N_10423,N_10383);
or U10705 (N_10705,N_10459,N_10331);
or U10706 (N_10706,N_10144,N_10427);
xnor U10707 (N_10707,N_10065,N_9973);
xnor U10708 (N_10708,N_9848,N_9958);
or U10709 (N_10709,N_10340,N_9941);
nand U10710 (N_10710,N_10245,N_9943);
nor U10711 (N_10711,N_10334,N_10299);
xor U10712 (N_10712,N_9859,N_10083);
nor U10713 (N_10713,N_9820,N_9936);
nand U10714 (N_10714,N_10230,N_10437);
or U10715 (N_10715,N_10433,N_10465);
xnor U10716 (N_10716,N_10031,N_9952);
xnor U10717 (N_10717,N_9990,N_10320);
nor U10718 (N_10718,N_9823,N_10452);
or U10719 (N_10719,N_9837,N_10431);
nand U10720 (N_10720,N_10451,N_9866);
xnor U10721 (N_10721,N_9850,N_9798);
xnor U10722 (N_10722,N_10173,N_9810);
nand U10723 (N_10723,N_10442,N_10417);
and U10724 (N_10724,N_9970,N_10007);
xnor U10725 (N_10725,N_10406,N_10489);
xnor U10726 (N_10726,N_10148,N_9904);
nand U10727 (N_10727,N_10313,N_10180);
and U10728 (N_10728,N_10064,N_10261);
or U10729 (N_10729,N_10008,N_10038);
nand U10730 (N_10730,N_10105,N_10298);
and U10731 (N_10731,N_10035,N_9764);
nor U10732 (N_10732,N_10019,N_10113);
nor U10733 (N_10733,N_10122,N_9778);
xnor U10734 (N_10734,N_10168,N_9942);
or U10735 (N_10735,N_9854,N_10094);
and U10736 (N_10736,N_9818,N_10369);
nor U10737 (N_10737,N_10259,N_10498);
xnor U10738 (N_10738,N_10329,N_10051);
and U10739 (N_10739,N_10058,N_9842);
nor U10740 (N_10740,N_10206,N_10272);
xor U10741 (N_10741,N_10281,N_10024);
or U10742 (N_10742,N_10275,N_10098);
or U10743 (N_10743,N_10182,N_10128);
nand U10744 (N_10744,N_10057,N_9873);
and U10745 (N_10745,N_10166,N_10067);
xor U10746 (N_10746,N_10356,N_10135);
nand U10747 (N_10747,N_10252,N_10193);
xor U10748 (N_10748,N_10251,N_10157);
nor U10749 (N_10749,N_9901,N_9861);
nor U10750 (N_10750,N_10131,N_9825);
nor U10751 (N_10751,N_10250,N_10179);
nor U10752 (N_10752,N_9797,N_10209);
xnor U10753 (N_10753,N_10396,N_9863);
and U10754 (N_10754,N_9976,N_10412);
nand U10755 (N_10755,N_10150,N_10042);
nor U10756 (N_10756,N_10183,N_10034);
and U10757 (N_10757,N_10071,N_9953);
or U10758 (N_10758,N_10372,N_9991);
or U10759 (N_10759,N_9905,N_9978);
xnor U10760 (N_10760,N_10258,N_10456);
nor U10761 (N_10761,N_10389,N_9931);
nand U10762 (N_10762,N_9750,N_9846);
nand U10763 (N_10763,N_10004,N_10146);
nand U10764 (N_10764,N_10184,N_10282);
nor U10765 (N_10765,N_10027,N_10126);
nand U10766 (N_10766,N_10366,N_10395);
xor U10767 (N_10767,N_9913,N_10097);
or U10768 (N_10768,N_9912,N_10158);
xnor U10769 (N_10769,N_9783,N_10257);
nor U10770 (N_10770,N_10385,N_10224);
and U10771 (N_10771,N_10203,N_10482);
and U10772 (N_10772,N_10336,N_10162);
xnor U10773 (N_10773,N_10278,N_9885);
nor U10774 (N_10774,N_9862,N_10294);
and U10775 (N_10775,N_10232,N_10346);
nand U10776 (N_10776,N_10185,N_10023);
and U10777 (N_10777,N_10289,N_10300);
and U10778 (N_10778,N_10025,N_9935);
xor U10779 (N_10779,N_10190,N_10364);
and U10780 (N_10780,N_9858,N_10010);
nand U10781 (N_10781,N_9790,N_10485);
xor U10782 (N_10782,N_10028,N_10005);
or U10783 (N_10783,N_10103,N_10438);
xnor U10784 (N_10784,N_10450,N_9884);
nor U10785 (N_10785,N_9999,N_10231);
nand U10786 (N_10786,N_10248,N_10068);
and U10787 (N_10787,N_9983,N_10443);
and U10788 (N_10788,N_10444,N_10290);
nand U10789 (N_10789,N_10009,N_9779);
or U10790 (N_10790,N_9755,N_9856);
or U10791 (N_10791,N_10243,N_10241);
xnor U10792 (N_10792,N_10274,N_9831);
xnor U10793 (N_10793,N_9937,N_10453);
xor U10794 (N_10794,N_10043,N_10416);
and U10795 (N_10795,N_10212,N_9752);
xnor U10796 (N_10796,N_9876,N_10381);
nor U10797 (N_10797,N_10207,N_9833);
nand U10798 (N_10798,N_9836,N_10040);
xor U10799 (N_10799,N_10109,N_10211);
or U10800 (N_10800,N_9803,N_10319);
xor U10801 (N_10801,N_9891,N_10410);
or U10802 (N_10802,N_10101,N_9996);
nor U10803 (N_10803,N_9839,N_10255);
nand U10804 (N_10804,N_10053,N_10161);
or U10805 (N_10805,N_10214,N_9794);
or U10806 (N_10806,N_9916,N_9775);
and U10807 (N_10807,N_10046,N_9975);
or U10808 (N_10808,N_9806,N_9997);
or U10809 (N_10809,N_10147,N_9981);
or U10810 (N_10810,N_10228,N_9998);
or U10811 (N_10811,N_9802,N_10000);
nand U10812 (N_10812,N_10011,N_9830);
or U10813 (N_10813,N_10090,N_9928);
xnor U10814 (N_10814,N_10304,N_10240);
nor U10815 (N_10815,N_10470,N_10187);
or U10816 (N_10816,N_10059,N_10265);
nand U10817 (N_10817,N_10063,N_9962);
or U10818 (N_10818,N_9826,N_10229);
and U10819 (N_10819,N_10428,N_9760);
or U10820 (N_10820,N_10473,N_9979);
nor U10821 (N_10821,N_9768,N_10195);
and U10822 (N_10822,N_10014,N_9898);
nand U10823 (N_10823,N_10411,N_9781);
nand U10824 (N_10824,N_10474,N_10018);
and U10825 (N_10825,N_9984,N_10220);
xnor U10826 (N_10826,N_9828,N_9766);
or U10827 (N_10827,N_10463,N_9948);
nand U10828 (N_10828,N_10016,N_10192);
and U10829 (N_10829,N_10420,N_10091);
nor U10830 (N_10830,N_10293,N_10447);
nand U10831 (N_10831,N_10208,N_10199);
and U10832 (N_10832,N_9907,N_9879);
and U10833 (N_10833,N_10491,N_9840);
nand U10834 (N_10834,N_9878,N_10468);
and U10835 (N_10835,N_9769,N_10330);
nor U10836 (N_10836,N_10210,N_10457);
or U10837 (N_10837,N_9841,N_10107);
xor U10838 (N_10838,N_10478,N_10114);
or U10839 (N_10839,N_9951,N_9772);
nor U10840 (N_10840,N_9834,N_10430);
nor U10841 (N_10841,N_9860,N_10352);
nor U10842 (N_10842,N_10216,N_10467);
xnor U10843 (N_10843,N_10390,N_10351);
nand U10844 (N_10844,N_9966,N_10376);
or U10845 (N_10845,N_10286,N_10492);
nand U10846 (N_10846,N_9829,N_9870);
xor U10847 (N_10847,N_10172,N_10432);
nand U10848 (N_10848,N_10120,N_9922);
nand U10849 (N_10849,N_10400,N_10403);
nor U10850 (N_10850,N_10191,N_10348);
and U10851 (N_10851,N_10170,N_9920);
nand U10852 (N_10852,N_10186,N_10268);
and U10853 (N_10853,N_10092,N_9874);
nor U10854 (N_10854,N_9960,N_9893);
nand U10855 (N_10855,N_10138,N_10339);
or U10856 (N_10856,N_9944,N_10365);
nand U10857 (N_10857,N_10291,N_9789);
and U10858 (N_10858,N_10333,N_10253);
nand U10859 (N_10859,N_10117,N_10421);
nor U10860 (N_10860,N_10095,N_10314);
xnor U10861 (N_10861,N_10361,N_10285);
nor U10862 (N_10862,N_10167,N_10266);
or U10863 (N_10863,N_10178,N_10226);
xor U10864 (N_10864,N_10497,N_10283);
nand U10865 (N_10865,N_10475,N_10484);
or U10866 (N_10866,N_10002,N_10371);
nor U10867 (N_10867,N_10435,N_10139);
and U10868 (N_10868,N_10380,N_10121);
or U10869 (N_10869,N_10088,N_10347);
and U10870 (N_10870,N_9773,N_9762);
or U10871 (N_10871,N_10377,N_10415);
nand U10872 (N_10872,N_10089,N_10076);
and U10873 (N_10873,N_10003,N_10487);
nand U10874 (N_10874,N_9855,N_10414);
xnor U10875 (N_10875,N_10142,N_10488);
and U10876 (N_10876,N_9843,N_10183);
nand U10877 (N_10877,N_10003,N_9884);
or U10878 (N_10878,N_10496,N_10178);
nand U10879 (N_10879,N_10110,N_9879);
nor U10880 (N_10880,N_10152,N_10196);
nor U10881 (N_10881,N_9977,N_9851);
nand U10882 (N_10882,N_10179,N_9804);
nand U10883 (N_10883,N_10379,N_10129);
nand U10884 (N_10884,N_10018,N_10099);
and U10885 (N_10885,N_10130,N_10064);
and U10886 (N_10886,N_10231,N_10465);
nor U10887 (N_10887,N_10106,N_10452);
xor U10888 (N_10888,N_10415,N_9855);
nor U10889 (N_10889,N_9861,N_9980);
and U10890 (N_10890,N_10391,N_10188);
nand U10891 (N_10891,N_9758,N_9802);
nand U10892 (N_10892,N_10277,N_9838);
nor U10893 (N_10893,N_9904,N_10235);
nand U10894 (N_10894,N_10376,N_9924);
xor U10895 (N_10895,N_9845,N_10255);
or U10896 (N_10896,N_10324,N_9874);
and U10897 (N_10897,N_10225,N_10307);
or U10898 (N_10898,N_10242,N_9842);
xnor U10899 (N_10899,N_9983,N_9940);
nand U10900 (N_10900,N_10183,N_10143);
or U10901 (N_10901,N_10022,N_9808);
xnor U10902 (N_10902,N_10324,N_9938);
and U10903 (N_10903,N_9858,N_9839);
xnor U10904 (N_10904,N_10361,N_10061);
nor U10905 (N_10905,N_10035,N_10153);
nand U10906 (N_10906,N_10397,N_9959);
nand U10907 (N_10907,N_10433,N_9757);
or U10908 (N_10908,N_9938,N_10414);
xnor U10909 (N_10909,N_10420,N_10249);
nand U10910 (N_10910,N_10139,N_10030);
nor U10911 (N_10911,N_9767,N_10358);
and U10912 (N_10912,N_9842,N_10275);
or U10913 (N_10913,N_9854,N_9841);
nor U10914 (N_10914,N_9955,N_10058);
and U10915 (N_10915,N_10489,N_10317);
xor U10916 (N_10916,N_9973,N_9892);
or U10917 (N_10917,N_10111,N_10350);
xor U10918 (N_10918,N_10330,N_10319);
xnor U10919 (N_10919,N_10337,N_9912);
xnor U10920 (N_10920,N_10247,N_10048);
nand U10921 (N_10921,N_10437,N_9839);
nand U10922 (N_10922,N_9884,N_9781);
or U10923 (N_10923,N_9840,N_10417);
nor U10924 (N_10924,N_9964,N_9983);
or U10925 (N_10925,N_9949,N_10438);
nor U10926 (N_10926,N_10296,N_10109);
or U10927 (N_10927,N_9883,N_9849);
xor U10928 (N_10928,N_10309,N_10409);
nand U10929 (N_10929,N_9845,N_9876);
nand U10930 (N_10930,N_10265,N_10015);
nor U10931 (N_10931,N_9893,N_10124);
xor U10932 (N_10932,N_10274,N_9779);
or U10933 (N_10933,N_10423,N_10313);
xor U10934 (N_10934,N_10079,N_10246);
nor U10935 (N_10935,N_10065,N_10266);
nor U10936 (N_10936,N_9857,N_9868);
or U10937 (N_10937,N_10028,N_10256);
or U10938 (N_10938,N_9902,N_9862);
nand U10939 (N_10939,N_10368,N_10351);
xor U10940 (N_10940,N_9781,N_9865);
or U10941 (N_10941,N_10465,N_10119);
nand U10942 (N_10942,N_10394,N_10466);
nor U10943 (N_10943,N_9920,N_9837);
and U10944 (N_10944,N_10144,N_10468);
nor U10945 (N_10945,N_9982,N_9955);
nor U10946 (N_10946,N_9862,N_10415);
or U10947 (N_10947,N_10488,N_10132);
nand U10948 (N_10948,N_10446,N_10238);
nor U10949 (N_10949,N_10233,N_9773);
nor U10950 (N_10950,N_10065,N_9983);
xnor U10951 (N_10951,N_9987,N_10315);
xnor U10952 (N_10952,N_10262,N_10043);
xnor U10953 (N_10953,N_9824,N_10080);
nor U10954 (N_10954,N_9921,N_10488);
and U10955 (N_10955,N_10160,N_9776);
and U10956 (N_10956,N_10225,N_10126);
xnor U10957 (N_10957,N_10090,N_10313);
and U10958 (N_10958,N_10365,N_9833);
xnor U10959 (N_10959,N_10069,N_10179);
nor U10960 (N_10960,N_9923,N_9986);
xnor U10961 (N_10961,N_9790,N_10384);
nor U10962 (N_10962,N_10222,N_10367);
xor U10963 (N_10963,N_9945,N_10394);
nand U10964 (N_10964,N_10098,N_9916);
xnor U10965 (N_10965,N_10383,N_10249);
xnor U10966 (N_10966,N_10183,N_10212);
nand U10967 (N_10967,N_10096,N_10047);
nor U10968 (N_10968,N_9921,N_10294);
or U10969 (N_10969,N_10484,N_10185);
nand U10970 (N_10970,N_9798,N_10474);
nor U10971 (N_10971,N_9978,N_10427);
or U10972 (N_10972,N_9888,N_10477);
and U10973 (N_10973,N_9797,N_9821);
xnor U10974 (N_10974,N_10486,N_9979);
and U10975 (N_10975,N_10030,N_10477);
nor U10976 (N_10976,N_10291,N_10242);
nor U10977 (N_10977,N_9751,N_10008);
nor U10978 (N_10978,N_9992,N_9795);
and U10979 (N_10979,N_10295,N_10288);
nand U10980 (N_10980,N_9783,N_9918);
or U10981 (N_10981,N_10034,N_10223);
nand U10982 (N_10982,N_10085,N_9822);
and U10983 (N_10983,N_10299,N_10401);
nand U10984 (N_10984,N_10058,N_9822);
nor U10985 (N_10985,N_10044,N_10482);
xor U10986 (N_10986,N_9981,N_10418);
xor U10987 (N_10987,N_9825,N_9771);
or U10988 (N_10988,N_9914,N_10086);
or U10989 (N_10989,N_9943,N_9975);
nor U10990 (N_10990,N_10321,N_9916);
nor U10991 (N_10991,N_10271,N_10415);
xor U10992 (N_10992,N_10015,N_10411);
xnor U10993 (N_10993,N_10351,N_9986);
nor U10994 (N_10994,N_10480,N_10457);
and U10995 (N_10995,N_10232,N_10157);
nand U10996 (N_10996,N_9845,N_10266);
xor U10997 (N_10997,N_10324,N_10212);
nand U10998 (N_10998,N_10057,N_10011);
or U10999 (N_10999,N_9788,N_10460);
and U11000 (N_11000,N_9973,N_9985);
nand U11001 (N_11001,N_9975,N_10415);
nor U11002 (N_11002,N_9856,N_10008);
or U11003 (N_11003,N_10319,N_10093);
nand U11004 (N_11004,N_9854,N_10270);
xnor U11005 (N_11005,N_10357,N_9852);
or U11006 (N_11006,N_10056,N_10298);
or U11007 (N_11007,N_10015,N_10075);
nand U11008 (N_11008,N_9887,N_9864);
xnor U11009 (N_11009,N_10197,N_10233);
or U11010 (N_11010,N_10237,N_10428);
nor U11011 (N_11011,N_10141,N_9958);
and U11012 (N_11012,N_10437,N_10295);
nand U11013 (N_11013,N_10082,N_10038);
nor U11014 (N_11014,N_10204,N_10385);
and U11015 (N_11015,N_9808,N_10165);
nand U11016 (N_11016,N_9827,N_10200);
nand U11017 (N_11017,N_9896,N_10125);
or U11018 (N_11018,N_10075,N_10066);
nor U11019 (N_11019,N_9760,N_10048);
nand U11020 (N_11020,N_9955,N_9776);
nand U11021 (N_11021,N_9775,N_10488);
nand U11022 (N_11022,N_10048,N_10065);
nor U11023 (N_11023,N_10097,N_10250);
nor U11024 (N_11024,N_10027,N_9916);
or U11025 (N_11025,N_9859,N_9893);
or U11026 (N_11026,N_9795,N_10482);
and U11027 (N_11027,N_9913,N_9865);
or U11028 (N_11028,N_9869,N_9948);
nand U11029 (N_11029,N_10200,N_10370);
xnor U11030 (N_11030,N_9901,N_9916);
nand U11031 (N_11031,N_10026,N_9768);
or U11032 (N_11032,N_10472,N_10090);
and U11033 (N_11033,N_9868,N_9848);
nor U11034 (N_11034,N_10240,N_10395);
xnor U11035 (N_11035,N_10399,N_10091);
or U11036 (N_11036,N_10049,N_10459);
nor U11037 (N_11037,N_10194,N_9980);
and U11038 (N_11038,N_10261,N_10074);
or U11039 (N_11039,N_10272,N_10119);
nand U11040 (N_11040,N_10190,N_9832);
nand U11041 (N_11041,N_10380,N_9909);
or U11042 (N_11042,N_10093,N_10156);
and U11043 (N_11043,N_10435,N_10484);
or U11044 (N_11044,N_10269,N_10115);
and U11045 (N_11045,N_10112,N_10138);
and U11046 (N_11046,N_9927,N_10368);
nor U11047 (N_11047,N_10376,N_10344);
and U11048 (N_11048,N_10142,N_10315);
nand U11049 (N_11049,N_10175,N_10481);
nand U11050 (N_11050,N_9806,N_10368);
nor U11051 (N_11051,N_9854,N_10314);
nor U11052 (N_11052,N_10247,N_9979);
and U11053 (N_11053,N_9891,N_10089);
nor U11054 (N_11054,N_10406,N_9965);
nand U11055 (N_11055,N_10271,N_10055);
and U11056 (N_11056,N_9754,N_9769);
or U11057 (N_11057,N_10446,N_10301);
and U11058 (N_11058,N_10437,N_9809);
and U11059 (N_11059,N_9945,N_9871);
xor U11060 (N_11060,N_9924,N_10207);
nor U11061 (N_11061,N_10374,N_9866);
xor U11062 (N_11062,N_10378,N_9754);
nor U11063 (N_11063,N_10287,N_9936);
nor U11064 (N_11064,N_10002,N_10423);
and U11065 (N_11065,N_10424,N_9770);
xor U11066 (N_11066,N_10140,N_9785);
xnor U11067 (N_11067,N_9833,N_9942);
nor U11068 (N_11068,N_10118,N_10430);
nand U11069 (N_11069,N_9843,N_10292);
xnor U11070 (N_11070,N_10347,N_10103);
nand U11071 (N_11071,N_10408,N_10412);
nor U11072 (N_11072,N_10369,N_10230);
and U11073 (N_11073,N_10184,N_9952);
nand U11074 (N_11074,N_10413,N_10130);
and U11075 (N_11075,N_10133,N_10447);
or U11076 (N_11076,N_10250,N_9855);
xnor U11077 (N_11077,N_10297,N_9981);
or U11078 (N_11078,N_10432,N_10387);
xor U11079 (N_11079,N_10174,N_9879);
or U11080 (N_11080,N_10168,N_10350);
xor U11081 (N_11081,N_9951,N_9882);
xor U11082 (N_11082,N_9899,N_9855);
or U11083 (N_11083,N_10302,N_10104);
or U11084 (N_11084,N_10096,N_9945);
or U11085 (N_11085,N_10269,N_9885);
nor U11086 (N_11086,N_10234,N_10304);
nor U11087 (N_11087,N_9804,N_10220);
nor U11088 (N_11088,N_9845,N_10123);
nand U11089 (N_11089,N_10489,N_10017);
nand U11090 (N_11090,N_9895,N_9869);
nor U11091 (N_11091,N_9976,N_9752);
and U11092 (N_11092,N_9871,N_10265);
nand U11093 (N_11093,N_10038,N_10060);
nand U11094 (N_11094,N_10340,N_10056);
or U11095 (N_11095,N_10459,N_10096);
nand U11096 (N_11096,N_10075,N_10473);
nor U11097 (N_11097,N_10408,N_9902);
xnor U11098 (N_11098,N_10368,N_10180);
or U11099 (N_11099,N_10081,N_9885);
and U11100 (N_11100,N_10162,N_9871);
xor U11101 (N_11101,N_10244,N_9869);
nor U11102 (N_11102,N_9815,N_9923);
and U11103 (N_11103,N_10448,N_9753);
and U11104 (N_11104,N_9906,N_9785);
nor U11105 (N_11105,N_9952,N_10342);
nor U11106 (N_11106,N_10455,N_10406);
or U11107 (N_11107,N_10073,N_10052);
nor U11108 (N_11108,N_10126,N_10207);
or U11109 (N_11109,N_10085,N_10022);
xor U11110 (N_11110,N_10458,N_10313);
or U11111 (N_11111,N_10154,N_9992);
and U11112 (N_11112,N_10267,N_9975);
xnor U11113 (N_11113,N_10204,N_9941);
or U11114 (N_11114,N_10080,N_10147);
xnor U11115 (N_11115,N_10313,N_10194);
nand U11116 (N_11116,N_9844,N_9984);
or U11117 (N_11117,N_10381,N_9760);
nand U11118 (N_11118,N_10315,N_9948);
nand U11119 (N_11119,N_10358,N_10149);
and U11120 (N_11120,N_10446,N_9953);
and U11121 (N_11121,N_10278,N_10492);
and U11122 (N_11122,N_10239,N_10204);
nor U11123 (N_11123,N_10075,N_10166);
nand U11124 (N_11124,N_10208,N_10235);
nor U11125 (N_11125,N_10246,N_10310);
nor U11126 (N_11126,N_9970,N_10158);
nand U11127 (N_11127,N_10010,N_10290);
or U11128 (N_11128,N_10358,N_9917);
or U11129 (N_11129,N_10258,N_10332);
and U11130 (N_11130,N_10128,N_10337);
xor U11131 (N_11131,N_10438,N_9882);
or U11132 (N_11132,N_10124,N_10354);
nor U11133 (N_11133,N_9858,N_9841);
nor U11134 (N_11134,N_10052,N_10248);
xnor U11135 (N_11135,N_9829,N_10235);
and U11136 (N_11136,N_9971,N_10413);
nand U11137 (N_11137,N_10338,N_10299);
nor U11138 (N_11138,N_10162,N_10265);
xnor U11139 (N_11139,N_10088,N_9887);
and U11140 (N_11140,N_9888,N_10398);
nor U11141 (N_11141,N_10498,N_10129);
nand U11142 (N_11142,N_10149,N_10231);
nor U11143 (N_11143,N_10151,N_9750);
or U11144 (N_11144,N_10267,N_10484);
or U11145 (N_11145,N_10064,N_9807);
nor U11146 (N_11146,N_10469,N_10027);
and U11147 (N_11147,N_10200,N_9974);
or U11148 (N_11148,N_9810,N_10225);
and U11149 (N_11149,N_9782,N_9834);
nor U11150 (N_11150,N_9801,N_10440);
nand U11151 (N_11151,N_9857,N_10028);
xor U11152 (N_11152,N_9900,N_9846);
nand U11153 (N_11153,N_10002,N_10184);
nor U11154 (N_11154,N_10197,N_10048);
nand U11155 (N_11155,N_10494,N_10007);
nand U11156 (N_11156,N_10432,N_10264);
nor U11157 (N_11157,N_10467,N_9811);
and U11158 (N_11158,N_10439,N_10097);
or U11159 (N_11159,N_10049,N_9786);
or U11160 (N_11160,N_10031,N_10264);
xnor U11161 (N_11161,N_10386,N_10012);
nor U11162 (N_11162,N_10130,N_10461);
and U11163 (N_11163,N_10074,N_10131);
nand U11164 (N_11164,N_10002,N_9968);
nor U11165 (N_11165,N_10169,N_10027);
nor U11166 (N_11166,N_10265,N_9843);
xnor U11167 (N_11167,N_10098,N_10267);
and U11168 (N_11168,N_9788,N_10326);
nor U11169 (N_11169,N_9912,N_9799);
xor U11170 (N_11170,N_10096,N_9785);
xnor U11171 (N_11171,N_10450,N_10115);
nand U11172 (N_11172,N_10107,N_9813);
and U11173 (N_11173,N_10257,N_10414);
nand U11174 (N_11174,N_9908,N_9986);
or U11175 (N_11175,N_9948,N_10181);
nor U11176 (N_11176,N_9901,N_10453);
or U11177 (N_11177,N_9991,N_10410);
and U11178 (N_11178,N_9807,N_10469);
xnor U11179 (N_11179,N_9916,N_10467);
nand U11180 (N_11180,N_10088,N_9771);
nor U11181 (N_11181,N_10234,N_9806);
nor U11182 (N_11182,N_10005,N_9936);
nor U11183 (N_11183,N_10256,N_10058);
nand U11184 (N_11184,N_10446,N_9899);
nand U11185 (N_11185,N_10258,N_9933);
nand U11186 (N_11186,N_10248,N_9869);
nand U11187 (N_11187,N_10095,N_9968);
nor U11188 (N_11188,N_9821,N_10284);
and U11189 (N_11189,N_10268,N_9868);
or U11190 (N_11190,N_10161,N_10493);
and U11191 (N_11191,N_10032,N_9754);
nand U11192 (N_11192,N_9783,N_9987);
and U11193 (N_11193,N_10245,N_10120);
or U11194 (N_11194,N_10302,N_10238);
xor U11195 (N_11195,N_9857,N_9996);
nand U11196 (N_11196,N_10028,N_10131);
xnor U11197 (N_11197,N_9922,N_9842);
and U11198 (N_11198,N_9768,N_10395);
nand U11199 (N_11199,N_10061,N_10300);
or U11200 (N_11200,N_10411,N_10453);
xor U11201 (N_11201,N_9873,N_9818);
nor U11202 (N_11202,N_10374,N_10281);
or U11203 (N_11203,N_10227,N_10305);
or U11204 (N_11204,N_9875,N_10159);
nor U11205 (N_11205,N_10233,N_9904);
nor U11206 (N_11206,N_10299,N_9891);
nor U11207 (N_11207,N_9972,N_10370);
and U11208 (N_11208,N_9953,N_10169);
nor U11209 (N_11209,N_9822,N_10452);
or U11210 (N_11210,N_9987,N_10118);
xnor U11211 (N_11211,N_9924,N_9932);
and U11212 (N_11212,N_10113,N_10394);
nor U11213 (N_11213,N_9998,N_9807);
nor U11214 (N_11214,N_9818,N_10016);
nor U11215 (N_11215,N_9866,N_10417);
and U11216 (N_11216,N_10176,N_10195);
or U11217 (N_11217,N_10159,N_9819);
nand U11218 (N_11218,N_9875,N_9752);
xnor U11219 (N_11219,N_10185,N_9902);
nor U11220 (N_11220,N_10426,N_9949);
nand U11221 (N_11221,N_10061,N_10401);
xor U11222 (N_11222,N_10458,N_10228);
nand U11223 (N_11223,N_9998,N_9862);
xor U11224 (N_11224,N_10110,N_10408);
or U11225 (N_11225,N_10342,N_10362);
nor U11226 (N_11226,N_10127,N_10447);
nor U11227 (N_11227,N_10207,N_10320);
or U11228 (N_11228,N_10225,N_9794);
or U11229 (N_11229,N_9795,N_10197);
and U11230 (N_11230,N_10322,N_9898);
nand U11231 (N_11231,N_10117,N_10133);
nor U11232 (N_11232,N_10499,N_10210);
nor U11233 (N_11233,N_9810,N_9954);
nand U11234 (N_11234,N_10099,N_10093);
nand U11235 (N_11235,N_9881,N_9886);
or U11236 (N_11236,N_10260,N_10068);
or U11237 (N_11237,N_9823,N_10168);
nor U11238 (N_11238,N_9753,N_10203);
or U11239 (N_11239,N_10010,N_9832);
nand U11240 (N_11240,N_10246,N_9908);
and U11241 (N_11241,N_10477,N_10349);
nand U11242 (N_11242,N_10370,N_10194);
nor U11243 (N_11243,N_9844,N_10397);
xnor U11244 (N_11244,N_10117,N_9771);
and U11245 (N_11245,N_9863,N_10452);
or U11246 (N_11246,N_10001,N_9789);
nand U11247 (N_11247,N_10406,N_9788);
nor U11248 (N_11248,N_9935,N_10304);
or U11249 (N_11249,N_10472,N_10101);
nor U11250 (N_11250,N_10621,N_10580);
nand U11251 (N_11251,N_10588,N_10637);
or U11252 (N_11252,N_10917,N_11120);
xor U11253 (N_11253,N_10968,N_10875);
or U11254 (N_11254,N_10925,N_10636);
nor U11255 (N_11255,N_11000,N_10523);
xor U11256 (N_11256,N_11169,N_10914);
and U11257 (N_11257,N_11221,N_10891);
or U11258 (N_11258,N_11190,N_10806);
xor U11259 (N_11259,N_10955,N_10851);
nor U11260 (N_11260,N_10660,N_10829);
and U11261 (N_11261,N_10900,N_10516);
nor U11262 (N_11262,N_11235,N_10513);
nor U11263 (N_11263,N_10929,N_11044);
nor U11264 (N_11264,N_10772,N_10840);
nor U11265 (N_11265,N_11213,N_10501);
xnor U11266 (N_11266,N_10850,N_10540);
nand U11267 (N_11267,N_11074,N_11089);
and U11268 (N_11268,N_10777,N_10833);
or U11269 (N_11269,N_10729,N_11162);
xor U11270 (N_11270,N_11116,N_10894);
xor U11271 (N_11271,N_10878,N_11129);
and U11272 (N_11272,N_11019,N_10932);
or U11273 (N_11273,N_10574,N_11094);
nand U11274 (N_11274,N_10532,N_10852);
nor U11275 (N_11275,N_10763,N_11037);
xor U11276 (N_11276,N_10794,N_10944);
xor U11277 (N_11277,N_11146,N_11036);
nor U11278 (N_11278,N_11052,N_10895);
or U11279 (N_11279,N_10896,N_10776);
nor U11280 (N_11280,N_10564,N_10521);
nor U11281 (N_11281,N_10774,N_11075);
and U11282 (N_11282,N_10593,N_11210);
nor U11283 (N_11283,N_11144,N_10718);
or U11284 (N_11284,N_11027,N_10893);
nor U11285 (N_11285,N_10957,N_10578);
and U11286 (N_11286,N_10611,N_10725);
and U11287 (N_11287,N_10535,N_11164);
or U11288 (N_11288,N_11200,N_11048);
and U11289 (N_11289,N_10715,N_11243);
xnor U11290 (N_11290,N_10815,N_10835);
xnor U11291 (N_11291,N_10541,N_11140);
and U11292 (N_11292,N_10619,N_11185);
nand U11293 (N_11293,N_10842,N_10868);
nor U11294 (N_11294,N_11077,N_10614);
and U11295 (N_11295,N_11108,N_11104);
xnor U11296 (N_11296,N_11125,N_11232);
nor U11297 (N_11297,N_10675,N_11192);
xor U11298 (N_11298,N_11087,N_10740);
nand U11299 (N_11299,N_11069,N_10522);
and U11300 (N_11300,N_10890,N_10988);
nand U11301 (N_11301,N_11004,N_10892);
nand U11302 (N_11302,N_11101,N_10762);
xor U11303 (N_11303,N_10809,N_11127);
and U11304 (N_11304,N_10814,N_10692);
nor U11305 (N_11305,N_11078,N_10935);
nand U11306 (N_11306,N_11092,N_10722);
and U11307 (N_11307,N_11156,N_10993);
or U11308 (N_11308,N_11006,N_10884);
and U11309 (N_11309,N_10834,N_11173);
nand U11310 (N_11310,N_10604,N_10951);
xnor U11311 (N_11311,N_10572,N_10671);
or U11312 (N_11312,N_11042,N_11241);
nor U11313 (N_11313,N_10606,N_11238);
or U11314 (N_11314,N_10888,N_11194);
and U11315 (N_11315,N_11193,N_10537);
nand U11316 (N_11316,N_11188,N_10727);
or U11317 (N_11317,N_10986,N_10886);
or U11318 (N_11318,N_11109,N_11060);
and U11319 (N_11319,N_10802,N_10934);
nand U11320 (N_11320,N_11072,N_11240);
or U11321 (N_11321,N_10966,N_10976);
nand U11322 (N_11322,N_10629,N_11033);
nand U11323 (N_11323,N_11136,N_10573);
or U11324 (N_11324,N_10755,N_10939);
xnor U11325 (N_11325,N_10870,N_10652);
nand U11326 (N_11326,N_10643,N_10552);
nor U11327 (N_11327,N_10743,N_11132);
xnor U11328 (N_11328,N_10947,N_10674);
or U11329 (N_11329,N_10563,N_11008);
nand U11330 (N_11330,N_10577,N_11047);
xor U11331 (N_11331,N_10529,N_10766);
xnor U11332 (N_11332,N_10867,N_11028);
nor U11333 (N_11333,N_10985,N_10817);
nand U11334 (N_11334,N_10634,N_10848);
or U11335 (N_11335,N_10942,N_10977);
and U11336 (N_11336,N_11198,N_10964);
or U11337 (N_11337,N_11001,N_10555);
and U11338 (N_11338,N_10994,N_10758);
xnor U11339 (N_11339,N_10707,N_11152);
and U11340 (N_11340,N_10741,N_11212);
xnor U11341 (N_11341,N_10981,N_10667);
nor U11342 (N_11342,N_10754,N_10769);
nor U11343 (N_11343,N_11216,N_10841);
xor U11344 (N_11344,N_10723,N_11218);
nor U11345 (N_11345,N_11070,N_10873);
and U11346 (N_11346,N_11141,N_10680);
nand U11347 (N_11347,N_10864,N_10686);
xor U11348 (N_11348,N_10681,N_10791);
and U11349 (N_11349,N_10736,N_11040);
or U11350 (N_11350,N_10823,N_11195);
nor U11351 (N_11351,N_10906,N_11021);
nand U11352 (N_11352,N_10733,N_11045);
nand U11353 (N_11353,N_10531,N_10519);
xor U11354 (N_11354,N_11172,N_11170);
or U11355 (N_11355,N_10633,N_10605);
nor U11356 (N_11356,N_10861,N_11026);
nand U11357 (N_11357,N_10688,N_11063);
or U11358 (N_11358,N_10926,N_10909);
xnor U11359 (N_11359,N_10609,N_10992);
and U11360 (N_11360,N_10553,N_10533);
and U11361 (N_11361,N_11211,N_11056);
nand U11362 (N_11362,N_10797,N_11180);
nand U11363 (N_11363,N_11154,N_11130);
nor U11364 (N_11364,N_10624,N_10590);
nor U11365 (N_11365,N_11208,N_10677);
and U11366 (N_11366,N_10607,N_10856);
or U11367 (N_11367,N_10732,N_10865);
nor U11368 (N_11368,N_10781,N_10941);
or U11369 (N_11369,N_10770,N_10931);
or U11370 (N_11370,N_11046,N_10622);
xnor U11371 (N_11371,N_10653,N_10560);
or U11372 (N_11372,N_10980,N_10698);
and U11373 (N_11373,N_10544,N_10728);
or U11374 (N_11374,N_10946,N_10584);
xor U11375 (N_11375,N_10846,N_10887);
or U11376 (N_11376,N_10627,N_10587);
xor U11377 (N_11377,N_11071,N_10921);
and U11378 (N_11378,N_10534,N_10617);
nor U11379 (N_11379,N_10596,N_10706);
nor U11380 (N_11380,N_11189,N_10821);
nand U11381 (N_11381,N_10928,N_10876);
xnor U11382 (N_11382,N_10717,N_11123);
or U11383 (N_11383,N_10866,N_11176);
xnor U11384 (N_11384,N_10649,N_10613);
xor U11385 (N_11385,N_11148,N_11002);
nor U11386 (N_11386,N_11088,N_10787);
or U11387 (N_11387,N_11203,N_10626);
or U11388 (N_11388,N_10549,N_10710);
nand U11389 (N_11389,N_10830,N_10703);
or U11390 (N_11390,N_10836,N_11206);
nor U11391 (N_11391,N_10704,N_11247);
xnor U11392 (N_11392,N_10881,N_10954);
or U11393 (N_11393,N_11233,N_10503);
nand U11394 (N_11394,N_10525,N_10602);
xnor U11395 (N_11395,N_11107,N_10752);
nand U11396 (N_11396,N_10709,N_10508);
nand U11397 (N_11397,N_10845,N_11005);
or U11398 (N_11398,N_10838,N_10880);
xor U11399 (N_11399,N_10586,N_10520);
xnor U11400 (N_11400,N_10975,N_10765);
nand U11401 (N_11401,N_10789,N_11058);
nand U11402 (N_11402,N_10872,N_11068);
nand U11403 (N_11403,N_10757,N_10664);
and U11404 (N_11404,N_10662,N_10625);
xor U11405 (N_11405,N_10623,N_10550);
or U11406 (N_11406,N_10601,N_11093);
nor U11407 (N_11407,N_11030,N_11017);
or U11408 (N_11408,N_11115,N_11034);
nor U11409 (N_11409,N_10663,N_10857);
or U11410 (N_11410,N_10665,N_10673);
or U11411 (N_11411,N_10788,N_11145);
or U11412 (N_11412,N_10701,N_10933);
xnor U11413 (N_11413,N_10991,N_10775);
or U11414 (N_11414,N_10656,N_11201);
xnor U11415 (N_11415,N_10764,N_11118);
or U11416 (N_11416,N_10554,N_10582);
or U11417 (N_11417,N_10889,N_11143);
nor U11418 (N_11418,N_10818,N_10877);
or U11419 (N_11419,N_10542,N_11237);
and U11420 (N_11420,N_10779,N_10970);
or U11421 (N_11421,N_11022,N_10798);
and U11422 (N_11422,N_10684,N_10545);
nand U11423 (N_11423,N_10509,N_10967);
and U11424 (N_11424,N_10915,N_10696);
xnor U11425 (N_11425,N_10863,N_11196);
and U11426 (N_11426,N_10882,N_11039);
xor U11427 (N_11427,N_11139,N_11090);
nand U11428 (N_11428,N_10902,N_11153);
and U11429 (N_11429,N_10828,N_11095);
and U11430 (N_11430,N_10989,N_10559);
and U11431 (N_11431,N_10569,N_10911);
nand U11432 (N_11432,N_10594,N_11029);
xnor U11433 (N_11433,N_10530,N_10803);
or U11434 (N_11434,N_10810,N_10747);
xor U11435 (N_11435,N_10517,N_10735);
xnor U11436 (N_11436,N_11003,N_10913);
xor U11437 (N_11437,N_10746,N_11084);
or U11438 (N_11438,N_10910,N_10953);
and U11439 (N_11439,N_10843,N_10855);
or U11440 (N_11440,N_10650,N_10753);
or U11441 (N_11441,N_10854,N_10641);
nor U11442 (N_11442,N_11219,N_10568);
or U11443 (N_11443,N_11174,N_10672);
nor U11444 (N_11444,N_10832,N_11049);
nor U11445 (N_11445,N_11245,N_10640);
and U11446 (N_11446,N_10571,N_10987);
or U11447 (N_11447,N_10585,N_10595);
or U11448 (N_11448,N_10603,N_10598);
nor U11449 (N_11449,N_11158,N_11227);
xor U11450 (N_11450,N_10796,N_11249);
nor U11451 (N_11451,N_10724,N_11099);
nand U11452 (N_11452,N_11166,N_10645);
nand U11453 (N_11453,N_10924,N_11137);
nor U11454 (N_11454,N_11182,N_10940);
nor U11455 (N_11455,N_11117,N_11128);
nand U11456 (N_11456,N_10731,N_11179);
and U11457 (N_11457,N_10514,N_10825);
or U11458 (N_11458,N_11014,N_11112);
nor U11459 (N_11459,N_10599,N_11124);
or U11460 (N_11460,N_11018,N_10804);
or U11461 (N_11461,N_10904,N_10635);
nand U11462 (N_11462,N_11224,N_10527);
nor U11463 (N_11463,N_11051,N_11106);
nor U11464 (N_11464,N_10901,N_10812);
and U11465 (N_11465,N_11100,N_11083);
and U11466 (N_11466,N_10759,N_10839);
nand U11467 (N_11467,N_10858,N_11012);
xnor U11468 (N_11468,N_10767,N_10507);
nand U11469 (N_11469,N_10918,N_10956);
xnor U11470 (N_11470,N_11151,N_10734);
nor U11471 (N_11471,N_10923,N_11102);
nand U11472 (N_11472,N_11248,N_11035);
nor U11473 (N_11473,N_10659,N_10853);
nand U11474 (N_11474,N_10642,N_11062);
and U11475 (N_11475,N_10936,N_11105);
or U11476 (N_11476,N_10515,N_10714);
xnor U11477 (N_11477,N_11065,N_10512);
nor U11478 (N_11478,N_10631,N_10971);
xor U11479 (N_11479,N_10801,N_10920);
or U11480 (N_11480,N_10963,N_10995);
and U11481 (N_11481,N_11142,N_10597);
and U11482 (N_11482,N_10807,N_11157);
or U11483 (N_11483,N_10600,N_10705);
and U11484 (N_11484,N_10615,N_10927);
xor U11485 (N_11485,N_11159,N_10974);
nor U11486 (N_11486,N_10778,N_11199);
xor U11487 (N_11487,N_10528,N_11187);
or U11488 (N_11488,N_11015,N_11114);
xor U11489 (N_11489,N_10742,N_11031);
xor U11490 (N_11490,N_11223,N_11214);
or U11491 (N_11491,N_11085,N_11082);
xor U11492 (N_11492,N_11121,N_10999);
nand U11493 (N_11493,N_11205,N_10819);
or U11494 (N_11494,N_10952,N_10518);
nand U11495 (N_11495,N_10849,N_10800);
or U11496 (N_11496,N_11009,N_10700);
and U11497 (N_11497,N_11041,N_10869);
or U11498 (N_11498,N_10500,N_11236);
and U11499 (N_11499,N_11186,N_10524);
or U11500 (N_11500,N_10996,N_11043);
nand U11501 (N_11501,N_10962,N_10561);
nand U11502 (N_11502,N_11225,N_10676);
or U11503 (N_11503,N_11010,N_10655);
and U11504 (N_11504,N_11081,N_10937);
nor U11505 (N_11505,N_11057,N_10546);
nand U11506 (N_11506,N_10938,N_10583);
and U11507 (N_11507,N_11230,N_10689);
and U11508 (N_11508,N_10945,N_11016);
nor U11509 (N_11509,N_10847,N_11079);
xor U11510 (N_11510,N_11020,N_11165);
nor U11511 (N_11511,N_11134,N_10756);
nand U11512 (N_11512,N_10874,N_10912);
and U11513 (N_11513,N_10502,N_10773);
nor U11514 (N_11514,N_10879,N_11023);
or U11515 (N_11515,N_10959,N_10871);
or U11516 (N_11516,N_10669,N_10793);
xor U11517 (N_11517,N_10712,N_10646);
xnor U11518 (N_11518,N_10897,N_10780);
nor U11519 (N_11519,N_10579,N_11091);
nor U11520 (N_11520,N_10687,N_10565);
and U11521 (N_11521,N_11025,N_10982);
nor U11522 (N_11522,N_10997,N_10784);
and U11523 (N_11523,N_10905,N_10651);
and U11524 (N_11524,N_11215,N_10506);
or U11525 (N_11525,N_10813,N_11234);
and U11526 (N_11526,N_11032,N_10983);
nand U11527 (N_11527,N_10575,N_10822);
and U11528 (N_11528,N_10682,N_10628);
nand U11529 (N_11529,N_10702,N_10771);
or U11530 (N_11530,N_10749,N_10737);
nand U11531 (N_11531,N_11067,N_10708);
nand U11532 (N_11532,N_10713,N_10750);
nor U11533 (N_11533,N_10683,N_10965);
and U11534 (N_11534,N_10539,N_11053);
nand U11535 (N_11535,N_11131,N_11181);
nor U11536 (N_11536,N_11138,N_11191);
and U11537 (N_11537,N_11231,N_10903);
and U11538 (N_11538,N_10510,N_10661);
and U11539 (N_11539,N_10562,N_10505);
or U11540 (N_11540,N_10526,N_11242);
nor U11541 (N_11541,N_11160,N_10551);
xor U11542 (N_11542,N_11055,N_10885);
and U11543 (N_11543,N_10536,N_10943);
or U11544 (N_11544,N_10973,N_10837);
nor U11545 (N_11545,N_10859,N_11226);
nor U11546 (N_11546,N_10930,N_10556);
xor U11547 (N_11547,N_10694,N_10998);
nand U11548 (N_11548,N_10760,N_10739);
or U11549 (N_11549,N_11133,N_11239);
nor U11550 (N_11550,N_10685,N_11080);
nand U11551 (N_11551,N_10695,N_10922);
xnor U11552 (N_11552,N_11103,N_10589);
or U11553 (N_11553,N_11168,N_11050);
or U11554 (N_11554,N_11155,N_10898);
nand U11555 (N_11555,N_11061,N_10979);
nor U11556 (N_11556,N_11096,N_11059);
or U11557 (N_11557,N_11161,N_10592);
and U11558 (N_11558,N_10748,N_10504);
or U11559 (N_11559,N_11244,N_10567);
nand U11560 (N_11560,N_11135,N_10969);
and U11561 (N_11561,N_11007,N_10576);
and U11562 (N_11562,N_10795,N_11149);
nor U11563 (N_11563,N_11013,N_10961);
nand U11564 (N_11564,N_10907,N_10608);
xnor U11565 (N_11565,N_10511,N_11126);
and U11566 (N_11566,N_10547,N_11111);
xor U11567 (N_11567,N_10805,N_11150);
and U11568 (N_11568,N_11207,N_10632);
or U11569 (N_11569,N_10711,N_11122);
and U11570 (N_11570,N_10648,N_10620);
xnor U11571 (N_11571,N_11076,N_10644);
or U11572 (N_11572,N_10949,N_11183);
xor U11573 (N_11573,N_10785,N_10978);
nor U11574 (N_11574,N_10657,N_11098);
nor U11575 (N_11575,N_11167,N_11024);
nor U11576 (N_11576,N_10690,N_11073);
xor U11577 (N_11577,N_10844,N_11222);
xor U11578 (N_11578,N_10699,N_10972);
and U11579 (N_11579,N_11178,N_11197);
and U11580 (N_11580,N_11217,N_10826);
nor U11581 (N_11581,N_10558,N_11184);
nand U11582 (N_11582,N_10782,N_10883);
nand U11583 (N_11583,N_10726,N_11054);
nand U11584 (N_11584,N_10827,N_11086);
nand U11585 (N_11585,N_10666,N_10899);
or U11586 (N_11586,N_10716,N_11229);
or U11587 (N_11587,N_10816,N_10916);
or U11588 (N_11588,N_10786,N_11113);
nor U11589 (N_11589,N_10638,N_10768);
xnor U11590 (N_11590,N_11209,N_10668);
nand U11591 (N_11591,N_10730,N_10720);
nand U11592 (N_11592,N_11147,N_10751);
and U11593 (N_11593,N_11228,N_10744);
xor U11594 (N_11594,N_10691,N_10738);
xnor U11595 (N_11595,N_11175,N_10908);
nand U11596 (N_11596,N_10548,N_10948);
nand U11597 (N_11597,N_10581,N_10678);
or U11598 (N_11598,N_10647,N_10630);
nor U11599 (N_11599,N_10658,N_10557);
nor U11600 (N_11600,N_10612,N_11038);
xor U11601 (N_11601,N_10745,N_10566);
xnor U11602 (N_11602,N_11202,N_11163);
nor U11603 (N_11603,N_10721,N_10543);
nor U11604 (N_11604,N_11011,N_10591);
nand U11605 (N_11605,N_10831,N_10792);
and U11606 (N_11606,N_10719,N_11246);
nor U11607 (N_11607,N_10761,N_11220);
nand U11608 (N_11608,N_10799,N_11171);
or U11609 (N_11609,N_10808,N_11110);
nand U11610 (N_11610,N_10783,N_10570);
nand U11611 (N_11611,N_10990,N_11204);
and U11612 (N_11612,N_10618,N_10950);
nor U11613 (N_11613,N_10538,N_10958);
nand U11614 (N_11614,N_10811,N_10790);
xnor U11615 (N_11615,N_10984,N_10862);
xor U11616 (N_11616,N_10960,N_11097);
or U11617 (N_11617,N_10697,N_11119);
or U11618 (N_11618,N_10616,N_10860);
or U11619 (N_11619,N_10670,N_10693);
or U11620 (N_11620,N_10639,N_11066);
and U11621 (N_11621,N_10610,N_10824);
nor U11622 (N_11622,N_10919,N_11064);
nand U11623 (N_11623,N_10679,N_10654);
nand U11624 (N_11624,N_10820,N_11177);
nor U11625 (N_11625,N_11189,N_10915);
or U11626 (N_11626,N_10505,N_11085);
nor U11627 (N_11627,N_11007,N_10979);
or U11628 (N_11628,N_10744,N_10782);
xnor U11629 (N_11629,N_10570,N_11111);
xor U11630 (N_11630,N_10906,N_11028);
nor U11631 (N_11631,N_11199,N_11217);
xor U11632 (N_11632,N_10813,N_10778);
nand U11633 (N_11633,N_10630,N_11017);
or U11634 (N_11634,N_11022,N_10563);
nand U11635 (N_11635,N_10661,N_10601);
and U11636 (N_11636,N_10744,N_10839);
nand U11637 (N_11637,N_10902,N_10904);
nor U11638 (N_11638,N_10894,N_10548);
nor U11639 (N_11639,N_10808,N_10961);
xor U11640 (N_11640,N_10891,N_11119);
xor U11641 (N_11641,N_10929,N_10579);
nand U11642 (N_11642,N_10819,N_11165);
and U11643 (N_11643,N_11078,N_10941);
or U11644 (N_11644,N_10780,N_10767);
nand U11645 (N_11645,N_11003,N_10789);
and U11646 (N_11646,N_11026,N_10891);
or U11647 (N_11647,N_10940,N_11096);
nor U11648 (N_11648,N_10886,N_11043);
xnor U11649 (N_11649,N_10581,N_10877);
nor U11650 (N_11650,N_11245,N_10748);
nand U11651 (N_11651,N_10908,N_10839);
nand U11652 (N_11652,N_11181,N_10548);
and U11653 (N_11653,N_11105,N_10769);
nor U11654 (N_11654,N_10745,N_10588);
nand U11655 (N_11655,N_10985,N_10673);
nand U11656 (N_11656,N_10657,N_10514);
and U11657 (N_11657,N_10854,N_10544);
nand U11658 (N_11658,N_10727,N_10688);
nand U11659 (N_11659,N_10554,N_10872);
and U11660 (N_11660,N_10547,N_10642);
or U11661 (N_11661,N_11207,N_10938);
nor U11662 (N_11662,N_10595,N_10879);
nand U11663 (N_11663,N_10830,N_10676);
nand U11664 (N_11664,N_10689,N_10761);
and U11665 (N_11665,N_10724,N_11197);
or U11666 (N_11666,N_10598,N_10586);
nor U11667 (N_11667,N_10640,N_10730);
nand U11668 (N_11668,N_10730,N_10849);
nor U11669 (N_11669,N_10726,N_10537);
nand U11670 (N_11670,N_10868,N_10821);
nand U11671 (N_11671,N_10948,N_10758);
nor U11672 (N_11672,N_11211,N_10744);
nand U11673 (N_11673,N_11120,N_11208);
nand U11674 (N_11674,N_10744,N_10740);
nor U11675 (N_11675,N_10920,N_11045);
or U11676 (N_11676,N_10828,N_11046);
or U11677 (N_11677,N_11218,N_10794);
and U11678 (N_11678,N_11155,N_11190);
or U11679 (N_11679,N_10951,N_10966);
xor U11680 (N_11680,N_10648,N_10705);
xor U11681 (N_11681,N_10722,N_10659);
nand U11682 (N_11682,N_10674,N_10535);
and U11683 (N_11683,N_10892,N_10590);
or U11684 (N_11684,N_10634,N_10600);
nand U11685 (N_11685,N_11215,N_10544);
nor U11686 (N_11686,N_10685,N_10772);
and U11687 (N_11687,N_11142,N_10911);
xor U11688 (N_11688,N_10891,N_10763);
and U11689 (N_11689,N_11170,N_11082);
or U11690 (N_11690,N_10905,N_11176);
nand U11691 (N_11691,N_11210,N_11043);
and U11692 (N_11692,N_11170,N_10914);
or U11693 (N_11693,N_11154,N_11093);
nand U11694 (N_11694,N_11022,N_10629);
nand U11695 (N_11695,N_10687,N_10523);
or U11696 (N_11696,N_10561,N_10734);
nand U11697 (N_11697,N_10812,N_11131);
xnor U11698 (N_11698,N_11124,N_11108);
and U11699 (N_11699,N_11202,N_10754);
or U11700 (N_11700,N_10978,N_11232);
nor U11701 (N_11701,N_10550,N_10793);
and U11702 (N_11702,N_10624,N_10809);
and U11703 (N_11703,N_11134,N_10674);
xor U11704 (N_11704,N_10701,N_10835);
nand U11705 (N_11705,N_11111,N_11121);
or U11706 (N_11706,N_11190,N_10517);
xor U11707 (N_11707,N_11020,N_10550);
xnor U11708 (N_11708,N_11038,N_10895);
nand U11709 (N_11709,N_11179,N_11155);
nor U11710 (N_11710,N_11246,N_10953);
or U11711 (N_11711,N_10555,N_11230);
nor U11712 (N_11712,N_10954,N_11230);
nor U11713 (N_11713,N_10935,N_10847);
nor U11714 (N_11714,N_10623,N_10988);
nor U11715 (N_11715,N_10914,N_11009);
or U11716 (N_11716,N_10619,N_10812);
xor U11717 (N_11717,N_11116,N_11101);
nand U11718 (N_11718,N_10531,N_10654);
and U11719 (N_11719,N_10634,N_10558);
nor U11720 (N_11720,N_10978,N_10999);
and U11721 (N_11721,N_11024,N_10737);
xnor U11722 (N_11722,N_11136,N_10670);
xor U11723 (N_11723,N_10969,N_11211);
nand U11724 (N_11724,N_10694,N_10561);
and U11725 (N_11725,N_10611,N_10676);
or U11726 (N_11726,N_10739,N_10721);
nor U11727 (N_11727,N_11234,N_10660);
or U11728 (N_11728,N_10961,N_11236);
or U11729 (N_11729,N_11005,N_10637);
and U11730 (N_11730,N_11016,N_11070);
nor U11731 (N_11731,N_10657,N_10763);
and U11732 (N_11732,N_10512,N_10802);
nand U11733 (N_11733,N_11023,N_11230);
xnor U11734 (N_11734,N_10836,N_10966);
and U11735 (N_11735,N_11248,N_10856);
nor U11736 (N_11736,N_10831,N_10549);
nand U11737 (N_11737,N_10634,N_10670);
nor U11738 (N_11738,N_10837,N_10782);
and U11739 (N_11739,N_10507,N_11178);
and U11740 (N_11740,N_10842,N_10851);
or U11741 (N_11741,N_10703,N_11114);
or U11742 (N_11742,N_10746,N_10578);
or U11743 (N_11743,N_10533,N_10667);
and U11744 (N_11744,N_10849,N_10645);
xnor U11745 (N_11745,N_11192,N_11164);
xor U11746 (N_11746,N_11048,N_10881);
nand U11747 (N_11747,N_10855,N_10717);
and U11748 (N_11748,N_11098,N_10920);
and U11749 (N_11749,N_10561,N_10767);
nand U11750 (N_11750,N_11131,N_10875);
nor U11751 (N_11751,N_10673,N_11102);
nand U11752 (N_11752,N_11184,N_10783);
nand U11753 (N_11753,N_10777,N_10705);
nand U11754 (N_11754,N_11158,N_10936);
nand U11755 (N_11755,N_10521,N_10616);
nor U11756 (N_11756,N_10944,N_10656);
nor U11757 (N_11757,N_10982,N_10578);
or U11758 (N_11758,N_10789,N_10941);
xor U11759 (N_11759,N_10557,N_10944);
xor U11760 (N_11760,N_10656,N_10916);
and U11761 (N_11761,N_11121,N_10875);
nand U11762 (N_11762,N_10575,N_10962);
nor U11763 (N_11763,N_11214,N_11144);
nor U11764 (N_11764,N_11008,N_10536);
xnor U11765 (N_11765,N_11092,N_10724);
xor U11766 (N_11766,N_10745,N_11040);
nand U11767 (N_11767,N_10517,N_10615);
or U11768 (N_11768,N_10867,N_11091);
and U11769 (N_11769,N_10610,N_11194);
nand U11770 (N_11770,N_10876,N_10604);
or U11771 (N_11771,N_10914,N_10729);
or U11772 (N_11772,N_11143,N_10707);
xnor U11773 (N_11773,N_10966,N_10938);
and U11774 (N_11774,N_11108,N_10668);
xnor U11775 (N_11775,N_10817,N_10997);
or U11776 (N_11776,N_10527,N_10923);
xnor U11777 (N_11777,N_10720,N_10709);
nand U11778 (N_11778,N_10546,N_10553);
or U11779 (N_11779,N_10588,N_10841);
xor U11780 (N_11780,N_11009,N_11133);
nand U11781 (N_11781,N_10616,N_10739);
and U11782 (N_11782,N_10773,N_10800);
nor U11783 (N_11783,N_11035,N_10847);
and U11784 (N_11784,N_11169,N_11230);
and U11785 (N_11785,N_10868,N_10654);
nor U11786 (N_11786,N_11034,N_10647);
nand U11787 (N_11787,N_10616,N_11007);
or U11788 (N_11788,N_11219,N_10948);
nand U11789 (N_11789,N_10959,N_10821);
and U11790 (N_11790,N_10525,N_11056);
nand U11791 (N_11791,N_10787,N_11022);
nor U11792 (N_11792,N_11056,N_11024);
xor U11793 (N_11793,N_11215,N_11184);
nor U11794 (N_11794,N_10725,N_10932);
and U11795 (N_11795,N_11074,N_10598);
nor U11796 (N_11796,N_10866,N_11023);
xnor U11797 (N_11797,N_10581,N_10870);
nor U11798 (N_11798,N_10658,N_11009);
xnor U11799 (N_11799,N_11023,N_11001);
and U11800 (N_11800,N_10978,N_11047);
xnor U11801 (N_11801,N_10870,N_10675);
and U11802 (N_11802,N_10548,N_10714);
and U11803 (N_11803,N_11218,N_10853);
or U11804 (N_11804,N_11165,N_10970);
or U11805 (N_11805,N_10652,N_11104);
nor U11806 (N_11806,N_10563,N_10662);
xor U11807 (N_11807,N_10593,N_10733);
or U11808 (N_11808,N_10623,N_10796);
nand U11809 (N_11809,N_11093,N_10925);
and U11810 (N_11810,N_11173,N_10970);
xnor U11811 (N_11811,N_10795,N_10830);
nor U11812 (N_11812,N_10986,N_11121);
and U11813 (N_11813,N_10672,N_10606);
xnor U11814 (N_11814,N_11150,N_10763);
xnor U11815 (N_11815,N_10727,N_10607);
xor U11816 (N_11816,N_10774,N_11160);
or U11817 (N_11817,N_10643,N_11164);
nor U11818 (N_11818,N_10536,N_11090);
nand U11819 (N_11819,N_11159,N_10976);
xor U11820 (N_11820,N_11018,N_11174);
and U11821 (N_11821,N_11119,N_10966);
xor U11822 (N_11822,N_11047,N_10972);
nand U11823 (N_11823,N_11097,N_11122);
xor U11824 (N_11824,N_11206,N_10680);
nor U11825 (N_11825,N_10630,N_10703);
and U11826 (N_11826,N_11081,N_10723);
and U11827 (N_11827,N_11011,N_10807);
and U11828 (N_11828,N_10658,N_10987);
or U11829 (N_11829,N_11050,N_10904);
and U11830 (N_11830,N_11061,N_10515);
nand U11831 (N_11831,N_10549,N_10895);
and U11832 (N_11832,N_10513,N_11027);
nand U11833 (N_11833,N_11223,N_11011);
nor U11834 (N_11834,N_10839,N_11175);
xor U11835 (N_11835,N_10911,N_10503);
xnor U11836 (N_11836,N_10888,N_10639);
and U11837 (N_11837,N_10831,N_11029);
xor U11838 (N_11838,N_11212,N_10997);
and U11839 (N_11839,N_10730,N_11190);
and U11840 (N_11840,N_11056,N_10658);
or U11841 (N_11841,N_11158,N_10699);
nor U11842 (N_11842,N_10848,N_10522);
nor U11843 (N_11843,N_11028,N_10790);
or U11844 (N_11844,N_11017,N_11075);
or U11845 (N_11845,N_11131,N_10948);
or U11846 (N_11846,N_11096,N_10886);
nor U11847 (N_11847,N_11194,N_10912);
nor U11848 (N_11848,N_10800,N_10917);
xor U11849 (N_11849,N_11154,N_11184);
nand U11850 (N_11850,N_10882,N_10566);
nor U11851 (N_11851,N_10593,N_10820);
xor U11852 (N_11852,N_11034,N_11009);
and U11853 (N_11853,N_10584,N_10890);
nor U11854 (N_11854,N_10721,N_10784);
and U11855 (N_11855,N_10631,N_11104);
and U11856 (N_11856,N_11133,N_10746);
nor U11857 (N_11857,N_10703,N_10577);
nand U11858 (N_11858,N_11006,N_10502);
or U11859 (N_11859,N_10573,N_10955);
nand U11860 (N_11860,N_11205,N_11198);
xor U11861 (N_11861,N_10729,N_10677);
nor U11862 (N_11862,N_11015,N_10562);
nor U11863 (N_11863,N_10575,N_11105);
xnor U11864 (N_11864,N_11093,N_10595);
or U11865 (N_11865,N_10707,N_10640);
nor U11866 (N_11866,N_10995,N_10610);
or U11867 (N_11867,N_10522,N_10916);
and U11868 (N_11868,N_10839,N_10856);
nor U11869 (N_11869,N_10502,N_10974);
and U11870 (N_11870,N_10607,N_11182);
nor U11871 (N_11871,N_11195,N_10881);
and U11872 (N_11872,N_10528,N_10825);
nor U11873 (N_11873,N_10937,N_11248);
or U11874 (N_11874,N_11000,N_10857);
and U11875 (N_11875,N_10554,N_10530);
nand U11876 (N_11876,N_11072,N_10563);
and U11877 (N_11877,N_11134,N_10621);
and U11878 (N_11878,N_10508,N_11239);
nor U11879 (N_11879,N_10857,N_10863);
nand U11880 (N_11880,N_10601,N_10753);
nor U11881 (N_11881,N_10704,N_10614);
nand U11882 (N_11882,N_10703,N_10926);
nand U11883 (N_11883,N_10907,N_10657);
xnor U11884 (N_11884,N_10815,N_11050);
or U11885 (N_11885,N_10810,N_10947);
nor U11886 (N_11886,N_11214,N_11018);
or U11887 (N_11887,N_11220,N_10993);
and U11888 (N_11888,N_11221,N_11209);
nand U11889 (N_11889,N_10766,N_10836);
or U11890 (N_11890,N_10780,N_10761);
and U11891 (N_11891,N_10837,N_11117);
or U11892 (N_11892,N_11005,N_10815);
or U11893 (N_11893,N_10975,N_10511);
nor U11894 (N_11894,N_11000,N_11096);
and U11895 (N_11895,N_11207,N_10857);
or U11896 (N_11896,N_11099,N_11238);
xnor U11897 (N_11897,N_10794,N_10943);
xor U11898 (N_11898,N_10606,N_10773);
nor U11899 (N_11899,N_11208,N_10966);
nor U11900 (N_11900,N_11243,N_10872);
nand U11901 (N_11901,N_10774,N_11020);
nand U11902 (N_11902,N_10594,N_11008);
or U11903 (N_11903,N_10980,N_10998);
or U11904 (N_11904,N_10711,N_10706);
or U11905 (N_11905,N_10776,N_10987);
and U11906 (N_11906,N_10773,N_10793);
xnor U11907 (N_11907,N_10790,N_11001);
nand U11908 (N_11908,N_10734,N_10838);
and U11909 (N_11909,N_11201,N_11227);
nor U11910 (N_11910,N_10990,N_10608);
or U11911 (N_11911,N_10962,N_11155);
and U11912 (N_11912,N_11081,N_10749);
nor U11913 (N_11913,N_11005,N_10951);
nor U11914 (N_11914,N_11128,N_10617);
nor U11915 (N_11915,N_10518,N_11227);
and U11916 (N_11916,N_10753,N_11171);
or U11917 (N_11917,N_10505,N_11016);
nand U11918 (N_11918,N_10626,N_10652);
nand U11919 (N_11919,N_10830,N_10775);
and U11920 (N_11920,N_10778,N_10705);
nand U11921 (N_11921,N_10780,N_10839);
xor U11922 (N_11922,N_10625,N_10587);
xnor U11923 (N_11923,N_10920,N_11050);
or U11924 (N_11924,N_10745,N_10907);
nor U11925 (N_11925,N_10955,N_10986);
xor U11926 (N_11926,N_11134,N_10529);
xor U11927 (N_11927,N_10669,N_10688);
or U11928 (N_11928,N_10797,N_10703);
nand U11929 (N_11929,N_10683,N_10648);
and U11930 (N_11930,N_10663,N_11200);
nor U11931 (N_11931,N_11243,N_10922);
nor U11932 (N_11932,N_10821,N_11169);
nor U11933 (N_11933,N_10593,N_10666);
nand U11934 (N_11934,N_11186,N_10642);
and U11935 (N_11935,N_10852,N_10705);
nor U11936 (N_11936,N_11042,N_10731);
nand U11937 (N_11937,N_10913,N_11041);
or U11938 (N_11938,N_10995,N_10678);
or U11939 (N_11939,N_10641,N_11173);
nand U11940 (N_11940,N_11071,N_10874);
nor U11941 (N_11941,N_10547,N_10622);
nor U11942 (N_11942,N_11191,N_10651);
xor U11943 (N_11943,N_10903,N_10573);
xor U11944 (N_11944,N_10944,N_10765);
and U11945 (N_11945,N_10669,N_10800);
xor U11946 (N_11946,N_10565,N_10747);
or U11947 (N_11947,N_11064,N_11075);
nand U11948 (N_11948,N_10694,N_10576);
xor U11949 (N_11949,N_11249,N_11154);
nor U11950 (N_11950,N_10699,N_10778);
nand U11951 (N_11951,N_10821,N_11206);
and U11952 (N_11952,N_10765,N_10671);
xnor U11953 (N_11953,N_10560,N_11225);
xnor U11954 (N_11954,N_10851,N_10585);
or U11955 (N_11955,N_10649,N_11150);
or U11956 (N_11956,N_10875,N_10575);
and U11957 (N_11957,N_10524,N_10804);
nor U11958 (N_11958,N_11080,N_11050);
or U11959 (N_11959,N_10559,N_11081);
nand U11960 (N_11960,N_11191,N_11205);
and U11961 (N_11961,N_10633,N_10654);
or U11962 (N_11962,N_11186,N_10559);
nand U11963 (N_11963,N_10694,N_10581);
or U11964 (N_11964,N_11006,N_10550);
nand U11965 (N_11965,N_10770,N_10765);
xnor U11966 (N_11966,N_11220,N_11170);
nand U11967 (N_11967,N_10552,N_11246);
xnor U11968 (N_11968,N_10907,N_10741);
xor U11969 (N_11969,N_10753,N_10750);
xnor U11970 (N_11970,N_10706,N_10615);
nand U11971 (N_11971,N_10874,N_11111);
and U11972 (N_11972,N_10602,N_10667);
or U11973 (N_11973,N_10718,N_10821);
and U11974 (N_11974,N_11192,N_10536);
xor U11975 (N_11975,N_10859,N_11082);
or U11976 (N_11976,N_10592,N_10632);
xnor U11977 (N_11977,N_11145,N_11090);
or U11978 (N_11978,N_11157,N_11042);
xnor U11979 (N_11979,N_11223,N_11113);
nand U11980 (N_11980,N_10761,N_10703);
xor U11981 (N_11981,N_10622,N_11206);
xnor U11982 (N_11982,N_10510,N_10633);
xnor U11983 (N_11983,N_11061,N_10766);
and U11984 (N_11984,N_11040,N_10981);
nand U11985 (N_11985,N_10730,N_11177);
and U11986 (N_11986,N_10898,N_10682);
and U11987 (N_11987,N_10665,N_11231);
nand U11988 (N_11988,N_10741,N_10927);
or U11989 (N_11989,N_11012,N_10528);
nand U11990 (N_11990,N_10573,N_11196);
xnor U11991 (N_11991,N_10869,N_10928);
and U11992 (N_11992,N_10627,N_10725);
xnor U11993 (N_11993,N_10653,N_11182);
nor U11994 (N_11994,N_10711,N_11185);
xnor U11995 (N_11995,N_10521,N_11118);
nor U11996 (N_11996,N_10510,N_10914);
and U11997 (N_11997,N_11056,N_11005);
or U11998 (N_11998,N_10625,N_10520);
or U11999 (N_11999,N_10508,N_10600);
nor U12000 (N_12000,N_11838,N_11903);
nor U12001 (N_12001,N_11440,N_11557);
nand U12002 (N_12002,N_11467,N_11839);
xnor U12003 (N_12003,N_11757,N_11494);
nand U12004 (N_12004,N_11894,N_11796);
nor U12005 (N_12005,N_11549,N_11954);
and U12006 (N_12006,N_11898,N_11939);
nand U12007 (N_12007,N_11957,N_11329);
and U12008 (N_12008,N_11765,N_11819);
nor U12009 (N_12009,N_11743,N_11454);
xor U12010 (N_12010,N_11418,N_11463);
nand U12011 (N_12011,N_11410,N_11717);
nand U12012 (N_12012,N_11659,N_11930);
xor U12013 (N_12013,N_11813,N_11651);
and U12014 (N_12014,N_11584,N_11676);
nand U12015 (N_12015,N_11871,N_11453);
or U12016 (N_12016,N_11464,N_11994);
and U12017 (N_12017,N_11374,N_11369);
nor U12018 (N_12018,N_11967,N_11755);
and U12019 (N_12019,N_11594,N_11846);
and U12020 (N_12020,N_11751,N_11526);
nor U12021 (N_12021,N_11548,N_11272);
nand U12022 (N_12022,N_11344,N_11711);
and U12023 (N_12023,N_11426,N_11791);
xnor U12024 (N_12024,N_11466,N_11539);
xnor U12025 (N_12025,N_11722,N_11968);
or U12026 (N_12026,N_11696,N_11781);
or U12027 (N_12027,N_11390,N_11383);
or U12028 (N_12028,N_11270,N_11976);
and U12029 (N_12029,N_11942,N_11474);
nand U12030 (N_12030,N_11462,N_11820);
xnor U12031 (N_12031,N_11621,N_11405);
xor U12032 (N_12032,N_11480,N_11725);
nand U12033 (N_12033,N_11766,N_11856);
nor U12034 (N_12034,N_11890,N_11528);
or U12035 (N_12035,N_11392,N_11875);
xnor U12036 (N_12036,N_11919,N_11830);
or U12037 (N_12037,N_11475,N_11646);
or U12038 (N_12038,N_11497,N_11363);
and U12039 (N_12039,N_11878,N_11896);
and U12040 (N_12040,N_11654,N_11909);
and U12041 (N_12041,N_11858,N_11885);
and U12042 (N_12042,N_11753,N_11362);
nor U12043 (N_12043,N_11705,N_11565);
xnor U12044 (N_12044,N_11785,N_11451);
xnor U12045 (N_12045,N_11786,N_11343);
xor U12046 (N_12046,N_11733,N_11851);
or U12047 (N_12047,N_11541,N_11776);
and U12048 (N_12048,N_11862,N_11368);
nor U12049 (N_12049,N_11568,N_11759);
or U12050 (N_12050,N_11652,N_11700);
xor U12051 (N_12051,N_11936,N_11436);
nor U12052 (N_12052,N_11727,N_11385);
and U12053 (N_12053,N_11800,N_11970);
or U12054 (N_12054,N_11570,N_11938);
nor U12055 (N_12055,N_11997,N_11389);
nand U12056 (N_12056,N_11545,N_11556);
nand U12057 (N_12057,N_11459,N_11406);
or U12058 (N_12058,N_11310,N_11435);
and U12059 (N_12059,N_11394,N_11694);
xnor U12060 (N_12060,N_11470,N_11378);
nor U12061 (N_12061,N_11840,N_11790);
xor U12062 (N_12062,N_11419,N_11865);
or U12063 (N_12063,N_11981,N_11834);
nor U12064 (N_12064,N_11625,N_11905);
or U12065 (N_12065,N_11639,N_11973);
and U12066 (N_12066,N_11253,N_11407);
or U12067 (N_12067,N_11376,N_11281);
xnor U12068 (N_12068,N_11417,N_11724);
and U12069 (N_12069,N_11635,N_11305);
nand U12070 (N_12070,N_11443,N_11349);
or U12071 (N_12071,N_11876,N_11506);
nand U12072 (N_12072,N_11465,N_11802);
and U12073 (N_12073,N_11689,N_11914);
nand U12074 (N_12074,N_11461,N_11302);
and U12075 (N_12075,N_11500,N_11317);
nor U12076 (N_12076,N_11409,N_11354);
nor U12077 (N_12077,N_11874,N_11437);
nand U12078 (N_12078,N_11615,N_11931);
nand U12079 (N_12079,N_11699,N_11821);
xor U12080 (N_12080,N_11276,N_11300);
and U12081 (N_12081,N_11708,N_11313);
nor U12082 (N_12082,N_11256,N_11804);
and U12083 (N_12083,N_11948,N_11469);
nand U12084 (N_12084,N_11398,N_11596);
nand U12085 (N_12085,N_11514,N_11673);
or U12086 (N_12086,N_11684,N_11562);
nand U12087 (N_12087,N_11803,N_11932);
and U12088 (N_12088,N_11853,N_11325);
and U12089 (N_12089,N_11384,N_11925);
and U12090 (N_12090,N_11430,N_11799);
and U12091 (N_12091,N_11609,N_11775);
nand U12092 (N_12092,N_11663,N_11697);
nor U12093 (N_12093,N_11287,N_11262);
nor U12094 (N_12094,N_11411,N_11792);
and U12095 (N_12095,N_11702,N_11863);
nand U12096 (N_12096,N_11729,N_11788);
and U12097 (N_12097,N_11522,N_11380);
nand U12098 (N_12098,N_11636,N_11664);
or U12099 (N_12099,N_11665,N_11546);
and U12100 (N_12100,N_11706,N_11251);
nand U12101 (N_12101,N_11543,N_11685);
nand U12102 (N_12102,N_11558,N_11472);
xor U12103 (N_12103,N_11601,N_11943);
and U12104 (N_12104,N_11715,N_11597);
and U12105 (N_12105,N_11987,N_11333);
xor U12106 (N_12106,N_11534,N_11946);
nor U12107 (N_12107,N_11319,N_11628);
or U12108 (N_12108,N_11739,N_11855);
xnor U12109 (N_12109,N_11415,N_11688);
or U12110 (N_12110,N_11575,N_11616);
or U12111 (N_12111,N_11823,N_11686);
or U12112 (N_12112,N_11810,N_11624);
nor U12113 (N_12113,N_11330,N_11872);
nor U12114 (N_12114,N_11586,N_11986);
nand U12115 (N_12115,N_11769,N_11709);
or U12116 (N_12116,N_11529,N_11752);
xor U12117 (N_12117,N_11393,N_11585);
and U12118 (N_12118,N_11395,N_11842);
or U12119 (N_12119,N_11250,N_11476);
nand U12120 (N_12120,N_11952,N_11701);
nor U12121 (N_12121,N_11666,N_11648);
and U12122 (N_12122,N_11927,N_11990);
nand U12123 (N_12123,N_11761,N_11365);
xor U12124 (N_12124,N_11959,N_11582);
and U12125 (N_12125,N_11814,N_11303);
xor U12126 (N_12126,N_11531,N_11295);
nand U12127 (N_12127,N_11749,N_11589);
or U12128 (N_12128,N_11487,N_11947);
xor U12129 (N_12129,N_11563,N_11397);
xor U12130 (N_12130,N_11844,N_11297);
nor U12131 (N_12131,N_11593,N_11483);
xor U12132 (N_12132,N_11351,N_11587);
xnor U12133 (N_12133,N_11951,N_11737);
nor U12134 (N_12134,N_11672,N_11771);
nand U12135 (N_12135,N_11446,N_11353);
xnor U12136 (N_12136,N_11518,N_11292);
or U12137 (N_12137,N_11493,N_11818);
xor U12138 (N_12138,N_11371,N_11763);
xnor U12139 (N_12139,N_11566,N_11261);
nor U12140 (N_12140,N_11502,N_11716);
and U12141 (N_12141,N_11316,N_11772);
nor U12142 (N_12142,N_11267,N_11561);
nor U12143 (N_12143,N_11963,N_11540);
nand U12144 (N_12144,N_11504,N_11832);
nand U12145 (N_12145,N_11883,N_11598);
and U12146 (N_12146,N_11895,N_11795);
or U12147 (N_12147,N_11857,N_11404);
xnor U12148 (N_12148,N_11797,N_11906);
nor U12149 (N_12149,N_11600,N_11798);
xnor U12150 (N_12150,N_11693,N_11745);
xor U12151 (N_12151,N_11320,N_11728);
xor U12152 (N_12152,N_11843,N_11632);
nor U12153 (N_12153,N_11252,N_11793);
nand U12154 (N_12154,N_11692,N_11547);
nor U12155 (N_12155,N_11294,N_11377);
and U12156 (N_12156,N_11860,N_11399);
nor U12157 (N_12157,N_11690,N_11762);
and U12158 (N_12158,N_11519,N_11817);
xnor U12159 (N_12159,N_11520,N_11622);
xnor U12160 (N_12160,N_11327,N_11660);
nand U12161 (N_12161,N_11731,N_11386);
xnor U12162 (N_12162,N_11884,N_11841);
or U12163 (N_12163,N_11640,N_11278);
nand U12164 (N_12164,N_11388,N_11675);
nand U12165 (N_12165,N_11880,N_11311);
and U12166 (N_12166,N_11611,N_11495);
and U12167 (N_12167,N_11460,N_11695);
and U12168 (N_12168,N_11760,N_11859);
nor U12169 (N_12169,N_11503,N_11698);
or U12170 (N_12170,N_11828,N_11805);
and U12171 (N_12171,N_11301,N_11431);
or U12172 (N_12172,N_11989,N_11551);
or U12173 (N_12173,N_11998,N_11555);
nand U12174 (N_12174,N_11870,N_11630);
and U12175 (N_12175,N_11811,N_11535);
nor U12176 (N_12176,N_11269,N_11413);
nor U12177 (N_12177,N_11271,N_11641);
nor U12178 (N_12178,N_11360,N_11682);
and U12179 (N_12179,N_11553,N_11361);
nor U12180 (N_12180,N_11336,N_11758);
and U12181 (N_12181,N_11434,N_11649);
xor U12182 (N_12182,N_11421,N_11726);
and U12183 (N_12183,N_11279,N_11783);
xnor U12184 (N_12184,N_11356,N_11642);
or U12185 (N_12185,N_11991,N_11835);
nand U12186 (N_12186,N_11707,N_11736);
xnor U12187 (N_12187,N_11339,N_11512);
xor U12188 (N_12188,N_11687,N_11816);
or U12189 (N_12189,N_11658,N_11933);
or U12190 (N_12190,N_11770,N_11444);
nor U12191 (N_12191,N_11254,N_11741);
nand U12192 (N_12192,N_11370,N_11629);
or U12193 (N_12193,N_11414,N_11794);
xnor U12194 (N_12194,N_11920,N_11911);
or U12195 (N_12195,N_11908,N_11321);
xnor U12196 (N_12196,N_11445,N_11789);
xnor U12197 (N_12197,N_11573,N_11581);
and U12198 (N_12198,N_11975,N_11979);
nor U12199 (N_12199,N_11677,N_11602);
and U12200 (N_12200,N_11940,N_11985);
nand U12201 (N_12201,N_11536,N_11929);
or U12202 (N_12202,N_11877,N_11427);
and U12203 (N_12203,N_11273,N_11260);
xor U12204 (N_12204,N_11286,N_11507);
nor U12205 (N_12205,N_11485,N_11774);
nor U12206 (N_12206,N_11777,N_11852);
nand U12207 (N_12207,N_11479,N_11671);
nor U12208 (N_12208,N_11825,N_11678);
nor U12209 (N_12209,N_11901,N_11669);
or U12210 (N_12210,N_11498,N_11918);
xnor U12211 (N_12211,N_11433,N_11482);
or U12212 (N_12212,N_11481,N_11449);
nand U12213 (N_12213,N_11645,N_11289);
nand U12214 (N_12214,N_11787,N_11620);
nor U12215 (N_12215,N_11734,N_11868);
nor U12216 (N_12216,N_11505,N_11450);
and U12217 (N_12217,N_11264,N_11599);
xor U12218 (N_12218,N_11879,N_11255);
and U12219 (N_12219,N_11366,N_11403);
and U12220 (N_12220,N_11348,N_11424);
xnor U12221 (N_12221,N_11337,N_11338);
xor U12222 (N_12222,N_11899,N_11744);
and U12223 (N_12223,N_11357,N_11691);
nand U12224 (N_12224,N_11661,N_11928);
nor U12225 (N_12225,N_11471,N_11552);
and U12226 (N_12226,N_11773,N_11326);
and U12227 (N_12227,N_11559,N_11972);
nor U12228 (N_12228,N_11275,N_11263);
nand U12229 (N_12229,N_11710,N_11680);
or U12230 (N_12230,N_11304,N_11416);
nor U12231 (N_12231,N_11809,N_11779);
or U12232 (N_12232,N_11937,N_11854);
nand U12233 (N_12233,N_11882,N_11334);
xnor U12234 (N_12234,N_11647,N_11283);
xor U12235 (N_12235,N_11496,N_11992);
xnor U12236 (N_12236,N_11439,N_11342);
xnor U12237 (N_12237,N_11274,N_11754);
or U12238 (N_12238,N_11867,N_11308);
and U12239 (N_12239,N_11668,N_11412);
nor U12240 (N_12240,N_11532,N_11574);
nand U12241 (N_12241,N_11468,N_11740);
nor U12242 (N_12242,N_11447,N_11259);
nor U12243 (N_12243,N_11341,N_11523);
nand U12244 (N_12244,N_11291,N_11923);
xnor U12245 (N_12245,N_11257,N_11517);
or U12246 (N_12246,N_11950,N_11554);
or U12247 (N_12247,N_11429,N_11812);
xor U12248 (N_12248,N_11966,N_11969);
or U12249 (N_12249,N_11346,N_11610);
or U12250 (N_12250,N_11627,N_11623);
nor U12251 (N_12251,N_11735,N_11511);
or U12252 (N_12252,N_11993,N_11323);
or U12253 (N_12253,N_11605,N_11538);
nand U12254 (N_12254,N_11352,N_11355);
nand U12255 (N_12255,N_11299,N_11836);
nand U12256 (N_12256,N_11530,N_11941);
nand U12257 (N_12257,N_11917,N_11533);
or U12258 (N_12258,N_11962,N_11924);
nand U12259 (N_12259,N_11367,N_11747);
nor U12260 (N_12260,N_11347,N_11400);
nor U12261 (N_12261,N_11432,N_11527);
nand U12262 (N_12262,N_11679,N_11888);
nor U12263 (N_12263,N_11569,N_11606);
nand U12264 (N_12264,N_11644,N_11509);
nand U12265 (N_12265,N_11478,N_11980);
xor U12266 (N_12266,N_11550,N_11332);
xor U12267 (N_12267,N_11491,N_11730);
or U12268 (N_12268,N_11815,N_11714);
nor U12269 (N_12269,N_11490,N_11588);
xnor U12270 (N_12270,N_11704,N_11662);
and U12271 (N_12271,N_11750,N_11655);
and U12272 (N_12272,N_11501,N_11583);
nor U12273 (N_12273,N_11309,N_11258);
and U12274 (N_12274,N_11742,N_11571);
nand U12275 (N_12275,N_11340,N_11379);
xor U12276 (N_12276,N_11955,N_11542);
nor U12277 (N_12277,N_11848,N_11983);
nor U12278 (N_12278,N_11977,N_11608);
nor U12279 (N_12279,N_11322,N_11891);
and U12280 (N_12280,N_11721,N_11827);
nor U12281 (N_12281,N_11387,N_11956);
and U12282 (N_12282,N_11960,N_11907);
or U12283 (N_12283,N_11808,N_11359);
xor U12284 (N_12284,N_11614,N_11382);
xor U12285 (N_12285,N_11350,N_11723);
nand U12286 (N_12286,N_11784,N_11458);
nand U12287 (N_12287,N_11964,N_11881);
and U12288 (N_12288,N_11580,N_11978);
and U12289 (N_12289,N_11576,N_11422);
and U12290 (N_12290,N_11280,N_11372);
xor U12291 (N_12291,N_11293,N_11277);
nor U12292 (N_12292,N_11612,N_11634);
or U12293 (N_12293,N_11578,N_11513);
nand U12294 (N_12294,N_11613,N_11674);
or U12295 (N_12295,N_11579,N_11958);
xnor U12296 (N_12296,N_11448,N_11656);
nand U12297 (N_12297,N_11780,N_11306);
nand U12298 (N_12298,N_11265,N_11971);
and U12299 (N_12299,N_11849,N_11886);
nor U12300 (N_12300,N_11893,N_11650);
or U12301 (N_12301,N_11944,N_11484);
nor U12302 (N_12302,N_11375,N_11607);
or U12303 (N_12303,N_11457,N_11298);
xor U12304 (N_12304,N_11913,N_11489);
nand U12305 (N_12305,N_11525,N_11910);
xnor U12306 (N_12306,N_11455,N_11829);
nor U12307 (N_12307,N_11683,N_11515);
and U12308 (N_12308,N_11510,N_11892);
or U12309 (N_12309,N_11831,N_11767);
xor U12310 (N_12310,N_11900,N_11953);
and U12311 (N_12311,N_11288,N_11845);
nor U12312 (N_12312,N_11560,N_11373);
or U12313 (N_12313,N_11764,N_11984);
nand U12314 (N_12314,N_11401,N_11364);
nor U12315 (N_12315,N_11887,N_11996);
xor U12316 (N_12316,N_11324,N_11402);
and U12317 (N_12317,N_11420,N_11328);
and U12318 (N_12318,N_11314,N_11738);
and U12319 (N_12319,N_11391,N_11423);
or U12320 (N_12320,N_11902,N_11284);
and U12321 (N_12321,N_11748,N_11837);
xnor U12322 (N_12322,N_11516,N_11591);
nand U12323 (N_12323,N_11861,N_11486);
nor U12324 (N_12324,N_11806,N_11441);
nor U12325 (N_12325,N_11603,N_11266);
and U12326 (N_12326,N_11961,N_11473);
nand U12327 (N_12327,N_11521,N_11756);
xnor U12328 (N_12328,N_11619,N_11873);
and U12329 (N_12329,N_11567,N_11408);
nand U12330 (N_12330,N_11782,N_11312);
nor U12331 (N_12331,N_11866,N_11626);
or U12332 (N_12332,N_11912,N_11703);
or U12333 (N_12333,N_11847,N_11618);
or U12334 (N_12334,N_11982,N_11999);
nor U12335 (N_12335,N_11438,N_11657);
xor U12336 (N_12336,N_11670,N_11801);
nand U12337 (N_12337,N_11282,N_11577);
xor U12338 (N_12338,N_11922,N_11916);
nor U12339 (N_12339,N_11719,N_11331);
nand U12340 (N_12340,N_11572,N_11643);
and U12341 (N_12341,N_11335,N_11477);
and U12342 (N_12342,N_11488,N_11296);
and U12343 (N_12343,N_11592,N_11889);
nor U12344 (N_12344,N_11712,N_11564);
nand U12345 (N_12345,N_11826,N_11442);
nor U12346 (N_12346,N_11456,N_11864);
nor U12347 (N_12347,N_11824,N_11949);
nor U12348 (N_12348,N_11307,N_11396);
nor U12349 (N_12349,N_11508,N_11428);
or U12350 (N_12350,N_11897,N_11988);
nor U12351 (N_12351,N_11524,N_11807);
nand U12352 (N_12352,N_11713,N_11921);
nor U12353 (N_12353,N_11850,N_11544);
nand U12354 (N_12354,N_11833,N_11974);
nor U12355 (N_12355,N_11345,N_11778);
or U12356 (N_12356,N_11631,N_11318);
or U12357 (N_12357,N_11425,N_11285);
nor U12358 (N_12358,N_11768,N_11945);
and U12359 (N_12359,N_11381,N_11681);
nand U12360 (N_12360,N_11935,N_11358);
or U12361 (N_12361,N_11633,N_11315);
xor U12362 (N_12362,N_11638,N_11926);
xnor U12363 (N_12363,N_11965,N_11452);
nor U12364 (N_12364,N_11537,N_11718);
nand U12365 (N_12365,N_11995,N_11934);
nand U12366 (N_12366,N_11617,N_11720);
nor U12367 (N_12367,N_11604,N_11653);
nor U12368 (N_12368,N_11268,N_11499);
or U12369 (N_12369,N_11492,N_11746);
nor U12370 (N_12370,N_11904,N_11869);
or U12371 (N_12371,N_11732,N_11590);
and U12372 (N_12372,N_11595,N_11667);
nor U12373 (N_12373,N_11822,N_11290);
nor U12374 (N_12374,N_11637,N_11915);
and U12375 (N_12375,N_11373,N_11464);
or U12376 (N_12376,N_11589,N_11601);
nor U12377 (N_12377,N_11362,N_11998);
or U12378 (N_12378,N_11569,N_11717);
nor U12379 (N_12379,N_11255,N_11491);
nand U12380 (N_12380,N_11800,N_11470);
nand U12381 (N_12381,N_11854,N_11312);
nand U12382 (N_12382,N_11275,N_11577);
nor U12383 (N_12383,N_11348,N_11577);
and U12384 (N_12384,N_11655,N_11305);
nor U12385 (N_12385,N_11794,N_11957);
xor U12386 (N_12386,N_11539,N_11869);
xnor U12387 (N_12387,N_11780,N_11389);
nor U12388 (N_12388,N_11812,N_11551);
nor U12389 (N_12389,N_11401,N_11460);
nand U12390 (N_12390,N_11593,N_11900);
nand U12391 (N_12391,N_11802,N_11734);
or U12392 (N_12392,N_11637,N_11611);
and U12393 (N_12393,N_11294,N_11821);
and U12394 (N_12394,N_11593,N_11638);
xor U12395 (N_12395,N_11844,N_11363);
nand U12396 (N_12396,N_11815,N_11807);
and U12397 (N_12397,N_11914,N_11940);
and U12398 (N_12398,N_11927,N_11759);
or U12399 (N_12399,N_11579,N_11385);
and U12400 (N_12400,N_11961,N_11487);
and U12401 (N_12401,N_11497,N_11500);
and U12402 (N_12402,N_11628,N_11541);
or U12403 (N_12403,N_11284,N_11624);
nand U12404 (N_12404,N_11780,N_11526);
nand U12405 (N_12405,N_11450,N_11745);
or U12406 (N_12406,N_11694,N_11329);
nor U12407 (N_12407,N_11702,N_11590);
nand U12408 (N_12408,N_11740,N_11570);
or U12409 (N_12409,N_11359,N_11255);
xor U12410 (N_12410,N_11807,N_11711);
and U12411 (N_12411,N_11916,N_11446);
xor U12412 (N_12412,N_11870,N_11277);
nor U12413 (N_12413,N_11812,N_11669);
nand U12414 (N_12414,N_11769,N_11757);
xor U12415 (N_12415,N_11846,N_11905);
xor U12416 (N_12416,N_11398,N_11369);
and U12417 (N_12417,N_11983,N_11851);
or U12418 (N_12418,N_11472,N_11491);
and U12419 (N_12419,N_11671,N_11560);
nand U12420 (N_12420,N_11707,N_11776);
nand U12421 (N_12421,N_11459,N_11326);
and U12422 (N_12422,N_11509,N_11682);
nor U12423 (N_12423,N_11843,N_11783);
and U12424 (N_12424,N_11655,N_11851);
and U12425 (N_12425,N_11857,N_11632);
xnor U12426 (N_12426,N_11815,N_11425);
xnor U12427 (N_12427,N_11616,N_11625);
and U12428 (N_12428,N_11459,N_11538);
or U12429 (N_12429,N_11369,N_11364);
xor U12430 (N_12430,N_11790,N_11335);
nor U12431 (N_12431,N_11425,N_11523);
and U12432 (N_12432,N_11531,N_11443);
and U12433 (N_12433,N_11466,N_11964);
nand U12434 (N_12434,N_11266,N_11413);
or U12435 (N_12435,N_11949,N_11754);
nand U12436 (N_12436,N_11430,N_11999);
xor U12437 (N_12437,N_11806,N_11722);
nand U12438 (N_12438,N_11854,N_11669);
nand U12439 (N_12439,N_11949,N_11758);
xnor U12440 (N_12440,N_11952,N_11568);
nor U12441 (N_12441,N_11742,N_11549);
or U12442 (N_12442,N_11675,N_11917);
xor U12443 (N_12443,N_11755,N_11906);
nor U12444 (N_12444,N_11555,N_11406);
or U12445 (N_12445,N_11907,N_11323);
nand U12446 (N_12446,N_11518,N_11912);
nand U12447 (N_12447,N_11604,N_11491);
nor U12448 (N_12448,N_11429,N_11261);
or U12449 (N_12449,N_11478,N_11841);
nor U12450 (N_12450,N_11915,N_11606);
nand U12451 (N_12451,N_11942,N_11956);
or U12452 (N_12452,N_11688,N_11358);
nand U12453 (N_12453,N_11438,N_11541);
xor U12454 (N_12454,N_11617,N_11998);
and U12455 (N_12455,N_11544,N_11830);
nand U12456 (N_12456,N_11593,N_11644);
nor U12457 (N_12457,N_11535,N_11980);
or U12458 (N_12458,N_11934,N_11867);
and U12459 (N_12459,N_11768,N_11875);
nor U12460 (N_12460,N_11424,N_11268);
or U12461 (N_12461,N_11968,N_11345);
nand U12462 (N_12462,N_11277,N_11420);
nand U12463 (N_12463,N_11447,N_11615);
xor U12464 (N_12464,N_11712,N_11275);
xnor U12465 (N_12465,N_11496,N_11861);
or U12466 (N_12466,N_11789,N_11466);
nand U12467 (N_12467,N_11277,N_11967);
nor U12468 (N_12468,N_11604,N_11906);
and U12469 (N_12469,N_11483,N_11512);
xor U12470 (N_12470,N_11488,N_11452);
or U12471 (N_12471,N_11846,N_11870);
nor U12472 (N_12472,N_11381,N_11847);
nor U12473 (N_12473,N_11288,N_11979);
xnor U12474 (N_12474,N_11454,N_11666);
or U12475 (N_12475,N_11788,N_11968);
xnor U12476 (N_12476,N_11913,N_11533);
xnor U12477 (N_12477,N_11499,N_11880);
or U12478 (N_12478,N_11920,N_11615);
or U12479 (N_12479,N_11397,N_11964);
nor U12480 (N_12480,N_11524,N_11369);
and U12481 (N_12481,N_11901,N_11924);
nor U12482 (N_12482,N_11259,N_11405);
or U12483 (N_12483,N_11691,N_11487);
or U12484 (N_12484,N_11477,N_11934);
and U12485 (N_12485,N_11911,N_11707);
or U12486 (N_12486,N_11460,N_11720);
and U12487 (N_12487,N_11863,N_11354);
nor U12488 (N_12488,N_11650,N_11483);
and U12489 (N_12489,N_11638,N_11886);
nor U12490 (N_12490,N_11717,N_11652);
nand U12491 (N_12491,N_11265,N_11308);
xor U12492 (N_12492,N_11914,N_11328);
and U12493 (N_12493,N_11482,N_11682);
and U12494 (N_12494,N_11330,N_11967);
nand U12495 (N_12495,N_11354,N_11520);
nand U12496 (N_12496,N_11499,N_11720);
xnor U12497 (N_12497,N_11558,N_11614);
nand U12498 (N_12498,N_11458,N_11429);
xnor U12499 (N_12499,N_11786,N_11888);
nand U12500 (N_12500,N_11882,N_11935);
nor U12501 (N_12501,N_11421,N_11601);
nand U12502 (N_12502,N_11914,N_11735);
xnor U12503 (N_12503,N_11452,N_11589);
nand U12504 (N_12504,N_11796,N_11771);
nand U12505 (N_12505,N_11407,N_11367);
nand U12506 (N_12506,N_11254,N_11690);
or U12507 (N_12507,N_11254,N_11549);
and U12508 (N_12508,N_11722,N_11884);
nor U12509 (N_12509,N_11906,N_11640);
nand U12510 (N_12510,N_11612,N_11799);
nor U12511 (N_12511,N_11733,N_11659);
nor U12512 (N_12512,N_11287,N_11294);
and U12513 (N_12513,N_11889,N_11942);
nand U12514 (N_12514,N_11705,N_11331);
xnor U12515 (N_12515,N_11972,N_11776);
and U12516 (N_12516,N_11809,N_11387);
or U12517 (N_12517,N_11473,N_11834);
or U12518 (N_12518,N_11778,N_11739);
xor U12519 (N_12519,N_11281,N_11864);
or U12520 (N_12520,N_11718,N_11373);
or U12521 (N_12521,N_11617,N_11681);
or U12522 (N_12522,N_11550,N_11641);
or U12523 (N_12523,N_11482,N_11509);
xor U12524 (N_12524,N_11347,N_11341);
or U12525 (N_12525,N_11338,N_11956);
nand U12526 (N_12526,N_11838,N_11455);
xor U12527 (N_12527,N_11794,N_11793);
nand U12528 (N_12528,N_11682,N_11770);
nand U12529 (N_12529,N_11285,N_11730);
or U12530 (N_12530,N_11447,N_11957);
nand U12531 (N_12531,N_11831,N_11437);
nand U12532 (N_12532,N_11760,N_11908);
or U12533 (N_12533,N_11928,N_11906);
nor U12534 (N_12534,N_11384,N_11705);
nor U12535 (N_12535,N_11490,N_11392);
nand U12536 (N_12536,N_11688,N_11621);
or U12537 (N_12537,N_11714,N_11334);
or U12538 (N_12538,N_11992,N_11972);
nor U12539 (N_12539,N_11435,N_11441);
and U12540 (N_12540,N_11733,N_11324);
or U12541 (N_12541,N_11363,N_11825);
nand U12542 (N_12542,N_11900,N_11594);
xor U12543 (N_12543,N_11718,N_11386);
or U12544 (N_12544,N_11431,N_11943);
or U12545 (N_12545,N_11518,N_11622);
nor U12546 (N_12546,N_11677,N_11908);
nand U12547 (N_12547,N_11279,N_11839);
or U12548 (N_12548,N_11320,N_11871);
xor U12549 (N_12549,N_11570,N_11826);
or U12550 (N_12550,N_11525,N_11504);
and U12551 (N_12551,N_11957,N_11639);
nor U12552 (N_12552,N_11591,N_11843);
or U12553 (N_12553,N_11648,N_11434);
nor U12554 (N_12554,N_11997,N_11325);
nand U12555 (N_12555,N_11911,N_11643);
nand U12556 (N_12556,N_11761,N_11768);
nand U12557 (N_12557,N_11533,N_11304);
xnor U12558 (N_12558,N_11287,N_11430);
or U12559 (N_12559,N_11858,N_11647);
xor U12560 (N_12560,N_11486,N_11432);
nand U12561 (N_12561,N_11385,N_11512);
and U12562 (N_12562,N_11273,N_11834);
or U12563 (N_12563,N_11856,N_11887);
nand U12564 (N_12564,N_11571,N_11840);
xor U12565 (N_12565,N_11352,N_11601);
and U12566 (N_12566,N_11255,N_11948);
nor U12567 (N_12567,N_11896,N_11623);
nor U12568 (N_12568,N_11272,N_11595);
nand U12569 (N_12569,N_11442,N_11733);
and U12570 (N_12570,N_11282,N_11837);
nor U12571 (N_12571,N_11322,N_11859);
nand U12572 (N_12572,N_11314,N_11914);
and U12573 (N_12573,N_11963,N_11827);
nor U12574 (N_12574,N_11700,N_11287);
nand U12575 (N_12575,N_11935,N_11944);
nor U12576 (N_12576,N_11821,N_11706);
and U12577 (N_12577,N_11645,N_11332);
xnor U12578 (N_12578,N_11743,N_11686);
nand U12579 (N_12579,N_11648,N_11851);
nor U12580 (N_12580,N_11432,N_11625);
nor U12581 (N_12581,N_11911,N_11285);
nor U12582 (N_12582,N_11726,N_11625);
or U12583 (N_12583,N_11557,N_11405);
and U12584 (N_12584,N_11558,N_11952);
nand U12585 (N_12585,N_11555,N_11543);
nor U12586 (N_12586,N_11968,N_11433);
or U12587 (N_12587,N_11865,N_11384);
and U12588 (N_12588,N_11558,N_11953);
nor U12589 (N_12589,N_11685,N_11360);
or U12590 (N_12590,N_11667,N_11458);
xnor U12591 (N_12591,N_11780,N_11537);
xnor U12592 (N_12592,N_11884,N_11437);
or U12593 (N_12593,N_11866,N_11516);
nand U12594 (N_12594,N_11302,N_11846);
and U12595 (N_12595,N_11302,N_11500);
nand U12596 (N_12596,N_11882,N_11592);
and U12597 (N_12597,N_11499,N_11997);
nand U12598 (N_12598,N_11885,N_11812);
and U12599 (N_12599,N_11734,N_11641);
and U12600 (N_12600,N_11597,N_11991);
nand U12601 (N_12601,N_11444,N_11316);
nand U12602 (N_12602,N_11857,N_11866);
nand U12603 (N_12603,N_11463,N_11979);
nor U12604 (N_12604,N_11548,N_11504);
nand U12605 (N_12605,N_11620,N_11531);
and U12606 (N_12606,N_11734,N_11603);
xor U12607 (N_12607,N_11635,N_11375);
and U12608 (N_12608,N_11337,N_11322);
and U12609 (N_12609,N_11538,N_11681);
nand U12610 (N_12610,N_11383,N_11534);
nor U12611 (N_12611,N_11536,N_11334);
nand U12612 (N_12612,N_11940,N_11724);
or U12613 (N_12613,N_11680,N_11910);
nor U12614 (N_12614,N_11269,N_11965);
xor U12615 (N_12615,N_11337,N_11932);
nand U12616 (N_12616,N_11491,N_11712);
or U12617 (N_12617,N_11519,N_11911);
xor U12618 (N_12618,N_11686,N_11367);
xor U12619 (N_12619,N_11465,N_11927);
and U12620 (N_12620,N_11660,N_11563);
and U12621 (N_12621,N_11356,N_11809);
nand U12622 (N_12622,N_11662,N_11575);
xor U12623 (N_12623,N_11906,N_11371);
or U12624 (N_12624,N_11789,N_11679);
and U12625 (N_12625,N_11635,N_11654);
or U12626 (N_12626,N_11413,N_11606);
xor U12627 (N_12627,N_11270,N_11318);
nor U12628 (N_12628,N_11558,N_11894);
nor U12629 (N_12629,N_11848,N_11905);
xnor U12630 (N_12630,N_11959,N_11924);
xnor U12631 (N_12631,N_11419,N_11996);
nor U12632 (N_12632,N_11968,N_11475);
nand U12633 (N_12633,N_11479,N_11315);
nand U12634 (N_12634,N_11271,N_11431);
and U12635 (N_12635,N_11585,N_11807);
and U12636 (N_12636,N_11938,N_11412);
and U12637 (N_12637,N_11965,N_11683);
xnor U12638 (N_12638,N_11449,N_11973);
xor U12639 (N_12639,N_11769,N_11529);
nor U12640 (N_12640,N_11405,N_11276);
and U12641 (N_12641,N_11482,N_11733);
nor U12642 (N_12642,N_11590,N_11459);
nand U12643 (N_12643,N_11547,N_11720);
and U12644 (N_12644,N_11432,N_11681);
nor U12645 (N_12645,N_11933,N_11935);
nand U12646 (N_12646,N_11453,N_11491);
and U12647 (N_12647,N_11341,N_11715);
nor U12648 (N_12648,N_11819,N_11636);
or U12649 (N_12649,N_11519,N_11884);
nand U12650 (N_12650,N_11919,N_11251);
and U12651 (N_12651,N_11605,N_11712);
or U12652 (N_12652,N_11546,N_11461);
xor U12653 (N_12653,N_11921,N_11494);
or U12654 (N_12654,N_11428,N_11682);
xnor U12655 (N_12655,N_11403,N_11282);
and U12656 (N_12656,N_11514,N_11769);
xor U12657 (N_12657,N_11295,N_11774);
or U12658 (N_12658,N_11366,N_11342);
xor U12659 (N_12659,N_11601,N_11714);
xnor U12660 (N_12660,N_11415,N_11863);
or U12661 (N_12661,N_11271,N_11950);
nand U12662 (N_12662,N_11896,N_11879);
and U12663 (N_12663,N_11904,N_11469);
or U12664 (N_12664,N_11672,N_11694);
or U12665 (N_12665,N_11458,N_11542);
and U12666 (N_12666,N_11256,N_11715);
or U12667 (N_12667,N_11950,N_11453);
xor U12668 (N_12668,N_11921,N_11800);
and U12669 (N_12669,N_11572,N_11375);
nor U12670 (N_12670,N_11968,N_11872);
or U12671 (N_12671,N_11789,N_11536);
xor U12672 (N_12672,N_11655,N_11695);
nand U12673 (N_12673,N_11701,N_11738);
nor U12674 (N_12674,N_11529,N_11503);
nand U12675 (N_12675,N_11421,N_11555);
xnor U12676 (N_12676,N_11341,N_11556);
xnor U12677 (N_12677,N_11683,N_11901);
or U12678 (N_12678,N_11434,N_11253);
nand U12679 (N_12679,N_11652,N_11559);
xnor U12680 (N_12680,N_11360,N_11585);
and U12681 (N_12681,N_11578,N_11547);
and U12682 (N_12682,N_11290,N_11697);
or U12683 (N_12683,N_11313,N_11589);
xnor U12684 (N_12684,N_11323,N_11756);
and U12685 (N_12685,N_11449,N_11321);
and U12686 (N_12686,N_11849,N_11549);
and U12687 (N_12687,N_11429,N_11502);
nor U12688 (N_12688,N_11971,N_11940);
or U12689 (N_12689,N_11682,N_11838);
nor U12690 (N_12690,N_11529,N_11854);
nor U12691 (N_12691,N_11440,N_11559);
nand U12692 (N_12692,N_11357,N_11528);
xnor U12693 (N_12693,N_11914,N_11571);
xnor U12694 (N_12694,N_11681,N_11626);
xor U12695 (N_12695,N_11965,N_11858);
or U12696 (N_12696,N_11883,N_11435);
nor U12697 (N_12697,N_11534,N_11469);
xor U12698 (N_12698,N_11747,N_11938);
xnor U12699 (N_12699,N_11991,N_11892);
nor U12700 (N_12700,N_11469,N_11674);
nor U12701 (N_12701,N_11535,N_11562);
xor U12702 (N_12702,N_11698,N_11684);
xor U12703 (N_12703,N_11399,N_11635);
nand U12704 (N_12704,N_11943,N_11354);
nand U12705 (N_12705,N_11887,N_11335);
nor U12706 (N_12706,N_11849,N_11430);
and U12707 (N_12707,N_11683,N_11698);
xnor U12708 (N_12708,N_11818,N_11317);
nand U12709 (N_12709,N_11429,N_11559);
nor U12710 (N_12710,N_11917,N_11788);
nor U12711 (N_12711,N_11277,N_11333);
nand U12712 (N_12712,N_11570,N_11777);
and U12713 (N_12713,N_11558,N_11537);
and U12714 (N_12714,N_11918,N_11854);
nor U12715 (N_12715,N_11649,N_11256);
nand U12716 (N_12716,N_11670,N_11507);
and U12717 (N_12717,N_11562,N_11681);
nand U12718 (N_12718,N_11583,N_11505);
and U12719 (N_12719,N_11997,N_11885);
nand U12720 (N_12720,N_11998,N_11315);
nor U12721 (N_12721,N_11706,N_11500);
or U12722 (N_12722,N_11583,N_11419);
xor U12723 (N_12723,N_11645,N_11417);
nor U12724 (N_12724,N_11316,N_11465);
and U12725 (N_12725,N_11545,N_11757);
xnor U12726 (N_12726,N_11533,N_11288);
nor U12727 (N_12727,N_11358,N_11255);
and U12728 (N_12728,N_11490,N_11393);
xnor U12729 (N_12729,N_11824,N_11429);
or U12730 (N_12730,N_11630,N_11832);
nor U12731 (N_12731,N_11708,N_11780);
nor U12732 (N_12732,N_11589,N_11811);
or U12733 (N_12733,N_11523,N_11917);
or U12734 (N_12734,N_11451,N_11996);
nand U12735 (N_12735,N_11484,N_11331);
or U12736 (N_12736,N_11321,N_11520);
and U12737 (N_12737,N_11787,N_11744);
xnor U12738 (N_12738,N_11326,N_11509);
nand U12739 (N_12739,N_11582,N_11250);
nand U12740 (N_12740,N_11726,N_11884);
and U12741 (N_12741,N_11643,N_11645);
nand U12742 (N_12742,N_11642,N_11836);
xor U12743 (N_12743,N_11901,N_11925);
and U12744 (N_12744,N_11596,N_11779);
xor U12745 (N_12745,N_11312,N_11543);
or U12746 (N_12746,N_11362,N_11287);
and U12747 (N_12747,N_11922,N_11917);
nor U12748 (N_12748,N_11658,N_11353);
xor U12749 (N_12749,N_11692,N_11911);
nand U12750 (N_12750,N_12387,N_12615);
nand U12751 (N_12751,N_12281,N_12317);
or U12752 (N_12752,N_12645,N_12115);
nor U12753 (N_12753,N_12063,N_12324);
xor U12754 (N_12754,N_12584,N_12284);
and U12755 (N_12755,N_12233,N_12206);
nor U12756 (N_12756,N_12350,N_12680);
nor U12757 (N_12757,N_12430,N_12376);
nor U12758 (N_12758,N_12023,N_12503);
nand U12759 (N_12759,N_12030,N_12444);
or U12760 (N_12760,N_12704,N_12014);
nand U12761 (N_12761,N_12577,N_12170);
nor U12762 (N_12762,N_12223,N_12360);
and U12763 (N_12763,N_12139,N_12517);
or U12764 (N_12764,N_12679,N_12307);
nand U12765 (N_12765,N_12555,N_12187);
or U12766 (N_12766,N_12055,N_12156);
nor U12767 (N_12767,N_12639,N_12747);
or U12768 (N_12768,N_12609,N_12658);
nand U12769 (N_12769,N_12237,N_12621);
nand U12770 (N_12770,N_12379,N_12670);
nor U12771 (N_12771,N_12560,N_12611);
or U12772 (N_12772,N_12031,N_12336);
xnor U12773 (N_12773,N_12147,N_12678);
and U12774 (N_12774,N_12054,N_12294);
xnor U12775 (N_12775,N_12586,N_12086);
xnor U12776 (N_12776,N_12238,N_12343);
or U12777 (N_12777,N_12509,N_12576);
nand U12778 (N_12778,N_12537,N_12362);
and U12779 (N_12779,N_12202,N_12308);
nand U12780 (N_12780,N_12268,N_12518);
xnor U12781 (N_12781,N_12501,N_12441);
or U12782 (N_12782,N_12231,N_12447);
nand U12783 (N_12783,N_12296,N_12392);
xor U12784 (N_12784,N_12065,N_12458);
nand U12785 (N_12785,N_12389,N_12559);
or U12786 (N_12786,N_12456,N_12262);
or U12787 (N_12787,N_12278,N_12465);
nor U12788 (N_12788,N_12071,N_12532);
xor U12789 (N_12789,N_12097,N_12190);
and U12790 (N_12790,N_12005,N_12269);
nand U12791 (N_12791,N_12736,N_12128);
or U12792 (N_12792,N_12689,N_12393);
xnor U12793 (N_12793,N_12104,N_12654);
or U12794 (N_12794,N_12561,N_12650);
nand U12795 (N_12795,N_12046,N_12460);
nand U12796 (N_12796,N_12204,N_12085);
or U12797 (N_12797,N_12466,N_12478);
or U12798 (N_12798,N_12333,N_12397);
or U12799 (N_12799,N_12527,N_12676);
nor U12800 (N_12800,N_12511,N_12148);
nand U12801 (N_12801,N_12042,N_12207);
nand U12802 (N_12802,N_12215,N_12058);
xnor U12803 (N_12803,N_12677,N_12717);
nor U12804 (N_12804,N_12123,N_12475);
nand U12805 (N_12805,N_12052,N_12361);
and U12806 (N_12806,N_12109,N_12339);
nor U12807 (N_12807,N_12468,N_12287);
or U12808 (N_12808,N_12493,N_12320);
and U12809 (N_12809,N_12276,N_12174);
nand U12810 (N_12810,N_12270,N_12606);
and U12811 (N_12811,N_12175,N_12089);
nor U12812 (N_12812,N_12210,N_12574);
or U12813 (N_12813,N_12247,N_12558);
nand U12814 (N_12814,N_12303,N_12041);
nor U12815 (N_12815,N_12154,N_12136);
nand U12816 (N_12816,N_12267,N_12453);
xor U12817 (N_12817,N_12483,N_12044);
nor U12818 (N_12818,N_12079,N_12024);
xnor U12819 (N_12819,N_12243,N_12193);
nand U12820 (N_12820,N_12127,N_12626);
nor U12821 (N_12821,N_12033,N_12640);
nand U12822 (N_12822,N_12731,N_12330);
nand U12823 (N_12823,N_12486,N_12675);
nand U12824 (N_12824,N_12533,N_12335);
nand U12825 (N_12825,N_12029,N_12107);
nand U12826 (N_12826,N_12334,N_12363);
xor U12827 (N_12827,N_12668,N_12045);
nand U12828 (N_12828,N_12399,N_12498);
or U12829 (N_12829,N_12290,N_12516);
or U12830 (N_12830,N_12013,N_12575);
nand U12831 (N_12831,N_12003,N_12607);
and U12832 (N_12832,N_12665,N_12250);
nor U12833 (N_12833,N_12552,N_12329);
or U12834 (N_12834,N_12698,N_12649);
or U12835 (N_12835,N_12573,N_12443);
and U12836 (N_12836,N_12007,N_12341);
or U12837 (N_12837,N_12508,N_12612);
nor U12838 (N_12838,N_12216,N_12484);
nand U12839 (N_12839,N_12548,N_12534);
or U12840 (N_12840,N_12218,N_12496);
xnor U12841 (N_12841,N_12017,N_12631);
nor U12842 (N_12842,N_12690,N_12239);
or U12843 (N_12843,N_12053,N_12227);
nand U12844 (N_12844,N_12211,N_12347);
or U12845 (N_12845,N_12624,N_12212);
or U12846 (N_12846,N_12248,N_12179);
nand U12847 (N_12847,N_12246,N_12356);
or U12848 (N_12848,N_12536,N_12372);
and U12849 (N_12849,N_12050,N_12126);
nor U12850 (N_12850,N_12157,N_12634);
and U12851 (N_12851,N_12070,N_12332);
xor U12852 (N_12852,N_12219,N_12488);
nor U12853 (N_12853,N_12378,N_12129);
xor U12854 (N_12854,N_12403,N_12208);
xor U12855 (N_12855,N_12656,N_12283);
and U12856 (N_12856,N_12472,N_12748);
xor U12857 (N_12857,N_12348,N_12681);
nor U12858 (N_12858,N_12662,N_12192);
nor U12859 (N_12859,N_12401,N_12171);
and U12860 (N_12860,N_12588,N_12744);
nor U12861 (N_12861,N_12742,N_12714);
xor U12862 (N_12862,N_12735,N_12661);
nand U12863 (N_12863,N_12370,N_12598);
and U12864 (N_12864,N_12669,N_12608);
xor U12865 (N_12865,N_12630,N_12386);
or U12866 (N_12866,N_12209,N_12112);
or U12867 (N_12867,N_12375,N_12181);
xor U12868 (N_12868,N_12095,N_12168);
xor U12869 (N_12869,N_12032,N_12718);
nor U12870 (N_12870,N_12295,N_12382);
nor U12871 (N_12871,N_12314,N_12197);
nand U12872 (N_12872,N_12277,N_12140);
and U12873 (N_12873,N_12073,N_12191);
or U12874 (N_12874,N_12686,N_12436);
nand U12875 (N_12875,N_12566,N_12494);
xor U12876 (N_12876,N_12617,N_12602);
and U12877 (N_12877,N_12522,N_12141);
or U12878 (N_12878,N_12728,N_12727);
nand U12879 (N_12879,N_12342,N_12489);
nor U12880 (N_12880,N_12265,N_12492);
nand U12881 (N_12881,N_12414,N_12049);
xnor U12882 (N_12882,N_12084,N_12235);
or U12883 (N_12883,N_12367,N_12463);
or U12884 (N_12884,N_12069,N_12582);
nand U12885 (N_12885,N_12258,N_12217);
and U12886 (N_12886,N_12051,N_12523);
and U12887 (N_12887,N_12520,N_12499);
nand U12888 (N_12888,N_12257,N_12571);
nand U12889 (N_12889,N_12528,N_12476);
xor U12890 (N_12890,N_12143,N_12180);
nand U12891 (N_12891,N_12599,N_12707);
nor U12892 (N_12892,N_12315,N_12705);
xor U12893 (N_12893,N_12732,N_12596);
nor U12894 (N_12894,N_12687,N_12729);
nand U12895 (N_12895,N_12064,N_12122);
xnor U12896 (N_12896,N_12477,N_12564);
or U12897 (N_12897,N_12539,N_12591);
nor U12898 (N_12898,N_12309,N_12697);
and U12899 (N_12899,N_12556,N_12442);
and U12900 (N_12900,N_12618,N_12568);
nor U12901 (N_12901,N_12098,N_12725);
nand U12902 (N_12902,N_12279,N_12060);
nand U12903 (N_12903,N_12435,N_12244);
nor U12904 (N_12904,N_12490,N_12225);
nand U12905 (N_12905,N_12485,N_12726);
nor U12906 (N_12906,N_12708,N_12629);
or U12907 (N_12907,N_12310,N_12312);
xor U12908 (N_12908,N_12423,N_12462);
and U12909 (N_12909,N_12711,N_12415);
nand U12910 (N_12910,N_12316,N_12578);
nand U12911 (N_12911,N_12119,N_12043);
xnor U12912 (N_12912,N_12094,N_12337);
and U12913 (N_12913,N_12567,N_12201);
nand U12914 (N_12914,N_12185,N_12530);
nand U12915 (N_12915,N_12396,N_12701);
xor U12916 (N_12916,N_12224,N_12454);
xor U12917 (N_12917,N_12006,N_12450);
xor U12918 (N_12918,N_12251,N_12565);
or U12919 (N_12919,N_12652,N_12724);
and U12920 (N_12920,N_12538,N_12021);
xnor U12921 (N_12921,N_12359,N_12167);
or U12922 (N_12922,N_12255,N_12205);
nand U12923 (N_12923,N_12001,N_12505);
or U12924 (N_12924,N_12660,N_12015);
xnor U12925 (N_12925,N_12616,N_12145);
or U12926 (N_12926,N_12637,N_12010);
nand U12927 (N_12927,N_12405,N_12721);
or U12928 (N_12928,N_12083,N_12614);
nand U12929 (N_12929,N_12331,N_12383);
and U12930 (N_12930,N_12152,N_12081);
nand U12931 (N_12931,N_12682,N_12402);
xnor U12932 (N_12932,N_12025,N_12076);
xnor U12933 (N_12933,N_12749,N_12713);
nand U12934 (N_12934,N_12432,N_12182);
nand U12935 (N_12935,N_12504,N_12229);
or U12936 (N_12936,N_12457,N_12090);
or U12937 (N_12937,N_12417,N_12271);
and U12938 (N_12938,N_12222,N_12221);
nand U12939 (N_12939,N_12035,N_12108);
nor U12940 (N_12940,N_12480,N_12072);
nand U12941 (N_12941,N_12091,N_12080);
nand U12942 (N_12942,N_12155,N_12743);
nand U12943 (N_12943,N_12018,N_12394);
nor U12944 (N_12944,N_12117,N_12026);
xnor U12945 (N_12945,N_12651,N_12666);
xor U12946 (N_12946,N_12138,N_12695);
and U12947 (N_12947,N_12028,N_12646);
and U12948 (N_12948,N_12293,N_12663);
or U12949 (N_12949,N_12694,N_12407);
or U12950 (N_12950,N_12427,N_12165);
or U12951 (N_12951,N_12068,N_12643);
xor U12952 (N_12952,N_12381,N_12635);
nor U12953 (N_12953,N_12413,N_12000);
nand U12954 (N_12954,N_12358,N_12338);
and U12955 (N_12955,N_12719,N_12059);
xnor U12956 (N_12956,N_12524,N_12481);
and U12957 (N_12957,N_12700,N_12589);
or U12958 (N_12958,N_12535,N_12422);
xnor U12959 (N_12959,N_12286,N_12737);
or U12960 (N_12960,N_12240,N_12592);
or U12961 (N_12961,N_12446,N_12706);
or U12962 (N_12962,N_12364,N_12692);
and U12963 (N_12963,N_12048,N_12377);
or U12964 (N_12964,N_12664,N_12703);
xnor U12965 (N_12965,N_12425,N_12604);
nor U12966 (N_12966,N_12543,N_12506);
nor U12967 (N_12967,N_12424,N_12088);
xnor U12968 (N_12968,N_12723,N_12467);
and U12969 (N_12969,N_12325,N_12684);
nor U12970 (N_12970,N_12730,N_12470);
nand U12971 (N_12971,N_12622,N_12572);
nand U12972 (N_12972,N_12605,N_12385);
nor U12973 (N_12973,N_12172,N_12092);
and U12974 (N_12974,N_12445,N_12259);
nand U12975 (N_12975,N_12437,N_12236);
nand U12976 (N_12976,N_12502,N_12159);
nor U12977 (N_12977,N_12228,N_12162);
xor U12978 (N_12978,N_12121,N_12234);
nor U12979 (N_12979,N_12304,N_12298);
and U12980 (N_12980,N_12184,N_12292);
nor U12981 (N_12981,N_12196,N_12547);
xnor U12982 (N_12982,N_12449,N_12693);
or U12983 (N_12983,N_12487,N_12100);
and U12984 (N_12984,N_12340,N_12620);
and U12985 (N_12985,N_12551,N_12553);
nor U12986 (N_12986,N_12130,N_12512);
and U12987 (N_12987,N_12638,N_12521);
and U12988 (N_12988,N_12513,N_12497);
or U12989 (N_12989,N_12408,N_12419);
nand U12990 (N_12990,N_12254,N_12570);
nor U12991 (N_12991,N_12173,N_12653);
or U12992 (N_12992,N_12299,N_12261);
or U12993 (N_12993,N_12531,N_12715);
nor U12994 (N_12994,N_12554,N_12297);
nor U12995 (N_12995,N_12289,N_12313);
nand U12996 (N_12996,N_12373,N_12074);
xor U12997 (N_12997,N_12352,N_12636);
and U12998 (N_12998,N_12149,N_12132);
nor U12999 (N_12999,N_12411,N_12507);
xor U13000 (N_13000,N_12011,N_12696);
xor U13001 (N_13001,N_12428,N_12491);
or U13002 (N_13002,N_12510,N_12452);
nand U13003 (N_13003,N_12199,N_12047);
or U13004 (N_13004,N_12544,N_12186);
nand U13005 (N_13005,N_12256,N_12305);
and U13006 (N_13006,N_12116,N_12061);
or U13007 (N_13007,N_12388,N_12264);
xnor U13008 (N_13008,N_12036,N_12124);
xor U13009 (N_13009,N_12365,N_12328);
or U13010 (N_13010,N_12291,N_12557);
nand U13011 (N_13011,N_12353,N_12710);
nand U13012 (N_13012,N_12434,N_12214);
nand U13013 (N_13013,N_12322,N_12702);
and U13014 (N_13014,N_12280,N_12406);
nand U13015 (N_13015,N_12648,N_12194);
nand U13016 (N_13016,N_12672,N_12323);
nor U13017 (N_13017,N_12716,N_12288);
or U13018 (N_13018,N_12078,N_12067);
xor U13019 (N_13019,N_12739,N_12549);
xor U13020 (N_13020,N_12722,N_12357);
nand U13021 (N_13021,N_12242,N_12657);
nor U13022 (N_13022,N_12161,N_12627);
or U13023 (N_13023,N_12495,N_12595);
nor U13024 (N_13024,N_12345,N_12075);
xor U13025 (N_13025,N_12683,N_12087);
or U13026 (N_13026,N_12623,N_12285);
xor U13027 (N_13027,N_12245,N_12355);
xnor U13028 (N_13028,N_12597,N_12712);
nor U13029 (N_13029,N_12164,N_12158);
nand U13030 (N_13030,N_12540,N_12579);
and U13031 (N_13031,N_12374,N_12593);
nand U13032 (N_13032,N_12034,N_12641);
or U13033 (N_13033,N_12009,N_12351);
nor U13034 (N_13034,N_12421,N_12318);
nand U13035 (N_13035,N_12213,N_12603);
or U13036 (N_13036,N_12390,N_12004);
xnor U13037 (N_13037,N_12688,N_12195);
or U13038 (N_13038,N_12169,N_12273);
xnor U13039 (N_13039,N_12368,N_12380);
nor U13040 (N_13040,N_12252,N_12327);
or U13041 (N_13041,N_12057,N_12022);
and U13042 (N_13042,N_12249,N_12633);
nor U13043 (N_13043,N_12581,N_12093);
nand U13044 (N_13044,N_12398,N_12569);
nor U13045 (N_13045,N_12198,N_12601);
xor U13046 (N_13046,N_12200,N_12272);
nand U13047 (N_13047,N_12241,N_12461);
nor U13048 (N_13048,N_12514,N_12118);
or U13049 (N_13049,N_12166,N_12134);
or U13050 (N_13050,N_12153,N_12188);
or U13051 (N_13051,N_12410,N_12594);
and U13052 (N_13052,N_12300,N_12220);
xor U13053 (N_13053,N_12404,N_12482);
xor U13054 (N_13054,N_12311,N_12178);
xnor U13055 (N_13055,N_12137,N_12203);
and U13056 (N_13056,N_12420,N_12619);
nor U13057 (N_13057,N_12082,N_12691);
and U13058 (N_13058,N_12176,N_12562);
xnor U13059 (N_13059,N_12580,N_12448);
or U13060 (N_13060,N_12189,N_12409);
and U13061 (N_13061,N_12451,N_12102);
nor U13062 (N_13062,N_12349,N_12738);
nor U13063 (N_13063,N_12099,N_12183);
xor U13064 (N_13064,N_12302,N_12671);
nor U13065 (N_13065,N_12418,N_12667);
nand U13066 (N_13066,N_12226,N_12741);
nor U13067 (N_13067,N_12439,N_12301);
and U13068 (N_13068,N_12734,N_12354);
or U13069 (N_13069,N_12369,N_12120);
nor U13070 (N_13070,N_12583,N_12125);
and U13071 (N_13071,N_12038,N_12039);
or U13072 (N_13072,N_12142,N_12344);
xor U13073 (N_13073,N_12647,N_12037);
nand U13074 (N_13074,N_12391,N_12019);
nand U13075 (N_13075,N_12529,N_12585);
nand U13076 (N_13076,N_12459,N_12135);
nor U13077 (N_13077,N_12266,N_12160);
or U13078 (N_13078,N_12455,N_12642);
nand U13079 (N_13079,N_12012,N_12674);
or U13080 (N_13080,N_12366,N_12306);
and U13081 (N_13081,N_12500,N_12101);
or U13082 (N_13082,N_12144,N_12590);
nand U13083 (N_13083,N_12321,N_12110);
nor U13084 (N_13084,N_12745,N_12066);
or U13085 (N_13085,N_12733,N_12008);
and U13086 (N_13086,N_12610,N_12525);
nand U13087 (N_13087,N_12709,N_12177);
nand U13088 (N_13088,N_12479,N_12746);
or U13089 (N_13089,N_12096,N_12163);
nand U13090 (N_13090,N_12546,N_12111);
xnor U13091 (N_13091,N_12105,N_12395);
nor U13092 (N_13092,N_12426,N_12282);
nor U13093 (N_13093,N_12440,N_12253);
and U13094 (N_13094,N_12438,N_12274);
nand U13095 (N_13095,N_12062,N_12655);
and U13096 (N_13096,N_12659,N_12230);
nor U13097 (N_13097,N_12346,N_12699);
and U13098 (N_13098,N_12474,N_12469);
and U13099 (N_13099,N_12114,N_12473);
or U13100 (N_13100,N_12685,N_12027);
nand U13101 (N_13101,N_12545,N_12002);
or U13102 (N_13102,N_12150,N_12587);
and U13103 (N_13103,N_12020,N_12550);
or U13104 (N_13104,N_12384,N_12644);
nand U13105 (N_13105,N_12326,N_12232);
xnor U13106 (N_13106,N_12400,N_12146);
nand U13107 (N_13107,N_12433,N_12515);
and U13108 (N_13108,N_12613,N_12519);
and U13109 (N_13109,N_12464,N_12632);
or U13110 (N_13110,N_12319,N_12416);
xor U13111 (N_13111,N_12431,N_12151);
nand U13112 (N_13112,N_12526,N_12740);
or U13113 (N_13113,N_12541,N_12263);
and U13114 (N_13114,N_12628,N_12542);
nor U13115 (N_13115,N_12563,N_12371);
and U13116 (N_13116,N_12600,N_12471);
nand U13117 (N_13117,N_12133,N_12625);
xor U13118 (N_13118,N_12103,N_12673);
or U13119 (N_13119,N_12056,N_12260);
nand U13120 (N_13120,N_12077,N_12040);
or U13121 (N_13121,N_12275,N_12113);
and U13122 (N_13122,N_12720,N_12412);
or U13123 (N_13123,N_12106,N_12131);
or U13124 (N_13124,N_12016,N_12429);
xor U13125 (N_13125,N_12522,N_12363);
or U13126 (N_13126,N_12282,N_12474);
or U13127 (N_13127,N_12682,N_12056);
nor U13128 (N_13128,N_12488,N_12363);
nor U13129 (N_13129,N_12275,N_12539);
nand U13130 (N_13130,N_12301,N_12583);
and U13131 (N_13131,N_12120,N_12003);
nand U13132 (N_13132,N_12715,N_12013);
nand U13133 (N_13133,N_12596,N_12135);
xnor U13134 (N_13134,N_12375,N_12525);
nand U13135 (N_13135,N_12116,N_12099);
or U13136 (N_13136,N_12015,N_12718);
nand U13137 (N_13137,N_12485,N_12270);
xor U13138 (N_13138,N_12042,N_12104);
nand U13139 (N_13139,N_12158,N_12191);
and U13140 (N_13140,N_12131,N_12246);
xor U13141 (N_13141,N_12525,N_12335);
or U13142 (N_13142,N_12534,N_12650);
or U13143 (N_13143,N_12046,N_12356);
xor U13144 (N_13144,N_12701,N_12660);
nor U13145 (N_13145,N_12612,N_12739);
or U13146 (N_13146,N_12309,N_12584);
nor U13147 (N_13147,N_12509,N_12079);
nand U13148 (N_13148,N_12070,N_12212);
or U13149 (N_13149,N_12397,N_12515);
or U13150 (N_13150,N_12526,N_12556);
nor U13151 (N_13151,N_12223,N_12371);
and U13152 (N_13152,N_12411,N_12340);
or U13153 (N_13153,N_12499,N_12514);
nor U13154 (N_13154,N_12252,N_12558);
or U13155 (N_13155,N_12117,N_12014);
and U13156 (N_13156,N_12296,N_12352);
xnor U13157 (N_13157,N_12360,N_12283);
nor U13158 (N_13158,N_12164,N_12430);
nor U13159 (N_13159,N_12608,N_12557);
nor U13160 (N_13160,N_12232,N_12637);
nand U13161 (N_13161,N_12634,N_12442);
nand U13162 (N_13162,N_12382,N_12622);
and U13163 (N_13163,N_12723,N_12633);
and U13164 (N_13164,N_12463,N_12145);
nor U13165 (N_13165,N_12617,N_12586);
or U13166 (N_13166,N_12337,N_12579);
nand U13167 (N_13167,N_12701,N_12277);
and U13168 (N_13168,N_12260,N_12161);
or U13169 (N_13169,N_12441,N_12367);
nor U13170 (N_13170,N_12469,N_12566);
and U13171 (N_13171,N_12581,N_12135);
and U13172 (N_13172,N_12654,N_12618);
and U13173 (N_13173,N_12398,N_12180);
and U13174 (N_13174,N_12289,N_12710);
nor U13175 (N_13175,N_12601,N_12716);
and U13176 (N_13176,N_12257,N_12058);
xor U13177 (N_13177,N_12168,N_12704);
nand U13178 (N_13178,N_12246,N_12084);
and U13179 (N_13179,N_12654,N_12240);
nand U13180 (N_13180,N_12242,N_12662);
and U13181 (N_13181,N_12606,N_12209);
nor U13182 (N_13182,N_12349,N_12584);
xor U13183 (N_13183,N_12382,N_12377);
xnor U13184 (N_13184,N_12108,N_12623);
xnor U13185 (N_13185,N_12524,N_12410);
xnor U13186 (N_13186,N_12158,N_12071);
nor U13187 (N_13187,N_12341,N_12077);
nand U13188 (N_13188,N_12190,N_12575);
or U13189 (N_13189,N_12319,N_12297);
xnor U13190 (N_13190,N_12574,N_12443);
nor U13191 (N_13191,N_12495,N_12557);
or U13192 (N_13192,N_12028,N_12077);
nand U13193 (N_13193,N_12086,N_12062);
or U13194 (N_13194,N_12231,N_12332);
nand U13195 (N_13195,N_12186,N_12053);
and U13196 (N_13196,N_12651,N_12056);
and U13197 (N_13197,N_12480,N_12519);
and U13198 (N_13198,N_12075,N_12645);
nand U13199 (N_13199,N_12293,N_12255);
nor U13200 (N_13200,N_12044,N_12516);
nand U13201 (N_13201,N_12553,N_12617);
and U13202 (N_13202,N_12429,N_12382);
nand U13203 (N_13203,N_12568,N_12284);
or U13204 (N_13204,N_12322,N_12051);
xor U13205 (N_13205,N_12388,N_12567);
nor U13206 (N_13206,N_12247,N_12298);
nand U13207 (N_13207,N_12116,N_12118);
and U13208 (N_13208,N_12261,N_12283);
xnor U13209 (N_13209,N_12642,N_12689);
nor U13210 (N_13210,N_12405,N_12737);
nor U13211 (N_13211,N_12295,N_12439);
nand U13212 (N_13212,N_12629,N_12565);
or U13213 (N_13213,N_12424,N_12274);
or U13214 (N_13214,N_12502,N_12557);
or U13215 (N_13215,N_12619,N_12299);
xor U13216 (N_13216,N_12403,N_12008);
or U13217 (N_13217,N_12378,N_12576);
xnor U13218 (N_13218,N_12655,N_12646);
or U13219 (N_13219,N_12748,N_12439);
nor U13220 (N_13220,N_12230,N_12452);
xnor U13221 (N_13221,N_12014,N_12017);
and U13222 (N_13222,N_12554,N_12325);
nand U13223 (N_13223,N_12116,N_12280);
nand U13224 (N_13224,N_12438,N_12426);
xnor U13225 (N_13225,N_12359,N_12361);
xor U13226 (N_13226,N_12082,N_12138);
nand U13227 (N_13227,N_12139,N_12466);
or U13228 (N_13228,N_12015,N_12498);
nor U13229 (N_13229,N_12637,N_12141);
xor U13230 (N_13230,N_12603,N_12410);
nand U13231 (N_13231,N_12115,N_12740);
or U13232 (N_13232,N_12677,N_12076);
xor U13233 (N_13233,N_12637,N_12105);
nor U13234 (N_13234,N_12114,N_12014);
nand U13235 (N_13235,N_12572,N_12195);
nor U13236 (N_13236,N_12533,N_12028);
xor U13237 (N_13237,N_12250,N_12000);
nor U13238 (N_13238,N_12098,N_12202);
nand U13239 (N_13239,N_12106,N_12053);
and U13240 (N_13240,N_12434,N_12285);
or U13241 (N_13241,N_12595,N_12093);
xor U13242 (N_13242,N_12196,N_12567);
or U13243 (N_13243,N_12552,N_12270);
xnor U13244 (N_13244,N_12165,N_12702);
xnor U13245 (N_13245,N_12547,N_12538);
and U13246 (N_13246,N_12058,N_12392);
nor U13247 (N_13247,N_12693,N_12537);
xor U13248 (N_13248,N_12748,N_12533);
or U13249 (N_13249,N_12690,N_12602);
xnor U13250 (N_13250,N_12104,N_12168);
or U13251 (N_13251,N_12369,N_12233);
nor U13252 (N_13252,N_12362,N_12495);
xor U13253 (N_13253,N_12202,N_12332);
nor U13254 (N_13254,N_12299,N_12467);
nor U13255 (N_13255,N_12610,N_12258);
nor U13256 (N_13256,N_12056,N_12727);
or U13257 (N_13257,N_12284,N_12687);
nand U13258 (N_13258,N_12731,N_12200);
nor U13259 (N_13259,N_12062,N_12526);
and U13260 (N_13260,N_12107,N_12596);
or U13261 (N_13261,N_12494,N_12472);
or U13262 (N_13262,N_12290,N_12544);
and U13263 (N_13263,N_12648,N_12647);
nand U13264 (N_13264,N_12553,N_12343);
xor U13265 (N_13265,N_12112,N_12022);
xor U13266 (N_13266,N_12423,N_12001);
or U13267 (N_13267,N_12632,N_12508);
nand U13268 (N_13268,N_12539,N_12571);
xnor U13269 (N_13269,N_12236,N_12146);
xor U13270 (N_13270,N_12049,N_12138);
nand U13271 (N_13271,N_12335,N_12324);
and U13272 (N_13272,N_12203,N_12240);
nand U13273 (N_13273,N_12500,N_12641);
xnor U13274 (N_13274,N_12341,N_12120);
nor U13275 (N_13275,N_12333,N_12480);
or U13276 (N_13276,N_12355,N_12242);
nor U13277 (N_13277,N_12493,N_12013);
nor U13278 (N_13278,N_12709,N_12328);
xnor U13279 (N_13279,N_12123,N_12340);
nand U13280 (N_13280,N_12087,N_12550);
or U13281 (N_13281,N_12271,N_12389);
and U13282 (N_13282,N_12560,N_12296);
or U13283 (N_13283,N_12046,N_12373);
and U13284 (N_13284,N_12263,N_12383);
nand U13285 (N_13285,N_12130,N_12556);
or U13286 (N_13286,N_12407,N_12597);
nor U13287 (N_13287,N_12345,N_12314);
nand U13288 (N_13288,N_12183,N_12292);
nor U13289 (N_13289,N_12289,N_12493);
nor U13290 (N_13290,N_12139,N_12048);
and U13291 (N_13291,N_12587,N_12231);
xnor U13292 (N_13292,N_12213,N_12098);
xor U13293 (N_13293,N_12457,N_12464);
xor U13294 (N_13294,N_12558,N_12423);
nor U13295 (N_13295,N_12515,N_12562);
xor U13296 (N_13296,N_12386,N_12273);
nand U13297 (N_13297,N_12438,N_12016);
or U13298 (N_13298,N_12208,N_12184);
and U13299 (N_13299,N_12243,N_12167);
xnor U13300 (N_13300,N_12223,N_12534);
nand U13301 (N_13301,N_12160,N_12454);
xor U13302 (N_13302,N_12081,N_12025);
nand U13303 (N_13303,N_12346,N_12313);
or U13304 (N_13304,N_12362,N_12582);
xor U13305 (N_13305,N_12336,N_12462);
nand U13306 (N_13306,N_12151,N_12516);
or U13307 (N_13307,N_12338,N_12501);
nor U13308 (N_13308,N_12170,N_12261);
or U13309 (N_13309,N_12232,N_12330);
nand U13310 (N_13310,N_12146,N_12054);
nand U13311 (N_13311,N_12495,N_12406);
nor U13312 (N_13312,N_12159,N_12668);
nor U13313 (N_13313,N_12445,N_12075);
and U13314 (N_13314,N_12290,N_12409);
nor U13315 (N_13315,N_12359,N_12203);
or U13316 (N_13316,N_12205,N_12111);
nand U13317 (N_13317,N_12633,N_12413);
nand U13318 (N_13318,N_12153,N_12513);
xnor U13319 (N_13319,N_12022,N_12028);
nand U13320 (N_13320,N_12494,N_12712);
or U13321 (N_13321,N_12614,N_12430);
and U13322 (N_13322,N_12626,N_12739);
and U13323 (N_13323,N_12706,N_12274);
nand U13324 (N_13324,N_12549,N_12238);
nand U13325 (N_13325,N_12059,N_12142);
nor U13326 (N_13326,N_12320,N_12381);
and U13327 (N_13327,N_12219,N_12429);
nor U13328 (N_13328,N_12316,N_12030);
and U13329 (N_13329,N_12515,N_12480);
xnor U13330 (N_13330,N_12256,N_12020);
xnor U13331 (N_13331,N_12114,N_12551);
xnor U13332 (N_13332,N_12276,N_12516);
nand U13333 (N_13333,N_12158,N_12324);
nor U13334 (N_13334,N_12635,N_12006);
and U13335 (N_13335,N_12716,N_12643);
nand U13336 (N_13336,N_12701,N_12037);
nand U13337 (N_13337,N_12565,N_12250);
xor U13338 (N_13338,N_12575,N_12057);
nand U13339 (N_13339,N_12366,N_12190);
and U13340 (N_13340,N_12502,N_12311);
or U13341 (N_13341,N_12588,N_12686);
nor U13342 (N_13342,N_12350,N_12001);
nor U13343 (N_13343,N_12296,N_12300);
or U13344 (N_13344,N_12488,N_12304);
nand U13345 (N_13345,N_12526,N_12275);
and U13346 (N_13346,N_12444,N_12395);
and U13347 (N_13347,N_12092,N_12575);
nand U13348 (N_13348,N_12506,N_12191);
nand U13349 (N_13349,N_12438,N_12193);
nand U13350 (N_13350,N_12283,N_12448);
nor U13351 (N_13351,N_12603,N_12602);
xor U13352 (N_13352,N_12194,N_12584);
or U13353 (N_13353,N_12651,N_12658);
nand U13354 (N_13354,N_12525,N_12271);
and U13355 (N_13355,N_12519,N_12195);
xnor U13356 (N_13356,N_12021,N_12462);
and U13357 (N_13357,N_12293,N_12625);
xnor U13358 (N_13358,N_12175,N_12395);
xnor U13359 (N_13359,N_12278,N_12712);
or U13360 (N_13360,N_12298,N_12212);
nand U13361 (N_13361,N_12191,N_12098);
nor U13362 (N_13362,N_12749,N_12628);
or U13363 (N_13363,N_12034,N_12107);
nand U13364 (N_13364,N_12386,N_12154);
or U13365 (N_13365,N_12046,N_12500);
nor U13366 (N_13366,N_12323,N_12260);
nand U13367 (N_13367,N_12520,N_12036);
or U13368 (N_13368,N_12317,N_12626);
or U13369 (N_13369,N_12438,N_12313);
nor U13370 (N_13370,N_12162,N_12205);
and U13371 (N_13371,N_12204,N_12594);
xor U13372 (N_13372,N_12385,N_12581);
nand U13373 (N_13373,N_12322,N_12565);
xnor U13374 (N_13374,N_12182,N_12394);
nor U13375 (N_13375,N_12211,N_12560);
and U13376 (N_13376,N_12394,N_12546);
nor U13377 (N_13377,N_12355,N_12722);
xnor U13378 (N_13378,N_12702,N_12041);
and U13379 (N_13379,N_12357,N_12481);
nor U13380 (N_13380,N_12124,N_12434);
xnor U13381 (N_13381,N_12388,N_12576);
and U13382 (N_13382,N_12628,N_12546);
and U13383 (N_13383,N_12157,N_12147);
nor U13384 (N_13384,N_12132,N_12458);
and U13385 (N_13385,N_12541,N_12027);
nor U13386 (N_13386,N_12152,N_12586);
nor U13387 (N_13387,N_12650,N_12603);
nor U13388 (N_13388,N_12494,N_12032);
or U13389 (N_13389,N_12298,N_12592);
xor U13390 (N_13390,N_12179,N_12568);
nor U13391 (N_13391,N_12285,N_12518);
and U13392 (N_13392,N_12538,N_12693);
nand U13393 (N_13393,N_12345,N_12003);
xnor U13394 (N_13394,N_12220,N_12140);
xnor U13395 (N_13395,N_12201,N_12012);
or U13396 (N_13396,N_12194,N_12087);
nand U13397 (N_13397,N_12006,N_12217);
or U13398 (N_13398,N_12223,N_12550);
or U13399 (N_13399,N_12178,N_12435);
nor U13400 (N_13400,N_12511,N_12675);
or U13401 (N_13401,N_12242,N_12473);
or U13402 (N_13402,N_12438,N_12029);
nand U13403 (N_13403,N_12633,N_12739);
xor U13404 (N_13404,N_12727,N_12402);
nand U13405 (N_13405,N_12342,N_12109);
or U13406 (N_13406,N_12010,N_12355);
xor U13407 (N_13407,N_12170,N_12014);
and U13408 (N_13408,N_12396,N_12522);
nand U13409 (N_13409,N_12318,N_12049);
or U13410 (N_13410,N_12384,N_12222);
or U13411 (N_13411,N_12407,N_12579);
nand U13412 (N_13412,N_12683,N_12579);
and U13413 (N_13413,N_12195,N_12652);
nor U13414 (N_13414,N_12114,N_12257);
nor U13415 (N_13415,N_12368,N_12628);
nand U13416 (N_13416,N_12103,N_12373);
nor U13417 (N_13417,N_12070,N_12083);
nor U13418 (N_13418,N_12246,N_12531);
nand U13419 (N_13419,N_12363,N_12441);
nand U13420 (N_13420,N_12441,N_12582);
nor U13421 (N_13421,N_12477,N_12541);
nand U13422 (N_13422,N_12214,N_12436);
nor U13423 (N_13423,N_12159,N_12602);
nand U13424 (N_13424,N_12712,N_12398);
nand U13425 (N_13425,N_12403,N_12264);
nand U13426 (N_13426,N_12707,N_12670);
nor U13427 (N_13427,N_12586,N_12244);
or U13428 (N_13428,N_12305,N_12573);
nand U13429 (N_13429,N_12737,N_12340);
and U13430 (N_13430,N_12546,N_12664);
or U13431 (N_13431,N_12113,N_12696);
xnor U13432 (N_13432,N_12033,N_12165);
and U13433 (N_13433,N_12222,N_12102);
or U13434 (N_13434,N_12075,N_12156);
xnor U13435 (N_13435,N_12250,N_12288);
nand U13436 (N_13436,N_12165,N_12699);
or U13437 (N_13437,N_12489,N_12699);
xor U13438 (N_13438,N_12117,N_12720);
or U13439 (N_13439,N_12607,N_12316);
and U13440 (N_13440,N_12316,N_12311);
nand U13441 (N_13441,N_12190,N_12383);
or U13442 (N_13442,N_12357,N_12673);
and U13443 (N_13443,N_12724,N_12522);
nand U13444 (N_13444,N_12302,N_12282);
or U13445 (N_13445,N_12391,N_12424);
and U13446 (N_13446,N_12202,N_12660);
and U13447 (N_13447,N_12227,N_12391);
xnor U13448 (N_13448,N_12166,N_12250);
and U13449 (N_13449,N_12344,N_12075);
nor U13450 (N_13450,N_12051,N_12656);
xnor U13451 (N_13451,N_12294,N_12358);
nand U13452 (N_13452,N_12223,N_12614);
xor U13453 (N_13453,N_12207,N_12287);
nor U13454 (N_13454,N_12065,N_12309);
nand U13455 (N_13455,N_12077,N_12317);
nor U13456 (N_13456,N_12642,N_12188);
nand U13457 (N_13457,N_12584,N_12464);
xnor U13458 (N_13458,N_12386,N_12476);
xnor U13459 (N_13459,N_12322,N_12045);
nand U13460 (N_13460,N_12171,N_12634);
xnor U13461 (N_13461,N_12735,N_12692);
or U13462 (N_13462,N_12372,N_12627);
xnor U13463 (N_13463,N_12719,N_12287);
or U13464 (N_13464,N_12144,N_12265);
and U13465 (N_13465,N_12249,N_12041);
and U13466 (N_13466,N_12315,N_12280);
nand U13467 (N_13467,N_12166,N_12227);
and U13468 (N_13468,N_12525,N_12503);
nor U13469 (N_13469,N_12213,N_12310);
nor U13470 (N_13470,N_12744,N_12626);
and U13471 (N_13471,N_12448,N_12270);
or U13472 (N_13472,N_12712,N_12720);
and U13473 (N_13473,N_12523,N_12408);
or U13474 (N_13474,N_12053,N_12269);
xnor U13475 (N_13475,N_12447,N_12078);
or U13476 (N_13476,N_12368,N_12233);
xnor U13477 (N_13477,N_12562,N_12294);
xor U13478 (N_13478,N_12171,N_12168);
and U13479 (N_13479,N_12686,N_12505);
nor U13480 (N_13480,N_12252,N_12660);
or U13481 (N_13481,N_12204,N_12030);
and U13482 (N_13482,N_12100,N_12179);
xnor U13483 (N_13483,N_12637,N_12393);
xnor U13484 (N_13484,N_12506,N_12442);
and U13485 (N_13485,N_12217,N_12276);
nand U13486 (N_13486,N_12432,N_12004);
nor U13487 (N_13487,N_12247,N_12245);
nor U13488 (N_13488,N_12242,N_12717);
or U13489 (N_13489,N_12319,N_12605);
or U13490 (N_13490,N_12471,N_12307);
nand U13491 (N_13491,N_12118,N_12705);
nand U13492 (N_13492,N_12019,N_12212);
or U13493 (N_13493,N_12223,N_12673);
xor U13494 (N_13494,N_12521,N_12642);
or U13495 (N_13495,N_12690,N_12331);
or U13496 (N_13496,N_12617,N_12729);
and U13497 (N_13497,N_12618,N_12076);
xnor U13498 (N_13498,N_12398,N_12024);
and U13499 (N_13499,N_12459,N_12058);
or U13500 (N_13500,N_13195,N_13426);
nand U13501 (N_13501,N_13105,N_13266);
nand U13502 (N_13502,N_13427,N_13245);
or U13503 (N_13503,N_13039,N_13060);
nor U13504 (N_13504,N_13433,N_12886);
nor U13505 (N_13505,N_13488,N_12903);
nand U13506 (N_13506,N_13406,N_13010);
xnor U13507 (N_13507,N_13100,N_13282);
or U13508 (N_13508,N_13000,N_13411);
and U13509 (N_13509,N_13090,N_13064);
nand U13510 (N_13510,N_13115,N_13131);
and U13511 (N_13511,N_12891,N_13168);
or U13512 (N_13512,N_13289,N_13377);
xor U13513 (N_13513,N_12775,N_13235);
xnor U13514 (N_13514,N_13112,N_12956);
nor U13515 (N_13515,N_13466,N_12796);
nand U13516 (N_13516,N_13357,N_12983);
and U13517 (N_13517,N_13445,N_13418);
nor U13518 (N_13518,N_13033,N_13422);
nor U13519 (N_13519,N_13181,N_13085);
xnor U13520 (N_13520,N_13253,N_13485);
xnor U13521 (N_13521,N_13149,N_12791);
or U13522 (N_13522,N_12830,N_13217);
nor U13523 (N_13523,N_12925,N_13356);
nand U13524 (N_13524,N_12911,N_13304);
nand U13525 (N_13525,N_13031,N_12974);
nor U13526 (N_13526,N_12959,N_12900);
nor U13527 (N_13527,N_13446,N_12902);
nor U13528 (N_13528,N_13080,N_13172);
nand U13529 (N_13529,N_13230,N_13143);
and U13530 (N_13530,N_12751,N_13331);
and U13531 (N_13531,N_12880,N_13099);
and U13532 (N_13532,N_13015,N_13117);
or U13533 (N_13533,N_13041,N_12767);
xor U13534 (N_13534,N_13258,N_13145);
and U13535 (N_13535,N_13447,N_12946);
nand U13536 (N_13536,N_13065,N_12894);
nand U13537 (N_13537,N_13081,N_13464);
and U13538 (N_13538,N_13495,N_12957);
or U13539 (N_13539,N_12968,N_13016);
nand U13540 (N_13540,N_12833,N_13469);
and U13541 (N_13541,N_13063,N_12826);
nor U13542 (N_13542,N_13297,N_13006);
xnor U13543 (N_13543,N_12843,N_13315);
nand U13544 (N_13544,N_13037,N_12770);
and U13545 (N_13545,N_13451,N_13483);
nand U13546 (N_13546,N_13075,N_13291);
or U13547 (N_13547,N_13110,N_13147);
and U13548 (N_13548,N_13102,N_12860);
xnor U13549 (N_13549,N_12982,N_12922);
xor U13550 (N_13550,N_13026,N_12892);
and U13551 (N_13551,N_12972,N_13299);
nor U13552 (N_13552,N_13129,N_13409);
and U13553 (N_13553,N_13474,N_13278);
nand U13554 (N_13554,N_12807,N_13313);
and U13555 (N_13555,N_13214,N_13259);
xor U13556 (N_13556,N_13206,N_12918);
and U13557 (N_13557,N_13255,N_13458);
nor U13558 (N_13558,N_12904,N_12781);
xor U13559 (N_13559,N_13240,N_12944);
and U13560 (N_13560,N_12761,N_13330);
nand U13561 (N_13561,N_12810,N_13173);
or U13562 (N_13562,N_13202,N_13155);
nor U13563 (N_13563,N_13076,N_12871);
nand U13564 (N_13564,N_12786,N_13398);
xor U13565 (N_13565,N_12965,N_12857);
and U13566 (N_13566,N_13449,N_12862);
nor U13567 (N_13567,N_12850,N_13264);
nand U13568 (N_13568,N_13349,N_13124);
or U13569 (N_13569,N_13092,N_13023);
and U13570 (N_13570,N_13316,N_13070);
nor U13571 (N_13571,N_13360,N_13327);
nand U13572 (N_13572,N_13222,N_13492);
nor U13573 (N_13573,N_13159,N_13152);
or U13574 (N_13574,N_13385,N_13400);
xor U13575 (N_13575,N_12960,N_12861);
nand U13576 (N_13576,N_13482,N_13002);
nor U13577 (N_13577,N_13397,N_13269);
and U13578 (N_13578,N_13061,N_12766);
and U13579 (N_13579,N_13233,N_13444);
or U13580 (N_13580,N_13440,N_13036);
or U13581 (N_13581,N_13054,N_13227);
xnor U13582 (N_13582,N_12869,N_13087);
nand U13583 (N_13583,N_13490,N_13365);
or U13584 (N_13584,N_12979,N_13103);
nor U13585 (N_13585,N_12962,N_13265);
xnor U13586 (N_13586,N_13186,N_12881);
or U13587 (N_13587,N_13093,N_13438);
nand U13588 (N_13588,N_13275,N_13216);
and U13589 (N_13589,N_12952,N_13012);
xnor U13590 (N_13590,N_13337,N_13040);
xor U13591 (N_13591,N_13188,N_13096);
and U13592 (N_13592,N_12805,N_12993);
nor U13593 (N_13593,N_13176,N_13234);
nor U13594 (N_13594,N_12831,N_13237);
or U13595 (N_13595,N_13208,N_12909);
or U13596 (N_13596,N_12859,N_13180);
xnor U13597 (N_13597,N_13004,N_12819);
nor U13598 (N_13598,N_13309,N_12936);
xor U13599 (N_13599,N_13138,N_13321);
or U13600 (N_13600,N_13396,N_13261);
xor U13601 (N_13601,N_13044,N_13118);
xnor U13602 (N_13602,N_13200,N_13342);
and U13603 (N_13603,N_12795,N_12759);
nand U13604 (N_13604,N_13194,N_12858);
nor U13605 (N_13605,N_13229,N_13336);
nor U13606 (N_13606,N_12836,N_13457);
nand U13607 (N_13607,N_13305,N_13161);
nor U13608 (N_13608,N_13276,N_12921);
and U13609 (N_13609,N_12799,N_12920);
or U13610 (N_13610,N_13371,N_12794);
nand U13611 (N_13611,N_12844,N_13473);
and U13612 (N_13612,N_12887,N_12899);
nor U13613 (N_13613,N_13462,N_13057);
nand U13614 (N_13614,N_13476,N_13211);
and U13615 (N_13615,N_13280,N_13153);
nor U13616 (N_13616,N_13496,N_13013);
and U13617 (N_13617,N_13011,N_12914);
and U13618 (N_13618,N_12879,N_13479);
nor U13619 (N_13619,N_13056,N_13192);
and U13620 (N_13620,N_13319,N_13437);
and U13621 (N_13621,N_13094,N_12809);
or U13622 (N_13622,N_13324,N_13442);
or U13623 (N_13623,N_13106,N_12874);
or U13624 (N_13624,N_12997,N_12910);
xor U13625 (N_13625,N_13018,N_12852);
xnor U13626 (N_13626,N_12923,N_13020);
or U13627 (N_13627,N_13286,N_13239);
nor U13628 (N_13628,N_13421,N_13114);
xnor U13629 (N_13629,N_12878,N_12950);
and U13630 (N_13630,N_13136,N_13133);
nand U13631 (N_13631,N_13210,N_12931);
and U13632 (N_13632,N_13032,N_13287);
xor U13633 (N_13633,N_13373,N_13379);
and U13634 (N_13634,N_13158,N_13499);
nor U13635 (N_13635,N_13363,N_13390);
xnor U13636 (N_13636,N_13244,N_13395);
or U13637 (N_13637,N_13215,N_13220);
or U13638 (N_13638,N_13046,N_13402);
nor U13639 (N_13639,N_12798,N_12981);
xor U13640 (N_13640,N_13189,N_13471);
xnor U13641 (N_13641,N_12930,N_12969);
and U13642 (N_13642,N_13213,N_12884);
or U13643 (N_13643,N_13197,N_13055);
xnor U13644 (N_13644,N_13104,N_12764);
and U13645 (N_13645,N_13480,N_12829);
and U13646 (N_13646,N_13248,N_13338);
and U13647 (N_13647,N_13370,N_13263);
and U13648 (N_13648,N_12973,N_12812);
nor U13649 (N_13649,N_12890,N_13311);
and U13650 (N_13650,N_13497,N_12938);
or U13651 (N_13651,N_13027,N_13095);
nor U13652 (N_13652,N_13272,N_13157);
or U13653 (N_13653,N_13074,N_12951);
or U13654 (N_13654,N_12929,N_12793);
nor U13655 (N_13655,N_12961,N_12937);
nand U13656 (N_13656,N_12995,N_13389);
or U13657 (N_13657,N_13268,N_12901);
nand U13658 (N_13658,N_13128,N_13163);
xnor U13659 (N_13659,N_13169,N_12953);
nand U13660 (N_13660,N_13450,N_13049);
and U13661 (N_13661,N_13439,N_12898);
xnor U13662 (N_13662,N_13212,N_13267);
nor U13663 (N_13663,N_13302,N_13467);
and U13664 (N_13664,N_13257,N_12855);
nor U13665 (N_13665,N_13205,N_13050);
or U13666 (N_13666,N_13294,N_12987);
nor U13667 (N_13667,N_12753,N_13201);
nor U13668 (N_13668,N_12964,N_13150);
xor U13669 (N_13669,N_13007,N_13303);
nor U13670 (N_13670,N_12877,N_13077);
nor U13671 (N_13671,N_13098,N_13366);
nor U13672 (N_13672,N_13034,N_13408);
nor U13673 (N_13673,N_13281,N_13290);
or U13674 (N_13674,N_12967,N_13463);
or U13675 (N_13675,N_12897,N_13394);
or U13676 (N_13676,N_13340,N_13160);
or U13677 (N_13677,N_13486,N_13254);
nor U13678 (N_13678,N_12822,N_12845);
nor U13679 (N_13679,N_12846,N_12814);
nand U13680 (N_13680,N_13154,N_13251);
nand U13681 (N_13681,N_13089,N_12977);
nor U13682 (N_13682,N_13226,N_12986);
nor U13683 (N_13683,N_13380,N_13196);
nor U13684 (N_13684,N_13417,N_12940);
nor U13685 (N_13685,N_13456,N_13284);
xnor U13686 (N_13686,N_13242,N_13224);
xnor U13687 (N_13687,N_12863,N_13475);
nand U13688 (N_13688,N_12966,N_13003);
xor U13689 (N_13689,N_13009,N_12989);
nor U13690 (N_13690,N_13454,N_13381);
nor U13691 (N_13691,N_13403,N_13329);
and U13692 (N_13692,N_13307,N_13119);
or U13693 (N_13693,N_13481,N_13300);
and U13694 (N_13694,N_13127,N_12917);
nand U13695 (N_13695,N_13353,N_13393);
nand U13696 (N_13696,N_13260,N_13101);
or U13697 (N_13697,N_13318,N_13148);
or U13698 (N_13698,N_13135,N_13292);
xor U13699 (N_13699,N_13301,N_13405);
xor U13700 (N_13700,N_13335,N_12851);
nor U13701 (N_13701,N_13218,N_13345);
nor U13702 (N_13702,N_12970,N_12971);
nand U13703 (N_13703,N_13174,N_12928);
xor U13704 (N_13704,N_13182,N_13484);
or U13705 (N_13705,N_12991,N_12943);
nand U13706 (N_13706,N_13035,N_12872);
nor U13707 (N_13707,N_13053,N_12856);
nor U13708 (N_13708,N_13191,N_13171);
xor U13709 (N_13709,N_12760,N_12808);
nor U13710 (N_13710,N_12954,N_13024);
or U13711 (N_13711,N_13107,N_12769);
xor U13712 (N_13712,N_12754,N_13066);
and U13713 (N_13713,N_13151,N_13341);
nor U13714 (N_13714,N_13051,N_12768);
or U13715 (N_13715,N_13392,N_12924);
and U13716 (N_13716,N_12750,N_12818);
and U13717 (N_13717,N_12849,N_12820);
xor U13718 (N_13718,N_13428,N_13452);
and U13719 (N_13719,N_13088,N_13415);
nand U13720 (N_13720,N_12867,N_12998);
and U13721 (N_13721,N_13320,N_13375);
or U13722 (N_13722,N_13332,N_12876);
nor U13723 (N_13723,N_12932,N_12756);
and U13724 (N_13724,N_13108,N_12915);
nand U13725 (N_13725,N_12763,N_12806);
nor U13726 (N_13726,N_13354,N_13178);
nor U13727 (N_13727,N_12824,N_12823);
nor U13728 (N_13728,N_13091,N_13014);
xnor U13729 (N_13729,N_12813,N_13071);
xnor U13730 (N_13730,N_12839,N_13052);
xnor U13731 (N_13731,N_13468,N_13472);
nor U13732 (N_13732,N_13019,N_13310);
xor U13733 (N_13733,N_13241,N_13126);
nand U13734 (N_13734,N_12840,N_13042);
xnor U13735 (N_13735,N_12975,N_13420);
nor U13736 (N_13736,N_13325,N_13435);
or U13737 (N_13737,N_13461,N_13339);
nand U13738 (N_13738,N_12771,N_13317);
xnor U13739 (N_13739,N_13223,N_13142);
or U13740 (N_13740,N_12948,N_13460);
or U13741 (N_13741,N_12792,N_13207);
and U13742 (N_13742,N_12803,N_13384);
or U13743 (N_13743,N_13141,N_12817);
xnor U13744 (N_13744,N_13121,N_13005);
xnor U13745 (N_13745,N_13491,N_12841);
and U13746 (N_13746,N_13184,N_13021);
xor U13747 (N_13747,N_13123,N_12958);
xnor U13748 (N_13748,N_13277,N_12868);
and U13749 (N_13749,N_12847,N_12828);
xor U13750 (N_13750,N_12802,N_12815);
or U13751 (N_13751,N_12801,N_13022);
xnor U13752 (N_13752,N_12895,N_13477);
and U13753 (N_13753,N_12865,N_13111);
nand U13754 (N_13754,N_13079,N_13203);
or U13755 (N_13755,N_13073,N_13025);
and U13756 (N_13756,N_13225,N_13132);
or U13757 (N_13757,N_13465,N_13298);
nor U13758 (N_13758,N_13185,N_13249);
and U13759 (N_13759,N_13498,N_13137);
nor U13760 (N_13760,N_13347,N_12908);
nand U13761 (N_13761,N_13165,N_13362);
xnor U13762 (N_13762,N_13164,N_13130);
or U13763 (N_13763,N_13274,N_12800);
nand U13764 (N_13764,N_13493,N_13270);
nor U13765 (N_13765,N_13334,N_13293);
and U13766 (N_13766,N_12864,N_12832);
xor U13767 (N_13767,N_12999,N_13062);
or U13768 (N_13768,N_12853,N_12757);
nand U13769 (N_13769,N_12939,N_12934);
and U13770 (N_13770,N_13116,N_12787);
nor U13771 (N_13771,N_12949,N_12835);
and U13772 (N_13772,N_12797,N_12883);
nand U13773 (N_13773,N_13391,N_12752);
nand U13774 (N_13774,N_12912,N_13047);
or U13775 (N_13775,N_12882,N_13441);
nand U13776 (N_13776,N_13029,N_13350);
xor U13777 (N_13777,N_12947,N_12777);
or U13778 (N_13778,N_13431,N_13401);
and U13779 (N_13779,N_12889,N_13068);
and U13780 (N_13780,N_12784,N_12785);
nor U13781 (N_13781,N_13043,N_13346);
xnor U13782 (N_13782,N_13288,N_12926);
nand U13783 (N_13783,N_13410,N_12789);
xnor U13784 (N_13784,N_13361,N_12827);
nor U13785 (N_13785,N_12854,N_13008);
nor U13786 (N_13786,N_13238,N_13448);
or U13787 (N_13787,N_13256,N_13372);
nand U13788 (N_13788,N_12919,N_13030);
nor U13789 (N_13789,N_12780,N_13199);
or U13790 (N_13790,N_13167,N_12913);
nand U13791 (N_13791,N_13364,N_13413);
nand U13792 (N_13792,N_13459,N_13387);
nor U13793 (N_13793,N_13312,N_13017);
nor U13794 (N_13794,N_13146,N_13236);
nand U13795 (N_13795,N_13399,N_13376);
xnor U13796 (N_13796,N_13209,N_13084);
or U13797 (N_13797,N_13028,N_13414);
xor U13798 (N_13798,N_12825,N_13175);
and U13799 (N_13799,N_13429,N_12990);
nand U13800 (N_13800,N_12955,N_13314);
nand U13801 (N_13801,N_12821,N_13228);
xor U13802 (N_13802,N_13295,N_13478);
nor U13803 (N_13803,N_12945,N_13424);
nand U13804 (N_13804,N_12838,N_13344);
nor U13805 (N_13805,N_13404,N_13083);
and U13806 (N_13806,N_12942,N_12875);
or U13807 (N_13807,N_13232,N_13359);
and U13808 (N_13808,N_13306,N_13134);
xor U13809 (N_13809,N_13069,N_13140);
nand U13810 (N_13810,N_12996,N_13072);
or U13811 (N_13811,N_12779,N_13470);
and U13812 (N_13812,N_13348,N_13416);
xor U13813 (N_13813,N_13378,N_13097);
or U13814 (N_13814,N_12933,N_12788);
nand U13815 (N_13815,N_13204,N_12873);
nor U13816 (N_13816,N_12762,N_13243);
nor U13817 (N_13817,N_12782,N_13283);
xor U13818 (N_13818,N_13343,N_13374);
or U13819 (N_13819,N_12790,N_13045);
xor U13820 (N_13820,N_12834,N_12842);
and U13821 (N_13821,N_13082,N_13308);
nor U13822 (N_13822,N_13388,N_12907);
nor U13823 (N_13823,N_13407,N_13271);
nand U13824 (N_13824,N_12896,N_13434);
nand U13825 (N_13825,N_13183,N_13455);
and U13826 (N_13826,N_12837,N_13179);
and U13827 (N_13827,N_13162,N_13323);
nor U13828 (N_13828,N_13193,N_13369);
and U13829 (N_13829,N_12870,N_13419);
and U13830 (N_13830,N_13273,N_12935);
nand U13831 (N_13831,N_12783,N_13086);
nor U13832 (N_13832,N_13368,N_13067);
nand U13833 (N_13833,N_13423,N_13487);
and U13834 (N_13834,N_12776,N_13494);
and U13835 (N_13835,N_12976,N_13383);
and U13836 (N_13836,N_13001,N_13190);
or U13837 (N_13837,N_13177,N_13412);
or U13838 (N_13838,N_12992,N_13078);
and U13839 (N_13839,N_12984,N_12893);
or U13840 (N_13840,N_12988,N_13386);
xor U13841 (N_13841,N_12773,N_13430);
or U13842 (N_13842,N_13144,N_13326);
nand U13843 (N_13843,N_13246,N_13425);
nand U13844 (N_13844,N_12758,N_13296);
xnor U13845 (N_13845,N_12941,N_13120);
and U13846 (N_13846,N_13453,N_13221);
nor U13847 (N_13847,N_12811,N_12848);
nor U13848 (N_13848,N_12816,N_12978);
xor U13849 (N_13849,N_13322,N_13285);
and U13850 (N_13850,N_13355,N_13109);
xnor U13851 (N_13851,N_13489,N_13328);
nand U13852 (N_13852,N_13352,N_12804);
nand U13853 (N_13853,N_12927,N_13048);
xnor U13854 (N_13854,N_13432,N_13122);
nand U13855 (N_13855,N_12980,N_13113);
and U13856 (N_13856,N_13382,N_12755);
and U13857 (N_13857,N_13252,N_12778);
xor U13858 (N_13858,N_13219,N_13333);
xnor U13859 (N_13859,N_13358,N_12774);
or U13860 (N_13860,N_13170,N_13058);
nor U13861 (N_13861,N_12765,N_12888);
or U13862 (N_13862,N_13038,N_13125);
or U13863 (N_13863,N_12905,N_13187);
nor U13864 (N_13864,N_12906,N_13436);
nor U13865 (N_13865,N_13367,N_13250);
and U13866 (N_13866,N_13279,N_12994);
nand U13867 (N_13867,N_12885,N_13139);
xnor U13868 (N_13868,N_13262,N_13351);
or U13869 (N_13869,N_13443,N_12963);
and U13870 (N_13870,N_12772,N_13247);
and U13871 (N_13871,N_12916,N_12866);
nor U13872 (N_13872,N_13166,N_13059);
xor U13873 (N_13873,N_13156,N_12985);
nand U13874 (N_13874,N_13198,N_13231);
xor U13875 (N_13875,N_12874,N_13145);
and U13876 (N_13876,N_13333,N_12884);
nand U13877 (N_13877,N_13098,N_13457);
and U13878 (N_13878,N_12878,N_13188);
and U13879 (N_13879,N_13348,N_12943);
nand U13880 (N_13880,N_12879,N_12894);
xnor U13881 (N_13881,N_12930,N_13440);
nand U13882 (N_13882,N_13369,N_13086);
xor U13883 (N_13883,N_13413,N_13470);
and U13884 (N_13884,N_12968,N_12903);
nor U13885 (N_13885,N_13496,N_13339);
nand U13886 (N_13886,N_12759,N_12752);
and U13887 (N_13887,N_12846,N_12949);
xnor U13888 (N_13888,N_12878,N_13115);
nor U13889 (N_13889,N_12761,N_13461);
xor U13890 (N_13890,N_13156,N_13152);
nor U13891 (N_13891,N_13210,N_13192);
and U13892 (N_13892,N_13189,N_13473);
or U13893 (N_13893,N_13389,N_13359);
or U13894 (N_13894,N_13071,N_12774);
or U13895 (N_13895,N_13138,N_13165);
nor U13896 (N_13896,N_13113,N_12926);
or U13897 (N_13897,N_12765,N_13157);
nor U13898 (N_13898,N_13403,N_13301);
xor U13899 (N_13899,N_12786,N_12902);
or U13900 (N_13900,N_13098,N_13085);
xor U13901 (N_13901,N_12949,N_13133);
nand U13902 (N_13902,N_12774,N_13122);
or U13903 (N_13903,N_12952,N_13270);
or U13904 (N_13904,N_13245,N_13019);
or U13905 (N_13905,N_13405,N_12761);
nor U13906 (N_13906,N_13421,N_13407);
xnor U13907 (N_13907,N_12790,N_13403);
and U13908 (N_13908,N_13334,N_12754);
and U13909 (N_13909,N_13177,N_13260);
nand U13910 (N_13910,N_13086,N_13265);
or U13911 (N_13911,N_13227,N_13218);
or U13912 (N_13912,N_12791,N_13333);
nand U13913 (N_13913,N_12876,N_13313);
nor U13914 (N_13914,N_13286,N_13192);
and U13915 (N_13915,N_12966,N_13122);
and U13916 (N_13916,N_13370,N_12763);
and U13917 (N_13917,N_12750,N_12843);
and U13918 (N_13918,N_13380,N_13184);
and U13919 (N_13919,N_13142,N_12984);
or U13920 (N_13920,N_13270,N_13079);
nor U13921 (N_13921,N_13024,N_12805);
xnor U13922 (N_13922,N_12980,N_13437);
and U13923 (N_13923,N_13213,N_13104);
nand U13924 (N_13924,N_13324,N_13477);
and U13925 (N_13925,N_12788,N_12782);
nor U13926 (N_13926,N_12764,N_13191);
xnor U13927 (N_13927,N_12908,N_12795);
xor U13928 (N_13928,N_13244,N_12932);
or U13929 (N_13929,N_12849,N_12857);
nor U13930 (N_13930,N_12965,N_13054);
xnor U13931 (N_13931,N_13113,N_13409);
nand U13932 (N_13932,N_13392,N_13420);
xor U13933 (N_13933,N_13147,N_13399);
nand U13934 (N_13934,N_13455,N_12814);
nor U13935 (N_13935,N_13312,N_13374);
nand U13936 (N_13936,N_12829,N_12985);
and U13937 (N_13937,N_13108,N_13090);
and U13938 (N_13938,N_12999,N_13392);
nor U13939 (N_13939,N_13149,N_13460);
and U13940 (N_13940,N_12964,N_13220);
or U13941 (N_13941,N_13011,N_13390);
xor U13942 (N_13942,N_13027,N_12783);
xnor U13943 (N_13943,N_12993,N_12830);
xnor U13944 (N_13944,N_13076,N_13277);
or U13945 (N_13945,N_13046,N_12881);
xnor U13946 (N_13946,N_13437,N_12873);
nor U13947 (N_13947,N_12900,N_13424);
and U13948 (N_13948,N_13219,N_12842);
or U13949 (N_13949,N_12992,N_12759);
xor U13950 (N_13950,N_12867,N_13325);
or U13951 (N_13951,N_13420,N_12991);
xor U13952 (N_13952,N_13365,N_12998);
or U13953 (N_13953,N_13490,N_13358);
and U13954 (N_13954,N_13179,N_12862);
xor U13955 (N_13955,N_13314,N_13238);
xor U13956 (N_13956,N_12781,N_13302);
and U13957 (N_13957,N_12768,N_13367);
nand U13958 (N_13958,N_13268,N_13043);
xor U13959 (N_13959,N_12863,N_13398);
or U13960 (N_13960,N_13126,N_12884);
or U13961 (N_13961,N_13455,N_13426);
nand U13962 (N_13962,N_13387,N_12949);
nand U13963 (N_13963,N_12994,N_13262);
xor U13964 (N_13964,N_13359,N_13473);
and U13965 (N_13965,N_13224,N_13128);
and U13966 (N_13966,N_13494,N_13462);
nor U13967 (N_13967,N_13365,N_13023);
nand U13968 (N_13968,N_13321,N_13198);
xor U13969 (N_13969,N_13212,N_13283);
or U13970 (N_13970,N_13044,N_13159);
xor U13971 (N_13971,N_13375,N_13487);
nor U13972 (N_13972,N_12861,N_12918);
nand U13973 (N_13973,N_13185,N_12788);
nor U13974 (N_13974,N_13481,N_13490);
nand U13975 (N_13975,N_13073,N_13300);
and U13976 (N_13976,N_12957,N_13016);
xor U13977 (N_13977,N_13097,N_12827);
nand U13978 (N_13978,N_13316,N_13172);
nor U13979 (N_13979,N_12759,N_13342);
nand U13980 (N_13980,N_13058,N_13182);
and U13981 (N_13981,N_13293,N_13156);
nor U13982 (N_13982,N_13327,N_13153);
and U13983 (N_13983,N_13241,N_13233);
or U13984 (N_13984,N_12786,N_13079);
nor U13985 (N_13985,N_13453,N_13477);
xnor U13986 (N_13986,N_13005,N_12803);
nand U13987 (N_13987,N_13090,N_13163);
nand U13988 (N_13988,N_13122,N_12874);
nand U13989 (N_13989,N_13148,N_12998);
nand U13990 (N_13990,N_13145,N_13021);
nand U13991 (N_13991,N_13278,N_13130);
nand U13992 (N_13992,N_13328,N_12764);
nor U13993 (N_13993,N_13239,N_13142);
and U13994 (N_13994,N_12939,N_13062);
nand U13995 (N_13995,N_13048,N_13215);
and U13996 (N_13996,N_13322,N_13057);
or U13997 (N_13997,N_12979,N_13362);
xor U13998 (N_13998,N_12851,N_13414);
or U13999 (N_13999,N_13088,N_13203);
xor U14000 (N_14000,N_13344,N_12966);
nand U14001 (N_14001,N_12789,N_13059);
and U14002 (N_14002,N_13345,N_13444);
xor U14003 (N_14003,N_12821,N_13485);
and U14004 (N_14004,N_12778,N_13452);
and U14005 (N_14005,N_13386,N_12971);
nand U14006 (N_14006,N_13432,N_12835);
or U14007 (N_14007,N_13287,N_13478);
or U14008 (N_14008,N_12825,N_13407);
or U14009 (N_14009,N_13148,N_13210);
nor U14010 (N_14010,N_12904,N_13322);
nand U14011 (N_14011,N_13377,N_13266);
and U14012 (N_14012,N_13087,N_13267);
nand U14013 (N_14013,N_13498,N_13295);
xor U14014 (N_14014,N_13359,N_12825);
or U14015 (N_14015,N_13330,N_13154);
nor U14016 (N_14016,N_13062,N_12922);
nand U14017 (N_14017,N_13022,N_13152);
nor U14018 (N_14018,N_12785,N_13270);
nand U14019 (N_14019,N_13411,N_12847);
and U14020 (N_14020,N_13239,N_13232);
nor U14021 (N_14021,N_13106,N_12924);
nor U14022 (N_14022,N_12957,N_13143);
nor U14023 (N_14023,N_13262,N_13268);
and U14024 (N_14024,N_13049,N_13424);
and U14025 (N_14025,N_13442,N_12865);
and U14026 (N_14026,N_13216,N_13033);
or U14027 (N_14027,N_13483,N_12900);
nor U14028 (N_14028,N_13263,N_13220);
nand U14029 (N_14029,N_13356,N_13068);
nor U14030 (N_14030,N_13029,N_13460);
xnor U14031 (N_14031,N_13436,N_13298);
and U14032 (N_14032,N_13335,N_13443);
nand U14033 (N_14033,N_12791,N_13007);
and U14034 (N_14034,N_12962,N_13231);
nor U14035 (N_14035,N_13385,N_12844);
nor U14036 (N_14036,N_13298,N_13464);
or U14037 (N_14037,N_13474,N_13197);
and U14038 (N_14038,N_13219,N_13147);
or U14039 (N_14039,N_13394,N_12911);
and U14040 (N_14040,N_12902,N_12987);
xnor U14041 (N_14041,N_13158,N_12934);
or U14042 (N_14042,N_13295,N_12783);
xnor U14043 (N_14043,N_12826,N_13479);
and U14044 (N_14044,N_13026,N_13084);
or U14045 (N_14045,N_13428,N_13250);
xor U14046 (N_14046,N_12998,N_13494);
xnor U14047 (N_14047,N_13213,N_13287);
nand U14048 (N_14048,N_12951,N_12800);
or U14049 (N_14049,N_13164,N_13088);
or U14050 (N_14050,N_13172,N_13057);
nand U14051 (N_14051,N_13003,N_13129);
or U14052 (N_14052,N_12905,N_13073);
or U14053 (N_14053,N_13294,N_13034);
nor U14054 (N_14054,N_13227,N_12961);
and U14055 (N_14055,N_13437,N_12896);
or U14056 (N_14056,N_12767,N_13367);
or U14057 (N_14057,N_13211,N_13337);
xor U14058 (N_14058,N_13473,N_13191);
xnor U14059 (N_14059,N_13408,N_13010);
xor U14060 (N_14060,N_13149,N_13008);
and U14061 (N_14061,N_13267,N_13442);
nor U14062 (N_14062,N_13036,N_12777);
nor U14063 (N_14063,N_12885,N_13208);
xnor U14064 (N_14064,N_13169,N_13390);
and U14065 (N_14065,N_13321,N_12884);
and U14066 (N_14066,N_13006,N_13208);
nor U14067 (N_14067,N_12933,N_12919);
nor U14068 (N_14068,N_12937,N_13479);
xor U14069 (N_14069,N_13414,N_13118);
nand U14070 (N_14070,N_13003,N_13111);
xor U14071 (N_14071,N_13332,N_13384);
nand U14072 (N_14072,N_12820,N_13337);
nor U14073 (N_14073,N_12784,N_13258);
xnor U14074 (N_14074,N_13234,N_13429);
and U14075 (N_14075,N_13466,N_12792);
xor U14076 (N_14076,N_13432,N_12960);
nand U14077 (N_14077,N_13246,N_13496);
or U14078 (N_14078,N_13380,N_13284);
nor U14079 (N_14079,N_13032,N_12940);
xor U14080 (N_14080,N_13393,N_13472);
or U14081 (N_14081,N_13187,N_13287);
nor U14082 (N_14082,N_13324,N_13129);
xnor U14083 (N_14083,N_13238,N_13020);
nor U14084 (N_14084,N_13259,N_13347);
xnor U14085 (N_14085,N_13309,N_12758);
or U14086 (N_14086,N_13270,N_12968);
nand U14087 (N_14087,N_13098,N_12804);
nor U14088 (N_14088,N_12953,N_12917);
or U14089 (N_14089,N_12932,N_13296);
and U14090 (N_14090,N_12813,N_13415);
xor U14091 (N_14091,N_12816,N_13358);
xor U14092 (N_14092,N_12812,N_12845);
nand U14093 (N_14093,N_13253,N_12989);
nor U14094 (N_14094,N_13363,N_13094);
nor U14095 (N_14095,N_13104,N_12999);
and U14096 (N_14096,N_13045,N_12833);
nand U14097 (N_14097,N_12843,N_13346);
or U14098 (N_14098,N_13207,N_12795);
and U14099 (N_14099,N_12869,N_12935);
or U14100 (N_14100,N_13098,N_12874);
xnor U14101 (N_14101,N_13300,N_13249);
or U14102 (N_14102,N_13441,N_13296);
nand U14103 (N_14103,N_13070,N_13491);
xnor U14104 (N_14104,N_13166,N_13323);
nand U14105 (N_14105,N_12785,N_13031);
or U14106 (N_14106,N_12833,N_13167);
nor U14107 (N_14107,N_13029,N_13196);
nand U14108 (N_14108,N_12933,N_13216);
or U14109 (N_14109,N_12958,N_13144);
and U14110 (N_14110,N_13185,N_13242);
nand U14111 (N_14111,N_13070,N_12828);
xor U14112 (N_14112,N_13146,N_12826);
xor U14113 (N_14113,N_13426,N_12872);
or U14114 (N_14114,N_13385,N_12775);
xnor U14115 (N_14115,N_13366,N_13149);
nor U14116 (N_14116,N_13390,N_13160);
and U14117 (N_14117,N_13240,N_12946);
xor U14118 (N_14118,N_12763,N_13087);
xnor U14119 (N_14119,N_13121,N_12881);
nor U14120 (N_14120,N_13486,N_13228);
and U14121 (N_14121,N_12980,N_12953);
and U14122 (N_14122,N_13169,N_13231);
nor U14123 (N_14123,N_12874,N_13217);
nor U14124 (N_14124,N_13498,N_13475);
and U14125 (N_14125,N_13019,N_12974);
nor U14126 (N_14126,N_12802,N_13241);
xor U14127 (N_14127,N_13190,N_12908);
and U14128 (N_14128,N_12919,N_12889);
or U14129 (N_14129,N_13097,N_13019);
nor U14130 (N_14130,N_12839,N_13262);
or U14131 (N_14131,N_12908,N_13232);
xor U14132 (N_14132,N_12881,N_13169);
or U14133 (N_14133,N_12935,N_12933);
nand U14134 (N_14134,N_13219,N_12965);
nand U14135 (N_14135,N_13209,N_13146);
nand U14136 (N_14136,N_12801,N_13456);
xor U14137 (N_14137,N_12774,N_12946);
xor U14138 (N_14138,N_13068,N_13228);
xor U14139 (N_14139,N_13291,N_13197);
or U14140 (N_14140,N_13064,N_13479);
xnor U14141 (N_14141,N_12927,N_12999);
nor U14142 (N_14142,N_13437,N_13446);
nand U14143 (N_14143,N_13395,N_13271);
and U14144 (N_14144,N_13425,N_13418);
or U14145 (N_14145,N_13423,N_12772);
xor U14146 (N_14146,N_12758,N_13466);
nand U14147 (N_14147,N_13097,N_13266);
nand U14148 (N_14148,N_12813,N_13400);
or U14149 (N_14149,N_13139,N_13338);
nor U14150 (N_14150,N_13490,N_12965);
xnor U14151 (N_14151,N_13107,N_13101);
and U14152 (N_14152,N_13095,N_13285);
or U14153 (N_14153,N_13474,N_13084);
xor U14154 (N_14154,N_12978,N_13272);
or U14155 (N_14155,N_12887,N_12978);
xor U14156 (N_14156,N_13355,N_13087);
nor U14157 (N_14157,N_12884,N_13123);
nor U14158 (N_14158,N_13091,N_13050);
nor U14159 (N_14159,N_13206,N_13094);
xnor U14160 (N_14160,N_12930,N_12959);
nor U14161 (N_14161,N_13196,N_13277);
nand U14162 (N_14162,N_12866,N_13470);
nor U14163 (N_14163,N_13469,N_13394);
and U14164 (N_14164,N_12800,N_13115);
nor U14165 (N_14165,N_13204,N_13474);
nor U14166 (N_14166,N_13099,N_13486);
or U14167 (N_14167,N_12980,N_13407);
nand U14168 (N_14168,N_12751,N_13383);
nor U14169 (N_14169,N_12909,N_13095);
nor U14170 (N_14170,N_12867,N_13281);
nor U14171 (N_14171,N_13181,N_13459);
xor U14172 (N_14172,N_13248,N_13333);
and U14173 (N_14173,N_13417,N_13428);
and U14174 (N_14174,N_13233,N_13146);
nor U14175 (N_14175,N_13343,N_13193);
nand U14176 (N_14176,N_12903,N_13018);
xor U14177 (N_14177,N_12991,N_13274);
and U14178 (N_14178,N_13362,N_13344);
xnor U14179 (N_14179,N_12969,N_12767);
xnor U14180 (N_14180,N_12937,N_13172);
xnor U14181 (N_14181,N_13083,N_13079);
or U14182 (N_14182,N_12985,N_13246);
nand U14183 (N_14183,N_13484,N_12957);
nor U14184 (N_14184,N_13312,N_13238);
or U14185 (N_14185,N_12775,N_13148);
and U14186 (N_14186,N_12754,N_13333);
nor U14187 (N_14187,N_13443,N_12817);
and U14188 (N_14188,N_13379,N_13230);
or U14189 (N_14189,N_13402,N_12805);
nand U14190 (N_14190,N_13173,N_12841);
nand U14191 (N_14191,N_12980,N_12905);
nor U14192 (N_14192,N_13315,N_12985);
nand U14193 (N_14193,N_13399,N_12932);
xor U14194 (N_14194,N_13404,N_13230);
or U14195 (N_14195,N_12823,N_13457);
xor U14196 (N_14196,N_12911,N_13301);
nand U14197 (N_14197,N_13041,N_13154);
or U14198 (N_14198,N_13368,N_13455);
and U14199 (N_14199,N_12960,N_12949);
nor U14200 (N_14200,N_12938,N_12981);
nand U14201 (N_14201,N_13468,N_13214);
or U14202 (N_14202,N_13180,N_13136);
and U14203 (N_14203,N_13289,N_13221);
nor U14204 (N_14204,N_12798,N_12932);
and U14205 (N_14205,N_13222,N_13179);
xor U14206 (N_14206,N_12789,N_13137);
and U14207 (N_14207,N_12793,N_13155);
xnor U14208 (N_14208,N_13239,N_12878);
or U14209 (N_14209,N_12935,N_13241);
xnor U14210 (N_14210,N_13292,N_13016);
or U14211 (N_14211,N_13417,N_13139);
and U14212 (N_14212,N_13327,N_13297);
nand U14213 (N_14213,N_13021,N_13247);
or U14214 (N_14214,N_13411,N_13190);
or U14215 (N_14215,N_12886,N_13260);
xnor U14216 (N_14216,N_13302,N_13177);
or U14217 (N_14217,N_13119,N_13026);
or U14218 (N_14218,N_13269,N_13360);
xor U14219 (N_14219,N_12971,N_13074);
and U14220 (N_14220,N_13419,N_12771);
nand U14221 (N_14221,N_13103,N_12811);
nor U14222 (N_14222,N_13106,N_13137);
or U14223 (N_14223,N_12821,N_12849);
and U14224 (N_14224,N_13237,N_13215);
or U14225 (N_14225,N_12967,N_13180);
nor U14226 (N_14226,N_12956,N_13470);
nand U14227 (N_14227,N_12923,N_13237);
nand U14228 (N_14228,N_13066,N_13228);
nor U14229 (N_14229,N_12941,N_13031);
nor U14230 (N_14230,N_12768,N_13080);
xnor U14231 (N_14231,N_13113,N_12793);
and U14232 (N_14232,N_12997,N_13439);
or U14233 (N_14233,N_12873,N_13470);
nor U14234 (N_14234,N_13109,N_13351);
and U14235 (N_14235,N_13391,N_13368);
and U14236 (N_14236,N_13156,N_12952);
nand U14237 (N_14237,N_13288,N_13270);
and U14238 (N_14238,N_13371,N_13392);
nand U14239 (N_14239,N_12950,N_13398);
and U14240 (N_14240,N_13018,N_13072);
nand U14241 (N_14241,N_13447,N_13324);
or U14242 (N_14242,N_13449,N_12769);
xor U14243 (N_14243,N_13108,N_13272);
or U14244 (N_14244,N_13238,N_12797);
nand U14245 (N_14245,N_13053,N_13329);
or U14246 (N_14246,N_12846,N_13482);
xnor U14247 (N_14247,N_12854,N_13057);
nor U14248 (N_14248,N_13027,N_12960);
nand U14249 (N_14249,N_13087,N_13325);
xor U14250 (N_14250,N_13790,N_14159);
and U14251 (N_14251,N_14101,N_13953);
and U14252 (N_14252,N_13794,N_14177);
xor U14253 (N_14253,N_14171,N_14005);
nand U14254 (N_14254,N_13771,N_14071);
and U14255 (N_14255,N_14009,N_13957);
xnor U14256 (N_14256,N_14145,N_14070);
nor U14257 (N_14257,N_13975,N_14123);
nor U14258 (N_14258,N_13591,N_13672);
xor U14259 (N_14259,N_14209,N_13639);
xnor U14260 (N_14260,N_13653,N_13802);
nand U14261 (N_14261,N_13823,N_13819);
xor U14262 (N_14262,N_13960,N_13891);
xor U14263 (N_14263,N_14248,N_13764);
or U14264 (N_14264,N_13655,N_13734);
nand U14265 (N_14265,N_13544,N_13511);
xnor U14266 (N_14266,N_13660,N_13528);
nand U14267 (N_14267,N_13913,N_14193);
nand U14268 (N_14268,N_14239,N_13645);
xnor U14269 (N_14269,N_13559,N_13889);
xor U14270 (N_14270,N_13784,N_13663);
or U14271 (N_14271,N_14048,N_13786);
nor U14272 (N_14272,N_14165,N_14115);
nor U14273 (N_14273,N_14004,N_13785);
xnor U14274 (N_14274,N_13755,N_14208);
nand U14275 (N_14275,N_13615,N_13968);
xnor U14276 (N_14276,N_13512,N_13727);
xor U14277 (N_14277,N_13848,N_14100);
and U14278 (N_14278,N_14046,N_13732);
and U14279 (N_14279,N_13509,N_13898);
nor U14280 (N_14280,N_13564,N_13661);
nand U14281 (N_14281,N_13656,N_14204);
nand U14282 (N_14282,N_13706,N_13871);
nor U14283 (N_14283,N_14189,N_13859);
nand U14284 (N_14284,N_13638,N_13557);
nand U14285 (N_14285,N_13990,N_13590);
nor U14286 (N_14286,N_13804,N_13574);
and U14287 (N_14287,N_14039,N_13515);
and U14288 (N_14288,N_13955,N_13806);
xnor U14289 (N_14289,N_13846,N_13807);
xor U14290 (N_14290,N_13626,N_14121);
or U14291 (N_14291,N_13984,N_13799);
nor U14292 (N_14292,N_13715,N_13675);
nand U14293 (N_14293,N_13780,N_13685);
nor U14294 (N_14294,N_13593,N_13912);
and U14295 (N_14295,N_13828,N_13622);
or U14296 (N_14296,N_14133,N_13772);
and U14297 (N_14297,N_13884,N_14003);
and U14298 (N_14298,N_13861,N_13890);
nor U14299 (N_14299,N_13555,N_13698);
or U14300 (N_14300,N_14215,N_14103);
and U14301 (N_14301,N_14181,N_13627);
or U14302 (N_14302,N_13707,N_13752);
nor U14303 (N_14303,N_13852,N_13911);
and U14304 (N_14304,N_13944,N_14201);
or U14305 (N_14305,N_13991,N_14116);
nor U14306 (N_14306,N_13820,N_13778);
nand U14307 (N_14307,N_14111,N_13952);
nor U14308 (N_14308,N_13974,N_13601);
nand U14309 (N_14309,N_13940,N_13554);
and U14310 (N_14310,N_13762,N_13548);
xor U14311 (N_14311,N_13980,N_13523);
or U14312 (N_14312,N_13905,N_13553);
or U14313 (N_14313,N_14151,N_13753);
nand U14314 (N_14314,N_13603,N_13666);
and U14315 (N_14315,N_13741,N_13759);
nor U14316 (N_14316,N_13943,N_13518);
and U14317 (N_14317,N_13896,N_13765);
or U14318 (N_14318,N_13572,N_14026);
and U14319 (N_14319,N_14162,N_13853);
nor U14320 (N_14320,N_13766,N_14086);
nand U14321 (N_14321,N_13678,N_13737);
or U14322 (N_14322,N_14090,N_13623);
or U14323 (N_14323,N_14170,N_14186);
and U14324 (N_14324,N_13740,N_13935);
nand U14325 (N_14325,N_14016,N_14220);
and U14326 (N_14326,N_14043,N_14141);
nand U14327 (N_14327,N_13586,N_14188);
nand U14328 (N_14328,N_14053,N_13792);
and U14329 (N_14329,N_14148,N_13878);
nand U14330 (N_14330,N_14038,N_13970);
nor U14331 (N_14331,N_14112,N_13662);
xor U14332 (N_14332,N_14032,N_13504);
nand U14333 (N_14333,N_13947,N_13691);
or U14334 (N_14334,N_14125,N_14076);
or U14335 (N_14335,N_14183,N_13526);
or U14336 (N_14336,N_13702,N_13966);
or U14337 (N_14337,N_13761,N_13694);
and U14338 (N_14338,N_13812,N_14142);
and U14339 (N_14339,N_13686,N_14191);
or U14340 (N_14340,N_13810,N_13735);
and U14341 (N_14341,N_13892,N_13893);
or U14342 (N_14342,N_13923,N_13719);
nor U14343 (N_14343,N_13883,N_13547);
xor U14344 (N_14344,N_14238,N_14099);
or U14345 (N_14345,N_13864,N_13865);
nand U14346 (N_14346,N_14221,N_14027);
nand U14347 (N_14347,N_13815,N_14054);
and U14348 (N_14348,N_13556,N_14233);
or U14349 (N_14349,N_13689,N_13900);
or U14350 (N_14350,N_13817,N_14205);
xnor U14351 (N_14351,N_13730,N_13972);
nand U14352 (N_14352,N_13500,N_14109);
nor U14353 (N_14353,N_13897,N_14033);
xor U14354 (N_14354,N_14001,N_13711);
nand U14355 (N_14355,N_13614,N_13998);
xor U14356 (N_14356,N_14018,N_14200);
nand U14357 (N_14357,N_13606,N_14147);
and U14358 (N_14358,N_13524,N_13709);
or U14359 (N_14359,N_14124,N_13566);
nor U14360 (N_14360,N_13797,N_14129);
and U14361 (N_14361,N_13543,N_13822);
nor U14362 (N_14362,N_13576,N_14045);
xor U14363 (N_14363,N_13985,N_13997);
or U14364 (N_14364,N_13522,N_13868);
or U14365 (N_14365,N_13774,N_13726);
nand U14366 (N_14366,N_14216,N_13647);
and U14367 (N_14367,N_13641,N_14120);
nand U14368 (N_14368,N_14131,N_13605);
xor U14369 (N_14369,N_13835,N_13742);
and U14370 (N_14370,N_13650,N_14047);
nand U14371 (N_14371,N_13869,N_13830);
nand U14372 (N_14372,N_13783,N_14073);
nor U14373 (N_14373,N_13542,N_13673);
xor U14374 (N_14374,N_13775,N_14069);
xor U14375 (N_14375,N_13757,N_13763);
xnor U14376 (N_14376,N_14114,N_14021);
and U14377 (N_14377,N_13959,N_13800);
and U14378 (N_14378,N_13825,N_14113);
nand U14379 (N_14379,N_13872,N_13895);
or U14380 (N_14380,N_14044,N_13643);
nand U14381 (N_14381,N_14082,N_13696);
or U14382 (N_14382,N_14227,N_13979);
xor U14383 (N_14383,N_13803,N_13926);
and U14384 (N_14384,N_14138,N_13527);
nor U14385 (N_14385,N_13733,N_13722);
or U14386 (N_14386,N_14210,N_14206);
xnor U14387 (N_14387,N_13779,N_13560);
and U14388 (N_14388,N_13978,N_14107);
nand U14389 (N_14389,N_14173,N_13743);
nand U14390 (N_14390,N_13705,N_13613);
nand U14391 (N_14391,N_13791,N_13608);
nand U14392 (N_14392,N_14187,N_14011);
or U14393 (N_14393,N_14196,N_13862);
nand U14394 (N_14394,N_13592,N_14092);
and U14395 (N_14395,N_14185,N_13583);
or U14396 (N_14396,N_13716,N_13501);
or U14397 (N_14397,N_14058,N_14085);
xnor U14398 (N_14398,N_14158,N_14130);
and U14399 (N_14399,N_13637,N_13899);
or U14400 (N_14400,N_14197,N_14153);
nor U14401 (N_14401,N_13505,N_13551);
or U14402 (N_14402,N_13721,N_13876);
or U14403 (N_14403,N_14091,N_13939);
and U14404 (N_14404,N_14061,N_14110);
or U14405 (N_14405,N_13826,N_13594);
xnor U14406 (N_14406,N_13860,N_14140);
nand U14407 (N_14407,N_13531,N_13677);
nor U14408 (N_14408,N_14034,N_13747);
nor U14409 (N_14409,N_13654,N_13886);
nand U14410 (N_14410,N_14022,N_13834);
nor U14411 (N_14411,N_14237,N_14137);
and U14412 (N_14412,N_13633,N_13618);
xnor U14413 (N_14413,N_13649,N_13910);
nor U14414 (N_14414,N_13628,N_14156);
and U14415 (N_14415,N_14136,N_13679);
and U14416 (N_14416,N_13611,N_13983);
nand U14417 (N_14417,N_14154,N_13934);
nor U14418 (N_14418,N_13575,N_13971);
xnor U14419 (N_14419,N_13680,N_14064);
nand U14420 (N_14420,N_13665,N_14066);
nand U14421 (N_14421,N_14134,N_13840);
nand U14422 (N_14422,N_14228,N_14122);
nor U14423 (N_14423,N_14169,N_13933);
or U14424 (N_14424,N_13577,N_13658);
and U14425 (N_14425,N_13671,N_13648);
nand U14426 (N_14426,N_13728,N_14242);
nor U14427 (N_14427,N_14119,N_13915);
or U14428 (N_14428,N_13579,N_14176);
xnor U14429 (N_14429,N_13720,N_14231);
nor U14430 (N_14430,N_13877,N_14015);
or U14431 (N_14431,N_13824,N_14190);
nor U14432 (N_14432,N_13965,N_13992);
or U14433 (N_14433,N_13703,N_14094);
or U14434 (N_14434,N_13525,N_13813);
xor U14435 (N_14435,N_14088,N_13712);
nand U14436 (N_14436,N_14065,N_13602);
or U14437 (N_14437,N_13773,N_13777);
or U14438 (N_14438,N_13903,N_13636);
xor U14439 (N_14439,N_14063,N_13536);
or U14440 (N_14440,N_13514,N_13558);
xor U14441 (N_14441,N_13879,N_13634);
nor U14442 (N_14442,N_13600,N_14075);
and U14443 (N_14443,N_13798,N_14182);
nand U14444 (N_14444,N_14059,N_14017);
nor U14445 (N_14445,N_13858,N_13616);
nor U14446 (N_14446,N_14164,N_13760);
nor U14447 (N_14447,N_13863,N_13919);
and U14448 (N_14448,N_13659,N_14068);
or U14449 (N_14449,N_14178,N_13967);
nor U14450 (N_14450,N_13539,N_13838);
or U14451 (N_14451,N_13697,N_14002);
xnor U14452 (N_14452,N_14050,N_13669);
and U14453 (N_14453,N_13776,N_13521);
xor U14454 (N_14454,N_13928,N_13738);
or U14455 (N_14455,N_13744,N_13963);
nor U14456 (N_14456,N_13842,N_13612);
nand U14457 (N_14457,N_13750,N_13567);
nor U14458 (N_14458,N_14230,N_14249);
and U14459 (N_14459,N_14149,N_14105);
and U14460 (N_14460,N_14223,N_13570);
and U14461 (N_14461,N_13902,N_13731);
xor U14462 (N_14462,N_14037,N_13552);
nand U14463 (N_14463,N_13918,N_14235);
nor U14464 (N_14464,N_14042,N_14020);
and U14465 (N_14465,N_14040,N_14051);
and U14466 (N_14466,N_13710,N_13629);
and U14467 (N_14467,N_13958,N_14072);
xnor U14468 (N_14468,N_14095,N_13517);
and U14469 (N_14469,N_13580,N_13847);
nand U14470 (N_14470,N_13818,N_14207);
nor U14471 (N_14471,N_13725,N_13969);
nor U14472 (N_14472,N_13751,N_13909);
or U14473 (N_14473,N_13922,N_13881);
or U14474 (N_14474,N_13585,N_13945);
xnor U14475 (N_14475,N_14117,N_13758);
xor U14476 (N_14476,N_13788,N_13995);
nor U14477 (N_14477,N_13831,N_13569);
nor U14478 (N_14478,N_14087,N_14195);
and U14479 (N_14479,N_14055,N_13787);
nor U14480 (N_14480,N_13956,N_13814);
or U14481 (N_14481,N_14062,N_13924);
nor U14482 (N_14482,N_14180,N_14166);
or U14483 (N_14483,N_13836,N_13635);
nand U14484 (N_14484,N_13982,N_14160);
nand U14485 (N_14485,N_14078,N_13821);
nand U14486 (N_14486,N_14202,N_13855);
nor U14487 (N_14487,N_13699,N_13851);
xor U14488 (N_14488,N_13519,N_14143);
xor U14489 (N_14489,N_13988,N_13816);
xor U14490 (N_14490,N_13961,N_14218);
nand U14491 (N_14491,N_13989,N_13901);
and U14492 (N_14492,N_13598,N_13950);
or U14493 (N_14493,N_13739,N_13805);
nor U14494 (N_14494,N_13954,N_13704);
nor U14495 (N_14495,N_13565,N_13692);
nand U14496 (N_14496,N_14139,N_13561);
or U14497 (N_14497,N_13538,N_13829);
nor U14498 (N_14498,N_14175,N_13917);
xor U14499 (N_14499,N_13857,N_13885);
nor U14500 (N_14500,N_13888,N_13746);
and U14501 (N_14501,N_14184,N_13941);
nor U14502 (N_14502,N_14041,N_13768);
nand U14503 (N_14503,N_13964,N_13651);
xnor U14504 (N_14504,N_14052,N_13845);
xor U14505 (N_14505,N_14098,N_13529);
nand U14506 (N_14506,N_13748,N_14106);
or U14507 (N_14507,N_13503,N_13767);
xnor U14508 (N_14508,N_13808,N_14012);
and U14509 (N_14509,N_13630,N_14225);
nand U14510 (N_14510,N_13880,N_14127);
nand U14511 (N_14511,N_13921,N_14203);
nor U14512 (N_14512,N_13723,N_13793);
nand U14513 (N_14513,N_13502,N_13621);
nand U14514 (N_14514,N_13789,N_13907);
or U14515 (N_14515,N_13644,N_14030);
nand U14516 (N_14516,N_13535,N_13582);
and U14517 (N_14517,N_14192,N_13631);
nand U14518 (N_14518,N_13596,N_13796);
or U14519 (N_14519,N_13801,N_14028);
xnor U14520 (N_14520,N_13625,N_14146);
xor U14521 (N_14521,N_14007,N_13908);
nor U14522 (N_14522,N_13942,N_14243);
and U14523 (N_14523,N_14013,N_13508);
nor U14524 (N_14524,N_14157,N_14161);
or U14525 (N_14525,N_14081,N_14144);
xor U14526 (N_14526,N_13640,N_13973);
xor U14527 (N_14527,N_13676,N_13713);
or U14528 (N_14528,N_14168,N_13770);
or U14529 (N_14529,N_13581,N_13718);
or U14530 (N_14530,N_13510,N_14104);
xor U14531 (N_14531,N_14135,N_13904);
and U14532 (N_14532,N_13930,N_13916);
or U14533 (N_14533,N_13782,N_14067);
or U14534 (N_14534,N_13674,N_13646);
nor U14535 (N_14535,N_13701,N_14049);
and U14536 (N_14536,N_13599,N_13533);
nand U14537 (N_14537,N_13549,N_13589);
and U14538 (N_14538,N_13987,N_13513);
nand U14539 (N_14539,N_13850,N_13695);
nor U14540 (N_14540,N_14213,N_14240);
and U14541 (N_14541,N_14031,N_13620);
nor U14542 (N_14542,N_13670,N_13844);
nand U14543 (N_14543,N_14172,N_13516);
nor U14544 (N_14544,N_13948,N_14163);
xor U14545 (N_14545,N_13882,N_14096);
and U14546 (N_14546,N_14089,N_13693);
nor U14547 (N_14547,N_14212,N_14057);
or U14548 (N_14548,N_14010,N_14167);
and U14549 (N_14549,N_13563,N_13936);
and U14550 (N_14550,N_13931,N_13520);
xor U14551 (N_14551,N_14214,N_13914);
nor U14552 (N_14552,N_13932,N_14080);
nor U14553 (N_14553,N_14102,N_14150);
xor U14554 (N_14554,N_13687,N_13700);
or U14555 (N_14555,N_14083,N_13745);
nor U14556 (N_14556,N_13873,N_13999);
nor U14557 (N_14557,N_14226,N_13610);
or U14558 (N_14558,N_14077,N_13854);
and U14559 (N_14559,N_14118,N_13977);
or U14560 (N_14560,N_13870,N_13927);
nor U14561 (N_14561,N_13587,N_13920);
nand U14562 (N_14562,N_13993,N_13976);
and U14563 (N_14563,N_14222,N_13684);
xor U14564 (N_14564,N_13595,N_13597);
nor U14565 (N_14565,N_14232,N_14084);
nand U14566 (N_14566,N_13534,N_14006);
nand U14567 (N_14567,N_13832,N_14241);
and U14568 (N_14568,N_14245,N_13874);
nor U14569 (N_14569,N_14097,N_13867);
nor U14570 (N_14570,N_13736,N_14056);
nor U14571 (N_14571,N_14211,N_14024);
xor U14572 (N_14572,N_14000,N_13754);
nand U14573 (N_14573,N_13540,N_13624);
or U14574 (N_14574,N_13937,N_13781);
nor U14575 (N_14575,N_13584,N_13568);
and U14576 (N_14576,N_14229,N_14219);
or U14577 (N_14577,N_13550,N_13530);
nand U14578 (N_14578,N_13833,N_13690);
xor U14579 (N_14579,N_13609,N_13607);
or U14580 (N_14580,N_14025,N_13769);
xnor U14581 (N_14581,N_14019,N_13546);
xnor U14582 (N_14582,N_14060,N_13652);
nand U14583 (N_14583,N_14132,N_13841);
xnor U14584 (N_14584,N_13507,N_14217);
nand U14585 (N_14585,N_14128,N_13951);
and U14586 (N_14586,N_13827,N_14247);
nand U14587 (N_14587,N_13729,N_13894);
xor U14588 (N_14588,N_13604,N_13724);
and U14589 (N_14589,N_13619,N_13996);
nor U14590 (N_14590,N_14023,N_13632);
xor U14591 (N_14591,N_13938,N_13962);
and U14592 (N_14592,N_13929,N_13875);
and U14593 (N_14593,N_14014,N_14224);
nor U14594 (N_14594,N_13749,N_14008);
or U14595 (N_14595,N_13811,N_14035);
xor U14596 (N_14596,N_13537,N_14199);
and U14597 (N_14597,N_13949,N_14108);
or U14598 (N_14598,N_13708,N_13856);
or U14599 (N_14599,N_13849,N_13795);
nor U14600 (N_14600,N_14126,N_13986);
xor U14601 (N_14601,N_13682,N_13617);
nand U14602 (N_14602,N_13545,N_14198);
nand U14603 (N_14603,N_13981,N_13756);
or U14604 (N_14604,N_14244,N_14179);
and U14605 (N_14605,N_13887,N_13839);
nand U14606 (N_14606,N_14194,N_14029);
nand U14607 (N_14607,N_13946,N_13562);
and U14608 (N_14608,N_13837,N_14074);
or U14609 (N_14609,N_14234,N_14246);
xnor U14610 (N_14610,N_13925,N_13668);
nor U14611 (N_14611,N_13571,N_13717);
or U14612 (N_14612,N_13657,N_13541);
xnor U14613 (N_14613,N_13683,N_13809);
or U14614 (N_14614,N_13667,N_14152);
and U14615 (N_14615,N_13642,N_13906);
and U14616 (N_14616,N_13681,N_13664);
nor U14617 (N_14617,N_13994,N_13688);
nor U14618 (N_14618,N_14236,N_14093);
xnor U14619 (N_14619,N_14174,N_13843);
xor U14620 (N_14620,N_13573,N_13506);
nand U14621 (N_14621,N_13578,N_13532);
and U14622 (N_14622,N_14036,N_14155);
and U14623 (N_14623,N_13714,N_13866);
nand U14624 (N_14624,N_13588,N_14079);
nand U14625 (N_14625,N_13702,N_13744);
or U14626 (N_14626,N_13780,N_13517);
or U14627 (N_14627,N_14211,N_13536);
xnor U14628 (N_14628,N_14033,N_13981);
xnor U14629 (N_14629,N_13726,N_13533);
nand U14630 (N_14630,N_13580,N_13935);
and U14631 (N_14631,N_13688,N_13758);
or U14632 (N_14632,N_14080,N_13862);
nand U14633 (N_14633,N_13583,N_14142);
nor U14634 (N_14634,N_13695,N_14106);
or U14635 (N_14635,N_13762,N_13616);
xor U14636 (N_14636,N_14058,N_14079);
and U14637 (N_14637,N_13680,N_13919);
or U14638 (N_14638,N_13677,N_13755);
nand U14639 (N_14639,N_13723,N_13785);
nor U14640 (N_14640,N_13856,N_13681);
xor U14641 (N_14641,N_13959,N_13743);
nor U14642 (N_14642,N_14123,N_14131);
or U14643 (N_14643,N_13571,N_13868);
and U14644 (N_14644,N_13906,N_13926);
xnor U14645 (N_14645,N_13992,N_13787);
nor U14646 (N_14646,N_14067,N_13599);
nand U14647 (N_14647,N_14011,N_13903);
nand U14648 (N_14648,N_13967,N_13901);
nor U14649 (N_14649,N_13876,N_13591);
or U14650 (N_14650,N_14198,N_13572);
or U14651 (N_14651,N_13761,N_13645);
nor U14652 (N_14652,N_13736,N_13840);
xor U14653 (N_14653,N_14090,N_14006);
or U14654 (N_14654,N_14222,N_13774);
and U14655 (N_14655,N_14017,N_13747);
nor U14656 (N_14656,N_14013,N_13705);
nand U14657 (N_14657,N_14146,N_13996);
or U14658 (N_14658,N_14024,N_13620);
or U14659 (N_14659,N_14094,N_13907);
xnor U14660 (N_14660,N_13909,N_14048);
xnor U14661 (N_14661,N_14023,N_14204);
xnor U14662 (N_14662,N_13975,N_14103);
and U14663 (N_14663,N_13898,N_13792);
or U14664 (N_14664,N_14060,N_13607);
nor U14665 (N_14665,N_13770,N_14054);
and U14666 (N_14666,N_13554,N_13995);
nor U14667 (N_14667,N_13638,N_13753);
or U14668 (N_14668,N_13890,N_13904);
nand U14669 (N_14669,N_14011,N_13658);
nor U14670 (N_14670,N_13608,N_14053);
nor U14671 (N_14671,N_14238,N_14085);
nor U14672 (N_14672,N_13709,N_14057);
or U14673 (N_14673,N_13502,N_14102);
and U14674 (N_14674,N_14125,N_14192);
xnor U14675 (N_14675,N_13715,N_14083);
nand U14676 (N_14676,N_13891,N_14031);
nand U14677 (N_14677,N_13845,N_14207);
nand U14678 (N_14678,N_13964,N_13520);
xor U14679 (N_14679,N_13776,N_13566);
and U14680 (N_14680,N_13540,N_14085);
and U14681 (N_14681,N_13639,N_14108);
xor U14682 (N_14682,N_13905,N_13866);
xnor U14683 (N_14683,N_14113,N_14176);
and U14684 (N_14684,N_13680,N_13814);
or U14685 (N_14685,N_13520,N_13734);
or U14686 (N_14686,N_13998,N_14247);
and U14687 (N_14687,N_14118,N_13652);
or U14688 (N_14688,N_14226,N_13994);
xnor U14689 (N_14689,N_13529,N_14104);
or U14690 (N_14690,N_13955,N_14207);
nand U14691 (N_14691,N_13677,N_13660);
or U14692 (N_14692,N_13696,N_13832);
and U14693 (N_14693,N_13900,N_14158);
or U14694 (N_14694,N_13723,N_14136);
nor U14695 (N_14695,N_13933,N_13892);
nand U14696 (N_14696,N_14059,N_13700);
xnor U14697 (N_14697,N_13848,N_13867);
nand U14698 (N_14698,N_13716,N_14188);
xor U14699 (N_14699,N_13807,N_14068);
nor U14700 (N_14700,N_13765,N_13771);
xnor U14701 (N_14701,N_13527,N_14107);
or U14702 (N_14702,N_13512,N_13729);
xor U14703 (N_14703,N_13635,N_13582);
nor U14704 (N_14704,N_14161,N_14178);
xnor U14705 (N_14705,N_13516,N_14003);
or U14706 (N_14706,N_13654,N_14064);
and U14707 (N_14707,N_14073,N_13695);
and U14708 (N_14708,N_13622,N_13907);
and U14709 (N_14709,N_13857,N_14065);
nor U14710 (N_14710,N_13893,N_13679);
xnor U14711 (N_14711,N_14243,N_14086);
xor U14712 (N_14712,N_13781,N_13554);
nor U14713 (N_14713,N_13877,N_13597);
and U14714 (N_14714,N_13780,N_13819);
xor U14715 (N_14715,N_13787,N_14070);
nand U14716 (N_14716,N_13752,N_14029);
nand U14717 (N_14717,N_13888,N_14219);
and U14718 (N_14718,N_13821,N_14144);
and U14719 (N_14719,N_13741,N_13948);
xor U14720 (N_14720,N_14169,N_13963);
or U14721 (N_14721,N_13536,N_13539);
nand U14722 (N_14722,N_14075,N_13578);
and U14723 (N_14723,N_13590,N_13950);
xor U14724 (N_14724,N_13809,N_13572);
nor U14725 (N_14725,N_13859,N_13786);
nor U14726 (N_14726,N_14045,N_13930);
and U14727 (N_14727,N_14115,N_14019);
and U14728 (N_14728,N_13905,N_13949);
nand U14729 (N_14729,N_14108,N_13695);
or U14730 (N_14730,N_14014,N_13814);
or U14731 (N_14731,N_13568,N_13669);
or U14732 (N_14732,N_14055,N_13578);
nor U14733 (N_14733,N_13945,N_13745);
and U14734 (N_14734,N_13637,N_13521);
and U14735 (N_14735,N_14029,N_13589);
and U14736 (N_14736,N_13516,N_13810);
nor U14737 (N_14737,N_13936,N_13732);
and U14738 (N_14738,N_13518,N_13515);
nor U14739 (N_14739,N_13898,N_13566);
and U14740 (N_14740,N_13687,N_14242);
or U14741 (N_14741,N_13899,N_13833);
nor U14742 (N_14742,N_13659,N_13704);
and U14743 (N_14743,N_13845,N_13543);
xnor U14744 (N_14744,N_13542,N_14014);
and U14745 (N_14745,N_14119,N_13999);
xnor U14746 (N_14746,N_13580,N_13808);
and U14747 (N_14747,N_13545,N_13877);
nand U14748 (N_14748,N_13786,N_14058);
xor U14749 (N_14749,N_14112,N_14211);
nand U14750 (N_14750,N_13631,N_13715);
or U14751 (N_14751,N_13513,N_13907);
or U14752 (N_14752,N_13575,N_13892);
nor U14753 (N_14753,N_13775,N_14094);
nand U14754 (N_14754,N_14186,N_14157);
nor U14755 (N_14755,N_13542,N_14007);
and U14756 (N_14756,N_13694,N_13820);
and U14757 (N_14757,N_13742,N_13515);
and U14758 (N_14758,N_14085,N_13670);
xor U14759 (N_14759,N_13502,N_14076);
xor U14760 (N_14760,N_14088,N_13897);
or U14761 (N_14761,N_14227,N_13704);
and U14762 (N_14762,N_13756,N_13925);
or U14763 (N_14763,N_14142,N_13512);
and U14764 (N_14764,N_14003,N_14050);
nor U14765 (N_14765,N_14105,N_13627);
or U14766 (N_14766,N_14030,N_14175);
and U14767 (N_14767,N_14180,N_13956);
or U14768 (N_14768,N_13968,N_13619);
nor U14769 (N_14769,N_14157,N_13816);
nor U14770 (N_14770,N_14070,N_13542);
or U14771 (N_14771,N_13791,N_13962);
nand U14772 (N_14772,N_14116,N_14019);
xnor U14773 (N_14773,N_13976,N_13951);
and U14774 (N_14774,N_13560,N_13819);
and U14775 (N_14775,N_13879,N_13654);
nand U14776 (N_14776,N_14203,N_14071);
nand U14777 (N_14777,N_13739,N_14225);
or U14778 (N_14778,N_13923,N_13728);
xnor U14779 (N_14779,N_13786,N_14209);
nand U14780 (N_14780,N_13684,N_13590);
xor U14781 (N_14781,N_14236,N_13695);
or U14782 (N_14782,N_13621,N_13659);
nand U14783 (N_14783,N_13839,N_14187);
nor U14784 (N_14784,N_13654,N_14050);
nor U14785 (N_14785,N_13877,N_14016);
nor U14786 (N_14786,N_13990,N_13905);
and U14787 (N_14787,N_13650,N_14159);
or U14788 (N_14788,N_14098,N_13942);
xnor U14789 (N_14789,N_14178,N_13626);
xor U14790 (N_14790,N_14205,N_13692);
nor U14791 (N_14791,N_13987,N_13887);
or U14792 (N_14792,N_13550,N_14040);
xor U14793 (N_14793,N_14073,N_13879);
nand U14794 (N_14794,N_13986,N_13779);
and U14795 (N_14795,N_14003,N_14058);
and U14796 (N_14796,N_13585,N_14085);
or U14797 (N_14797,N_13885,N_14063);
nor U14798 (N_14798,N_14145,N_13788);
nor U14799 (N_14799,N_14058,N_14158);
and U14800 (N_14800,N_14194,N_14169);
nor U14801 (N_14801,N_13808,N_13563);
or U14802 (N_14802,N_14052,N_13525);
xnor U14803 (N_14803,N_14169,N_14022);
nor U14804 (N_14804,N_14018,N_13868);
nand U14805 (N_14805,N_13877,N_13815);
nand U14806 (N_14806,N_14136,N_14187);
xnor U14807 (N_14807,N_14136,N_14182);
nand U14808 (N_14808,N_13794,N_14234);
or U14809 (N_14809,N_13970,N_13573);
nand U14810 (N_14810,N_13761,N_13669);
nor U14811 (N_14811,N_13596,N_14248);
or U14812 (N_14812,N_14108,N_14046);
nor U14813 (N_14813,N_13638,N_14206);
and U14814 (N_14814,N_13544,N_14025);
or U14815 (N_14815,N_13828,N_13844);
nand U14816 (N_14816,N_13612,N_14028);
nor U14817 (N_14817,N_14217,N_13835);
xnor U14818 (N_14818,N_13529,N_13868);
xor U14819 (N_14819,N_13674,N_13954);
nor U14820 (N_14820,N_14192,N_13594);
nand U14821 (N_14821,N_13572,N_14089);
xor U14822 (N_14822,N_14051,N_13970);
and U14823 (N_14823,N_14244,N_13550);
xor U14824 (N_14824,N_13911,N_13990);
nor U14825 (N_14825,N_13901,N_14128);
xor U14826 (N_14826,N_13859,N_13922);
nor U14827 (N_14827,N_14014,N_13979);
nor U14828 (N_14828,N_13626,N_13686);
nor U14829 (N_14829,N_14214,N_14028);
or U14830 (N_14830,N_13738,N_14004);
and U14831 (N_14831,N_14190,N_14160);
and U14832 (N_14832,N_13567,N_13568);
or U14833 (N_14833,N_14027,N_13688);
and U14834 (N_14834,N_14161,N_13608);
nor U14835 (N_14835,N_14236,N_13950);
nor U14836 (N_14836,N_13951,N_13618);
or U14837 (N_14837,N_13519,N_14119);
nand U14838 (N_14838,N_13578,N_14039);
or U14839 (N_14839,N_13802,N_13915);
nand U14840 (N_14840,N_13791,N_14079);
and U14841 (N_14841,N_14249,N_13806);
nand U14842 (N_14842,N_13877,N_14045);
nor U14843 (N_14843,N_13841,N_14034);
or U14844 (N_14844,N_13862,N_13961);
nor U14845 (N_14845,N_13648,N_13755);
and U14846 (N_14846,N_13681,N_14082);
and U14847 (N_14847,N_14204,N_13983);
nand U14848 (N_14848,N_13830,N_14107);
nor U14849 (N_14849,N_14119,N_13910);
xor U14850 (N_14850,N_13703,N_13885);
and U14851 (N_14851,N_13992,N_13675);
xor U14852 (N_14852,N_14044,N_13771);
xnor U14853 (N_14853,N_14047,N_14154);
nor U14854 (N_14854,N_13824,N_14236);
nor U14855 (N_14855,N_14112,N_13978);
and U14856 (N_14856,N_13851,N_13665);
or U14857 (N_14857,N_14129,N_14185);
nor U14858 (N_14858,N_14096,N_13911);
nor U14859 (N_14859,N_14120,N_13770);
and U14860 (N_14860,N_13674,N_14195);
nand U14861 (N_14861,N_13668,N_14014);
or U14862 (N_14862,N_14061,N_13789);
nand U14863 (N_14863,N_13898,N_13777);
or U14864 (N_14864,N_14020,N_13702);
and U14865 (N_14865,N_14005,N_14133);
or U14866 (N_14866,N_13682,N_13821);
nor U14867 (N_14867,N_13522,N_14024);
xor U14868 (N_14868,N_14129,N_13823);
or U14869 (N_14869,N_14119,N_14064);
nand U14870 (N_14870,N_13580,N_14134);
nor U14871 (N_14871,N_14044,N_13892);
and U14872 (N_14872,N_13725,N_13740);
or U14873 (N_14873,N_14209,N_14143);
or U14874 (N_14874,N_13641,N_14099);
nor U14875 (N_14875,N_13974,N_14225);
nor U14876 (N_14876,N_14220,N_13850);
or U14877 (N_14877,N_14101,N_14157);
and U14878 (N_14878,N_13934,N_13928);
or U14879 (N_14879,N_13937,N_13772);
and U14880 (N_14880,N_13772,N_14083);
and U14881 (N_14881,N_14204,N_13589);
and U14882 (N_14882,N_14087,N_13876);
and U14883 (N_14883,N_14019,N_14079);
or U14884 (N_14884,N_13576,N_13891);
or U14885 (N_14885,N_13763,N_13729);
nand U14886 (N_14886,N_13729,N_14035);
and U14887 (N_14887,N_14146,N_14128);
xnor U14888 (N_14888,N_14068,N_13815);
or U14889 (N_14889,N_13581,N_13804);
nand U14890 (N_14890,N_14138,N_13858);
nor U14891 (N_14891,N_14046,N_13527);
or U14892 (N_14892,N_13821,N_13645);
and U14893 (N_14893,N_13866,N_13959);
and U14894 (N_14894,N_14192,N_14001);
or U14895 (N_14895,N_13546,N_13948);
nor U14896 (N_14896,N_13837,N_13562);
and U14897 (N_14897,N_14154,N_13977);
xnor U14898 (N_14898,N_13997,N_14023);
xnor U14899 (N_14899,N_13624,N_13866);
nor U14900 (N_14900,N_14013,N_13796);
and U14901 (N_14901,N_13510,N_13573);
nor U14902 (N_14902,N_14204,N_13837);
nand U14903 (N_14903,N_14044,N_13733);
or U14904 (N_14904,N_13920,N_14147);
and U14905 (N_14905,N_13589,N_13853);
nor U14906 (N_14906,N_14139,N_13643);
and U14907 (N_14907,N_14080,N_13719);
and U14908 (N_14908,N_14033,N_14112);
nor U14909 (N_14909,N_14103,N_14085);
xnor U14910 (N_14910,N_13504,N_14158);
nand U14911 (N_14911,N_13772,N_13576);
nand U14912 (N_14912,N_14183,N_14018);
and U14913 (N_14913,N_13566,N_13510);
nand U14914 (N_14914,N_14081,N_13847);
xor U14915 (N_14915,N_13623,N_13965);
and U14916 (N_14916,N_13976,N_14071);
and U14917 (N_14917,N_13898,N_14200);
nand U14918 (N_14918,N_13597,N_14107);
nand U14919 (N_14919,N_14139,N_13506);
and U14920 (N_14920,N_13881,N_13995);
nand U14921 (N_14921,N_13810,N_13948);
xor U14922 (N_14922,N_13866,N_13876);
nand U14923 (N_14923,N_14156,N_14115);
nor U14924 (N_14924,N_14188,N_13767);
nor U14925 (N_14925,N_13546,N_13643);
xnor U14926 (N_14926,N_13591,N_14068);
xor U14927 (N_14927,N_13509,N_13946);
or U14928 (N_14928,N_13881,N_14227);
xor U14929 (N_14929,N_13806,N_13942);
xnor U14930 (N_14930,N_13609,N_13912);
xnor U14931 (N_14931,N_13613,N_13676);
nand U14932 (N_14932,N_14166,N_13654);
and U14933 (N_14933,N_13747,N_13535);
nand U14934 (N_14934,N_13509,N_13582);
nor U14935 (N_14935,N_13806,N_13823);
xor U14936 (N_14936,N_13576,N_13686);
and U14937 (N_14937,N_14116,N_13990);
and U14938 (N_14938,N_13826,N_14218);
nand U14939 (N_14939,N_13994,N_14163);
xor U14940 (N_14940,N_14013,N_13632);
and U14941 (N_14941,N_13683,N_13581);
nor U14942 (N_14942,N_13786,N_13837);
nor U14943 (N_14943,N_13808,N_14147);
nor U14944 (N_14944,N_13835,N_13727);
or U14945 (N_14945,N_13580,N_13688);
nor U14946 (N_14946,N_13942,N_13830);
nand U14947 (N_14947,N_13501,N_13699);
nor U14948 (N_14948,N_14192,N_14212);
or U14949 (N_14949,N_13938,N_13782);
and U14950 (N_14950,N_13812,N_13752);
nand U14951 (N_14951,N_13659,N_14199);
or U14952 (N_14952,N_14109,N_14232);
nor U14953 (N_14953,N_14137,N_14016);
xnor U14954 (N_14954,N_13888,N_13883);
and U14955 (N_14955,N_13945,N_14054);
or U14956 (N_14956,N_13825,N_14000);
and U14957 (N_14957,N_13822,N_13717);
and U14958 (N_14958,N_14147,N_14125);
nor U14959 (N_14959,N_13954,N_13843);
xnor U14960 (N_14960,N_14008,N_13813);
xor U14961 (N_14961,N_13595,N_13690);
or U14962 (N_14962,N_14188,N_14029);
or U14963 (N_14963,N_13536,N_14024);
nor U14964 (N_14964,N_13637,N_14134);
nand U14965 (N_14965,N_14095,N_14189);
xnor U14966 (N_14966,N_13969,N_13561);
and U14967 (N_14967,N_13810,N_13614);
xnor U14968 (N_14968,N_13605,N_14133);
or U14969 (N_14969,N_13765,N_13531);
nand U14970 (N_14970,N_13558,N_13568);
or U14971 (N_14971,N_13759,N_14009);
xor U14972 (N_14972,N_13601,N_14105);
or U14973 (N_14973,N_13679,N_13809);
nor U14974 (N_14974,N_13614,N_13755);
xor U14975 (N_14975,N_14133,N_13818);
or U14976 (N_14976,N_13971,N_13774);
xor U14977 (N_14977,N_14063,N_13692);
nand U14978 (N_14978,N_14045,N_14190);
nand U14979 (N_14979,N_13936,N_13932);
and U14980 (N_14980,N_13540,N_13814);
nor U14981 (N_14981,N_14235,N_14049);
nor U14982 (N_14982,N_14140,N_13744);
xnor U14983 (N_14983,N_13989,N_13819);
and U14984 (N_14984,N_13647,N_13699);
and U14985 (N_14985,N_13913,N_13828);
nor U14986 (N_14986,N_13794,N_14182);
and U14987 (N_14987,N_13825,N_13686);
nand U14988 (N_14988,N_14239,N_13839);
or U14989 (N_14989,N_14000,N_14246);
or U14990 (N_14990,N_14084,N_13740);
or U14991 (N_14991,N_13812,N_13845);
xor U14992 (N_14992,N_14246,N_14216);
or U14993 (N_14993,N_14101,N_14137);
and U14994 (N_14994,N_14007,N_13856);
and U14995 (N_14995,N_14091,N_13503);
nand U14996 (N_14996,N_13787,N_14033);
or U14997 (N_14997,N_13769,N_13995);
nor U14998 (N_14998,N_14246,N_13851);
nor U14999 (N_14999,N_13995,N_13713);
nand UO_0 (O_0,N_14499,N_14776);
xnor UO_1 (O_1,N_14384,N_14362);
or UO_2 (O_2,N_14507,N_14434);
nor UO_3 (O_3,N_14536,N_14686);
xnor UO_4 (O_4,N_14259,N_14888);
and UO_5 (O_5,N_14967,N_14291);
xnor UO_6 (O_6,N_14335,N_14938);
xnor UO_7 (O_7,N_14425,N_14275);
nor UO_8 (O_8,N_14783,N_14504);
nor UO_9 (O_9,N_14266,N_14726);
and UO_10 (O_10,N_14803,N_14532);
or UO_11 (O_11,N_14908,N_14325);
xnor UO_12 (O_12,N_14278,N_14934);
nand UO_13 (O_13,N_14792,N_14882);
xor UO_14 (O_14,N_14415,N_14595);
nor UO_15 (O_15,N_14963,N_14703);
nor UO_16 (O_16,N_14736,N_14567);
nor UO_17 (O_17,N_14288,N_14483);
and UO_18 (O_18,N_14932,N_14765);
nor UO_19 (O_19,N_14825,N_14323);
and UO_20 (O_20,N_14639,N_14664);
nand UO_21 (O_21,N_14740,N_14894);
nor UO_22 (O_22,N_14777,N_14674);
xor UO_23 (O_23,N_14443,N_14535);
nand UO_24 (O_24,N_14844,N_14402);
or UO_25 (O_25,N_14555,N_14418);
and UO_26 (O_26,N_14807,N_14702);
xnor UO_27 (O_27,N_14472,N_14440);
and UO_28 (O_28,N_14345,N_14978);
or UO_29 (O_29,N_14837,N_14454);
xnor UO_30 (O_30,N_14294,N_14329);
xor UO_31 (O_31,N_14917,N_14606);
or UO_32 (O_32,N_14574,N_14871);
nor UO_33 (O_33,N_14983,N_14289);
xor UO_34 (O_34,N_14467,N_14557);
xnor UO_35 (O_35,N_14346,N_14993);
nand UO_36 (O_36,N_14945,N_14793);
or UO_37 (O_37,N_14263,N_14265);
nand UO_38 (O_38,N_14319,N_14794);
and UO_39 (O_39,N_14848,N_14572);
xor UO_40 (O_40,N_14757,N_14342);
and UO_41 (O_41,N_14748,N_14753);
nor UO_42 (O_42,N_14430,N_14261);
or UO_43 (O_43,N_14782,N_14274);
nand UO_44 (O_44,N_14722,N_14786);
or UO_45 (O_45,N_14920,N_14845);
nand UO_46 (O_46,N_14324,N_14859);
nor UO_47 (O_47,N_14930,N_14608);
and UO_48 (O_48,N_14889,N_14691);
nor UO_49 (O_49,N_14490,N_14601);
or UO_50 (O_50,N_14252,N_14644);
and UO_51 (O_51,N_14290,N_14449);
nor UO_52 (O_52,N_14743,N_14376);
nor UO_53 (O_53,N_14568,N_14824);
and UO_54 (O_54,N_14396,N_14577);
xnor UO_55 (O_55,N_14571,N_14999);
and UO_56 (O_56,N_14598,N_14328);
nor UO_57 (O_57,N_14511,N_14818);
nand UO_58 (O_58,N_14481,N_14593);
or UO_59 (O_59,N_14370,N_14984);
xnor UO_60 (O_60,N_14399,N_14907);
and UO_61 (O_61,N_14355,N_14688);
or UO_62 (O_62,N_14305,N_14976);
and UO_63 (O_63,N_14995,N_14708);
and UO_64 (O_64,N_14353,N_14521);
and UO_65 (O_65,N_14506,N_14985);
or UO_66 (O_66,N_14735,N_14312);
or UO_67 (O_67,N_14961,N_14855);
or UO_68 (O_68,N_14322,N_14262);
nand UO_69 (O_69,N_14501,N_14698);
xnor UO_70 (O_70,N_14847,N_14956);
nor UO_71 (O_71,N_14914,N_14651);
xor UO_72 (O_72,N_14613,N_14633);
nand UO_73 (O_73,N_14800,N_14692);
nand UO_74 (O_74,N_14841,N_14380);
nor UO_75 (O_75,N_14895,N_14604);
and UO_76 (O_76,N_14971,N_14675);
and UO_77 (O_77,N_14401,N_14822);
xor UO_78 (O_78,N_14751,N_14948);
and UO_79 (O_79,N_14758,N_14546);
xnor UO_80 (O_80,N_14681,N_14709);
and UO_81 (O_81,N_14939,N_14271);
xnor UO_82 (O_82,N_14517,N_14282);
or UO_83 (O_83,N_14877,N_14890);
xnor UO_84 (O_84,N_14612,N_14417);
and UO_85 (O_85,N_14257,N_14497);
or UO_86 (O_86,N_14853,N_14697);
xor UO_87 (O_87,N_14419,N_14699);
xor UO_88 (O_88,N_14875,N_14918);
or UO_89 (O_89,N_14655,N_14409);
and UO_90 (O_90,N_14515,N_14911);
xor UO_91 (O_91,N_14696,N_14831);
xnor UO_92 (O_92,N_14772,N_14727);
or UO_93 (O_93,N_14879,N_14496);
nand UO_94 (O_94,N_14931,N_14404);
nand UO_95 (O_95,N_14363,N_14784);
nor UO_96 (O_96,N_14292,N_14585);
and UO_97 (O_97,N_14922,N_14545);
xnor UO_98 (O_98,N_14400,N_14336);
nand UO_99 (O_99,N_14638,N_14348);
nand UO_100 (O_100,N_14806,N_14494);
or UO_101 (O_101,N_14884,N_14421);
or UO_102 (O_102,N_14333,N_14277);
nor UO_103 (O_103,N_14789,N_14587);
or UO_104 (O_104,N_14398,N_14713);
and UO_105 (O_105,N_14343,N_14969);
and UO_106 (O_106,N_14405,N_14318);
nor UO_107 (O_107,N_14565,N_14795);
or UO_108 (O_108,N_14817,N_14919);
or UO_109 (O_109,N_14308,N_14293);
and UO_110 (O_110,N_14886,N_14367);
nor UO_111 (O_111,N_14617,N_14634);
nor UO_112 (O_112,N_14742,N_14827);
xnor UO_113 (O_113,N_14926,N_14547);
nand UO_114 (O_114,N_14774,N_14317);
nor UO_115 (O_115,N_14579,N_14474);
nor UO_116 (O_116,N_14512,N_14332);
xnor UO_117 (O_117,N_14739,N_14341);
xnor UO_118 (O_118,N_14330,N_14637);
xnor UO_119 (O_119,N_14858,N_14607);
and UO_120 (O_120,N_14386,N_14670);
nand UO_121 (O_121,N_14731,N_14390);
or UO_122 (O_122,N_14570,N_14986);
or UO_123 (O_123,N_14469,N_14628);
or UO_124 (O_124,N_14331,N_14991);
nor UO_125 (O_125,N_14937,N_14462);
xnor UO_126 (O_126,N_14798,N_14520);
nor UO_127 (O_127,N_14899,N_14927);
or UO_128 (O_128,N_14533,N_14668);
and UO_129 (O_129,N_14754,N_14987);
and UO_130 (O_130,N_14964,N_14428);
or UO_131 (O_131,N_14372,N_14647);
or UO_132 (O_132,N_14470,N_14368);
and UO_133 (O_133,N_14590,N_14750);
or UO_134 (O_134,N_14925,N_14620);
xnor UO_135 (O_135,N_14885,N_14359);
nand UO_136 (O_136,N_14661,N_14869);
xnor UO_137 (O_137,N_14498,N_14900);
or UO_138 (O_138,N_14870,N_14745);
xnor UO_139 (O_139,N_14276,N_14482);
nand UO_140 (O_140,N_14729,N_14821);
or UO_141 (O_141,N_14452,N_14588);
nor UO_142 (O_142,N_14599,N_14600);
and UO_143 (O_143,N_14551,N_14273);
nor UO_144 (O_144,N_14923,N_14780);
xor UO_145 (O_145,N_14720,N_14997);
nor UO_146 (O_146,N_14351,N_14673);
xor UO_147 (O_147,N_14279,N_14662);
or UO_148 (O_148,N_14829,N_14868);
xnor UO_149 (O_149,N_14867,N_14575);
or UO_150 (O_150,N_14435,N_14423);
and UO_151 (O_151,N_14251,N_14724);
or UO_152 (O_152,N_14788,N_14935);
and UO_153 (O_153,N_14801,N_14815);
nand UO_154 (O_154,N_14410,N_14326);
nor UO_155 (O_155,N_14752,N_14365);
or UO_156 (O_156,N_14422,N_14854);
xor UO_157 (O_157,N_14896,N_14744);
or UO_158 (O_158,N_14671,N_14687);
xnor UO_159 (O_159,N_14962,N_14349);
xor UO_160 (O_160,N_14830,N_14310);
nand UO_161 (O_161,N_14463,N_14645);
and UO_162 (O_162,N_14429,N_14377);
nor UO_163 (O_163,N_14759,N_14843);
nand UO_164 (O_164,N_14992,N_14672);
and UO_165 (O_165,N_14340,N_14493);
nor UO_166 (O_166,N_14471,N_14910);
nor UO_167 (O_167,N_14933,N_14819);
and UO_168 (O_168,N_14959,N_14385);
and UO_169 (O_169,N_14678,N_14849);
nor UO_170 (O_170,N_14952,N_14500);
or UO_171 (O_171,N_14611,N_14465);
or UO_172 (O_172,N_14796,N_14479);
or UO_173 (O_173,N_14828,N_14865);
or UO_174 (O_174,N_14610,N_14438);
xnor UO_175 (O_175,N_14912,N_14510);
and UO_176 (O_176,N_14812,N_14432);
nand UO_177 (O_177,N_14287,N_14619);
or UO_178 (O_178,N_14297,N_14977);
or UO_179 (O_179,N_14767,N_14450);
nor UO_180 (O_180,N_14475,N_14576);
nand UO_181 (O_181,N_14876,N_14556);
and UO_182 (O_182,N_14835,N_14458);
and UO_183 (O_183,N_14640,N_14898);
or UO_184 (O_184,N_14264,N_14408);
or UO_185 (O_185,N_14970,N_14397);
or UO_186 (O_186,N_14769,N_14666);
xor UO_187 (O_187,N_14569,N_14958);
or UO_188 (O_188,N_14791,N_14563);
or UO_189 (O_189,N_14646,N_14393);
nor UO_190 (O_190,N_14823,N_14761);
nor UO_191 (O_191,N_14455,N_14597);
or UO_192 (O_192,N_14989,N_14804);
nand UO_193 (O_193,N_14538,N_14609);
xnor UO_194 (O_194,N_14411,N_14477);
nor UO_195 (O_195,N_14591,N_14584);
and UO_196 (O_196,N_14439,N_14625);
nand UO_197 (O_197,N_14354,N_14679);
nor UO_198 (O_198,N_14300,N_14542);
xor UO_199 (O_199,N_14560,N_14809);
or UO_200 (O_200,N_14453,N_14272);
nor UO_201 (O_201,N_14446,N_14808);
or UO_202 (O_202,N_14860,N_14667);
xnor UO_203 (O_203,N_14526,N_14487);
and UO_204 (O_204,N_14658,N_14578);
nor UO_205 (O_205,N_14375,N_14424);
nor UO_206 (O_206,N_14878,N_14712);
and UO_207 (O_207,N_14764,N_14840);
nand UO_208 (O_208,N_14839,N_14659);
or UO_209 (O_209,N_14892,N_14285);
or UO_210 (O_210,N_14657,N_14371);
nor UO_211 (O_211,N_14778,N_14998);
and UO_212 (O_212,N_14361,N_14719);
xor UO_213 (O_213,N_14905,N_14857);
nand UO_214 (O_214,N_14623,N_14383);
and UO_215 (O_215,N_14773,N_14909);
or UO_216 (O_216,N_14650,N_14957);
nor UO_217 (O_217,N_14311,N_14605);
nor UO_218 (O_218,N_14596,N_14763);
nor UO_219 (O_219,N_14842,N_14513);
nor UO_220 (O_220,N_14781,N_14451);
and UO_221 (O_221,N_14880,N_14344);
xnor UO_222 (O_222,N_14785,N_14315);
or UO_223 (O_223,N_14381,N_14615);
and UO_224 (O_224,N_14592,N_14391);
nor UO_225 (O_225,N_14941,N_14669);
or UO_226 (O_226,N_14954,N_14717);
nor UO_227 (O_227,N_14387,N_14725);
or UO_228 (O_228,N_14947,N_14975);
or UO_229 (O_229,N_14581,N_14820);
xor UO_230 (O_230,N_14447,N_14721);
nor UO_231 (O_231,N_14485,N_14732);
nor UO_232 (O_232,N_14856,N_14460);
nand UO_233 (O_233,N_14643,N_14929);
nor UO_234 (O_234,N_14530,N_14988);
or UO_235 (O_235,N_14250,N_14942);
and UO_236 (O_236,N_14586,N_14347);
xor UO_237 (O_237,N_14255,N_14531);
nor UO_238 (O_238,N_14389,N_14799);
or UO_239 (O_239,N_14682,N_14901);
xnor UO_240 (O_240,N_14269,N_14339);
and UO_241 (O_241,N_14356,N_14392);
and UO_242 (O_242,N_14406,N_14522);
xor UO_243 (O_243,N_14337,N_14779);
nor UO_244 (O_244,N_14473,N_14529);
and UO_245 (O_245,N_14524,N_14771);
and UO_246 (O_246,N_14738,N_14874);
nand UO_247 (O_247,N_14427,N_14616);
or UO_248 (O_248,N_14559,N_14756);
xnor UO_249 (O_249,N_14676,N_14583);
nand UO_250 (O_250,N_14648,N_14629);
xor UO_251 (O_251,N_14833,N_14836);
nand UO_252 (O_252,N_14968,N_14951);
and UO_253 (O_253,N_14502,N_14445);
xor UO_254 (O_254,N_14979,N_14810);
nand UO_255 (O_255,N_14913,N_14805);
nor UO_256 (O_256,N_14286,N_14940);
or UO_257 (O_257,N_14694,N_14893);
and UO_258 (O_258,N_14495,N_14295);
or UO_259 (O_259,N_14838,N_14352);
or UO_260 (O_260,N_14505,N_14928);
and UO_261 (O_261,N_14811,N_14755);
xnor UO_262 (O_262,N_14516,N_14701);
nor UO_263 (O_263,N_14695,N_14582);
nor UO_264 (O_264,N_14420,N_14614);
and UO_265 (O_265,N_14350,N_14790);
xor UO_266 (O_266,N_14746,N_14514);
nand UO_267 (O_267,N_14834,N_14630);
xor UO_268 (O_268,N_14921,N_14906);
nor UO_269 (O_269,N_14741,N_14730);
nor UO_270 (O_270,N_14562,N_14544);
nand UO_271 (O_271,N_14656,N_14749);
nor UO_272 (O_272,N_14254,N_14814);
nand UO_273 (O_273,N_14589,N_14768);
and UO_274 (O_274,N_14525,N_14314);
or UO_275 (O_275,N_14523,N_14413);
or UO_276 (O_276,N_14663,N_14734);
or UO_277 (O_277,N_14594,N_14946);
nand UO_278 (O_278,N_14258,N_14407);
xnor UO_279 (O_279,N_14466,N_14321);
xnor UO_280 (O_280,N_14897,N_14573);
nor UO_281 (O_281,N_14456,N_14728);
or UO_282 (O_282,N_14541,N_14327);
or UO_283 (O_283,N_14284,N_14881);
nand UO_284 (O_284,N_14762,N_14710);
xnor UO_285 (O_285,N_14394,N_14540);
nor UO_286 (O_286,N_14373,N_14564);
nand UO_287 (O_287,N_14972,N_14464);
xnor UO_288 (O_288,N_14851,N_14723);
nor UO_289 (O_289,N_14832,N_14973);
or UO_290 (O_290,N_14902,N_14503);
nor UO_291 (O_291,N_14296,N_14558);
xor UO_292 (O_292,N_14635,N_14436);
and UO_293 (O_293,N_14622,N_14379);
or UO_294 (O_294,N_14338,N_14626);
or UO_295 (O_295,N_14684,N_14816);
nor UO_296 (O_296,N_14864,N_14299);
or UO_297 (O_297,N_14281,N_14426);
nor UO_298 (O_298,N_14537,N_14554);
and UO_299 (O_299,N_14685,N_14943);
nor UO_300 (O_300,N_14457,N_14680);
or UO_301 (O_301,N_14309,N_14715);
nor UO_302 (O_302,N_14260,N_14862);
and UO_303 (O_303,N_14395,N_14488);
xor UO_304 (O_304,N_14760,N_14364);
nor UO_305 (O_305,N_14459,N_14256);
and UO_306 (O_306,N_14618,N_14509);
nor UO_307 (O_307,N_14304,N_14334);
xnor UO_308 (O_308,N_14298,N_14561);
nand UO_309 (O_309,N_14303,N_14965);
and UO_310 (O_310,N_14480,N_14378);
or UO_311 (O_311,N_14268,N_14621);
or UO_312 (O_312,N_14448,N_14747);
or UO_313 (O_313,N_14549,N_14861);
xor UO_314 (O_314,N_14949,N_14552);
nand UO_315 (O_315,N_14766,N_14548);
nand UO_316 (O_316,N_14916,N_14508);
xnor UO_317 (O_317,N_14433,N_14707);
nand UO_318 (O_318,N_14476,N_14280);
or UO_319 (O_319,N_14491,N_14270);
nand UO_320 (O_320,N_14580,N_14374);
nand UO_321 (O_321,N_14627,N_14478);
or UO_322 (O_322,N_14631,N_14653);
or UO_323 (O_323,N_14700,N_14283);
xor UO_324 (O_324,N_14974,N_14936);
and UO_325 (O_325,N_14519,N_14950);
nor UO_326 (O_326,N_14775,N_14307);
or UO_327 (O_327,N_14437,N_14904);
nor UO_328 (O_328,N_14733,N_14534);
nand UO_329 (O_329,N_14431,N_14320);
and UO_330 (O_330,N_14718,N_14873);
nand UO_331 (O_331,N_14690,N_14492);
nand UO_332 (O_332,N_14850,N_14846);
xnor UO_333 (O_333,N_14444,N_14716);
nand UO_334 (O_334,N_14489,N_14654);
xor UO_335 (O_335,N_14802,N_14649);
or UO_336 (O_336,N_14403,N_14677);
xor UO_337 (O_337,N_14787,N_14903);
nand UO_338 (O_338,N_14414,N_14813);
nand UO_339 (O_339,N_14360,N_14693);
xnor UO_340 (O_340,N_14388,N_14737);
xnor UO_341 (O_341,N_14641,N_14366);
and UO_342 (O_342,N_14528,N_14484);
nor UO_343 (O_343,N_14704,N_14382);
nor UO_344 (O_344,N_14539,N_14883);
xnor UO_345 (O_345,N_14253,N_14550);
nor UO_346 (O_346,N_14797,N_14852);
nand UO_347 (O_347,N_14955,N_14891);
xor UO_348 (O_348,N_14996,N_14980);
or UO_349 (O_349,N_14826,N_14602);
nand UO_350 (O_350,N_14683,N_14953);
nand UO_351 (O_351,N_14527,N_14863);
nor UO_352 (O_352,N_14924,N_14770);
nand UO_353 (O_353,N_14665,N_14543);
nor UO_354 (O_354,N_14960,N_14313);
or UO_355 (O_355,N_14994,N_14711);
xnor UO_356 (O_356,N_14369,N_14966);
nor UO_357 (O_357,N_14714,N_14461);
nand UO_358 (O_358,N_14632,N_14441);
or UO_359 (O_359,N_14944,N_14982);
nand UO_360 (O_360,N_14302,N_14990);
and UO_361 (O_361,N_14306,N_14915);
nand UO_362 (O_362,N_14652,N_14486);
and UO_363 (O_363,N_14301,N_14887);
xnor UO_364 (O_364,N_14357,N_14872);
and UO_365 (O_365,N_14636,N_14689);
xnor UO_366 (O_366,N_14660,N_14553);
or UO_367 (O_367,N_14316,N_14412);
nand UO_368 (O_368,N_14416,N_14705);
or UO_369 (O_369,N_14603,N_14706);
xnor UO_370 (O_370,N_14468,N_14642);
nor UO_371 (O_371,N_14566,N_14518);
and UO_372 (O_372,N_14624,N_14267);
or UO_373 (O_373,N_14442,N_14981);
and UO_374 (O_374,N_14866,N_14358);
nor UO_375 (O_375,N_14445,N_14891);
xnor UO_376 (O_376,N_14748,N_14400);
and UO_377 (O_377,N_14304,N_14288);
nor UO_378 (O_378,N_14694,N_14668);
or UO_379 (O_379,N_14895,N_14803);
and UO_380 (O_380,N_14768,N_14752);
xnor UO_381 (O_381,N_14489,N_14544);
and UO_382 (O_382,N_14925,N_14720);
and UO_383 (O_383,N_14829,N_14554);
nand UO_384 (O_384,N_14845,N_14281);
nand UO_385 (O_385,N_14581,N_14611);
or UO_386 (O_386,N_14343,N_14279);
or UO_387 (O_387,N_14263,N_14314);
and UO_388 (O_388,N_14956,N_14288);
and UO_389 (O_389,N_14527,N_14377);
nand UO_390 (O_390,N_14799,N_14437);
or UO_391 (O_391,N_14631,N_14326);
xnor UO_392 (O_392,N_14964,N_14672);
or UO_393 (O_393,N_14867,N_14553);
xnor UO_394 (O_394,N_14757,N_14253);
nor UO_395 (O_395,N_14258,N_14857);
and UO_396 (O_396,N_14430,N_14591);
xnor UO_397 (O_397,N_14771,N_14419);
xnor UO_398 (O_398,N_14405,N_14797);
nor UO_399 (O_399,N_14308,N_14418);
and UO_400 (O_400,N_14589,N_14969);
or UO_401 (O_401,N_14429,N_14341);
nand UO_402 (O_402,N_14990,N_14284);
nor UO_403 (O_403,N_14640,N_14263);
or UO_404 (O_404,N_14929,N_14599);
nand UO_405 (O_405,N_14721,N_14307);
or UO_406 (O_406,N_14679,N_14847);
or UO_407 (O_407,N_14344,N_14945);
and UO_408 (O_408,N_14426,N_14340);
or UO_409 (O_409,N_14487,N_14371);
xor UO_410 (O_410,N_14630,N_14365);
and UO_411 (O_411,N_14728,N_14923);
nand UO_412 (O_412,N_14626,N_14625);
or UO_413 (O_413,N_14446,N_14355);
nor UO_414 (O_414,N_14926,N_14997);
xnor UO_415 (O_415,N_14683,N_14743);
or UO_416 (O_416,N_14575,N_14624);
nor UO_417 (O_417,N_14971,N_14324);
or UO_418 (O_418,N_14842,N_14462);
nand UO_419 (O_419,N_14839,N_14644);
nand UO_420 (O_420,N_14726,N_14951);
and UO_421 (O_421,N_14890,N_14843);
and UO_422 (O_422,N_14553,N_14406);
nand UO_423 (O_423,N_14749,N_14937);
nand UO_424 (O_424,N_14688,N_14764);
and UO_425 (O_425,N_14634,N_14321);
and UO_426 (O_426,N_14792,N_14950);
nand UO_427 (O_427,N_14508,N_14519);
or UO_428 (O_428,N_14291,N_14539);
xor UO_429 (O_429,N_14855,N_14959);
nand UO_430 (O_430,N_14256,N_14842);
or UO_431 (O_431,N_14260,N_14596);
or UO_432 (O_432,N_14569,N_14741);
nor UO_433 (O_433,N_14359,N_14745);
nand UO_434 (O_434,N_14600,N_14869);
and UO_435 (O_435,N_14337,N_14303);
xor UO_436 (O_436,N_14429,N_14997);
and UO_437 (O_437,N_14297,N_14712);
nand UO_438 (O_438,N_14465,N_14621);
nor UO_439 (O_439,N_14627,N_14323);
nand UO_440 (O_440,N_14648,N_14945);
nand UO_441 (O_441,N_14526,N_14608);
xor UO_442 (O_442,N_14340,N_14588);
and UO_443 (O_443,N_14363,N_14443);
nor UO_444 (O_444,N_14598,N_14506);
xnor UO_445 (O_445,N_14809,N_14305);
and UO_446 (O_446,N_14324,N_14839);
xnor UO_447 (O_447,N_14544,N_14859);
xor UO_448 (O_448,N_14455,N_14784);
nor UO_449 (O_449,N_14882,N_14770);
nor UO_450 (O_450,N_14580,N_14521);
xor UO_451 (O_451,N_14294,N_14390);
nor UO_452 (O_452,N_14817,N_14718);
or UO_453 (O_453,N_14852,N_14370);
nor UO_454 (O_454,N_14957,N_14893);
xnor UO_455 (O_455,N_14364,N_14914);
and UO_456 (O_456,N_14270,N_14980);
xnor UO_457 (O_457,N_14594,N_14728);
nand UO_458 (O_458,N_14505,N_14504);
xor UO_459 (O_459,N_14582,N_14830);
nor UO_460 (O_460,N_14433,N_14355);
nand UO_461 (O_461,N_14968,N_14375);
nand UO_462 (O_462,N_14448,N_14740);
nor UO_463 (O_463,N_14548,N_14530);
or UO_464 (O_464,N_14897,N_14571);
or UO_465 (O_465,N_14350,N_14383);
or UO_466 (O_466,N_14642,N_14617);
nor UO_467 (O_467,N_14504,N_14709);
or UO_468 (O_468,N_14924,N_14619);
and UO_469 (O_469,N_14771,N_14462);
nor UO_470 (O_470,N_14562,N_14365);
or UO_471 (O_471,N_14927,N_14658);
xor UO_472 (O_472,N_14512,N_14397);
and UO_473 (O_473,N_14446,N_14472);
xor UO_474 (O_474,N_14269,N_14353);
and UO_475 (O_475,N_14632,N_14875);
and UO_476 (O_476,N_14773,N_14696);
or UO_477 (O_477,N_14436,N_14629);
and UO_478 (O_478,N_14543,N_14656);
nor UO_479 (O_479,N_14768,N_14484);
xnor UO_480 (O_480,N_14848,N_14496);
nor UO_481 (O_481,N_14970,N_14740);
or UO_482 (O_482,N_14982,N_14926);
nand UO_483 (O_483,N_14849,N_14870);
nand UO_484 (O_484,N_14895,N_14793);
nor UO_485 (O_485,N_14413,N_14276);
nor UO_486 (O_486,N_14942,N_14359);
nor UO_487 (O_487,N_14683,N_14914);
xnor UO_488 (O_488,N_14884,N_14686);
and UO_489 (O_489,N_14910,N_14634);
or UO_490 (O_490,N_14397,N_14984);
xnor UO_491 (O_491,N_14979,N_14884);
nor UO_492 (O_492,N_14495,N_14353);
nand UO_493 (O_493,N_14367,N_14908);
or UO_494 (O_494,N_14515,N_14459);
nand UO_495 (O_495,N_14586,N_14744);
nand UO_496 (O_496,N_14614,N_14813);
xor UO_497 (O_497,N_14807,N_14967);
and UO_498 (O_498,N_14861,N_14894);
or UO_499 (O_499,N_14991,N_14532);
and UO_500 (O_500,N_14300,N_14724);
nor UO_501 (O_501,N_14310,N_14841);
and UO_502 (O_502,N_14539,N_14688);
xnor UO_503 (O_503,N_14939,N_14502);
xor UO_504 (O_504,N_14846,N_14882);
or UO_505 (O_505,N_14338,N_14892);
nand UO_506 (O_506,N_14813,N_14711);
or UO_507 (O_507,N_14852,N_14387);
nand UO_508 (O_508,N_14687,N_14251);
nor UO_509 (O_509,N_14570,N_14699);
nor UO_510 (O_510,N_14978,N_14623);
and UO_511 (O_511,N_14348,N_14944);
nand UO_512 (O_512,N_14600,N_14936);
and UO_513 (O_513,N_14603,N_14771);
nand UO_514 (O_514,N_14469,N_14880);
or UO_515 (O_515,N_14304,N_14841);
nor UO_516 (O_516,N_14827,N_14544);
nand UO_517 (O_517,N_14582,N_14979);
nand UO_518 (O_518,N_14796,N_14331);
nand UO_519 (O_519,N_14806,N_14985);
and UO_520 (O_520,N_14945,N_14725);
or UO_521 (O_521,N_14611,N_14362);
nand UO_522 (O_522,N_14746,N_14969);
nor UO_523 (O_523,N_14365,N_14403);
nand UO_524 (O_524,N_14632,N_14662);
xnor UO_525 (O_525,N_14595,N_14326);
or UO_526 (O_526,N_14963,N_14664);
and UO_527 (O_527,N_14529,N_14523);
nand UO_528 (O_528,N_14265,N_14390);
and UO_529 (O_529,N_14373,N_14411);
and UO_530 (O_530,N_14992,N_14538);
nor UO_531 (O_531,N_14502,N_14946);
or UO_532 (O_532,N_14800,N_14923);
and UO_533 (O_533,N_14903,N_14943);
nor UO_534 (O_534,N_14550,N_14351);
nand UO_535 (O_535,N_14829,N_14250);
or UO_536 (O_536,N_14620,N_14903);
and UO_537 (O_537,N_14562,N_14414);
nor UO_538 (O_538,N_14470,N_14904);
or UO_539 (O_539,N_14478,N_14544);
or UO_540 (O_540,N_14648,N_14437);
and UO_541 (O_541,N_14929,N_14856);
xor UO_542 (O_542,N_14427,N_14934);
and UO_543 (O_543,N_14859,N_14807);
nor UO_544 (O_544,N_14867,N_14796);
nand UO_545 (O_545,N_14989,N_14599);
nor UO_546 (O_546,N_14680,N_14866);
nor UO_547 (O_547,N_14821,N_14379);
or UO_548 (O_548,N_14336,N_14719);
or UO_549 (O_549,N_14603,N_14898);
and UO_550 (O_550,N_14562,N_14910);
nor UO_551 (O_551,N_14466,N_14819);
nand UO_552 (O_552,N_14657,N_14683);
nand UO_553 (O_553,N_14296,N_14674);
or UO_554 (O_554,N_14833,N_14846);
and UO_555 (O_555,N_14593,N_14649);
or UO_556 (O_556,N_14397,N_14252);
xor UO_557 (O_557,N_14537,N_14722);
nor UO_558 (O_558,N_14651,N_14528);
xnor UO_559 (O_559,N_14413,N_14272);
or UO_560 (O_560,N_14909,N_14296);
nand UO_561 (O_561,N_14680,N_14613);
nor UO_562 (O_562,N_14785,N_14310);
nand UO_563 (O_563,N_14730,N_14596);
or UO_564 (O_564,N_14270,N_14942);
or UO_565 (O_565,N_14354,N_14777);
xnor UO_566 (O_566,N_14636,N_14754);
and UO_567 (O_567,N_14389,N_14878);
or UO_568 (O_568,N_14774,N_14682);
or UO_569 (O_569,N_14670,N_14569);
nor UO_570 (O_570,N_14452,N_14426);
or UO_571 (O_571,N_14956,N_14838);
nor UO_572 (O_572,N_14776,N_14903);
xor UO_573 (O_573,N_14395,N_14674);
nand UO_574 (O_574,N_14542,N_14436);
and UO_575 (O_575,N_14488,N_14591);
or UO_576 (O_576,N_14369,N_14955);
and UO_577 (O_577,N_14560,N_14692);
nor UO_578 (O_578,N_14629,N_14808);
nand UO_579 (O_579,N_14885,N_14694);
nand UO_580 (O_580,N_14913,N_14934);
xor UO_581 (O_581,N_14384,N_14701);
nor UO_582 (O_582,N_14791,N_14923);
nand UO_583 (O_583,N_14810,N_14279);
nand UO_584 (O_584,N_14259,N_14276);
xnor UO_585 (O_585,N_14441,N_14537);
nor UO_586 (O_586,N_14806,N_14566);
xnor UO_587 (O_587,N_14339,N_14401);
xor UO_588 (O_588,N_14589,N_14573);
nor UO_589 (O_589,N_14575,N_14951);
nand UO_590 (O_590,N_14402,N_14978);
nand UO_591 (O_591,N_14901,N_14609);
and UO_592 (O_592,N_14994,N_14745);
nor UO_593 (O_593,N_14950,N_14720);
xnor UO_594 (O_594,N_14935,N_14460);
or UO_595 (O_595,N_14392,N_14294);
nand UO_596 (O_596,N_14396,N_14480);
or UO_597 (O_597,N_14615,N_14940);
nor UO_598 (O_598,N_14563,N_14464);
xnor UO_599 (O_599,N_14421,N_14809);
nand UO_600 (O_600,N_14930,N_14431);
and UO_601 (O_601,N_14504,N_14876);
and UO_602 (O_602,N_14630,N_14499);
xnor UO_603 (O_603,N_14915,N_14336);
nand UO_604 (O_604,N_14781,N_14652);
and UO_605 (O_605,N_14890,N_14786);
or UO_606 (O_606,N_14875,N_14769);
and UO_607 (O_607,N_14935,N_14413);
nor UO_608 (O_608,N_14621,N_14326);
or UO_609 (O_609,N_14639,N_14297);
and UO_610 (O_610,N_14655,N_14674);
nand UO_611 (O_611,N_14782,N_14740);
xor UO_612 (O_612,N_14299,N_14957);
or UO_613 (O_613,N_14439,N_14621);
and UO_614 (O_614,N_14433,N_14888);
and UO_615 (O_615,N_14278,N_14697);
nand UO_616 (O_616,N_14920,N_14496);
nor UO_617 (O_617,N_14934,N_14867);
or UO_618 (O_618,N_14348,N_14643);
nor UO_619 (O_619,N_14890,N_14373);
nand UO_620 (O_620,N_14413,N_14855);
xnor UO_621 (O_621,N_14666,N_14473);
xnor UO_622 (O_622,N_14547,N_14472);
nor UO_623 (O_623,N_14305,N_14844);
and UO_624 (O_624,N_14495,N_14467);
xnor UO_625 (O_625,N_14346,N_14948);
and UO_626 (O_626,N_14278,N_14790);
and UO_627 (O_627,N_14881,N_14521);
or UO_628 (O_628,N_14317,N_14813);
nand UO_629 (O_629,N_14805,N_14322);
nand UO_630 (O_630,N_14921,N_14305);
xnor UO_631 (O_631,N_14718,N_14726);
nor UO_632 (O_632,N_14528,N_14966);
or UO_633 (O_633,N_14351,N_14438);
xnor UO_634 (O_634,N_14785,N_14676);
nor UO_635 (O_635,N_14257,N_14780);
or UO_636 (O_636,N_14483,N_14897);
xnor UO_637 (O_637,N_14592,N_14786);
and UO_638 (O_638,N_14558,N_14560);
and UO_639 (O_639,N_14894,N_14566);
or UO_640 (O_640,N_14366,N_14424);
nor UO_641 (O_641,N_14381,N_14546);
and UO_642 (O_642,N_14681,N_14332);
or UO_643 (O_643,N_14453,N_14531);
and UO_644 (O_644,N_14797,N_14388);
and UO_645 (O_645,N_14517,N_14426);
or UO_646 (O_646,N_14649,N_14850);
nand UO_647 (O_647,N_14297,N_14364);
and UO_648 (O_648,N_14832,N_14944);
or UO_649 (O_649,N_14684,N_14558);
and UO_650 (O_650,N_14562,N_14640);
and UO_651 (O_651,N_14601,N_14917);
and UO_652 (O_652,N_14760,N_14922);
xor UO_653 (O_653,N_14796,N_14748);
xnor UO_654 (O_654,N_14710,N_14445);
xor UO_655 (O_655,N_14480,N_14726);
xor UO_656 (O_656,N_14627,N_14340);
nand UO_657 (O_657,N_14366,N_14460);
nand UO_658 (O_658,N_14731,N_14940);
and UO_659 (O_659,N_14523,N_14601);
and UO_660 (O_660,N_14441,N_14578);
nor UO_661 (O_661,N_14318,N_14447);
xnor UO_662 (O_662,N_14842,N_14764);
nor UO_663 (O_663,N_14423,N_14983);
nand UO_664 (O_664,N_14979,N_14718);
xor UO_665 (O_665,N_14721,N_14986);
nand UO_666 (O_666,N_14383,N_14862);
xor UO_667 (O_667,N_14670,N_14341);
xnor UO_668 (O_668,N_14326,N_14458);
nor UO_669 (O_669,N_14297,N_14531);
and UO_670 (O_670,N_14466,N_14620);
and UO_671 (O_671,N_14280,N_14574);
or UO_672 (O_672,N_14556,N_14776);
nor UO_673 (O_673,N_14986,N_14418);
xnor UO_674 (O_674,N_14910,N_14304);
nor UO_675 (O_675,N_14470,N_14260);
xnor UO_676 (O_676,N_14869,N_14662);
nand UO_677 (O_677,N_14265,N_14276);
nand UO_678 (O_678,N_14300,N_14339);
nor UO_679 (O_679,N_14973,N_14362);
nor UO_680 (O_680,N_14361,N_14763);
and UO_681 (O_681,N_14716,N_14665);
nor UO_682 (O_682,N_14536,N_14485);
xnor UO_683 (O_683,N_14345,N_14657);
and UO_684 (O_684,N_14697,N_14762);
xnor UO_685 (O_685,N_14252,N_14474);
nand UO_686 (O_686,N_14926,N_14531);
or UO_687 (O_687,N_14707,N_14462);
xnor UO_688 (O_688,N_14739,N_14417);
or UO_689 (O_689,N_14611,N_14722);
and UO_690 (O_690,N_14538,N_14314);
nor UO_691 (O_691,N_14394,N_14880);
or UO_692 (O_692,N_14852,N_14956);
or UO_693 (O_693,N_14870,N_14712);
nor UO_694 (O_694,N_14919,N_14522);
nor UO_695 (O_695,N_14309,N_14743);
nand UO_696 (O_696,N_14851,N_14558);
xor UO_697 (O_697,N_14833,N_14572);
xor UO_698 (O_698,N_14291,N_14547);
nor UO_699 (O_699,N_14451,N_14544);
nand UO_700 (O_700,N_14585,N_14582);
and UO_701 (O_701,N_14272,N_14728);
and UO_702 (O_702,N_14422,N_14393);
and UO_703 (O_703,N_14636,N_14711);
nor UO_704 (O_704,N_14485,N_14959);
or UO_705 (O_705,N_14326,N_14332);
and UO_706 (O_706,N_14254,N_14651);
xnor UO_707 (O_707,N_14549,N_14892);
nand UO_708 (O_708,N_14900,N_14266);
and UO_709 (O_709,N_14853,N_14406);
and UO_710 (O_710,N_14771,N_14601);
or UO_711 (O_711,N_14504,N_14945);
nand UO_712 (O_712,N_14809,N_14637);
and UO_713 (O_713,N_14716,N_14451);
xor UO_714 (O_714,N_14366,N_14429);
nor UO_715 (O_715,N_14784,N_14672);
nand UO_716 (O_716,N_14390,N_14564);
xor UO_717 (O_717,N_14754,N_14849);
nor UO_718 (O_718,N_14361,N_14949);
and UO_719 (O_719,N_14803,N_14288);
or UO_720 (O_720,N_14999,N_14322);
nor UO_721 (O_721,N_14587,N_14297);
nand UO_722 (O_722,N_14317,N_14479);
nand UO_723 (O_723,N_14326,N_14420);
xnor UO_724 (O_724,N_14504,N_14359);
and UO_725 (O_725,N_14255,N_14827);
and UO_726 (O_726,N_14593,N_14297);
xnor UO_727 (O_727,N_14263,N_14973);
xor UO_728 (O_728,N_14318,N_14696);
nor UO_729 (O_729,N_14815,N_14662);
or UO_730 (O_730,N_14522,N_14839);
or UO_731 (O_731,N_14948,N_14855);
nand UO_732 (O_732,N_14346,N_14395);
or UO_733 (O_733,N_14954,N_14615);
nand UO_734 (O_734,N_14713,N_14558);
and UO_735 (O_735,N_14929,N_14892);
nor UO_736 (O_736,N_14803,N_14416);
nor UO_737 (O_737,N_14360,N_14653);
nor UO_738 (O_738,N_14548,N_14669);
and UO_739 (O_739,N_14438,N_14825);
and UO_740 (O_740,N_14730,N_14276);
xor UO_741 (O_741,N_14493,N_14419);
xor UO_742 (O_742,N_14469,N_14464);
nor UO_743 (O_743,N_14907,N_14396);
nor UO_744 (O_744,N_14561,N_14694);
xnor UO_745 (O_745,N_14930,N_14878);
xnor UO_746 (O_746,N_14726,N_14856);
nand UO_747 (O_747,N_14960,N_14487);
or UO_748 (O_748,N_14563,N_14543);
nand UO_749 (O_749,N_14398,N_14610);
and UO_750 (O_750,N_14721,N_14863);
nand UO_751 (O_751,N_14351,N_14656);
xor UO_752 (O_752,N_14958,N_14824);
nand UO_753 (O_753,N_14614,N_14401);
and UO_754 (O_754,N_14484,N_14984);
nand UO_755 (O_755,N_14397,N_14837);
xor UO_756 (O_756,N_14572,N_14379);
and UO_757 (O_757,N_14789,N_14871);
xnor UO_758 (O_758,N_14594,N_14857);
and UO_759 (O_759,N_14618,N_14746);
or UO_760 (O_760,N_14360,N_14485);
xor UO_761 (O_761,N_14416,N_14989);
nor UO_762 (O_762,N_14268,N_14577);
or UO_763 (O_763,N_14276,N_14995);
or UO_764 (O_764,N_14645,N_14416);
or UO_765 (O_765,N_14288,N_14579);
nand UO_766 (O_766,N_14883,N_14547);
nor UO_767 (O_767,N_14924,N_14939);
nor UO_768 (O_768,N_14820,N_14605);
and UO_769 (O_769,N_14598,N_14628);
or UO_770 (O_770,N_14567,N_14852);
xnor UO_771 (O_771,N_14301,N_14905);
nor UO_772 (O_772,N_14522,N_14787);
and UO_773 (O_773,N_14800,N_14519);
or UO_774 (O_774,N_14801,N_14322);
and UO_775 (O_775,N_14829,N_14545);
and UO_776 (O_776,N_14877,N_14286);
or UO_777 (O_777,N_14448,N_14601);
xor UO_778 (O_778,N_14796,N_14499);
or UO_779 (O_779,N_14264,N_14917);
or UO_780 (O_780,N_14520,N_14283);
nor UO_781 (O_781,N_14852,N_14722);
nand UO_782 (O_782,N_14781,N_14378);
or UO_783 (O_783,N_14585,N_14813);
and UO_784 (O_784,N_14857,N_14604);
nor UO_785 (O_785,N_14802,N_14869);
xor UO_786 (O_786,N_14692,N_14542);
and UO_787 (O_787,N_14936,N_14910);
or UO_788 (O_788,N_14603,N_14288);
or UO_789 (O_789,N_14336,N_14440);
nand UO_790 (O_790,N_14926,N_14384);
nor UO_791 (O_791,N_14356,N_14941);
nor UO_792 (O_792,N_14598,N_14408);
xnor UO_793 (O_793,N_14424,N_14446);
and UO_794 (O_794,N_14873,N_14952);
nand UO_795 (O_795,N_14395,N_14472);
xor UO_796 (O_796,N_14413,N_14734);
nor UO_797 (O_797,N_14318,N_14284);
nand UO_798 (O_798,N_14586,N_14253);
nand UO_799 (O_799,N_14331,N_14541);
nor UO_800 (O_800,N_14806,N_14745);
xnor UO_801 (O_801,N_14690,N_14871);
nand UO_802 (O_802,N_14492,N_14770);
and UO_803 (O_803,N_14651,N_14812);
xnor UO_804 (O_804,N_14401,N_14718);
nor UO_805 (O_805,N_14588,N_14320);
xnor UO_806 (O_806,N_14892,N_14264);
and UO_807 (O_807,N_14323,N_14264);
and UO_808 (O_808,N_14541,N_14536);
nor UO_809 (O_809,N_14634,N_14498);
or UO_810 (O_810,N_14357,N_14517);
or UO_811 (O_811,N_14601,N_14332);
or UO_812 (O_812,N_14961,N_14633);
and UO_813 (O_813,N_14859,N_14561);
and UO_814 (O_814,N_14737,N_14424);
xnor UO_815 (O_815,N_14336,N_14692);
or UO_816 (O_816,N_14281,N_14617);
xor UO_817 (O_817,N_14595,N_14308);
or UO_818 (O_818,N_14661,N_14806);
or UO_819 (O_819,N_14768,N_14524);
nand UO_820 (O_820,N_14893,N_14914);
or UO_821 (O_821,N_14880,N_14608);
nand UO_822 (O_822,N_14519,N_14497);
nor UO_823 (O_823,N_14390,N_14645);
xor UO_824 (O_824,N_14780,N_14553);
and UO_825 (O_825,N_14284,N_14790);
nand UO_826 (O_826,N_14911,N_14996);
xnor UO_827 (O_827,N_14310,N_14894);
nor UO_828 (O_828,N_14926,N_14263);
nand UO_829 (O_829,N_14640,N_14934);
nand UO_830 (O_830,N_14349,N_14987);
and UO_831 (O_831,N_14445,N_14683);
and UO_832 (O_832,N_14585,N_14872);
or UO_833 (O_833,N_14959,N_14729);
and UO_834 (O_834,N_14475,N_14548);
or UO_835 (O_835,N_14263,N_14401);
or UO_836 (O_836,N_14256,N_14720);
and UO_837 (O_837,N_14313,N_14966);
nor UO_838 (O_838,N_14576,N_14483);
nand UO_839 (O_839,N_14433,N_14942);
and UO_840 (O_840,N_14727,N_14811);
nand UO_841 (O_841,N_14255,N_14965);
or UO_842 (O_842,N_14985,N_14827);
or UO_843 (O_843,N_14261,N_14509);
or UO_844 (O_844,N_14633,N_14978);
and UO_845 (O_845,N_14878,N_14600);
xor UO_846 (O_846,N_14562,N_14781);
nand UO_847 (O_847,N_14716,N_14847);
and UO_848 (O_848,N_14385,N_14553);
xor UO_849 (O_849,N_14815,N_14602);
nor UO_850 (O_850,N_14606,N_14352);
xor UO_851 (O_851,N_14354,N_14914);
xor UO_852 (O_852,N_14831,N_14713);
and UO_853 (O_853,N_14806,N_14367);
xnor UO_854 (O_854,N_14686,N_14397);
and UO_855 (O_855,N_14945,N_14477);
and UO_856 (O_856,N_14403,N_14597);
nand UO_857 (O_857,N_14746,N_14295);
xor UO_858 (O_858,N_14693,N_14400);
nor UO_859 (O_859,N_14294,N_14854);
nor UO_860 (O_860,N_14871,N_14944);
xnor UO_861 (O_861,N_14831,N_14388);
xor UO_862 (O_862,N_14420,N_14446);
xor UO_863 (O_863,N_14315,N_14823);
and UO_864 (O_864,N_14407,N_14751);
or UO_865 (O_865,N_14553,N_14451);
xnor UO_866 (O_866,N_14572,N_14314);
and UO_867 (O_867,N_14322,N_14571);
nor UO_868 (O_868,N_14412,N_14643);
or UO_869 (O_869,N_14555,N_14957);
nor UO_870 (O_870,N_14813,N_14898);
and UO_871 (O_871,N_14923,N_14746);
nand UO_872 (O_872,N_14373,N_14345);
or UO_873 (O_873,N_14636,N_14368);
or UO_874 (O_874,N_14983,N_14638);
and UO_875 (O_875,N_14277,N_14517);
and UO_876 (O_876,N_14356,N_14254);
nor UO_877 (O_877,N_14743,N_14684);
or UO_878 (O_878,N_14717,N_14373);
xnor UO_879 (O_879,N_14335,N_14263);
xnor UO_880 (O_880,N_14517,N_14604);
xnor UO_881 (O_881,N_14431,N_14395);
nand UO_882 (O_882,N_14319,N_14765);
or UO_883 (O_883,N_14609,N_14383);
xor UO_884 (O_884,N_14538,N_14423);
nand UO_885 (O_885,N_14507,N_14793);
nor UO_886 (O_886,N_14615,N_14529);
nor UO_887 (O_887,N_14602,N_14643);
or UO_888 (O_888,N_14591,N_14684);
xor UO_889 (O_889,N_14484,N_14850);
xor UO_890 (O_890,N_14995,N_14662);
and UO_891 (O_891,N_14418,N_14566);
and UO_892 (O_892,N_14728,N_14386);
or UO_893 (O_893,N_14659,N_14874);
and UO_894 (O_894,N_14688,N_14761);
xnor UO_895 (O_895,N_14601,N_14673);
nor UO_896 (O_896,N_14970,N_14328);
or UO_897 (O_897,N_14545,N_14767);
xnor UO_898 (O_898,N_14872,N_14823);
xnor UO_899 (O_899,N_14544,N_14764);
xnor UO_900 (O_900,N_14345,N_14754);
nand UO_901 (O_901,N_14899,N_14981);
nand UO_902 (O_902,N_14658,N_14369);
xnor UO_903 (O_903,N_14984,N_14319);
nor UO_904 (O_904,N_14896,N_14863);
nor UO_905 (O_905,N_14685,N_14859);
nand UO_906 (O_906,N_14982,N_14546);
nand UO_907 (O_907,N_14401,N_14649);
and UO_908 (O_908,N_14583,N_14933);
or UO_909 (O_909,N_14846,N_14765);
nand UO_910 (O_910,N_14880,N_14396);
or UO_911 (O_911,N_14297,N_14522);
and UO_912 (O_912,N_14450,N_14806);
nor UO_913 (O_913,N_14635,N_14778);
xnor UO_914 (O_914,N_14977,N_14725);
nor UO_915 (O_915,N_14857,N_14690);
nor UO_916 (O_916,N_14681,N_14459);
or UO_917 (O_917,N_14254,N_14637);
and UO_918 (O_918,N_14994,N_14473);
nand UO_919 (O_919,N_14922,N_14763);
nand UO_920 (O_920,N_14451,N_14749);
xor UO_921 (O_921,N_14275,N_14545);
or UO_922 (O_922,N_14497,N_14820);
and UO_923 (O_923,N_14467,N_14650);
or UO_924 (O_924,N_14814,N_14376);
or UO_925 (O_925,N_14386,N_14281);
and UO_926 (O_926,N_14989,N_14699);
nand UO_927 (O_927,N_14558,N_14548);
nor UO_928 (O_928,N_14341,N_14890);
or UO_929 (O_929,N_14792,N_14886);
nor UO_930 (O_930,N_14968,N_14319);
and UO_931 (O_931,N_14510,N_14266);
or UO_932 (O_932,N_14540,N_14380);
nand UO_933 (O_933,N_14770,N_14909);
xor UO_934 (O_934,N_14448,N_14741);
nand UO_935 (O_935,N_14523,N_14833);
nor UO_936 (O_936,N_14575,N_14985);
and UO_937 (O_937,N_14955,N_14951);
xnor UO_938 (O_938,N_14475,N_14877);
or UO_939 (O_939,N_14483,N_14590);
and UO_940 (O_940,N_14749,N_14263);
and UO_941 (O_941,N_14847,N_14892);
xnor UO_942 (O_942,N_14935,N_14390);
or UO_943 (O_943,N_14680,N_14829);
nor UO_944 (O_944,N_14794,N_14979);
and UO_945 (O_945,N_14640,N_14386);
and UO_946 (O_946,N_14764,N_14456);
nor UO_947 (O_947,N_14549,N_14632);
nand UO_948 (O_948,N_14585,N_14645);
and UO_949 (O_949,N_14323,N_14477);
and UO_950 (O_950,N_14487,N_14546);
and UO_951 (O_951,N_14443,N_14337);
and UO_952 (O_952,N_14296,N_14833);
nor UO_953 (O_953,N_14701,N_14768);
xor UO_954 (O_954,N_14664,N_14569);
and UO_955 (O_955,N_14485,N_14630);
xor UO_956 (O_956,N_14654,N_14548);
nor UO_957 (O_957,N_14540,N_14880);
nor UO_958 (O_958,N_14277,N_14457);
nor UO_959 (O_959,N_14924,N_14334);
xnor UO_960 (O_960,N_14339,N_14752);
xnor UO_961 (O_961,N_14545,N_14555);
xor UO_962 (O_962,N_14375,N_14624);
nor UO_963 (O_963,N_14269,N_14731);
nand UO_964 (O_964,N_14347,N_14707);
and UO_965 (O_965,N_14877,N_14820);
and UO_966 (O_966,N_14763,N_14856);
and UO_967 (O_967,N_14604,N_14270);
nor UO_968 (O_968,N_14800,N_14375);
or UO_969 (O_969,N_14749,N_14638);
or UO_970 (O_970,N_14442,N_14469);
nand UO_971 (O_971,N_14723,N_14473);
or UO_972 (O_972,N_14748,N_14387);
or UO_973 (O_973,N_14556,N_14948);
nor UO_974 (O_974,N_14336,N_14531);
xor UO_975 (O_975,N_14897,N_14544);
nand UO_976 (O_976,N_14738,N_14380);
xnor UO_977 (O_977,N_14509,N_14402);
and UO_978 (O_978,N_14684,N_14616);
or UO_979 (O_979,N_14702,N_14283);
and UO_980 (O_980,N_14553,N_14617);
nor UO_981 (O_981,N_14789,N_14323);
nor UO_982 (O_982,N_14563,N_14986);
nand UO_983 (O_983,N_14404,N_14760);
nor UO_984 (O_984,N_14903,N_14289);
nand UO_985 (O_985,N_14492,N_14484);
and UO_986 (O_986,N_14879,N_14416);
nor UO_987 (O_987,N_14844,N_14385);
and UO_988 (O_988,N_14504,N_14385);
or UO_989 (O_989,N_14594,N_14546);
and UO_990 (O_990,N_14759,N_14391);
or UO_991 (O_991,N_14288,N_14654);
and UO_992 (O_992,N_14728,N_14776);
nand UO_993 (O_993,N_14491,N_14350);
or UO_994 (O_994,N_14411,N_14338);
or UO_995 (O_995,N_14705,N_14687);
or UO_996 (O_996,N_14717,N_14822);
or UO_997 (O_997,N_14931,N_14952);
nand UO_998 (O_998,N_14610,N_14903);
nor UO_999 (O_999,N_14632,N_14386);
xor UO_1000 (O_1000,N_14879,N_14726);
nand UO_1001 (O_1001,N_14509,N_14556);
xor UO_1002 (O_1002,N_14333,N_14527);
xor UO_1003 (O_1003,N_14929,N_14781);
nor UO_1004 (O_1004,N_14480,N_14283);
or UO_1005 (O_1005,N_14671,N_14442);
nor UO_1006 (O_1006,N_14673,N_14332);
and UO_1007 (O_1007,N_14783,N_14802);
nor UO_1008 (O_1008,N_14735,N_14473);
nand UO_1009 (O_1009,N_14662,N_14837);
or UO_1010 (O_1010,N_14292,N_14544);
xor UO_1011 (O_1011,N_14279,N_14733);
xor UO_1012 (O_1012,N_14406,N_14684);
nand UO_1013 (O_1013,N_14820,N_14705);
xnor UO_1014 (O_1014,N_14842,N_14929);
nor UO_1015 (O_1015,N_14780,N_14395);
or UO_1016 (O_1016,N_14522,N_14632);
nand UO_1017 (O_1017,N_14859,N_14757);
nand UO_1018 (O_1018,N_14577,N_14366);
nor UO_1019 (O_1019,N_14456,N_14495);
nor UO_1020 (O_1020,N_14586,N_14525);
and UO_1021 (O_1021,N_14981,N_14465);
or UO_1022 (O_1022,N_14587,N_14752);
or UO_1023 (O_1023,N_14486,N_14338);
nor UO_1024 (O_1024,N_14324,N_14379);
nand UO_1025 (O_1025,N_14576,N_14552);
and UO_1026 (O_1026,N_14666,N_14890);
nor UO_1027 (O_1027,N_14295,N_14914);
nor UO_1028 (O_1028,N_14883,N_14299);
and UO_1029 (O_1029,N_14906,N_14372);
or UO_1030 (O_1030,N_14686,N_14419);
nand UO_1031 (O_1031,N_14858,N_14647);
xnor UO_1032 (O_1032,N_14480,N_14660);
nor UO_1033 (O_1033,N_14689,N_14629);
and UO_1034 (O_1034,N_14667,N_14816);
xnor UO_1035 (O_1035,N_14668,N_14531);
nor UO_1036 (O_1036,N_14363,N_14886);
xor UO_1037 (O_1037,N_14580,N_14995);
nor UO_1038 (O_1038,N_14927,N_14827);
or UO_1039 (O_1039,N_14715,N_14450);
nand UO_1040 (O_1040,N_14276,N_14549);
and UO_1041 (O_1041,N_14481,N_14426);
xor UO_1042 (O_1042,N_14674,N_14905);
nor UO_1043 (O_1043,N_14737,N_14621);
xnor UO_1044 (O_1044,N_14905,N_14445);
nand UO_1045 (O_1045,N_14521,N_14424);
nor UO_1046 (O_1046,N_14909,N_14698);
and UO_1047 (O_1047,N_14758,N_14631);
or UO_1048 (O_1048,N_14982,N_14580);
xnor UO_1049 (O_1049,N_14252,N_14499);
nor UO_1050 (O_1050,N_14321,N_14614);
nor UO_1051 (O_1051,N_14561,N_14660);
nand UO_1052 (O_1052,N_14795,N_14836);
nand UO_1053 (O_1053,N_14791,N_14981);
nand UO_1054 (O_1054,N_14986,N_14580);
xnor UO_1055 (O_1055,N_14803,N_14388);
nand UO_1056 (O_1056,N_14578,N_14830);
nor UO_1057 (O_1057,N_14589,N_14550);
and UO_1058 (O_1058,N_14389,N_14782);
nand UO_1059 (O_1059,N_14397,N_14874);
nand UO_1060 (O_1060,N_14929,N_14875);
nor UO_1061 (O_1061,N_14758,N_14912);
or UO_1062 (O_1062,N_14652,N_14602);
nand UO_1063 (O_1063,N_14377,N_14894);
or UO_1064 (O_1064,N_14843,N_14760);
xor UO_1065 (O_1065,N_14298,N_14721);
and UO_1066 (O_1066,N_14559,N_14421);
and UO_1067 (O_1067,N_14816,N_14694);
or UO_1068 (O_1068,N_14829,N_14439);
and UO_1069 (O_1069,N_14349,N_14449);
xor UO_1070 (O_1070,N_14345,N_14261);
nand UO_1071 (O_1071,N_14531,N_14541);
nand UO_1072 (O_1072,N_14711,N_14316);
or UO_1073 (O_1073,N_14804,N_14595);
or UO_1074 (O_1074,N_14954,N_14996);
and UO_1075 (O_1075,N_14606,N_14431);
or UO_1076 (O_1076,N_14538,N_14605);
nor UO_1077 (O_1077,N_14733,N_14516);
and UO_1078 (O_1078,N_14311,N_14808);
nand UO_1079 (O_1079,N_14686,N_14687);
nand UO_1080 (O_1080,N_14644,N_14409);
or UO_1081 (O_1081,N_14415,N_14571);
xnor UO_1082 (O_1082,N_14797,N_14952);
and UO_1083 (O_1083,N_14898,N_14573);
nand UO_1084 (O_1084,N_14991,N_14721);
nor UO_1085 (O_1085,N_14402,N_14653);
xnor UO_1086 (O_1086,N_14799,N_14788);
or UO_1087 (O_1087,N_14737,N_14734);
xnor UO_1088 (O_1088,N_14355,N_14826);
xor UO_1089 (O_1089,N_14272,N_14968);
nand UO_1090 (O_1090,N_14828,N_14257);
and UO_1091 (O_1091,N_14693,N_14891);
nor UO_1092 (O_1092,N_14423,N_14613);
nand UO_1093 (O_1093,N_14653,N_14664);
nand UO_1094 (O_1094,N_14560,N_14264);
nand UO_1095 (O_1095,N_14345,N_14948);
and UO_1096 (O_1096,N_14885,N_14417);
nor UO_1097 (O_1097,N_14869,N_14885);
or UO_1098 (O_1098,N_14842,N_14960);
and UO_1099 (O_1099,N_14485,N_14842);
and UO_1100 (O_1100,N_14620,N_14915);
or UO_1101 (O_1101,N_14363,N_14931);
xnor UO_1102 (O_1102,N_14594,N_14344);
nor UO_1103 (O_1103,N_14502,N_14780);
nand UO_1104 (O_1104,N_14668,N_14355);
or UO_1105 (O_1105,N_14652,N_14439);
nand UO_1106 (O_1106,N_14448,N_14940);
nor UO_1107 (O_1107,N_14366,N_14979);
nand UO_1108 (O_1108,N_14752,N_14947);
xnor UO_1109 (O_1109,N_14271,N_14880);
xnor UO_1110 (O_1110,N_14698,N_14771);
xnor UO_1111 (O_1111,N_14360,N_14799);
and UO_1112 (O_1112,N_14265,N_14515);
nor UO_1113 (O_1113,N_14483,N_14585);
nor UO_1114 (O_1114,N_14924,N_14911);
or UO_1115 (O_1115,N_14479,N_14871);
nand UO_1116 (O_1116,N_14540,N_14624);
nor UO_1117 (O_1117,N_14984,N_14972);
or UO_1118 (O_1118,N_14528,N_14797);
xnor UO_1119 (O_1119,N_14974,N_14381);
nor UO_1120 (O_1120,N_14830,N_14382);
nor UO_1121 (O_1121,N_14280,N_14460);
and UO_1122 (O_1122,N_14809,N_14610);
or UO_1123 (O_1123,N_14729,N_14560);
nand UO_1124 (O_1124,N_14960,N_14676);
xor UO_1125 (O_1125,N_14637,N_14669);
xnor UO_1126 (O_1126,N_14889,N_14698);
and UO_1127 (O_1127,N_14658,N_14430);
or UO_1128 (O_1128,N_14628,N_14525);
nand UO_1129 (O_1129,N_14566,N_14395);
and UO_1130 (O_1130,N_14395,N_14609);
nor UO_1131 (O_1131,N_14349,N_14973);
and UO_1132 (O_1132,N_14717,N_14515);
nand UO_1133 (O_1133,N_14655,N_14620);
xnor UO_1134 (O_1134,N_14923,N_14299);
or UO_1135 (O_1135,N_14911,N_14966);
and UO_1136 (O_1136,N_14783,N_14378);
or UO_1137 (O_1137,N_14679,N_14439);
xor UO_1138 (O_1138,N_14949,N_14699);
and UO_1139 (O_1139,N_14790,N_14834);
or UO_1140 (O_1140,N_14400,N_14785);
and UO_1141 (O_1141,N_14927,N_14879);
nor UO_1142 (O_1142,N_14716,N_14898);
xor UO_1143 (O_1143,N_14464,N_14788);
or UO_1144 (O_1144,N_14845,N_14927);
and UO_1145 (O_1145,N_14560,N_14542);
xor UO_1146 (O_1146,N_14777,N_14866);
and UO_1147 (O_1147,N_14800,N_14644);
and UO_1148 (O_1148,N_14869,N_14924);
and UO_1149 (O_1149,N_14969,N_14712);
or UO_1150 (O_1150,N_14571,N_14299);
nor UO_1151 (O_1151,N_14771,N_14797);
and UO_1152 (O_1152,N_14556,N_14814);
nand UO_1153 (O_1153,N_14281,N_14436);
nor UO_1154 (O_1154,N_14728,N_14447);
and UO_1155 (O_1155,N_14295,N_14543);
nand UO_1156 (O_1156,N_14638,N_14414);
nor UO_1157 (O_1157,N_14251,N_14899);
nand UO_1158 (O_1158,N_14628,N_14863);
nor UO_1159 (O_1159,N_14405,N_14430);
xor UO_1160 (O_1160,N_14759,N_14624);
or UO_1161 (O_1161,N_14724,N_14310);
nor UO_1162 (O_1162,N_14884,N_14493);
xnor UO_1163 (O_1163,N_14611,N_14700);
nor UO_1164 (O_1164,N_14968,N_14556);
nand UO_1165 (O_1165,N_14793,N_14526);
and UO_1166 (O_1166,N_14523,N_14291);
or UO_1167 (O_1167,N_14930,N_14985);
and UO_1168 (O_1168,N_14834,N_14866);
nand UO_1169 (O_1169,N_14792,N_14472);
nor UO_1170 (O_1170,N_14734,N_14931);
nand UO_1171 (O_1171,N_14308,N_14618);
and UO_1172 (O_1172,N_14773,N_14266);
nand UO_1173 (O_1173,N_14429,N_14363);
and UO_1174 (O_1174,N_14311,N_14801);
xnor UO_1175 (O_1175,N_14528,N_14821);
nand UO_1176 (O_1176,N_14489,N_14355);
xnor UO_1177 (O_1177,N_14618,N_14530);
nor UO_1178 (O_1178,N_14551,N_14770);
and UO_1179 (O_1179,N_14939,N_14552);
and UO_1180 (O_1180,N_14361,N_14776);
and UO_1181 (O_1181,N_14520,N_14289);
nor UO_1182 (O_1182,N_14475,N_14462);
nand UO_1183 (O_1183,N_14323,N_14968);
nor UO_1184 (O_1184,N_14438,N_14289);
nor UO_1185 (O_1185,N_14993,N_14977);
xor UO_1186 (O_1186,N_14603,N_14258);
or UO_1187 (O_1187,N_14694,N_14834);
nor UO_1188 (O_1188,N_14313,N_14543);
nand UO_1189 (O_1189,N_14337,N_14713);
nor UO_1190 (O_1190,N_14964,N_14915);
xnor UO_1191 (O_1191,N_14708,N_14335);
nand UO_1192 (O_1192,N_14750,N_14723);
nand UO_1193 (O_1193,N_14352,N_14633);
nand UO_1194 (O_1194,N_14946,N_14314);
nand UO_1195 (O_1195,N_14476,N_14947);
nand UO_1196 (O_1196,N_14292,N_14576);
nand UO_1197 (O_1197,N_14987,N_14566);
and UO_1198 (O_1198,N_14822,N_14734);
or UO_1199 (O_1199,N_14773,N_14677);
or UO_1200 (O_1200,N_14395,N_14869);
or UO_1201 (O_1201,N_14404,N_14674);
nand UO_1202 (O_1202,N_14377,N_14974);
and UO_1203 (O_1203,N_14320,N_14371);
xor UO_1204 (O_1204,N_14910,N_14484);
nor UO_1205 (O_1205,N_14401,N_14816);
nand UO_1206 (O_1206,N_14645,N_14743);
or UO_1207 (O_1207,N_14569,N_14696);
or UO_1208 (O_1208,N_14269,N_14489);
nor UO_1209 (O_1209,N_14634,N_14743);
nor UO_1210 (O_1210,N_14797,N_14815);
nor UO_1211 (O_1211,N_14718,N_14877);
nand UO_1212 (O_1212,N_14821,N_14925);
nor UO_1213 (O_1213,N_14373,N_14837);
xor UO_1214 (O_1214,N_14793,N_14429);
or UO_1215 (O_1215,N_14877,N_14369);
nand UO_1216 (O_1216,N_14613,N_14281);
or UO_1217 (O_1217,N_14845,N_14672);
nand UO_1218 (O_1218,N_14992,N_14323);
nor UO_1219 (O_1219,N_14925,N_14536);
and UO_1220 (O_1220,N_14919,N_14643);
nor UO_1221 (O_1221,N_14995,N_14919);
or UO_1222 (O_1222,N_14497,N_14926);
xor UO_1223 (O_1223,N_14905,N_14842);
and UO_1224 (O_1224,N_14480,N_14918);
nor UO_1225 (O_1225,N_14404,N_14483);
and UO_1226 (O_1226,N_14868,N_14271);
xor UO_1227 (O_1227,N_14873,N_14732);
nor UO_1228 (O_1228,N_14997,N_14290);
xnor UO_1229 (O_1229,N_14931,N_14523);
and UO_1230 (O_1230,N_14403,N_14372);
xor UO_1231 (O_1231,N_14375,N_14720);
nor UO_1232 (O_1232,N_14920,N_14319);
and UO_1233 (O_1233,N_14675,N_14947);
or UO_1234 (O_1234,N_14383,N_14627);
nand UO_1235 (O_1235,N_14541,N_14254);
and UO_1236 (O_1236,N_14834,N_14728);
or UO_1237 (O_1237,N_14724,N_14462);
xnor UO_1238 (O_1238,N_14533,N_14474);
and UO_1239 (O_1239,N_14782,N_14745);
and UO_1240 (O_1240,N_14371,N_14592);
nor UO_1241 (O_1241,N_14799,N_14971);
or UO_1242 (O_1242,N_14306,N_14526);
and UO_1243 (O_1243,N_14534,N_14809);
nor UO_1244 (O_1244,N_14253,N_14589);
and UO_1245 (O_1245,N_14692,N_14665);
or UO_1246 (O_1246,N_14345,N_14442);
xor UO_1247 (O_1247,N_14615,N_14814);
or UO_1248 (O_1248,N_14933,N_14648);
xnor UO_1249 (O_1249,N_14909,N_14798);
nand UO_1250 (O_1250,N_14548,N_14353);
and UO_1251 (O_1251,N_14383,N_14800);
nand UO_1252 (O_1252,N_14600,N_14852);
nand UO_1253 (O_1253,N_14458,N_14537);
nor UO_1254 (O_1254,N_14693,N_14885);
and UO_1255 (O_1255,N_14392,N_14907);
and UO_1256 (O_1256,N_14547,N_14899);
or UO_1257 (O_1257,N_14432,N_14940);
xor UO_1258 (O_1258,N_14970,N_14402);
nor UO_1259 (O_1259,N_14367,N_14407);
xnor UO_1260 (O_1260,N_14733,N_14592);
nor UO_1261 (O_1261,N_14495,N_14799);
xnor UO_1262 (O_1262,N_14702,N_14291);
nor UO_1263 (O_1263,N_14883,N_14718);
nand UO_1264 (O_1264,N_14265,N_14744);
or UO_1265 (O_1265,N_14495,N_14641);
xor UO_1266 (O_1266,N_14647,N_14946);
nor UO_1267 (O_1267,N_14685,N_14281);
or UO_1268 (O_1268,N_14423,N_14804);
nand UO_1269 (O_1269,N_14403,N_14778);
nor UO_1270 (O_1270,N_14547,N_14293);
nand UO_1271 (O_1271,N_14962,N_14790);
and UO_1272 (O_1272,N_14417,N_14817);
nor UO_1273 (O_1273,N_14472,N_14450);
nand UO_1274 (O_1274,N_14675,N_14328);
and UO_1275 (O_1275,N_14985,N_14330);
xnor UO_1276 (O_1276,N_14575,N_14291);
or UO_1277 (O_1277,N_14549,N_14721);
and UO_1278 (O_1278,N_14509,N_14457);
nand UO_1279 (O_1279,N_14517,N_14893);
xnor UO_1280 (O_1280,N_14982,N_14545);
xor UO_1281 (O_1281,N_14792,N_14880);
xor UO_1282 (O_1282,N_14883,N_14861);
or UO_1283 (O_1283,N_14315,N_14867);
nor UO_1284 (O_1284,N_14370,N_14818);
and UO_1285 (O_1285,N_14715,N_14308);
xor UO_1286 (O_1286,N_14856,N_14935);
nor UO_1287 (O_1287,N_14790,N_14685);
nor UO_1288 (O_1288,N_14966,N_14296);
nor UO_1289 (O_1289,N_14268,N_14790);
xor UO_1290 (O_1290,N_14749,N_14273);
or UO_1291 (O_1291,N_14613,N_14951);
xor UO_1292 (O_1292,N_14766,N_14997);
nor UO_1293 (O_1293,N_14422,N_14721);
xnor UO_1294 (O_1294,N_14789,N_14711);
and UO_1295 (O_1295,N_14853,N_14625);
and UO_1296 (O_1296,N_14922,N_14859);
and UO_1297 (O_1297,N_14496,N_14820);
and UO_1298 (O_1298,N_14893,N_14824);
nor UO_1299 (O_1299,N_14540,N_14289);
or UO_1300 (O_1300,N_14350,N_14252);
nor UO_1301 (O_1301,N_14334,N_14664);
nand UO_1302 (O_1302,N_14683,N_14624);
xnor UO_1303 (O_1303,N_14251,N_14471);
or UO_1304 (O_1304,N_14575,N_14818);
and UO_1305 (O_1305,N_14727,N_14649);
or UO_1306 (O_1306,N_14710,N_14373);
nand UO_1307 (O_1307,N_14920,N_14262);
xor UO_1308 (O_1308,N_14888,N_14585);
and UO_1309 (O_1309,N_14905,N_14817);
nand UO_1310 (O_1310,N_14263,N_14612);
or UO_1311 (O_1311,N_14256,N_14493);
nand UO_1312 (O_1312,N_14923,N_14572);
and UO_1313 (O_1313,N_14331,N_14554);
and UO_1314 (O_1314,N_14665,N_14731);
nor UO_1315 (O_1315,N_14554,N_14555);
xnor UO_1316 (O_1316,N_14709,N_14291);
nor UO_1317 (O_1317,N_14652,N_14570);
or UO_1318 (O_1318,N_14964,N_14620);
nor UO_1319 (O_1319,N_14895,N_14324);
and UO_1320 (O_1320,N_14316,N_14319);
and UO_1321 (O_1321,N_14286,N_14437);
xnor UO_1322 (O_1322,N_14902,N_14415);
xor UO_1323 (O_1323,N_14967,N_14447);
or UO_1324 (O_1324,N_14829,N_14488);
nor UO_1325 (O_1325,N_14464,N_14967);
and UO_1326 (O_1326,N_14638,N_14402);
and UO_1327 (O_1327,N_14833,N_14321);
nand UO_1328 (O_1328,N_14748,N_14778);
and UO_1329 (O_1329,N_14669,N_14590);
and UO_1330 (O_1330,N_14353,N_14550);
nand UO_1331 (O_1331,N_14821,N_14676);
nand UO_1332 (O_1332,N_14949,N_14612);
or UO_1333 (O_1333,N_14435,N_14522);
nand UO_1334 (O_1334,N_14432,N_14795);
xnor UO_1335 (O_1335,N_14619,N_14330);
or UO_1336 (O_1336,N_14800,N_14468);
nor UO_1337 (O_1337,N_14312,N_14273);
nand UO_1338 (O_1338,N_14295,N_14843);
and UO_1339 (O_1339,N_14471,N_14920);
and UO_1340 (O_1340,N_14817,N_14684);
nor UO_1341 (O_1341,N_14528,N_14426);
nand UO_1342 (O_1342,N_14645,N_14386);
and UO_1343 (O_1343,N_14259,N_14538);
and UO_1344 (O_1344,N_14278,N_14736);
or UO_1345 (O_1345,N_14390,N_14744);
nand UO_1346 (O_1346,N_14731,N_14280);
nand UO_1347 (O_1347,N_14627,N_14687);
xor UO_1348 (O_1348,N_14398,N_14933);
or UO_1349 (O_1349,N_14745,N_14748);
nor UO_1350 (O_1350,N_14590,N_14822);
xor UO_1351 (O_1351,N_14868,N_14537);
nand UO_1352 (O_1352,N_14778,N_14543);
xor UO_1353 (O_1353,N_14353,N_14632);
or UO_1354 (O_1354,N_14415,N_14290);
xor UO_1355 (O_1355,N_14669,N_14638);
and UO_1356 (O_1356,N_14344,N_14853);
xor UO_1357 (O_1357,N_14646,N_14361);
nand UO_1358 (O_1358,N_14483,N_14586);
nor UO_1359 (O_1359,N_14490,N_14607);
and UO_1360 (O_1360,N_14547,N_14972);
nor UO_1361 (O_1361,N_14398,N_14515);
and UO_1362 (O_1362,N_14575,N_14678);
or UO_1363 (O_1363,N_14841,N_14405);
xor UO_1364 (O_1364,N_14578,N_14488);
xnor UO_1365 (O_1365,N_14924,N_14793);
or UO_1366 (O_1366,N_14781,N_14695);
nor UO_1367 (O_1367,N_14825,N_14943);
nand UO_1368 (O_1368,N_14727,N_14965);
or UO_1369 (O_1369,N_14494,N_14644);
and UO_1370 (O_1370,N_14870,N_14924);
or UO_1371 (O_1371,N_14575,N_14660);
xnor UO_1372 (O_1372,N_14259,N_14939);
nand UO_1373 (O_1373,N_14353,N_14591);
xnor UO_1374 (O_1374,N_14331,N_14556);
nor UO_1375 (O_1375,N_14437,N_14941);
xor UO_1376 (O_1376,N_14444,N_14250);
xor UO_1377 (O_1377,N_14368,N_14538);
nor UO_1378 (O_1378,N_14791,N_14826);
nand UO_1379 (O_1379,N_14835,N_14417);
nand UO_1380 (O_1380,N_14500,N_14621);
nor UO_1381 (O_1381,N_14630,N_14492);
or UO_1382 (O_1382,N_14960,N_14852);
nor UO_1383 (O_1383,N_14804,N_14646);
nand UO_1384 (O_1384,N_14601,N_14745);
or UO_1385 (O_1385,N_14669,N_14811);
and UO_1386 (O_1386,N_14427,N_14295);
nand UO_1387 (O_1387,N_14367,N_14737);
nor UO_1388 (O_1388,N_14272,N_14493);
nand UO_1389 (O_1389,N_14471,N_14345);
and UO_1390 (O_1390,N_14440,N_14983);
and UO_1391 (O_1391,N_14734,N_14920);
nand UO_1392 (O_1392,N_14759,N_14293);
and UO_1393 (O_1393,N_14750,N_14250);
or UO_1394 (O_1394,N_14473,N_14914);
or UO_1395 (O_1395,N_14995,N_14689);
xnor UO_1396 (O_1396,N_14272,N_14823);
or UO_1397 (O_1397,N_14659,N_14970);
xnor UO_1398 (O_1398,N_14953,N_14401);
xor UO_1399 (O_1399,N_14527,N_14961);
nor UO_1400 (O_1400,N_14633,N_14813);
or UO_1401 (O_1401,N_14469,N_14334);
and UO_1402 (O_1402,N_14403,N_14396);
or UO_1403 (O_1403,N_14844,N_14643);
xor UO_1404 (O_1404,N_14994,N_14993);
xnor UO_1405 (O_1405,N_14488,N_14749);
nor UO_1406 (O_1406,N_14387,N_14851);
xnor UO_1407 (O_1407,N_14987,N_14340);
nor UO_1408 (O_1408,N_14380,N_14726);
and UO_1409 (O_1409,N_14325,N_14826);
or UO_1410 (O_1410,N_14574,N_14559);
nor UO_1411 (O_1411,N_14458,N_14628);
xnor UO_1412 (O_1412,N_14553,N_14651);
nand UO_1413 (O_1413,N_14334,N_14817);
nand UO_1414 (O_1414,N_14364,N_14528);
or UO_1415 (O_1415,N_14873,N_14562);
and UO_1416 (O_1416,N_14981,N_14809);
and UO_1417 (O_1417,N_14704,N_14482);
nor UO_1418 (O_1418,N_14679,N_14516);
nand UO_1419 (O_1419,N_14635,N_14333);
nor UO_1420 (O_1420,N_14837,N_14769);
nor UO_1421 (O_1421,N_14754,N_14392);
nor UO_1422 (O_1422,N_14290,N_14984);
nand UO_1423 (O_1423,N_14285,N_14635);
nand UO_1424 (O_1424,N_14887,N_14401);
nor UO_1425 (O_1425,N_14489,N_14469);
or UO_1426 (O_1426,N_14254,N_14464);
or UO_1427 (O_1427,N_14691,N_14999);
or UO_1428 (O_1428,N_14761,N_14270);
or UO_1429 (O_1429,N_14293,N_14898);
nand UO_1430 (O_1430,N_14269,N_14263);
or UO_1431 (O_1431,N_14485,N_14602);
xnor UO_1432 (O_1432,N_14295,N_14705);
xnor UO_1433 (O_1433,N_14602,N_14513);
or UO_1434 (O_1434,N_14883,N_14631);
xor UO_1435 (O_1435,N_14673,N_14471);
xnor UO_1436 (O_1436,N_14517,N_14256);
and UO_1437 (O_1437,N_14374,N_14645);
and UO_1438 (O_1438,N_14932,N_14591);
and UO_1439 (O_1439,N_14974,N_14872);
nand UO_1440 (O_1440,N_14949,N_14429);
xnor UO_1441 (O_1441,N_14867,N_14509);
nand UO_1442 (O_1442,N_14325,N_14448);
nand UO_1443 (O_1443,N_14629,N_14613);
nand UO_1444 (O_1444,N_14782,N_14775);
xor UO_1445 (O_1445,N_14714,N_14999);
or UO_1446 (O_1446,N_14676,N_14432);
xor UO_1447 (O_1447,N_14608,N_14902);
xor UO_1448 (O_1448,N_14756,N_14370);
nor UO_1449 (O_1449,N_14775,N_14886);
nand UO_1450 (O_1450,N_14389,N_14430);
nand UO_1451 (O_1451,N_14827,N_14298);
nand UO_1452 (O_1452,N_14255,N_14503);
xor UO_1453 (O_1453,N_14378,N_14758);
nand UO_1454 (O_1454,N_14814,N_14731);
and UO_1455 (O_1455,N_14486,N_14318);
nor UO_1456 (O_1456,N_14984,N_14523);
nor UO_1457 (O_1457,N_14348,N_14349);
or UO_1458 (O_1458,N_14567,N_14448);
nand UO_1459 (O_1459,N_14631,N_14643);
or UO_1460 (O_1460,N_14803,N_14521);
or UO_1461 (O_1461,N_14835,N_14890);
or UO_1462 (O_1462,N_14682,N_14658);
and UO_1463 (O_1463,N_14958,N_14675);
and UO_1464 (O_1464,N_14827,N_14988);
and UO_1465 (O_1465,N_14794,N_14887);
nand UO_1466 (O_1466,N_14994,N_14685);
xnor UO_1467 (O_1467,N_14800,N_14447);
and UO_1468 (O_1468,N_14486,N_14869);
nand UO_1469 (O_1469,N_14414,N_14496);
and UO_1470 (O_1470,N_14851,N_14907);
nand UO_1471 (O_1471,N_14536,N_14821);
or UO_1472 (O_1472,N_14379,N_14750);
xor UO_1473 (O_1473,N_14271,N_14263);
and UO_1474 (O_1474,N_14850,N_14349);
and UO_1475 (O_1475,N_14387,N_14577);
or UO_1476 (O_1476,N_14500,N_14526);
xnor UO_1477 (O_1477,N_14288,N_14897);
nand UO_1478 (O_1478,N_14944,N_14335);
nor UO_1479 (O_1479,N_14410,N_14605);
xor UO_1480 (O_1480,N_14307,N_14825);
nor UO_1481 (O_1481,N_14891,N_14388);
nand UO_1482 (O_1482,N_14827,N_14731);
nand UO_1483 (O_1483,N_14855,N_14774);
and UO_1484 (O_1484,N_14745,N_14426);
xor UO_1485 (O_1485,N_14822,N_14992);
nand UO_1486 (O_1486,N_14275,N_14952);
nor UO_1487 (O_1487,N_14726,N_14557);
nand UO_1488 (O_1488,N_14822,N_14995);
nor UO_1489 (O_1489,N_14997,N_14932);
and UO_1490 (O_1490,N_14782,N_14560);
nor UO_1491 (O_1491,N_14977,N_14443);
or UO_1492 (O_1492,N_14796,N_14305);
and UO_1493 (O_1493,N_14397,N_14610);
and UO_1494 (O_1494,N_14289,N_14891);
xor UO_1495 (O_1495,N_14893,N_14412);
nand UO_1496 (O_1496,N_14616,N_14510);
or UO_1497 (O_1497,N_14462,N_14898);
or UO_1498 (O_1498,N_14954,N_14983);
xor UO_1499 (O_1499,N_14796,N_14615);
and UO_1500 (O_1500,N_14658,N_14843);
nor UO_1501 (O_1501,N_14521,N_14411);
or UO_1502 (O_1502,N_14585,N_14316);
xnor UO_1503 (O_1503,N_14280,N_14285);
and UO_1504 (O_1504,N_14909,N_14697);
or UO_1505 (O_1505,N_14733,N_14265);
or UO_1506 (O_1506,N_14631,N_14615);
or UO_1507 (O_1507,N_14916,N_14993);
nor UO_1508 (O_1508,N_14500,N_14815);
nor UO_1509 (O_1509,N_14744,N_14551);
nor UO_1510 (O_1510,N_14429,N_14737);
and UO_1511 (O_1511,N_14537,N_14672);
nand UO_1512 (O_1512,N_14634,N_14823);
xor UO_1513 (O_1513,N_14771,N_14346);
and UO_1514 (O_1514,N_14840,N_14465);
or UO_1515 (O_1515,N_14993,N_14974);
xnor UO_1516 (O_1516,N_14633,N_14630);
nand UO_1517 (O_1517,N_14768,N_14603);
nor UO_1518 (O_1518,N_14851,N_14848);
xnor UO_1519 (O_1519,N_14470,N_14506);
xnor UO_1520 (O_1520,N_14261,N_14908);
and UO_1521 (O_1521,N_14551,N_14882);
nor UO_1522 (O_1522,N_14943,N_14505);
xnor UO_1523 (O_1523,N_14623,N_14417);
xnor UO_1524 (O_1524,N_14376,N_14355);
nor UO_1525 (O_1525,N_14251,N_14996);
and UO_1526 (O_1526,N_14814,N_14759);
nor UO_1527 (O_1527,N_14528,N_14787);
nand UO_1528 (O_1528,N_14879,N_14329);
or UO_1529 (O_1529,N_14836,N_14806);
nor UO_1530 (O_1530,N_14648,N_14741);
xor UO_1531 (O_1531,N_14511,N_14847);
and UO_1532 (O_1532,N_14332,N_14429);
and UO_1533 (O_1533,N_14296,N_14693);
or UO_1534 (O_1534,N_14284,N_14349);
and UO_1535 (O_1535,N_14725,N_14988);
nand UO_1536 (O_1536,N_14868,N_14845);
nor UO_1537 (O_1537,N_14383,N_14790);
or UO_1538 (O_1538,N_14794,N_14790);
xnor UO_1539 (O_1539,N_14733,N_14882);
or UO_1540 (O_1540,N_14432,N_14648);
nand UO_1541 (O_1541,N_14623,N_14784);
and UO_1542 (O_1542,N_14572,N_14349);
nand UO_1543 (O_1543,N_14451,N_14439);
and UO_1544 (O_1544,N_14624,N_14364);
or UO_1545 (O_1545,N_14666,N_14406);
or UO_1546 (O_1546,N_14481,N_14512);
or UO_1547 (O_1547,N_14982,N_14477);
nand UO_1548 (O_1548,N_14911,N_14346);
and UO_1549 (O_1549,N_14882,N_14642);
or UO_1550 (O_1550,N_14549,N_14698);
xnor UO_1551 (O_1551,N_14605,N_14596);
nand UO_1552 (O_1552,N_14723,N_14757);
nor UO_1553 (O_1553,N_14418,N_14588);
nand UO_1554 (O_1554,N_14892,N_14804);
and UO_1555 (O_1555,N_14893,N_14431);
or UO_1556 (O_1556,N_14433,N_14467);
and UO_1557 (O_1557,N_14589,N_14856);
and UO_1558 (O_1558,N_14920,N_14619);
or UO_1559 (O_1559,N_14850,N_14302);
nor UO_1560 (O_1560,N_14390,N_14487);
and UO_1561 (O_1561,N_14749,N_14409);
xor UO_1562 (O_1562,N_14976,N_14674);
and UO_1563 (O_1563,N_14930,N_14850);
or UO_1564 (O_1564,N_14471,N_14818);
nand UO_1565 (O_1565,N_14703,N_14542);
and UO_1566 (O_1566,N_14620,N_14870);
nor UO_1567 (O_1567,N_14913,N_14306);
xor UO_1568 (O_1568,N_14713,N_14897);
nand UO_1569 (O_1569,N_14340,N_14380);
nand UO_1570 (O_1570,N_14998,N_14799);
xor UO_1571 (O_1571,N_14631,N_14639);
nor UO_1572 (O_1572,N_14910,N_14613);
nor UO_1573 (O_1573,N_14602,N_14395);
nand UO_1574 (O_1574,N_14863,N_14484);
and UO_1575 (O_1575,N_14826,N_14264);
and UO_1576 (O_1576,N_14923,N_14317);
or UO_1577 (O_1577,N_14815,N_14425);
or UO_1578 (O_1578,N_14579,N_14969);
nor UO_1579 (O_1579,N_14581,N_14318);
and UO_1580 (O_1580,N_14839,N_14837);
and UO_1581 (O_1581,N_14405,N_14846);
nand UO_1582 (O_1582,N_14637,N_14283);
xnor UO_1583 (O_1583,N_14661,N_14673);
or UO_1584 (O_1584,N_14472,N_14872);
nand UO_1585 (O_1585,N_14976,N_14964);
nor UO_1586 (O_1586,N_14409,N_14768);
xnor UO_1587 (O_1587,N_14380,N_14279);
xor UO_1588 (O_1588,N_14773,N_14655);
and UO_1589 (O_1589,N_14695,N_14679);
and UO_1590 (O_1590,N_14635,N_14552);
or UO_1591 (O_1591,N_14290,N_14584);
or UO_1592 (O_1592,N_14392,N_14513);
and UO_1593 (O_1593,N_14556,N_14411);
or UO_1594 (O_1594,N_14864,N_14909);
nor UO_1595 (O_1595,N_14412,N_14662);
xor UO_1596 (O_1596,N_14422,N_14810);
nand UO_1597 (O_1597,N_14275,N_14613);
nor UO_1598 (O_1598,N_14695,N_14546);
or UO_1599 (O_1599,N_14913,N_14633);
xnor UO_1600 (O_1600,N_14825,N_14954);
nand UO_1601 (O_1601,N_14511,N_14335);
nand UO_1602 (O_1602,N_14721,N_14253);
nor UO_1603 (O_1603,N_14520,N_14731);
or UO_1604 (O_1604,N_14368,N_14638);
nor UO_1605 (O_1605,N_14477,N_14916);
xnor UO_1606 (O_1606,N_14516,N_14649);
and UO_1607 (O_1607,N_14957,N_14640);
and UO_1608 (O_1608,N_14557,N_14501);
and UO_1609 (O_1609,N_14786,N_14588);
or UO_1610 (O_1610,N_14569,N_14828);
or UO_1611 (O_1611,N_14602,N_14659);
and UO_1612 (O_1612,N_14960,N_14994);
nand UO_1613 (O_1613,N_14927,N_14301);
nand UO_1614 (O_1614,N_14606,N_14302);
or UO_1615 (O_1615,N_14332,N_14609);
or UO_1616 (O_1616,N_14580,N_14663);
and UO_1617 (O_1617,N_14879,N_14338);
xnor UO_1618 (O_1618,N_14942,N_14899);
nand UO_1619 (O_1619,N_14652,N_14884);
nand UO_1620 (O_1620,N_14924,N_14642);
nand UO_1621 (O_1621,N_14458,N_14924);
or UO_1622 (O_1622,N_14331,N_14666);
and UO_1623 (O_1623,N_14641,N_14699);
and UO_1624 (O_1624,N_14968,N_14307);
nor UO_1625 (O_1625,N_14307,N_14426);
nand UO_1626 (O_1626,N_14538,N_14723);
and UO_1627 (O_1627,N_14846,N_14839);
xnor UO_1628 (O_1628,N_14838,N_14593);
xnor UO_1629 (O_1629,N_14327,N_14917);
and UO_1630 (O_1630,N_14595,N_14366);
nand UO_1631 (O_1631,N_14946,N_14351);
xor UO_1632 (O_1632,N_14427,N_14342);
xnor UO_1633 (O_1633,N_14333,N_14561);
nor UO_1634 (O_1634,N_14561,N_14795);
or UO_1635 (O_1635,N_14628,N_14553);
xnor UO_1636 (O_1636,N_14282,N_14608);
nor UO_1637 (O_1637,N_14390,N_14364);
and UO_1638 (O_1638,N_14960,N_14837);
nor UO_1639 (O_1639,N_14951,N_14621);
nand UO_1640 (O_1640,N_14984,N_14569);
or UO_1641 (O_1641,N_14392,N_14279);
nand UO_1642 (O_1642,N_14948,N_14490);
or UO_1643 (O_1643,N_14741,N_14531);
or UO_1644 (O_1644,N_14900,N_14693);
xor UO_1645 (O_1645,N_14911,N_14735);
nor UO_1646 (O_1646,N_14774,N_14902);
or UO_1647 (O_1647,N_14787,N_14301);
xor UO_1648 (O_1648,N_14983,N_14681);
nor UO_1649 (O_1649,N_14589,N_14675);
and UO_1650 (O_1650,N_14869,N_14317);
xnor UO_1651 (O_1651,N_14496,N_14822);
nand UO_1652 (O_1652,N_14985,N_14395);
xnor UO_1653 (O_1653,N_14901,N_14641);
xor UO_1654 (O_1654,N_14368,N_14796);
xor UO_1655 (O_1655,N_14588,N_14339);
or UO_1656 (O_1656,N_14635,N_14272);
nor UO_1657 (O_1657,N_14427,N_14367);
nand UO_1658 (O_1658,N_14943,N_14935);
nor UO_1659 (O_1659,N_14256,N_14457);
nand UO_1660 (O_1660,N_14613,N_14318);
or UO_1661 (O_1661,N_14800,N_14758);
nor UO_1662 (O_1662,N_14511,N_14930);
and UO_1663 (O_1663,N_14983,N_14331);
or UO_1664 (O_1664,N_14501,N_14899);
or UO_1665 (O_1665,N_14616,N_14710);
and UO_1666 (O_1666,N_14282,N_14643);
nand UO_1667 (O_1667,N_14769,N_14528);
or UO_1668 (O_1668,N_14573,N_14866);
nand UO_1669 (O_1669,N_14377,N_14798);
or UO_1670 (O_1670,N_14779,N_14590);
or UO_1671 (O_1671,N_14352,N_14444);
nand UO_1672 (O_1672,N_14361,N_14373);
or UO_1673 (O_1673,N_14286,N_14599);
nand UO_1674 (O_1674,N_14749,N_14572);
nand UO_1675 (O_1675,N_14486,N_14402);
nor UO_1676 (O_1676,N_14610,N_14469);
and UO_1677 (O_1677,N_14573,N_14793);
nor UO_1678 (O_1678,N_14427,N_14417);
and UO_1679 (O_1679,N_14769,N_14652);
nor UO_1680 (O_1680,N_14956,N_14909);
nor UO_1681 (O_1681,N_14457,N_14971);
or UO_1682 (O_1682,N_14533,N_14616);
nor UO_1683 (O_1683,N_14820,N_14427);
xnor UO_1684 (O_1684,N_14652,N_14910);
xor UO_1685 (O_1685,N_14971,N_14669);
nor UO_1686 (O_1686,N_14387,N_14617);
or UO_1687 (O_1687,N_14768,N_14593);
or UO_1688 (O_1688,N_14761,N_14943);
and UO_1689 (O_1689,N_14276,N_14947);
or UO_1690 (O_1690,N_14757,N_14682);
or UO_1691 (O_1691,N_14744,N_14994);
or UO_1692 (O_1692,N_14260,N_14915);
nor UO_1693 (O_1693,N_14643,N_14663);
nor UO_1694 (O_1694,N_14669,N_14926);
nor UO_1695 (O_1695,N_14842,N_14798);
or UO_1696 (O_1696,N_14815,N_14574);
or UO_1697 (O_1697,N_14493,N_14549);
and UO_1698 (O_1698,N_14520,N_14759);
and UO_1699 (O_1699,N_14889,N_14661);
or UO_1700 (O_1700,N_14625,N_14312);
nand UO_1701 (O_1701,N_14517,N_14537);
xor UO_1702 (O_1702,N_14486,N_14831);
and UO_1703 (O_1703,N_14746,N_14549);
or UO_1704 (O_1704,N_14731,N_14773);
nand UO_1705 (O_1705,N_14914,N_14287);
nand UO_1706 (O_1706,N_14591,N_14521);
and UO_1707 (O_1707,N_14519,N_14912);
xor UO_1708 (O_1708,N_14898,N_14798);
xnor UO_1709 (O_1709,N_14874,N_14388);
and UO_1710 (O_1710,N_14902,N_14798);
nand UO_1711 (O_1711,N_14962,N_14704);
xnor UO_1712 (O_1712,N_14527,N_14905);
or UO_1713 (O_1713,N_14334,N_14646);
nand UO_1714 (O_1714,N_14888,N_14995);
or UO_1715 (O_1715,N_14671,N_14902);
xnor UO_1716 (O_1716,N_14483,N_14458);
xnor UO_1717 (O_1717,N_14506,N_14306);
nor UO_1718 (O_1718,N_14661,N_14769);
xor UO_1719 (O_1719,N_14648,N_14927);
nor UO_1720 (O_1720,N_14650,N_14978);
nor UO_1721 (O_1721,N_14714,N_14284);
nand UO_1722 (O_1722,N_14465,N_14965);
xnor UO_1723 (O_1723,N_14479,N_14363);
nor UO_1724 (O_1724,N_14798,N_14933);
or UO_1725 (O_1725,N_14303,N_14960);
or UO_1726 (O_1726,N_14286,N_14611);
xor UO_1727 (O_1727,N_14648,N_14975);
and UO_1728 (O_1728,N_14857,N_14725);
and UO_1729 (O_1729,N_14250,N_14601);
nor UO_1730 (O_1730,N_14265,N_14404);
and UO_1731 (O_1731,N_14448,N_14887);
and UO_1732 (O_1732,N_14816,N_14721);
xnor UO_1733 (O_1733,N_14863,N_14699);
xor UO_1734 (O_1734,N_14687,N_14780);
nor UO_1735 (O_1735,N_14978,N_14602);
and UO_1736 (O_1736,N_14261,N_14698);
nand UO_1737 (O_1737,N_14363,N_14635);
and UO_1738 (O_1738,N_14756,N_14493);
and UO_1739 (O_1739,N_14666,N_14587);
nor UO_1740 (O_1740,N_14931,N_14403);
nor UO_1741 (O_1741,N_14381,N_14882);
nand UO_1742 (O_1742,N_14679,N_14625);
nor UO_1743 (O_1743,N_14269,N_14587);
nand UO_1744 (O_1744,N_14973,N_14336);
or UO_1745 (O_1745,N_14763,N_14713);
and UO_1746 (O_1746,N_14542,N_14488);
nand UO_1747 (O_1747,N_14297,N_14982);
nor UO_1748 (O_1748,N_14579,N_14752);
and UO_1749 (O_1749,N_14927,N_14382);
and UO_1750 (O_1750,N_14655,N_14428);
nand UO_1751 (O_1751,N_14654,N_14979);
and UO_1752 (O_1752,N_14727,N_14823);
and UO_1753 (O_1753,N_14705,N_14626);
xnor UO_1754 (O_1754,N_14514,N_14711);
xor UO_1755 (O_1755,N_14380,N_14363);
nand UO_1756 (O_1756,N_14929,N_14834);
or UO_1757 (O_1757,N_14397,N_14942);
and UO_1758 (O_1758,N_14373,N_14303);
nand UO_1759 (O_1759,N_14778,N_14649);
or UO_1760 (O_1760,N_14866,N_14983);
and UO_1761 (O_1761,N_14867,N_14383);
and UO_1762 (O_1762,N_14951,N_14353);
xor UO_1763 (O_1763,N_14548,N_14918);
nand UO_1764 (O_1764,N_14319,N_14661);
xnor UO_1765 (O_1765,N_14601,N_14911);
and UO_1766 (O_1766,N_14491,N_14610);
nor UO_1767 (O_1767,N_14922,N_14691);
nor UO_1768 (O_1768,N_14580,N_14980);
and UO_1769 (O_1769,N_14750,N_14999);
nor UO_1770 (O_1770,N_14967,N_14868);
or UO_1771 (O_1771,N_14381,N_14528);
nor UO_1772 (O_1772,N_14897,N_14953);
or UO_1773 (O_1773,N_14943,N_14755);
nand UO_1774 (O_1774,N_14826,N_14489);
or UO_1775 (O_1775,N_14676,N_14470);
nand UO_1776 (O_1776,N_14465,N_14445);
or UO_1777 (O_1777,N_14657,N_14304);
xnor UO_1778 (O_1778,N_14428,N_14509);
nand UO_1779 (O_1779,N_14251,N_14900);
and UO_1780 (O_1780,N_14809,N_14910);
or UO_1781 (O_1781,N_14577,N_14892);
xor UO_1782 (O_1782,N_14671,N_14879);
and UO_1783 (O_1783,N_14484,N_14784);
or UO_1784 (O_1784,N_14417,N_14547);
xor UO_1785 (O_1785,N_14896,N_14821);
xor UO_1786 (O_1786,N_14398,N_14988);
nand UO_1787 (O_1787,N_14940,N_14825);
nor UO_1788 (O_1788,N_14792,N_14947);
nand UO_1789 (O_1789,N_14821,N_14356);
nor UO_1790 (O_1790,N_14967,N_14650);
and UO_1791 (O_1791,N_14667,N_14720);
xnor UO_1792 (O_1792,N_14477,N_14420);
or UO_1793 (O_1793,N_14810,N_14797);
xnor UO_1794 (O_1794,N_14885,N_14430);
nor UO_1795 (O_1795,N_14717,N_14473);
or UO_1796 (O_1796,N_14446,N_14315);
and UO_1797 (O_1797,N_14664,N_14724);
xor UO_1798 (O_1798,N_14819,N_14507);
nand UO_1799 (O_1799,N_14319,N_14777);
or UO_1800 (O_1800,N_14255,N_14759);
and UO_1801 (O_1801,N_14925,N_14490);
nand UO_1802 (O_1802,N_14822,N_14867);
and UO_1803 (O_1803,N_14287,N_14498);
nand UO_1804 (O_1804,N_14954,N_14269);
xnor UO_1805 (O_1805,N_14475,N_14434);
nor UO_1806 (O_1806,N_14807,N_14573);
nor UO_1807 (O_1807,N_14269,N_14993);
nand UO_1808 (O_1808,N_14571,N_14461);
nand UO_1809 (O_1809,N_14666,N_14656);
nor UO_1810 (O_1810,N_14606,N_14826);
nor UO_1811 (O_1811,N_14751,N_14798);
nand UO_1812 (O_1812,N_14424,N_14769);
nor UO_1813 (O_1813,N_14792,N_14428);
nand UO_1814 (O_1814,N_14740,N_14482);
and UO_1815 (O_1815,N_14434,N_14827);
xnor UO_1816 (O_1816,N_14484,N_14648);
nand UO_1817 (O_1817,N_14982,N_14737);
xor UO_1818 (O_1818,N_14508,N_14999);
xnor UO_1819 (O_1819,N_14906,N_14607);
and UO_1820 (O_1820,N_14374,N_14260);
nand UO_1821 (O_1821,N_14344,N_14618);
or UO_1822 (O_1822,N_14530,N_14968);
nand UO_1823 (O_1823,N_14672,N_14328);
xnor UO_1824 (O_1824,N_14435,N_14307);
xnor UO_1825 (O_1825,N_14528,N_14827);
xnor UO_1826 (O_1826,N_14494,N_14430);
nand UO_1827 (O_1827,N_14689,N_14506);
and UO_1828 (O_1828,N_14261,N_14710);
nand UO_1829 (O_1829,N_14800,N_14685);
xor UO_1830 (O_1830,N_14833,N_14507);
nor UO_1831 (O_1831,N_14391,N_14980);
or UO_1832 (O_1832,N_14349,N_14522);
xor UO_1833 (O_1833,N_14338,N_14594);
and UO_1834 (O_1834,N_14962,N_14884);
nor UO_1835 (O_1835,N_14347,N_14533);
nor UO_1836 (O_1836,N_14619,N_14655);
nor UO_1837 (O_1837,N_14864,N_14450);
and UO_1838 (O_1838,N_14385,N_14980);
nand UO_1839 (O_1839,N_14787,N_14565);
xnor UO_1840 (O_1840,N_14886,N_14928);
nand UO_1841 (O_1841,N_14628,N_14705);
nor UO_1842 (O_1842,N_14752,N_14407);
nor UO_1843 (O_1843,N_14331,N_14403);
xor UO_1844 (O_1844,N_14848,N_14459);
nand UO_1845 (O_1845,N_14707,N_14370);
nor UO_1846 (O_1846,N_14549,N_14330);
nor UO_1847 (O_1847,N_14708,N_14806);
or UO_1848 (O_1848,N_14866,N_14823);
or UO_1849 (O_1849,N_14805,N_14850);
nor UO_1850 (O_1850,N_14681,N_14894);
nand UO_1851 (O_1851,N_14766,N_14954);
and UO_1852 (O_1852,N_14904,N_14484);
and UO_1853 (O_1853,N_14318,N_14756);
nor UO_1854 (O_1854,N_14804,N_14539);
nand UO_1855 (O_1855,N_14273,N_14795);
nor UO_1856 (O_1856,N_14772,N_14300);
nor UO_1857 (O_1857,N_14818,N_14664);
and UO_1858 (O_1858,N_14544,N_14558);
and UO_1859 (O_1859,N_14503,N_14304);
and UO_1860 (O_1860,N_14789,N_14539);
nor UO_1861 (O_1861,N_14420,N_14887);
nand UO_1862 (O_1862,N_14849,N_14321);
xor UO_1863 (O_1863,N_14834,N_14252);
nor UO_1864 (O_1864,N_14839,N_14308);
nand UO_1865 (O_1865,N_14474,N_14695);
or UO_1866 (O_1866,N_14709,N_14669);
and UO_1867 (O_1867,N_14859,N_14834);
xor UO_1868 (O_1868,N_14428,N_14555);
or UO_1869 (O_1869,N_14500,N_14587);
nor UO_1870 (O_1870,N_14683,N_14870);
nor UO_1871 (O_1871,N_14606,N_14975);
and UO_1872 (O_1872,N_14492,N_14664);
nor UO_1873 (O_1873,N_14668,N_14441);
and UO_1874 (O_1874,N_14650,N_14508);
xnor UO_1875 (O_1875,N_14771,N_14831);
nor UO_1876 (O_1876,N_14497,N_14889);
xnor UO_1877 (O_1877,N_14791,N_14264);
nor UO_1878 (O_1878,N_14643,N_14964);
nor UO_1879 (O_1879,N_14307,N_14718);
or UO_1880 (O_1880,N_14734,N_14279);
xnor UO_1881 (O_1881,N_14898,N_14774);
nor UO_1882 (O_1882,N_14318,N_14476);
nor UO_1883 (O_1883,N_14569,N_14876);
nor UO_1884 (O_1884,N_14649,N_14287);
nand UO_1885 (O_1885,N_14760,N_14743);
xor UO_1886 (O_1886,N_14538,N_14396);
nor UO_1887 (O_1887,N_14621,N_14534);
and UO_1888 (O_1888,N_14955,N_14912);
or UO_1889 (O_1889,N_14583,N_14593);
or UO_1890 (O_1890,N_14432,N_14502);
or UO_1891 (O_1891,N_14381,N_14770);
and UO_1892 (O_1892,N_14682,N_14328);
and UO_1893 (O_1893,N_14765,N_14734);
and UO_1894 (O_1894,N_14639,N_14738);
nand UO_1895 (O_1895,N_14431,N_14305);
xnor UO_1896 (O_1896,N_14581,N_14400);
nor UO_1897 (O_1897,N_14759,N_14924);
or UO_1898 (O_1898,N_14328,N_14846);
and UO_1899 (O_1899,N_14778,N_14607);
xor UO_1900 (O_1900,N_14264,N_14552);
nor UO_1901 (O_1901,N_14490,N_14536);
xnor UO_1902 (O_1902,N_14998,N_14511);
nor UO_1903 (O_1903,N_14726,N_14563);
or UO_1904 (O_1904,N_14323,N_14562);
nor UO_1905 (O_1905,N_14627,N_14572);
xnor UO_1906 (O_1906,N_14504,N_14899);
xnor UO_1907 (O_1907,N_14330,N_14487);
or UO_1908 (O_1908,N_14623,N_14332);
nand UO_1909 (O_1909,N_14578,N_14916);
or UO_1910 (O_1910,N_14589,N_14957);
xor UO_1911 (O_1911,N_14609,N_14840);
nor UO_1912 (O_1912,N_14674,N_14888);
nand UO_1913 (O_1913,N_14888,N_14493);
or UO_1914 (O_1914,N_14720,N_14682);
nand UO_1915 (O_1915,N_14272,N_14889);
and UO_1916 (O_1916,N_14733,N_14952);
nand UO_1917 (O_1917,N_14830,N_14380);
or UO_1918 (O_1918,N_14486,N_14724);
or UO_1919 (O_1919,N_14333,N_14688);
nand UO_1920 (O_1920,N_14459,N_14587);
and UO_1921 (O_1921,N_14984,N_14796);
nand UO_1922 (O_1922,N_14437,N_14379);
and UO_1923 (O_1923,N_14659,N_14812);
and UO_1924 (O_1924,N_14481,N_14566);
nand UO_1925 (O_1925,N_14872,N_14307);
nand UO_1926 (O_1926,N_14495,N_14668);
nor UO_1927 (O_1927,N_14252,N_14478);
nand UO_1928 (O_1928,N_14556,N_14702);
and UO_1929 (O_1929,N_14384,N_14309);
nor UO_1930 (O_1930,N_14462,N_14951);
xor UO_1931 (O_1931,N_14520,N_14315);
nand UO_1932 (O_1932,N_14826,N_14906);
and UO_1933 (O_1933,N_14779,N_14988);
and UO_1934 (O_1934,N_14270,N_14287);
xnor UO_1935 (O_1935,N_14442,N_14966);
and UO_1936 (O_1936,N_14973,N_14420);
nor UO_1937 (O_1937,N_14565,N_14744);
or UO_1938 (O_1938,N_14452,N_14493);
xor UO_1939 (O_1939,N_14582,N_14375);
nand UO_1940 (O_1940,N_14916,N_14814);
and UO_1941 (O_1941,N_14499,N_14271);
xnor UO_1942 (O_1942,N_14869,N_14315);
and UO_1943 (O_1943,N_14596,N_14713);
xor UO_1944 (O_1944,N_14736,N_14445);
or UO_1945 (O_1945,N_14638,N_14269);
or UO_1946 (O_1946,N_14480,N_14664);
or UO_1947 (O_1947,N_14453,N_14918);
and UO_1948 (O_1948,N_14588,N_14349);
nor UO_1949 (O_1949,N_14579,N_14526);
or UO_1950 (O_1950,N_14370,N_14503);
xor UO_1951 (O_1951,N_14820,N_14778);
and UO_1952 (O_1952,N_14350,N_14334);
and UO_1953 (O_1953,N_14301,N_14958);
xor UO_1954 (O_1954,N_14515,N_14927);
nor UO_1955 (O_1955,N_14848,N_14310);
and UO_1956 (O_1956,N_14497,N_14890);
nand UO_1957 (O_1957,N_14409,N_14571);
nand UO_1958 (O_1958,N_14546,N_14356);
nand UO_1959 (O_1959,N_14945,N_14445);
nand UO_1960 (O_1960,N_14991,N_14676);
or UO_1961 (O_1961,N_14628,N_14632);
or UO_1962 (O_1962,N_14740,N_14393);
or UO_1963 (O_1963,N_14306,N_14631);
xor UO_1964 (O_1964,N_14913,N_14527);
nor UO_1965 (O_1965,N_14460,N_14858);
or UO_1966 (O_1966,N_14846,N_14909);
nor UO_1967 (O_1967,N_14897,N_14671);
nor UO_1968 (O_1968,N_14840,N_14504);
or UO_1969 (O_1969,N_14646,N_14567);
or UO_1970 (O_1970,N_14657,N_14703);
or UO_1971 (O_1971,N_14306,N_14538);
nand UO_1972 (O_1972,N_14454,N_14658);
xor UO_1973 (O_1973,N_14661,N_14424);
xnor UO_1974 (O_1974,N_14742,N_14276);
xnor UO_1975 (O_1975,N_14267,N_14833);
nor UO_1976 (O_1976,N_14293,N_14477);
and UO_1977 (O_1977,N_14272,N_14898);
nor UO_1978 (O_1978,N_14657,N_14332);
or UO_1979 (O_1979,N_14996,N_14770);
nand UO_1980 (O_1980,N_14464,N_14627);
nor UO_1981 (O_1981,N_14688,N_14315);
nand UO_1982 (O_1982,N_14945,N_14400);
or UO_1983 (O_1983,N_14334,N_14957);
nand UO_1984 (O_1984,N_14777,N_14581);
or UO_1985 (O_1985,N_14901,N_14511);
or UO_1986 (O_1986,N_14252,N_14999);
nand UO_1987 (O_1987,N_14690,N_14352);
xor UO_1988 (O_1988,N_14364,N_14594);
or UO_1989 (O_1989,N_14456,N_14498);
or UO_1990 (O_1990,N_14791,N_14297);
or UO_1991 (O_1991,N_14871,N_14458);
or UO_1992 (O_1992,N_14599,N_14258);
nand UO_1993 (O_1993,N_14347,N_14277);
or UO_1994 (O_1994,N_14949,N_14800);
nor UO_1995 (O_1995,N_14401,N_14429);
or UO_1996 (O_1996,N_14970,N_14817);
nand UO_1997 (O_1997,N_14844,N_14442);
or UO_1998 (O_1998,N_14456,N_14351);
nand UO_1999 (O_1999,N_14678,N_14942);
endmodule