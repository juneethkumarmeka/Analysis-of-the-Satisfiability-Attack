module basic_1000_10000_1500_5_levels_1xor_1(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999;
xor U0 (N_0,In_61,In_351);
and U1 (N_1,In_659,In_909);
and U2 (N_2,In_560,In_486);
nor U3 (N_3,In_704,In_869);
nor U4 (N_4,In_160,In_209);
and U5 (N_5,In_628,In_271);
nor U6 (N_6,In_763,In_754);
nor U7 (N_7,In_948,In_641);
nand U8 (N_8,In_432,In_158);
nand U9 (N_9,In_205,In_278);
nor U10 (N_10,In_377,In_988);
or U11 (N_11,In_855,In_56);
nand U12 (N_12,In_602,In_630);
nor U13 (N_13,In_406,In_940);
nor U14 (N_14,In_256,In_541);
nand U15 (N_15,In_171,In_549);
xnor U16 (N_16,In_424,In_725);
or U17 (N_17,In_224,In_885);
nor U18 (N_18,In_305,In_149);
or U19 (N_19,In_287,In_732);
or U20 (N_20,In_671,In_814);
or U21 (N_21,In_748,In_753);
and U22 (N_22,In_186,In_874);
or U23 (N_23,In_567,In_657);
nor U24 (N_24,In_309,In_78);
nand U25 (N_25,In_901,In_579);
or U26 (N_26,In_756,In_174);
nor U27 (N_27,In_41,In_584);
and U28 (N_28,In_286,In_841);
and U29 (N_29,In_319,In_267);
or U30 (N_30,In_582,In_290);
nor U31 (N_31,In_871,In_606);
and U32 (N_32,In_53,In_744);
and U33 (N_33,In_137,In_778);
nor U34 (N_34,In_735,In_288);
nor U35 (N_35,In_879,In_345);
nand U36 (N_36,In_572,In_955);
or U37 (N_37,In_875,In_935);
or U38 (N_38,In_957,In_916);
nand U39 (N_39,In_244,In_85);
and U40 (N_40,In_552,In_525);
and U41 (N_41,In_425,In_636);
nor U42 (N_42,In_777,In_787);
nor U43 (N_43,In_326,In_383);
nor U44 (N_44,In_682,In_890);
nor U45 (N_45,In_862,In_76);
and U46 (N_46,In_20,In_173);
and U47 (N_47,In_699,In_611);
and U48 (N_48,In_485,In_896);
and U49 (N_49,In_818,In_736);
nand U50 (N_50,In_134,In_164);
or U51 (N_51,In_446,In_551);
and U52 (N_52,In_713,In_369);
nand U53 (N_53,In_973,In_404);
and U54 (N_54,In_831,In_431);
or U55 (N_55,In_182,In_124);
and U56 (N_56,In_811,In_22);
nand U57 (N_57,In_199,In_632);
nor U58 (N_58,In_429,In_302);
or U59 (N_59,In_996,In_58);
or U60 (N_60,In_332,In_907);
nor U61 (N_61,In_846,In_29);
and U62 (N_62,In_557,In_556);
nand U63 (N_63,In_615,In_532);
nor U64 (N_64,In_791,In_21);
or U65 (N_65,In_655,In_397);
nor U66 (N_66,In_511,In_422);
nand U67 (N_67,In_553,In_263);
or U68 (N_68,In_2,In_788);
or U69 (N_69,In_453,In_361);
or U70 (N_70,In_71,In_410);
nor U71 (N_71,In_497,In_133);
and U72 (N_72,In_707,In_842);
nand U73 (N_73,In_917,In_922);
nor U74 (N_74,In_793,In_587);
and U75 (N_75,In_508,In_280);
and U76 (N_76,In_574,In_747);
and U77 (N_77,In_172,In_884);
nor U78 (N_78,In_543,In_334);
nand U79 (N_79,In_324,In_591);
or U80 (N_80,In_703,In_38);
and U81 (N_81,In_573,In_755);
nand U82 (N_82,In_784,In_765);
nand U83 (N_83,In_733,In_315);
or U84 (N_84,In_32,In_720);
and U85 (N_85,In_193,In_110);
nand U86 (N_86,In_63,In_986);
xor U87 (N_87,In_356,In_154);
and U88 (N_88,In_605,In_570);
or U89 (N_89,In_537,In_692);
nor U90 (N_90,In_207,In_662);
nand U91 (N_91,In_65,In_336);
nor U92 (N_92,In_937,In_761);
and U93 (N_93,In_312,In_254);
or U94 (N_94,In_604,In_48);
or U95 (N_95,In_652,In_499);
and U96 (N_96,In_740,In_146);
nor U97 (N_97,In_34,In_766);
and U98 (N_98,In_318,In_64);
and U99 (N_99,In_418,In_168);
and U100 (N_100,In_536,In_170);
nand U101 (N_101,In_35,In_125);
nor U102 (N_102,In_350,In_459);
or U103 (N_103,In_179,In_304);
or U104 (N_104,In_313,In_514);
or U105 (N_105,In_321,In_638);
nand U106 (N_106,In_214,In_307);
or U107 (N_107,In_129,In_365);
nor U108 (N_108,In_165,In_196);
or U109 (N_109,In_674,In_946);
or U110 (N_110,In_27,In_46);
or U111 (N_111,In_565,In_741);
or U112 (N_112,In_442,In_643);
or U113 (N_113,In_999,In_989);
or U114 (N_114,In_598,In_443);
nor U115 (N_115,In_140,In_7);
and U116 (N_116,In_650,In_681);
or U117 (N_117,In_633,In_200);
or U118 (N_118,In_191,In_337);
xor U119 (N_119,In_131,In_440);
nand U120 (N_120,In_272,In_329);
and U121 (N_121,In_858,In_863);
nand U122 (N_122,In_283,In_822);
and U123 (N_123,In_669,In_163);
and U124 (N_124,In_375,In_931);
nand U125 (N_125,In_436,In_184);
or U126 (N_126,In_281,In_159);
and U127 (N_127,In_227,In_127);
nand U128 (N_128,In_435,In_969);
nor U129 (N_129,In_419,In_757);
nor U130 (N_130,In_112,In_434);
nand U131 (N_131,In_387,In_391);
nor U132 (N_132,In_107,In_210);
and U133 (N_133,In_603,In_300);
nand U134 (N_134,In_684,In_796);
nand U135 (N_135,In_547,In_496);
or U136 (N_136,In_92,In_839);
nor U137 (N_137,In_555,In_672);
nor U138 (N_138,In_379,In_843);
or U139 (N_139,In_36,In_382);
nand U140 (N_140,In_428,In_881);
or U141 (N_141,In_228,In_359);
and U142 (N_142,In_562,In_18);
nand U143 (N_143,In_403,In_201);
or U144 (N_144,In_62,In_762);
nand U145 (N_145,In_771,In_490);
or U146 (N_146,In_117,In_780);
nor U147 (N_147,In_866,In_581);
nor U148 (N_148,In_226,In_677);
and U149 (N_149,In_921,In_729);
nand U150 (N_150,In_792,In_625);
nand U151 (N_151,In_120,In_223);
nand U152 (N_152,In_631,In_279);
and U153 (N_153,In_231,In_348);
nor U154 (N_154,In_390,In_489);
nand U155 (N_155,In_507,In_370);
nand U156 (N_156,In_724,In_772);
and U157 (N_157,In_232,In_9);
or U158 (N_158,In_229,In_142);
nand U159 (N_159,In_847,In_526);
nor U160 (N_160,In_666,In_971);
nor U161 (N_161,In_143,In_972);
or U162 (N_162,In_743,In_688);
nor U163 (N_163,In_798,In_904);
nor U164 (N_164,In_530,In_84);
nand U165 (N_165,In_456,In_487);
or U166 (N_166,In_396,In_820);
and U167 (N_167,In_686,In_920);
nor U168 (N_168,In_706,In_39);
nor U169 (N_169,In_248,In_953);
nand U170 (N_170,In_176,In_910);
or U171 (N_171,In_538,In_306);
or U172 (N_172,In_468,In_457);
nor U173 (N_173,In_190,In_658);
nand U174 (N_174,In_601,In_216);
nand U175 (N_175,In_647,In_644);
or U176 (N_176,In_482,In_401);
nor U177 (N_177,In_219,In_276);
and U178 (N_178,In_258,In_634);
nor U179 (N_179,In_180,In_296);
or U180 (N_180,In_333,In_421);
nand U181 (N_181,In_696,In_141);
or U182 (N_182,In_540,In_376);
or U183 (N_183,In_919,In_926);
or U184 (N_184,In_883,In_640);
nand U185 (N_185,In_451,In_979);
or U186 (N_186,In_455,In_402);
nor U187 (N_187,In_575,In_42);
and U188 (N_188,In_308,In_806);
nor U189 (N_189,In_646,In_15);
nand U190 (N_190,In_578,In_568);
nor U191 (N_191,In_670,In_262);
and U192 (N_192,In_607,In_167);
nor U193 (N_193,In_259,In_995);
and U194 (N_194,In_779,In_679);
or U195 (N_195,In_651,In_810);
or U196 (N_196,In_360,In_566);
and U197 (N_197,In_135,In_510);
nand U198 (N_198,In_477,In_89);
nor U199 (N_199,In_983,In_664);
nand U200 (N_200,In_970,In_548);
or U201 (N_201,In_119,In_204);
nor U202 (N_202,In_534,In_93);
nor U203 (N_203,In_524,In_785);
nor U204 (N_204,In_824,In_82);
and U205 (N_205,In_389,In_962);
and U206 (N_206,In_801,In_592);
or U207 (N_207,In_899,In_518);
nor U208 (N_208,In_840,In_100);
and U209 (N_209,In_794,In_963);
nand U210 (N_210,In_430,In_569);
or U211 (N_211,In_83,In_246);
or U212 (N_212,In_407,In_113);
or U213 (N_213,In_411,In_997);
or U214 (N_214,In_195,In_166);
or U215 (N_215,In_817,In_230);
nand U216 (N_216,In_466,In_414);
or U217 (N_217,In_177,In_799);
or U218 (N_218,In_412,In_114);
or U219 (N_219,In_265,In_234);
or U220 (N_220,In_752,In_576);
nor U221 (N_221,In_738,In_994);
nor U222 (N_222,In_803,In_284);
and U223 (N_223,In_225,In_75);
or U224 (N_224,In_366,In_484);
and U225 (N_225,In_493,In_938);
nor U226 (N_226,In_268,In_739);
and U227 (N_227,In_197,In_624);
nand U228 (N_228,In_54,In_836);
or U229 (N_229,In_106,In_895);
and U230 (N_230,In_373,In_368);
or U231 (N_231,In_861,In_721);
or U232 (N_232,In_14,In_249);
nor U233 (N_233,In_545,In_723);
and U234 (N_234,In_586,In_878);
nand U235 (N_235,In_104,In_668);
nor U236 (N_236,In_797,In_608);
and U237 (N_237,In_903,In_610);
and U238 (N_238,In_161,In_807);
nand U239 (N_239,In_597,In_564);
xor U240 (N_240,In_790,In_138);
and U241 (N_241,In_915,In_795);
or U242 (N_242,In_472,In_423);
nor U243 (N_243,In_709,In_561);
nor U244 (N_244,In_452,In_645);
nor U245 (N_245,In_469,In_891);
nor U246 (N_246,In_90,In_449);
nand U247 (N_247,In_894,In_868);
nor U248 (N_248,In_372,In_23);
or U249 (N_249,In_417,In_257);
or U250 (N_250,In_123,In_388);
and U251 (N_251,In_954,In_776);
and U252 (N_252,In_447,In_491);
nor U253 (N_253,In_595,In_947);
nor U254 (N_254,In_355,In_620);
and U255 (N_255,In_266,In_8);
nand U256 (N_256,In_661,In_936);
and U257 (N_257,In_301,In_4);
or U258 (N_258,In_458,In_212);
nor U259 (N_259,In_950,In_531);
nor U260 (N_260,In_533,In_67);
nor U261 (N_261,In_28,In_589);
or U262 (N_262,In_5,In_585);
nor U263 (N_263,In_465,In_642);
or U264 (N_264,In_52,In_464);
and U265 (N_265,In_69,In_719);
nand U266 (N_266,In_588,In_888);
and U267 (N_267,In_208,In_660);
or U268 (N_268,In_439,In_450);
and U269 (N_269,In_235,In_619);
nor U270 (N_270,In_978,In_77);
and U271 (N_271,In_832,In_789);
or U272 (N_272,In_653,In_854);
or U273 (N_273,In_277,In_74);
nand U274 (N_274,In_57,In_448);
nor U275 (N_275,In_714,In_539);
or U276 (N_276,In_162,In_101);
or U277 (N_277,In_577,In_949);
or U278 (N_278,In_136,In_51);
nand U279 (N_279,In_317,In_483);
nand U280 (N_280,In_88,In_804);
nor U281 (N_281,In_364,In_151);
nor U282 (N_282,In_700,In_813);
nor U283 (N_283,In_961,In_520);
or U284 (N_284,In_665,In_902);
nor U285 (N_285,In_678,In_600);
nor U286 (N_286,In_908,In_928);
or U287 (N_287,In_358,In_467);
nand U288 (N_288,In_498,In_378);
nand U289 (N_289,In_764,In_105);
or U290 (N_290,In_691,In_19);
and U291 (N_291,In_217,In_852);
and U292 (N_292,In_60,In_405);
nor U293 (N_293,In_758,In_6);
and U294 (N_294,In_261,In_775);
nand U295 (N_295,In_590,In_274);
nand U296 (N_296,In_941,In_716);
nand U297 (N_297,In_320,In_238);
nor U298 (N_298,In_649,In_66);
nand U299 (N_299,In_900,In_596);
and U300 (N_300,In_374,In_500);
nand U301 (N_301,In_346,In_509);
nor U302 (N_302,In_966,In_745);
nand U303 (N_303,In_685,In_623);
or U304 (N_304,In_148,In_815);
or U305 (N_305,In_175,In_275);
nor U306 (N_306,In_139,In_96);
and U307 (N_307,In_689,In_87);
nand U308 (N_308,In_50,In_825);
and U309 (N_309,In_37,In_132);
nand U310 (N_310,In_192,In_635);
and U311 (N_311,In_55,In_952);
nand U312 (N_312,In_554,In_914);
nor U313 (N_313,In_654,In_897);
nor U314 (N_314,In_357,In_233);
nand U315 (N_315,In_558,In_478);
nor U316 (N_316,In_857,In_701);
and U317 (N_317,In_715,In_918);
or U318 (N_318,In_844,In_294);
nor U319 (N_319,In_583,In_43);
and U320 (N_320,In_49,In_338);
nor U321 (N_321,In_956,In_220);
or U322 (N_322,In_959,In_599);
and U323 (N_323,In_222,In_945);
and U324 (N_324,In_951,In_354);
nor U325 (N_325,In_639,In_16);
and U326 (N_326,In_121,In_399);
nand U327 (N_327,In_853,In_236);
nand U328 (N_328,In_929,In_991);
or U329 (N_329,In_103,In_98);
or U330 (N_330,In_710,In_479);
nor U331 (N_331,In_363,In_86);
or U332 (N_332,In_218,In_697);
and U333 (N_333,In_958,In_981);
nand U334 (N_334,In_297,In_471);
and U335 (N_335,In_802,In_718);
or U336 (N_336,In_827,In_816);
or U337 (N_337,In_830,In_282);
nand U338 (N_338,In_728,In_693);
nand U339 (N_339,In_616,In_512);
and U340 (N_340,In_990,In_473);
nor U341 (N_341,In_749,In_144);
or U342 (N_342,In_385,In_698);
nand U343 (N_343,In_157,In_726);
or U344 (N_344,In_829,In_310);
and U345 (N_345,In_504,In_759);
or U346 (N_346,In_99,In_325);
and U347 (N_347,In_426,In_993);
nand U348 (N_348,In_438,In_108);
and U349 (N_349,In_571,In_445);
nand U350 (N_350,In_934,In_960);
and U351 (N_351,In_240,In_476);
or U352 (N_352,In_343,In_559);
nand U353 (N_353,In_837,In_712);
nor U354 (N_354,In_349,In_239);
nor U355 (N_355,In_147,In_462);
nand U356 (N_356,In_59,In_45);
nor U357 (N_357,In_155,In_40);
and U358 (N_358,In_250,In_328);
or U359 (N_359,In_474,In_933);
nand U360 (N_360,In_913,In_683);
nor U361 (N_361,In_344,In_269);
or U362 (N_362,In_594,In_202);
nor U363 (N_363,In_94,In_911);
and U364 (N_364,In_347,In_152);
and U365 (N_365,In_188,In_260);
nor U366 (N_366,In_505,In_734);
and U367 (N_367,In_339,In_834);
nor U368 (N_368,In_11,In_626);
nand U369 (N_369,In_408,In_394);
and U370 (N_370,In_109,In_398);
and U371 (N_371,In_433,In_31);
nand U372 (N_372,In_495,In_609);
nand U373 (N_373,In_169,In_116);
and U374 (N_374,In_835,In_47);
or U375 (N_375,In_331,In_289);
and U376 (N_376,In_675,In_877);
and U377 (N_377,In_711,In_461);
nor U378 (N_378,In_145,In_515);
nand U379 (N_379,In_905,In_912);
nand U380 (N_380,In_245,In_115);
and U381 (N_381,In_695,In_298);
nor U382 (N_382,In_156,In_44);
nor U383 (N_383,In_295,In_24);
or U384 (N_384,In_550,In_821);
nor U385 (N_385,In_415,In_242);
and U386 (N_386,In_30,In_544);
nor U387 (N_387,In_270,In_454);
or U388 (N_388,In_867,In_393);
nor U389 (N_389,In_705,In_965);
nor U390 (N_390,In_189,In_181);
or U391 (N_391,In_26,In_864);
nor U392 (N_392,In_676,In_1);
nand U393 (N_393,In_335,In_845);
or U394 (N_394,In_255,In_826);
or U395 (N_395,In_314,In_648);
or U396 (N_396,In_898,In_870);
nand U397 (N_397,In_859,In_656);
or U398 (N_398,In_980,In_198);
nand U399 (N_399,In_828,In_95);
and U400 (N_400,In_542,In_72);
nand U401 (N_401,In_667,In_617);
nand U402 (N_402,In_808,In_621);
or U403 (N_403,In_494,In_805);
nor U404 (N_404,In_0,In_717);
nor U405 (N_405,In_273,In_441);
or U406 (N_406,In_91,In_800);
or U407 (N_407,In_985,In_727);
nand U408 (N_408,In_774,In_856);
nor U409 (N_409,In_687,In_944);
and U410 (N_410,In_968,In_342);
nor U411 (N_411,In_786,In_247);
and U412 (N_412,In_243,In_722);
or U413 (N_413,In_241,In_882);
nand U414 (N_414,In_481,In_211);
or U415 (N_415,In_923,In_111);
or U416 (N_416,In_849,In_593);
or U417 (N_417,In_976,In_444);
nand U418 (N_418,In_299,In_3);
nand U419 (N_419,In_975,In_291);
nor U420 (N_420,In_81,In_880);
nand U421 (N_421,In_984,In_409);
or U422 (N_422,In_506,In_130);
and U423 (N_423,In_128,In_460);
nor U424 (N_424,In_618,In_386);
nor U425 (N_425,In_939,In_519);
nand U426 (N_426,In_527,In_833);
or U427 (N_427,In_237,In_528);
nor U428 (N_428,In_702,In_475);
nor U429 (N_429,In_708,In_927);
nand U430 (N_430,In_742,In_185);
nand U431 (N_431,In_889,In_352);
and U432 (N_432,In_535,In_783);
or U433 (N_433,In_876,In_860);
nand U434 (N_434,In_663,In_851);
and U435 (N_435,In_673,In_812);
nor U436 (N_436,In_427,In_153);
or U437 (N_437,In_637,In_694);
and U438 (N_438,In_327,In_150);
nor U439 (N_439,In_760,In_68);
and U440 (N_440,In_480,In_213);
nand U441 (N_441,In_420,In_215);
or U442 (N_442,In_400,In_384);
nor U443 (N_443,In_513,In_942);
or U444 (N_444,In_886,In_178);
or U445 (N_445,In_930,In_292);
and U446 (N_446,In_353,In_768);
nor U447 (N_447,In_80,In_967);
and U448 (N_448,In_848,In_850);
and U449 (N_449,In_492,In_503);
nand U450 (N_450,In_629,In_982);
or U451 (N_451,In_680,In_380);
and U452 (N_452,In_887,In_769);
nor U453 (N_453,In_964,In_122);
nor U454 (N_454,In_516,In_470);
nand U455 (N_455,In_70,In_322);
nor U456 (N_456,In_79,In_341);
or U457 (N_457,In_872,In_819);
or U458 (N_458,In_529,In_770);
nand U459 (N_459,In_194,In_906);
or U460 (N_460,In_17,In_251);
or U461 (N_461,In_612,In_463);
and U462 (N_462,In_932,In_622);
or U463 (N_463,In_838,In_523);
and U464 (N_464,In_746,In_118);
and U465 (N_465,In_252,In_943);
nand U466 (N_466,In_781,In_187);
nand U467 (N_467,In_285,In_340);
or U468 (N_468,In_737,In_751);
nor U469 (N_469,In_413,In_311);
nor U470 (N_470,In_102,In_97);
nor U471 (N_471,In_893,In_362);
or U472 (N_472,In_614,In_416);
nor U473 (N_473,In_330,In_782);
and U474 (N_474,In_998,In_323);
nand U475 (N_475,In_627,In_750);
nand U476 (N_476,In_13,In_206);
nor U477 (N_477,In_367,In_73);
nand U478 (N_478,In_731,In_865);
xnor U479 (N_479,In_264,In_126);
or U480 (N_480,In_521,In_580);
or U481 (N_481,In_253,In_546);
nand U482 (N_482,In_977,In_183);
nand U483 (N_483,In_987,In_773);
or U484 (N_484,In_809,In_974);
and U485 (N_485,In_873,In_892);
nand U486 (N_486,In_613,In_501);
or U487 (N_487,In_517,In_502);
and U488 (N_488,In_316,In_12);
nand U489 (N_489,In_767,In_33);
nor U490 (N_490,In_823,In_293);
and U491 (N_491,In_392,In_381);
nand U492 (N_492,In_488,In_303);
and U493 (N_493,In_924,In_437);
and U494 (N_494,In_221,In_925);
nand U495 (N_495,In_522,In_371);
or U496 (N_496,In_563,In_25);
nand U497 (N_497,In_10,In_690);
and U498 (N_498,In_395,In_992);
nor U499 (N_499,In_203,In_730);
or U500 (N_500,In_887,In_790);
and U501 (N_501,In_662,In_564);
or U502 (N_502,In_166,In_449);
xnor U503 (N_503,In_433,In_122);
nor U504 (N_504,In_149,In_932);
or U505 (N_505,In_838,In_229);
or U506 (N_506,In_975,In_907);
and U507 (N_507,In_52,In_891);
nand U508 (N_508,In_695,In_248);
or U509 (N_509,In_651,In_522);
nor U510 (N_510,In_748,In_732);
nand U511 (N_511,In_653,In_296);
nor U512 (N_512,In_671,In_683);
nor U513 (N_513,In_36,In_332);
and U514 (N_514,In_216,In_457);
or U515 (N_515,In_21,In_15);
nand U516 (N_516,In_148,In_260);
or U517 (N_517,In_818,In_12);
or U518 (N_518,In_576,In_50);
nor U519 (N_519,In_187,In_904);
and U520 (N_520,In_752,In_412);
and U521 (N_521,In_9,In_236);
or U522 (N_522,In_598,In_406);
and U523 (N_523,In_695,In_759);
nand U524 (N_524,In_315,In_888);
or U525 (N_525,In_452,In_560);
nand U526 (N_526,In_242,In_523);
or U527 (N_527,In_739,In_738);
nor U528 (N_528,In_900,In_796);
nand U529 (N_529,In_537,In_7);
and U530 (N_530,In_323,In_440);
and U531 (N_531,In_231,In_737);
nand U532 (N_532,In_453,In_5);
nand U533 (N_533,In_935,In_191);
or U534 (N_534,In_174,In_919);
and U535 (N_535,In_710,In_942);
or U536 (N_536,In_562,In_956);
or U537 (N_537,In_534,In_616);
nand U538 (N_538,In_152,In_797);
nor U539 (N_539,In_726,In_284);
nor U540 (N_540,In_797,In_123);
and U541 (N_541,In_339,In_247);
or U542 (N_542,In_153,In_117);
and U543 (N_543,In_421,In_293);
or U544 (N_544,In_704,In_845);
and U545 (N_545,In_460,In_538);
nor U546 (N_546,In_146,In_937);
and U547 (N_547,In_249,In_473);
nor U548 (N_548,In_358,In_603);
and U549 (N_549,In_701,In_876);
or U550 (N_550,In_792,In_698);
nor U551 (N_551,In_539,In_518);
nand U552 (N_552,In_885,In_165);
nand U553 (N_553,In_220,In_911);
and U554 (N_554,In_486,In_878);
nor U555 (N_555,In_595,In_676);
nand U556 (N_556,In_940,In_56);
nand U557 (N_557,In_101,In_147);
nor U558 (N_558,In_628,In_807);
or U559 (N_559,In_842,In_515);
or U560 (N_560,In_0,In_466);
nor U561 (N_561,In_382,In_731);
nand U562 (N_562,In_225,In_432);
nor U563 (N_563,In_310,In_801);
nand U564 (N_564,In_831,In_769);
and U565 (N_565,In_538,In_546);
or U566 (N_566,In_30,In_128);
nor U567 (N_567,In_255,In_440);
nor U568 (N_568,In_736,In_873);
nand U569 (N_569,In_949,In_505);
or U570 (N_570,In_46,In_698);
and U571 (N_571,In_144,In_68);
nand U572 (N_572,In_137,In_187);
nor U573 (N_573,In_77,In_293);
nor U574 (N_574,In_623,In_92);
nor U575 (N_575,In_885,In_251);
nand U576 (N_576,In_862,In_425);
or U577 (N_577,In_239,In_33);
or U578 (N_578,In_24,In_468);
or U579 (N_579,In_455,In_683);
and U580 (N_580,In_938,In_595);
nand U581 (N_581,In_693,In_880);
or U582 (N_582,In_832,In_831);
or U583 (N_583,In_254,In_902);
nor U584 (N_584,In_887,In_570);
or U585 (N_585,In_750,In_616);
and U586 (N_586,In_109,In_448);
nor U587 (N_587,In_580,In_371);
or U588 (N_588,In_313,In_755);
or U589 (N_589,In_729,In_900);
nor U590 (N_590,In_655,In_59);
and U591 (N_591,In_695,In_299);
and U592 (N_592,In_456,In_848);
nand U593 (N_593,In_969,In_800);
nor U594 (N_594,In_130,In_708);
and U595 (N_595,In_741,In_83);
or U596 (N_596,In_765,In_817);
nor U597 (N_597,In_873,In_707);
nand U598 (N_598,In_847,In_366);
nor U599 (N_599,In_678,In_261);
nor U600 (N_600,In_790,In_888);
nor U601 (N_601,In_52,In_208);
or U602 (N_602,In_824,In_966);
nor U603 (N_603,In_166,In_509);
nor U604 (N_604,In_822,In_101);
and U605 (N_605,In_539,In_255);
nor U606 (N_606,In_821,In_737);
xor U607 (N_607,In_142,In_109);
and U608 (N_608,In_929,In_425);
or U609 (N_609,In_52,In_245);
nor U610 (N_610,In_194,In_886);
nor U611 (N_611,In_111,In_486);
nand U612 (N_612,In_109,In_477);
nand U613 (N_613,In_915,In_162);
or U614 (N_614,In_714,In_98);
or U615 (N_615,In_526,In_527);
nor U616 (N_616,In_673,In_616);
nor U617 (N_617,In_67,In_153);
nor U618 (N_618,In_756,In_982);
nand U619 (N_619,In_521,In_971);
nor U620 (N_620,In_258,In_92);
or U621 (N_621,In_157,In_806);
nor U622 (N_622,In_921,In_736);
or U623 (N_623,In_672,In_883);
and U624 (N_624,In_65,In_143);
nor U625 (N_625,In_200,In_260);
or U626 (N_626,In_865,In_613);
or U627 (N_627,In_72,In_235);
nor U628 (N_628,In_448,In_94);
nand U629 (N_629,In_791,In_273);
nand U630 (N_630,In_938,In_20);
or U631 (N_631,In_603,In_294);
and U632 (N_632,In_137,In_249);
nor U633 (N_633,In_950,In_642);
or U634 (N_634,In_901,In_284);
or U635 (N_635,In_484,In_175);
nor U636 (N_636,In_720,In_493);
and U637 (N_637,In_98,In_505);
and U638 (N_638,In_569,In_195);
nor U639 (N_639,In_64,In_74);
nor U640 (N_640,In_950,In_272);
or U641 (N_641,In_451,In_603);
nand U642 (N_642,In_337,In_178);
nand U643 (N_643,In_985,In_641);
or U644 (N_644,In_409,In_635);
nor U645 (N_645,In_711,In_915);
and U646 (N_646,In_689,In_16);
and U647 (N_647,In_731,In_394);
or U648 (N_648,In_45,In_903);
and U649 (N_649,In_642,In_344);
nor U650 (N_650,In_508,In_332);
nand U651 (N_651,In_544,In_272);
nor U652 (N_652,In_855,In_131);
or U653 (N_653,In_84,In_201);
and U654 (N_654,In_858,In_229);
or U655 (N_655,In_313,In_607);
or U656 (N_656,In_932,In_797);
nand U657 (N_657,In_140,In_550);
and U658 (N_658,In_598,In_843);
nor U659 (N_659,In_677,In_802);
or U660 (N_660,In_462,In_282);
or U661 (N_661,In_160,In_499);
nor U662 (N_662,In_890,In_560);
nand U663 (N_663,In_836,In_167);
nor U664 (N_664,In_612,In_381);
nor U665 (N_665,In_909,In_472);
or U666 (N_666,In_838,In_665);
and U667 (N_667,In_359,In_78);
nor U668 (N_668,In_807,In_849);
nand U669 (N_669,In_455,In_309);
or U670 (N_670,In_747,In_144);
nand U671 (N_671,In_818,In_371);
nand U672 (N_672,In_376,In_115);
and U673 (N_673,In_594,In_250);
nor U674 (N_674,In_226,In_434);
and U675 (N_675,In_890,In_270);
or U676 (N_676,In_787,In_58);
or U677 (N_677,In_89,In_532);
nand U678 (N_678,In_496,In_423);
or U679 (N_679,In_658,In_86);
nand U680 (N_680,In_602,In_103);
nand U681 (N_681,In_678,In_454);
or U682 (N_682,In_666,In_468);
nor U683 (N_683,In_494,In_2);
nand U684 (N_684,In_961,In_896);
or U685 (N_685,In_55,In_973);
nor U686 (N_686,In_124,In_839);
nor U687 (N_687,In_319,In_664);
or U688 (N_688,In_639,In_46);
or U689 (N_689,In_34,In_515);
or U690 (N_690,In_102,In_110);
and U691 (N_691,In_970,In_740);
or U692 (N_692,In_359,In_475);
and U693 (N_693,In_576,In_310);
nor U694 (N_694,In_875,In_774);
nand U695 (N_695,In_632,In_574);
nand U696 (N_696,In_621,In_728);
and U697 (N_697,In_280,In_363);
nor U698 (N_698,In_985,In_347);
and U699 (N_699,In_642,In_20);
and U700 (N_700,In_217,In_763);
nor U701 (N_701,In_493,In_134);
or U702 (N_702,In_255,In_960);
nor U703 (N_703,In_165,In_618);
nand U704 (N_704,In_140,In_497);
or U705 (N_705,In_168,In_73);
or U706 (N_706,In_136,In_544);
nor U707 (N_707,In_453,In_339);
or U708 (N_708,In_210,In_496);
or U709 (N_709,In_917,In_840);
nand U710 (N_710,In_153,In_696);
and U711 (N_711,In_215,In_228);
nor U712 (N_712,In_206,In_466);
or U713 (N_713,In_288,In_197);
nor U714 (N_714,In_845,In_380);
nand U715 (N_715,In_703,In_786);
and U716 (N_716,In_217,In_992);
or U717 (N_717,In_75,In_861);
or U718 (N_718,In_958,In_114);
nor U719 (N_719,In_821,In_238);
and U720 (N_720,In_679,In_995);
or U721 (N_721,In_981,In_116);
nand U722 (N_722,In_786,In_930);
or U723 (N_723,In_840,In_483);
and U724 (N_724,In_632,In_895);
or U725 (N_725,In_376,In_685);
xnor U726 (N_726,In_168,In_295);
nor U727 (N_727,In_144,In_250);
or U728 (N_728,In_325,In_40);
nor U729 (N_729,In_288,In_203);
xor U730 (N_730,In_260,In_293);
nor U731 (N_731,In_341,In_652);
nor U732 (N_732,In_444,In_203);
or U733 (N_733,In_629,In_666);
or U734 (N_734,In_462,In_216);
or U735 (N_735,In_347,In_105);
xor U736 (N_736,In_825,In_29);
and U737 (N_737,In_272,In_992);
or U738 (N_738,In_342,In_745);
and U739 (N_739,In_109,In_408);
or U740 (N_740,In_719,In_76);
nand U741 (N_741,In_905,In_853);
nor U742 (N_742,In_115,In_619);
nor U743 (N_743,In_149,In_644);
or U744 (N_744,In_695,In_823);
or U745 (N_745,In_787,In_758);
xnor U746 (N_746,In_891,In_278);
or U747 (N_747,In_907,In_968);
or U748 (N_748,In_582,In_842);
nand U749 (N_749,In_886,In_298);
and U750 (N_750,In_328,In_307);
and U751 (N_751,In_212,In_761);
and U752 (N_752,In_642,In_408);
nand U753 (N_753,In_201,In_704);
or U754 (N_754,In_376,In_35);
or U755 (N_755,In_833,In_856);
or U756 (N_756,In_760,In_689);
nand U757 (N_757,In_670,In_629);
and U758 (N_758,In_912,In_368);
and U759 (N_759,In_993,In_103);
nand U760 (N_760,In_672,In_919);
or U761 (N_761,In_537,In_974);
and U762 (N_762,In_121,In_43);
or U763 (N_763,In_485,In_181);
xnor U764 (N_764,In_146,In_105);
nand U765 (N_765,In_296,In_46);
nor U766 (N_766,In_281,In_491);
or U767 (N_767,In_111,In_928);
or U768 (N_768,In_294,In_575);
nand U769 (N_769,In_38,In_168);
or U770 (N_770,In_261,In_51);
nor U771 (N_771,In_535,In_751);
or U772 (N_772,In_604,In_59);
nor U773 (N_773,In_798,In_669);
nand U774 (N_774,In_552,In_721);
and U775 (N_775,In_208,In_76);
nand U776 (N_776,In_269,In_949);
nand U777 (N_777,In_405,In_660);
nand U778 (N_778,In_973,In_672);
nand U779 (N_779,In_890,In_700);
and U780 (N_780,In_22,In_414);
or U781 (N_781,In_663,In_549);
and U782 (N_782,In_242,In_269);
or U783 (N_783,In_780,In_663);
and U784 (N_784,In_548,In_342);
nor U785 (N_785,In_944,In_536);
and U786 (N_786,In_417,In_654);
and U787 (N_787,In_703,In_969);
or U788 (N_788,In_418,In_946);
or U789 (N_789,In_161,In_48);
nand U790 (N_790,In_11,In_903);
nand U791 (N_791,In_180,In_885);
nand U792 (N_792,In_604,In_205);
and U793 (N_793,In_511,In_175);
nand U794 (N_794,In_490,In_894);
or U795 (N_795,In_776,In_597);
nor U796 (N_796,In_847,In_35);
nand U797 (N_797,In_170,In_105);
nor U798 (N_798,In_952,In_296);
nand U799 (N_799,In_55,In_585);
and U800 (N_800,In_604,In_369);
or U801 (N_801,In_413,In_960);
nor U802 (N_802,In_382,In_197);
nand U803 (N_803,In_592,In_632);
and U804 (N_804,In_822,In_896);
nand U805 (N_805,In_320,In_227);
nand U806 (N_806,In_232,In_924);
or U807 (N_807,In_966,In_838);
nand U808 (N_808,In_697,In_539);
and U809 (N_809,In_367,In_961);
nor U810 (N_810,In_957,In_259);
or U811 (N_811,In_490,In_841);
or U812 (N_812,In_676,In_102);
and U813 (N_813,In_773,In_411);
and U814 (N_814,In_484,In_474);
and U815 (N_815,In_665,In_33);
nand U816 (N_816,In_334,In_450);
and U817 (N_817,In_148,In_487);
nand U818 (N_818,In_108,In_482);
xor U819 (N_819,In_613,In_517);
nor U820 (N_820,In_199,In_984);
nand U821 (N_821,In_260,In_938);
nand U822 (N_822,In_651,In_829);
and U823 (N_823,In_637,In_98);
nand U824 (N_824,In_769,In_566);
or U825 (N_825,In_704,In_284);
nand U826 (N_826,In_521,In_830);
nand U827 (N_827,In_813,In_337);
nand U828 (N_828,In_643,In_267);
nor U829 (N_829,In_917,In_550);
nand U830 (N_830,In_662,In_213);
nand U831 (N_831,In_917,In_277);
or U832 (N_832,In_100,In_723);
nor U833 (N_833,In_683,In_962);
nand U834 (N_834,In_35,In_853);
nor U835 (N_835,In_856,In_999);
nand U836 (N_836,In_25,In_605);
nor U837 (N_837,In_274,In_458);
and U838 (N_838,In_206,In_575);
nor U839 (N_839,In_535,In_888);
nor U840 (N_840,In_89,In_983);
or U841 (N_841,In_685,In_95);
or U842 (N_842,In_121,In_402);
nand U843 (N_843,In_183,In_596);
nor U844 (N_844,In_207,In_149);
nand U845 (N_845,In_388,In_786);
nor U846 (N_846,In_674,In_854);
nand U847 (N_847,In_618,In_326);
or U848 (N_848,In_586,In_861);
nor U849 (N_849,In_861,In_905);
nor U850 (N_850,In_75,In_41);
nand U851 (N_851,In_682,In_423);
nand U852 (N_852,In_213,In_720);
or U853 (N_853,In_185,In_670);
nand U854 (N_854,In_144,In_426);
or U855 (N_855,In_654,In_982);
and U856 (N_856,In_332,In_868);
nor U857 (N_857,In_796,In_433);
nor U858 (N_858,In_947,In_491);
or U859 (N_859,In_388,In_7);
nor U860 (N_860,In_81,In_256);
nor U861 (N_861,In_367,In_322);
and U862 (N_862,In_107,In_929);
or U863 (N_863,In_457,In_346);
nand U864 (N_864,In_853,In_631);
nor U865 (N_865,In_287,In_416);
or U866 (N_866,In_607,In_835);
or U867 (N_867,In_168,In_642);
nand U868 (N_868,In_738,In_976);
or U869 (N_869,In_734,In_768);
nor U870 (N_870,In_73,In_496);
or U871 (N_871,In_566,In_240);
and U872 (N_872,In_212,In_856);
and U873 (N_873,In_417,In_974);
nand U874 (N_874,In_374,In_532);
nor U875 (N_875,In_719,In_377);
nand U876 (N_876,In_130,In_628);
or U877 (N_877,In_835,In_420);
or U878 (N_878,In_605,In_959);
or U879 (N_879,In_88,In_604);
or U880 (N_880,In_695,In_961);
or U881 (N_881,In_159,In_926);
and U882 (N_882,In_734,In_462);
nand U883 (N_883,In_706,In_598);
or U884 (N_884,In_999,In_269);
or U885 (N_885,In_893,In_751);
or U886 (N_886,In_750,In_312);
or U887 (N_887,In_12,In_505);
or U888 (N_888,In_922,In_464);
and U889 (N_889,In_30,In_735);
nor U890 (N_890,In_142,In_562);
nand U891 (N_891,In_458,In_146);
nand U892 (N_892,In_579,In_229);
nor U893 (N_893,In_309,In_301);
nor U894 (N_894,In_739,In_270);
nor U895 (N_895,In_228,In_508);
and U896 (N_896,In_357,In_644);
and U897 (N_897,In_838,In_13);
nand U898 (N_898,In_945,In_225);
and U899 (N_899,In_572,In_545);
nor U900 (N_900,In_10,In_819);
nor U901 (N_901,In_537,In_0);
nor U902 (N_902,In_267,In_333);
or U903 (N_903,In_366,In_145);
or U904 (N_904,In_378,In_89);
and U905 (N_905,In_83,In_448);
nand U906 (N_906,In_992,In_481);
nor U907 (N_907,In_132,In_696);
nor U908 (N_908,In_817,In_23);
xor U909 (N_909,In_677,In_460);
nand U910 (N_910,In_504,In_349);
xor U911 (N_911,In_673,In_936);
nand U912 (N_912,In_495,In_768);
and U913 (N_913,In_891,In_892);
nand U914 (N_914,In_294,In_505);
xor U915 (N_915,In_865,In_661);
or U916 (N_916,In_930,In_18);
nand U917 (N_917,In_464,In_986);
and U918 (N_918,In_812,In_469);
nor U919 (N_919,In_743,In_813);
and U920 (N_920,In_521,In_604);
nand U921 (N_921,In_111,In_200);
and U922 (N_922,In_990,In_332);
nand U923 (N_923,In_129,In_639);
nand U924 (N_924,In_834,In_126);
xnor U925 (N_925,In_592,In_306);
or U926 (N_926,In_727,In_382);
or U927 (N_927,In_457,In_509);
and U928 (N_928,In_467,In_105);
and U929 (N_929,In_570,In_479);
and U930 (N_930,In_400,In_995);
nand U931 (N_931,In_936,In_35);
nor U932 (N_932,In_236,In_888);
nor U933 (N_933,In_534,In_670);
or U934 (N_934,In_87,In_906);
nor U935 (N_935,In_634,In_912);
nor U936 (N_936,In_539,In_318);
nand U937 (N_937,In_665,In_110);
nand U938 (N_938,In_525,In_553);
nand U939 (N_939,In_550,In_378);
nand U940 (N_940,In_248,In_973);
nor U941 (N_941,In_762,In_351);
nor U942 (N_942,In_942,In_455);
nand U943 (N_943,In_305,In_52);
xnor U944 (N_944,In_407,In_102);
nand U945 (N_945,In_864,In_710);
and U946 (N_946,In_240,In_397);
nand U947 (N_947,In_355,In_145);
nor U948 (N_948,In_857,In_881);
nor U949 (N_949,In_210,In_154);
nor U950 (N_950,In_975,In_626);
nor U951 (N_951,In_66,In_21);
nand U952 (N_952,In_454,In_168);
nand U953 (N_953,In_919,In_96);
nand U954 (N_954,In_347,In_245);
or U955 (N_955,In_270,In_710);
or U956 (N_956,In_920,In_862);
nor U957 (N_957,In_903,In_986);
and U958 (N_958,In_613,In_637);
nor U959 (N_959,In_38,In_403);
and U960 (N_960,In_514,In_251);
and U961 (N_961,In_985,In_713);
nor U962 (N_962,In_786,In_700);
nor U963 (N_963,In_142,In_430);
and U964 (N_964,In_629,In_485);
or U965 (N_965,In_917,In_769);
or U966 (N_966,In_992,In_942);
nand U967 (N_967,In_30,In_693);
or U968 (N_968,In_867,In_359);
and U969 (N_969,In_814,In_484);
nand U970 (N_970,In_850,In_975);
or U971 (N_971,In_500,In_472);
nand U972 (N_972,In_787,In_244);
nor U973 (N_973,In_712,In_747);
nand U974 (N_974,In_395,In_669);
nand U975 (N_975,In_505,In_120);
and U976 (N_976,In_904,In_87);
or U977 (N_977,In_117,In_62);
nor U978 (N_978,In_725,In_759);
and U979 (N_979,In_565,In_880);
and U980 (N_980,In_848,In_287);
nor U981 (N_981,In_737,In_523);
nand U982 (N_982,In_712,In_791);
or U983 (N_983,In_71,In_616);
and U984 (N_984,In_258,In_133);
and U985 (N_985,In_351,In_855);
or U986 (N_986,In_583,In_23);
or U987 (N_987,In_239,In_162);
nor U988 (N_988,In_63,In_768);
or U989 (N_989,In_983,In_276);
nand U990 (N_990,In_366,In_262);
or U991 (N_991,In_932,In_408);
xnor U992 (N_992,In_168,In_850);
nand U993 (N_993,In_649,In_722);
nor U994 (N_994,In_539,In_85);
nand U995 (N_995,In_330,In_911);
nor U996 (N_996,In_68,In_540);
and U997 (N_997,In_9,In_116);
or U998 (N_998,In_180,In_347);
or U999 (N_999,In_944,In_265);
and U1000 (N_1000,In_638,In_752);
nand U1001 (N_1001,In_633,In_279);
and U1002 (N_1002,In_106,In_243);
nor U1003 (N_1003,In_827,In_99);
nand U1004 (N_1004,In_203,In_780);
nor U1005 (N_1005,In_86,In_846);
or U1006 (N_1006,In_168,In_244);
nor U1007 (N_1007,In_549,In_910);
nor U1008 (N_1008,In_263,In_114);
or U1009 (N_1009,In_747,In_270);
nand U1010 (N_1010,In_290,In_491);
or U1011 (N_1011,In_389,In_695);
nor U1012 (N_1012,In_568,In_600);
nand U1013 (N_1013,In_325,In_117);
nor U1014 (N_1014,In_127,In_157);
and U1015 (N_1015,In_326,In_697);
nor U1016 (N_1016,In_660,In_101);
nor U1017 (N_1017,In_866,In_522);
nor U1018 (N_1018,In_281,In_576);
or U1019 (N_1019,In_305,In_775);
nor U1020 (N_1020,In_888,In_494);
nand U1021 (N_1021,In_10,In_594);
nor U1022 (N_1022,In_445,In_102);
and U1023 (N_1023,In_195,In_254);
nand U1024 (N_1024,In_412,In_170);
and U1025 (N_1025,In_143,In_170);
or U1026 (N_1026,In_371,In_632);
nand U1027 (N_1027,In_722,In_84);
nand U1028 (N_1028,In_288,In_37);
nor U1029 (N_1029,In_831,In_709);
or U1030 (N_1030,In_689,In_381);
nand U1031 (N_1031,In_114,In_221);
or U1032 (N_1032,In_8,In_419);
or U1033 (N_1033,In_453,In_50);
or U1034 (N_1034,In_251,In_269);
and U1035 (N_1035,In_389,In_753);
nor U1036 (N_1036,In_335,In_48);
or U1037 (N_1037,In_149,In_573);
nand U1038 (N_1038,In_159,In_355);
or U1039 (N_1039,In_398,In_174);
or U1040 (N_1040,In_928,In_523);
or U1041 (N_1041,In_940,In_227);
or U1042 (N_1042,In_596,In_86);
and U1043 (N_1043,In_545,In_94);
and U1044 (N_1044,In_32,In_275);
and U1045 (N_1045,In_771,In_704);
nand U1046 (N_1046,In_310,In_864);
and U1047 (N_1047,In_286,In_107);
nand U1048 (N_1048,In_846,In_17);
and U1049 (N_1049,In_316,In_131);
and U1050 (N_1050,In_738,In_488);
nor U1051 (N_1051,In_18,In_618);
and U1052 (N_1052,In_745,In_740);
or U1053 (N_1053,In_162,In_933);
nor U1054 (N_1054,In_584,In_770);
or U1055 (N_1055,In_802,In_928);
and U1056 (N_1056,In_283,In_806);
nor U1057 (N_1057,In_307,In_281);
or U1058 (N_1058,In_781,In_147);
and U1059 (N_1059,In_122,In_868);
nor U1060 (N_1060,In_100,In_682);
or U1061 (N_1061,In_300,In_455);
nand U1062 (N_1062,In_5,In_139);
nor U1063 (N_1063,In_521,In_120);
or U1064 (N_1064,In_806,In_961);
nor U1065 (N_1065,In_412,In_274);
xor U1066 (N_1066,In_762,In_829);
nor U1067 (N_1067,In_908,In_462);
or U1068 (N_1068,In_778,In_743);
or U1069 (N_1069,In_909,In_84);
nand U1070 (N_1070,In_407,In_333);
nand U1071 (N_1071,In_889,In_886);
nand U1072 (N_1072,In_258,In_738);
nor U1073 (N_1073,In_934,In_293);
and U1074 (N_1074,In_692,In_301);
nand U1075 (N_1075,In_611,In_601);
nand U1076 (N_1076,In_645,In_430);
nor U1077 (N_1077,In_701,In_845);
nand U1078 (N_1078,In_435,In_573);
and U1079 (N_1079,In_850,In_439);
nor U1080 (N_1080,In_716,In_44);
nand U1081 (N_1081,In_517,In_23);
and U1082 (N_1082,In_15,In_400);
nand U1083 (N_1083,In_792,In_451);
nand U1084 (N_1084,In_705,In_562);
and U1085 (N_1085,In_40,In_982);
nor U1086 (N_1086,In_831,In_72);
nand U1087 (N_1087,In_961,In_324);
and U1088 (N_1088,In_488,In_858);
nand U1089 (N_1089,In_808,In_525);
nand U1090 (N_1090,In_240,In_888);
nor U1091 (N_1091,In_13,In_533);
nor U1092 (N_1092,In_33,In_586);
xor U1093 (N_1093,In_632,In_527);
or U1094 (N_1094,In_415,In_108);
and U1095 (N_1095,In_741,In_284);
nor U1096 (N_1096,In_41,In_397);
and U1097 (N_1097,In_852,In_365);
or U1098 (N_1098,In_789,In_356);
nor U1099 (N_1099,In_844,In_521);
or U1100 (N_1100,In_540,In_942);
nor U1101 (N_1101,In_890,In_40);
nand U1102 (N_1102,In_431,In_144);
nand U1103 (N_1103,In_759,In_957);
nor U1104 (N_1104,In_161,In_73);
or U1105 (N_1105,In_194,In_874);
and U1106 (N_1106,In_599,In_680);
or U1107 (N_1107,In_299,In_407);
nand U1108 (N_1108,In_403,In_901);
nand U1109 (N_1109,In_684,In_664);
nand U1110 (N_1110,In_104,In_348);
nor U1111 (N_1111,In_976,In_489);
nor U1112 (N_1112,In_660,In_231);
or U1113 (N_1113,In_348,In_821);
and U1114 (N_1114,In_919,In_553);
nor U1115 (N_1115,In_589,In_566);
or U1116 (N_1116,In_845,In_21);
nor U1117 (N_1117,In_889,In_907);
or U1118 (N_1118,In_956,In_828);
nor U1119 (N_1119,In_404,In_603);
or U1120 (N_1120,In_416,In_587);
or U1121 (N_1121,In_552,In_462);
nor U1122 (N_1122,In_849,In_37);
nor U1123 (N_1123,In_709,In_751);
and U1124 (N_1124,In_482,In_648);
or U1125 (N_1125,In_122,In_904);
nand U1126 (N_1126,In_587,In_251);
nor U1127 (N_1127,In_222,In_347);
nor U1128 (N_1128,In_355,In_33);
nand U1129 (N_1129,In_819,In_132);
nand U1130 (N_1130,In_278,In_378);
and U1131 (N_1131,In_123,In_239);
nand U1132 (N_1132,In_587,In_881);
and U1133 (N_1133,In_807,In_84);
and U1134 (N_1134,In_162,In_664);
nand U1135 (N_1135,In_578,In_923);
and U1136 (N_1136,In_91,In_757);
and U1137 (N_1137,In_177,In_538);
nand U1138 (N_1138,In_87,In_266);
nand U1139 (N_1139,In_41,In_334);
or U1140 (N_1140,In_28,In_992);
nand U1141 (N_1141,In_235,In_585);
and U1142 (N_1142,In_318,In_750);
and U1143 (N_1143,In_318,In_886);
nand U1144 (N_1144,In_633,In_851);
or U1145 (N_1145,In_236,In_845);
or U1146 (N_1146,In_163,In_852);
nand U1147 (N_1147,In_298,In_52);
nand U1148 (N_1148,In_727,In_646);
nor U1149 (N_1149,In_303,In_986);
nor U1150 (N_1150,In_939,In_309);
or U1151 (N_1151,In_882,In_377);
nor U1152 (N_1152,In_479,In_622);
xnor U1153 (N_1153,In_386,In_551);
nand U1154 (N_1154,In_377,In_604);
and U1155 (N_1155,In_318,In_176);
or U1156 (N_1156,In_114,In_823);
nand U1157 (N_1157,In_222,In_382);
and U1158 (N_1158,In_680,In_378);
or U1159 (N_1159,In_70,In_847);
nor U1160 (N_1160,In_989,In_492);
nand U1161 (N_1161,In_929,In_912);
nand U1162 (N_1162,In_282,In_460);
nand U1163 (N_1163,In_162,In_582);
and U1164 (N_1164,In_379,In_461);
or U1165 (N_1165,In_815,In_76);
and U1166 (N_1166,In_429,In_418);
nand U1167 (N_1167,In_140,In_763);
or U1168 (N_1168,In_707,In_500);
or U1169 (N_1169,In_91,In_447);
nand U1170 (N_1170,In_99,In_589);
nand U1171 (N_1171,In_568,In_6);
nor U1172 (N_1172,In_283,In_708);
or U1173 (N_1173,In_634,In_488);
and U1174 (N_1174,In_33,In_104);
or U1175 (N_1175,In_592,In_413);
nand U1176 (N_1176,In_886,In_810);
nand U1177 (N_1177,In_95,In_271);
nor U1178 (N_1178,In_587,In_312);
and U1179 (N_1179,In_431,In_980);
xor U1180 (N_1180,In_826,In_219);
and U1181 (N_1181,In_303,In_725);
and U1182 (N_1182,In_255,In_919);
nor U1183 (N_1183,In_142,In_620);
nor U1184 (N_1184,In_432,In_181);
and U1185 (N_1185,In_310,In_372);
and U1186 (N_1186,In_112,In_17);
nor U1187 (N_1187,In_617,In_405);
xor U1188 (N_1188,In_157,In_118);
and U1189 (N_1189,In_906,In_424);
nand U1190 (N_1190,In_192,In_27);
nand U1191 (N_1191,In_583,In_384);
and U1192 (N_1192,In_34,In_76);
nor U1193 (N_1193,In_343,In_453);
and U1194 (N_1194,In_324,In_730);
nor U1195 (N_1195,In_69,In_81);
or U1196 (N_1196,In_862,In_507);
nand U1197 (N_1197,In_298,In_71);
nor U1198 (N_1198,In_652,In_316);
nand U1199 (N_1199,In_533,In_257);
and U1200 (N_1200,In_14,In_936);
or U1201 (N_1201,In_900,In_955);
nor U1202 (N_1202,In_94,In_13);
nor U1203 (N_1203,In_510,In_6);
nand U1204 (N_1204,In_578,In_105);
and U1205 (N_1205,In_765,In_561);
and U1206 (N_1206,In_883,In_639);
or U1207 (N_1207,In_938,In_389);
and U1208 (N_1208,In_710,In_997);
nand U1209 (N_1209,In_52,In_499);
nor U1210 (N_1210,In_921,In_142);
nand U1211 (N_1211,In_94,In_302);
or U1212 (N_1212,In_547,In_150);
nand U1213 (N_1213,In_689,In_593);
nand U1214 (N_1214,In_293,In_355);
or U1215 (N_1215,In_82,In_374);
and U1216 (N_1216,In_633,In_285);
nand U1217 (N_1217,In_621,In_946);
nor U1218 (N_1218,In_491,In_427);
nor U1219 (N_1219,In_26,In_548);
or U1220 (N_1220,In_422,In_300);
nand U1221 (N_1221,In_932,In_439);
and U1222 (N_1222,In_196,In_119);
nor U1223 (N_1223,In_25,In_890);
nand U1224 (N_1224,In_290,In_869);
or U1225 (N_1225,In_980,In_577);
and U1226 (N_1226,In_716,In_962);
or U1227 (N_1227,In_714,In_767);
nand U1228 (N_1228,In_808,In_495);
nand U1229 (N_1229,In_307,In_55);
or U1230 (N_1230,In_172,In_365);
or U1231 (N_1231,In_245,In_126);
nor U1232 (N_1232,In_154,In_969);
or U1233 (N_1233,In_541,In_364);
or U1234 (N_1234,In_535,In_473);
nand U1235 (N_1235,In_679,In_411);
nor U1236 (N_1236,In_360,In_715);
nor U1237 (N_1237,In_707,In_510);
nand U1238 (N_1238,In_982,In_560);
nand U1239 (N_1239,In_455,In_413);
and U1240 (N_1240,In_136,In_801);
or U1241 (N_1241,In_500,In_725);
nand U1242 (N_1242,In_443,In_134);
nor U1243 (N_1243,In_843,In_436);
nor U1244 (N_1244,In_999,In_252);
nor U1245 (N_1245,In_453,In_580);
nand U1246 (N_1246,In_16,In_163);
and U1247 (N_1247,In_137,In_772);
nor U1248 (N_1248,In_1,In_423);
nand U1249 (N_1249,In_738,In_88);
or U1250 (N_1250,In_3,In_371);
or U1251 (N_1251,In_464,In_796);
nand U1252 (N_1252,In_247,In_965);
or U1253 (N_1253,In_84,In_558);
and U1254 (N_1254,In_35,In_369);
nand U1255 (N_1255,In_756,In_337);
or U1256 (N_1256,In_908,In_231);
and U1257 (N_1257,In_79,In_803);
nor U1258 (N_1258,In_399,In_203);
or U1259 (N_1259,In_983,In_835);
nor U1260 (N_1260,In_297,In_362);
nor U1261 (N_1261,In_294,In_86);
nand U1262 (N_1262,In_124,In_5);
nand U1263 (N_1263,In_654,In_705);
or U1264 (N_1264,In_396,In_405);
nor U1265 (N_1265,In_311,In_97);
nand U1266 (N_1266,In_436,In_597);
nand U1267 (N_1267,In_870,In_125);
nor U1268 (N_1268,In_34,In_636);
nand U1269 (N_1269,In_151,In_340);
nor U1270 (N_1270,In_165,In_405);
nor U1271 (N_1271,In_439,In_2);
or U1272 (N_1272,In_288,In_27);
nand U1273 (N_1273,In_614,In_929);
nor U1274 (N_1274,In_922,In_705);
or U1275 (N_1275,In_353,In_185);
nor U1276 (N_1276,In_735,In_252);
nand U1277 (N_1277,In_466,In_154);
and U1278 (N_1278,In_773,In_339);
or U1279 (N_1279,In_550,In_619);
nor U1280 (N_1280,In_806,In_281);
nor U1281 (N_1281,In_569,In_514);
nor U1282 (N_1282,In_676,In_489);
nand U1283 (N_1283,In_529,In_498);
nand U1284 (N_1284,In_775,In_253);
or U1285 (N_1285,In_969,In_701);
nand U1286 (N_1286,In_732,In_301);
or U1287 (N_1287,In_747,In_344);
nor U1288 (N_1288,In_488,In_188);
and U1289 (N_1289,In_809,In_876);
nand U1290 (N_1290,In_941,In_101);
nand U1291 (N_1291,In_269,In_230);
nand U1292 (N_1292,In_368,In_137);
nor U1293 (N_1293,In_83,In_531);
and U1294 (N_1294,In_302,In_59);
nor U1295 (N_1295,In_264,In_371);
and U1296 (N_1296,In_983,In_318);
xor U1297 (N_1297,In_697,In_327);
and U1298 (N_1298,In_822,In_467);
nand U1299 (N_1299,In_119,In_922);
nand U1300 (N_1300,In_820,In_139);
or U1301 (N_1301,In_132,In_812);
nor U1302 (N_1302,In_250,In_44);
nand U1303 (N_1303,In_469,In_647);
nor U1304 (N_1304,In_769,In_205);
and U1305 (N_1305,In_979,In_18);
nand U1306 (N_1306,In_501,In_732);
nand U1307 (N_1307,In_216,In_712);
or U1308 (N_1308,In_502,In_40);
nand U1309 (N_1309,In_839,In_760);
and U1310 (N_1310,In_417,In_781);
and U1311 (N_1311,In_369,In_643);
or U1312 (N_1312,In_743,In_974);
nand U1313 (N_1313,In_495,In_280);
and U1314 (N_1314,In_360,In_519);
or U1315 (N_1315,In_725,In_443);
nand U1316 (N_1316,In_570,In_739);
nor U1317 (N_1317,In_610,In_28);
or U1318 (N_1318,In_710,In_878);
or U1319 (N_1319,In_595,In_579);
and U1320 (N_1320,In_922,In_95);
and U1321 (N_1321,In_704,In_829);
nor U1322 (N_1322,In_53,In_786);
nor U1323 (N_1323,In_86,In_350);
and U1324 (N_1324,In_951,In_115);
or U1325 (N_1325,In_406,In_705);
and U1326 (N_1326,In_773,In_940);
nand U1327 (N_1327,In_705,In_677);
nor U1328 (N_1328,In_944,In_656);
or U1329 (N_1329,In_159,In_106);
and U1330 (N_1330,In_963,In_859);
nand U1331 (N_1331,In_449,In_350);
and U1332 (N_1332,In_196,In_909);
or U1333 (N_1333,In_6,In_287);
nand U1334 (N_1334,In_240,In_156);
nor U1335 (N_1335,In_747,In_99);
or U1336 (N_1336,In_923,In_954);
and U1337 (N_1337,In_95,In_858);
nand U1338 (N_1338,In_520,In_559);
nand U1339 (N_1339,In_592,In_340);
nor U1340 (N_1340,In_748,In_191);
or U1341 (N_1341,In_363,In_27);
or U1342 (N_1342,In_504,In_296);
or U1343 (N_1343,In_703,In_589);
nor U1344 (N_1344,In_703,In_884);
or U1345 (N_1345,In_428,In_910);
nand U1346 (N_1346,In_302,In_535);
or U1347 (N_1347,In_26,In_179);
and U1348 (N_1348,In_133,In_655);
or U1349 (N_1349,In_958,In_16);
nand U1350 (N_1350,In_914,In_346);
nor U1351 (N_1351,In_673,In_375);
nand U1352 (N_1352,In_229,In_484);
nor U1353 (N_1353,In_938,In_16);
nand U1354 (N_1354,In_207,In_329);
and U1355 (N_1355,In_946,In_461);
nor U1356 (N_1356,In_295,In_251);
or U1357 (N_1357,In_270,In_358);
nand U1358 (N_1358,In_262,In_193);
nor U1359 (N_1359,In_590,In_289);
nor U1360 (N_1360,In_169,In_245);
and U1361 (N_1361,In_590,In_679);
nand U1362 (N_1362,In_269,In_118);
nand U1363 (N_1363,In_192,In_149);
nand U1364 (N_1364,In_843,In_967);
nand U1365 (N_1365,In_258,In_726);
nor U1366 (N_1366,In_143,In_936);
nand U1367 (N_1367,In_503,In_980);
and U1368 (N_1368,In_717,In_553);
nor U1369 (N_1369,In_629,In_290);
and U1370 (N_1370,In_980,In_391);
nand U1371 (N_1371,In_592,In_703);
or U1372 (N_1372,In_112,In_640);
and U1373 (N_1373,In_35,In_198);
nor U1374 (N_1374,In_472,In_708);
or U1375 (N_1375,In_708,In_988);
nand U1376 (N_1376,In_401,In_971);
nand U1377 (N_1377,In_804,In_197);
nor U1378 (N_1378,In_795,In_928);
or U1379 (N_1379,In_593,In_786);
nand U1380 (N_1380,In_872,In_845);
or U1381 (N_1381,In_875,In_662);
or U1382 (N_1382,In_395,In_668);
or U1383 (N_1383,In_866,In_212);
nor U1384 (N_1384,In_189,In_672);
nor U1385 (N_1385,In_862,In_970);
nand U1386 (N_1386,In_292,In_890);
and U1387 (N_1387,In_265,In_165);
nand U1388 (N_1388,In_759,In_328);
nand U1389 (N_1389,In_573,In_511);
nor U1390 (N_1390,In_843,In_246);
nor U1391 (N_1391,In_160,In_724);
or U1392 (N_1392,In_575,In_947);
or U1393 (N_1393,In_360,In_16);
or U1394 (N_1394,In_572,In_13);
or U1395 (N_1395,In_198,In_972);
nand U1396 (N_1396,In_819,In_278);
nand U1397 (N_1397,In_346,In_166);
and U1398 (N_1398,In_370,In_516);
and U1399 (N_1399,In_7,In_352);
nor U1400 (N_1400,In_534,In_497);
and U1401 (N_1401,In_880,In_446);
nand U1402 (N_1402,In_972,In_565);
or U1403 (N_1403,In_601,In_461);
and U1404 (N_1404,In_85,In_274);
and U1405 (N_1405,In_428,In_278);
and U1406 (N_1406,In_653,In_38);
nand U1407 (N_1407,In_751,In_635);
nor U1408 (N_1408,In_634,In_393);
and U1409 (N_1409,In_468,In_334);
or U1410 (N_1410,In_504,In_159);
nand U1411 (N_1411,In_169,In_532);
nand U1412 (N_1412,In_661,In_402);
nor U1413 (N_1413,In_22,In_568);
and U1414 (N_1414,In_319,In_754);
nor U1415 (N_1415,In_399,In_765);
nor U1416 (N_1416,In_266,In_800);
or U1417 (N_1417,In_866,In_904);
nor U1418 (N_1418,In_53,In_377);
nand U1419 (N_1419,In_716,In_979);
nand U1420 (N_1420,In_461,In_752);
and U1421 (N_1421,In_681,In_263);
nand U1422 (N_1422,In_221,In_206);
and U1423 (N_1423,In_529,In_376);
or U1424 (N_1424,In_381,In_526);
nand U1425 (N_1425,In_237,In_559);
or U1426 (N_1426,In_881,In_485);
nor U1427 (N_1427,In_724,In_648);
or U1428 (N_1428,In_794,In_863);
nor U1429 (N_1429,In_518,In_139);
and U1430 (N_1430,In_882,In_132);
or U1431 (N_1431,In_570,In_319);
nor U1432 (N_1432,In_629,In_402);
or U1433 (N_1433,In_851,In_255);
and U1434 (N_1434,In_136,In_924);
or U1435 (N_1435,In_918,In_78);
and U1436 (N_1436,In_599,In_132);
or U1437 (N_1437,In_876,In_544);
nor U1438 (N_1438,In_445,In_732);
or U1439 (N_1439,In_267,In_816);
nor U1440 (N_1440,In_14,In_921);
and U1441 (N_1441,In_415,In_813);
or U1442 (N_1442,In_119,In_570);
or U1443 (N_1443,In_478,In_104);
and U1444 (N_1444,In_123,In_992);
and U1445 (N_1445,In_29,In_414);
nand U1446 (N_1446,In_491,In_923);
or U1447 (N_1447,In_918,In_606);
nor U1448 (N_1448,In_252,In_990);
and U1449 (N_1449,In_775,In_655);
and U1450 (N_1450,In_257,In_613);
nand U1451 (N_1451,In_321,In_943);
or U1452 (N_1452,In_895,In_508);
nand U1453 (N_1453,In_262,In_563);
or U1454 (N_1454,In_107,In_701);
nor U1455 (N_1455,In_553,In_614);
nor U1456 (N_1456,In_832,In_437);
and U1457 (N_1457,In_675,In_340);
nor U1458 (N_1458,In_135,In_250);
or U1459 (N_1459,In_969,In_471);
or U1460 (N_1460,In_110,In_957);
xor U1461 (N_1461,In_587,In_529);
nand U1462 (N_1462,In_131,In_718);
xnor U1463 (N_1463,In_803,In_781);
or U1464 (N_1464,In_798,In_791);
nor U1465 (N_1465,In_760,In_514);
or U1466 (N_1466,In_77,In_41);
nand U1467 (N_1467,In_142,In_628);
and U1468 (N_1468,In_752,In_896);
nand U1469 (N_1469,In_881,In_578);
and U1470 (N_1470,In_672,In_184);
nor U1471 (N_1471,In_709,In_569);
nand U1472 (N_1472,In_272,In_928);
nor U1473 (N_1473,In_103,In_882);
and U1474 (N_1474,In_368,In_11);
or U1475 (N_1475,In_627,In_821);
nand U1476 (N_1476,In_500,In_923);
and U1477 (N_1477,In_530,In_896);
nor U1478 (N_1478,In_923,In_566);
and U1479 (N_1479,In_496,In_614);
or U1480 (N_1480,In_452,In_166);
or U1481 (N_1481,In_6,In_489);
and U1482 (N_1482,In_919,In_146);
and U1483 (N_1483,In_471,In_673);
nor U1484 (N_1484,In_428,In_825);
and U1485 (N_1485,In_838,In_860);
and U1486 (N_1486,In_985,In_907);
or U1487 (N_1487,In_983,In_592);
nor U1488 (N_1488,In_798,In_952);
and U1489 (N_1489,In_368,In_766);
nand U1490 (N_1490,In_880,In_194);
or U1491 (N_1491,In_417,In_648);
nand U1492 (N_1492,In_645,In_433);
and U1493 (N_1493,In_984,In_82);
or U1494 (N_1494,In_224,In_296);
and U1495 (N_1495,In_515,In_451);
and U1496 (N_1496,In_626,In_235);
nor U1497 (N_1497,In_999,In_801);
or U1498 (N_1498,In_862,In_328);
or U1499 (N_1499,In_259,In_802);
or U1500 (N_1500,In_75,In_11);
or U1501 (N_1501,In_656,In_373);
nor U1502 (N_1502,In_123,In_845);
and U1503 (N_1503,In_14,In_461);
or U1504 (N_1504,In_625,In_612);
or U1505 (N_1505,In_740,In_890);
or U1506 (N_1506,In_812,In_914);
nand U1507 (N_1507,In_227,In_437);
and U1508 (N_1508,In_475,In_911);
or U1509 (N_1509,In_148,In_471);
nor U1510 (N_1510,In_367,In_715);
and U1511 (N_1511,In_243,In_739);
nor U1512 (N_1512,In_113,In_268);
and U1513 (N_1513,In_779,In_104);
nor U1514 (N_1514,In_545,In_191);
or U1515 (N_1515,In_853,In_125);
nand U1516 (N_1516,In_375,In_118);
nand U1517 (N_1517,In_532,In_80);
nor U1518 (N_1518,In_503,In_153);
nand U1519 (N_1519,In_980,In_18);
or U1520 (N_1520,In_115,In_448);
nor U1521 (N_1521,In_684,In_305);
nand U1522 (N_1522,In_730,In_984);
and U1523 (N_1523,In_92,In_408);
nor U1524 (N_1524,In_39,In_610);
and U1525 (N_1525,In_415,In_469);
nand U1526 (N_1526,In_363,In_928);
and U1527 (N_1527,In_471,In_863);
or U1528 (N_1528,In_840,In_807);
nand U1529 (N_1529,In_886,In_144);
and U1530 (N_1530,In_139,In_975);
and U1531 (N_1531,In_135,In_713);
and U1532 (N_1532,In_237,In_969);
nand U1533 (N_1533,In_891,In_123);
or U1534 (N_1534,In_886,In_553);
nor U1535 (N_1535,In_421,In_193);
nand U1536 (N_1536,In_142,In_565);
nand U1537 (N_1537,In_105,In_248);
nand U1538 (N_1538,In_266,In_972);
or U1539 (N_1539,In_347,In_95);
and U1540 (N_1540,In_698,In_57);
nor U1541 (N_1541,In_38,In_495);
nand U1542 (N_1542,In_56,In_365);
nand U1543 (N_1543,In_704,In_328);
nor U1544 (N_1544,In_190,In_733);
nand U1545 (N_1545,In_359,In_122);
or U1546 (N_1546,In_480,In_604);
and U1547 (N_1547,In_842,In_905);
nor U1548 (N_1548,In_153,In_723);
nor U1549 (N_1549,In_260,In_342);
nand U1550 (N_1550,In_319,In_659);
nor U1551 (N_1551,In_538,In_702);
and U1552 (N_1552,In_460,In_280);
or U1553 (N_1553,In_224,In_557);
or U1554 (N_1554,In_976,In_488);
and U1555 (N_1555,In_894,In_843);
nor U1556 (N_1556,In_295,In_203);
nor U1557 (N_1557,In_260,In_43);
or U1558 (N_1558,In_551,In_27);
nand U1559 (N_1559,In_988,In_613);
and U1560 (N_1560,In_792,In_320);
nor U1561 (N_1561,In_368,In_806);
nand U1562 (N_1562,In_608,In_602);
nand U1563 (N_1563,In_399,In_126);
nand U1564 (N_1564,In_758,In_271);
or U1565 (N_1565,In_604,In_727);
or U1566 (N_1566,In_851,In_292);
or U1567 (N_1567,In_587,In_568);
nor U1568 (N_1568,In_242,In_378);
nand U1569 (N_1569,In_289,In_345);
nor U1570 (N_1570,In_441,In_5);
or U1571 (N_1571,In_315,In_124);
and U1572 (N_1572,In_588,In_503);
nand U1573 (N_1573,In_248,In_165);
nor U1574 (N_1574,In_60,In_901);
or U1575 (N_1575,In_659,In_190);
nand U1576 (N_1576,In_581,In_218);
nor U1577 (N_1577,In_865,In_225);
nand U1578 (N_1578,In_643,In_508);
nor U1579 (N_1579,In_93,In_521);
nand U1580 (N_1580,In_552,In_350);
nor U1581 (N_1581,In_843,In_388);
and U1582 (N_1582,In_664,In_333);
nand U1583 (N_1583,In_975,In_677);
nand U1584 (N_1584,In_11,In_606);
nand U1585 (N_1585,In_602,In_883);
nand U1586 (N_1586,In_885,In_817);
nand U1587 (N_1587,In_41,In_869);
nor U1588 (N_1588,In_245,In_652);
nand U1589 (N_1589,In_845,In_55);
nor U1590 (N_1590,In_383,In_918);
or U1591 (N_1591,In_492,In_582);
and U1592 (N_1592,In_938,In_382);
or U1593 (N_1593,In_792,In_888);
and U1594 (N_1594,In_63,In_384);
or U1595 (N_1595,In_509,In_149);
nand U1596 (N_1596,In_71,In_488);
nor U1597 (N_1597,In_714,In_908);
or U1598 (N_1598,In_253,In_219);
or U1599 (N_1599,In_344,In_971);
nor U1600 (N_1600,In_2,In_103);
nor U1601 (N_1601,In_219,In_151);
and U1602 (N_1602,In_349,In_82);
nand U1603 (N_1603,In_275,In_599);
or U1604 (N_1604,In_693,In_981);
nand U1605 (N_1605,In_650,In_860);
or U1606 (N_1606,In_299,In_820);
nand U1607 (N_1607,In_7,In_748);
or U1608 (N_1608,In_177,In_261);
nor U1609 (N_1609,In_482,In_141);
nand U1610 (N_1610,In_999,In_698);
nand U1611 (N_1611,In_843,In_99);
nor U1612 (N_1612,In_982,In_238);
nand U1613 (N_1613,In_441,In_841);
and U1614 (N_1614,In_816,In_187);
or U1615 (N_1615,In_453,In_393);
nor U1616 (N_1616,In_16,In_955);
or U1617 (N_1617,In_66,In_382);
nand U1618 (N_1618,In_361,In_82);
and U1619 (N_1619,In_555,In_805);
nor U1620 (N_1620,In_121,In_595);
nand U1621 (N_1621,In_188,In_832);
nand U1622 (N_1622,In_652,In_601);
or U1623 (N_1623,In_694,In_585);
nand U1624 (N_1624,In_519,In_124);
nand U1625 (N_1625,In_145,In_298);
nand U1626 (N_1626,In_297,In_140);
or U1627 (N_1627,In_474,In_664);
nand U1628 (N_1628,In_816,In_355);
nor U1629 (N_1629,In_718,In_316);
or U1630 (N_1630,In_596,In_765);
and U1631 (N_1631,In_673,In_158);
nor U1632 (N_1632,In_330,In_892);
or U1633 (N_1633,In_745,In_627);
nor U1634 (N_1634,In_433,In_870);
nand U1635 (N_1635,In_804,In_445);
or U1636 (N_1636,In_552,In_916);
nand U1637 (N_1637,In_69,In_489);
or U1638 (N_1638,In_392,In_183);
and U1639 (N_1639,In_424,In_404);
or U1640 (N_1640,In_46,In_304);
nor U1641 (N_1641,In_238,In_42);
nand U1642 (N_1642,In_925,In_563);
nor U1643 (N_1643,In_399,In_639);
nor U1644 (N_1644,In_196,In_281);
nand U1645 (N_1645,In_396,In_304);
nand U1646 (N_1646,In_732,In_589);
nor U1647 (N_1647,In_823,In_171);
nand U1648 (N_1648,In_999,In_773);
nor U1649 (N_1649,In_152,In_99);
or U1650 (N_1650,In_154,In_887);
nand U1651 (N_1651,In_520,In_33);
nand U1652 (N_1652,In_445,In_670);
nand U1653 (N_1653,In_109,In_93);
and U1654 (N_1654,In_429,In_40);
or U1655 (N_1655,In_130,In_200);
and U1656 (N_1656,In_1,In_104);
or U1657 (N_1657,In_237,In_155);
nand U1658 (N_1658,In_968,In_391);
nand U1659 (N_1659,In_906,In_747);
nor U1660 (N_1660,In_301,In_577);
nand U1661 (N_1661,In_64,In_441);
or U1662 (N_1662,In_322,In_156);
and U1663 (N_1663,In_914,In_427);
or U1664 (N_1664,In_318,In_106);
nor U1665 (N_1665,In_573,In_878);
and U1666 (N_1666,In_120,In_457);
or U1667 (N_1667,In_585,In_125);
and U1668 (N_1668,In_272,In_267);
and U1669 (N_1669,In_304,In_164);
and U1670 (N_1670,In_303,In_310);
nor U1671 (N_1671,In_55,In_342);
nor U1672 (N_1672,In_949,In_684);
nor U1673 (N_1673,In_160,In_318);
and U1674 (N_1674,In_124,In_486);
nand U1675 (N_1675,In_691,In_961);
nand U1676 (N_1676,In_810,In_709);
nand U1677 (N_1677,In_631,In_961);
and U1678 (N_1678,In_461,In_640);
or U1679 (N_1679,In_880,In_1);
and U1680 (N_1680,In_728,In_345);
nor U1681 (N_1681,In_290,In_49);
nand U1682 (N_1682,In_197,In_471);
and U1683 (N_1683,In_628,In_634);
nor U1684 (N_1684,In_664,In_387);
nor U1685 (N_1685,In_385,In_471);
xor U1686 (N_1686,In_987,In_390);
nand U1687 (N_1687,In_243,In_418);
and U1688 (N_1688,In_342,In_600);
nor U1689 (N_1689,In_261,In_517);
xnor U1690 (N_1690,In_378,In_46);
or U1691 (N_1691,In_152,In_133);
and U1692 (N_1692,In_455,In_491);
nand U1693 (N_1693,In_701,In_586);
nor U1694 (N_1694,In_905,In_997);
nand U1695 (N_1695,In_678,In_941);
and U1696 (N_1696,In_131,In_978);
nand U1697 (N_1697,In_223,In_258);
and U1698 (N_1698,In_372,In_750);
or U1699 (N_1699,In_982,In_693);
and U1700 (N_1700,In_163,In_528);
or U1701 (N_1701,In_544,In_39);
and U1702 (N_1702,In_280,In_671);
nor U1703 (N_1703,In_750,In_837);
and U1704 (N_1704,In_17,In_582);
nand U1705 (N_1705,In_381,In_739);
nand U1706 (N_1706,In_734,In_87);
and U1707 (N_1707,In_91,In_479);
nor U1708 (N_1708,In_751,In_65);
and U1709 (N_1709,In_978,In_585);
and U1710 (N_1710,In_74,In_19);
or U1711 (N_1711,In_698,In_143);
nand U1712 (N_1712,In_759,In_681);
nor U1713 (N_1713,In_961,In_260);
nor U1714 (N_1714,In_395,In_689);
nand U1715 (N_1715,In_895,In_390);
or U1716 (N_1716,In_198,In_416);
nor U1717 (N_1717,In_773,In_853);
xnor U1718 (N_1718,In_215,In_664);
or U1719 (N_1719,In_912,In_296);
nand U1720 (N_1720,In_70,In_382);
nand U1721 (N_1721,In_719,In_602);
nor U1722 (N_1722,In_35,In_469);
and U1723 (N_1723,In_751,In_112);
nor U1724 (N_1724,In_53,In_295);
nor U1725 (N_1725,In_443,In_962);
nor U1726 (N_1726,In_568,In_702);
nand U1727 (N_1727,In_664,In_137);
nand U1728 (N_1728,In_467,In_71);
nand U1729 (N_1729,In_405,In_143);
and U1730 (N_1730,In_122,In_847);
nand U1731 (N_1731,In_348,In_738);
or U1732 (N_1732,In_265,In_450);
and U1733 (N_1733,In_266,In_289);
nor U1734 (N_1734,In_890,In_348);
nand U1735 (N_1735,In_38,In_804);
or U1736 (N_1736,In_660,In_149);
or U1737 (N_1737,In_696,In_401);
or U1738 (N_1738,In_11,In_759);
or U1739 (N_1739,In_978,In_943);
and U1740 (N_1740,In_960,In_251);
nor U1741 (N_1741,In_695,In_790);
or U1742 (N_1742,In_224,In_672);
nor U1743 (N_1743,In_751,In_849);
or U1744 (N_1744,In_392,In_158);
or U1745 (N_1745,In_844,In_439);
and U1746 (N_1746,In_217,In_973);
xor U1747 (N_1747,In_148,In_628);
or U1748 (N_1748,In_657,In_209);
nor U1749 (N_1749,In_472,In_190);
and U1750 (N_1750,In_605,In_376);
or U1751 (N_1751,In_210,In_976);
and U1752 (N_1752,In_822,In_369);
nor U1753 (N_1753,In_772,In_541);
xnor U1754 (N_1754,In_153,In_789);
or U1755 (N_1755,In_156,In_989);
or U1756 (N_1756,In_986,In_998);
nand U1757 (N_1757,In_781,In_297);
or U1758 (N_1758,In_785,In_337);
or U1759 (N_1759,In_355,In_966);
or U1760 (N_1760,In_577,In_146);
or U1761 (N_1761,In_670,In_355);
nor U1762 (N_1762,In_833,In_903);
nand U1763 (N_1763,In_653,In_108);
or U1764 (N_1764,In_618,In_805);
and U1765 (N_1765,In_273,In_128);
or U1766 (N_1766,In_737,In_907);
or U1767 (N_1767,In_63,In_630);
and U1768 (N_1768,In_403,In_54);
and U1769 (N_1769,In_138,In_637);
nor U1770 (N_1770,In_422,In_166);
and U1771 (N_1771,In_839,In_750);
and U1772 (N_1772,In_54,In_595);
and U1773 (N_1773,In_213,In_171);
and U1774 (N_1774,In_136,In_933);
and U1775 (N_1775,In_360,In_727);
nand U1776 (N_1776,In_93,In_163);
or U1777 (N_1777,In_380,In_203);
nor U1778 (N_1778,In_287,In_498);
nand U1779 (N_1779,In_624,In_320);
nand U1780 (N_1780,In_496,In_50);
and U1781 (N_1781,In_154,In_554);
nand U1782 (N_1782,In_749,In_79);
nor U1783 (N_1783,In_744,In_432);
and U1784 (N_1784,In_357,In_68);
and U1785 (N_1785,In_201,In_605);
nor U1786 (N_1786,In_390,In_581);
nand U1787 (N_1787,In_475,In_484);
and U1788 (N_1788,In_355,In_397);
nand U1789 (N_1789,In_366,In_597);
nand U1790 (N_1790,In_806,In_671);
or U1791 (N_1791,In_628,In_798);
nor U1792 (N_1792,In_706,In_88);
or U1793 (N_1793,In_466,In_894);
nand U1794 (N_1794,In_574,In_41);
nor U1795 (N_1795,In_864,In_736);
nor U1796 (N_1796,In_945,In_564);
nand U1797 (N_1797,In_941,In_737);
and U1798 (N_1798,In_513,In_450);
nor U1799 (N_1799,In_5,In_4);
or U1800 (N_1800,In_573,In_339);
nand U1801 (N_1801,In_957,In_718);
nor U1802 (N_1802,In_115,In_5);
nand U1803 (N_1803,In_353,In_835);
or U1804 (N_1804,In_159,In_273);
and U1805 (N_1805,In_375,In_921);
nor U1806 (N_1806,In_284,In_245);
nand U1807 (N_1807,In_461,In_8);
nor U1808 (N_1808,In_14,In_204);
nand U1809 (N_1809,In_318,In_784);
and U1810 (N_1810,In_615,In_866);
or U1811 (N_1811,In_590,In_730);
nand U1812 (N_1812,In_450,In_577);
nand U1813 (N_1813,In_948,In_463);
xnor U1814 (N_1814,In_929,In_202);
or U1815 (N_1815,In_102,In_437);
nor U1816 (N_1816,In_575,In_657);
nand U1817 (N_1817,In_347,In_129);
nor U1818 (N_1818,In_867,In_388);
nand U1819 (N_1819,In_171,In_752);
nand U1820 (N_1820,In_617,In_600);
nor U1821 (N_1821,In_266,In_211);
nor U1822 (N_1822,In_348,In_557);
nor U1823 (N_1823,In_583,In_848);
and U1824 (N_1824,In_966,In_213);
nor U1825 (N_1825,In_429,In_634);
nor U1826 (N_1826,In_635,In_179);
nor U1827 (N_1827,In_155,In_574);
nand U1828 (N_1828,In_986,In_81);
nor U1829 (N_1829,In_514,In_228);
nor U1830 (N_1830,In_481,In_457);
and U1831 (N_1831,In_564,In_990);
and U1832 (N_1832,In_248,In_308);
nand U1833 (N_1833,In_103,In_32);
and U1834 (N_1834,In_897,In_983);
or U1835 (N_1835,In_277,In_548);
nor U1836 (N_1836,In_137,In_58);
nor U1837 (N_1837,In_789,In_486);
or U1838 (N_1838,In_338,In_403);
and U1839 (N_1839,In_639,In_637);
or U1840 (N_1840,In_822,In_800);
or U1841 (N_1841,In_703,In_468);
or U1842 (N_1842,In_421,In_91);
nand U1843 (N_1843,In_197,In_928);
nor U1844 (N_1844,In_561,In_815);
and U1845 (N_1845,In_686,In_291);
or U1846 (N_1846,In_963,In_441);
nor U1847 (N_1847,In_193,In_491);
or U1848 (N_1848,In_769,In_525);
or U1849 (N_1849,In_374,In_987);
nor U1850 (N_1850,In_247,In_701);
nand U1851 (N_1851,In_833,In_492);
and U1852 (N_1852,In_940,In_135);
and U1853 (N_1853,In_384,In_44);
nand U1854 (N_1854,In_567,In_719);
nand U1855 (N_1855,In_609,In_15);
and U1856 (N_1856,In_567,In_215);
and U1857 (N_1857,In_559,In_990);
or U1858 (N_1858,In_785,In_541);
xor U1859 (N_1859,In_717,In_317);
and U1860 (N_1860,In_168,In_203);
nor U1861 (N_1861,In_898,In_584);
nor U1862 (N_1862,In_408,In_722);
nand U1863 (N_1863,In_774,In_398);
nor U1864 (N_1864,In_914,In_194);
nor U1865 (N_1865,In_360,In_358);
or U1866 (N_1866,In_873,In_236);
nand U1867 (N_1867,In_217,In_698);
nand U1868 (N_1868,In_940,In_888);
nand U1869 (N_1869,In_520,In_653);
and U1870 (N_1870,In_471,In_712);
xnor U1871 (N_1871,In_982,In_476);
or U1872 (N_1872,In_508,In_358);
nand U1873 (N_1873,In_583,In_197);
and U1874 (N_1874,In_350,In_649);
nor U1875 (N_1875,In_861,In_864);
nor U1876 (N_1876,In_534,In_389);
nor U1877 (N_1877,In_999,In_131);
and U1878 (N_1878,In_369,In_2);
or U1879 (N_1879,In_290,In_52);
and U1880 (N_1880,In_324,In_941);
nor U1881 (N_1881,In_7,In_9);
or U1882 (N_1882,In_860,In_228);
and U1883 (N_1883,In_595,In_539);
nand U1884 (N_1884,In_766,In_44);
or U1885 (N_1885,In_438,In_97);
nand U1886 (N_1886,In_962,In_312);
xnor U1887 (N_1887,In_40,In_768);
or U1888 (N_1888,In_838,In_38);
nor U1889 (N_1889,In_222,In_517);
or U1890 (N_1890,In_518,In_534);
or U1891 (N_1891,In_774,In_408);
nor U1892 (N_1892,In_609,In_582);
or U1893 (N_1893,In_524,In_130);
or U1894 (N_1894,In_684,In_612);
nand U1895 (N_1895,In_497,In_287);
or U1896 (N_1896,In_410,In_607);
nand U1897 (N_1897,In_659,In_764);
nand U1898 (N_1898,In_842,In_343);
or U1899 (N_1899,In_260,In_703);
nand U1900 (N_1900,In_612,In_797);
nand U1901 (N_1901,In_733,In_935);
and U1902 (N_1902,In_733,In_555);
nor U1903 (N_1903,In_699,In_714);
or U1904 (N_1904,In_758,In_296);
or U1905 (N_1905,In_8,In_193);
and U1906 (N_1906,In_818,In_556);
nor U1907 (N_1907,In_724,In_868);
nand U1908 (N_1908,In_62,In_877);
nor U1909 (N_1909,In_347,In_375);
or U1910 (N_1910,In_496,In_425);
and U1911 (N_1911,In_140,In_950);
nand U1912 (N_1912,In_65,In_593);
and U1913 (N_1913,In_72,In_630);
or U1914 (N_1914,In_549,In_935);
nand U1915 (N_1915,In_60,In_58);
nor U1916 (N_1916,In_447,In_812);
or U1917 (N_1917,In_292,In_592);
nor U1918 (N_1918,In_334,In_907);
nor U1919 (N_1919,In_791,In_72);
or U1920 (N_1920,In_934,In_595);
nand U1921 (N_1921,In_105,In_766);
nor U1922 (N_1922,In_236,In_547);
or U1923 (N_1923,In_590,In_796);
nor U1924 (N_1924,In_745,In_391);
nor U1925 (N_1925,In_652,In_197);
nand U1926 (N_1926,In_910,In_740);
nand U1927 (N_1927,In_273,In_809);
or U1928 (N_1928,In_659,In_586);
and U1929 (N_1929,In_900,In_613);
and U1930 (N_1930,In_758,In_69);
or U1931 (N_1931,In_669,In_327);
and U1932 (N_1932,In_863,In_188);
and U1933 (N_1933,In_342,In_96);
and U1934 (N_1934,In_20,In_674);
nor U1935 (N_1935,In_443,In_834);
nand U1936 (N_1936,In_685,In_321);
or U1937 (N_1937,In_149,In_753);
nand U1938 (N_1938,In_199,In_497);
nor U1939 (N_1939,In_602,In_242);
nor U1940 (N_1940,In_913,In_429);
or U1941 (N_1941,In_37,In_832);
and U1942 (N_1942,In_501,In_972);
or U1943 (N_1943,In_454,In_571);
and U1944 (N_1944,In_444,In_419);
nor U1945 (N_1945,In_178,In_435);
or U1946 (N_1946,In_592,In_894);
or U1947 (N_1947,In_825,In_43);
and U1948 (N_1948,In_115,In_946);
nand U1949 (N_1949,In_768,In_351);
nand U1950 (N_1950,In_837,In_373);
nand U1951 (N_1951,In_71,In_854);
nand U1952 (N_1952,In_674,In_380);
nor U1953 (N_1953,In_634,In_448);
and U1954 (N_1954,In_371,In_129);
and U1955 (N_1955,In_266,In_177);
nor U1956 (N_1956,In_190,In_746);
and U1957 (N_1957,In_629,In_12);
nand U1958 (N_1958,In_500,In_665);
nand U1959 (N_1959,In_966,In_356);
nand U1960 (N_1960,In_314,In_873);
nand U1961 (N_1961,In_939,In_917);
or U1962 (N_1962,In_641,In_298);
or U1963 (N_1963,In_953,In_478);
nor U1964 (N_1964,In_671,In_191);
nor U1965 (N_1965,In_264,In_983);
or U1966 (N_1966,In_748,In_890);
or U1967 (N_1967,In_842,In_189);
nand U1968 (N_1968,In_330,In_93);
nand U1969 (N_1969,In_305,In_29);
nor U1970 (N_1970,In_3,In_910);
and U1971 (N_1971,In_898,In_23);
or U1972 (N_1972,In_694,In_294);
and U1973 (N_1973,In_259,In_358);
or U1974 (N_1974,In_468,In_140);
nand U1975 (N_1975,In_414,In_20);
nand U1976 (N_1976,In_776,In_81);
or U1977 (N_1977,In_142,In_893);
nor U1978 (N_1978,In_572,In_23);
and U1979 (N_1979,In_199,In_832);
nand U1980 (N_1980,In_752,In_543);
or U1981 (N_1981,In_555,In_334);
nand U1982 (N_1982,In_632,In_63);
nor U1983 (N_1983,In_349,In_946);
nand U1984 (N_1984,In_845,In_33);
nor U1985 (N_1985,In_307,In_547);
nand U1986 (N_1986,In_142,In_392);
nor U1987 (N_1987,In_228,In_194);
nand U1988 (N_1988,In_469,In_596);
nor U1989 (N_1989,In_880,In_416);
or U1990 (N_1990,In_798,In_836);
or U1991 (N_1991,In_217,In_761);
nor U1992 (N_1992,In_250,In_469);
nor U1993 (N_1993,In_630,In_452);
nor U1994 (N_1994,In_742,In_856);
nand U1995 (N_1995,In_366,In_330);
and U1996 (N_1996,In_486,In_127);
nand U1997 (N_1997,In_981,In_888);
or U1998 (N_1998,In_697,In_494);
nand U1999 (N_1999,In_334,In_319);
nor U2000 (N_2000,N_867,N_611);
or U2001 (N_2001,N_1796,N_1201);
or U2002 (N_2002,N_407,N_1671);
nor U2003 (N_2003,N_1681,N_1936);
or U2004 (N_2004,N_1085,N_314);
nand U2005 (N_2005,N_163,N_893);
nor U2006 (N_2006,N_1933,N_393);
or U2007 (N_2007,N_605,N_1321);
nand U2008 (N_2008,N_971,N_361);
nor U2009 (N_2009,N_500,N_1148);
nand U2010 (N_2010,N_995,N_984);
nand U2011 (N_2011,N_1239,N_1407);
nor U2012 (N_2012,N_733,N_1410);
nand U2013 (N_2013,N_1521,N_882);
or U2014 (N_2014,N_1856,N_1195);
nor U2015 (N_2015,N_531,N_746);
nand U2016 (N_2016,N_862,N_686);
nand U2017 (N_2017,N_217,N_1850);
or U2018 (N_2018,N_1534,N_1557);
nor U2019 (N_2019,N_1824,N_442);
nor U2020 (N_2020,N_320,N_175);
or U2021 (N_2021,N_1778,N_578);
and U2022 (N_2022,N_749,N_1795);
or U2023 (N_2023,N_69,N_1593);
nand U2024 (N_2024,N_515,N_929);
or U2025 (N_2025,N_728,N_813);
nand U2026 (N_2026,N_1971,N_1114);
nand U2027 (N_2027,N_732,N_927);
or U2028 (N_2028,N_181,N_276);
and U2029 (N_2029,N_1132,N_1399);
nor U2030 (N_2030,N_152,N_953);
nor U2031 (N_2031,N_1682,N_1319);
or U2032 (N_2032,N_891,N_1854);
xnor U2033 (N_2033,N_1324,N_1209);
nor U2034 (N_2034,N_1583,N_624);
and U2035 (N_2035,N_763,N_251);
or U2036 (N_2036,N_559,N_1898);
and U2037 (N_2037,N_1845,N_1490);
and U2038 (N_2038,N_794,N_873);
nand U2039 (N_2039,N_292,N_1269);
nand U2040 (N_2040,N_1282,N_1818);
nand U2041 (N_2041,N_94,N_297);
or U2042 (N_2042,N_1328,N_737);
or U2043 (N_2043,N_370,N_1683);
nand U2044 (N_2044,N_595,N_1147);
nand U2045 (N_2045,N_1296,N_1046);
nor U2046 (N_2046,N_1530,N_880);
or U2047 (N_2047,N_1851,N_59);
and U2048 (N_2048,N_1531,N_1591);
nor U2049 (N_2049,N_1720,N_1432);
nor U2050 (N_2050,N_757,N_1863);
nor U2051 (N_2051,N_114,N_825);
nor U2052 (N_2052,N_1464,N_702);
nor U2053 (N_2053,N_734,N_552);
nor U2054 (N_2054,N_1082,N_432);
nor U2055 (N_2055,N_1973,N_1672);
nor U2056 (N_2056,N_1451,N_863);
nor U2057 (N_2057,N_325,N_1077);
nand U2058 (N_2058,N_725,N_854);
or U2059 (N_2059,N_324,N_424);
or U2060 (N_2060,N_1317,N_1507);
nand U2061 (N_2061,N_601,N_530);
nand U2062 (N_2062,N_1520,N_1875);
or U2063 (N_2063,N_1900,N_1956);
nor U2064 (N_2064,N_437,N_745);
or U2065 (N_2065,N_1033,N_1295);
or U2066 (N_2066,N_486,N_1665);
nor U2067 (N_2067,N_538,N_980);
nor U2068 (N_2068,N_1895,N_1481);
nor U2069 (N_2069,N_1785,N_421);
or U2070 (N_2070,N_1897,N_289);
nand U2071 (N_2071,N_1752,N_456);
nor U2072 (N_2072,N_244,N_23);
and U2073 (N_2073,N_301,N_539);
nand U2074 (N_2074,N_1199,N_1709);
or U2075 (N_2075,N_1794,N_850);
or U2076 (N_2076,N_233,N_573);
nor U2077 (N_2077,N_579,N_21);
nor U2078 (N_2078,N_353,N_1646);
nand U2079 (N_2079,N_1375,N_985);
nand U2080 (N_2080,N_40,N_1702);
or U2081 (N_2081,N_1587,N_200);
nand U2082 (N_2082,N_489,N_748);
or U2083 (N_2083,N_920,N_731);
nand U2084 (N_2084,N_1453,N_379);
or U2085 (N_2085,N_1699,N_17);
or U2086 (N_2086,N_650,N_318);
nand U2087 (N_2087,N_380,N_693);
or U2088 (N_2088,N_1523,N_1804);
nand U2089 (N_2089,N_1142,N_1292);
xor U2090 (N_2090,N_1910,N_1013);
and U2091 (N_2091,N_1962,N_11);
nand U2092 (N_2092,N_1647,N_1967);
nand U2093 (N_2093,N_1164,N_1056);
and U2094 (N_2094,N_29,N_194);
nand U2095 (N_2095,N_1725,N_1345);
and U2096 (N_2096,N_1669,N_1303);
and U2097 (N_2097,N_1746,N_470);
and U2098 (N_2098,N_1182,N_1569);
and U2099 (N_2099,N_1940,N_857);
and U2100 (N_2100,N_1070,N_1457);
nand U2101 (N_2101,N_1981,N_1329);
nor U2102 (N_2102,N_336,N_1819);
and U2103 (N_2103,N_333,N_512);
and U2104 (N_2104,N_1073,N_1125);
and U2105 (N_2105,N_1828,N_34);
nand U2106 (N_2106,N_860,N_663);
nand U2107 (N_2107,N_1753,N_1734);
or U2108 (N_2108,N_1975,N_1458);
nor U2109 (N_2109,N_1678,N_309);
nor U2110 (N_2110,N_654,N_865);
nand U2111 (N_2111,N_1606,N_522);
nor U2112 (N_2112,N_323,N_1601);
nand U2113 (N_2113,N_188,N_1069);
or U2114 (N_2114,N_204,N_1730);
nor U2115 (N_2115,N_977,N_1740);
and U2116 (N_2116,N_20,N_1468);
or U2117 (N_2117,N_754,N_1389);
nor U2118 (N_2118,N_645,N_1318);
nor U2119 (N_2119,N_675,N_1728);
or U2120 (N_2120,N_394,N_1543);
or U2121 (N_2121,N_1486,N_43);
nor U2122 (N_2122,N_1123,N_229);
nand U2123 (N_2123,N_1765,N_1308);
and U2124 (N_2124,N_30,N_1629);
or U2125 (N_2125,N_682,N_1197);
nand U2126 (N_2126,N_1772,N_206);
and U2127 (N_2127,N_1686,N_1846);
and U2128 (N_2128,N_847,N_1739);
nor U2129 (N_2129,N_1304,N_1838);
nand U2130 (N_2130,N_1844,N_1149);
and U2131 (N_2131,N_1718,N_1234);
nand U2132 (N_2132,N_1146,N_1660);
nand U2133 (N_2133,N_429,N_1040);
and U2134 (N_2134,N_1829,N_1834);
nor U2135 (N_2135,N_439,N_507);
nand U2136 (N_2136,N_373,N_1045);
nand U2137 (N_2137,N_717,N_153);
and U2138 (N_2138,N_593,N_788);
and U2139 (N_2139,N_1293,N_449);
nand U2140 (N_2140,N_419,N_1948);
nor U2141 (N_2141,N_955,N_348);
or U2142 (N_2142,N_649,N_237);
nor U2143 (N_2143,N_298,N_287);
and U2144 (N_2144,N_1731,N_1110);
nor U2145 (N_2145,N_1256,N_716);
and U2146 (N_2146,N_304,N_1397);
nor U2147 (N_2147,N_1913,N_327);
nand U2148 (N_2148,N_1541,N_1249);
or U2149 (N_2149,N_1398,N_869);
and U2150 (N_2150,N_1489,N_602);
nand U2151 (N_2151,N_433,N_1836);
and U2152 (N_2152,N_1855,N_303);
nor U2153 (N_2153,N_1789,N_1221);
and U2154 (N_2154,N_1525,N_886);
and U2155 (N_2155,N_1265,N_1770);
and U2156 (N_2156,N_644,N_768);
or U2157 (N_2157,N_25,N_619);
nor U2158 (N_2158,N_32,N_1208);
nor U2159 (N_2159,N_575,N_1762);
or U2160 (N_2160,N_1381,N_387);
nor U2161 (N_2161,N_685,N_554);
or U2162 (N_2162,N_1416,N_260);
and U2163 (N_2163,N_646,N_473);
or U2164 (N_2164,N_553,N_1330);
or U2165 (N_2165,N_1176,N_1130);
nor U2166 (N_2166,N_1350,N_134);
nor U2167 (N_2167,N_1411,N_691);
and U2168 (N_2168,N_1966,N_284);
nor U2169 (N_2169,N_250,N_979);
nand U2170 (N_2170,N_293,N_1471);
or U2171 (N_2171,N_176,N_1436);
nor U2172 (N_2172,N_279,N_1021);
and U2173 (N_2173,N_1782,N_1885);
nand U2174 (N_2174,N_1611,N_747);
nor U2175 (N_2175,N_372,N_1032);
or U2176 (N_2176,N_1815,N_1947);
nand U2177 (N_2177,N_281,N_1786);
or U2178 (N_2178,N_377,N_463);
and U2179 (N_2179,N_275,N_819);
or U2180 (N_2180,N_981,N_990);
and U2181 (N_2181,N_1367,N_249);
and U2182 (N_2182,N_1577,N_368);
nand U2183 (N_2183,N_1989,N_992);
and U2184 (N_2184,N_885,N_54);
or U2185 (N_2185,N_881,N_1874);
or U2186 (N_2186,N_1093,N_1335);
nor U2187 (N_2187,N_1676,N_1509);
nand U2188 (N_2188,N_861,N_1492);
nand U2189 (N_2189,N_1325,N_1217);
nand U2190 (N_2190,N_896,N_1987);
nand U2191 (N_2191,N_1347,N_1086);
or U2192 (N_2192,N_1310,N_1336);
xnor U2193 (N_2193,N_1639,N_501);
nand U2194 (N_2194,N_228,N_1722);
or U2195 (N_2195,N_1424,N_1442);
or U2196 (N_2196,N_1379,N_256);
or U2197 (N_2197,N_680,N_332);
or U2198 (N_2198,N_606,N_1403);
and U2199 (N_2199,N_116,N_90);
or U2200 (N_2200,N_169,N_1995);
and U2201 (N_2201,N_1764,N_1480);
or U2202 (N_2202,N_317,N_77);
nor U2203 (N_2203,N_369,N_668);
nand U2204 (N_2204,N_105,N_678);
and U2205 (N_2205,N_1476,N_420);
nand U2206 (N_2206,N_1316,N_1886);
nor U2207 (N_2207,N_855,N_1359);
nand U2208 (N_2208,N_1128,N_753);
and U2209 (N_2209,N_8,N_366);
xnor U2210 (N_2210,N_1161,N_14);
nor U2211 (N_2211,N_799,N_83);
nand U2212 (N_2212,N_465,N_1503);
nand U2213 (N_2213,N_329,N_991);
nor U2214 (N_2214,N_612,N_817);
or U2215 (N_2215,N_779,N_1267);
nor U2216 (N_2216,N_359,N_1615);
or U2217 (N_2217,N_933,N_1004);
nand U2218 (N_2218,N_1435,N_681);
and U2219 (N_2219,N_986,N_1779);
and U2220 (N_2220,N_1165,N_1969);
nor U2221 (N_2221,N_1723,N_494);
and U2222 (N_2222,N_1858,N_598);
nand U2223 (N_2223,N_1354,N_1092);
or U2224 (N_2224,N_884,N_1276);
and U2225 (N_2225,N_1438,N_1690);
and U2226 (N_2226,N_1988,N_160);
or U2227 (N_2227,N_1036,N_919);
nor U2228 (N_2228,N_1558,N_775);
nand U2229 (N_2229,N_60,N_834);
and U2230 (N_2230,N_555,N_1384);
and U2231 (N_2231,N_1198,N_410);
or U2232 (N_2232,N_852,N_180);
xor U2233 (N_2233,N_776,N_1444);
or U2234 (N_2234,N_1250,N_750);
nand U2235 (N_2235,N_1602,N_613);
nor U2236 (N_2236,N_328,N_130);
nand U2237 (N_2237,N_1679,N_1302);
or U2238 (N_2238,N_1642,N_947);
nor U2239 (N_2239,N_1423,N_1826);
nor U2240 (N_2240,N_958,N_1320);
xor U2241 (N_2241,N_864,N_1160);
and U2242 (N_2242,N_626,N_1155);
nor U2243 (N_2243,N_563,N_633);
or U2244 (N_2244,N_313,N_434);
nand U2245 (N_2245,N_349,N_707);
nor U2246 (N_2246,N_1698,N_1305);
or U2247 (N_2247,N_155,N_1658);
or U2248 (N_2248,N_1213,N_1088);
or U2249 (N_2249,N_178,N_803);
or U2250 (N_2250,N_1907,N_634);
nor U2251 (N_2251,N_1264,N_1651);
and U2252 (N_2252,N_1491,N_1545);
nand U2253 (N_2253,N_1878,N_1691);
nand U2254 (N_2254,N_37,N_1645);
nand U2255 (N_2255,N_641,N_1225);
or U2256 (N_2256,N_1798,N_1235);
nor U2257 (N_2257,N_826,N_1505);
nor U2258 (N_2258,N_1284,N_1964);
nand U2259 (N_2259,N_1514,N_1382);
and U2260 (N_2260,N_647,N_1697);
and U2261 (N_2261,N_1127,N_1958);
nand U2262 (N_2262,N_55,N_1478);
nor U2263 (N_2263,N_263,N_1763);
nor U2264 (N_2264,N_1871,N_714);
nand U2265 (N_2265,N_1749,N_950);
nand U2266 (N_2266,N_976,N_27);
nand U2267 (N_2267,N_1797,N_1167);
or U2268 (N_2268,N_959,N_875);
nand U2269 (N_2269,N_252,N_78);
or U2270 (N_2270,N_1882,N_632);
nand U2271 (N_2271,N_1346,N_341);
or U2272 (N_2272,N_84,N_96);
nor U2273 (N_2273,N_255,N_389);
or U2274 (N_2274,N_112,N_792);
or U2275 (N_2275,N_1504,N_1605);
or U2276 (N_2276,N_1528,N_793);
or U2277 (N_2277,N_1810,N_1341);
nand U2278 (N_2278,N_1238,N_1242);
and U2279 (N_2279,N_1835,N_877);
nand U2280 (N_2280,N_1641,N_1777);
nand U2281 (N_2281,N_743,N_557);
nand U2282 (N_2282,N_1332,N_1972);
or U2283 (N_2283,N_1,N_49);
and U2284 (N_2284,N_1542,N_1050);
and U2285 (N_2285,N_242,N_836);
and U2286 (N_2286,N_905,N_898);
nor U2287 (N_2287,N_513,N_1982);
and U2288 (N_2288,N_761,N_1771);
or U2289 (N_2289,N_853,N_708);
and U2290 (N_2290,N_787,N_1735);
and U2291 (N_2291,N_452,N_1930);
nand U2292 (N_2292,N_608,N_1437);
or U2293 (N_2293,N_273,N_168);
nand U2294 (N_2294,N_558,N_1729);
nor U2295 (N_2295,N_345,N_784);
and U2296 (N_2296,N_1358,N_1757);
and U2297 (N_2297,N_1994,N_944);
and U2298 (N_2298,N_1756,N_1568);
or U2299 (N_2299,N_1944,N_1051);
and U2300 (N_2300,N_381,N_5);
and U2301 (N_2301,N_690,N_1852);
nor U2302 (N_2302,N_179,N_683);
nor U2303 (N_2303,N_1783,N_1177);
nor U2304 (N_2304,N_1570,N_783);
nand U2305 (N_2305,N_240,N_856);
nand U2306 (N_2306,N_639,N_245);
nand U2307 (N_2307,N_804,N_1376);
and U2308 (N_2308,N_1390,N_677);
xor U2309 (N_2309,N_1353,N_1290);
and U2310 (N_2310,N_268,N_1371);
nand U2311 (N_2311,N_1552,N_1278);
and U2312 (N_2312,N_514,N_1527);
xnor U2313 (N_2313,N_1113,N_189);
or U2314 (N_2314,N_523,N_148);
or U2315 (N_2315,N_1117,N_495);
and U2316 (N_2316,N_1080,N_1063);
and U2317 (N_2317,N_36,N_1842);
or U2318 (N_2318,N_1083,N_1768);
and U2319 (N_2319,N_830,N_1145);
or U2320 (N_2320,N_1924,N_1079);
or U2321 (N_2321,N_661,N_1750);
nor U2322 (N_2322,N_1011,N_1825);
and U2323 (N_2323,N_1044,N_1331);
and U2324 (N_2324,N_1386,N_1538);
nor U2325 (N_2325,N_1474,N_1151);
nor U2326 (N_2326,N_1584,N_1169);
and U2327 (N_2327,N_906,N_1214);
or U2328 (N_2328,N_700,N_1236);
and U2329 (N_2329,N_902,N_527);
or U2330 (N_2330,N_1904,N_588);
nor U2331 (N_2331,N_136,N_1456);
nor U2332 (N_2332,N_1294,N_1617);
and U2333 (N_2333,N_1189,N_1881);
or U2334 (N_2334,N_350,N_174);
nor U2335 (N_2335,N_948,N_1993);
or U2336 (N_2336,N_2,N_1065);
or U2337 (N_2337,N_729,N_1159);
nand U2338 (N_2338,N_1685,N_1263);
nand U2339 (N_2339,N_208,N_1551);
or U2340 (N_2340,N_1806,N_635);
or U2341 (N_2341,N_202,N_759);
nand U2342 (N_2342,N_1449,N_1612);
and U2343 (N_2343,N_128,N_1596);
or U2344 (N_2344,N_1941,N_1048);
and U2345 (N_2345,N_1550,N_648);
nand U2346 (N_2346,N_762,N_1738);
or U2347 (N_2347,N_42,N_1823);
or U2348 (N_2348,N_1932,N_492);
and U2349 (N_2349,N_147,N_1546);
and U2350 (N_2350,N_1893,N_664);
or U2351 (N_2351,N_1207,N_482);
and U2352 (N_2352,N_19,N_968);
nand U2353 (N_2353,N_257,N_103);
and U2354 (N_2354,N_278,N_506);
nand U2355 (N_2355,N_963,N_1905);
and U2356 (N_2356,N_1368,N_1119);
and U2357 (N_2357,N_85,N_1656);
or U2358 (N_2358,N_485,N_858);
nand U2359 (N_2359,N_541,N_978);
nor U2360 (N_2360,N_232,N_755);
and U2361 (N_2361,N_213,N_455);
or U2362 (N_2362,N_674,N_1495);
nand U2363 (N_2363,N_265,N_1780);
nor U2364 (N_2364,N_1903,N_1576);
and U2365 (N_2365,N_346,N_1865);
and U2366 (N_2366,N_1630,N_365);
nor U2367 (N_2367,N_907,N_534);
nand U2368 (N_2368,N_508,N_190);
xor U2369 (N_2369,N_1134,N_1868);
nor U2370 (N_2370,N_119,N_1517);
nand U2371 (N_2371,N_1340,N_720);
nand U2372 (N_2372,N_1053,N_931);
nand U2373 (N_2373,N_414,N_580);
and U2374 (N_2374,N_1003,N_1422);
or U2375 (N_2375,N_1120,N_1872);
nor U2376 (N_2376,N_171,N_71);
or U2377 (N_2377,N_436,N_165);
nor U2378 (N_2378,N_721,N_1742);
nand U2379 (N_2379,N_666,N_1673);
nand U2380 (N_2380,N_384,N_216);
nand U2381 (N_2381,N_302,N_1440);
or U2382 (N_2382,N_167,N_1559);
nor U2383 (N_2383,N_827,N_1488);
or U2384 (N_2384,N_1864,N_1532);
and U2385 (N_2385,N_604,N_548);
or U2386 (N_2386,N_493,N_688);
or U2387 (N_2387,N_1508,N_1255);
nand U2388 (N_2388,N_141,N_773);
nor U2389 (N_2389,N_343,N_88);
nand U2390 (N_2390,N_658,N_1467);
nand U2391 (N_2391,N_1412,N_1019);
or U2392 (N_2392,N_1748,N_1482);
or U2393 (N_2393,N_1101,N_1613);
nand U2394 (N_2394,N_848,N_1413);
nor U2395 (N_2395,N_1622,N_1774);
nor U2396 (N_2396,N_478,N_1377);
and U2397 (N_2397,N_1228,N_807);
nand U2398 (N_2398,N_1866,N_993);
or U2399 (N_2399,N_1983,N_1433);
nand U2400 (N_2400,N_1405,N_1816);
nand U2401 (N_2401,N_1166,N_1094);
and U2402 (N_2402,N_1938,N_477);
nand U2403 (N_2403,N_106,N_93);
or U2404 (N_2404,N_1415,N_375);
nand U2405 (N_2405,N_777,N_1873);
nor U2406 (N_2406,N_1091,N_1054);
nand U2407 (N_2407,N_1364,N_1574);
or U2408 (N_2408,N_435,N_226);
and U2409 (N_2409,N_614,N_1219);
or U2410 (N_2410,N_295,N_1581);
or U2411 (N_2411,N_568,N_1644);
nor U2412 (N_2412,N_464,N_797);
or U2413 (N_2413,N_1733,N_184);
nor U2414 (N_2414,N_209,N_73);
or U2415 (N_2415,N_271,N_417);
xnor U2416 (N_2416,N_207,N_79);
nor U2417 (N_2417,N_1803,N_1867);
or U2418 (N_2418,N_1706,N_1300);
or U2419 (N_2419,N_1713,N_684);
or U2420 (N_2420,N_544,N_294);
or U2421 (N_2421,N_735,N_44);
nand U2422 (N_2422,N_1190,N_550);
and U2423 (N_2423,N_592,N_914);
or U2424 (N_2424,N_1144,N_1957);
nor U2425 (N_2425,N_1839,N_1102);
nor U2426 (N_2426,N_1515,N_490);
nand U2427 (N_2427,N_599,N_1425);
and U2428 (N_2428,N_358,N_97);
and U2429 (N_2429,N_1025,N_1977);
nor U2430 (N_2430,N_1877,N_1240);
and U2431 (N_2431,N_291,N_1418);
nand U2432 (N_2432,N_1181,N_1378);
or U2433 (N_2433,N_1916,N_91);
and U2434 (N_2434,N_802,N_62);
and U2435 (N_2435,N_1883,N_203);
nand U2436 (N_2436,N_1920,N_930);
or U2437 (N_2437,N_1277,N_765);
and U2438 (N_2438,N_1628,N_998);
and U2439 (N_2439,N_832,N_1247);
or U2440 (N_2440,N_566,N_1979);
or U2441 (N_2441,N_1887,N_1754);
nand U2442 (N_2442,N_1500,N_1042);
or U2443 (N_2443,N_1890,N_440);
or U2444 (N_2444,N_1743,N_438);
and U2445 (N_2445,N_1652,N_225);
or U2446 (N_2446,N_589,N_925);
nor U2447 (N_2447,N_154,N_1588);
nor U2448 (N_2448,N_4,N_1674);
and U2449 (N_2449,N_471,N_461);
nor U2450 (N_2450,N_1573,N_876);
and U2451 (N_2451,N_220,N_342);
nor U2452 (N_2452,N_334,N_1648);
nand U2453 (N_2453,N_1485,N_1253);
nand U2454 (N_2454,N_1792,N_1626);
and U2455 (N_2455,N_1775,N_1275);
nor U2456 (N_2456,N_509,N_1349);
or U2457 (N_2457,N_1633,N_1103);
or U2458 (N_2458,N_1472,N_1635);
or U2459 (N_2459,N_1790,N_1459);
nor U2460 (N_2460,N_529,N_1880);
and U2461 (N_2461,N_1465,N_431);
or U2462 (N_2462,N_1516,N_138);
or U2463 (N_2463,N_1714,N_1272);
or U2464 (N_2464,N_866,N_1005);
or U2465 (N_2465,N_1108,N_1539);
nor U2466 (N_2466,N_331,N_1787);
or U2467 (N_2467,N_789,N_1607);
and U2468 (N_2468,N_888,N_1519);
and U2469 (N_2469,N_1809,N_625);
nor U2470 (N_2470,N_427,N_670);
nand U2471 (N_2471,N_874,N_806);
and U2472 (N_2472,N_395,N_542);
nand U2473 (N_2473,N_617,N_1443);
nor U2474 (N_2474,N_1374,N_1799);
or U2475 (N_2475,N_1529,N_1627);
nand U2476 (N_2476,N_701,N_423);
nor U2477 (N_2477,N_1580,N_1156);
nor U2478 (N_2478,N_1758,N_1248);
nor U2479 (N_2479,N_782,N_815);
or U2480 (N_2480,N_227,N_1097);
nand U2481 (N_2481,N_1100,N_1227);
nand U2482 (N_2482,N_808,N_1695);
and U2483 (N_2483,N_752,N_897);
nand U2484 (N_2484,N_1241,N_591);
or U2485 (N_2485,N_1366,N_310);
or U2486 (N_2486,N_185,N_1137);
nor U2487 (N_2487,N_472,N_526);
nand U2488 (N_2488,N_1163,N_1109);
nor U2489 (N_2489,N_1892,N_703);
and U2490 (N_2490,N_1649,N_972);
nand U2491 (N_2491,N_191,N_1662);
and U2492 (N_2492,N_31,N_47);
nand U2493 (N_2493,N_1037,N_1192);
or U2494 (N_2494,N_126,N_1355);
nand U2495 (N_2495,N_665,N_911);
nand U2496 (N_2496,N_1943,N_231);
or U2497 (N_2497,N_951,N_1406);
nor U2498 (N_2498,N_1847,N_6);
or U2499 (N_2499,N_822,N_296);
nor U2500 (N_2500,N_600,N_210);
or U2501 (N_2501,N_937,N_1902);
nand U2502 (N_2502,N_547,N_535);
nand U2503 (N_2503,N_406,N_1041);
nor U2504 (N_2504,N_790,N_1620);
and U2505 (N_2505,N_16,N_308);
nand U2506 (N_2506,N_151,N_164);
nand U2507 (N_2507,N_451,N_1830);
nor U2508 (N_2508,N_1285,N_1929);
xor U2509 (N_2509,N_890,N_767);
nor U2510 (N_2510,N_1499,N_50);
or U2511 (N_2511,N_710,N_704);
or U2512 (N_2512,N_476,N_1154);
nand U2513 (N_2513,N_1064,N_1362);
nor U2514 (N_2514,N_1894,N_934);
nor U2515 (N_2515,N_1935,N_1876);
nand U2516 (N_2516,N_1487,N_1429);
and U2517 (N_2517,N_214,N_1394);
nor U2518 (N_2518,N_1891,N_1965);
or U2519 (N_2519,N_1271,N_46);
nor U2520 (N_2520,N_1595,N_413);
or U2521 (N_2521,N_469,N_1210);
nand U2522 (N_2522,N_371,N_1215);
or U2523 (N_2523,N_1726,N_1946);
nand U2524 (N_2524,N_1206,N_567);
nor U2525 (N_2525,N_1513,N_936);
and U2526 (N_2526,N_525,N_1901);
or U2527 (N_2527,N_1002,N_1518);
nand U2528 (N_2528,N_1126,N_1802);
nor U2529 (N_2529,N_620,N_468);
or U2530 (N_2530,N_1172,N_238);
and U2531 (N_2531,N_1822,N_1879);
or U2532 (N_2532,N_1419,N_1357);
or U2533 (N_2533,N_157,N_1661);
and U2534 (N_2534,N_248,N_290);
nand U2535 (N_2535,N_669,N_528);
xor U2536 (N_2536,N_277,N_1344);
or U2537 (N_2537,N_967,N_652);
nand U2538 (N_2538,N_1018,N_1095);
and U2539 (N_2539,N_340,N_243);
or U2540 (N_2540,N_1060,N_68);
nand U2541 (N_2541,N_1252,N_1506);
and U2542 (N_2542,N_183,N_520);
nor U2543 (N_2543,N_846,N_1369);
and U2544 (N_2544,N_166,N_1084);
or U2545 (N_2545,N_1712,N_193);
and U2546 (N_2546,N_221,N_475);
or U2547 (N_2547,N_1254,N_1625);
or U2548 (N_2548,N_1719,N_1000);
nor U2549 (N_2549,N_1494,N_12);
nand U2550 (N_2550,N_628,N_1643);
and U2551 (N_2551,N_479,N_386);
nand U2552 (N_2552,N_61,N_1703);
nor U2553 (N_2553,N_1684,N_718);
nand U2554 (N_2554,N_1736,N_399);
nand U2555 (N_2555,N_1111,N_1640);
and U2556 (N_2556,N_1135,N_133);
nand U2557 (N_2557,N_1047,N_344);
or U2558 (N_2558,N_355,N_781);
nor U2559 (N_2559,N_1554,N_1062);
nand U2560 (N_2560,N_1006,N_339);
or U2561 (N_2561,N_1140,N_946);
or U2562 (N_2562,N_1755,N_1667);
nor U2563 (N_2563,N_1348,N_1751);
nor U2564 (N_2564,N_576,N_698);
nor U2565 (N_2565,N_1998,N_1270);
nand U2566 (N_2566,N_964,N_676);
nor U2567 (N_2567,N_1180,N_135);
xor U2568 (N_2568,N_1727,N_923);
nor U2569 (N_2569,N_1031,N_140);
xnor U2570 (N_2570,N_81,N_1841);
or U2571 (N_2571,N_247,N_659);
and U2572 (N_2572,N_1664,N_623);
and U2573 (N_2573,N_319,N_1937);
nor U2574 (N_2574,N_142,N_660);
nand U2575 (N_2575,N_657,N_1857);
nand U2576 (N_2576,N_1365,N_653);
or U2577 (N_2577,N_1016,N_1578);
and U2578 (N_2578,N_418,N_246);
nor U2579 (N_2579,N_945,N_1884);
nor U2580 (N_2580,N_1540,N_581);
or U2581 (N_2581,N_796,N_1363);
and U2582 (N_2582,N_1312,N_307);
and U2583 (N_2583,N_627,N_1980);
or U2584 (N_2584,N_337,N_392);
nor U2585 (N_2585,N_98,N_272);
nand U2586 (N_2586,N_1848,N_584);
and U2587 (N_2587,N_280,N_441);
xnor U2588 (N_2588,N_844,N_335);
or U2589 (N_2589,N_195,N_1408);
nor U2590 (N_2590,N_139,N_491);
and U2591 (N_2591,N_1136,N_1393);
or U2592 (N_2592,N_1402,N_1059);
and U2593 (N_2593,N_364,N_158);
and U2594 (N_2594,N_398,N_949);
nor U2595 (N_2595,N_1970,N_125);
and U2596 (N_2596,N_109,N_1636);
and U2597 (N_2597,N_887,N_480);
and U2598 (N_2598,N_1637,N_1445);
nor U2599 (N_2599,N_1955,N_1071);
nand U2600 (N_2600,N_1414,N_656);
nor U2601 (N_2601,N_1484,N_1566);
nand U2602 (N_2602,N_1522,N_935);
and U2603 (N_2603,N_1567,N_771);
and U2604 (N_2604,N_800,N_1976);
and U2605 (N_2605,N_488,N_1562);
nand U2606 (N_2606,N_1609,N_378);
or U2607 (N_2607,N_895,N_1261);
nand U2608 (N_2608,N_1619,N_253);
nand U2609 (N_2609,N_1614,N_1066);
nand U2610 (N_2610,N_230,N_1853);
or U2611 (N_2611,N_1537,N_182);
nor U2612 (N_2612,N_1216,N_1396);
nor U2613 (N_2613,N_838,N_1171);
or U2614 (N_2614,N_1237,N_1618);
and U2615 (N_2615,N_1928,N_1732);
nand U2616 (N_2616,N_982,N_453);
or U2617 (N_2617,N_1385,N_1991);
nor U2618 (N_2618,N_258,N_39);
xnor U2619 (N_2619,N_1087,N_1222);
nand U2620 (N_2620,N_562,N_121);
and U2621 (N_2621,N_474,N_1279);
or U2622 (N_2622,N_1211,N_288);
or U2623 (N_2623,N_1862,N_299);
or U2624 (N_2624,N_1843,N_0);
nor U2625 (N_2625,N_1820,N_415);
nor U2626 (N_2626,N_996,N_939);
or U2627 (N_2627,N_1483,N_1832);
nand U2628 (N_2628,N_26,N_57);
nor U2629 (N_2629,N_1544,N_1565);
and U2630 (N_2630,N_1224,N_564);
nand U2631 (N_2631,N_67,N_689);
nor U2632 (N_2632,N_1352,N_894);
or U2633 (N_2633,N_818,N_388);
or U2634 (N_2634,N_814,N_1373);
nor U2635 (N_2635,N_1974,N_828);
or U2636 (N_2636,N_1283,N_1417);
or U2637 (N_2637,N_74,N_259);
and U2638 (N_2638,N_396,N_1431);
and U2639 (N_2639,N_1921,N_261);
or U2640 (N_2640,N_1800,N_1395);
nand U2641 (N_2641,N_1131,N_1592);
nand U2642 (N_2642,N_1788,N_687);
nor U2643 (N_2643,N_1724,N_918);
and U2644 (N_2644,N_1138,N_610);
nand U2645 (N_2645,N_401,N_1984);
nand U2646 (N_2646,N_713,N_811);
nand U2647 (N_2647,N_1273,N_837);
nand U2648 (N_2648,N_3,N_1428);
or U2649 (N_2649,N_1585,N_86);
nor U2650 (N_2650,N_374,N_1589);
nor U2651 (N_2651,N_1188,N_1343);
nor U2652 (N_2652,N_405,N_821);
and U2653 (N_2653,N_409,N_1462);
and U2654 (N_2654,N_999,N_594);
and U2655 (N_2655,N_723,N_1143);
nor U2656 (N_2656,N_1670,N_615);
nor U2657 (N_2657,N_1711,N_1693);
or U2658 (N_2658,N_1229,N_487);
and U2659 (N_2659,N_1708,N_1663);
nand U2660 (N_2660,N_1502,N_322);
or U2661 (N_2661,N_1288,N_1315);
or U2662 (N_2662,N_502,N_397);
or U2663 (N_2663,N_33,N_812);
nor U2664 (N_2664,N_1590,N_940);
nand U2665 (N_2665,N_908,N_1023);
nor U2666 (N_2666,N_536,N_1960);
or U2667 (N_2667,N_1680,N_45);
and U2668 (N_2668,N_1870,N_1990);
and U2669 (N_2669,N_1466,N_1942);
nor U2670 (N_2670,N_1454,N_1582);
or U2671 (N_2671,N_1203,N_1026);
nand U2672 (N_2672,N_58,N_505);
nor U2673 (N_2673,N_1654,N_1479);
and U2674 (N_2674,N_621,N_1388);
and U2675 (N_2675,N_1931,N_201);
or U2676 (N_2676,N_1536,N_1017);
or U2677 (N_2677,N_922,N_1153);
and U2678 (N_2678,N_403,N_809);
nor U2679 (N_2679,N_145,N_351);
nor U2680 (N_2680,N_957,N_1963);
or U2681 (N_2681,N_454,N_1115);
xor U2682 (N_2682,N_1631,N_1533);
nor U2683 (N_2683,N_1380,N_738);
or U2684 (N_2684,N_1696,N_840);
nand U2685 (N_2685,N_1773,N_111);
or U2686 (N_2686,N_450,N_820);
nor U2687 (N_2687,N_124,N_1204);
or U2688 (N_2688,N_1477,N_1391);
and U2689 (N_2689,N_1030,N_1561);
and U2690 (N_2690,N_1556,N_1688);
nand U2691 (N_2691,N_697,N_1677);
or U2692 (N_2692,N_122,N_1027);
nor U2693 (N_2693,N_943,N_651);
or U2694 (N_2694,N_643,N_15);
nor U2695 (N_2695,N_1007,N_871);
and U2696 (N_2696,N_239,N_889);
nand U2697 (N_2697,N_1555,N_915);
or U2698 (N_2698,N_1896,N_842);
nor U2699 (N_2699,N_107,N_13);
or U2700 (N_2700,N_1737,N_1849);
nand U2701 (N_2701,N_1721,N_1401);
and U2702 (N_2702,N_1058,N_1926);
nand U2703 (N_2703,N_774,N_1889);
nand U2704 (N_2704,N_267,N_460);
nand U2705 (N_2705,N_1173,N_618);
xnor U2706 (N_2706,N_311,N_1266);
or U2707 (N_2707,N_131,N_1497);
nand U2708 (N_2708,N_662,N_1511);
nand U2709 (N_2709,N_1572,N_1187);
and U2710 (N_2710,N_66,N_845);
nor U2711 (N_2711,N_516,N_1009);
or U2712 (N_2712,N_583,N_1427);
and U2713 (N_2713,N_1246,N_462);
and U2714 (N_2714,N_1333,N_510);
or U2715 (N_2715,N_574,N_1473);
or U2716 (N_2716,N_315,N_1212);
or U2717 (N_2717,N_1493,N_1911);
or U2718 (N_2718,N_1231,N_569);
and U2719 (N_2719,N_1243,N_823);
nand U2720 (N_2720,N_543,N_285);
nand U2721 (N_2721,N_363,N_511);
and U2722 (N_2722,N_1997,N_444);
and U2723 (N_2723,N_1370,N_282);
nand U2724 (N_2724,N_1840,N_408);
or U2725 (N_2725,N_571,N_269);
or U2726 (N_2726,N_1194,N_1951);
or U2727 (N_2727,N_667,N_952);
nand U2728 (N_2728,N_80,N_1869);
xnor U2729 (N_2729,N_904,N_402);
and U2730 (N_2730,N_1139,N_362);
or U2731 (N_2731,N_1262,N_1233);
or U2732 (N_2732,N_1121,N_1659);
or U2733 (N_2733,N_1434,N_1978);
nor U2734 (N_2734,N_1043,N_1028);
or U2735 (N_2735,N_924,N_637);
or U2736 (N_2736,N_810,N_422);
or U2737 (N_2737,N_942,N_696);
nand U2738 (N_2738,N_622,N_1311);
or U2739 (N_2739,N_1888,N_695);
and U2740 (N_2740,N_1553,N_1986);
nor U2741 (N_2741,N_1289,N_642);
or U2742 (N_2742,N_70,N_1745);
or U2743 (N_2743,N_521,N_772);
nand U2744 (N_2744,N_916,N_1461);
or U2745 (N_2745,N_1859,N_448);
or U2746 (N_2746,N_1174,N_577);
nor U2747 (N_2747,N_549,N_970);
nand U2748 (N_2748,N_903,N_300);
nor U2749 (N_2749,N_51,N_1925);
nand U2750 (N_2750,N_560,N_1666);
or U2751 (N_2751,N_144,N_426);
and U2752 (N_2752,N_1298,N_1950);
nand U2753 (N_2753,N_1096,N_503);
or U2754 (N_2754,N_1548,N_205);
or U2755 (N_2755,N_416,N_899);
nand U2756 (N_2756,N_376,N_445);
nand U2757 (N_2757,N_254,N_1001);
or U2758 (N_2758,N_938,N_961);
xor U2759 (N_2759,N_1291,N_1081);
nand U2760 (N_2760,N_312,N_1074);
nor U2761 (N_2761,N_1535,N_672);
or U2762 (N_2762,N_1624,N_1334);
nor U2763 (N_2763,N_187,N_824);
or U2764 (N_2764,N_484,N_1949);
or U2765 (N_2765,N_222,N_1934);
and U2766 (N_2766,N_1475,N_1860);
or U2767 (N_2767,N_616,N_412);
or U2768 (N_2768,N_7,N_962);
and U2769 (N_2769,N_570,N_400);
or U2770 (N_2770,N_590,N_1057);
nand U2771 (N_2771,N_357,N_1232);
or U2772 (N_2772,N_878,N_1668);
nor U2773 (N_2773,N_517,N_1811);
and U2774 (N_2774,N_211,N_726);
nor U2775 (N_2775,N_1014,N_829);
nor U2776 (N_2776,N_117,N_705);
and U2777 (N_2777,N_123,N_1498);
nor U2778 (N_2778,N_18,N_954);
or U2779 (N_2779,N_1309,N_1704);
nand U2780 (N_2780,N_586,N_928);
nand U2781 (N_2781,N_496,N_631);
and U2782 (N_2782,N_22,N_102);
and U2783 (N_2783,N_430,N_1603);
and U2784 (N_2784,N_1769,N_997);
nand U2785 (N_2785,N_1687,N_63);
xor U2786 (N_2786,N_1638,N_988);
or U2787 (N_2787,N_540,N_1791);
nor U2788 (N_2788,N_41,N_1906);
or U2789 (N_2789,N_709,N_1078);
nor U2790 (N_2790,N_270,N_872);
nor U2791 (N_2791,N_1157,N_572);
and U2792 (N_2792,N_1061,N_1226);
nand U2793 (N_2793,N_912,N_921);
or U2794 (N_2794,N_177,N_1692);
nand U2795 (N_2795,N_306,N_1075);
nor U2796 (N_2796,N_913,N_994);
nand U2797 (N_2797,N_197,N_1701);
and U2798 (N_2798,N_1599,N_831);
nor U2799 (N_2799,N_795,N_638);
and U2800 (N_2800,N_1833,N_497);
or U2801 (N_2801,N_1917,N_1813);
and U2802 (N_2802,N_1179,N_1259);
nand U2803 (N_2803,N_966,N_715);
or U2804 (N_2804,N_1314,N_360);
nor U2805 (N_2805,N_1072,N_446);
or U2806 (N_2806,N_1996,N_1805);
nor U2807 (N_2807,N_974,N_1650);
or U2808 (N_2808,N_212,N_1579);
or U2809 (N_2809,N_879,N_1012);
and U2810 (N_2810,N_1919,N_1441);
nand U2811 (N_2811,N_1409,N_587);
or U2812 (N_2812,N_1716,N_1524);
nor U2813 (N_2813,N_1939,N_1952);
nor U2814 (N_2814,N_1469,N_565);
nand U2815 (N_2815,N_1116,N_969);
or U2816 (N_2816,N_956,N_582);
nand U2817 (N_2817,N_694,N_724);
or U2818 (N_2818,N_706,N_118);
and U2819 (N_2819,N_99,N_286);
and U2820 (N_2820,N_766,N_356);
and U2821 (N_2821,N_1322,N_162);
nor U2822 (N_2822,N_739,N_143);
nor U2823 (N_2823,N_1383,N_1597);
nor U2824 (N_2824,N_1992,N_1175);
nor U2825 (N_2825,N_1327,N_1717);
and U2826 (N_2826,N_1245,N_532);
nand U2827 (N_2827,N_1124,N_1526);
nor U2828 (N_2828,N_1760,N_1448);
or U2829 (N_2829,N_1313,N_1600);
and U2830 (N_2830,N_780,N_192);
nand U2831 (N_2831,N_236,N_1781);
nor U2832 (N_2832,N_382,N_1193);
and U2833 (N_2833,N_1392,N_1257);
nand U2834 (N_2834,N_1715,N_1744);
and U2835 (N_2835,N_137,N_1251);
or U2836 (N_2836,N_1372,N_1118);
or U2837 (N_2837,N_973,N_95);
nand U2838 (N_2838,N_1784,N_910);
and U2839 (N_2839,N_699,N_1326);
nand U2840 (N_2840,N_223,N_1387);
nor U2841 (N_2841,N_1024,N_1052);
or U2842 (N_2842,N_127,N_132);
or U2843 (N_2843,N_1776,N_1421);
and U2844 (N_2844,N_751,N_1133);
nor U2845 (N_2845,N_1338,N_603);
and U2846 (N_2846,N_48,N_1927);
nor U2847 (N_2847,N_108,N_1510);
nor U2848 (N_2848,N_367,N_120);
nand U2849 (N_2849,N_352,N_404);
or U2850 (N_2850,N_1741,N_932);
nand U2851 (N_2851,N_769,N_1961);
nor U2852 (N_2852,N_965,N_1178);
nand U2853 (N_2853,N_1586,N_1099);
nand U2854 (N_2854,N_218,N_851);
and U2855 (N_2855,N_1560,N_1287);
or U2856 (N_2856,N_1608,N_744);
or U2857 (N_2857,N_82,N_1339);
nor U2858 (N_2858,N_199,N_391);
nand U2859 (N_2859,N_110,N_1501);
or U2860 (N_2860,N_1985,N_1653);
nor U2861 (N_2861,N_900,N_87);
nand U2862 (N_2862,N_1400,N_892);
nand U2863 (N_2863,N_1306,N_1694);
and U2864 (N_2864,N_149,N_1915);
or U2865 (N_2865,N_38,N_1220);
and U2866 (N_2866,N_1205,N_785);
and U2867 (N_2867,N_758,N_326);
nand U2868 (N_2868,N_1183,N_283);
and U2869 (N_2869,N_1604,N_524);
or U2870 (N_2870,N_428,N_1634);
xor U2871 (N_2871,N_1223,N_989);
or U2872 (N_2872,N_883,N_161);
nor U2873 (N_2873,N_28,N_1230);
nor U2874 (N_2874,N_64,N_1909);
and U2875 (N_2875,N_1076,N_52);
or U2876 (N_2876,N_1152,N_1446);
nand U2877 (N_2877,N_546,N_960);
and U2878 (N_2878,N_1450,N_447);
and U2879 (N_2879,N_1747,N_1038);
nor U2880 (N_2880,N_1049,N_1426);
nand U2881 (N_2881,N_499,N_839);
nor U2882 (N_2882,N_736,N_1186);
and U2883 (N_2883,N_1034,N_1861);
nand U2884 (N_2884,N_640,N_347);
nand U2885 (N_2885,N_1361,N_224);
nor U2886 (N_2886,N_241,N_778);
nand U2887 (N_2887,N_1707,N_791);
nand U2888 (N_2888,N_305,N_466);
nor U2889 (N_2889,N_101,N_1112);
nand U2890 (N_2890,N_1170,N_1914);
or U2891 (N_2891,N_1141,N_1549);
nand U2892 (N_2892,N_1035,N_719);
nor U2893 (N_2893,N_1812,N_816);
nor U2894 (N_2894,N_609,N_1105);
or U2895 (N_2895,N_727,N_170);
and U2896 (N_2896,N_1184,N_354);
nand U2897 (N_2897,N_1020,N_740);
and U2898 (N_2898,N_1821,N_1705);
nor U2899 (N_2899,N_987,N_756);
or U2900 (N_2900,N_1022,N_1571);
and U2901 (N_2901,N_596,N_53);
nand U2902 (N_2902,N_385,N_1185);
nor U2903 (N_2903,N_730,N_1761);
nor U2904 (N_2904,N_1281,N_1129);
nand U2905 (N_2905,N_1953,N_316);
nand U2906 (N_2906,N_1470,N_215);
and U2907 (N_2907,N_835,N_1616);
or U2908 (N_2908,N_1817,N_1356);
nor U2909 (N_2909,N_585,N_1447);
nor U2910 (N_2910,N_338,N_1808);
nor U2911 (N_2911,N_1623,N_186);
nand U2912 (N_2912,N_104,N_870);
nor U2913 (N_2913,N_630,N_1959);
or U2914 (N_2914,N_636,N_1793);
and U2915 (N_2915,N_498,N_150);
nand U2916 (N_2916,N_1286,N_561);
or U2917 (N_2917,N_801,N_711);
or U2918 (N_2918,N_1547,N_1297);
nand U2919 (N_2919,N_1575,N_741);
and U2920 (N_2920,N_671,N_443);
or U2921 (N_2921,N_425,N_1015);
and U2922 (N_2922,N_1337,N_975);
or U2923 (N_2923,N_1945,N_1610);
or U2924 (N_2924,N_457,N_1801);
and U2925 (N_2925,N_262,N_742);
nand U2926 (N_2926,N_1202,N_1908);
nor U2927 (N_2927,N_1191,N_1351);
nor U2928 (N_2928,N_219,N_1675);
or U2929 (N_2929,N_1323,N_235);
and U2930 (N_2930,N_1831,N_655);
and U2931 (N_2931,N_917,N_692);
nand U2932 (N_2932,N_56,N_390);
and U2933 (N_2933,N_483,N_1439);
nand U2934 (N_2934,N_9,N_113);
nand U2935 (N_2935,N_159,N_1594);
nor U2936 (N_2936,N_868,N_72);
nand U2937 (N_2937,N_983,N_1455);
nand U2938 (N_2938,N_1700,N_1452);
or U2939 (N_2939,N_1657,N_849);
nor U2940 (N_2940,N_1158,N_533);
nand U2941 (N_2941,N_1268,N_234);
and U2942 (N_2942,N_24,N_76);
and U2943 (N_2943,N_597,N_941);
and U2944 (N_2944,N_1837,N_383);
nor U2945 (N_2945,N_764,N_909);
nand U2946 (N_2946,N_1055,N_770);
or U2947 (N_2947,N_1598,N_35);
nand U2948 (N_2948,N_1299,N_607);
and U2949 (N_2949,N_673,N_1098);
or U2950 (N_2950,N_1563,N_115);
and U2951 (N_2951,N_859,N_1162);
nor U2952 (N_2952,N_1244,N_1463);
and U2953 (N_2953,N_196,N_760);
nand U2954 (N_2954,N_1107,N_1200);
and U2955 (N_2955,N_100,N_1404);
and U2956 (N_2956,N_1655,N_1260);
or U2957 (N_2957,N_1918,N_1807);
nor U2958 (N_2958,N_1496,N_146);
nor U2959 (N_2959,N_1430,N_926);
and U2960 (N_2960,N_1008,N_1766);
nand U2961 (N_2961,N_843,N_1689);
nor U2962 (N_2962,N_411,N_1912);
or U2963 (N_2963,N_198,N_556);
nor U2964 (N_2964,N_551,N_833);
nor U2965 (N_2965,N_1122,N_264);
or U2966 (N_2966,N_1621,N_518);
nor U2967 (N_2967,N_1814,N_330);
nor U2968 (N_2968,N_1710,N_129);
nor U2969 (N_2969,N_1089,N_1010);
or U2970 (N_2970,N_629,N_1632);
and U2971 (N_2971,N_89,N_1301);
nand U2972 (N_2972,N_1923,N_1922);
nor U2973 (N_2973,N_156,N_274);
nand U2974 (N_2974,N_1767,N_1168);
and U2975 (N_2975,N_519,N_1274);
or U2976 (N_2976,N_1150,N_75);
nand U2977 (N_2977,N_712,N_798);
nand U2978 (N_2978,N_321,N_173);
or U2979 (N_2979,N_805,N_1039);
nor U2980 (N_2980,N_1104,N_1280);
or U2981 (N_2981,N_458,N_172);
or U2982 (N_2982,N_481,N_1999);
or U2983 (N_2983,N_841,N_537);
or U2984 (N_2984,N_1564,N_1307);
and U2985 (N_2985,N_1420,N_1827);
and U2986 (N_2986,N_1090,N_1360);
nand U2987 (N_2987,N_722,N_467);
and U2988 (N_2988,N_1460,N_1218);
nand U2989 (N_2989,N_1954,N_679);
or U2990 (N_2990,N_65,N_786);
and U2991 (N_2991,N_266,N_459);
or U2992 (N_2992,N_1029,N_92);
and U2993 (N_2993,N_1342,N_1759);
nor U2994 (N_2994,N_504,N_1068);
or U2995 (N_2995,N_1196,N_901);
nand U2996 (N_2996,N_1106,N_1067);
nor U2997 (N_2997,N_1968,N_545);
and U2998 (N_2998,N_10,N_1512);
nor U2999 (N_2999,N_1258,N_1899);
and U3000 (N_3000,N_684,N_876);
nor U3001 (N_3001,N_697,N_831);
nor U3002 (N_3002,N_1447,N_701);
or U3003 (N_3003,N_945,N_919);
or U3004 (N_3004,N_387,N_751);
and U3005 (N_3005,N_1841,N_742);
and U3006 (N_3006,N_471,N_1525);
and U3007 (N_3007,N_1751,N_367);
and U3008 (N_3008,N_757,N_411);
nor U3009 (N_3009,N_1762,N_1131);
nor U3010 (N_3010,N_1452,N_102);
or U3011 (N_3011,N_1653,N_396);
nor U3012 (N_3012,N_690,N_1840);
and U3013 (N_3013,N_1426,N_1616);
nand U3014 (N_3014,N_1663,N_500);
or U3015 (N_3015,N_689,N_1461);
nand U3016 (N_3016,N_1113,N_1322);
nand U3017 (N_3017,N_416,N_1357);
or U3018 (N_3018,N_936,N_931);
or U3019 (N_3019,N_1974,N_991);
or U3020 (N_3020,N_1337,N_375);
and U3021 (N_3021,N_1076,N_985);
or U3022 (N_3022,N_1433,N_1339);
or U3023 (N_3023,N_1287,N_1188);
and U3024 (N_3024,N_1123,N_1458);
or U3025 (N_3025,N_1015,N_1567);
nor U3026 (N_3026,N_1657,N_1371);
and U3027 (N_3027,N_1664,N_1484);
nand U3028 (N_3028,N_836,N_621);
and U3029 (N_3029,N_59,N_147);
or U3030 (N_3030,N_1323,N_562);
and U3031 (N_3031,N_1352,N_364);
nor U3032 (N_3032,N_481,N_1701);
nand U3033 (N_3033,N_1856,N_445);
nor U3034 (N_3034,N_1142,N_609);
or U3035 (N_3035,N_796,N_1016);
nand U3036 (N_3036,N_1313,N_1881);
nand U3037 (N_3037,N_1998,N_1329);
nor U3038 (N_3038,N_460,N_328);
nor U3039 (N_3039,N_98,N_413);
and U3040 (N_3040,N_943,N_251);
or U3041 (N_3041,N_1556,N_1176);
and U3042 (N_3042,N_621,N_694);
and U3043 (N_3043,N_707,N_1572);
and U3044 (N_3044,N_1461,N_1271);
nand U3045 (N_3045,N_85,N_220);
or U3046 (N_3046,N_1952,N_5);
nor U3047 (N_3047,N_107,N_1637);
or U3048 (N_3048,N_1152,N_1450);
or U3049 (N_3049,N_1737,N_612);
nand U3050 (N_3050,N_132,N_1681);
nor U3051 (N_3051,N_985,N_1264);
nand U3052 (N_3052,N_1338,N_428);
nor U3053 (N_3053,N_1,N_1426);
and U3054 (N_3054,N_261,N_1783);
and U3055 (N_3055,N_507,N_488);
nor U3056 (N_3056,N_401,N_1910);
nor U3057 (N_3057,N_802,N_1580);
nor U3058 (N_3058,N_958,N_1465);
and U3059 (N_3059,N_298,N_1316);
nor U3060 (N_3060,N_1036,N_749);
and U3061 (N_3061,N_1600,N_519);
nor U3062 (N_3062,N_1594,N_336);
nor U3063 (N_3063,N_26,N_886);
nor U3064 (N_3064,N_761,N_10);
or U3065 (N_3065,N_258,N_941);
nor U3066 (N_3066,N_626,N_1166);
and U3067 (N_3067,N_1041,N_452);
or U3068 (N_3068,N_21,N_1269);
and U3069 (N_3069,N_220,N_5);
and U3070 (N_3070,N_980,N_1505);
nor U3071 (N_3071,N_1577,N_1106);
or U3072 (N_3072,N_312,N_924);
or U3073 (N_3073,N_1397,N_1658);
or U3074 (N_3074,N_171,N_645);
nand U3075 (N_3075,N_620,N_252);
nor U3076 (N_3076,N_1318,N_1333);
and U3077 (N_3077,N_1417,N_1652);
nand U3078 (N_3078,N_1550,N_1834);
nand U3079 (N_3079,N_1546,N_1334);
and U3080 (N_3080,N_1311,N_901);
nand U3081 (N_3081,N_1217,N_1543);
or U3082 (N_3082,N_875,N_1793);
or U3083 (N_3083,N_916,N_928);
nor U3084 (N_3084,N_649,N_19);
nor U3085 (N_3085,N_209,N_1642);
or U3086 (N_3086,N_617,N_183);
and U3087 (N_3087,N_93,N_324);
and U3088 (N_3088,N_1184,N_1601);
or U3089 (N_3089,N_826,N_100);
nor U3090 (N_3090,N_338,N_802);
and U3091 (N_3091,N_285,N_1449);
nand U3092 (N_3092,N_139,N_1726);
nand U3093 (N_3093,N_1516,N_1639);
or U3094 (N_3094,N_987,N_1540);
xnor U3095 (N_3095,N_560,N_1039);
or U3096 (N_3096,N_1541,N_1279);
and U3097 (N_3097,N_140,N_810);
or U3098 (N_3098,N_1735,N_213);
nor U3099 (N_3099,N_1967,N_104);
or U3100 (N_3100,N_163,N_1574);
and U3101 (N_3101,N_1700,N_1623);
and U3102 (N_3102,N_1806,N_653);
nor U3103 (N_3103,N_407,N_159);
nand U3104 (N_3104,N_336,N_861);
nor U3105 (N_3105,N_1463,N_1353);
xnor U3106 (N_3106,N_51,N_956);
nand U3107 (N_3107,N_307,N_1482);
nor U3108 (N_3108,N_1283,N_1254);
and U3109 (N_3109,N_321,N_1382);
xor U3110 (N_3110,N_1155,N_923);
and U3111 (N_3111,N_1897,N_885);
nand U3112 (N_3112,N_546,N_1266);
and U3113 (N_3113,N_560,N_1618);
nor U3114 (N_3114,N_1527,N_815);
and U3115 (N_3115,N_377,N_470);
nand U3116 (N_3116,N_257,N_1874);
nor U3117 (N_3117,N_1362,N_832);
nor U3118 (N_3118,N_792,N_1801);
nand U3119 (N_3119,N_406,N_1161);
nor U3120 (N_3120,N_739,N_60);
or U3121 (N_3121,N_507,N_1510);
nand U3122 (N_3122,N_674,N_590);
or U3123 (N_3123,N_874,N_214);
nor U3124 (N_3124,N_41,N_1376);
and U3125 (N_3125,N_757,N_77);
or U3126 (N_3126,N_1111,N_1893);
nand U3127 (N_3127,N_435,N_1968);
and U3128 (N_3128,N_1319,N_360);
nand U3129 (N_3129,N_420,N_108);
and U3130 (N_3130,N_846,N_1322);
or U3131 (N_3131,N_1619,N_561);
or U3132 (N_3132,N_1011,N_1177);
nor U3133 (N_3133,N_804,N_167);
and U3134 (N_3134,N_795,N_1361);
nand U3135 (N_3135,N_513,N_1890);
nand U3136 (N_3136,N_1889,N_385);
nor U3137 (N_3137,N_1658,N_1528);
nor U3138 (N_3138,N_475,N_1615);
nor U3139 (N_3139,N_535,N_823);
nand U3140 (N_3140,N_917,N_1475);
nand U3141 (N_3141,N_922,N_1355);
and U3142 (N_3142,N_460,N_682);
nand U3143 (N_3143,N_1526,N_1858);
nand U3144 (N_3144,N_317,N_1333);
nand U3145 (N_3145,N_10,N_1164);
or U3146 (N_3146,N_579,N_1061);
or U3147 (N_3147,N_1657,N_612);
nor U3148 (N_3148,N_1068,N_317);
and U3149 (N_3149,N_1223,N_1182);
nand U3150 (N_3150,N_1836,N_1602);
nand U3151 (N_3151,N_1502,N_1123);
nand U3152 (N_3152,N_1464,N_261);
and U3153 (N_3153,N_664,N_998);
and U3154 (N_3154,N_14,N_1942);
nor U3155 (N_3155,N_233,N_1551);
nand U3156 (N_3156,N_523,N_1332);
nor U3157 (N_3157,N_1809,N_1772);
and U3158 (N_3158,N_1082,N_269);
nand U3159 (N_3159,N_852,N_398);
and U3160 (N_3160,N_1793,N_125);
nor U3161 (N_3161,N_480,N_1598);
nor U3162 (N_3162,N_1670,N_1693);
and U3163 (N_3163,N_119,N_1991);
nor U3164 (N_3164,N_54,N_148);
nand U3165 (N_3165,N_1376,N_1212);
and U3166 (N_3166,N_1217,N_950);
or U3167 (N_3167,N_906,N_1339);
or U3168 (N_3168,N_636,N_682);
nand U3169 (N_3169,N_732,N_3);
nand U3170 (N_3170,N_448,N_1407);
nand U3171 (N_3171,N_1015,N_205);
or U3172 (N_3172,N_1675,N_185);
or U3173 (N_3173,N_1172,N_1301);
nor U3174 (N_3174,N_880,N_1403);
xor U3175 (N_3175,N_846,N_1454);
or U3176 (N_3176,N_1816,N_979);
nand U3177 (N_3177,N_1415,N_664);
nor U3178 (N_3178,N_735,N_1593);
xor U3179 (N_3179,N_996,N_1384);
or U3180 (N_3180,N_1669,N_348);
or U3181 (N_3181,N_489,N_696);
nor U3182 (N_3182,N_1433,N_719);
or U3183 (N_3183,N_1685,N_388);
or U3184 (N_3184,N_369,N_1424);
nor U3185 (N_3185,N_380,N_968);
nand U3186 (N_3186,N_1239,N_1971);
nor U3187 (N_3187,N_855,N_680);
nor U3188 (N_3188,N_32,N_1710);
and U3189 (N_3189,N_1077,N_1348);
or U3190 (N_3190,N_849,N_795);
nand U3191 (N_3191,N_74,N_501);
nand U3192 (N_3192,N_1875,N_1675);
or U3193 (N_3193,N_1573,N_1021);
nor U3194 (N_3194,N_906,N_1144);
and U3195 (N_3195,N_262,N_781);
nand U3196 (N_3196,N_1296,N_953);
nor U3197 (N_3197,N_314,N_1407);
or U3198 (N_3198,N_1779,N_164);
nand U3199 (N_3199,N_880,N_1943);
or U3200 (N_3200,N_99,N_310);
or U3201 (N_3201,N_134,N_7);
nand U3202 (N_3202,N_187,N_816);
nor U3203 (N_3203,N_1154,N_1156);
nor U3204 (N_3204,N_1212,N_1700);
or U3205 (N_3205,N_1212,N_1341);
and U3206 (N_3206,N_974,N_634);
and U3207 (N_3207,N_642,N_1642);
and U3208 (N_3208,N_1999,N_801);
xor U3209 (N_3209,N_61,N_480);
and U3210 (N_3210,N_1361,N_1802);
nor U3211 (N_3211,N_816,N_228);
nand U3212 (N_3212,N_796,N_68);
nor U3213 (N_3213,N_1033,N_651);
nor U3214 (N_3214,N_1887,N_1988);
and U3215 (N_3215,N_309,N_1768);
nand U3216 (N_3216,N_1619,N_134);
nor U3217 (N_3217,N_1395,N_39);
nor U3218 (N_3218,N_1453,N_1983);
and U3219 (N_3219,N_1751,N_630);
nand U3220 (N_3220,N_1492,N_1135);
or U3221 (N_3221,N_1228,N_406);
nand U3222 (N_3222,N_400,N_343);
or U3223 (N_3223,N_187,N_115);
or U3224 (N_3224,N_490,N_77);
or U3225 (N_3225,N_1379,N_980);
or U3226 (N_3226,N_411,N_758);
nand U3227 (N_3227,N_1510,N_1770);
or U3228 (N_3228,N_154,N_1164);
nor U3229 (N_3229,N_55,N_1939);
nor U3230 (N_3230,N_1337,N_831);
nor U3231 (N_3231,N_1745,N_1502);
nor U3232 (N_3232,N_1494,N_237);
and U3233 (N_3233,N_1546,N_1734);
nor U3234 (N_3234,N_833,N_1611);
nor U3235 (N_3235,N_1205,N_452);
nand U3236 (N_3236,N_595,N_1913);
nor U3237 (N_3237,N_1470,N_1110);
nor U3238 (N_3238,N_905,N_1750);
and U3239 (N_3239,N_390,N_1250);
nor U3240 (N_3240,N_893,N_618);
nor U3241 (N_3241,N_712,N_1849);
or U3242 (N_3242,N_1545,N_1790);
nor U3243 (N_3243,N_1711,N_1472);
and U3244 (N_3244,N_987,N_1816);
and U3245 (N_3245,N_1027,N_175);
and U3246 (N_3246,N_1144,N_464);
and U3247 (N_3247,N_715,N_962);
and U3248 (N_3248,N_388,N_1884);
nand U3249 (N_3249,N_1055,N_1977);
nand U3250 (N_3250,N_400,N_86);
and U3251 (N_3251,N_237,N_1212);
nor U3252 (N_3252,N_270,N_1802);
or U3253 (N_3253,N_484,N_1317);
and U3254 (N_3254,N_1045,N_812);
nand U3255 (N_3255,N_1701,N_5);
and U3256 (N_3256,N_885,N_1147);
nor U3257 (N_3257,N_1482,N_1426);
xor U3258 (N_3258,N_1552,N_176);
or U3259 (N_3259,N_64,N_854);
nor U3260 (N_3260,N_1976,N_904);
or U3261 (N_3261,N_1908,N_976);
or U3262 (N_3262,N_1316,N_1726);
nand U3263 (N_3263,N_416,N_1153);
and U3264 (N_3264,N_1937,N_1316);
nand U3265 (N_3265,N_433,N_1374);
nand U3266 (N_3266,N_1036,N_117);
and U3267 (N_3267,N_1631,N_1497);
or U3268 (N_3268,N_451,N_1627);
nand U3269 (N_3269,N_30,N_400);
and U3270 (N_3270,N_755,N_1360);
nor U3271 (N_3271,N_106,N_267);
and U3272 (N_3272,N_1658,N_391);
and U3273 (N_3273,N_955,N_1774);
or U3274 (N_3274,N_1118,N_1325);
nand U3275 (N_3275,N_178,N_914);
nor U3276 (N_3276,N_1852,N_1752);
nor U3277 (N_3277,N_805,N_1706);
or U3278 (N_3278,N_1425,N_648);
and U3279 (N_3279,N_646,N_694);
nor U3280 (N_3280,N_1446,N_1595);
nand U3281 (N_3281,N_427,N_311);
and U3282 (N_3282,N_359,N_1553);
and U3283 (N_3283,N_1512,N_928);
nor U3284 (N_3284,N_1666,N_1949);
or U3285 (N_3285,N_1226,N_182);
nand U3286 (N_3286,N_490,N_367);
or U3287 (N_3287,N_1564,N_73);
nand U3288 (N_3288,N_1707,N_1561);
or U3289 (N_3289,N_360,N_676);
nand U3290 (N_3290,N_1045,N_644);
nand U3291 (N_3291,N_1515,N_303);
xor U3292 (N_3292,N_1885,N_1487);
nand U3293 (N_3293,N_1979,N_450);
nor U3294 (N_3294,N_1562,N_158);
nor U3295 (N_3295,N_487,N_1276);
or U3296 (N_3296,N_327,N_510);
nand U3297 (N_3297,N_74,N_557);
nor U3298 (N_3298,N_1321,N_1724);
xnor U3299 (N_3299,N_495,N_1143);
xnor U3300 (N_3300,N_645,N_29);
and U3301 (N_3301,N_813,N_172);
and U3302 (N_3302,N_1283,N_831);
nor U3303 (N_3303,N_688,N_429);
nand U3304 (N_3304,N_1402,N_823);
nor U3305 (N_3305,N_1755,N_1866);
and U3306 (N_3306,N_496,N_1528);
nand U3307 (N_3307,N_1779,N_1967);
and U3308 (N_3308,N_874,N_1214);
or U3309 (N_3309,N_599,N_170);
and U3310 (N_3310,N_1744,N_758);
and U3311 (N_3311,N_945,N_1654);
nand U3312 (N_3312,N_468,N_1718);
or U3313 (N_3313,N_1560,N_36);
or U3314 (N_3314,N_1823,N_1307);
and U3315 (N_3315,N_1210,N_344);
nor U3316 (N_3316,N_383,N_695);
and U3317 (N_3317,N_157,N_1664);
nor U3318 (N_3318,N_713,N_970);
and U3319 (N_3319,N_1035,N_84);
nor U3320 (N_3320,N_104,N_1451);
nand U3321 (N_3321,N_1953,N_406);
nor U3322 (N_3322,N_1723,N_1040);
xnor U3323 (N_3323,N_1518,N_471);
nor U3324 (N_3324,N_378,N_1754);
or U3325 (N_3325,N_540,N_1852);
and U3326 (N_3326,N_1565,N_907);
or U3327 (N_3327,N_619,N_351);
or U3328 (N_3328,N_1778,N_1270);
nand U3329 (N_3329,N_513,N_1519);
and U3330 (N_3330,N_920,N_1694);
or U3331 (N_3331,N_808,N_589);
nand U3332 (N_3332,N_1996,N_1851);
or U3333 (N_3333,N_693,N_499);
nand U3334 (N_3334,N_1626,N_953);
nor U3335 (N_3335,N_464,N_1635);
and U3336 (N_3336,N_532,N_796);
or U3337 (N_3337,N_1577,N_1551);
and U3338 (N_3338,N_1674,N_530);
and U3339 (N_3339,N_865,N_529);
or U3340 (N_3340,N_1361,N_895);
and U3341 (N_3341,N_404,N_699);
nor U3342 (N_3342,N_489,N_1913);
or U3343 (N_3343,N_1303,N_944);
nand U3344 (N_3344,N_37,N_308);
and U3345 (N_3345,N_1275,N_1764);
and U3346 (N_3346,N_1339,N_1603);
or U3347 (N_3347,N_923,N_177);
or U3348 (N_3348,N_1744,N_1116);
nor U3349 (N_3349,N_278,N_202);
and U3350 (N_3350,N_390,N_1311);
nand U3351 (N_3351,N_646,N_537);
nand U3352 (N_3352,N_157,N_1307);
nand U3353 (N_3353,N_438,N_354);
or U3354 (N_3354,N_1473,N_1105);
and U3355 (N_3355,N_637,N_1545);
or U3356 (N_3356,N_1053,N_430);
or U3357 (N_3357,N_1309,N_623);
nor U3358 (N_3358,N_889,N_1960);
or U3359 (N_3359,N_1506,N_1515);
nor U3360 (N_3360,N_346,N_1406);
and U3361 (N_3361,N_285,N_1559);
and U3362 (N_3362,N_1511,N_373);
or U3363 (N_3363,N_1880,N_1572);
or U3364 (N_3364,N_1091,N_566);
nand U3365 (N_3365,N_1897,N_523);
nand U3366 (N_3366,N_220,N_773);
or U3367 (N_3367,N_1900,N_440);
and U3368 (N_3368,N_1219,N_749);
nor U3369 (N_3369,N_1850,N_1249);
nand U3370 (N_3370,N_270,N_1509);
or U3371 (N_3371,N_576,N_1512);
nor U3372 (N_3372,N_603,N_821);
and U3373 (N_3373,N_500,N_1007);
nor U3374 (N_3374,N_541,N_1472);
xnor U3375 (N_3375,N_91,N_1623);
nand U3376 (N_3376,N_801,N_1475);
nor U3377 (N_3377,N_1497,N_1763);
nor U3378 (N_3378,N_1966,N_201);
nor U3379 (N_3379,N_1580,N_424);
nand U3380 (N_3380,N_1846,N_489);
nor U3381 (N_3381,N_1426,N_504);
or U3382 (N_3382,N_1763,N_1293);
and U3383 (N_3383,N_865,N_1727);
or U3384 (N_3384,N_471,N_1498);
nand U3385 (N_3385,N_1197,N_1393);
and U3386 (N_3386,N_1850,N_387);
or U3387 (N_3387,N_762,N_24);
nand U3388 (N_3388,N_971,N_321);
and U3389 (N_3389,N_1493,N_854);
and U3390 (N_3390,N_1268,N_318);
and U3391 (N_3391,N_622,N_115);
nand U3392 (N_3392,N_1930,N_1672);
and U3393 (N_3393,N_1562,N_247);
or U3394 (N_3394,N_713,N_634);
nor U3395 (N_3395,N_1497,N_260);
nand U3396 (N_3396,N_1052,N_1614);
nand U3397 (N_3397,N_494,N_1232);
and U3398 (N_3398,N_613,N_1745);
nand U3399 (N_3399,N_494,N_1269);
and U3400 (N_3400,N_1663,N_651);
nand U3401 (N_3401,N_1348,N_1927);
and U3402 (N_3402,N_87,N_389);
and U3403 (N_3403,N_991,N_476);
nand U3404 (N_3404,N_1757,N_322);
and U3405 (N_3405,N_1239,N_94);
and U3406 (N_3406,N_25,N_1291);
and U3407 (N_3407,N_1156,N_1193);
nand U3408 (N_3408,N_241,N_1664);
or U3409 (N_3409,N_738,N_61);
and U3410 (N_3410,N_738,N_1523);
nand U3411 (N_3411,N_1393,N_188);
or U3412 (N_3412,N_111,N_993);
nand U3413 (N_3413,N_653,N_1913);
or U3414 (N_3414,N_1859,N_1700);
and U3415 (N_3415,N_1556,N_1762);
or U3416 (N_3416,N_270,N_1823);
or U3417 (N_3417,N_506,N_1941);
nand U3418 (N_3418,N_503,N_1527);
nand U3419 (N_3419,N_613,N_389);
or U3420 (N_3420,N_389,N_924);
nor U3421 (N_3421,N_1154,N_1337);
nor U3422 (N_3422,N_631,N_106);
or U3423 (N_3423,N_627,N_605);
nand U3424 (N_3424,N_1538,N_1834);
nand U3425 (N_3425,N_1708,N_782);
nand U3426 (N_3426,N_138,N_1029);
and U3427 (N_3427,N_936,N_1963);
nand U3428 (N_3428,N_13,N_473);
and U3429 (N_3429,N_112,N_1741);
and U3430 (N_3430,N_1671,N_776);
and U3431 (N_3431,N_946,N_681);
or U3432 (N_3432,N_1668,N_482);
nor U3433 (N_3433,N_602,N_596);
nor U3434 (N_3434,N_136,N_1291);
nor U3435 (N_3435,N_1566,N_1848);
nor U3436 (N_3436,N_744,N_1176);
nand U3437 (N_3437,N_635,N_463);
and U3438 (N_3438,N_239,N_303);
nor U3439 (N_3439,N_491,N_1074);
nor U3440 (N_3440,N_486,N_344);
or U3441 (N_3441,N_504,N_1596);
nor U3442 (N_3442,N_1865,N_1427);
nand U3443 (N_3443,N_1432,N_763);
nor U3444 (N_3444,N_701,N_965);
and U3445 (N_3445,N_555,N_620);
and U3446 (N_3446,N_660,N_1655);
nor U3447 (N_3447,N_293,N_1301);
or U3448 (N_3448,N_535,N_1406);
or U3449 (N_3449,N_142,N_340);
nand U3450 (N_3450,N_91,N_832);
or U3451 (N_3451,N_1729,N_125);
nand U3452 (N_3452,N_939,N_248);
and U3453 (N_3453,N_1380,N_341);
or U3454 (N_3454,N_850,N_648);
nand U3455 (N_3455,N_266,N_1179);
nand U3456 (N_3456,N_1455,N_954);
and U3457 (N_3457,N_436,N_751);
or U3458 (N_3458,N_1972,N_1028);
and U3459 (N_3459,N_195,N_1754);
and U3460 (N_3460,N_1578,N_1767);
nor U3461 (N_3461,N_776,N_378);
nand U3462 (N_3462,N_80,N_1406);
nor U3463 (N_3463,N_1525,N_1419);
nand U3464 (N_3464,N_864,N_1300);
nand U3465 (N_3465,N_1833,N_576);
nor U3466 (N_3466,N_446,N_1545);
nand U3467 (N_3467,N_1591,N_1696);
or U3468 (N_3468,N_312,N_1524);
nor U3469 (N_3469,N_1796,N_311);
nand U3470 (N_3470,N_869,N_1494);
nand U3471 (N_3471,N_295,N_4);
and U3472 (N_3472,N_78,N_1104);
nand U3473 (N_3473,N_1881,N_855);
nor U3474 (N_3474,N_1814,N_1521);
or U3475 (N_3475,N_1896,N_1997);
and U3476 (N_3476,N_64,N_765);
nor U3477 (N_3477,N_1753,N_237);
and U3478 (N_3478,N_1531,N_1748);
nor U3479 (N_3479,N_1781,N_1698);
and U3480 (N_3480,N_263,N_1532);
and U3481 (N_3481,N_1270,N_1154);
or U3482 (N_3482,N_1970,N_346);
or U3483 (N_3483,N_468,N_414);
and U3484 (N_3484,N_974,N_13);
nor U3485 (N_3485,N_631,N_1804);
or U3486 (N_3486,N_1880,N_202);
or U3487 (N_3487,N_392,N_1988);
and U3488 (N_3488,N_851,N_1747);
or U3489 (N_3489,N_1366,N_206);
nand U3490 (N_3490,N_785,N_1560);
or U3491 (N_3491,N_1794,N_1776);
or U3492 (N_3492,N_1923,N_267);
nand U3493 (N_3493,N_1412,N_1361);
nor U3494 (N_3494,N_1799,N_1161);
nand U3495 (N_3495,N_1075,N_1929);
or U3496 (N_3496,N_945,N_335);
or U3497 (N_3497,N_1822,N_969);
and U3498 (N_3498,N_550,N_209);
and U3499 (N_3499,N_497,N_309);
nand U3500 (N_3500,N_881,N_928);
nor U3501 (N_3501,N_776,N_1710);
or U3502 (N_3502,N_401,N_1700);
or U3503 (N_3503,N_20,N_1088);
nor U3504 (N_3504,N_866,N_1459);
nand U3505 (N_3505,N_1418,N_676);
or U3506 (N_3506,N_805,N_527);
nand U3507 (N_3507,N_23,N_887);
nor U3508 (N_3508,N_1035,N_1501);
or U3509 (N_3509,N_1243,N_361);
and U3510 (N_3510,N_910,N_1840);
nor U3511 (N_3511,N_1229,N_18);
or U3512 (N_3512,N_1612,N_1690);
nor U3513 (N_3513,N_796,N_264);
nor U3514 (N_3514,N_1610,N_1033);
xnor U3515 (N_3515,N_1079,N_90);
nor U3516 (N_3516,N_1507,N_1375);
nand U3517 (N_3517,N_383,N_1774);
nand U3518 (N_3518,N_1605,N_1660);
and U3519 (N_3519,N_1564,N_1088);
and U3520 (N_3520,N_267,N_1253);
nor U3521 (N_3521,N_1676,N_881);
or U3522 (N_3522,N_1632,N_149);
nor U3523 (N_3523,N_1401,N_1197);
or U3524 (N_3524,N_1469,N_183);
or U3525 (N_3525,N_765,N_1525);
or U3526 (N_3526,N_1605,N_1523);
and U3527 (N_3527,N_1302,N_1060);
nand U3528 (N_3528,N_1687,N_221);
xor U3529 (N_3529,N_340,N_788);
nand U3530 (N_3530,N_1380,N_630);
nand U3531 (N_3531,N_972,N_411);
nand U3532 (N_3532,N_1414,N_621);
nor U3533 (N_3533,N_601,N_1069);
and U3534 (N_3534,N_1843,N_778);
nor U3535 (N_3535,N_430,N_1997);
nand U3536 (N_3536,N_1979,N_379);
nor U3537 (N_3537,N_91,N_1295);
nand U3538 (N_3538,N_1150,N_607);
nor U3539 (N_3539,N_71,N_383);
or U3540 (N_3540,N_534,N_1506);
or U3541 (N_3541,N_1043,N_1064);
nand U3542 (N_3542,N_1603,N_221);
or U3543 (N_3543,N_389,N_1106);
and U3544 (N_3544,N_1256,N_1262);
or U3545 (N_3545,N_809,N_766);
or U3546 (N_3546,N_1131,N_1365);
nor U3547 (N_3547,N_30,N_1745);
and U3548 (N_3548,N_741,N_99);
and U3549 (N_3549,N_646,N_770);
nor U3550 (N_3550,N_51,N_1370);
and U3551 (N_3551,N_1517,N_699);
or U3552 (N_3552,N_215,N_1058);
nand U3553 (N_3553,N_377,N_1766);
nand U3554 (N_3554,N_1538,N_1406);
nand U3555 (N_3555,N_1928,N_867);
nor U3556 (N_3556,N_1719,N_1951);
nor U3557 (N_3557,N_1968,N_307);
and U3558 (N_3558,N_265,N_692);
nand U3559 (N_3559,N_598,N_950);
nor U3560 (N_3560,N_1585,N_423);
nor U3561 (N_3561,N_283,N_933);
nand U3562 (N_3562,N_1780,N_1708);
nand U3563 (N_3563,N_1292,N_367);
nand U3564 (N_3564,N_1473,N_1214);
nand U3565 (N_3565,N_776,N_391);
nand U3566 (N_3566,N_1937,N_1031);
or U3567 (N_3567,N_1094,N_1789);
nor U3568 (N_3568,N_936,N_898);
nand U3569 (N_3569,N_942,N_1653);
nand U3570 (N_3570,N_1547,N_1746);
and U3571 (N_3571,N_1200,N_263);
nor U3572 (N_3572,N_157,N_1946);
nand U3573 (N_3573,N_287,N_530);
nor U3574 (N_3574,N_1112,N_57);
or U3575 (N_3575,N_1125,N_1767);
nor U3576 (N_3576,N_695,N_1984);
and U3577 (N_3577,N_1426,N_497);
and U3578 (N_3578,N_403,N_1626);
and U3579 (N_3579,N_1464,N_463);
and U3580 (N_3580,N_1099,N_464);
or U3581 (N_3581,N_997,N_489);
nor U3582 (N_3582,N_241,N_1700);
or U3583 (N_3583,N_1719,N_1973);
nand U3584 (N_3584,N_1930,N_1704);
nor U3585 (N_3585,N_813,N_651);
or U3586 (N_3586,N_1535,N_1996);
nand U3587 (N_3587,N_843,N_193);
and U3588 (N_3588,N_914,N_757);
nand U3589 (N_3589,N_1480,N_1587);
nand U3590 (N_3590,N_748,N_488);
and U3591 (N_3591,N_807,N_1336);
or U3592 (N_3592,N_500,N_1517);
nor U3593 (N_3593,N_237,N_207);
and U3594 (N_3594,N_539,N_1958);
and U3595 (N_3595,N_350,N_1333);
and U3596 (N_3596,N_223,N_1625);
or U3597 (N_3597,N_841,N_1026);
nor U3598 (N_3598,N_1747,N_1974);
nand U3599 (N_3599,N_1697,N_1094);
or U3600 (N_3600,N_1937,N_1038);
or U3601 (N_3601,N_1227,N_1112);
nor U3602 (N_3602,N_166,N_1961);
and U3603 (N_3603,N_346,N_200);
or U3604 (N_3604,N_1760,N_222);
xnor U3605 (N_3605,N_735,N_979);
nand U3606 (N_3606,N_1714,N_1362);
and U3607 (N_3607,N_1145,N_1827);
nand U3608 (N_3608,N_1438,N_1651);
or U3609 (N_3609,N_231,N_1399);
nand U3610 (N_3610,N_1479,N_232);
or U3611 (N_3611,N_1446,N_1287);
or U3612 (N_3612,N_1019,N_1635);
and U3613 (N_3613,N_1434,N_374);
nor U3614 (N_3614,N_1184,N_1248);
and U3615 (N_3615,N_959,N_1948);
nand U3616 (N_3616,N_1778,N_1554);
and U3617 (N_3617,N_1748,N_813);
nor U3618 (N_3618,N_1199,N_880);
nand U3619 (N_3619,N_1746,N_249);
and U3620 (N_3620,N_1458,N_1281);
or U3621 (N_3621,N_1232,N_677);
nor U3622 (N_3622,N_805,N_660);
or U3623 (N_3623,N_437,N_802);
or U3624 (N_3624,N_1692,N_787);
nor U3625 (N_3625,N_447,N_1522);
or U3626 (N_3626,N_1366,N_1600);
or U3627 (N_3627,N_726,N_198);
nor U3628 (N_3628,N_1362,N_1342);
or U3629 (N_3629,N_1092,N_1995);
nand U3630 (N_3630,N_1709,N_1735);
nor U3631 (N_3631,N_1611,N_574);
and U3632 (N_3632,N_645,N_1426);
nor U3633 (N_3633,N_1632,N_1106);
or U3634 (N_3634,N_573,N_266);
nand U3635 (N_3635,N_1615,N_1656);
nor U3636 (N_3636,N_889,N_1855);
nand U3637 (N_3637,N_581,N_1234);
and U3638 (N_3638,N_1730,N_710);
nand U3639 (N_3639,N_1996,N_1059);
nand U3640 (N_3640,N_1229,N_1312);
or U3641 (N_3641,N_962,N_1403);
and U3642 (N_3642,N_1669,N_723);
and U3643 (N_3643,N_1500,N_260);
nor U3644 (N_3644,N_1179,N_36);
nor U3645 (N_3645,N_1910,N_369);
or U3646 (N_3646,N_1973,N_1428);
nor U3647 (N_3647,N_1410,N_694);
nand U3648 (N_3648,N_1367,N_1735);
nand U3649 (N_3649,N_1902,N_262);
nand U3650 (N_3650,N_137,N_1740);
nor U3651 (N_3651,N_1014,N_1627);
nor U3652 (N_3652,N_1069,N_318);
and U3653 (N_3653,N_1947,N_359);
nand U3654 (N_3654,N_1147,N_611);
nor U3655 (N_3655,N_29,N_185);
and U3656 (N_3656,N_1956,N_784);
and U3657 (N_3657,N_1035,N_1138);
nand U3658 (N_3658,N_1202,N_1962);
or U3659 (N_3659,N_1966,N_1471);
or U3660 (N_3660,N_1846,N_1596);
nor U3661 (N_3661,N_292,N_1582);
and U3662 (N_3662,N_1730,N_1625);
nor U3663 (N_3663,N_281,N_277);
nor U3664 (N_3664,N_210,N_786);
or U3665 (N_3665,N_989,N_352);
xnor U3666 (N_3666,N_616,N_1748);
or U3667 (N_3667,N_1946,N_1943);
and U3668 (N_3668,N_471,N_1283);
and U3669 (N_3669,N_1188,N_1959);
nor U3670 (N_3670,N_295,N_1277);
nand U3671 (N_3671,N_1900,N_896);
and U3672 (N_3672,N_1553,N_320);
nor U3673 (N_3673,N_96,N_997);
nand U3674 (N_3674,N_1480,N_415);
or U3675 (N_3675,N_224,N_287);
and U3676 (N_3676,N_859,N_1394);
nand U3677 (N_3677,N_324,N_1310);
and U3678 (N_3678,N_406,N_432);
nand U3679 (N_3679,N_556,N_1961);
or U3680 (N_3680,N_1900,N_1114);
nor U3681 (N_3681,N_1052,N_693);
xnor U3682 (N_3682,N_1610,N_355);
nor U3683 (N_3683,N_1071,N_632);
nand U3684 (N_3684,N_849,N_1677);
or U3685 (N_3685,N_1174,N_1176);
nand U3686 (N_3686,N_51,N_1143);
nand U3687 (N_3687,N_682,N_1973);
nor U3688 (N_3688,N_1961,N_1039);
nand U3689 (N_3689,N_1715,N_1324);
nand U3690 (N_3690,N_581,N_955);
nor U3691 (N_3691,N_559,N_210);
nor U3692 (N_3692,N_1370,N_1645);
and U3693 (N_3693,N_1982,N_348);
nor U3694 (N_3694,N_815,N_1267);
nor U3695 (N_3695,N_715,N_229);
nand U3696 (N_3696,N_1716,N_1116);
nand U3697 (N_3697,N_617,N_688);
nand U3698 (N_3698,N_645,N_661);
or U3699 (N_3699,N_105,N_1702);
nor U3700 (N_3700,N_1086,N_1984);
or U3701 (N_3701,N_1368,N_964);
xnor U3702 (N_3702,N_1655,N_692);
or U3703 (N_3703,N_659,N_449);
nand U3704 (N_3704,N_1924,N_1785);
nor U3705 (N_3705,N_1607,N_302);
and U3706 (N_3706,N_1884,N_922);
and U3707 (N_3707,N_983,N_1909);
and U3708 (N_3708,N_576,N_1869);
and U3709 (N_3709,N_412,N_447);
nor U3710 (N_3710,N_436,N_31);
nand U3711 (N_3711,N_979,N_1915);
nor U3712 (N_3712,N_1895,N_1279);
or U3713 (N_3713,N_1331,N_1882);
and U3714 (N_3714,N_498,N_220);
nand U3715 (N_3715,N_1528,N_1886);
nand U3716 (N_3716,N_727,N_1513);
nor U3717 (N_3717,N_673,N_1619);
or U3718 (N_3718,N_1975,N_1677);
or U3719 (N_3719,N_1909,N_1448);
nor U3720 (N_3720,N_1247,N_5);
nor U3721 (N_3721,N_416,N_161);
or U3722 (N_3722,N_70,N_1723);
and U3723 (N_3723,N_1347,N_1026);
and U3724 (N_3724,N_491,N_1281);
nand U3725 (N_3725,N_1389,N_1032);
xor U3726 (N_3726,N_1762,N_164);
nor U3727 (N_3727,N_1677,N_633);
nor U3728 (N_3728,N_870,N_400);
and U3729 (N_3729,N_111,N_1090);
or U3730 (N_3730,N_1379,N_14);
or U3731 (N_3731,N_1142,N_920);
or U3732 (N_3732,N_1453,N_583);
nor U3733 (N_3733,N_1019,N_119);
or U3734 (N_3734,N_806,N_825);
nor U3735 (N_3735,N_1445,N_880);
nand U3736 (N_3736,N_1482,N_1781);
or U3737 (N_3737,N_1676,N_1507);
or U3738 (N_3738,N_1142,N_891);
nand U3739 (N_3739,N_1933,N_486);
nand U3740 (N_3740,N_1944,N_1465);
nor U3741 (N_3741,N_918,N_148);
or U3742 (N_3742,N_412,N_282);
nand U3743 (N_3743,N_1096,N_1869);
xnor U3744 (N_3744,N_297,N_376);
nor U3745 (N_3745,N_1641,N_1219);
nand U3746 (N_3746,N_1837,N_1162);
nand U3747 (N_3747,N_1951,N_547);
or U3748 (N_3748,N_847,N_1607);
nor U3749 (N_3749,N_1923,N_104);
nor U3750 (N_3750,N_1431,N_416);
or U3751 (N_3751,N_1960,N_1782);
or U3752 (N_3752,N_1036,N_1291);
and U3753 (N_3753,N_756,N_1829);
nor U3754 (N_3754,N_1719,N_845);
nor U3755 (N_3755,N_1274,N_34);
nand U3756 (N_3756,N_192,N_1450);
nand U3757 (N_3757,N_527,N_1690);
nand U3758 (N_3758,N_856,N_1592);
nand U3759 (N_3759,N_74,N_840);
nor U3760 (N_3760,N_1052,N_1453);
and U3761 (N_3761,N_1413,N_1813);
and U3762 (N_3762,N_113,N_1262);
nor U3763 (N_3763,N_473,N_1851);
or U3764 (N_3764,N_1559,N_193);
or U3765 (N_3765,N_1729,N_1061);
nor U3766 (N_3766,N_1044,N_536);
nand U3767 (N_3767,N_1335,N_994);
nor U3768 (N_3768,N_1818,N_1849);
nand U3769 (N_3769,N_953,N_105);
and U3770 (N_3770,N_1508,N_121);
nand U3771 (N_3771,N_513,N_798);
and U3772 (N_3772,N_1786,N_1899);
or U3773 (N_3773,N_1805,N_1973);
nor U3774 (N_3774,N_765,N_244);
and U3775 (N_3775,N_1116,N_959);
and U3776 (N_3776,N_768,N_1109);
and U3777 (N_3777,N_1501,N_756);
and U3778 (N_3778,N_1248,N_1157);
nand U3779 (N_3779,N_1256,N_908);
and U3780 (N_3780,N_1272,N_1168);
or U3781 (N_3781,N_460,N_1272);
or U3782 (N_3782,N_1385,N_428);
and U3783 (N_3783,N_855,N_15);
nor U3784 (N_3784,N_88,N_874);
and U3785 (N_3785,N_1989,N_1202);
and U3786 (N_3786,N_1527,N_1327);
or U3787 (N_3787,N_1199,N_623);
and U3788 (N_3788,N_1842,N_595);
or U3789 (N_3789,N_1823,N_1583);
nor U3790 (N_3790,N_1675,N_515);
or U3791 (N_3791,N_1409,N_1281);
nand U3792 (N_3792,N_72,N_490);
or U3793 (N_3793,N_1930,N_1810);
or U3794 (N_3794,N_188,N_1832);
or U3795 (N_3795,N_1142,N_486);
or U3796 (N_3796,N_1311,N_594);
nor U3797 (N_3797,N_932,N_769);
or U3798 (N_3798,N_1752,N_1673);
or U3799 (N_3799,N_220,N_608);
or U3800 (N_3800,N_310,N_145);
nand U3801 (N_3801,N_675,N_885);
and U3802 (N_3802,N_631,N_1143);
nor U3803 (N_3803,N_644,N_1389);
and U3804 (N_3804,N_184,N_537);
or U3805 (N_3805,N_1741,N_1649);
nand U3806 (N_3806,N_1556,N_1445);
nor U3807 (N_3807,N_907,N_1256);
nor U3808 (N_3808,N_799,N_1707);
nand U3809 (N_3809,N_590,N_1970);
and U3810 (N_3810,N_1689,N_86);
or U3811 (N_3811,N_1010,N_414);
nand U3812 (N_3812,N_332,N_909);
nor U3813 (N_3813,N_350,N_1478);
xnor U3814 (N_3814,N_1150,N_896);
or U3815 (N_3815,N_487,N_1812);
nor U3816 (N_3816,N_133,N_1363);
and U3817 (N_3817,N_16,N_1919);
or U3818 (N_3818,N_827,N_1370);
nor U3819 (N_3819,N_623,N_619);
and U3820 (N_3820,N_1512,N_807);
nor U3821 (N_3821,N_1301,N_454);
nor U3822 (N_3822,N_542,N_105);
nand U3823 (N_3823,N_1899,N_698);
or U3824 (N_3824,N_814,N_951);
nand U3825 (N_3825,N_1113,N_984);
or U3826 (N_3826,N_1791,N_1034);
nand U3827 (N_3827,N_1974,N_1912);
nand U3828 (N_3828,N_1939,N_1188);
nand U3829 (N_3829,N_1634,N_856);
nand U3830 (N_3830,N_845,N_1190);
nor U3831 (N_3831,N_684,N_1093);
and U3832 (N_3832,N_1756,N_923);
and U3833 (N_3833,N_878,N_298);
nand U3834 (N_3834,N_1992,N_1853);
and U3835 (N_3835,N_762,N_262);
nand U3836 (N_3836,N_46,N_68);
nor U3837 (N_3837,N_873,N_521);
nand U3838 (N_3838,N_634,N_1711);
nand U3839 (N_3839,N_283,N_749);
nand U3840 (N_3840,N_1538,N_1411);
and U3841 (N_3841,N_96,N_1927);
and U3842 (N_3842,N_480,N_936);
or U3843 (N_3843,N_1470,N_1693);
and U3844 (N_3844,N_564,N_1649);
nand U3845 (N_3845,N_799,N_1806);
nand U3846 (N_3846,N_1935,N_1147);
and U3847 (N_3847,N_465,N_1987);
and U3848 (N_3848,N_1238,N_956);
and U3849 (N_3849,N_142,N_192);
nand U3850 (N_3850,N_1996,N_1015);
and U3851 (N_3851,N_1412,N_838);
nor U3852 (N_3852,N_707,N_1003);
or U3853 (N_3853,N_780,N_549);
or U3854 (N_3854,N_646,N_367);
and U3855 (N_3855,N_58,N_726);
nor U3856 (N_3856,N_436,N_1315);
nand U3857 (N_3857,N_1267,N_294);
or U3858 (N_3858,N_1961,N_1521);
or U3859 (N_3859,N_887,N_1540);
nand U3860 (N_3860,N_832,N_664);
nor U3861 (N_3861,N_110,N_819);
or U3862 (N_3862,N_1932,N_307);
nand U3863 (N_3863,N_160,N_1969);
and U3864 (N_3864,N_1139,N_978);
nor U3865 (N_3865,N_1461,N_300);
and U3866 (N_3866,N_1246,N_492);
and U3867 (N_3867,N_50,N_506);
nand U3868 (N_3868,N_1833,N_42);
nor U3869 (N_3869,N_488,N_1242);
or U3870 (N_3870,N_267,N_1855);
nand U3871 (N_3871,N_1848,N_213);
and U3872 (N_3872,N_1118,N_1652);
or U3873 (N_3873,N_121,N_226);
nand U3874 (N_3874,N_365,N_575);
or U3875 (N_3875,N_592,N_1349);
or U3876 (N_3876,N_1404,N_1770);
nand U3877 (N_3877,N_186,N_9);
or U3878 (N_3878,N_82,N_330);
nand U3879 (N_3879,N_666,N_416);
and U3880 (N_3880,N_1246,N_1581);
or U3881 (N_3881,N_252,N_637);
and U3882 (N_3882,N_1924,N_807);
and U3883 (N_3883,N_1467,N_662);
or U3884 (N_3884,N_1139,N_1685);
nor U3885 (N_3885,N_1270,N_1352);
or U3886 (N_3886,N_178,N_1590);
nand U3887 (N_3887,N_1459,N_256);
and U3888 (N_3888,N_749,N_418);
nand U3889 (N_3889,N_929,N_918);
or U3890 (N_3890,N_1500,N_1279);
nand U3891 (N_3891,N_325,N_1856);
or U3892 (N_3892,N_1000,N_61);
nand U3893 (N_3893,N_1735,N_1939);
nand U3894 (N_3894,N_832,N_1713);
and U3895 (N_3895,N_1704,N_1249);
and U3896 (N_3896,N_1951,N_249);
and U3897 (N_3897,N_1786,N_1749);
nand U3898 (N_3898,N_1163,N_40);
or U3899 (N_3899,N_124,N_1535);
nand U3900 (N_3900,N_669,N_164);
nor U3901 (N_3901,N_805,N_1910);
nand U3902 (N_3902,N_145,N_862);
and U3903 (N_3903,N_14,N_352);
nand U3904 (N_3904,N_1339,N_68);
nor U3905 (N_3905,N_736,N_940);
and U3906 (N_3906,N_783,N_1536);
nand U3907 (N_3907,N_337,N_13);
nor U3908 (N_3908,N_1577,N_5);
or U3909 (N_3909,N_1940,N_120);
or U3910 (N_3910,N_352,N_814);
or U3911 (N_3911,N_50,N_338);
or U3912 (N_3912,N_1252,N_1682);
nand U3913 (N_3913,N_588,N_1673);
or U3914 (N_3914,N_504,N_542);
nand U3915 (N_3915,N_1355,N_1645);
nor U3916 (N_3916,N_1910,N_472);
nor U3917 (N_3917,N_1183,N_1075);
nand U3918 (N_3918,N_1712,N_984);
or U3919 (N_3919,N_344,N_412);
and U3920 (N_3920,N_1438,N_564);
and U3921 (N_3921,N_1474,N_455);
nand U3922 (N_3922,N_142,N_248);
nor U3923 (N_3923,N_1158,N_913);
nor U3924 (N_3924,N_850,N_74);
nand U3925 (N_3925,N_540,N_33);
nand U3926 (N_3926,N_861,N_1324);
nor U3927 (N_3927,N_1106,N_1836);
nor U3928 (N_3928,N_882,N_1218);
nor U3929 (N_3929,N_390,N_310);
nor U3930 (N_3930,N_1105,N_138);
or U3931 (N_3931,N_482,N_964);
nand U3932 (N_3932,N_381,N_493);
and U3933 (N_3933,N_67,N_130);
xnor U3934 (N_3934,N_1186,N_893);
nor U3935 (N_3935,N_944,N_1506);
nor U3936 (N_3936,N_1861,N_1325);
nor U3937 (N_3937,N_131,N_1911);
nand U3938 (N_3938,N_291,N_229);
nand U3939 (N_3939,N_696,N_594);
nor U3940 (N_3940,N_606,N_421);
xor U3941 (N_3941,N_1747,N_232);
nor U3942 (N_3942,N_546,N_1829);
nor U3943 (N_3943,N_1758,N_1898);
and U3944 (N_3944,N_1557,N_1751);
or U3945 (N_3945,N_1182,N_528);
and U3946 (N_3946,N_707,N_553);
and U3947 (N_3947,N_69,N_709);
or U3948 (N_3948,N_1755,N_645);
nor U3949 (N_3949,N_1155,N_945);
nand U3950 (N_3950,N_1172,N_1671);
nand U3951 (N_3951,N_1889,N_1794);
or U3952 (N_3952,N_1503,N_1938);
and U3953 (N_3953,N_1516,N_1675);
nand U3954 (N_3954,N_1945,N_205);
nand U3955 (N_3955,N_82,N_1705);
nor U3956 (N_3956,N_1320,N_422);
nor U3957 (N_3957,N_1285,N_1170);
nand U3958 (N_3958,N_629,N_332);
nand U3959 (N_3959,N_410,N_1563);
nor U3960 (N_3960,N_1835,N_1334);
and U3961 (N_3961,N_1480,N_1907);
or U3962 (N_3962,N_62,N_1584);
nand U3963 (N_3963,N_1581,N_442);
nand U3964 (N_3964,N_1602,N_1147);
and U3965 (N_3965,N_1745,N_1757);
nand U3966 (N_3966,N_800,N_281);
nor U3967 (N_3967,N_1917,N_1516);
or U3968 (N_3968,N_264,N_1720);
or U3969 (N_3969,N_1039,N_884);
and U3970 (N_3970,N_1281,N_1627);
nand U3971 (N_3971,N_1583,N_190);
and U3972 (N_3972,N_621,N_785);
or U3973 (N_3973,N_611,N_815);
or U3974 (N_3974,N_1516,N_489);
nand U3975 (N_3975,N_1151,N_742);
or U3976 (N_3976,N_1833,N_638);
nor U3977 (N_3977,N_1110,N_1239);
or U3978 (N_3978,N_1692,N_931);
and U3979 (N_3979,N_1839,N_41);
or U3980 (N_3980,N_603,N_1790);
nor U3981 (N_3981,N_501,N_1389);
and U3982 (N_3982,N_946,N_1005);
nor U3983 (N_3983,N_1768,N_402);
nor U3984 (N_3984,N_1061,N_1547);
or U3985 (N_3985,N_719,N_1712);
and U3986 (N_3986,N_210,N_807);
and U3987 (N_3987,N_615,N_1900);
or U3988 (N_3988,N_869,N_182);
and U3989 (N_3989,N_1005,N_812);
and U3990 (N_3990,N_765,N_844);
or U3991 (N_3991,N_541,N_1042);
or U3992 (N_3992,N_812,N_0);
or U3993 (N_3993,N_168,N_1724);
nand U3994 (N_3994,N_1542,N_1788);
or U3995 (N_3995,N_138,N_1180);
nand U3996 (N_3996,N_1900,N_783);
or U3997 (N_3997,N_1496,N_1233);
and U3998 (N_3998,N_438,N_905);
nand U3999 (N_3999,N_1011,N_406);
nor U4000 (N_4000,N_2927,N_3699);
or U4001 (N_4001,N_2808,N_2455);
and U4002 (N_4002,N_2029,N_3879);
or U4003 (N_4003,N_3423,N_2889);
or U4004 (N_4004,N_2350,N_3963);
nor U4005 (N_4005,N_3462,N_3696);
or U4006 (N_4006,N_3992,N_2212);
and U4007 (N_4007,N_3933,N_2098);
nor U4008 (N_4008,N_2088,N_2483);
nand U4009 (N_4009,N_3981,N_3336);
nor U4010 (N_4010,N_2108,N_3072);
or U4011 (N_4011,N_3746,N_3216);
and U4012 (N_4012,N_3431,N_2067);
and U4013 (N_4013,N_3800,N_3526);
xnor U4014 (N_4014,N_2140,N_2886);
nor U4015 (N_4015,N_3536,N_2295);
xnor U4016 (N_4016,N_2262,N_3817);
nand U4017 (N_4017,N_3109,N_3138);
nand U4018 (N_4018,N_3183,N_3214);
nand U4019 (N_4019,N_3913,N_3795);
and U4020 (N_4020,N_2096,N_3297);
nand U4021 (N_4021,N_2965,N_3627);
or U4022 (N_4022,N_3157,N_3130);
and U4023 (N_4023,N_2118,N_2122);
nand U4024 (N_4024,N_3483,N_3167);
or U4025 (N_4025,N_2534,N_2837);
nor U4026 (N_4026,N_3146,N_2620);
nand U4027 (N_4027,N_2637,N_3465);
nand U4028 (N_4028,N_3801,N_3751);
nand U4029 (N_4029,N_2725,N_2780);
nand U4030 (N_4030,N_3281,N_3850);
nand U4031 (N_4031,N_3613,N_2908);
nor U4032 (N_4032,N_3286,N_2244);
nor U4033 (N_4033,N_2762,N_2080);
or U4034 (N_4034,N_3032,N_2922);
nand U4035 (N_4035,N_3652,N_2025);
or U4036 (N_4036,N_2665,N_3796);
and U4037 (N_4037,N_2175,N_2801);
and U4038 (N_4038,N_2659,N_2042);
nand U4039 (N_4039,N_3532,N_2806);
or U4040 (N_4040,N_3759,N_3365);
and U4041 (N_4041,N_2490,N_2256);
and U4042 (N_4042,N_2263,N_2103);
nand U4043 (N_4043,N_3397,N_3371);
nor U4044 (N_4044,N_2905,N_2340);
or U4045 (N_4045,N_3271,N_2346);
and U4046 (N_4046,N_2440,N_3260);
nand U4047 (N_4047,N_2744,N_2773);
or U4048 (N_4048,N_2882,N_3961);
nor U4049 (N_4049,N_3847,N_3680);
nor U4050 (N_4050,N_2273,N_3363);
nor U4051 (N_4051,N_2537,N_3623);
nor U4052 (N_4052,N_3421,N_2997);
nor U4053 (N_4053,N_2297,N_3047);
or U4054 (N_4054,N_2960,N_2125);
nand U4055 (N_4055,N_3055,N_2131);
nand U4056 (N_4056,N_3201,N_3313);
nand U4057 (N_4057,N_2755,N_2944);
and U4058 (N_4058,N_3486,N_3162);
nor U4059 (N_4059,N_2402,N_2688);
or U4060 (N_4060,N_3856,N_3059);
or U4061 (N_4061,N_2290,N_2929);
or U4062 (N_4062,N_2028,N_2609);
or U4063 (N_4063,N_3975,N_3158);
and U4064 (N_4064,N_2251,N_3422);
and U4065 (N_4065,N_2723,N_2472);
nand U4066 (N_4066,N_2893,N_3539);
and U4067 (N_4067,N_2265,N_3663);
nand U4068 (N_4068,N_3579,N_2660);
and U4069 (N_4069,N_2648,N_2538);
or U4070 (N_4070,N_3614,N_3448);
nand U4071 (N_4071,N_3775,N_3124);
nor U4072 (N_4072,N_3394,N_3892);
nand U4073 (N_4073,N_3122,N_2159);
and U4074 (N_4074,N_2686,N_3996);
and U4075 (N_4075,N_2985,N_3487);
nor U4076 (N_4076,N_2489,N_3332);
or U4077 (N_4077,N_3156,N_2511);
or U4078 (N_4078,N_3435,N_3895);
or U4079 (N_4079,N_2014,N_3776);
nor U4080 (N_4080,N_3247,N_3596);
or U4081 (N_4081,N_3338,N_2287);
nor U4082 (N_4082,N_3301,N_3037);
and U4083 (N_4083,N_3459,N_2570);
and U4084 (N_4084,N_2624,N_3026);
and U4085 (N_4085,N_3269,N_3238);
nand U4086 (N_4086,N_2520,N_3855);
or U4087 (N_4087,N_3973,N_2388);
nor U4088 (N_4088,N_3711,N_3098);
nand U4089 (N_4089,N_3867,N_2890);
and U4090 (N_4090,N_3656,N_3246);
and U4091 (N_4091,N_3919,N_3331);
or U4092 (N_4092,N_2249,N_3950);
or U4093 (N_4093,N_3102,N_2493);
nand U4094 (N_4094,N_2496,N_3642);
nand U4095 (N_4095,N_3608,N_2216);
and U4096 (N_4096,N_3785,N_3419);
nor U4097 (N_4097,N_3547,N_2284);
xnor U4098 (N_4098,N_2236,N_3993);
nand U4099 (N_4099,N_2454,N_2474);
xnor U4100 (N_4100,N_3083,N_3794);
and U4101 (N_4101,N_2794,N_2279);
nand U4102 (N_4102,N_3706,N_2091);
and U4103 (N_4103,N_2195,N_3306);
or U4104 (N_4104,N_2319,N_3921);
nand U4105 (N_4105,N_2838,N_3144);
nand U4106 (N_4106,N_3493,N_3900);
or U4107 (N_4107,N_2250,N_3779);
and U4108 (N_4108,N_3094,N_3510);
nand U4109 (N_4109,N_2618,N_2583);
and U4110 (N_4110,N_2733,N_2895);
nor U4111 (N_4111,N_2711,N_3418);
or U4112 (N_4112,N_2527,N_3215);
and U4113 (N_4113,N_3182,N_3282);
nor U4114 (N_4114,N_2649,N_2348);
or U4115 (N_4115,N_2689,N_3834);
and U4116 (N_4116,N_2463,N_2937);
nand U4117 (N_4117,N_3770,N_3545);
nor U4118 (N_4118,N_3716,N_2602);
nand U4119 (N_4119,N_3385,N_3844);
and U4120 (N_4120,N_2010,N_3780);
nand U4121 (N_4121,N_2831,N_3113);
nand U4122 (N_4122,N_3771,N_3799);
nor U4123 (N_4123,N_3004,N_3342);
nand U4124 (N_4124,N_2399,N_2062);
and U4125 (N_4125,N_3988,N_2207);
and U4126 (N_4126,N_2215,N_3087);
and U4127 (N_4127,N_2549,N_2741);
nor U4128 (N_4128,N_3051,N_2541);
nand U4129 (N_4129,N_3831,N_2656);
and U4130 (N_4130,N_2529,N_3858);
nand U4131 (N_4131,N_3236,N_2226);
nor U4132 (N_4132,N_2799,N_2781);
and U4133 (N_4133,N_2850,N_3965);
nor U4134 (N_4134,N_2083,N_3703);
nor U4135 (N_4135,N_2685,N_2591);
and U4136 (N_4136,N_3432,N_3184);
or U4137 (N_4137,N_2151,N_2242);
nand U4138 (N_4138,N_2726,N_2971);
or U4139 (N_4139,N_2338,N_2724);
nor U4140 (N_4140,N_2015,N_2961);
and U4141 (N_4141,N_3626,N_2593);
nor U4142 (N_4142,N_3581,N_3350);
and U4143 (N_4143,N_3505,N_2912);
nor U4144 (N_4144,N_2757,N_3232);
and U4145 (N_4145,N_2045,N_3682);
or U4146 (N_4146,N_2381,N_2863);
and U4147 (N_4147,N_3388,N_2401);
or U4148 (N_4148,N_2243,N_3253);
or U4149 (N_4149,N_2238,N_2946);
and U4150 (N_4150,N_2819,N_2524);
nand U4151 (N_4151,N_2482,N_3689);
or U4152 (N_4152,N_2606,N_2146);
nand U4153 (N_4153,N_2331,N_3212);
nor U4154 (N_4154,N_3120,N_3669);
or U4155 (N_4155,N_3335,N_2460);
nand U4156 (N_4156,N_2953,N_2547);
nand U4157 (N_4157,N_2434,N_3748);
or U4158 (N_4158,N_2873,N_2704);
nor U4159 (N_4159,N_2322,N_3035);
nor U4160 (N_4160,N_2261,N_3005);
and U4161 (N_4161,N_2558,N_2132);
or U4162 (N_4162,N_2707,N_3570);
nand U4163 (N_4163,N_2239,N_3381);
or U4164 (N_4164,N_2608,N_3242);
and U4165 (N_4165,N_2866,N_2750);
and U4166 (N_4166,N_2364,N_2170);
nor U4167 (N_4167,N_3139,N_3828);
nand U4168 (N_4168,N_2019,N_2793);
and U4169 (N_4169,N_3861,N_2258);
and U4170 (N_4170,N_3500,N_3274);
nand U4171 (N_4171,N_3029,N_3808);
and U4172 (N_4172,N_3071,N_3323);
or U4173 (N_4173,N_3966,N_2502);
nand U4174 (N_4174,N_3885,N_2877);
nand U4175 (N_4175,N_3792,N_2567);
nor U4176 (N_4176,N_3722,N_3538);
and U4177 (N_4177,N_2840,N_3129);
and U4178 (N_4178,N_2610,N_2016);
or U4179 (N_4179,N_2335,N_3901);
or U4180 (N_4180,N_3890,N_3117);
nand U4181 (N_4181,N_3709,N_2803);
or U4182 (N_4182,N_3470,N_2975);
or U4183 (N_4183,N_3293,N_3906);
and U4184 (N_4184,N_2945,N_2134);
or U4185 (N_4185,N_2257,N_3445);
nor U4186 (N_4186,N_2625,N_2836);
nor U4187 (N_4187,N_2714,N_3079);
nand U4188 (N_4188,N_3307,N_2457);
nand U4189 (N_4189,N_2821,N_2275);
nand U4190 (N_4190,N_3220,N_2420);
and U4191 (N_4191,N_2491,N_2484);
nor U4192 (N_4192,N_3917,N_3284);
or U4193 (N_4193,N_2375,N_2136);
nor U4194 (N_4194,N_2772,N_2081);
nor U4195 (N_4195,N_2109,N_2693);
nor U4196 (N_4196,N_3252,N_3718);
and U4197 (N_4197,N_3628,N_2931);
and U4198 (N_4198,N_3620,N_2674);
nor U4199 (N_4199,N_3469,N_3386);
and U4200 (N_4200,N_3761,N_3686);
or U4201 (N_4201,N_2052,N_2349);
nand U4202 (N_4202,N_3121,N_3474);
and U4203 (N_4203,N_3401,N_2951);
nor U4204 (N_4204,N_3936,N_3108);
nor U4205 (N_4205,N_2954,N_3409);
nor U4206 (N_4206,N_2106,N_3560);
or U4207 (N_4207,N_3968,N_3104);
and U4208 (N_4208,N_3278,N_2892);
nand U4209 (N_4209,N_2414,N_3592);
and U4210 (N_4210,N_3151,N_2470);
and U4211 (N_4211,N_2386,N_3967);
nand U4212 (N_4212,N_2814,N_3352);
nand U4213 (N_4213,N_2763,N_2069);
or U4214 (N_4214,N_3272,N_2544);
and U4215 (N_4215,N_3612,N_3233);
nor U4216 (N_4216,N_3179,N_3717);
nand U4217 (N_4217,N_2993,N_2580);
nand U4218 (N_4218,N_2980,N_2355);
or U4219 (N_4219,N_2037,N_2650);
nor U4220 (N_4220,N_2669,N_2400);
or U4221 (N_4221,N_2044,N_2681);
nand U4222 (N_4222,N_2237,N_2252);
xnor U4223 (N_4223,N_3499,N_2049);
nand U4224 (N_4224,N_3577,N_2370);
and U4225 (N_4225,N_3725,N_3768);
and U4226 (N_4226,N_3877,N_2079);
and U4227 (N_4227,N_2556,N_3078);
or U4228 (N_4228,N_3617,N_2839);
or U4229 (N_4229,N_3829,N_3523);
nand U4230 (N_4230,N_2309,N_3513);
or U4231 (N_4231,N_2754,N_2783);
xor U4232 (N_4232,N_2898,N_3142);
or U4233 (N_4233,N_3887,N_3664);
nand U4234 (N_4234,N_2816,N_3390);
and U4235 (N_4235,N_2588,N_2706);
nand U4236 (N_4236,N_2712,N_2043);
nor U4237 (N_4237,N_2532,N_2915);
nand U4238 (N_4238,N_2802,N_2135);
or U4239 (N_4239,N_2771,N_3466);
nand U4240 (N_4240,N_2156,N_2976);
and U4241 (N_4241,N_3020,N_3683);
or U4242 (N_4242,N_2565,N_3195);
nand U4243 (N_4243,N_2790,N_3145);
nor U4244 (N_4244,N_2202,N_2767);
nand U4245 (N_4245,N_3197,N_3046);
or U4246 (N_4246,N_3629,N_2487);
or U4247 (N_4247,N_2746,N_2942);
nor U4248 (N_4248,N_3865,N_3165);
and U4249 (N_4249,N_3727,N_2110);
and U4250 (N_4250,N_2306,N_3672);
nor U4251 (N_4251,N_3149,N_2291);
or U4252 (N_4252,N_2872,N_3349);
and U4253 (N_4253,N_2183,N_2813);
nor U4254 (N_4254,N_3533,N_3908);
and U4255 (N_4255,N_2281,N_2901);
nand U4256 (N_4256,N_2046,N_2345);
and U4257 (N_4257,N_2531,N_3852);
and U4258 (N_4258,N_3943,N_3011);
nor U4259 (N_4259,N_3033,N_3690);
nor U4260 (N_4260,N_2476,N_2318);
or U4261 (N_4261,N_2023,N_2030);
xor U4262 (N_4262,N_3075,N_3827);
nand U4263 (N_4263,N_2259,N_2005);
and U4264 (N_4264,N_2418,N_3235);
nand U4265 (N_4265,N_3695,N_2533);
or U4266 (N_4266,N_2479,N_3942);
nor U4267 (N_4267,N_3436,N_2939);
nand U4268 (N_4268,N_2353,N_2779);
nand U4269 (N_4269,N_3633,N_2990);
nor U4270 (N_4270,N_2357,N_2050);
and U4271 (N_4271,N_3554,N_2933);
nand U4272 (N_4272,N_2234,N_3911);
and U4273 (N_4273,N_3366,N_2546);
nor U4274 (N_4274,N_3137,N_2094);
or U4275 (N_4275,N_3140,N_3555);
nor U4276 (N_4276,N_3914,N_3954);
nor U4277 (N_4277,N_2329,N_3518);
nor U4278 (N_4278,N_2424,N_3873);
nor U4279 (N_4279,N_2209,N_2646);
nand U4280 (N_4280,N_2930,N_2983);
or U4281 (N_4281,N_3168,N_3128);
nand U4282 (N_4282,N_3076,N_2371);
or U4283 (N_4283,N_3638,N_3008);
nand U4284 (N_4284,N_3084,N_3553);
or U4285 (N_4285,N_3881,N_3791);
xor U4286 (N_4286,N_3821,N_2989);
and U4287 (N_4287,N_3684,N_2006);
and U4288 (N_4288,N_2661,N_2663);
or U4289 (N_4289,N_3659,N_2341);
xor U4290 (N_4290,N_3781,N_2920);
nor U4291 (N_4291,N_3615,N_3417);
nand U4292 (N_4292,N_2086,N_3199);
xnor U4293 (N_4293,N_2114,N_3039);
nand U4294 (N_4294,N_2708,N_3316);
nand U4295 (N_4295,N_3893,N_3951);
or U4296 (N_4296,N_2283,N_2488);
nand U4297 (N_4297,N_2582,N_2737);
nor U4298 (N_4298,N_3442,N_3223);
nand U4299 (N_4299,N_2766,N_3645);
or U4300 (N_4300,N_2082,N_2720);
nand U4301 (N_4301,N_3647,N_2126);
nand U4302 (N_4302,N_3089,N_3133);
nand U4303 (N_4303,N_3732,N_3279);
or U4304 (N_4304,N_3876,N_3840);
nand U4305 (N_4305,N_3757,N_3986);
or U4306 (N_4306,N_3820,N_3014);
or U4307 (N_4307,N_3670,N_2760);
nor U4308 (N_4308,N_2959,N_3790);
nand U4309 (N_4309,N_2880,N_2092);
or U4310 (N_4310,N_3502,N_3531);
nor U4311 (N_4311,N_2730,N_2373);
nor U4312 (N_4312,N_2260,N_2087);
or U4313 (N_4313,N_2224,N_2492);
and U4314 (N_4314,N_3926,N_3164);
nor U4315 (N_4315,N_3481,N_2495);
nor U4316 (N_4316,N_2431,N_3042);
xor U4317 (N_4317,N_3327,N_3530);
or U4318 (N_4318,N_2991,N_3760);
nor U4319 (N_4319,N_2825,N_2498);
or U4320 (N_4320,N_2964,N_2382);
xor U4321 (N_4321,N_3754,N_2557);
or U4322 (N_4322,N_3472,N_3292);
or U4323 (N_4323,N_3974,N_3163);
or U4324 (N_4324,N_3549,N_3863);
or U4325 (N_4325,N_2826,N_2060);
nor U4326 (N_4326,N_3449,N_3243);
nand U4327 (N_4327,N_2143,N_2392);
and U4328 (N_4328,N_2447,N_3728);
and U4329 (N_4329,N_3275,N_2519);
nand U4330 (N_4330,N_3362,N_2769);
and U4331 (N_4331,N_2503,N_3310);
or U4332 (N_4332,N_2078,N_3333);
nor U4333 (N_4333,N_3221,N_3050);
or U4334 (N_4334,N_3907,N_3949);
and U4335 (N_4335,N_3063,N_2830);
or U4336 (N_4336,N_3685,N_2363);
nand U4337 (N_4337,N_2138,N_3657);
nand U4338 (N_4338,N_2102,N_2336);
nor U4339 (N_4339,N_3229,N_2996);
nand U4340 (N_4340,N_2459,N_2627);
or U4341 (N_4341,N_2128,N_2032);
or U4342 (N_4342,N_2633,N_2137);
or U4343 (N_4343,N_2026,N_3028);
nor U4344 (N_4344,N_3681,N_3372);
nor U4345 (N_4345,N_2415,N_3111);
and U4346 (N_4346,N_2906,N_2594);
and U4347 (N_4347,N_3290,N_3302);
nor U4348 (N_4348,N_3240,N_2184);
nand U4349 (N_4349,N_3583,N_3648);
or U4350 (N_4350,N_3103,N_3153);
nand U4351 (N_4351,N_2747,N_2792);
nor U4352 (N_4352,N_2304,N_3482);
and U4353 (N_4353,N_2426,N_2849);
or U4354 (N_4354,N_3070,N_3096);
or U4355 (N_4355,N_2148,N_3254);
nor U4356 (N_4356,N_2918,N_2982);
nor U4357 (N_4357,N_3793,N_3248);
and U4358 (N_4358,N_3068,N_2584);
nand U4359 (N_4359,N_2378,N_2333);
and U4360 (N_4360,N_2278,N_2073);
nand U4361 (N_4361,N_3957,N_3994);
nor U4362 (N_4362,N_2913,N_3131);
or U4363 (N_4363,N_2542,N_3213);
nor U4364 (N_4364,N_2956,N_2181);
nor U4365 (N_4365,N_3489,N_3360);
nand U4366 (N_4366,N_3081,N_3920);
nand U4367 (N_4367,N_2694,N_3172);
nand U4368 (N_4368,N_3517,N_2116);
or U4369 (N_4369,N_2323,N_3446);
or U4370 (N_4370,N_2411,N_3619);
nor U4371 (N_4371,N_3319,N_2123);
or U4372 (N_4372,N_3389,N_3516);
or U4373 (N_4373,N_3527,N_2478);
and U4374 (N_4374,N_2652,N_3180);
nor U4375 (N_4375,N_2450,N_3773);
or U4376 (N_4376,N_3479,N_3255);
and U4377 (N_4377,N_3878,N_2815);
or U4378 (N_4378,N_3267,N_3208);
or U4379 (N_4379,N_3875,N_3705);
nor U4380 (N_4380,N_3447,N_2743);
and U4381 (N_4381,N_3762,N_3640);
and U4382 (N_4382,N_3196,N_2395);
or U4383 (N_4383,N_2267,N_3374);
nor U4384 (N_4384,N_2332,N_2651);
or U4385 (N_4385,N_2903,N_3105);
and U4386 (N_4386,N_2528,N_3378);
or U4387 (N_4387,N_3057,N_3610);
and U4388 (N_4388,N_3230,N_2630);
or U4389 (N_4389,N_2093,N_2327);
and U4390 (N_4390,N_2421,N_3224);
and U4391 (N_4391,N_3529,N_2210);
nor U4392 (N_4392,N_3354,N_2384);
and U4393 (N_4393,N_3507,N_3200);
and U4394 (N_4394,N_2469,N_3406);
and U4395 (N_4395,N_3673,N_3148);
or U4396 (N_4396,N_2233,N_2921);
and U4397 (N_4397,N_3691,N_3118);
nand U4398 (N_4398,N_2999,N_2786);
and U4399 (N_4399,N_3774,N_2505);
and U4400 (N_4400,N_3136,N_2040);
nor U4401 (N_4401,N_2330,N_3107);
nor U4402 (N_4402,N_3152,N_3999);
nand U4403 (N_4403,N_2687,N_3514);
nor U4404 (N_4404,N_2775,N_2853);
nor U4405 (N_4405,N_3763,N_3150);
nand U4406 (N_4406,N_3928,N_2798);
and U4407 (N_4407,N_2645,N_3600);
nand U4408 (N_4408,N_3842,N_2286);
nor U4409 (N_4409,N_3185,N_2604);
or U4410 (N_4410,N_2623,N_2899);
nor U4411 (N_4411,N_3739,N_3439);
and U4412 (N_4412,N_2870,N_2578);
or U4413 (N_4413,N_3740,N_2288);
or U4414 (N_4414,N_2867,N_3484);
or U4415 (N_4415,N_3326,N_3512);
nor U4416 (N_4416,N_2406,N_3896);
nor U4417 (N_4417,N_3702,N_2680);
or U4418 (N_4418,N_2589,N_3015);
nand U4419 (N_4419,N_2884,N_2752);
and U4420 (N_4420,N_2075,N_3341);
xor U4421 (N_4421,N_3368,N_2676);
nand U4422 (N_4422,N_3041,N_2177);
nand U4423 (N_4423,N_2955,N_2012);
or U4424 (N_4424,N_3524,N_2590);
nand U4425 (N_4425,N_2429,N_2343);
nand U4426 (N_4426,N_3375,N_2229);
or U4427 (N_4427,N_2756,N_2142);
and U4428 (N_4428,N_3766,N_3457);
and U4429 (N_4429,N_2316,N_3730);
and U4430 (N_4430,N_3591,N_2448);
or U4431 (N_4431,N_2227,N_2809);
nand U4432 (N_4432,N_3707,N_3601);
nor U4433 (N_4433,N_3383,N_3067);
and U4434 (N_4434,N_2344,N_3053);
nand U4435 (N_4435,N_2410,N_3045);
nor U4436 (N_4436,N_2059,N_3080);
nand U4437 (N_4437,N_2857,N_3427);
or U4438 (N_4438,N_3723,N_3285);
and U4439 (N_4439,N_3241,N_2936);
and U4440 (N_4440,N_2439,N_3305);
nand U4441 (N_4441,N_3458,N_2719);
or U4442 (N_4442,N_2888,N_3810);
nand U4443 (N_4443,N_2246,N_2540);
or U4444 (N_4444,N_3376,N_3295);
nor U4445 (N_4445,N_2198,N_3049);
or U4446 (N_4446,N_3115,N_3983);
nand U4447 (N_4447,N_2186,N_2453);
and U4448 (N_4448,N_3328,N_2807);
nand U4449 (N_4449,N_3298,N_2515);
nand U4450 (N_4450,N_2805,N_3693);
and U4451 (N_4451,N_2876,N_2764);
nand U4452 (N_4452,N_3724,N_3915);
nor U4453 (N_4453,N_2058,N_3463);
and U4454 (N_4454,N_3424,N_2366);
nor U4455 (N_4455,N_2709,N_3219);
and U4456 (N_4456,N_3337,N_3937);
nand U4457 (N_4457,N_3320,N_3597);
nor U4458 (N_4458,N_3309,N_2387);
or U4459 (N_4459,N_2768,N_2220);
nor U4460 (N_4460,N_2810,N_2626);
or U4461 (N_4461,N_2471,N_2302);
nand U4462 (N_4462,N_3783,N_3273);
or U4463 (N_4463,N_3343,N_3634);
nor U4464 (N_4464,N_2413,N_2940);
nor U4465 (N_4465,N_2765,N_3927);
nand U4466 (N_4466,N_3537,N_3490);
and U4467 (N_4467,N_2612,N_2716);
and U4468 (N_4468,N_2161,N_2280);
nand U4469 (N_4469,N_3382,N_3351);
and U4470 (N_4470,N_2662,N_3169);
nand U4471 (N_4471,N_2268,N_3270);
nand U4472 (N_4472,N_3398,N_3916);
nand U4473 (N_4473,N_2169,N_2616);
and U4474 (N_4474,N_2848,N_2981);
nand U4475 (N_4475,N_2587,N_3441);
or U4476 (N_4476,N_2317,N_2509);
nor U4477 (N_4477,N_3329,N_2368);
nor U4478 (N_4478,N_3340,N_3317);
nor U4479 (N_4479,N_2966,N_3891);
or U4480 (N_4480,N_3013,N_3772);
and U4481 (N_4481,N_3888,N_2120);
nand U4482 (N_4482,N_3346,N_2254);
and U4483 (N_4483,N_3520,N_3123);
nor U4484 (N_4484,N_3007,N_2718);
xnor U4485 (N_4485,N_2666,N_2947);
nor U4486 (N_4486,N_3979,N_2795);
or U4487 (N_4487,N_3789,N_3859);
or U4488 (N_4488,N_3807,N_2352);
or U4489 (N_4489,N_2225,N_3226);
nor U4490 (N_4490,N_3618,N_3173);
or U4491 (N_4491,N_3835,N_2844);
nand U4492 (N_4492,N_3939,N_2064);
nand U4493 (N_4493,N_3719,N_3978);
and U4494 (N_4494,N_3426,N_3589);
and U4495 (N_4495,N_2354,N_3704);
and U4496 (N_4496,N_2222,N_2577);
or U4497 (N_4497,N_2213,N_3948);
nor U4498 (N_4498,N_3824,N_2068);
or U4499 (N_4499,N_3712,N_2512);
nand U4500 (N_4500,N_2791,N_3959);
or U4501 (N_4501,N_3575,N_3822);
nand U4502 (N_4502,N_3621,N_2938);
and U4503 (N_4503,N_2811,N_3189);
nand U4504 (N_4504,N_3982,N_2444);
nor U4505 (N_4505,N_3956,N_3303);
nand U4506 (N_4506,N_2066,N_3752);
nor U4507 (N_4507,N_3519,N_3373);
nor U4508 (N_4508,N_2530,N_2314);
or U4509 (N_4509,N_3475,N_3631);
or U4510 (N_4510,N_2745,N_2449);
and U4511 (N_4511,N_3909,N_3412);
or U4512 (N_4512,N_3116,N_3980);
nand U4513 (N_4513,N_2562,N_2008);
nand U4514 (N_4514,N_3665,N_2145);
nor U4515 (N_4515,N_2581,N_3453);
nor U4516 (N_4516,N_2740,N_2510);
or U4517 (N_4517,N_3677,N_2232);
nand U4518 (N_4518,N_3522,N_2405);
and U4519 (N_4519,N_2804,N_2300);
nand U4520 (N_4520,N_2822,N_3866);
xnor U4521 (N_4521,N_2168,N_3987);
nor U4522 (N_4522,N_3905,N_2572);
and U4523 (N_4523,N_3886,N_3225);
and U4524 (N_4524,N_3099,N_3100);
and U4525 (N_4525,N_2334,N_3676);
nor U4526 (N_4526,N_3603,N_2228);
nand U4527 (N_4527,N_3440,N_3995);
nand U4528 (N_4528,N_3300,N_2173);
nand U4529 (N_4529,N_2879,N_2596);
and U4530 (N_4530,N_2231,N_3085);
or U4531 (N_4531,N_2513,N_3477);
and U4532 (N_4532,N_3357,N_2568);
or U4533 (N_4533,N_2869,N_3324);
or U4534 (N_4534,N_3880,N_2605);
nand U4535 (N_4535,N_3806,N_3141);
or U4536 (N_4536,N_3315,N_2535);
or U4537 (N_4537,N_3000,N_3438);
or U4538 (N_4538,N_2180,N_2036);
and U4539 (N_4539,N_2600,N_3869);
or U4540 (N_4540,N_3587,N_2221);
and U4541 (N_4541,N_2705,N_3204);
nand U4542 (N_4542,N_2241,N_2855);
or U4543 (N_4543,N_2313,N_3234);
or U4544 (N_4544,N_2099,N_3125);
or U4545 (N_4545,N_3984,N_3093);
nor U4546 (N_4546,N_2285,N_3239);
nand U4547 (N_4547,N_2007,N_3720);
nand U4548 (N_4548,N_2270,N_2298);
nor U4549 (N_4549,N_2729,N_3002);
and U4550 (N_4550,N_3870,N_3434);
and U4551 (N_4551,N_2928,N_3661);
nand U4552 (N_4552,N_2409,N_3653);
or U4553 (N_4553,N_2129,N_2619);
nor U4554 (N_4554,N_2009,N_3334);
and U4555 (N_4555,N_3468,N_2571);
nand U4556 (N_4556,N_2742,N_3650);
or U4557 (N_4557,N_3250,N_3461);
or U4558 (N_4558,N_3803,N_2292);
nor U4559 (N_4559,N_3548,N_3668);
nand U4560 (N_4560,N_2022,N_2564);
and U4561 (N_4561,N_3485,N_3060);
and U4562 (N_4562,N_2678,N_3062);
or U4563 (N_4563,N_3192,N_3710);
nor U4564 (N_4564,N_3450,N_3864);
and U4565 (N_4565,N_2289,N_2559);
nor U4566 (N_4566,N_2201,N_2647);
and U4567 (N_4567,N_2759,N_2230);
and U4568 (N_4568,N_3494,N_2628);
and U4569 (N_4569,N_3454,N_3506);
or U4570 (N_4570,N_3700,N_3871);
or U4571 (N_4571,N_2601,N_2035);
nor U4572 (N_4572,N_3654,N_2374);
and U4573 (N_4573,N_2248,N_2501);
or U4574 (N_4574,N_2033,N_3912);
nand U4575 (N_4575,N_2379,N_2365);
nand U4576 (N_4576,N_3813,N_2218);
and U4577 (N_4577,N_3787,N_2900);
nor U4578 (N_4578,N_2885,N_3001);
nand U4579 (N_4579,N_2321,N_2607);
nand U4580 (N_4580,N_2165,N_2774);
and U4581 (N_4581,N_2778,N_3862);
and U4582 (N_4582,N_3283,N_3798);
and U4583 (N_4583,N_3321,N_2521);
nand U4584 (N_4584,N_3480,N_2446);
nand U4585 (N_4585,N_3637,N_2917);
nor U4586 (N_4586,N_2518,N_3742);
nand U4587 (N_4587,N_2090,N_3646);
and U4588 (N_4588,N_3599,N_3017);
nand U4589 (N_4589,N_2728,N_3392);
and U4590 (N_4590,N_3266,N_3127);
or U4591 (N_4591,N_3433,N_3814);
nand U4592 (N_4592,N_3585,N_2301);
or U4593 (N_4593,N_3582,N_2902);
nand U4594 (N_4594,N_2308,N_2970);
nand U4595 (N_4595,N_3359,N_2700);
or U4596 (N_4596,N_2957,N_3802);
or U4597 (N_4597,N_2673,N_3218);
nor U4598 (N_4598,N_3291,N_3171);
and U4599 (N_4599,N_2315,N_3198);
or U4600 (N_4600,N_2253,N_3643);
nand U4601 (N_4601,N_3367,N_2638);
and U4602 (N_4602,N_2174,N_3030);
and U4603 (N_4603,N_3402,N_3764);
nor U4604 (N_4604,N_2155,N_3540);
or U4605 (N_4605,N_3733,N_3399);
nor U4606 (N_4606,N_3625,N_2682);
or U4607 (N_4607,N_2896,N_2051);
or U4608 (N_4608,N_3588,N_2130);
and U4609 (N_4609,N_2787,N_3058);
or U4610 (N_4610,N_2111,N_2749);
nand U4611 (N_4611,N_3938,N_2948);
nand U4612 (N_4612,N_2962,N_2061);
nand U4613 (N_4613,N_2425,N_3280);
or U4614 (N_4614,N_2144,N_3541);
or U4615 (N_4615,N_2690,N_3175);
nor U4616 (N_4616,N_2024,N_2897);
and U4617 (N_4617,N_3159,N_3649);
or U4618 (N_4618,N_3052,N_2149);
or U4619 (N_4619,N_2859,N_2191);
nor U4620 (N_4620,N_2085,N_3767);
or U4621 (N_4621,N_2466,N_2271);
and U4622 (N_4622,N_3430,N_2435);
nor U4623 (N_4623,N_2621,N_2194);
and U4624 (N_4624,N_2018,N_3155);
and U4625 (N_4625,N_3651,N_2133);
nor U4626 (N_4626,N_3040,N_2824);
nor U4627 (N_4627,N_3688,N_2214);
or U4628 (N_4628,N_3955,N_3176);
and U4629 (N_4629,N_2188,N_3964);
or U4630 (N_4630,N_3202,N_2555);
or U4631 (N_4631,N_3816,N_2785);
and U4632 (N_4632,N_3091,N_3503);
or U4633 (N_4633,N_2823,N_2179);
nor U4634 (N_4634,N_2397,N_2039);
or U4635 (N_4635,N_2858,N_2834);
nor U4636 (N_4636,N_2671,N_2445);
and U4637 (N_4637,N_3747,N_2545);
and U4638 (N_4638,N_2910,N_2963);
nor U4639 (N_4639,N_2995,N_2097);
or U4640 (N_4640,N_3846,N_2390);
or U4641 (N_4641,N_3393,N_3925);
or U4642 (N_4642,N_2784,N_2176);
and U4643 (N_4643,N_2679,N_2441);
and U4644 (N_4644,N_3404,N_3788);
nor U4645 (N_4645,N_2727,N_2100);
nor U4646 (N_4646,N_2702,N_2312);
or U4647 (N_4647,N_2211,N_2843);
nand U4648 (N_4648,N_2011,N_2603);
and U4649 (N_4649,N_3003,N_3542);
and U4650 (N_4650,N_2820,N_2196);
or U4651 (N_4651,N_3838,N_3743);
nor U4652 (N_4652,N_2699,N_3826);
nand U4653 (N_4653,N_2423,N_2452);
nand U4654 (N_4654,N_2561,N_3132);
and U4655 (N_4655,N_3410,N_3391);
nor U4656 (N_4656,N_3990,N_3777);
nor U4657 (N_4657,N_2480,N_2428);
and U4658 (N_4658,N_3515,N_2860);
nor U4659 (N_4659,N_3194,N_3674);
or U4660 (N_4660,N_2171,N_3923);
or U4661 (N_4661,N_3845,N_2883);
or U4662 (N_4662,N_3737,N_2691);
nor U4663 (N_4663,N_3413,N_3977);
nor U4664 (N_4664,N_2266,N_2828);
nor U4665 (N_4665,N_3188,N_2632);
or U4666 (N_4666,N_2077,N_2552);
nand U4667 (N_4667,N_3191,N_3687);
or U4668 (N_4668,N_2851,N_2695);
nand U4669 (N_4669,N_2736,N_3174);
nor U4670 (N_4670,N_2703,N_3797);
nand U4671 (N_4671,N_3495,N_2433);
nand U4672 (N_4672,N_3209,N_2294);
and U4673 (N_4673,N_2788,N_3947);
nor U4674 (N_4674,N_2634,N_2655);
nor U4675 (N_4675,N_2115,N_2597);
nand U4676 (N_4676,N_3698,N_3641);
or U4677 (N_4677,N_3666,N_2548);
or U4678 (N_4678,N_3786,N_3380);
nor U4679 (N_4679,N_3556,N_3066);
nor U4680 (N_4680,N_3325,N_3217);
nor U4681 (N_4681,N_3578,N_2832);
or U4682 (N_4682,N_3395,N_3244);
nand U4683 (N_4683,N_2310,N_3935);
or U4684 (N_4684,N_3187,N_3312);
nor U4685 (N_4685,N_3428,N_3511);
and U4686 (N_4686,N_3736,N_2984);
nand U4687 (N_4687,N_2987,N_3501);
and U4688 (N_4688,N_3848,N_2299);
or U4689 (N_4689,N_3090,N_2124);
and U4690 (N_4690,N_2941,N_2675);
or U4691 (N_4691,N_3504,N_2777);
nor U4692 (N_4692,N_2560,N_3566);
and U4693 (N_4693,N_2670,N_2383);
or U4694 (N_4694,N_3114,N_3289);
nand U4695 (N_4695,N_2868,N_3384);
nor U4696 (N_4696,N_2430,N_2084);
nand U4697 (N_4697,N_2543,N_3941);
and U4698 (N_4698,N_2972,N_3815);
nand U4699 (N_4699,N_2398,N_2551);
nor U4700 (N_4700,N_2553,N_3211);
nor U4701 (N_4701,N_2739,N_2573);
and U4702 (N_4702,N_3958,N_2197);
and U4703 (N_4703,N_3205,N_2141);
nand U4704 (N_4704,N_3154,N_2157);
nand U4705 (N_4705,N_2911,N_3177);
nor U4706 (N_4706,N_2361,N_2127);
nand U4707 (N_4707,N_3231,N_3353);
or U4708 (N_4708,N_3809,N_3658);
or U4709 (N_4709,N_3662,N_2121);
nor U4710 (N_4710,N_3488,N_2968);
and U4711 (N_4711,N_2481,N_2852);
nand U4712 (N_4712,N_3819,N_2154);
or U4713 (N_4713,N_3952,N_3632);
or U4714 (N_4714,N_3715,N_3407);
or U4715 (N_4715,N_2874,N_3110);
or U4716 (N_4716,N_3135,N_2376);
nor U4717 (N_4717,N_3679,N_2697);
nand U4718 (N_4718,N_3894,N_2958);
nor U4719 (N_4719,N_2417,N_3755);
nor U4720 (N_4720,N_2926,N_3160);
nor U4721 (N_4721,N_2817,N_2031);
nand U4722 (N_4722,N_2935,N_2904);
and U4723 (N_4723,N_2163,N_3745);
or U4724 (N_4724,N_3311,N_2475);
nand U4725 (N_4725,N_3416,N_3604);
and U4726 (N_4726,N_2119,N_3043);
or U4727 (N_4727,N_2187,N_2751);
and U4728 (N_4728,N_3143,N_3726);
and U4729 (N_4729,N_3476,N_3314);
nand U4730 (N_4730,N_2089,N_2320);
nand U4731 (N_4731,N_3019,N_3496);
nand U4732 (N_4732,N_3263,N_3823);
xor U4733 (N_4733,N_3897,N_3287);
or U4734 (N_4734,N_2247,N_2342);
and U4735 (N_4735,N_2667,N_2998);
nor U4736 (N_4736,N_2057,N_2875);
or U4737 (N_4737,N_3491,N_3021);
and U4738 (N_4738,N_3095,N_3639);
and U4739 (N_4739,N_2465,N_3249);
nor U4740 (N_4740,N_3605,N_3379);
and U4741 (N_4741,N_2812,N_3753);
nor U4742 (N_4742,N_2497,N_2047);
and U4743 (N_4743,N_2485,N_3170);
and U4744 (N_4744,N_3929,N_2003);
nor U4745 (N_4745,N_2393,N_3074);
nand U4746 (N_4746,N_3924,N_3203);
nand U4747 (N_4747,N_2574,N_3088);
nand U4748 (N_4748,N_2192,N_2027);
nor U4749 (N_4749,N_2004,N_2443);
nor U4750 (N_4750,N_3369,N_2506);
nand U4751 (N_4751,N_3595,N_3069);
nor U4752 (N_4752,N_2846,N_2919);
nand U4753 (N_4753,N_2585,N_2592);
and U4754 (N_4754,N_3318,N_2636);
nand U4755 (N_4755,N_3497,N_3010);
nand U4756 (N_4756,N_3414,N_2507);
nor U4757 (N_4757,N_2514,N_2622);
or U4758 (N_4758,N_3784,N_3471);
nand U4759 (N_4759,N_3969,N_2658);
and U4760 (N_4760,N_2789,N_3609);
nand U4761 (N_4761,N_2422,N_2701);
nor U4762 (N_4762,N_2887,N_2525);
and U4763 (N_4763,N_2891,N_3837);
or U4764 (N_4764,N_3697,N_2916);
and U4765 (N_4765,N_2934,N_2635);
nor U4766 (N_4766,N_3918,N_3778);
nand U4767 (N_4767,N_3678,N_2734);
nand U4768 (N_4768,N_3805,N_2326);
nand U4769 (N_4769,N_3265,N_3345);
or U4770 (N_4770,N_3227,N_2611);
nor U4771 (N_4771,N_3902,N_2845);
nand U4772 (N_4772,N_3571,N_2722);
or U4773 (N_4773,N_3508,N_2178);
and U4774 (N_4774,N_3299,N_2881);
and U4775 (N_4775,N_3106,N_2847);
and U4776 (N_4776,N_2282,N_2973);
or U4777 (N_4777,N_2841,N_3884);
and U4778 (N_4778,N_2385,N_3400);
and U4779 (N_4779,N_2160,N_2644);
or U4780 (N_4780,N_2770,N_3868);
or U4781 (N_4781,N_2494,N_3903);
nand U4782 (N_4782,N_3960,N_3564);
or U4783 (N_4783,N_2468,N_2536);
and U4784 (N_4784,N_2500,N_3944);
nor U4785 (N_4785,N_3358,N_3889);
xor U4786 (N_4786,N_2101,N_2193);
and U4787 (N_4787,N_3874,N_3860);
nand U4788 (N_4788,N_3635,N_3245);
and U4789 (N_4789,N_2677,N_3854);
nand U4790 (N_4790,N_2245,N_2829);
and U4791 (N_4791,N_2753,N_2217);
nand U4792 (N_4792,N_3024,N_3729);
nand U4793 (N_4793,N_2684,N_3097);
nand U4794 (N_4794,N_3016,N_3985);
nor U4795 (N_4795,N_3976,N_3825);
nand U4796 (N_4796,N_3811,N_3756);
xor U4797 (N_4797,N_3038,N_3451);
or U4798 (N_4798,N_2575,N_2153);
nand U4799 (N_4799,N_2324,N_3945);
and U4800 (N_4800,N_2436,N_2296);
and U4801 (N_4801,N_3857,N_3535);
nand U4802 (N_4802,N_2276,N_3065);
and U4803 (N_4803,N_2107,N_3744);
nor U4804 (N_4804,N_2328,N_3559);
nor U4805 (N_4805,N_3568,N_2150);
nand U4806 (N_4806,N_3843,N_3023);
nor U4807 (N_4807,N_2054,N_3576);
nor U4808 (N_4808,N_2969,N_3660);
or U4809 (N_4809,N_2579,N_2683);
or U4810 (N_4810,N_3092,N_3841);
nor U4811 (N_4811,N_2360,N_3953);
or U4812 (N_4812,N_2522,N_3735);
nor U4813 (N_4813,N_2698,N_3473);
nand U4814 (N_4814,N_2878,N_3064);
or U4815 (N_4815,N_3544,N_3832);
nand U4816 (N_4816,N_3222,N_2827);
nand U4817 (N_4817,N_2629,N_2657);
and U4818 (N_4818,N_2613,N_3355);
nand U4819 (N_4819,N_2372,N_2643);
nand U4820 (N_4820,N_2208,N_2391);
and U4821 (N_4821,N_2113,N_2642);
and U4822 (N_4822,N_2223,N_3721);
or U4823 (N_4823,N_3962,N_3006);
and U4824 (N_4824,N_2437,N_3590);
nand U4825 (N_4825,N_3569,N_3396);
nand U4826 (N_4826,N_3027,N_3558);
or U4827 (N_4827,N_3607,N_2293);
and U4828 (N_4828,N_3022,N_3818);
nand U4829 (N_4829,N_3552,N_2835);
nor U4830 (N_4830,N_3713,N_3611);
or U4831 (N_4831,N_2641,N_2732);
or U4832 (N_4832,N_2796,N_3403);
nor U4833 (N_4833,N_2190,N_2311);
nand U4834 (N_4834,N_2095,N_3166);
or U4835 (N_4835,N_3972,N_2654);
nand U4836 (N_4836,N_2074,N_2923);
nand U4837 (N_4837,N_2517,N_2854);
or U4838 (N_4838,N_3061,N_2427);
or U4839 (N_4839,N_2664,N_2339);
nand U4840 (N_4840,N_3602,N_3922);
or U4841 (N_4841,N_2986,N_2924);
nor U4842 (N_4842,N_3562,N_2182);
nand U4843 (N_4843,N_3971,N_2462);
or U4844 (N_4844,N_2800,N_3054);
nor U4845 (N_4845,N_3572,N_2950);
nor U4846 (N_4846,N_3056,N_2396);
or U4847 (N_4847,N_2065,N_3898);
nand U4848 (N_4848,N_2598,N_2034);
or U4849 (N_4849,N_2949,N_2377);
and U4850 (N_4850,N_2979,N_2200);
nor U4851 (N_4851,N_2269,N_2419);
nand U4852 (N_4852,N_2856,N_2071);
or U4853 (N_4853,N_2105,N_3765);
and U4854 (N_4854,N_2076,N_2053);
nand U4855 (N_4855,N_3251,N_2761);
nand U4856 (N_4856,N_3584,N_2925);
or U4857 (N_4857,N_2554,N_2412);
and U4858 (N_4858,N_3408,N_3836);
nand U4859 (N_4859,N_3671,N_3478);
or U4860 (N_4860,N_2977,N_3181);
or U4861 (N_4861,N_3464,N_3940);
or U4862 (N_4862,N_2516,N_2871);
nor U4863 (N_4863,N_3330,N_2235);
and U4864 (N_4864,N_2464,N_2992);
nand U4865 (N_4865,N_3931,N_2461);
or U4866 (N_4866,N_2738,N_2362);
and U4867 (N_4867,N_2442,N_3851);
nor U4868 (N_4868,N_3534,N_3586);
and U4869 (N_4869,N_3437,N_2072);
and U4870 (N_4870,N_2978,N_2162);
nand U4871 (N_4871,N_3749,N_3258);
nand U4872 (N_4872,N_2152,N_3429);
nor U4873 (N_4873,N_3883,N_2380);
nor U4874 (N_4874,N_2347,N_3675);
nor U4875 (N_4875,N_3573,N_2204);
and U4876 (N_4876,N_3574,N_2952);
nor U4877 (N_4877,N_3904,N_2403);
or U4878 (N_4878,N_3207,N_2408);
nand U4879 (N_4879,N_3361,N_2861);
nand U4880 (N_4880,N_2255,N_3812);
nand U4881 (N_4881,N_2199,N_2595);
nor U4882 (N_4882,N_2932,N_3498);
nand U4883 (N_4883,N_3882,N_2523);
or U4884 (N_4884,N_2696,N_2563);
and U4885 (N_4885,N_2782,N_2566);
or U4886 (N_4886,N_3991,N_2865);
and U4887 (N_4887,N_3387,N_2205);
nand U4888 (N_4888,N_2438,N_2303);
nor U4889 (N_4889,N_3701,N_3758);
and U4890 (N_4890,N_3738,N_3044);
and U4891 (N_4891,N_2914,N_3567);
or U4892 (N_4892,N_2056,N_2272);
and U4893 (N_4893,N_3344,N_2539);
nor U4894 (N_4894,N_3237,N_2550);
and U4895 (N_4895,N_2147,N_3804);
nor U4896 (N_4896,N_3119,N_2206);
nand U4897 (N_4897,N_2367,N_2710);
or U4898 (N_4898,N_2586,N_3708);
nor U4899 (N_4899,N_2504,N_3339);
or U4900 (N_4900,N_2776,N_3970);
nor U4901 (N_4901,N_2758,N_2717);
or U4902 (N_4902,N_3899,N_3025);
and U4903 (N_4903,N_2456,N_3624);
or U4904 (N_4904,N_3420,N_3186);
nand U4905 (N_4905,N_2277,N_2640);
nand U4906 (N_4906,N_3750,N_2576);
nor U4907 (N_4907,N_3193,N_2432);
or U4908 (N_4908,N_3934,N_3031);
or U4909 (N_4909,N_3276,N_3086);
and U4910 (N_4910,N_3731,N_3849);
nor U4911 (N_4911,N_3101,N_2041);
and U4912 (N_4912,N_3161,N_3456);
nor U4913 (N_4913,N_3565,N_3012);
xor U4914 (N_4914,N_3036,N_2021);
or U4915 (N_4915,N_2818,N_3347);
nor U4916 (N_4916,N_2473,N_2988);
and U4917 (N_4917,N_2748,N_2189);
or U4918 (N_4918,N_2164,N_3593);
and U4919 (N_4919,N_2731,N_3830);
or U4920 (N_4920,N_3667,N_2172);
or U4921 (N_4921,N_2020,N_3048);
and U4922 (N_4922,N_3932,N_3550);
and U4923 (N_4923,N_3630,N_2974);
and U4924 (N_4924,N_2264,N_2668);
nand U4925 (N_4925,N_3563,N_2721);
nand U4926 (N_4926,N_3734,N_3206);
nor U4927 (N_4927,N_2185,N_2167);
nand U4928 (N_4928,N_2166,N_3989);
or U4929 (N_4929,N_2797,N_2862);
nand U4930 (N_4930,N_2337,N_3509);
nand U4931 (N_4931,N_3112,N_3546);
nand U4932 (N_4932,N_2842,N_2416);
or U4933 (N_4933,N_3551,N_2499);
nor U4934 (N_4934,N_2907,N_3082);
and U4935 (N_4935,N_2358,N_3521);
and U4936 (N_4936,N_2055,N_3443);
or U4937 (N_4937,N_3018,N_3557);
nor U4938 (N_4938,N_2735,N_3598);
nand U4939 (N_4939,N_3714,N_2359);
or U4940 (N_4940,N_2070,N_3525);
nand U4941 (N_4941,N_3126,N_3228);
or U4942 (N_4942,N_3308,N_3268);
nand U4943 (N_4943,N_3304,N_3415);
nand U4944 (N_4944,N_2407,N_2614);
or U4945 (N_4945,N_3769,N_3543);
nand U4946 (N_4946,N_2139,N_3655);
nand U4947 (N_4947,N_2219,N_2615);
nand U4948 (N_4948,N_3009,N_2943);
nor U4949 (N_4949,N_3261,N_3839);
and U4950 (N_4950,N_2325,N_3594);
and U4951 (N_4951,N_3561,N_3694);
nand U4952 (N_4952,N_3257,N_2715);
or U4953 (N_4953,N_3277,N_3998);
and U4954 (N_4954,N_2653,N_3370);
and U4955 (N_4955,N_3580,N_3782);
and U4956 (N_4956,N_2864,N_2274);
or U4957 (N_4957,N_3178,N_2639);
nor U4958 (N_4958,N_2967,N_2389);
nand U4959 (N_4959,N_2404,N_3528);
and U4960 (N_4960,N_2631,N_3460);
nor U4961 (N_4961,N_2477,N_2833);
and U4962 (N_4962,N_3405,N_2569);
or U4963 (N_4963,N_3348,N_3444);
nor U4964 (N_4964,N_3467,N_3741);
nor U4965 (N_4965,N_3356,N_3322);
or U4966 (N_4966,N_3616,N_3997);
and U4967 (N_4967,N_3256,N_3377);
and U4968 (N_4968,N_2112,N_3411);
and U4969 (N_4969,N_2356,N_3134);
and U4970 (N_4970,N_2307,N_2508);
nand U4971 (N_4971,N_3077,N_2467);
nand U4972 (N_4972,N_2692,N_3606);
and U4973 (N_4973,N_2369,N_3294);
and U4974 (N_4974,N_2203,N_3946);
nor U4975 (N_4975,N_2013,N_3034);
or U4976 (N_4976,N_2001,N_3455);
and U4977 (N_4977,N_3288,N_3622);
nand U4978 (N_4978,N_2104,N_2038);
nand U4979 (N_4979,N_3644,N_2451);
nand U4980 (N_4980,N_2458,N_2351);
and U4981 (N_4981,N_3853,N_3210);
nand U4982 (N_4982,N_2000,N_2002);
nor U4983 (N_4983,N_2063,N_2048);
nand U4984 (N_4984,N_2909,N_3636);
nand U4985 (N_4985,N_2486,N_3073);
and U4986 (N_4986,N_3425,N_3262);
or U4987 (N_4987,N_3147,N_3833);
nor U4988 (N_4988,N_3259,N_2117);
nand U4989 (N_4989,N_3872,N_2672);
nand U4990 (N_4990,N_3452,N_2240);
or U4991 (N_4991,N_3296,N_3190);
nor U4992 (N_4992,N_2713,N_2617);
or U4993 (N_4993,N_2994,N_2394);
nand U4994 (N_4994,N_2017,N_3930);
or U4995 (N_4995,N_2894,N_2305);
nor U4996 (N_4996,N_3910,N_3364);
and U4997 (N_4997,N_2599,N_3492);
nand U4998 (N_4998,N_2158,N_3692);
and U4999 (N_4999,N_3264,N_2526);
and U5000 (N_5000,N_2124,N_3526);
or U5001 (N_5001,N_3491,N_3798);
nand U5002 (N_5002,N_3103,N_2904);
or U5003 (N_5003,N_2369,N_2143);
or U5004 (N_5004,N_3739,N_2232);
or U5005 (N_5005,N_2671,N_2097);
and U5006 (N_5006,N_3793,N_3911);
nand U5007 (N_5007,N_2004,N_3715);
or U5008 (N_5008,N_3565,N_2917);
and U5009 (N_5009,N_2318,N_3090);
nor U5010 (N_5010,N_3764,N_2479);
and U5011 (N_5011,N_3335,N_2298);
nand U5012 (N_5012,N_2273,N_3051);
or U5013 (N_5013,N_3521,N_3465);
nand U5014 (N_5014,N_3931,N_2535);
and U5015 (N_5015,N_3255,N_3510);
nand U5016 (N_5016,N_2625,N_2944);
nand U5017 (N_5017,N_2043,N_3330);
nor U5018 (N_5018,N_3700,N_3413);
nand U5019 (N_5019,N_2050,N_3577);
or U5020 (N_5020,N_2913,N_3155);
and U5021 (N_5021,N_3812,N_2574);
and U5022 (N_5022,N_3295,N_2665);
nand U5023 (N_5023,N_3631,N_2966);
or U5024 (N_5024,N_3878,N_3499);
or U5025 (N_5025,N_2138,N_3238);
or U5026 (N_5026,N_2792,N_3063);
or U5027 (N_5027,N_3099,N_2780);
or U5028 (N_5028,N_3848,N_2345);
nor U5029 (N_5029,N_2200,N_3998);
nor U5030 (N_5030,N_2185,N_3221);
or U5031 (N_5031,N_3441,N_3675);
or U5032 (N_5032,N_2689,N_3641);
and U5033 (N_5033,N_2426,N_2960);
nor U5034 (N_5034,N_3815,N_3916);
or U5035 (N_5035,N_2122,N_2153);
and U5036 (N_5036,N_2746,N_3899);
xor U5037 (N_5037,N_3754,N_3230);
nand U5038 (N_5038,N_3614,N_3413);
or U5039 (N_5039,N_2829,N_2142);
nand U5040 (N_5040,N_3337,N_3176);
or U5041 (N_5041,N_2095,N_2480);
nand U5042 (N_5042,N_3040,N_2754);
nand U5043 (N_5043,N_2910,N_3045);
nand U5044 (N_5044,N_2287,N_2205);
nor U5045 (N_5045,N_2839,N_2837);
or U5046 (N_5046,N_2481,N_2003);
nand U5047 (N_5047,N_3754,N_2332);
and U5048 (N_5048,N_3336,N_2335);
and U5049 (N_5049,N_2709,N_2007);
and U5050 (N_5050,N_2880,N_2039);
and U5051 (N_5051,N_3768,N_3565);
and U5052 (N_5052,N_3035,N_3950);
nand U5053 (N_5053,N_3911,N_2901);
nand U5054 (N_5054,N_3916,N_2570);
nor U5055 (N_5055,N_2645,N_2043);
or U5056 (N_5056,N_3978,N_3417);
nand U5057 (N_5057,N_3083,N_2621);
nand U5058 (N_5058,N_2299,N_3568);
nand U5059 (N_5059,N_3898,N_2029);
or U5060 (N_5060,N_3878,N_2950);
or U5061 (N_5061,N_3830,N_3272);
nor U5062 (N_5062,N_2949,N_2341);
and U5063 (N_5063,N_2426,N_3257);
nor U5064 (N_5064,N_3401,N_2677);
or U5065 (N_5065,N_2120,N_3575);
nor U5066 (N_5066,N_2144,N_2989);
or U5067 (N_5067,N_2114,N_3213);
nand U5068 (N_5068,N_3454,N_2591);
nor U5069 (N_5069,N_2550,N_3167);
nand U5070 (N_5070,N_3720,N_2219);
nor U5071 (N_5071,N_3478,N_2815);
or U5072 (N_5072,N_3128,N_2039);
or U5073 (N_5073,N_3006,N_3702);
and U5074 (N_5074,N_2933,N_3216);
nor U5075 (N_5075,N_3916,N_2482);
nor U5076 (N_5076,N_3751,N_2084);
or U5077 (N_5077,N_3251,N_2782);
or U5078 (N_5078,N_3072,N_3425);
nor U5079 (N_5079,N_2686,N_2840);
nand U5080 (N_5080,N_3219,N_3509);
and U5081 (N_5081,N_3441,N_3553);
and U5082 (N_5082,N_2791,N_3312);
or U5083 (N_5083,N_3822,N_3633);
and U5084 (N_5084,N_2934,N_2663);
or U5085 (N_5085,N_3233,N_2671);
and U5086 (N_5086,N_2752,N_3397);
or U5087 (N_5087,N_2108,N_3267);
nor U5088 (N_5088,N_2878,N_2024);
and U5089 (N_5089,N_3094,N_3408);
and U5090 (N_5090,N_2470,N_3250);
or U5091 (N_5091,N_2892,N_2194);
nand U5092 (N_5092,N_2627,N_3882);
and U5093 (N_5093,N_2578,N_2698);
nor U5094 (N_5094,N_3440,N_3935);
nor U5095 (N_5095,N_2849,N_2620);
and U5096 (N_5096,N_2520,N_3745);
or U5097 (N_5097,N_2697,N_3571);
nor U5098 (N_5098,N_3100,N_2818);
nand U5099 (N_5099,N_2319,N_3162);
nor U5100 (N_5100,N_3789,N_2474);
nand U5101 (N_5101,N_3981,N_3945);
nand U5102 (N_5102,N_2363,N_3282);
or U5103 (N_5103,N_2273,N_2166);
or U5104 (N_5104,N_3889,N_3642);
or U5105 (N_5105,N_2443,N_3392);
nand U5106 (N_5106,N_2732,N_3268);
and U5107 (N_5107,N_2584,N_2184);
or U5108 (N_5108,N_3114,N_3684);
or U5109 (N_5109,N_2331,N_2171);
nand U5110 (N_5110,N_3517,N_2819);
nor U5111 (N_5111,N_3302,N_3816);
and U5112 (N_5112,N_3233,N_3774);
or U5113 (N_5113,N_3755,N_2357);
or U5114 (N_5114,N_3279,N_2549);
and U5115 (N_5115,N_2688,N_2949);
and U5116 (N_5116,N_3322,N_3323);
nor U5117 (N_5117,N_2988,N_2949);
nor U5118 (N_5118,N_2229,N_3071);
nor U5119 (N_5119,N_3625,N_3782);
nor U5120 (N_5120,N_2846,N_2949);
or U5121 (N_5121,N_3097,N_3797);
or U5122 (N_5122,N_2960,N_2002);
and U5123 (N_5123,N_2687,N_3248);
and U5124 (N_5124,N_2766,N_2908);
nor U5125 (N_5125,N_2947,N_3813);
and U5126 (N_5126,N_2028,N_3237);
or U5127 (N_5127,N_3330,N_3352);
or U5128 (N_5128,N_3298,N_2169);
nand U5129 (N_5129,N_3907,N_2366);
or U5130 (N_5130,N_3868,N_3843);
or U5131 (N_5131,N_3672,N_3137);
nand U5132 (N_5132,N_3174,N_3534);
and U5133 (N_5133,N_3012,N_3234);
nand U5134 (N_5134,N_2910,N_3745);
nor U5135 (N_5135,N_3224,N_2605);
nor U5136 (N_5136,N_2275,N_3611);
nor U5137 (N_5137,N_3064,N_3015);
or U5138 (N_5138,N_3872,N_3442);
nor U5139 (N_5139,N_3258,N_3549);
nor U5140 (N_5140,N_2356,N_3045);
and U5141 (N_5141,N_2383,N_3549);
nand U5142 (N_5142,N_2732,N_2812);
or U5143 (N_5143,N_3007,N_3168);
nand U5144 (N_5144,N_2625,N_3611);
or U5145 (N_5145,N_2906,N_2648);
or U5146 (N_5146,N_3290,N_2505);
nor U5147 (N_5147,N_2843,N_3523);
nor U5148 (N_5148,N_2394,N_2918);
nor U5149 (N_5149,N_2815,N_3934);
nand U5150 (N_5150,N_2704,N_2499);
or U5151 (N_5151,N_3680,N_3307);
nor U5152 (N_5152,N_2983,N_2490);
and U5153 (N_5153,N_2215,N_3311);
nand U5154 (N_5154,N_2152,N_3769);
and U5155 (N_5155,N_3689,N_2058);
nor U5156 (N_5156,N_2513,N_3713);
and U5157 (N_5157,N_3834,N_3736);
nor U5158 (N_5158,N_3941,N_2646);
and U5159 (N_5159,N_2665,N_2973);
nor U5160 (N_5160,N_2609,N_2281);
nand U5161 (N_5161,N_2159,N_2134);
and U5162 (N_5162,N_3915,N_2023);
nand U5163 (N_5163,N_2736,N_3467);
nand U5164 (N_5164,N_3318,N_3330);
nand U5165 (N_5165,N_2033,N_3151);
xor U5166 (N_5166,N_2768,N_3027);
nor U5167 (N_5167,N_3687,N_2050);
nor U5168 (N_5168,N_3110,N_3003);
nand U5169 (N_5169,N_3273,N_2105);
or U5170 (N_5170,N_2066,N_2674);
or U5171 (N_5171,N_3190,N_3186);
or U5172 (N_5172,N_3932,N_2122);
and U5173 (N_5173,N_3068,N_2489);
or U5174 (N_5174,N_2791,N_2173);
and U5175 (N_5175,N_2182,N_2759);
nand U5176 (N_5176,N_3705,N_3786);
or U5177 (N_5177,N_2137,N_2468);
and U5178 (N_5178,N_3620,N_2808);
nand U5179 (N_5179,N_2323,N_2645);
and U5180 (N_5180,N_3637,N_2629);
and U5181 (N_5181,N_2170,N_2098);
or U5182 (N_5182,N_2842,N_3874);
nand U5183 (N_5183,N_2508,N_2120);
and U5184 (N_5184,N_2048,N_3900);
nand U5185 (N_5185,N_3797,N_2864);
nand U5186 (N_5186,N_2596,N_3786);
nor U5187 (N_5187,N_2402,N_3832);
xor U5188 (N_5188,N_2514,N_3118);
nand U5189 (N_5189,N_3114,N_2436);
or U5190 (N_5190,N_3553,N_2792);
xnor U5191 (N_5191,N_2154,N_3293);
nand U5192 (N_5192,N_3590,N_3559);
and U5193 (N_5193,N_2311,N_3196);
or U5194 (N_5194,N_3755,N_3685);
or U5195 (N_5195,N_3055,N_2641);
and U5196 (N_5196,N_3257,N_3216);
nand U5197 (N_5197,N_2056,N_3802);
nand U5198 (N_5198,N_2970,N_3872);
or U5199 (N_5199,N_2693,N_3766);
xor U5200 (N_5200,N_3158,N_2069);
or U5201 (N_5201,N_2603,N_2311);
or U5202 (N_5202,N_2007,N_2724);
and U5203 (N_5203,N_2465,N_2641);
and U5204 (N_5204,N_3429,N_3501);
nor U5205 (N_5205,N_3784,N_3386);
or U5206 (N_5206,N_3808,N_3856);
nor U5207 (N_5207,N_2992,N_3802);
or U5208 (N_5208,N_3034,N_3629);
nand U5209 (N_5209,N_3217,N_3927);
and U5210 (N_5210,N_3921,N_2608);
or U5211 (N_5211,N_2257,N_2821);
and U5212 (N_5212,N_2467,N_2698);
and U5213 (N_5213,N_2807,N_3329);
and U5214 (N_5214,N_3323,N_2317);
nor U5215 (N_5215,N_3643,N_2107);
nand U5216 (N_5216,N_3021,N_2746);
nand U5217 (N_5217,N_3458,N_2732);
nor U5218 (N_5218,N_3963,N_2936);
or U5219 (N_5219,N_2009,N_3966);
and U5220 (N_5220,N_2065,N_2789);
or U5221 (N_5221,N_2319,N_3196);
nor U5222 (N_5222,N_3545,N_3807);
or U5223 (N_5223,N_2923,N_3771);
nor U5224 (N_5224,N_3190,N_2814);
nand U5225 (N_5225,N_2261,N_3539);
nor U5226 (N_5226,N_3925,N_2939);
nor U5227 (N_5227,N_3568,N_3386);
nor U5228 (N_5228,N_3387,N_3471);
nand U5229 (N_5229,N_3864,N_2473);
nand U5230 (N_5230,N_2865,N_2027);
or U5231 (N_5231,N_3345,N_2118);
nor U5232 (N_5232,N_3771,N_2601);
nand U5233 (N_5233,N_3292,N_3000);
nand U5234 (N_5234,N_3602,N_2925);
nor U5235 (N_5235,N_2748,N_3307);
nand U5236 (N_5236,N_3032,N_2077);
and U5237 (N_5237,N_3082,N_3317);
nor U5238 (N_5238,N_3134,N_3121);
nor U5239 (N_5239,N_2784,N_3949);
or U5240 (N_5240,N_2480,N_3521);
nor U5241 (N_5241,N_3166,N_3011);
nand U5242 (N_5242,N_2056,N_3640);
nor U5243 (N_5243,N_3509,N_2682);
or U5244 (N_5244,N_3083,N_2058);
and U5245 (N_5245,N_3920,N_2541);
or U5246 (N_5246,N_2335,N_2122);
nand U5247 (N_5247,N_3653,N_3745);
or U5248 (N_5248,N_2979,N_2377);
nand U5249 (N_5249,N_2821,N_2044);
and U5250 (N_5250,N_3003,N_2959);
and U5251 (N_5251,N_3715,N_2759);
nand U5252 (N_5252,N_2944,N_2844);
or U5253 (N_5253,N_2258,N_3734);
nand U5254 (N_5254,N_2990,N_3684);
nor U5255 (N_5255,N_2298,N_2867);
nand U5256 (N_5256,N_3020,N_2555);
or U5257 (N_5257,N_2223,N_2264);
or U5258 (N_5258,N_2004,N_3667);
nor U5259 (N_5259,N_3434,N_2909);
nor U5260 (N_5260,N_2524,N_3151);
or U5261 (N_5261,N_2971,N_3406);
or U5262 (N_5262,N_3143,N_2438);
or U5263 (N_5263,N_3499,N_3768);
nand U5264 (N_5264,N_2323,N_3717);
and U5265 (N_5265,N_3029,N_2248);
or U5266 (N_5266,N_3262,N_3819);
nand U5267 (N_5267,N_3004,N_2736);
and U5268 (N_5268,N_3500,N_3607);
nand U5269 (N_5269,N_2451,N_2187);
nor U5270 (N_5270,N_2771,N_3431);
nor U5271 (N_5271,N_2983,N_3704);
or U5272 (N_5272,N_2982,N_2362);
and U5273 (N_5273,N_3677,N_2035);
nor U5274 (N_5274,N_3694,N_3153);
or U5275 (N_5275,N_3978,N_2649);
and U5276 (N_5276,N_2955,N_2056);
or U5277 (N_5277,N_2964,N_3562);
nor U5278 (N_5278,N_3051,N_2469);
nand U5279 (N_5279,N_3692,N_3326);
nand U5280 (N_5280,N_2103,N_2222);
nor U5281 (N_5281,N_3478,N_2173);
nand U5282 (N_5282,N_2471,N_3633);
or U5283 (N_5283,N_3172,N_3450);
or U5284 (N_5284,N_3909,N_3484);
nor U5285 (N_5285,N_2536,N_2810);
nand U5286 (N_5286,N_2300,N_3361);
nor U5287 (N_5287,N_2937,N_2200);
nor U5288 (N_5288,N_3924,N_2190);
and U5289 (N_5289,N_3198,N_2111);
and U5290 (N_5290,N_3639,N_2803);
nand U5291 (N_5291,N_3463,N_3317);
nor U5292 (N_5292,N_3721,N_3806);
nor U5293 (N_5293,N_3587,N_3696);
nor U5294 (N_5294,N_2795,N_2061);
or U5295 (N_5295,N_3962,N_2562);
and U5296 (N_5296,N_2619,N_2251);
and U5297 (N_5297,N_3162,N_2981);
nor U5298 (N_5298,N_2173,N_2542);
nor U5299 (N_5299,N_2663,N_2560);
and U5300 (N_5300,N_2638,N_3733);
or U5301 (N_5301,N_3029,N_2527);
or U5302 (N_5302,N_2226,N_3909);
and U5303 (N_5303,N_3268,N_3203);
and U5304 (N_5304,N_3665,N_3301);
nand U5305 (N_5305,N_3045,N_2105);
nand U5306 (N_5306,N_2721,N_3265);
nand U5307 (N_5307,N_3144,N_3129);
or U5308 (N_5308,N_3030,N_2027);
and U5309 (N_5309,N_3762,N_2776);
nor U5310 (N_5310,N_2384,N_3719);
or U5311 (N_5311,N_3831,N_2886);
and U5312 (N_5312,N_2056,N_2667);
nor U5313 (N_5313,N_2832,N_2249);
nand U5314 (N_5314,N_3566,N_2135);
nand U5315 (N_5315,N_3723,N_3435);
nor U5316 (N_5316,N_3919,N_2051);
nand U5317 (N_5317,N_2338,N_2522);
or U5318 (N_5318,N_2758,N_2865);
or U5319 (N_5319,N_2068,N_2760);
and U5320 (N_5320,N_2823,N_2502);
and U5321 (N_5321,N_2898,N_3685);
nor U5322 (N_5322,N_2445,N_2138);
and U5323 (N_5323,N_3265,N_3349);
or U5324 (N_5324,N_2958,N_2766);
nor U5325 (N_5325,N_3553,N_2400);
or U5326 (N_5326,N_2383,N_2992);
nand U5327 (N_5327,N_2161,N_2302);
and U5328 (N_5328,N_2962,N_3317);
and U5329 (N_5329,N_3068,N_3880);
nor U5330 (N_5330,N_3551,N_3539);
or U5331 (N_5331,N_3614,N_2036);
nand U5332 (N_5332,N_2328,N_2303);
or U5333 (N_5333,N_3976,N_3814);
and U5334 (N_5334,N_2801,N_3092);
or U5335 (N_5335,N_2125,N_2182);
and U5336 (N_5336,N_2873,N_2650);
or U5337 (N_5337,N_2292,N_2227);
or U5338 (N_5338,N_2015,N_2109);
nand U5339 (N_5339,N_2070,N_3382);
and U5340 (N_5340,N_3818,N_2724);
nor U5341 (N_5341,N_3150,N_2151);
and U5342 (N_5342,N_3066,N_2728);
and U5343 (N_5343,N_2279,N_3420);
and U5344 (N_5344,N_2283,N_2141);
and U5345 (N_5345,N_2066,N_2296);
nor U5346 (N_5346,N_3389,N_3648);
or U5347 (N_5347,N_3983,N_2133);
nand U5348 (N_5348,N_2083,N_3239);
nor U5349 (N_5349,N_2730,N_3699);
nand U5350 (N_5350,N_2570,N_2941);
nand U5351 (N_5351,N_2739,N_2847);
and U5352 (N_5352,N_2806,N_3751);
nand U5353 (N_5353,N_2744,N_3856);
or U5354 (N_5354,N_2247,N_3246);
or U5355 (N_5355,N_3106,N_2125);
nor U5356 (N_5356,N_2044,N_2390);
and U5357 (N_5357,N_2349,N_3257);
and U5358 (N_5358,N_3023,N_2592);
and U5359 (N_5359,N_3078,N_2959);
nand U5360 (N_5360,N_2854,N_2425);
nor U5361 (N_5361,N_3575,N_3817);
nand U5362 (N_5362,N_3919,N_3418);
and U5363 (N_5363,N_3781,N_3683);
and U5364 (N_5364,N_3765,N_2350);
nand U5365 (N_5365,N_2677,N_3781);
and U5366 (N_5366,N_3160,N_2256);
nor U5367 (N_5367,N_3778,N_2492);
nor U5368 (N_5368,N_2635,N_2340);
or U5369 (N_5369,N_3041,N_2054);
or U5370 (N_5370,N_3434,N_3696);
nand U5371 (N_5371,N_2967,N_2975);
nor U5372 (N_5372,N_2197,N_3069);
or U5373 (N_5373,N_2252,N_3553);
nand U5374 (N_5374,N_2456,N_2476);
nand U5375 (N_5375,N_2160,N_3856);
nand U5376 (N_5376,N_2526,N_3684);
nor U5377 (N_5377,N_3280,N_3976);
and U5378 (N_5378,N_3896,N_2668);
or U5379 (N_5379,N_3344,N_3794);
nor U5380 (N_5380,N_3277,N_2377);
and U5381 (N_5381,N_3770,N_3552);
nor U5382 (N_5382,N_3527,N_3164);
and U5383 (N_5383,N_3174,N_2548);
nand U5384 (N_5384,N_3476,N_2164);
and U5385 (N_5385,N_3092,N_3288);
or U5386 (N_5386,N_3377,N_2956);
and U5387 (N_5387,N_3370,N_2636);
and U5388 (N_5388,N_3567,N_2645);
nor U5389 (N_5389,N_3880,N_3912);
or U5390 (N_5390,N_2560,N_3816);
or U5391 (N_5391,N_3367,N_3569);
nand U5392 (N_5392,N_2350,N_2067);
nand U5393 (N_5393,N_2805,N_2282);
or U5394 (N_5394,N_3111,N_2692);
and U5395 (N_5395,N_2123,N_2364);
and U5396 (N_5396,N_3907,N_2490);
nand U5397 (N_5397,N_3255,N_2862);
nor U5398 (N_5398,N_3279,N_3193);
nand U5399 (N_5399,N_2917,N_2501);
nand U5400 (N_5400,N_2711,N_2516);
nand U5401 (N_5401,N_2173,N_2113);
nor U5402 (N_5402,N_2147,N_3969);
or U5403 (N_5403,N_2569,N_3539);
or U5404 (N_5404,N_2323,N_2654);
or U5405 (N_5405,N_3795,N_3573);
or U5406 (N_5406,N_3055,N_2378);
nor U5407 (N_5407,N_2174,N_2088);
nor U5408 (N_5408,N_3877,N_2801);
nand U5409 (N_5409,N_3936,N_2339);
nand U5410 (N_5410,N_2979,N_2291);
nor U5411 (N_5411,N_2663,N_2717);
nor U5412 (N_5412,N_3111,N_3239);
or U5413 (N_5413,N_2545,N_2013);
nor U5414 (N_5414,N_2484,N_3480);
and U5415 (N_5415,N_3165,N_2027);
nand U5416 (N_5416,N_2213,N_3100);
and U5417 (N_5417,N_3272,N_2823);
nor U5418 (N_5418,N_3736,N_2832);
and U5419 (N_5419,N_3194,N_2213);
nor U5420 (N_5420,N_2548,N_2710);
nand U5421 (N_5421,N_2225,N_3706);
or U5422 (N_5422,N_2846,N_3497);
nor U5423 (N_5423,N_2823,N_3599);
nand U5424 (N_5424,N_2988,N_3841);
or U5425 (N_5425,N_3364,N_3365);
nand U5426 (N_5426,N_3945,N_3772);
nand U5427 (N_5427,N_2895,N_2875);
nand U5428 (N_5428,N_2996,N_2530);
nor U5429 (N_5429,N_3457,N_2513);
nand U5430 (N_5430,N_3985,N_2125);
nand U5431 (N_5431,N_3109,N_3408);
or U5432 (N_5432,N_3084,N_2461);
or U5433 (N_5433,N_3711,N_3100);
nand U5434 (N_5434,N_2838,N_3918);
nand U5435 (N_5435,N_3791,N_3284);
nand U5436 (N_5436,N_3290,N_3813);
or U5437 (N_5437,N_3283,N_3672);
nand U5438 (N_5438,N_2249,N_2236);
nand U5439 (N_5439,N_3887,N_2826);
nor U5440 (N_5440,N_2999,N_2997);
or U5441 (N_5441,N_3418,N_3578);
or U5442 (N_5442,N_3012,N_2279);
nor U5443 (N_5443,N_3586,N_3137);
nand U5444 (N_5444,N_2128,N_2670);
xnor U5445 (N_5445,N_2600,N_3462);
or U5446 (N_5446,N_2223,N_3414);
nand U5447 (N_5447,N_3191,N_2950);
and U5448 (N_5448,N_2932,N_2962);
or U5449 (N_5449,N_2720,N_3510);
and U5450 (N_5450,N_3708,N_3152);
nand U5451 (N_5451,N_2205,N_2371);
and U5452 (N_5452,N_3918,N_3813);
and U5453 (N_5453,N_2276,N_2877);
nand U5454 (N_5454,N_2958,N_2780);
nor U5455 (N_5455,N_2591,N_3865);
nor U5456 (N_5456,N_2982,N_3391);
nor U5457 (N_5457,N_2933,N_3138);
or U5458 (N_5458,N_2701,N_3230);
nand U5459 (N_5459,N_3350,N_2712);
or U5460 (N_5460,N_2659,N_2447);
nand U5461 (N_5461,N_3730,N_3461);
nand U5462 (N_5462,N_2360,N_2882);
or U5463 (N_5463,N_2595,N_2405);
and U5464 (N_5464,N_2119,N_2281);
and U5465 (N_5465,N_2044,N_2312);
nand U5466 (N_5466,N_2654,N_3072);
nand U5467 (N_5467,N_3876,N_3043);
nor U5468 (N_5468,N_2241,N_2111);
nor U5469 (N_5469,N_3834,N_3222);
and U5470 (N_5470,N_2787,N_3639);
or U5471 (N_5471,N_2314,N_2204);
or U5472 (N_5472,N_3573,N_3812);
or U5473 (N_5473,N_3078,N_2900);
and U5474 (N_5474,N_2685,N_3394);
nand U5475 (N_5475,N_2066,N_2374);
nor U5476 (N_5476,N_2281,N_3217);
or U5477 (N_5477,N_3762,N_2152);
or U5478 (N_5478,N_3725,N_2602);
nand U5479 (N_5479,N_2514,N_3688);
nor U5480 (N_5480,N_2273,N_2203);
nor U5481 (N_5481,N_3219,N_2738);
or U5482 (N_5482,N_3161,N_3454);
or U5483 (N_5483,N_3079,N_3892);
and U5484 (N_5484,N_2430,N_2408);
or U5485 (N_5485,N_2161,N_2017);
nor U5486 (N_5486,N_3511,N_2447);
nor U5487 (N_5487,N_2518,N_2279);
and U5488 (N_5488,N_3933,N_3543);
nor U5489 (N_5489,N_3849,N_3762);
and U5490 (N_5490,N_2528,N_2272);
nor U5491 (N_5491,N_3506,N_2283);
or U5492 (N_5492,N_2451,N_2462);
nand U5493 (N_5493,N_3138,N_3861);
or U5494 (N_5494,N_3102,N_2826);
nand U5495 (N_5495,N_2928,N_2500);
or U5496 (N_5496,N_2383,N_3673);
and U5497 (N_5497,N_3201,N_3727);
nand U5498 (N_5498,N_3783,N_3282);
nor U5499 (N_5499,N_2271,N_3715);
nand U5500 (N_5500,N_3141,N_3995);
nand U5501 (N_5501,N_3260,N_3503);
nor U5502 (N_5502,N_3790,N_3551);
and U5503 (N_5503,N_2422,N_3279);
and U5504 (N_5504,N_2849,N_3794);
and U5505 (N_5505,N_3467,N_2554);
or U5506 (N_5506,N_2341,N_3847);
nor U5507 (N_5507,N_2829,N_2857);
nand U5508 (N_5508,N_3143,N_3401);
or U5509 (N_5509,N_2335,N_2597);
and U5510 (N_5510,N_3604,N_2991);
or U5511 (N_5511,N_3295,N_3929);
nand U5512 (N_5512,N_3128,N_2287);
or U5513 (N_5513,N_2002,N_3745);
and U5514 (N_5514,N_2388,N_3317);
and U5515 (N_5515,N_2745,N_2699);
or U5516 (N_5516,N_2637,N_3713);
nor U5517 (N_5517,N_2920,N_2005);
or U5518 (N_5518,N_2524,N_3624);
and U5519 (N_5519,N_2610,N_3517);
nor U5520 (N_5520,N_3893,N_2107);
nor U5521 (N_5521,N_2401,N_2418);
or U5522 (N_5522,N_3627,N_2110);
and U5523 (N_5523,N_3879,N_3982);
nor U5524 (N_5524,N_3136,N_3277);
nand U5525 (N_5525,N_3105,N_2069);
or U5526 (N_5526,N_3957,N_3169);
xor U5527 (N_5527,N_3362,N_3282);
or U5528 (N_5528,N_3770,N_2211);
and U5529 (N_5529,N_2953,N_3182);
nor U5530 (N_5530,N_2505,N_2460);
nand U5531 (N_5531,N_2557,N_3846);
and U5532 (N_5532,N_2565,N_2271);
and U5533 (N_5533,N_3365,N_2628);
nand U5534 (N_5534,N_2619,N_3392);
nor U5535 (N_5535,N_2458,N_2679);
and U5536 (N_5536,N_3125,N_2745);
and U5537 (N_5537,N_2876,N_3113);
nand U5538 (N_5538,N_3071,N_3582);
and U5539 (N_5539,N_2009,N_3147);
nor U5540 (N_5540,N_2411,N_3413);
or U5541 (N_5541,N_2204,N_2277);
nor U5542 (N_5542,N_2710,N_2389);
and U5543 (N_5543,N_2569,N_2637);
and U5544 (N_5544,N_2081,N_2995);
nand U5545 (N_5545,N_3742,N_2209);
and U5546 (N_5546,N_3175,N_3703);
nand U5547 (N_5547,N_3637,N_3104);
or U5548 (N_5548,N_3997,N_2531);
and U5549 (N_5549,N_2872,N_2462);
and U5550 (N_5550,N_3590,N_3631);
nand U5551 (N_5551,N_2624,N_3077);
nor U5552 (N_5552,N_3048,N_3051);
nor U5553 (N_5553,N_2570,N_2850);
nor U5554 (N_5554,N_2148,N_2537);
and U5555 (N_5555,N_3069,N_3957);
nand U5556 (N_5556,N_3903,N_3758);
and U5557 (N_5557,N_3220,N_2743);
xor U5558 (N_5558,N_3191,N_2721);
nor U5559 (N_5559,N_2172,N_2738);
nor U5560 (N_5560,N_3469,N_2452);
or U5561 (N_5561,N_2256,N_2760);
and U5562 (N_5562,N_2544,N_3672);
or U5563 (N_5563,N_3825,N_3317);
or U5564 (N_5564,N_3606,N_2806);
and U5565 (N_5565,N_3794,N_2585);
nand U5566 (N_5566,N_3762,N_2409);
nor U5567 (N_5567,N_3170,N_2746);
or U5568 (N_5568,N_3138,N_2094);
nand U5569 (N_5569,N_3498,N_2442);
nand U5570 (N_5570,N_3100,N_3080);
or U5571 (N_5571,N_2580,N_3903);
nor U5572 (N_5572,N_2320,N_3802);
or U5573 (N_5573,N_2099,N_2904);
and U5574 (N_5574,N_3250,N_3004);
nand U5575 (N_5575,N_3698,N_3938);
or U5576 (N_5576,N_2561,N_2034);
nand U5577 (N_5577,N_3389,N_2806);
or U5578 (N_5578,N_2663,N_2825);
nor U5579 (N_5579,N_2532,N_3253);
or U5580 (N_5580,N_3807,N_2121);
nand U5581 (N_5581,N_2568,N_3668);
nand U5582 (N_5582,N_2848,N_3561);
nand U5583 (N_5583,N_2745,N_2413);
or U5584 (N_5584,N_2611,N_3149);
xnor U5585 (N_5585,N_2701,N_2776);
or U5586 (N_5586,N_3827,N_2370);
nand U5587 (N_5587,N_2096,N_3368);
and U5588 (N_5588,N_2209,N_2371);
or U5589 (N_5589,N_2472,N_2729);
nor U5590 (N_5590,N_2825,N_2874);
nor U5591 (N_5591,N_2899,N_2167);
or U5592 (N_5592,N_3263,N_2943);
or U5593 (N_5593,N_3047,N_3369);
nand U5594 (N_5594,N_2332,N_2927);
nor U5595 (N_5595,N_3553,N_3955);
xor U5596 (N_5596,N_3897,N_2956);
or U5597 (N_5597,N_2776,N_3619);
nor U5598 (N_5598,N_3989,N_2193);
or U5599 (N_5599,N_3499,N_2189);
or U5600 (N_5600,N_3940,N_3397);
or U5601 (N_5601,N_3088,N_3916);
or U5602 (N_5602,N_2713,N_3630);
and U5603 (N_5603,N_2969,N_3729);
nand U5604 (N_5604,N_3724,N_2869);
xor U5605 (N_5605,N_3127,N_2943);
or U5606 (N_5606,N_3716,N_3921);
nor U5607 (N_5607,N_2415,N_3863);
nand U5608 (N_5608,N_3557,N_2434);
and U5609 (N_5609,N_2845,N_2554);
nand U5610 (N_5610,N_3515,N_2457);
nor U5611 (N_5611,N_3397,N_3197);
and U5612 (N_5612,N_2031,N_3220);
nand U5613 (N_5613,N_2702,N_2720);
nor U5614 (N_5614,N_2907,N_2954);
and U5615 (N_5615,N_2984,N_3947);
nand U5616 (N_5616,N_3682,N_2988);
or U5617 (N_5617,N_3332,N_2264);
nand U5618 (N_5618,N_3847,N_3912);
nand U5619 (N_5619,N_3830,N_2341);
and U5620 (N_5620,N_3537,N_2315);
and U5621 (N_5621,N_2034,N_3667);
or U5622 (N_5622,N_3888,N_3964);
or U5623 (N_5623,N_2145,N_2433);
nand U5624 (N_5624,N_2021,N_2635);
or U5625 (N_5625,N_2689,N_2323);
and U5626 (N_5626,N_3608,N_2283);
and U5627 (N_5627,N_2295,N_2625);
nor U5628 (N_5628,N_2515,N_3904);
or U5629 (N_5629,N_2482,N_2347);
nand U5630 (N_5630,N_2665,N_2869);
and U5631 (N_5631,N_3049,N_2896);
nand U5632 (N_5632,N_3591,N_2396);
and U5633 (N_5633,N_3555,N_2207);
or U5634 (N_5634,N_2255,N_3939);
nand U5635 (N_5635,N_2760,N_3792);
nand U5636 (N_5636,N_2319,N_2682);
nor U5637 (N_5637,N_2940,N_2713);
nand U5638 (N_5638,N_3668,N_2028);
or U5639 (N_5639,N_3220,N_2963);
nand U5640 (N_5640,N_2028,N_2063);
nor U5641 (N_5641,N_3109,N_3908);
nor U5642 (N_5642,N_2588,N_3547);
or U5643 (N_5643,N_3817,N_3465);
nand U5644 (N_5644,N_2495,N_3538);
nand U5645 (N_5645,N_3582,N_2286);
nand U5646 (N_5646,N_2611,N_2990);
and U5647 (N_5647,N_3376,N_3731);
nand U5648 (N_5648,N_2214,N_2843);
nor U5649 (N_5649,N_3091,N_3561);
or U5650 (N_5650,N_3802,N_3725);
or U5651 (N_5651,N_3761,N_2248);
nand U5652 (N_5652,N_3860,N_2314);
nor U5653 (N_5653,N_3222,N_2288);
nor U5654 (N_5654,N_3654,N_2506);
nand U5655 (N_5655,N_3141,N_2169);
or U5656 (N_5656,N_2442,N_3408);
nand U5657 (N_5657,N_2771,N_3679);
and U5658 (N_5658,N_3084,N_2078);
and U5659 (N_5659,N_3163,N_2422);
nand U5660 (N_5660,N_3881,N_2108);
or U5661 (N_5661,N_2211,N_3467);
nand U5662 (N_5662,N_2831,N_3692);
nand U5663 (N_5663,N_3252,N_3551);
nand U5664 (N_5664,N_3477,N_2430);
and U5665 (N_5665,N_3370,N_3523);
or U5666 (N_5666,N_2606,N_3508);
and U5667 (N_5667,N_3433,N_2257);
and U5668 (N_5668,N_2946,N_2826);
or U5669 (N_5669,N_3268,N_2150);
and U5670 (N_5670,N_2151,N_3555);
nand U5671 (N_5671,N_2358,N_2381);
nand U5672 (N_5672,N_3110,N_3291);
nor U5673 (N_5673,N_3400,N_3597);
and U5674 (N_5674,N_2618,N_3880);
nor U5675 (N_5675,N_3136,N_3502);
and U5676 (N_5676,N_2327,N_2934);
nor U5677 (N_5677,N_3018,N_2049);
or U5678 (N_5678,N_3422,N_2541);
nand U5679 (N_5679,N_3653,N_3096);
nor U5680 (N_5680,N_3452,N_2366);
and U5681 (N_5681,N_3937,N_2513);
or U5682 (N_5682,N_2260,N_2821);
or U5683 (N_5683,N_2672,N_2978);
nand U5684 (N_5684,N_3955,N_2489);
and U5685 (N_5685,N_3245,N_2834);
nor U5686 (N_5686,N_3320,N_2289);
nor U5687 (N_5687,N_2485,N_3032);
or U5688 (N_5688,N_3795,N_2337);
or U5689 (N_5689,N_2892,N_3091);
nand U5690 (N_5690,N_2502,N_3875);
nand U5691 (N_5691,N_3501,N_2590);
nor U5692 (N_5692,N_2336,N_3746);
or U5693 (N_5693,N_3329,N_2738);
or U5694 (N_5694,N_3285,N_2591);
and U5695 (N_5695,N_2405,N_2188);
and U5696 (N_5696,N_2799,N_3279);
or U5697 (N_5697,N_3997,N_3243);
nor U5698 (N_5698,N_2845,N_2959);
nand U5699 (N_5699,N_2217,N_3995);
and U5700 (N_5700,N_3164,N_3358);
nor U5701 (N_5701,N_2506,N_3865);
nand U5702 (N_5702,N_2696,N_2608);
xnor U5703 (N_5703,N_2879,N_2742);
and U5704 (N_5704,N_3107,N_3433);
and U5705 (N_5705,N_2545,N_2184);
nor U5706 (N_5706,N_3062,N_2021);
or U5707 (N_5707,N_2239,N_3568);
or U5708 (N_5708,N_2365,N_3549);
nand U5709 (N_5709,N_2666,N_2076);
or U5710 (N_5710,N_3598,N_2276);
nand U5711 (N_5711,N_3576,N_3439);
nand U5712 (N_5712,N_3988,N_3414);
nor U5713 (N_5713,N_2454,N_3511);
and U5714 (N_5714,N_2324,N_2866);
or U5715 (N_5715,N_3553,N_3033);
nand U5716 (N_5716,N_3316,N_3967);
and U5717 (N_5717,N_3713,N_2430);
nand U5718 (N_5718,N_3988,N_3269);
or U5719 (N_5719,N_2241,N_2717);
nand U5720 (N_5720,N_2459,N_3375);
or U5721 (N_5721,N_3839,N_2365);
and U5722 (N_5722,N_2918,N_2978);
nand U5723 (N_5723,N_3971,N_3056);
and U5724 (N_5724,N_2093,N_2168);
nand U5725 (N_5725,N_2407,N_3248);
or U5726 (N_5726,N_2522,N_3864);
or U5727 (N_5727,N_3740,N_2759);
nor U5728 (N_5728,N_3398,N_2428);
and U5729 (N_5729,N_3861,N_2574);
or U5730 (N_5730,N_2216,N_3776);
nand U5731 (N_5731,N_3377,N_3152);
nand U5732 (N_5732,N_3233,N_3296);
nand U5733 (N_5733,N_2689,N_2555);
and U5734 (N_5734,N_2619,N_3692);
or U5735 (N_5735,N_2122,N_2145);
nand U5736 (N_5736,N_2448,N_3709);
or U5737 (N_5737,N_3949,N_3724);
nand U5738 (N_5738,N_3314,N_3022);
nand U5739 (N_5739,N_2163,N_2241);
or U5740 (N_5740,N_2546,N_2007);
and U5741 (N_5741,N_2385,N_3189);
and U5742 (N_5742,N_3995,N_3198);
nand U5743 (N_5743,N_3942,N_3870);
or U5744 (N_5744,N_2924,N_2367);
nand U5745 (N_5745,N_3417,N_2357);
nor U5746 (N_5746,N_3792,N_3737);
nand U5747 (N_5747,N_2526,N_2882);
nand U5748 (N_5748,N_3449,N_2999);
nand U5749 (N_5749,N_3433,N_2157);
or U5750 (N_5750,N_3632,N_3757);
nor U5751 (N_5751,N_2611,N_2005);
or U5752 (N_5752,N_2466,N_3408);
or U5753 (N_5753,N_3938,N_3849);
nor U5754 (N_5754,N_3590,N_2933);
or U5755 (N_5755,N_3272,N_2466);
or U5756 (N_5756,N_2501,N_2511);
or U5757 (N_5757,N_2756,N_2185);
nand U5758 (N_5758,N_2651,N_3674);
nand U5759 (N_5759,N_2746,N_2188);
or U5760 (N_5760,N_3437,N_3121);
and U5761 (N_5761,N_2914,N_2437);
and U5762 (N_5762,N_2791,N_2366);
nor U5763 (N_5763,N_2711,N_3826);
nand U5764 (N_5764,N_3899,N_2842);
or U5765 (N_5765,N_2582,N_3091);
and U5766 (N_5766,N_3623,N_2252);
and U5767 (N_5767,N_2794,N_3498);
nand U5768 (N_5768,N_2971,N_2335);
or U5769 (N_5769,N_3066,N_3259);
and U5770 (N_5770,N_3363,N_2886);
or U5771 (N_5771,N_2312,N_2414);
nor U5772 (N_5772,N_3252,N_3959);
nand U5773 (N_5773,N_2196,N_2838);
nand U5774 (N_5774,N_2381,N_3673);
or U5775 (N_5775,N_3134,N_2084);
and U5776 (N_5776,N_3451,N_2412);
and U5777 (N_5777,N_3506,N_2822);
nand U5778 (N_5778,N_3264,N_3747);
and U5779 (N_5779,N_3745,N_2335);
nor U5780 (N_5780,N_2063,N_2520);
and U5781 (N_5781,N_3856,N_2942);
nand U5782 (N_5782,N_2389,N_2067);
or U5783 (N_5783,N_2313,N_3076);
or U5784 (N_5784,N_2136,N_3328);
nor U5785 (N_5785,N_3781,N_2471);
and U5786 (N_5786,N_2417,N_3970);
nand U5787 (N_5787,N_2820,N_3476);
and U5788 (N_5788,N_2629,N_2485);
or U5789 (N_5789,N_2818,N_3056);
nor U5790 (N_5790,N_2477,N_2570);
and U5791 (N_5791,N_2770,N_3243);
or U5792 (N_5792,N_2001,N_2302);
nor U5793 (N_5793,N_3058,N_2275);
nand U5794 (N_5794,N_3046,N_2852);
and U5795 (N_5795,N_3385,N_3090);
nand U5796 (N_5796,N_2806,N_2743);
and U5797 (N_5797,N_2797,N_2147);
or U5798 (N_5798,N_2715,N_2999);
nand U5799 (N_5799,N_2592,N_3564);
nor U5800 (N_5800,N_2852,N_3303);
nor U5801 (N_5801,N_3798,N_3796);
nand U5802 (N_5802,N_2380,N_3332);
and U5803 (N_5803,N_2030,N_3906);
and U5804 (N_5804,N_2265,N_2717);
nor U5805 (N_5805,N_3798,N_3763);
or U5806 (N_5806,N_2806,N_2412);
nand U5807 (N_5807,N_2491,N_2019);
nand U5808 (N_5808,N_2287,N_3890);
and U5809 (N_5809,N_3347,N_3223);
nor U5810 (N_5810,N_2549,N_2953);
or U5811 (N_5811,N_3616,N_3779);
nand U5812 (N_5812,N_2990,N_3787);
nand U5813 (N_5813,N_2452,N_3555);
nor U5814 (N_5814,N_2864,N_3691);
nor U5815 (N_5815,N_2818,N_2492);
nor U5816 (N_5816,N_3120,N_2044);
nor U5817 (N_5817,N_2408,N_2759);
nand U5818 (N_5818,N_2999,N_2871);
nand U5819 (N_5819,N_2117,N_3363);
nor U5820 (N_5820,N_3399,N_3997);
nand U5821 (N_5821,N_3754,N_3418);
nor U5822 (N_5822,N_2197,N_2615);
nor U5823 (N_5823,N_2872,N_3096);
and U5824 (N_5824,N_3703,N_2099);
nand U5825 (N_5825,N_2045,N_3115);
nor U5826 (N_5826,N_2692,N_3403);
and U5827 (N_5827,N_3007,N_3735);
nor U5828 (N_5828,N_2450,N_3574);
or U5829 (N_5829,N_2852,N_3607);
or U5830 (N_5830,N_3226,N_2423);
and U5831 (N_5831,N_2078,N_2410);
nand U5832 (N_5832,N_3810,N_3171);
and U5833 (N_5833,N_3200,N_3085);
or U5834 (N_5834,N_3940,N_2765);
and U5835 (N_5835,N_3540,N_3647);
and U5836 (N_5836,N_3967,N_2572);
nor U5837 (N_5837,N_3933,N_3127);
nand U5838 (N_5838,N_2301,N_3053);
nor U5839 (N_5839,N_2835,N_2258);
nor U5840 (N_5840,N_2430,N_2935);
nor U5841 (N_5841,N_3356,N_2617);
nor U5842 (N_5842,N_2423,N_2414);
and U5843 (N_5843,N_3698,N_3030);
nand U5844 (N_5844,N_2873,N_3267);
or U5845 (N_5845,N_2408,N_3539);
nor U5846 (N_5846,N_2978,N_2409);
nor U5847 (N_5847,N_3143,N_2791);
nor U5848 (N_5848,N_2393,N_3792);
or U5849 (N_5849,N_3227,N_2909);
nand U5850 (N_5850,N_3351,N_3410);
or U5851 (N_5851,N_3821,N_2491);
nand U5852 (N_5852,N_3611,N_3393);
xor U5853 (N_5853,N_3027,N_3318);
and U5854 (N_5854,N_2614,N_3465);
nor U5855 (N_5855,N_3676,N_2522);
nor U5856 (N_5856,N_2812,N_2761);
and U5857 (N_5857,N_2872,N_2505);
nand U5858 (N_5858,N_2180,N_3963);
and U5859 (N_5859,N_2985,N_3098);
nand U5860 (N_5860,N_3982,N_3932);
nand U5861 (N_5861,N_2879,N_3614);
and U5862 (N_5862,N_2147,N_2430);
and U5863 (N_5863,N_2711,N_3483);
nand U5864 (N_5864,N_2530,N_3887);
or U5865 (N_5865,N_2803,N_2679);
or U5866 (N_5866,N_2830,N_2162);
and U5867 (N_5867,N_2269,N_2416);
and U5868 (N_5868,N_2316,N_3820);
and U5869 (N_5869,N_2446,N_3471);
nand U5870 (N_5870,N_3603,N_3255);
or U5871 (N_5871,N_3573,N_3415);
and U5872 (N_5872,N_3645,N_2580);
or U5873 (N_5873,N_2344,N_3432);
nor U5874 (N_5874,N_2790,N_2019);
nand U5875 (N_5875,N_2065,N_3390);
nor U5876 (N_5876,N_3472,N_3951);
and U5877 (N_5877,N_3860,N_2341);
nand U5878 (N_5878,N_2951,N_3759);
nor U5879 (N_5879,N_3508,N_3829);
or U5880 (N_5880,N_3513,N_2512);
nor U5881 (N_5881,N_2627,N_2296);
or U5882 (N_5882,N_3213,N_3263);
and U5883 (N_5883,N_2248,N_2357);
nand U5884 (N_5884,N_2938,N_2652);
and U5885 (N_5885,N_2294,N_2476);
or U5886 (N_5886,N_2349,N_3625);
nand U5887 (N_5887,N_3364,N_3926);
nand U5888 (N_5888,N_2499,N_3234);
nand U5889 (N_5889,N_3506,N_2633);
nand U5890 (N_5890,N_2010,N_2463);
nor U5891 (N_5891,N_2350,N_2426);
nand U5892 (N_5892,N_2424,N_3805);
or U5893 (N_5893,N_3621,N_3091);
nand U5894 (N_5894,N_3735,N_2452);
nand U5895 (N_5895,N_3509,N_2800);
and U5896 (N_5896,N_3078,N_2960);
or U5897 (N_5897,N_3642,N_3096);
nor U5898 (N_5898,N_3426,N_2417);
and U5899 (N_5899,N_2684,N_3602);
and U5900 (N_5900,N_3299,N_3318);
or U5901 (N_5901,N_3571,N_2097);
nor U5902 (N_5902,N_3241,N_3611);
or U5903 (N_5903,N_2333,N_2988);
nand U5904 (N_5904,N_3627,N_3144);
and U5905 (N_5905,N_2638,N_3047);
nand U5906 (N_5906,N_2313,N_3951);
or U5907 (N_5907,N_2493,N_3157);
or U5908 (N_5908,N_3859,N_2861);
and U5909 (N_5909,N_2641,N_3825);
nor U5910 (N_5910,N_2573,N_2854);
and U5911 (N_5911,N_3634,N_2192);
nand U5912 (N_5912,N_3809,N_2151);
nor U5913 (N_5913,N_3746,N_3096);
nand U5914 (N_5914,N_2844,N_2657);
nand U5915 (N_5915,N_2080,N_3996);
and U5916 (N_5916,N_2836,N_3348);
and U5917 (N_5917,N_2442,N_3438);
and U5918 (N_5918,N_2717,N_2017);
or U5919 (N_5919,N_2542,N_2756);
nor U5920 (N_5920,N_3750,N_3547);
nor U5921 (N_5921,N_2473,N_3723);
nand U5922 (N_5922,N_3091,N_3317);
or U5923 (N_5923,N_3406,N_2215);
and U5924 (N_5924,N_3708,N_2918);
nand U5925 (N_5925,N_2700,N_2176);
nor U5926 (N_5926,N_3587,N_3187);
or U5927 (N_5927,N_3593,N_2240);
and U5928 (N_5928,N_2841,N_3116);
nand U5929 (N_5929,N_2335,N_3908);
and U5930 (N_5930,N_3099,N_2808);
and U5931 (N_5931,N_3661,N_2999);
or U5932 (N_5932,N_2966,N_3287);
or U5933 (N_5933,N_3792,N_2442);
nand U5934 (N_5934,N_3343,N_3825);
or U5935 (N_5935,N_3684,N_3269);
nor U5936 (N_5936,N_2626,N_2103);
nand U5937 (N_5937,N_3426,N_3652);
nand U5938 (N_5938,N_3461,N_3003);
or U5939 (N_5939,N_2245,N_2403);
nand U5940 (N_5940,N_2384,N_2421);
and U5941 (N_5941,N_3256,N_3880);
and U5942 (N_5942,N_3562,N_2415);
or U5943 (N_5943,N_2171,N_3620);
and U5944 (N_5944,N_2826,N_3620);
nand U5945 (N_5945,N_2328,N_3135);
nor U5946 (N_5946,N_3083,N_2530);
and U5947 (N_5947,N_3106,N_3807);
or U5948 (N_5948,N_2353,N_2493);
nand U5949 (N_5949,N_3877,N_2335);
and U5950 (N_5950,N_2702,N_2168);
or U5951 (N_5951,N_2197,N_2893);
or U5952 (N_5952,N_3054,N_2059);
or U5953 (N_5953,N_3817,N_3336);
and U5954 (N_5954,N_3442,N_3537);
nand U5955 (N_5955,N_3348,N_3342);
and U5956 (N_5956,N_2086,N_3233);
and U5957 (N_5957,N_3696,N_2004);
and U5958 (N_5958,N_2560,N_3967);
nand U5959 (N_5959,N_3376,N_2351);
and U5960 (N_5960,N_2527,N_2839);
or U5961 (N_5961,N_2400,N_2001);
nand U5962 (N_5962,N_3032,N_2941);
nand U5963 (N_5963,N_2980,N_3855);
nand U5964 (N_5964,N_2391,N_2790);
nor U5965 (N_5965,N_3341,N_3734);
nor U5966 (N_5966,N_3418,N_3476);
or U5967 (N_5967,N_3447,N_2890);
and U5968 (N_5968,N_3675,N_3826);
or U5969 (N_5969,N_3820,N_2764);
and U5970 (N_5970,N_3598,N_2440);
and U5971 (N_5971,N_3555,N_2625);
nor U5972 (N_5972,N_3940,N_3680);
or U5973 (N_5973,N_3178,N_2355);
and U5974 (N_5974,N_3757,N_2502);
nand U5975 (N_5975,N_2031,N_3946);
nor U5976 (N_5976,N_2229,N_2949);
or U5977 (N_5977,N_3266,N_3142);
nand U5978 (N_5978,N_2384,N_2947);
nor U5979 (N_5979,N_2851,N_3463);
nand U5980 (N_5980,N_2999,N_3219);
nand U5981 (N_5981,N_2383,N_2351);
and U5982 (N_5982,N_2674,N_3635);
and U5983 (N_5983,N_3633,N_2910);
nand U5984 (N_5984,N_2607,N_2097);
or U5985 (N_5985,N_3293,N_2922);
nand U5986 (N_5986,N_3386,N_2746);
nor U5987 (N_5987,N_2397,N_3268);
nand U5988 (N_5988,N_2621,N_3227);
xor U5989 (N_5989,N_3358,N_2139);
or U5990 (N_5990,N_3002,N_2797);
nor U5991 (N_5991,N_2611,N_2248);
or U5992 (N_5992,N_2077,N_3391);
nor U5993 (N_5993,N_3808,N_3113);
and U5994 (N_5994,N_2770,N_2098);
nor U5995 (N_5995,N_3834,N_2147);
and U5996 (N_5996,N_2383,N_3321);
and U5997 (N_5997,N_2827,N_2915);
nor U5998 (N_5998,N_2606,N_2511);
nand U5999 (N_5999,N_3691,N_3163);
or U6000 (N_6000,N_4348,N_5513);
nor U6001 (N_6001,N_5618,N_5966);
nand U6002 (N_6002,N_4145,N_5954);
or U6003 (N_6003,N_5327,N_4117);
nor U6004 (N_6004,N_5294,N_5114);
or U6005 (N_6005,N_5497,N_5910);
nand U6006 (N_6006,N_4116,N_5462);
or U6007 (N_6007,N_4052,N_4974);
or U6008 (N_6008,N_4012,N_5061);
or U6009 (N_6009,N_5325,N_4254);
and U6010 (N_6010,N_4747,N_4204);
or U6011 (N_6011,N_4397,N_4272);
and U6012 (N_6012,N_4139,N_5806);
nor U6013 (N_6013,N_5382,N_5243);
nand U6014 (N_6014,N_5430,N_5745);
and U6015 (N_6015,N_4080,N_5053);
xor U6016 (N_6016,N_4409,N_4276);
and U6017 (N_6017,N_4508,N_4279);
or U6018 (N_6018,N_4487,N_5718);
or U6019 (N_6019,N_5579,N_5669);
nor U6020 (N_6020,N_5581,N_4365);
and U6021 (N_6021,N_5833,N_4362);
and U6022 (N_6022,N_4370,N_5627);
nor U6023 (N_6023,N_5181,N_4283);
or U6024 (N_6024,N_5438,N_5839);
nor U6025 (N_6025,N_5088,N_4374);
nand U6026 (N_6026,N_4024,N_5974);
nor U6027 (N_6027,N_5008,N_4927);
and U6028 (N_6028,N_5595,N_5597);
or U6029 (N_6029,N_4547,N_5388);
nor U6030 (N_6030,N_4431,N_4320);
nand U6031 (N_6031,N_5896,N_4242);
and U6032 (N_6032,N_4767,N_4981);
nand U6033 (N_6033,N_4522,N_5744);
nand U6034 (N_6034,N_4137,N_5429);
nand U6035 (N_6035,N_4349,N_4863);
or U6036 (N_6036,N_4836,N_5561);
or U6037 (N_6037,N_5081,N_4783);
nor U6038 (N_6038,N_5790,N_5856);
nor U6039 (N_6039,N_5370,N_5979);
and U6040 (N_6040,N_5989,N_5862);
nor U6041 (N_6041,N_5242,N_5315);
and U6042 (N_6042,N_4401,N_4147);
or U6043 (N_6043,N_5919,N_5024);
or U6044 (N_6044,N_4623,N_4748);
or U6045 (N_6045,N_5741,N_4607);
nand U6046 (N_6046,N_4909,N_5555);
or U6047 (N_6047,N_4011,N_5336);
and U6048 (N_6048,N_5365,N_4679);
and U6049 (N_6049,N_5940,N_5480);
nor U6050 (N_6050,N_5519,N_4674);
nor U6051 (N_6051,N_5638,N_4962);
and U6052 (N_6052,N_5870,N_4959);
nor U6053 (N_6053,N_4700,N_4448);
nor U6054 (N_6054,N_4449,N_5028);
or U6055 (N_6055,N_4838,N_4288);
nor U6056 (N_6056,N_5076,N_5157);
nand U6057 (N_6057,N_5845,N_5409);
nand U6058 (N_6058,N_4926,N_5149);
nand U6059 (N_6059,N_5252,N_5947);
or U6060 (N_6060,N_4030,N_4219);
and U6061 (N_6061,N_4619,N_4539);
and U6062 (N_6062,N_4026,N_4994);
and U6063 (N_6063,N_5923,N_4657);
and U6064 (N_6064,N_5971,N_5539);
nor U6065 (N_6065,N_5318,N_5861);
nand U6066 (N_6066,N_5660,N_5316);
or U6067 (N_6067,N_5713,N_4692);
nor U6068 (N_6068,N_4207,N_5568);
nor U6069 (N_6069,N_5494,N_4779);
and U6070 (N_6070,N_5363,N_5569);
nor U6071 (N_6071,N_5803,N_4742);
or U6072 (N_6072,N_5355,N_5570);
nor U6073 (N_6073,N_5523,N_4193);
nor U6074 (N_6074,N_4495,N_5554);
or U6075 (N_6075,N_4014,N_4939);
nand U6076 (N_6076,N_5521,N_5460);
nand U6077 (N_6077,N_4354,N_5935);
and U6078 (N_6078,N_5909,N_5606);
nor U6079 (N_6079,N_5714,N_4820);
nand U6080 (N_6080,N_4895,N_5276);
nor U6081 (N_6081,N_5267,N_5587);
or U6082 (N_6082,N_4726,N_4070);
nor U6083 (N_6083,N_4466,N_4109);
and U6084 (N_6084,N_5347,N_5083);
xor U6085 (N_6085,N_5859,N_4424);
nand U6086 (N_6086,N_4652,N_4531);
nor U6087 (N_6087,N_5217,N_4253);
nor U6088 (N_6088,N_5179,N_5021);
nand U6089 (N_6089,N_4339,N_5077);
or U6090 (N_6090,N_5826,N_4453);
or U6091 (N_6091,N_4853,N_4824);
nor U6092 (N_6092,N_5025,N_4074);
and U6093 (N_6093,N_4661,N_4220);
nor U6094 (N_6094,N_5942,N_5485);
nand U6095 (N_6095,N_5778,N_4061);
and U6096 (N_6096,N_5122,N_5377);
nand U6097 (N_6097,N_4690,N_5035);
and U6098 (N_6098,N_5273,N_4650);
nor U6099 (N_6099,N_4319,N_5361);
nand U6100 (N_6100,N_5189,N_4773);
nand U6101 (N_6101,N_5876,N_5257);
or U6102 (N_6102,N_5020,N_4032);
or U6103 (N_6103,N_5868,N_4439);
or U6104 (N_6104,N_4513,N_5216);
and U6105 (N_6105,N_5924,N_4822);
and U6106 (N_6106,N_4544,N_4287);
or U6107 (N_6107,N_5624,N_4901);
nor U6108 (N_6108,N_5586,N_4473);
nand U6109 (N_6109,N_5457,N_5755);
nand U6110 (N_6110,N_5001,N_4073);
and U6111 (N_6111,N_5930,N_5925);
nand U6112 (N_6112,N_5095,N_4442);
and U6113 (N_6113,N_4684,N_4016);
nand U6114 (N_6114,N_5598,N_4815);
and U6115 (N_6115,N_5372,N_5481);
nor U6116 (N_6116,N_5793,N_4251);
nor U6117 (N_6117,N_5702,N_4880);
and U6118 (N_6118,N_5014,N_4878);
nor U6119 (N_6119,N_5248,N_4877);
nand U6120 (N_6120,N_4239,N_5400);
and U6121 (N_6121,N_4372,N_5023);
or U6122 (N_6122,N_4325,N_5982);
and U6123 (N_6123,N_4788,N_4752);
nand U6124 (N_6124,N_4810,N_5373);
nor U6125 (N_6125,N_5929,N_4102);
nor U6126 (N_6126,N_4525,N_4699);
nand U6127 (N_6127,N_5906,N_4617);
nand U6128 (N_6128,N_4977,N_5220);
and U6129 (N_6129,N_5453,N_5708);
nor U6130 (N_6130,N_5013,N_4757);
or U6131 (N_6131,N_4947,N_4993);
nand U6132 (N_6132,N_5685,N_5652);
nand U6133 (N_6133,N_5063,N_5402);
or U6134 (N_6134,N_5734,N_5064);
or U6135 (N_6135,N_4714,N_4867);
or U6136 (N_6136,N_4437,N_4567);
and U6137 (N_6137,N_5324,N_4414);
nand U6138 (N_6138,N_5823,N_4015);
nor U6139 (N_6139,N_5703,N_5849);
nand U6140 (N_6140,N_4955,N_5011);
nor U6141 (N_6141,N_5346,N_4653);
or U6142 (N_6142,N_4092,N_4006);
nand U6143 (N_6143,N_4655,N_5461);
and U6144 (N_6144,N_4645,N_4925);
and U6145 (N_6145,N_5050,N_5293);
nor U6146 (N_6146,N_4526,N_4432);
nor U6147 (N_6147,N_4676,N_4938);
nand U6148 (N_6148,N_4702,N_4605);
nand U6149 (N_6149,N_4184,N_4392);
nand U6150 (N_6150,N_4943,N_4935);
nand U6151 (N_6151,N_5829,N_4924);
or U6152 (N_6152,N_5265,N_5514);
and U6153 (N_6153,N_4769,N_5903);
and U6154 (N_6154,N_4530,N_4045);
nand U6155 (N_6155,N_5807,N_5464);
or U6156 (N_6156,N_5834,N_5368);
or U6157 (N_6157,N_5302,N_4459);
or U6158 (N_6158,N_5697,N_5091);
and U6159 (N_6159,N_4126,N_5663);
nor U6160 (N_6160,N_5976,N_5912);
or U6161 (N_6161,N_4727,N_4274);
and U6162 (N_6162,N_5204,N_5997);
and U6163 (N_6163,N_5477,N_5310);
or U6164 (N_6164,N_5757,N_4507);
or U6165 (N_6165,N_4611,N_4599);
nand U6166 (N_6166,N_4469,N_4851);
and U6167 (N_6167,N_4845,N_5482);
or U6168 (N_6168,N_4464,N_4831);
and U6169 (N_6169,N_5884,N_5214);
or U6170 (N_6170,N_4462,N_4330);
or U6171 (N_6171,N_5374,N_4527);
nor U6172 (N_6172,N_5203,N_4781);
and U6173 (N_6173,N_4436,N_4956);
nor U6174 (N_6174,N_5185,N_5335);
nor U6175 (N_6175,N_5235,N_5719);
nor U6176 (N_6176,N_4375,N_4755);
nor U6177 (N_6177,N_5705,N_4721);
and U6178 (N_6178,N_4160,N_4476);
nor U6179 (N_6179,N_5169,N_4123);
or U6180 (N_6180,N_4166,N_4581);
or U6181 (N_6181,N_4963,N_4310);
nand U6182 (N_6182,N_4896,N_4179);
or U6183 (N_6183,N_5017,N_4686);
and U6184 (N_6184,N_4404,N_5292);
or U6185 (N_6185,N_5193,N_5710);
and U6186 (N_6186,N_4488,N_4717);
nand U6187 (N_6187,N_4989,N_5751);
or U6188 (N_6188,N_5917,N_4558);
or U6189 (N_6189,N_4647,N_4622);
and U6190 (N_6190,N_5977,N_5197);
nand U6191 (N_6191,N_5218,N_4534);
and U6192 (N_6192,N_5754,N_4545);
xor U6193 (N_6193,N_5578,N_5634);
nand U6194 (N_6194,N_4860,N_5175);
nor U6195 (N_6195,N_5244,N_5738);
nor U6196 (N_6196,N_4218,N_5591);
nand U6197 (N_6197,N_4698,N_5796);
nand U6198 (N_6198,N_4398,N_4406);
nor U6199 (N_6199,N_5228,N_5222);
nand U6200 (N_6200,N_5186,N_5413);
nand U6201 (N_6201,N_5147,N_4746);
or U6202 (N_6202,N_4520,N_4814);
nor U6203 (N_6203,N_4990,N_5167);
and U6204 (N_6204,N_5756,N_5448);
and U6205 (N_6205,N_5840,N_5074);
nor U6206 (N_6206,N_4708,N_5852);
nor U6207 (N_6207,N_5678,N_5151);
and U6208 (N_6208,N_5253,N_4793);
and U6209 (N_6209,N_5812,N_4008);
and U6210 (N_6210,N_5145,N_4625);
nand U6211 (N_6211,N_5455,N_4563);
and U6212 (N_6212,N_5677,N_5103);
and U6213 (N_6213,N_5245,N_4723);
or U6214 (N_6214,N_5658,N_4912);
or U6215 (N_6215,N_4130,N_4118);
nand U6216 (N_6216,N_5915,N_4506);
and U6217 (N_6217,N_5854,N_4480);
nand U6218 (N_6218,N_4468,N_5225);
and U6219 (N_6219,N_5015,N_4837);
or U6220 (N_6220,N_4396,N_5306);
or U6221 (N_6221,N_5196,N_5934);
nand U6222 (N_6222,N_5978,N_4969);
or U6223 (N_6223,N_4094,N_5106);
and U6224 (N_6224,N_4445,N_4157);
nor U6225 (N_6225,N_4601,N_4433);
nor U6226 (N_6226,N_5308,N_5951);
nor U6227 (N_6227,N_4856,N_5936);
or U6228 (N_6228,N_4069,N_5067);
and U6229 (N_6229,N_4019,N_4232);
and U6230 (N_6230,N_5736,N_4076);
nor U6231 (N_6231,N_5300,N_4422);
or U6232 (N_6232,N_4483,N_4651);
nor U6233 (N_6233,N_5577,N_5282);
nor U6234 (N_6234,N_5992,N_5715);
and U6235 (N_6235,N_4238,N_4930);
or U6236 (N_6236,N_4311,N_5527);
nor U6237 (N_6237,N_5219,N_5125);
or U6238 (N_6238,N_5297,N_4874);
and U6239 (N_6239,N_4532,N_5511);
nand U6240 (N_6240,N_4825,N_4791);
nand U6241 (N_6241,N_5842,N_4983);
and U6242 (N_6242,N_5055,N_4854);
nand U6243 (N_6243,N_4150,N_5105);
nor U6244 (N_6244,N_4919,N_5544);
or U6245 (N_6245,N_5899,N_4072);
nor U6246 (N_6246,N_4178,N_4371);
or U6247 (N_6247,N_5999,N_5993);
nor U6248 (N_6248,N_4946,N_5068);
nor U6249 (N_6249,N_5501,N_4916);
or U6250 (N_6250,N_5323,N_4022);
and U6251 (N_6251,N_4904,N_5330);
or U6252 (N_6252,N_4865,N_4666);
nor U6253 (N_6253,N_4594,N_5440);
and U6254 (N_6254,N_4753,N_5092);
nor U6255 (N_6255,N_4872,N_5442);
or U6256 (N_6256,N_4040,N_5237);
and U6257 (N_6257,N_4264,N_5616);
or U6258 (N_6258,N_5120,N_4987);
or U6259 (N_6259,N_4952,N_5931);
nand U6260 (N_6260,N_4013,N_4095);
and U6261 (N_6261,N_4380,N_5512);
or U6262 (N_6262,N_4703,N_4941);
nor U6263 (N_6263,N_4479,N_4713);
or U6264 (N_6264,N_4002,N_5952);
nand U6265 (N_6265,N_4028,N_4113);
or U6266 (N_6266,N_4823,N_4082);
or U6267 (N_6267,N_4830,N_4934);
nand U6268 (N_6268,N_4606,N_5117);
nand U6269 (N_6269,N_5637,N_5768);
nand U6270 (N_6270,N_5333,N_4777);
nor U6271 (N_6271,N_5467,N_5726);
nor U6272 (N_6272,N_4988,N_4751);
and U6273 (N_6273,N_5797,N_5838);
nand U6274 (N_6274,N_5644,N_4120);
and U6275 (N_6275,N_5226,N_5969);
or U6276 (N_6276,N_5454,N_4053);
and U6277 (N_6277,N_5277,N_5086);
nand U6278 (N_6278,N_4602,N_5036);
and U6279 (N_6279,N_4195,N_5506);
and U6280 (N_6280,N_5562,N_4451);
nand U6281 (N_6281,N_5148,N_4633);
nand U6282 (N_6282,N_4187,N_4741);
or U6283 (N_6283,N_5988,N_4887);
nor U6284 (N_6284,N_5065,N_5419);
nand U6285 (N_6285,N_4868,N_4472);
nor U6286 (N_6286,N_4675,N_5881);
nor U6287 (N_6287,N_5320,N_5633);
nand U6288 (N_6288,N_5016,N_5609);
and U6289 (N_6289,N_5339,N_4503);
nand U6290 (N_6290,N_5853,N_5321);
nor U6291 (N_6291,N_5352,N_5432);
or U6292 (N_6292,N_4850,N_5835);
nor U6293 (N_6293,N_4629,N_5628);
or U6294 (N_6294,N_4308,N_4143);
nor U6295 (N_6295,N_4639,N_4075);
xor U6296 (N_6296,N_5532,N_4496);
nor U6297 (N_6297,N_4750,N_4132);
or U6298 (N_6298,N_5687,N_5777);
nand U6299 (N_6299,N_5192,N_4801);
nand U6300 (N_6300,N_4050,N_4360);
or U6301 (N_6301,N_4626,N_4720);
nand U6302 (N_6302,N_4331,N_4604);
nand U6303 (N_6303,N_4305,N_5255);
and U6304 (N_6304,N_5572,N_4226);
and U6305 (N_6305,N_5108,N_4548);
nor U6306 (N_6306,N_4097,N_4920);
nand U6307 (N_6307,N_5998,N_4083);
nand U6308 (N_6308,N_5421,N_4897);
nand U6309 (N_6309,N_4124,N_4275);
and U6310 (N_6310,N_5503,N_4217);
nand U6311 (N_6311,N_5588,N_4039);
and U6312 (N_6312,N_5094,N_4847);
and U6313 (N_6313,N_5709,N_4658);
or U6314 (N_6314,N_5201,N_4710);
nor U6315 (N_6315,N_5126,N_5887);
and U6316 (N_6316,N_4636,N_4689);
nor U6317 (N_6317,N_4996,N_5699);
or U6318 (N_6318,N_4500,N_5897);
and U6319 (N_6319,N_5776,N_4376);
or U6320 (N_6320,N_4174,N_5789);
nor U6321 (N_6321,N_4034,N_5371);
nor U6322 (N_6322,N_5066,N_4571);
or U6323 (N_6323,N_5119,N_4486);
nand U6324 (N_6324,N_4267,N_4388);
nand U6325 (N_6325,N_5502,N_4378);
and U6326 (N_6326,N_4361,N_5780);
nor U6327 (N_6327,N_4707,N_4314);
nor U6328 (N_6328,N_5882,N_4366);
nand U6329 (N_6329,N_4010,N_5518);
nand U6330 (N_6330,N_5112,N_4898);
nand U6331 (N_6331,N_5445,N_4294);
and U6332 (N_6332,N_5389,N_5168);
nor U6333 (N_6333,N_5256,N_5855);
nor U6334 (N_6334,N_4728,N_4694);
nand U6335 (N_6335,N_4512,N_4642);
or U6336 (N_6336,N_4031,N_5085);
and U6337 (N_6337,N_4299,N_5760);
nand U6338 (N_6338,N_5163,N_4491);
and U6339 (N_6339,N_5102,N_5417);
or U6340 (N_6340,N_5753,N_4923);
xnor U6341 (N_6341,N_4332,N_4509);
or U6342 (N_6342,N_4345,N_4493);
and U6343 (N_6343,N_4778,N_5720);
or U6344 (N_6344,N_5822,N_4133);
nand U6345 (N_6345,N_5799,N_5921);
nor U6346 (N_6346,N_5766,N_4761);
nand U6347 (N_6347,N_5090,N_4411);
xor U6348 (N_6348,N_4654,N_5913);
nor U6349 (N_6349,N_5198,N_4235);
nand U6350 (N_6350,N_4260,N_4271);
and U6351 (N_6351,N_4862,N_5212);
nor U6352 (N_6352,N_5546,N_4813);
and U6353 (N_6353,N_4816,N_4154);
nor U6354 (N_6354,N_4616,N_5551);
nor U6355 (N_6355,N_4886,N_4301);
nor U6356 (N_6356,N_4986,N_4541);
and U6357 (N_6357,N_4461,N_5392);
nor U6358 (N_6358,N_5968,N_4852);
nand U6359 (N_6359,N_5087,N_5060);
nand U6360 (N_6360,N_5594,N_5810);
or U6361 (N_6361,N_5161,N_5864);
nand U6362 (N_6362,N_5900,N_5611);
xor U6363 (N_6363,N_4044,N_5801);
nor U6364 (N_6364,N_5057,N_5390);
and U6365 (N_6365,N_5704,N_4327);
or U6366 (N_6366,N_4586,N_4682);
nor U6367 (N_6367,N_4960,N_4693);
and U6368 (N_6368,N_5492,N_5284);
nand U6369 (N_6369,N_5963,N_5174);
nor U6370 (N_6370,N_5444,N_4245);
and U6371 (N_6371,N_5111,N_4576);
or U6372 (N_6372,N_5844,N_5183);
xnor U6373 (N_6373,N_5622,N_4389);
xnor U6374 (N_6374,N_5332,N_5836);
nor U6375 (N_6375,N_5537,N_4671);
or U6376 (N_6376,N_5137,N_4200);
or U6377 (N_6377,N_5642,N_5795);
nor U6378 (N_6378,N_4163,N_4900);
or U6379 (N_6379,N_4441,N_5607);
nand U6380 (N_6380,N_4588,N_4165);
or U6381 (N_6381,N_4928,N_5231);
or U6382 (N_6382,N_4368,N_4065);
and U6383 (N_6383,N_5681,N_4447);
nand U6384 (N_6384,N_5961,N_5981);
nand U6385 (N_6385,N_4300,N_4965);
nor U6386 (N_6386,N_4907,N_4551);
or U6387 (N_6387,N_4338,N_5199);
or U6388 (N_6388,N_4931,N_4839);
and U6389 (N_6389,N_5635,N_5716);
or U6390 (N_6390,N_4478,N_5800);
nor U6391 (N_6391,N_5116,N_4049);
and U6392 (N_6392,N_4086,N_5535);
and U6393 (N_6393,N_5426,N_5655);
nand U6394 (N_6394,N_4192,N_4729);
nand U6395 (N_6395,N_4557,N_5348);
and U6396 (N_6396,N_4335,N_5032);
or U6397 (N_6397,N_5779,N_5033);
nand U6398 (N_6398,N_4964,N_4191);
and U6399 (N_6399,N_4701,N_5246);
and U6400 (N_6400,N_5808,N_5617);
nand U6401 (N_6401,N_4776,N_5556);
or U6402 (N_6402,N_5422,N_5656);
or U6403 (N_6403,N_4188,N_4077);
or U6404 (N_6404,N_5124,N_5831);
nand U6405 (N_6405,N_5794,N_4948);
and U6406 (N_6406,N_4434,N_5407);
and U6407 (N_6407,N_4786,N_5908);
and U6408 (N_6408,N_4902,N_4535);
and U6409 (N_6409,N_4662,N_4967);
or U6410 (N_6410,N_4555,N_5960);
and U6411 (N_6411,N_4932,N_4324);
nand U6412 (N_6412,N_5004,N_4937);
nor U6413 (N_6413,N_5888,N_4550);
nand U6414 (N_6414,N_4575,N_5775);
or U6415 (N_6415,N_5949,N_5383);
and U6416 (N_6416,N_5962,N_5058);
nand U6417 (N_6417,N_4377,N_5620);
or U6418 (N_6418,N_4582,N_5410);
nor U6419 (N_6419,N_4756,N_5639);
or U6420 (N_6420,N_5603,N_4246);
nand U6421 (N_6421,N_5843,N_5012);
nand U6422 (N_6422,N_5694,N_5159);
or U6423 (N_6423,N_4664,N_4731);
nor U6424 (N_6424,N_5229,N_5322);
nor U6425 (N_6425,N_4438,N_5397);
nand U6426 (N_6426,N_5973,N_5495);
or U6427 (N_6427,N_4792,N_4190);
nand U6428 (N_6428,N_4189,N_4475);
nor U6429 (N_6429,N_5451,N_5958);
nor U6430 (N_6430,N_4968,N_5580);
or U6431 (N_6431,N_5329,N_4344);
nand U6432 (N_6432,N_5287,N_5459);
nor U6433 (N_6433,N_4185,N_4574);
nand U6434 (N_6434,N_4322,N_5798);
or U6435 (N_6435,N_5643,N_5096);
and U6436 (N_6436,N_4060,N_5007);
and U6437 (N_6437,N_4067,N_5152);
nor U6438 (N_6438,N_4559,N_5414);
nor U6439 (N_6439,N_5805,N_4936);
nor U6440 (N_6440,N_5529,N_4807);
xor U6441 (N_6441,N_5700,N_5260);
or U6442 (N_6442,N_5771,N_4770);
nand U6443 (N_6443,N_5249,N_5251);
nand U6444 (N_6444,N_4585,N_4985);
and U6445 (N_6445,N_5288,N_5084);
nand U6446 (N_6446,N_4966,N_4659);
and U6447 (N_6447,N_5684,N_4161);
nand U6448 (N_6448,N_4614,N_4155);
and U6449 (N_6449,N_5489,N_4443);
nor U6450 (N_6450,N_5964,N_5671);
nor U6451 (N_6451,N_5274,N_4537);
nor U6452 (N_6452,N_4597,N_4600);
or U6453 (N_6453,N_4062,N_5911);
and U6454 (N_6454,N_5530,N_5605);
or U6455 (N_6455,N_4066,N_4316);
or U6456 (N_6456,N_4399,N_4691);
nor U6457 (N_6457,N_4482,N_5268);
or U6458 (N_6458,N_4270,N_5772);
nand U6459 (N_6459,N_4945,N_5943);
and U6460 (N_6460,N_5338,N_4855);
and U6461 (N_6461,N_5747,N_5184);
nor U6462 (N_6462,N_5010,N_4511);
xnor U6463 (N_6463,N_5567,N_4719);
or U6464 (N_6464,N_4148,N_4765);
nand U6465 (N_6465,N_5369,N_5080);
nor U6466 (N_6466,N_5783,N_4128);
or U6467 (N_6467,N_5127,N_4669);
nor U6468 (N_6468,N_5928,N_4259);
nor U6469 (N_6469,N_5224,N_5946);
or U6470 (N_6470,N_5585,N_5098);
and U6471 (N_6471,N_4739,N_4638);
nor U6472 (N_6472,N_4706,N_4549);
or U6473 (N_6473,N_5038,N_5679);
or U6474 (N_6474,N_5926,N_5047);
and U6475 (N_6475,N_4307,N_4467);
and U6476 (N_6476,N_5405,N_4334);
or U6477 (N_6477,N_4353,N_5877);
nor U6478 (N_6478,N_4819,N_4857);
or U6479 (N_6479,N_5782,N_4416);
nor U6480 (N_6480,N_4716,N_5337);
and U6481 (N_6481,N_5456,N_5233);
nor U6482 (N_6482,N_5848,N_5404);
nand U6483 (N_6483,N_4228,N_5841);
xor U6484 (N_6484,N_5176,N_5984);
nor U6485 (N_6485,N_5526,N_4269);
nor U6486 (N_6486,N_5416,N_4367);
and U6487 (N_6487,N_4673,N_4603);
nand U6488 (N_6488,N_5412,N_4685);
and U6489 (N_6489,N_4352,N_5764);
nor U6490 (N_6490,N_4151,N_5664);
nor U6491 (N_6491,N_5990,N_4805);
and U6492 (N_6492,N_5955,N_5904);
and U6493 (N_6493,N_4291,N_4250);
nor U6494 (N_6494,N_4997,N_5211);
or U6495 (N_6495,N_5089,N_4430);
or U6496 (N_6496,N_4042,N_4859);
or U6497 (N_6497,N_5263,N_4734);
nand U6498 (N_6498,N_4890,N_5515);
nand U6499 (N_6499,N_5230,N_5686);
nand U6500 (N_6500,N_4538,N_5724);
xor U6501 (N_6501,N_4340,N_5496);
nor U6502 (N_6502,N_5858,N_5072);
nor U6503 (N_6503,N_4180,N_4091);
nand U6504 (N_6504,N_5173,N_4420);
xor U6505 (N_6505,N_5781,N_5815);
or U6506 (N_6506,N_5309,N_5816);
nand U6507 (N_6507,N_5393,N_5427);
nand U6508 (N_6508,N_4152,N_4950);
and U6509 (N_6509,N_5970,N_5136);
nor U6510 (N_6510,N_4056,N_4304);
nor U6511 (N_6511,N_5941,N_4216);
nand U6512 (N_6512,N_5259,N_4921);
or U6513 (N_6513,N_5584,N_4224);
nand U6514 (N_6514,N_4210,N_4982);
nor U6515 (N_6515,N_4223,N_4146);
nand U6516 (N_6516,N_5463,N_5784);
and U6517 (N_6517,N_4518,N_5360);
nor U6518 (N_6518,N_4172,N_5592);
nor U6519 (N_6519,N_4632,N_4568);
nor U6520 (N_6520,N_4450,N_5140);
nor U6521 (N_6521,N_4884,N_4681);
and U6522 (N_6522,N_4976,N_4593);
nand U6523 (N_6523,N_4517,N_4231);
and U6524 (N_6524,N_5286,N_5610);
and U6525 (N_6525,N_5927,N_4875);
or U6526 (N_6526,N_5051,N_4408);
nor U6527 (N_6527,N_4381,N_5509);
and U6528 (N_6528,N_5118,N_4656);
nand U6529 (N_6529,N_4648,N_5396);
and U6530 (N_6530,N_5391,N_4168);
and U6531 (N_6531,N_5227,N_4005);
nand U6532 (N_6532,N_5510,N_4630);
and U6533 (N_6533,N_4444,N_4917);
nor U6534 (N_6534,N_4589,N_5746);
and U6535 (N_6535,N_5533,N_4543);
or U6536 (N_6536,N_5436,N_4615);
or U6537 (N_6537,N_4709,N_4252);
or U6538 (N_6538,N_5860,N_4149);
nor U6539 (N_6539,N_5340,N_4159);
and U6540 (N_6540,N_4782,N_4230);
or U6541 (N_6541,N_5558,N_5517);
and U6542 (N_6542,N_5825,N_4802);
and U6543 (N_6543,N_4999,N_4961);
or U6544 (N_6544,N_4027,N_4759);
or U6545 (N_6545,N_5027,N_4055);
and U6546 (N_6546,N_4735,N_4315);
and U6547 (N_6547,N_4725,N_4302);
nand U6548 (N_6548,N_4227,N_5948);
or U6549 (N_6549,N_5589,N_4081);
and U6550 (N_6550,N_5654,N_5264);
xnor U6551 (N_6551,N_5767,N_5447);
or U6552 (N_6552,N_5524,N_4899);
nor U6553 (N_6553,N_5632,N_4763);
and U6554 (N_6554,N_4524,N_4176);
nand U6555 (N_6555,N_4114,N_4347);
xnor U6556 (N_6556,N_4129,N_4336);
or U6557 (N_6557,N_5564,N_5814);
nor U6558 (N_6558,N_5049,N_4737);
nor U6559 (N_6559,N_5215,N_5944);
and U6560 (N_6560,N_4196,N_5765);
and U6561 (N_6561,N_4809,N_5353);
nor U6562 (N_6562,N_4047,N_4812);
nand U6563 (N_6563,N_4182,N_4456);
and U6564 (N_6564,N_5141,N_4323);
or U6565 (N_6565,N_5680,N_4084);
nand U6566 (N_6566,N_5345,N_4394);
and U6567 (N_6567,N_5006,N_5623);
or U6568 (N_6568,N_4208,N_5626);
and U6569 (N_6569,N_5701,N_5266);
nor U6570 (N_6570,N_5894,N_5641);
nor U6571 (N_6571,N_4905,N_5648);
or U6572 (N_6572,N_5596,N_4265);
and U6573 (N_6573,N_4222,N_5600);
nand U6574 (N_6574,N_4112,N_5194);
and U6575 (N_6575,N_5202,N_5824);
nand U6576 (N_6576,N_5073,N_4670);
and U6577 (N_6577,N_5560,N_4817);
or U6578 (N_6578,N_4046,N_4268);
nand U6579 (N_6579,N_5547,N_5059);
or U6580 (N_6580,N_4215,N_4870);
and U6581 (N_6581,N_5221,N_4906);
nor U6582 (N_6582,N_4089,N_4806);
nor U6583 (N_6583,N_4313,N_4552);
and U6584 (N_6584,N_5062,N_4293);
nor U6585 (N_6585,N_5791,N_4018);
nand U6586 (N_6586,N_4333,N_5557);
or U6587 (N_6587,N_5662,N_5439);
nor U6588 (N_6588,N_5743,N_5078);
or U6589 (N_6589,N_5905,N_4672);
nand U6590 (N_6590,N_5450,N_5953);
nor U6591 (N_6591,N_5657,N_5239);
and U6592 (N_6592,N_5508,N_4321);
nor U6593 (N_6593,N_4458,N_5434);
nand U6594 (N_6594,N_5313,N_4797);
nand U6595 (N_6595,N_5543,N_4641);
and U6596 (N_6596,N_5957,N_4828);
xnor U6597 (N_6597,N_4794,N_4958);
nand U6598 (N_6598,N_5357,N_5727);
nor U6599 (N_6599,N_4297,N_5281);
and U6600 (N_6600,N_4282,N_4627);
or U6601 (N_6601,N_4583,N_5907);
or U6602 (N_6602,N_5376,N_5759);
and U6603 (N_6603,N_5364,N_4186);
or U6604 (N_6604,N_5541,N_5150);
and U6605 (N_6605,N_4804,N_4631);
and U6606 (N_6606,N_5155,N_4980);
nand U6607 (N_6607,N_5138,N_5299);
and U6608 (N_6608,N_5991,N_4871);
nor U6609 (N_6609,N_4312,N_5487);
nand U6610 (N_6610,N_4020,N_5182);
nand U6611 (N_6611,N_4608,N_5188);
nand U6612 (N_6612,N_5980,N_4385);
or U6613 (N_6613,N_5732,N_5162);
and U6614 (N_6614,N_4384,N_5731);
nor U6615 (N_6615,N_5811,N_4876);
nand U6616 (N_6616,N_4490,N_4973);
nor U6617 (N_6617,N_4667,N_5254);
nand U6618 (N_6618,N_5056,N_5354);
nand U6619 (N_6619,N_4350,N_5180);
or U6620 (N_6620,N_5387,N_5420);
or U6621 (N_6621,N_4455,N_5104);
and U6622 (N_6622,N_4848,N_4564);
and U6623 (N_6623,N_5739,N_4835);
or U6624 (N_6624,N_5937,N_5030);
xnor U6625 (N_6625,N_5769,N_5466);
and U6626 (N_6626,N_4104,N_4068);
nand U6627 (N_6627,N_4100,N_5240);
nor U6628 (N_6628,N_5695,N_5446);
and U6629 (N_6629,N_5415,N_4021);
or U6630 (N_6630,N_5041,N_5075);
and U6631 (N_6631,N_5082,N_4866);
and U6632 (N_6632,N_4383,N_5054);
xor U6633 (N_6633,N_5207,N_4212);
or U6634 (N_6634,N_4953,N_5291);
nand U6635 (N_6635,N_5334,N_5717);
nand U6636 (N_6636,N_4356,N_4922);
and U6637 (N_6637,N_4369,N_4036);
or U6638 (N_6638,N_5378,N_4292);
nor U6639 (N_6639,N_5195,N_5331);
or U6640 (N_6640,N_4954,N_4079);
xnor U6641 (N_6641,N_4740,N_5762);
nand U6642 (N_6642,N_5002,N_4043);
nand U6643 (N_6643,N_5563,N_5933);
nand U6644 (N_6644,N_4127,N_4843);
or U6645 (N_6645,N_4306,N_4979);
or U6646 (N_6646,N_4529,N_4144);
nor U6647 (N_6647,N_5763,N_5191);
and U6648 (N_6648,N_4382,N_5548);
nor U6649 (N_6649,N_5311,N_5034);
or U6650 (N_6650,N_5590,N_4749);
or U6651 (N_6651,N_5153,N_5465);
nor U6652 (N_6652,N_4419,N_4596);
or U6653 (N_6653,N_4425,N_4914);
or U6654 (N_6654,N_5499,N_4101);
and U6655 (N_6655,N_5536,N_5305);
nand U6656 (N_6656,N_4093,N_4379);
and U6657 (N_6657,N_4829,N_5200);
nor U6658 (N_6658,N_5540,N_4273);
and U6659 (N_6659,N_4266,N_4435);
and U6660 (N_6660,N_5742,N_4844);
nand U6661 (N_6661,N_4821,N_4678);
nor U6662 (N_6662,N_4796,N_4704);
or U6663 (N_6663,N_4463,N_5351);
and U6664 (N_6664,N_4775,N_5735);
nand U6665 (N_6665,N_5343,N_5009);
nand U6666 (N_6666,N_4908,N_4054);
nand U6667 (N_6667,N_4351,N_5614);
nand U6668 (N_6668,N_4744,N_4136);
nor U6669 (N_6669,N_4718,N_4784);
or U6670 (N_6670,N_4164,N_4494);
nand U6671 (N_6671,N_5269,N_4454);
nor U6672 (N_6672,N_5278,N_4957);
and U6673 (N_6673,N_5918,N_4612);
and U6674 (N_6674,N_4236,N_5965);
nand U6675 (N_6675,N_4167,N_4465);
nand U6676 (N_6676,N_4918,N_5786);
nor U6677 (N_6677,N_5576,N_4004);
nor U6678 (N_6678,N_4841,N_4284);
and U6679 (N_6679,N_5139,N_5135);
xor U6680 (N_6680,N_5832,N_4099);
nand U6681 (N_6681,N_5223,N_5433);
nand U6682 (N_6682,N_4911,N_5468);
and U6683 (N_6683,N_4485,N_5052);
and U6684 (N_6684,N_4995,N_5398);
or U6685 (N_6685,N_4038,N_5728);
nand U6686 (N_6686,N_4158,N_5785);
nand U6687 (N_6687,N_4470,N_5093);
nor U6688 (N_6688,N_5690,N_4110);
and U6689 (N_6689,N_5885,N_5863);
or U6690 (N_6690,N_4405,N_4402);
xnor U6691 (N_6691,N_5956,N_5069);
and U6692 (N_6692,N_5711,N_4426);
or U6693 (N_6693,N_5018,N_5707);
nor U6694 (N_6694,N_4799,N_5131);
and U6695 (N_6695,N_4029,N_4722);
or U6696 (N_6696,N_4342,N_4971);
nand U6697 (N_6697,N_4785,N_5653);
xor U6698 (N_6698,N_5344,N_5406);
nor U6699 (N_6699,N_5646,N_4277);
and U6700 (N_6700,N_4309,N_5939);
nor U6701 (N_6701,N_5630,N_4197);
nor U6702 (N_6702,N_4649,N_4885);
and U6703 (N_6703,N_5166,N_5883);
nor U6704 (N_6704,N_5621,N_5381);
and U6705 (N_6705,N_5470,N_4141);
xnor U6706 (N_6706,N_4233,N_5042);
nand U6707 (N_6707,N_5250,N_5241);
and U6708 (N_6708,N_4764,N_4400);
nor U6709 (N_6709,N_5865,N_4849);
or U6710 (N_6710,N_4888,N_5932);
and U6711 (N_6711,N_5208,N_5000);
nor U6712 (N_6712,N_5403,N_4663);
or U6713 (N_6713,N_4628,N_5488);
nand U6714 (N_6714,N_4942,N_4359);
or U6715 (N_6715,N_4107,N_4944);
nor U6716 (N_6716,N_4562,N_5079);
nor U6717 (N_6717,N_4007,N_5820);
or U6718 (N_6718,N_5129,N_5319);
or U6719 (N_6719,N_5851,N_5258);
nand U6720 (N_6720,N_5867,N_5817);
nand U6721 (N_6721,N_4523,N_4579);
nand U6722 (N_6722,N_4337,N_5234);
nor U6723 (N_6723,N_4554,N_5566);
and U6724 (N_6724,N_5819,N_5675);
and U6725 (N_6725,N_4680,N_5994);
nand U6726 (N_6726,N_4194,N_5328);
nand U6727 (N_6727,N_4051,N_5522);
nand U6728 (N_6728,N_5818,N_5366);
nor U6729 (N_6729,N_5706,N_5100);
xnor U6730 (N_6730,N_5553,N_4637);
and U6731 (N_6731,N_5938,N_5608);
or U6732 (N_6732,N_5528,N_4162);
or U6733 (N_6733,N_5471,N_5493);
nor U6734 (N_6734,N_4240,N_4280);
nand U6735 (N_6735,N_5359,N_5437);
or U6736 (N_6736,N_5983,N_4000);
nand U6737 (N_6737,N_4546,N_5871);
nor U6738 (N_6738,N_4156,N_5478);
nor U6739 (N_6739,N_5737,N_4078);
and U6740 (N_6740,N_4712,N_5401);
nand U6741 (N_6741,N_4281,N_5425);
nor U6742 (N_6742,N_4566,N_4991);
and U6743 (N_6743,N_4115,N_5484);
nor U6744 (N_6744,N_5029,N_5483);
nand U6745 (N_6745,N_5170,N_5809);
nor U6746 (N_6746,N_5538,N_5748);
or U6747 (N_6747,N_4153,N_5171);
nand U6748 (N_6748,N_5692,N_4774);
and U6749 (N_6749,N_4428,N_4285);
and U6750 (N_6750,N_5891,N_5435);
nor U6751 (N_6751,N_5123,N_4592);
and U6752 (N_6752,N_5945,N_5879);
or U6753 (N_6753,N_5682,N_4504);
nand U6754 (N_6754,N_4992,N_4131);
or U6755 (N_6755,N_5996,N_4640);
nand U6756 (N_6756,N_4861,N_5550);
nand U6757 (N_6757,N_5665,N_5975);
or U6758 (N_6758,N_5574,N_5295);
and U6759 (N_6759,N_5670,N_4064);
and U6760 (N_6760,N_4440,N_5914);
nor U6761 (N_6761,N_4811,N_4800);
nor U6762 (N_6762,N_4346,N_4766);
nor U6763 (N_6763,N_5443,N_5847);
and U6764 (N_6764,N_5270,N_5046);
nand U6765 (N_6765,N_5474,N_5458);
nor U6766 (N_6766,N_4386,N_5044);
nor U6767 (N_6767,N_5723,N_4471);
nand U6768 (N_6768,N_5895,N_4057);
and U6769 (N_6769,N_4417,N_4243);
nand U6770 (N_6770,N_4893,N_4125);
nor U6771 (N_6771,N_4929,N_5285);
nor U6772 (N_6772,N_4058,N_4715);
nor U6773 (N_6773,N_4017,N_5395);
nand U6774 (N_6774,N_5985,N_4025);
and U6775 (N_6775,N_5599,N_4577);
or U6776 (N_6776,N_5133,N_5326);
and U6777 (N_6777,N_4474,N_5261);
nor U6778 (N_6778,N_5486,N_5649);
and U6779 (N_6779,N_5730,N_5901);
nand U6780 (N_6780,N_4387,N_5721);
and U6781 (N_6781,N_5613,N_4695);
nand U6782 (N_6782,N_5296,N_4170);
nand U6783 (N_6783,N_4827,N_5650);
nand U6784 (N_6784,N_4119,N_4041);
or U6785 (N_6785,N_4578,N_5750);
nor U6786 (N_6786,N_5615,N_5629);
nand U6787 (N_6787,N_4477,N_4003);
nand U6788 (N_6788,N_5101,N_5418);
and U6789 (N_6789,N_5232,N_4403);
or U6790 (N_6790,N_4913,N_5473);
and U6791 (N_6791,N_4668,N_4364);
and U6792 (N_6792,N_4949,N_4889);
nor U6793 (N_6793,N_5206,N_4289);
or U6794 (N_6794,N_4970,N_4978);
nor U6795 (N_6795,N_5950,N_5972);
or U6796 (N_6796,N_4933,N_4533);
nand U6797 (N_6797,N_4221,N_5107);
and U6798 (N_6798,N_5298,N_4733);
nand U6799 (N_6799,N_5573,N_4135);
nor U6800 (N_6800,N_5733,N_5156);
nor U6801 (N_6801,N_5729,N_4001);
nand U6802 (N_6802,N_4858,N_5475);
nand U6803 (N_6803,N_5802,N_4317);
nand U6804 (N_6804,N_4169,N_5916);
and U6805 (N_6805,N_5275,N_4951);
nor U6806 (N_6806,N_5431,N_4758);
or U6807 (N_6807,N_5099,N_5172);
or U6808 (N_6808,N_5602,N_5280);
or U6809 (N_6809,N_5872,N_5889);
and U6810 (N_6810,N_5469,N_4105);
nor U6811 (N_6811,N_5749,N_5110);
and U6812 (N_6812,N_5898,N_5774);
nor U6813 (N_6813,N_4063,N_4111);
or U6814 (N_6814,N_5869,N_4290);
nand U6815 (N_6815,N_4096,N_4229);
or U6816 (N_6816,N_4569,N_5037);
nor U6817 (N_6817,N_4711,N_4413);
nor U6818 (N_6818,N_4643,N_5142);
or U6819 (N_6819,N_5850,N_5830);
nand U6820 (N_6820,N_5031,N_4808);
nand U6821 (N_6821,N_5379,N_4318);
or U6822 (N_6822,N_4201,N_5279);
nand U6823 (N_6823,N_4696,N_4609);
nand U6824 (N_6824,N_4787,N_5048);
and U6825 (N_6825,N_5071,N_4358);
and U6826 (N_6826,N_4610,N_5674);
nand U6827 (N_6827,N_5476,N_5375);
and U6828 (N_6828,N_5143,N_4059);
or U6829 (N_6829,N_4121,N_4998);
or U6830 (N_6830,N_5902,N_5583);
nand U6831 (N_6831,N_5666,N_5892);
xor U6832 (N_6832,N_4572,N_4972);
or U6833 (N_6833,N_5045,N_4891);
or U6834 (N_6834,N_4528,N_4211);
nor U6835 (N_6835,N_4181,N_4457);
and U6836 (N_6836,N_4071,N_5428);
and U6837 (N_6837,N_4869,N_4515);
and U6838 (N_6838,N_5132,N_5575);
nor U6839 (N_6839,N_5209,N_4789);
and U6840 (N_6840,N_4199,N_5612);
nand U6841 (N_6841,N_5504,N_4561);
and U6842 (N_6842,N_4536,N_4138);
nor U6843 (N_6843,N_5205,N_5314);
and U6844 (N_6844,N_4501,N_4248);
or U6845 (N_6845,N_5283,N_4140);
or U6846 (N_6846,N_5312,N_4621);
and U6847 (N_6847,N_4296,N_4122);
nor U6848 (N_6848,N_4915,N_5349);
and U6849 (N_6849,N_4832,N_5121);
nand U6850 (N_6850,N_5647,N_5271);
nor U6851 (N_6851,N_4598,N_4343);
and U6852 (N_6852,N_4035,N_4037);
nand U6853 (N_6853,N_4206,N_5097);
and U6854 (N_6854,N_5317,N_5828);
nor U6855 (N_6855,N_4183,N_5113);
or U6856 (N_6856,N_5827,N_4446);
nor U6857 (N_6857,N_4743,N_4590);
nor U6858 (N_6858,N_5604,N_4261);
or U6859 (N_6859,N_5022,N_4570);
nand U6860 (N_6860,N_4171,N_4298);
and U6861 (N_6861,N_4175,N_5238);
nand U6862 (N_6862,N_5676,N_4754);
nand U6863 (N_6863,N_4882,N_4730);
nor U6864 (N_6864,N_4452,N_4412);
or U6865 (N_6865,N_4573,N_4634);
and U6866 (N_6866,N_5289,N_5441);
nand U6867 (N_6867,N_5262,N_5165);
nor U6868 (N_6868,N_5673,N_4618);
nor U6869 (N_6869,N_4881,N_4328);
and U6870 (N_6870,N_4418,N_4697);
nor U6871 (N_6871,N_4879,N_4732);
nor U6872 (N_6872,N_4103,N_4833);
and U6873 (N_6873,N_4873,N_5026);
nor U6874 (N_6874,N_5893,N_4247);
nand U6875 (N_6875,N_4940,N_5247);
nor U6876 (N_6876,N_5134,N_5384);
nor U6877 (N_6877,N_5890,N_4745);
or U6878 (N_6878,N_4591,N_5307);
or U6879 (N_6879,N_5667,N_5507);
and U6880 (N_6880,N_5959,N_4249);
and U6881 (N_6881,N_4108,N_4492);
or U6882 (N_6882,N_5631,N_4363);
and U6883 (N_6883,N_4214,N_4098);
or U6884 (N_6884,N_4198,N_5154);
or U6885 (N_6885,N_4768,N_4357);
nand U6886 (N_6886,N_4427,N_5866);
nand U6887 (N_6887,N_5761,N_5571);
nor U6888 (N_6888,N_4497,N_5804);
nor U6889 (N_6889,N_5472,N_4481);
or U6890 (N_6890,N_5003,N_4234);
or U6891 (N_6891,N_5995,N_5693);
or U6892 (N_6892,N_5813,N_5236);
and U6893 (N_6893,N_5668,N_5040);
nand U6894 (N_6894,N_5967,N_5423);
nor U6895 (N_6895,N_5770,N_5424);
nand U6896 (N_6896,N_5559,N_4262);
or U6897 (N_6897,N_4624,N_4258);
and U6898 (N_6898,N_5130,N_4278);
and U6899 (N_6899,N_4771,N_5873);
nand U6900 (N_6900,N_5019,N_4106);
or U6901 (N_6901,N_4407,N_4263);
nor U6902 (N_6902,N_4256,N_5342);
nor U6903 (N_6903,N_5787,N_4516);
nor U6904 (N_6904,N_4635,N_4209);
or U6905 (N_6905,N_4795,N_5399);
nor U6906 (N_6906,N_4203,N_5362);
nand U6907 (N_6907,N_5683,N_4177);
or U6908 (N_6908,N_5210,N_4205);
and U6909 (N_6909,N_5187,N_4087);
nand U6910 (N_6910,N_5109,N_4738);
and U6911 (N_6911,N_5531,N_5449);
nand U6912 (N_6912,N_4090,N_5986);
nand U6913 (N_6913,N_5651,N_5725);
or U6914 (N_6914,N_5479,N_4894);
and U6915 (N_6915,N_4225,N_5846);
and U6916 (N_6916,N_5886,N_4724);
nor U6917 (N_6917,N_4213,N_4423);
or U6918 (N_6918,N_5158,N_5408);
nand U6919 (N_6919,N_5490,N_5696);
nor U6920 (N_6920,N_5625,N_4910);
and U6921 (N_6921,N_5500,N_4683);
or U6922 (N_6922,N_5880,N_4565);
and U6923 (N_6923,N_4780,N_5070);
or U6924 (N_6924,N_5146,N_4142);
and U6925 (N_6925,N_5452,N_5115);
or U6926 (N_6926,N_5758,N_4736);
nand U6927 (N_6927,N_5792,N_5688);
nand U6928 (N_6928,N_5356,N_4790);
and U6929 (N_6929,N_4903,N_5837);
nor U6930 (N_6930,N_4772,N_5301);
nand U6931 (N_6931,N_4846,N_5178);
nor U6932 (N_6932,N_5712,N_5659);
and U6933 (N_6933,N_4510,N_5385);
or U6934 (N_6934,N_4255,N_4803);
and U6935 (N_6935,N_5636,N_4644);
and U6936 (N_6936,N_5689,N_4975);
nand U6937 (N_6937,N_5672,N_4237);
and U6938 (N_6938,N_5542,N_5043);
nor U6939 (N_6939,N_5788,N_5177);
or U6940 (N_6940,N_5358,N_4984);
nor U6941 (N_6941,N_5645,N_4033);
or U6942 (N_6942,N_4355,N_4329);
nand U6943 (N_6943,N_4286,N_4134);
or U6944 (N_6944,N_4760,N_5160);
and U6945 (N_6945,N_4415,N_5367);
or U6946 (N_6946,N_4341,N_5857);
and U6947 (N_6947,N_5565,N_5722);
nor U6948 (N_6948,N_4677,N_4514);
xor U6949 (N_6949,N_4244,N_5534);
or U6950 (N_6950,N_5773,N_5752);
or U6951 (N_6951,N_5005,N_4421);
nand U6952 (N_6952,N_4620,N_5878);
and U6953 (N_6953,N_5516,N_4241);
and U6954 (N_6954,N_4326,N_4818);
or U6955 (N_6955,N_4390,N_5987);
nand U6956 (N_6956,N_5619,N_4303);
nor U6957 (N_6957,N_4009,N_4410);
nor U6958 (N_6958,N_4864,N_5303);
and U6959 (N_6959,N_5593,N_4429);
or U6960 (N_6960,N_5304,N_5290);
or U6961 (N_6961,N_5640,N_5164);
nor U6962 (N_6962,N_4883,N_5505);
nor U6963 (N_6963,N_4688,N_4646);
or U6964 (N_6964,N_5691,N_5386);
or U6965 (N_6965,N_5582,N_5698);
nor U6966 (N_6966,N_4391,N_5491);
nand U6967 (N_6967,N_5545,N_4665);
nor U6968 (N_6968,N_5875,N_4553);
or U6969 (N_6969,N_4393,N_5411);
nor U6970 (N_6970,N_4173,N_5549);
nand U6971 (N_6971,N_4484,N_4519);
and U6972 (N_6972,N_5213,N_5601);
nor U6973 (N_6973,N_4595,N_4257);
nor U6974 (N_6974,N_4798,N_4202);
nor U6975 (N_6975,N_4834,N_4705);
nand U6976 (N_6976,N_5920,N_4395);
and U6977 (N_6977,N_5821,N_4762);
nor U6978 (N_6978,N_4542,N_4023);
or U6979 (N_6979,N_4540,N_4373);
or U6980 (N_6980,N_4687,N_5394);
or U6981 (N_6981,N_4580,N_4499);
nor U6982 (N_6982,N_5525,N_4460);
or U6983 (N_6983,N_5039,N_4613);
nand U6984 (N_6984,N_4088,N_4048);
and U6985 (N_6985,N_5341,N_4489);
nand U6986 (N_6986,N_4840,N_4560);
and U6987 (N_6987,N_4502,N_5498);
nor U6988 (N_6988,N_5190,N_4587);
and U6989 (N_6989,N_5350,N_4892);
nor U6990 (N_6990,N_4085,N_5922);
and U6991 (N_6991,N_4505,N_4842);
nor U6992 (N_6992,N_5552,N_5874);
nand U6993 (N_6993,N_4660,N_5380);
and U6994 (N_6994,N_5272,N_4498);
or U6995 (N_6995,N_4826,N_5520);
nor U6996 (N_6996,N_4295,N_5740);
and U6997 (N_6997,N_5661,N_5128);
and U6998 (N_6998,N_4556,N_4521);
and U6999 (N_6999,N_5144,N_4584);
and U7000 (N_7000,N_5821,N_4369);
or U7001 (N_7001,N_4875,N_5955);
xor U7002 (N_7002,N_4641,N_5701);
nand U7003 (N_7003,N_5678,N_4495);
nor U7004 (N_7004,N_4964,N_5647);
nor U7005 (N_7005,N_4869,N_4803);
and U7006 (N_7006,N_5077,N_5272);
nand U7007 (N_7007,N_5662,N_4429);
or U7008 (N_7008,N_4484,N_4248);
and U7009 (N_7009,N_4670,N_5449);
or U7010 (N_7010,N_4864,N_4588);
nor U7011 (N_7011,N_4026,N_4485);
or U7012 (N_7012,N_5672,N_4796);
and U7013 (N_7013,N_5932,N_4140);
and U7014 (N_7014,N_4845,N_4245);
and U7015 (N_7015,N_5487,N_5585);
nor U7016 (N_7016,N_4095,N_4659);
nand U7017 (N_7017,N_5252,N_5321);
nor U7018 (N_7018,N_5940,N_5363);
nand U7019 (N_7019,N_5333,N_5585);
nor U7020 (N_7020,N_4694,N_4253);
and U7021 (N_7021,N_5599,N_4664);
nand U7022 (N_7022,N_5543,N_5106);
and U7023 (N_7023,N_4689,N_4147);
nor U7024 (N_7024,N_4317,N_5422);
nand U7025 (N_7025,N_4698,N_5299);
nand U7026 (N_7026,N_5596,N_5233);
nand U7027 (N_7027,N_4930,N_4979);
nand U7028 (N_7028,N_4851,N_4383);
nor U7029 (N_7029,N_5390,N_4039);
or U7030 (N_7030,N_4701,N_4958);
and U7031 (N_7031,N_4587,N_5160);
and U7032 (N_7032,N_4744,N_5842);
nor U7033 (N_7033,N_4266,N_5994);
nor U7034 (N_7034,N_5200,N_5680);
and U7035 (N_7035,N_4138,N_5814);
or U7036 (N_7036,N_5167,N_5637);
nand U7037 (N_7037,N_4283,N_5345);
or U7038 (N_7038,N_4585,N_5573);
and U7039 (N_7039,N_5769,N_4889);
and U7040 (N_7040,N_5217,N_4518);
nor U7041 (N_7041,N_4408,N_4307);
nand U7042 (N_7042,N_4898,N_5198);
and U7043 (N_7043,N_5536,N_4924);
nand U7044 (N_7044,N_5424,N_5160);
or U7045 (N_7045,N_4270,N_5113);
and U7046 (N_7046,N_4497,N_4869);
and U7047 (N_7047,N_4230,N_4766);
or U7048 (N_7048,N_5898,N_4204);
nor U7049 (N_7049,N_5364,N_4594);
and U7050 (N_7050,N_5035,N_4763);
nand U7051 (N_7051,N_4409,N_5399);
nand U7052 (N_7052,N_4766,N_4360);
nor U7053 (N_7053,N_4612,N_5499);
or U7054 (N_7054,N_4226,N_5037);
and U7055 (N_7055,N_5674,N_4938);
or U7056 (N_7056,N_4762,N_5865);
and U7057 (N_7057,N_5158,N_4473);
and U7058 (N_7058,N_4303,N_4012);
and U7059 (N_7059,N_5208,N_4151);
or U7060 (N_7060,N_5609,N_5988);
or U7061 (N_7061,N_5502,N_4327);
or U7062 (N_7062,N_4526,N_4209);
nand U7063 (N_7063,N_4308,N_5262);
or U7064 (N_7064,N_4440,N_4487);
and U7065 (N_7065,N_4699,N_5074);
or U7066 (N_7066,N_5350,N_5637);
and U7067 (N_7067,N_4852,N_4614);
or U7068 (N_7068,N_4734,N_4528);
and U7069 (N_7069,N_5506,N_5247);
nor U7070 (N_7070,N_5591,N_5505);
nor U7071 (N_7071,N_5695,N_4081);
nand U7072 (N_7072,N_5343,N_5896);
and U7073 (N_7073,N_4859,N_5192);
or U7074 (N_7074,N_4415,N_4174);
and U7075 (N_7075,N_4593,N_5505);
and U7076 (N_7076,N_5687,N_5249);
and U7077 (N_7077,N_5375,N_4980);
and U7078 (N_7078,N_5362,N_5414);
nor U7079 (N_7079,N_5115,N_4205);
nand U7080 (N_7080,N_4924,N_5568);
and U7081 (N_7081,N_5478,N_4540);
and U7082 (N_7082,N_5344,N_4530);
or U7083 (N_7083,N_4370,N_4945);
nor U7084 (N_7084,N_5362,N_4466);
nor U7085 (N_7085,N_4564,N_4384);
nand U7086 (N_7086,N_5730,N_4506);
and U7087 (N_7087,N_4263,N_5818);
nor U7088 (N_7088,N_5391,N_5595);
and U7089 (N_7089,N_5856,N_5187);
xnor U7090 (N_7090,N_5936,N_5618);
or U7091 (N_7091,N_5262,N_4980);
nand U7092 (N_7092,N_4774,N_5588);
and U7093 (N_7093,N_5153,N_5963);
and U7094 (N_7094,N_4602,N_5325);
nor U7095 (N_7095,N_5155,N_4342);
nand U7096 (N_7096,N_4363,N_4975);
and U7097 (N_7097,N_4846,N_5212);
nand U7098 (N_7098,N_4236,N_4048);
nand U7099 (N_7099,N_4910,N_4543);
or U7100 (N_7100,N_4315,N_5741);
and U7101 (N_7101,N_4943,N_4228);
and U7102 (N_7102,N_4994,N_5847);
nor U7103 (N_7103,N_4758,N_4556);
nand U7104 (N_7104,N_4098,N_5279);
or U7105 (N_7105,N_4880,N_5474);
nor U7106 (N_7106,N_5707,N_4171);
or U7107 (N_7107,N_4668,N_5567);
and U7108 (N_7108,N_4819,N_4799);
nand U7109 (N_7109,N_4731,N_5898);
nand U7110 (N_7110,N_5122,N_5330);
and U7111 (N_7111,N_4032,N_4544);
nor U7112 (N_7112,N_5400,N_5489);
nand U7113 (N_7113,N_5740,N_4509);
nand U7114 (N_7114,N_5737,N_4225);
or U7115 (N_7115,N_5783,N_5239);
nand U7116 (N_7116,N_5614,N_5706);
or U7117 (N_7117,N_5579,N_5067);
nand U7118 (N_7118,N_4334,N_4745);
or U7119 (N_7119,N_5387,N_4301);
and U7120 (N_7120,N_4599,N_5345);
nand U7121 (N_7121,N_4284,N_4771);
nor U7122 (N_7122,N_4744,N_4498);
nand U7123 (N_7123,N_4762,N_5247);
nand U7124 (N_7124,N_5193,N_5541);
or U7125 (N_7125,N_4199,N_4983);
nor U7126 (N_7126,N_4271,N_4261);
nor U7127 (N_7127,N_4362,N_4758);
and U7128 (N_7128,N_5215,N_5319);
and U7129 (N_7129,N_4346,N_5560);
nor U7130 (N_7130,N_5644,N_4331);
or U7131 (N_7131,N_4342,N_5949);
nor U7132 (N_7132,N_5730,N_4745);
or U7133 (N_7133,N_4624,N_5109);
nor U7134 (N_7134,N_4228,N_4458);
or U7135 (N_7135,N_4974,N_4157);
xor U7136 (N_7136,N_4044,N_4689);
and U7137 (N_7137,N_5044,N_4127);
nor U7138 (N_7138,N_4288,N_5340);
nand U7139 (N_7139,N_4143,N_4891);
and U7140 (N_7140,N_4334,N_5106);
and U7141 (N_7141,N_5819,N_4667);
or U7142 (N_7142,N_5782,N_5628);
nand U7143 (N_7143,N_5263,N_4887);
nand U7144 (N_7144,N_4792,N_4817);
or U7145 (N_7145,N_5236,N_5572);
nand U7146 (N_7146,N_5028,N_4377);
nor U7147 (N_7147,N_4728,N_4989);
nand U7148 (N_7148,N_4912,N_4628);
nor U7149 (N_7149,N_5858,N_4347);
nor U7150 (N_7150,N_4265,N_4666);
or U7151 (N_7151,N_5222,N_5007);
and U7152 (N_7152,N_5503,N_4080);
nand U7153 (N_7153,N_4237,N_4602);
nand U7154 (N_7154,N_4310,N_4006);
and U7155 (N_7155,N_5491,N_4906);
and U7156 (N_7156,N_4254,N_5529);
or U7157 (N_7157,N_5650,N_5486);
nand U7158 (N_7158,N_4701,N_4117);
and U7159 (N_7159,N_5870,N_5430);
and U7160 (N_7160,N_5399,N_5587);
nand U7161 (N_7161,N_4158,N_4379);
or U7162 (N_7162,N_5337,N_4833);
or U7163 (N_7163,N_4329,N_5065);
nand U7164 (N_7164,N_5623,N_5370);
or U7165 (N_7165,N_4636,N_5451);
and U7166 (N_7166,N_4241,N_5315);
nor U7167 (N_7167,N_4077,N_5428);
nor U7168 (N_7168,N_5854,N_4584);
or U7169 (N_7169,N_5241,N_5028);
nand U7170 (N_7170,N_5838,N_4263);
nand U7171 (N_7171,N_4505,N_5356);
and U7172 (N_7172,N_4670,N_5224);
nand U7173 (N_7173,N_4721,N_5740);
xor U7174 (N_7174,N_5291,N_5056);
nand U7175 (N_7175,N_4670,N_5050);
nor U7176 (N_7176,N_4389,N_4240);
nand U7177 (N_7177,N_4287,N_4767);
and U7178 (N_7178,N_4074,N_5632);
and U7179 (N_7179,N_5262,N_5714);
nand U7180 (N_7180,N_5952,N_4485);
or U7181 (N_7181,N_4525,N_4077);
nor U7182 (N_7182,N_4945,N_5898);
nand U7183 (N_7183,N_5757,N_4552);
nor U7184 (N_7184,N_5072,N_4425);
nand U7185 (N_7185,N_5973,N_4659);
nor U7186 (N_7186,N_5972,N_5710);
nand U7187 (N_7187,N_5119,N_5950);
and U7188 (N_7188,N_4785,N_4946);
nand U7189 (N_7189,N_4823,N_4436);
or U7190 (N_7190,N_4347,N_4235);
nor U7191 (N_7191,N_4225,N_4235);
and U7192 (N_7192,N_4382,N_5793);
nand U7193 (N_7193,N_4820,N_4311);
nand U7194 (N_7194,N_5394,N_5873);
and U7195 (N_7195,N_4751,N_4277);
or U7196 (N_7196,N_5307,N_4651);
or U7197 (N_7197,N_5673,N_4837);
and U7198 (N_7198,N_4052,N_4934);
nand U7199 (N_7199,N_4361,N_4821);
nand U7200 (N_7200,N_5486,N_4413);
nand U7201 (N_7201,N_4934,N_5785);
and U7202 (N_7202,N_5592,N_4399);
or U7203 (N_7203,N_4850,N_5843);
nand U7204 (N_7204,N_4426,N_4083);
nand U7205 (N_7205,N_4933,N_4476);
nor U7206 (N_7206,N_5840,N_5813);
or U7207 (N_7207,N_5598,N_4012);
and U7208 (N_7208,N_4121,N_4248);
nor U7209 (N_7209,N_5172,N_4012);
nand U7210 (N_7210,N_4244,N_4438);
nand U7211 (N_7211,N_4929,N_5159);
or U7212 (N_7212,N_5645,N_5614);
nor U7213 (N_7213,N_4091,N_5595);
nor U7214 (N_7214,N_4067,N_4265);
nor U7215 (N_7215,N_5801,N_4480);
and U7216 (N_7216,N_5902,N_5038);
nand U7217 (N_7217,N_4439,N_5095);
nand U7218 (N_7218,N_4777,N_5339);
and U7219 (N_7219,N_5590,N_5697);
nand U7220 (N_7220,N_4991,N_5511);
or U7221 (N_7221,N_5771,N_5363);
nor U7222 (N_7222,N_4179,N_4959);
nand U7223 (N_7223,N_4117,N_5325);
or U7224 (N_7224,N_4643,N_5110);
nor U7225 (N_7225,N_5592,N_5577);
nor U7226 (N_7226,N_4704,N_4423);
and U7227 (N_7227,N_4661,N_4988);
or U7228 (N_7228,N_5148,N_4968);
or U7229 (N_7229,N_5994,N_4770);
and U7230 (N_7230,N_4172,N_4575);
nand U7231 (N_7231,N_5794,N_4326);
or U7232 (N_7232,N_4682,N_4177);
nand U7233 (N_7233,N_5100,N_4689);
nand U7234 (N_7234,N_4520,N_4087);
and U7235 (N_7235,N_4368,N_5671);
or U7236 (N_7236,N_4610,N_5123);
or U7237 (N_7237,N_5892,N_5328);
nand U7238 (N_7238,N_5646,N_4854);
nand U7239 (N_7239,N_5422,N_5444);
or U7240 (N_7240,N_4414,N_5583);
and U7241 (N_7241,N_5782,N_4039);
or U7242 (N_7242,N_5481,N_4518);
nand U7243 (N_7243,N_5420,N_4338);
nor U7244 (N_7244,N_5746,N_5661);
and U7245 (N_7245,N_5280,N_5962);
or U7246 (N_7246,N_4051,N_5629);
nand U7247 (N_7247,N_5584,N_5886);
or U7248 (N_7248,N_5812,N_5541);
nor U7249 (N_7249,N_4482,N_5132);
nor U7250 (N_7250,N_5626,N_4047);
or U7251 (N_7251,N_4028,N_5675);
nand U7252 (N_7252,N_4085,N_4653);
and U7253 (N_7253,N_5643,N_4463);
and U7254 (N_7254,N_5975,N_5840);
nor U7255 (N_7255,N_5174,N_5240);
or U7256 (N_7256,N_5910,N_4534);
nor U7257 (N_7257,N_4514,N_4157);
and U7258 (N_7258,N_5848,N_4756);
and U7259 (N_7259,N_5135,N_4471);
nand U7260 (N_7260,N_5050,N_4399);
nor U7261 (N_7261,N_5693,N_5910);
or U7262 (N_7262,N_4862,N_5073);
nand U7263 (N_7263,N_4888,N_5989);
nor U7264 (N_7264,N_5276,N_5860);
or U7265 (N_7265,N_5421,N_4409);
or U7266 (N_7266,N_4102,N_4277);
and U7267 (N_7267,N_5417,N_4580);
nand U7268 (N_7268,N_4754,N_5947);
nand U7269 (N_7269,N_5641,N_4390);
nor U7270 (N_7270,N_5442,N_5440);
nor U7271 (N_7271,N_5547,N_5496);
or U7272 (N_7272,N_5987,N_5599);
or U7273 (N_7273,N_4975,N_4156);
nor U7274 (N_7274,N_4802,N_4603);
nand U7275 (N_7275,N_5589,N_4489);
xor U7276 (N_7276,N_5117,N_4407);
nor U7277 (N_7277,N_5958,N_4909);
or U7278 (N_7278,N_5609,N_5863);
or U7279 (N_7279,N_5518,N_5036);
nor U7280 (N_7280,N_5539,N_5324);
nor U7281 (N_7281,N_5830,N_4465);
or U7282 (N_7282,N_5728,N_5643);
or U7283 (N_7283,N_4851,N_5495);
and U7284 (N_7284,N_5920,N_4828);
nand U7285 (N_7285,N_4825,N_5422);
and U7286 (N_7286,N_4656,N_4385);
nand U7287 (N_7287,N_4088,N_5070);
or U7288 (N_7288,N_4096,N_4781);
or U7289 (N_7289,N_5511,N_5316);
and U7290 (N_7290,N_4004,N_5030);
nand U7291 (N_7291,N_4767,N_4635);
and U7292 (N_7292,N_4426,N_4068);
or U7293 (N_7293,N_4352,N_4070);
nor U7294 (N_7294,N_5044,N_4757);
nand U7295 (N_7295,N_5934,N_4712);
nand U7296 (N_7296,N_4806,N_4870);
or U7297 (N_7297,N_5906,N_5849);
or U7298 (N_7298,N_5922,N_4214);
nand U7299 (N_7299,N_5024,N_5680);
and U7300 (N_7300,N_5710,N_4791);
and U7301 (N_7301,N_4507,N_5592);
and U7302 (N_7302,N_4916,N_4128);
and U7303 (N_7303,N_5905,N_4980);
nand U7304 (N_7304,N_4244,N_4578);
and U7305 (N_7305,N_4504,N_5720);
nor U7306 (N_7306,N_4184,N_4594);
or U7307 (N_7307,N_5838,N_4429);
nand U7308 (N_7308,N_5955,N_5564);
and U7309 (N_7309,N_5871,N_5854);
nand U7310 (N_7310,N_5969,N_5081);
or U7311 (N_7311,N_4497,N_4887);
nor U7312 (N_7312,N_4091,N_4354);
nand U7313 (N_7313,N_5104,N_5532);
nand U7314 (N_7314,N_4442,N_5107);
nor U7315 (N_7315,N_5104,N_5142);
nor U7316 (N_7316,N_5521,N_5060);
nand U7317 (N_7317,N_4770,N_4258);
nand U7318 (N_7318,N_4815,N_4493);
nand U7319 (N_7319,N_5258,N_5646);
and U7320 (N_7320,N_4440,N_4337);
and U7321 (N_7321,N_4468,N_5949);
nor U7322 (N_7322,N_5406,N_4677);
or U7323 (N_7323,N_4640,N_4592);
and U7324 (N_7324,N_4350,N_5639);
and U7325 (N_7325,N_5151,N_4825);
and U7326 (N_7326,N_4921,N_4532);
nor U7327 (N_7327,N_5136,N_4617);
and U7328 (N_7328,N_4183,N_5901);
or U7329 (N_7329,N_4781,N_5996);
or U7330 (N_7330,N_5305,N_4406);
nand U7331 (N_7331,N_5302,N_5993);
nor U7332 (N_7332,N_4676,N_5159);
and U7333 (N_7333,N_5054,N_5877);
or U7334 (N_7334,N_5675,N_5456);
nand U7335 (N_7335,N_4128,N_5832);
nor U7336 (N_7336,N_5037,N_5311);
nor U7337 (N_7337,N_5862,N_5071);
or U7338 (N_7338,N_5627,N_4985);
nor U7339 (N_7339,N_4174,N_4148);
and U7340 (N_7340,N_4420,N_4615);
nor U7341 (N_7341,N_4416,N_4126);
nor U7342 (N_7342,N_4506,N_4669);
nor U7343 (N_7343,N_5649,N_5237);
and U7344 (N_7344,N_4224,N_4370);
or U7345 (N_7345,N_4886,N_5634);
and U7346 (N_7346,N_4269,N_4356);
nand U7347 (N_7347,N_5946,N_5401);
and U7348 (N_7348,N_5865,N_5801);
nand U7349 (N_7349,N_5081,N_5835);
nor U7350 (N_7350,N_4584,N_4986);
nand U7351 (N_7351,N_5837,N_4783);
nand U7352 (N_7352,N_4077,N_5250);
and U7353 (N_7353,N_5160,N_5498);
nand U7354 (N_7354,N_4106,N_5015);
xor U7355 (N_7355,N_4568,N_4138);
xnor U7356 (N_7356,N_5840,N_4243);
nand U7357 (N_7357,N_4526,N_5995);
nand U7358 (N_7358,N_5771,N_5726);
nor U7359 (N_7359,N_5198,N_5661);
and U7360 (N_7360,N_4156,N_4960);
and U7361 (N_7361,N_5410,N_5839);
nor U7362 (N_7362,N_4655,N_4160);
nand U7363 (N_7363,N_4945,N_5791);
or U7364 (N_7364,N_4773,N_4246);
and U7365 (N_7365,N_5213,N_4003);
nand U7366 (N_7366,N_4114,N_5258);
or U7367 (N_7367,N_4744,N_5287);
and U7368 (N_7368,N_4175,N_5156);
nand U7369 (N_7369,N_4159,N_4517);
and U7370 (N_7370,N_4991,N_4969);
nor U7371 (N_7371,N_4750,N_4096);
and U7372 (N_7372,N_5596,N_5053);
nor U7373 (N_7373,N_5885,N_5047);
and U7374 (N_7374,N_4975,N_4453);
nor U7375 (N_7375,N_5154,N_4454);
nor U7376 (N_7376,N_4481,N_4838);
nor U7377 (N_7377,N_5599,N_5558);
nor U7378 (N_7378,N_5042,N_4093);
nor U7379 (N_7379,N_5878,N_5392);
nor U7380 (N_7380,N_5704,N_5532);
nor U7381 (N_7381,N_4189,N_4652);
or U7382 (N_7382,N_4668,N_5020);
and U7383 (N_7383,N_4242,N_5887);
and U7384 (N_7384,N_4338,N_5001);
nand U7385 (N_7385,N_5046,N_5751);
nor U7386 (N_7386,N_5707,N_5413);
nand U7387 (N_7387,N_5292,N_4446);
or U7388 (N_7388,N_5907,N_4955);
nor U7389 (N_7389,N_4021,N_5772);
nand U7390 (N_7390,N_5835,N_4993);
and U7391 (N_7391,N_4597,N_5892);
and U7392 (N_7392,N_5715,N_5202);
and U7393 (N_7393,N_4076,N_4501);
and U7394 (N_7394,N_4960,N_5203);
and U7395 (N_7395,N_5059,N_4262);
nand U7396 (N_7396,N_5210,N_5208);
or U7397 (N_7397,N_4159,N_4260);
nand U7398 (N_7398,N_5473,N_4906);
or U7399 (N_7399,N_4185,N_5254);
or U7400 (N_7400,N_5815,N_5375);
and U7401 (N_7401,N_5145,N_4698);
nand U7402 (N_7402,N_5269,N_5055);
and U7403 (N_7403,N_5373,N_4503);
and U7404 (N_7404,N_4753,N_4787);
nand U7405 (N_7405,N_5405,N_5271);
and U7406 (N_7406,N_5456,N_4356);
nand U7407 (N_7407,N_4125,N_5769);
or U7408 (N_7408,N_5514,N_4644);
nand U7409 (N_7409,N_5387,N_5911);
or U7410 (N_7410,N_4814,N_4922);
and U7411 (N_7411,N_4243,N_5266);
or U7412 (N_7412,N_5288,N_4059);
nor U7413 (N_7413,N_4827,N_5311);
nand U7414 (N_7414,N_4581,N_5468);
or U7415 (N_7415,N_4768,N_4183);
nor U7416 (N_7416,N_5048,N_4694);
or U7417 (N_7417,N_5913,N_5491);
or U7418 (N_7418,N_4524,N_4801);
nand U7419 (N_7419,N_4382,N_4203);
or U7420 (N_7420,N_4949,N_5901);
and U7421 (N_7421,N_4592,N_5395);
and U7422 (N_7422,N_5063,N_5514);
and U7423 (N_7423,N_5689,N_4453);
nor U7424 (N_7424,N_4032,N_4292);
and U7425 (N_7425,N_5943,N_5807);
or U7426 (N_7426,N_5617,N_4959);
and U7427 (N_7427,N_5449,N_5549);
and U7428 (N_7428,N_4597,N_5679);
nand U7429 (N_7429,N_4243,N_4770);
and U7430 (N_7430,N_5345,N_4734);
nand U7431 (N_7431,N_4154,N_5157);
and U7432 (N_7432,N_4910,N_5760);
nor U7433 (N_7433,N_5157,N_4507);
nand U7434 (N_7434,N_5304,N_5905);
or U7435 (N_7435,N_4740,N_4561);
nor U7436 (N_7436,N_4497,N_5369);
and U7437 (N_7437,N_5564,N_5544);
nor U7438 (N_7438,N_4058,N_5437);
nand U7439 (N_7439,N_4345,N_4389);
or U7440 (N_7440,N_4083,N_4551);
and U7441 (N_7441,N_4289,N_5376);
or U7442 (N_7442,N_4789,N_4122);
and U7443 (N_7443,N_5267,N_4883);
or U7444 (N_7444,N_5349,N_4928);
or U7445 (N_7445,N_5281,N_5300);
or U7446 (N_7446,N_5487,N_5462);
nand U7447 (N_7447,N_5793,N_4522);
nand U7448 (N_7448,N_5020,N_4559);
nand U7449 (N_7449,N_4407,N_4790);
and U7450 (N_7450,N_5397,N_5728);
nor U7451 (N_7451,N_4562,N_4698);
or U7452 (N_7452,N_4977,N_4709);
or U7453 (N_7453,N_4251,N_5322);
nor U7454 (N_7454,N_5771,N_5525);
nor U7455 (N_7455,N_5098,N_4716);
nand U7456 (N_7456,N_4253,N_4322);
nand U7457 (N_7457,N_5735,N_4286);
or U7458 (N_7458,N_4546,N_5299);
or U7459 (N_7459,N_5739,N_5426);
nor U7460 (N_7460,N_5867,N_5723);
or U7461 (N_7461,N_4212,N_4569);
nor U7462 (N_7462,N_5325,N_5254);
nand U7463 (N_7463,N_4123,N_5314);
and U7464 (N_7464,N_5175,N_5147);
nor U7465 (N_7465,N_5335,N_4533);
or U7466 (N_7466,N_5154,N_5116);
nor U7467 (N_7467,N_5677,N_5410);
nor U7468 (N_7468,N_5972,N_5802);
or U7469 (N_7469,N_4500,N_4315);
nor U7470 (N_7470,N_5001,N_4704);
and U7471 (N_7471,N_4815,N_4570);
nand U7472 (N_7472,N_4968,N_5888);
or U7473 (N_7473,N_5651,N_5760);
and U7474 (N_7474,N_5114,N_5403);
or U7475 (N_7475,N_5870,N_4035);
nand U7476 (N_7476,N_5177,N_5875);
and U7477 (N_7477,N_5061,N_4798);
nand U7478 (N_7478,N_4772,N_4326);
or U7479 (N_7479,N_4741,N_5235);
and U7480 (N_7480,N_4808,N_5026);
nor U7481 (N_7481,N_5698,N_4911);
nand U7482 (N_7482,N_4831,N_5496);
nor U7483 (N_7483,N_4865,N_4293);
and U7484 (N_7484,N_4386,N_5370);
and U7485 (N_7485,N_5148,N_5818);
and U7486 (N_7486,N_4873,N_5155);
nor U7487 (N_7487,N_4562,N_5420);
nor U7488 (N_7488,N_5520,N_5951);
and U7489 (N_7489,N_5333,N_5038);
and U7490 (N_7490,N_4842,N_4801);
and U7491 (N_7491,N_5039,N_4893);
or U7492 (N_7492,N_4893,N_5488);
or U7493 (N_7493,N_5499,N_4457);
and U7494 (N_7494,N_5753,N_4140);
nor U7495 (N_7495,N_5263,N_4369);
nand U7496 (N_7496,N_4176,N_5414);
and U7497 (N_7497,N_5453,N_4348);
or U7498 (N_7498,N_4032,N_4907);
nor U7499 (N_7499,N_4936,N_4620);
nand U7500 (N_7500,N_5066,N_4344);
or U7501 (N_7501,N_4131,N_4291);
nor U7502 (N_7502,N_5438,N_5524);
or U7503 (N_7503,N_5789,N_5254);
nor U7504 (N_7504,N_4992,N_5529);
nor U7505 (N_7505,N_4637,N_5022);
nor U7506 (N_7506,N_4091,N_4300);
or U7507 (N_7507,N_5534,N_4353);
nor U7508 (N_7508,N_5462,N_4713);
nor U7509 (N_7509,N_4177,N_4854);
nor U7510 (N_7510,N_5646,N_4853);
or U7511 (N_7511,N_5922,N_4965);
or U7512 (N_7512,N_5740,N_5501);
nor U7513 (N_7513,N_4540,N_4068);
nor U7514 (N_7514,N_5725,N_4748);
nand U7515 (N_7515,N_4748,N_5544);
and U7516 (N_7516,N_5633,N_4003);
xor U7517 (N_7517,N_4913,N_5888);
nand U7518 (N_7518,N_5140,N_4923);
and U7519 (N_7519,N_5760,N_5965);
and U7520 (N_7520,N_5028,N_4101);
or U7521 (N_7521,N_4814,N_5359);
nand U7522 (N_7522,N_4822,N_4700);
nor U7523 (N_7523,N_5366,N_4616);
or U7524 (N_7524,N_5554,N_5898);
nand U7525 (N_7525,N_5890,N_5501);
nand U7526 (N_7526,N_4155,N_5112);
nand U7527 (N_7527,N_5710,N_4693);
nor U7528 (N_7528,N_4148,N_5463);
or U7529 (N_7529,N_5204,N_5297);
nand U7530 (N_7530,N_4596,N_4996);
nor U7531 (N_7531,N_5420,N_4763);
or U7532 (N_7532,N_5135,N_4287);
or U7533 (N_7533,N_4677,N_4538);
or U7534 (N_7534,N_5361,N_4486);
nand U7535 (N_7535,N_5573,N_5764);
nand U7536 (N_7536,N_4329,N_5869);
nand U7537 (N_7537,N_5437,N_5759);
or U7538 (N_7538,N_5911,N_5454);
nor U7539 (N_7539,N_4289,N_5880);
and U7540 (N_7540,N_5339,N_4765);
or U7541 (N_7541,N_4231,N_5377);
nor U7542 (N_7542,N_5874,N_4959);
nor U7543 (N_7543,N_5470,N_5703);
nand U7544 (N_7544,N_4301,N_4752);
nor U7545 (N_7545,N_4909,N_4798);
nor U7546 (N_7546,N_5394,N_5775);
or U7547 (N_7547,N_5216,N_5023);
nor U7548 (N_7548,N_5581,N_5278);
nand U7549 (N_7549,N_5992,N_4861);
nor U7550 (N_7550,N_4937,N_5564);
and U7551 (N_7551,N_4260,N_4037);
and U7552 (N_7552,N_5026,N_4855);
or U7553 (N_7553,N_4116,N_5271);
nand U7554 (N_7554,N_5023,N_5321);
nor U7555 (N_7555,N_4781,N_5359);
nor U7556 (N_7556,N_5258,N_5619);
nor U7557 (N_7557,N_5820,N_4154);
nand U7558 (N_7558,N_4306,N_4462);
or U7559 (N_7559,N_5123,N_5686);
and U7560 (N_7560,N_5952,N_5532);
nor U7561 (N_7561,N_4281,N_5374);
or U7562 (N_7562,N_4403,N_4955);
nand U7563 (N_7563,N_5395,N_4198);
nor U7564 (N_7564,N_5819,N_4939);
and U7565 (N_7565,N_4059,N_5368);
nor U7566 (N_7566,N_5631,N_5708);
and U7567 (N_7567,N_4354,N_4523);
nand U7568 (N_7568,N_4607,N_4797);
and U7569 (N_7569,N_5505,N_5997);
or U7570 (N_7570,N_5642,N_5836);
and U7571 (N_7571,N_4683,N_4468);
nor U7572 (N_7572,N_4117,N_5035);
nand U7573 (N_7573,N_5975,N_5734);
and U7574 (N_7574,N_4125,N_5687);
nand U7575 (N_7575,N_4530,N_5345);
and U7576 (N_7576,N_4070,N_4019);
and U7577 (N_7577,N_4916,N_4858);
or U7578 (N_7578,N_5528,N_4565);
nor U7579 (N_7579,N_5518,N_4835);
or U7580 (N_7580,N_5485,N_5526);
nand U7581 (N_7581,N_4344,N_4632);
or U7582 (N_7582,N_5534,N_4847);
and U7583 (N_7583,N_4604,N_5840);
nand U7584 (N_7584,N_5520,N_4241);
or U7585 (N_7585,N_4084,N_4649);
or U7586 (N_7586,N_4118,N_5041);
or U7587 (N_7587,N_4135,N_5198);
nand U7588 (N_7588,N_5554,N_5707);
and U7589 (N_7589,N_4253,N_4935);
and U7590 (N_7590,N_4956,N_5482);
or U7591 (N_7591,N_5853,N_5124);
or U7592 (N_7592,N_5628,N_4971);
or U7593 (N_7593,N_5393,N_4189);
nor U7594 (N_7594,N_4939,N_5271);
and U7595 (N_7595,N_4226,N_5197);
nand U7596 (N_7596,N_4138,N_5957);
nand U7597 (N_7597,N_5702,N_5032);
or U7598 (N_7598,N_4238,N_5175);
nor U7599 (N_7599,N_5125,N_4770);
or U7600 (N_7600,N_4646,N_4660);
nor U7601 (N_7601,N_5540,N_4839);
or U7602 (N_7602,N_5491,N_5289);
xnor U7603 (N_7603,N_4768,N_5575);
or U7604 (N_7604,N_4098,N_4734);
nor U7605 (N_7605,N_4754,N_5673);
nor U7606 (N_7606,N_4776,N_5028);
and U7607 (N_7607,N_4497,N_4493);
nor U7608 (N_7608,N_4789,N_5458);
nor U7609 (N_7609,N_4166,N_4448);
and U7610 (N_7610,N_5136,N_4490);
and U7611 (N_7611,N_4880,N_5201);
nor U7612 (N_7612,N_5182,N_4045);
or U7613 (N_7613,N_4052,N_4312);
xnor U7614 (N_7614,N_4959,N_4098);
nor U7615 (N_7615,N_4222,N_5003);
and U7616 (N_7616,N_5041,N_5162);
and U7617 (N_7617,N_4218,N_5953);
nand U7618 (N_7618,N_4766,N_5720);
or U7619 (N_7619,N_4137,N_5106);
nor U7620 (N_7620,N_4458,N_4214);
nand U7621 (N_7621,N_4260,N_4034);
nand U7622 (N_7622,N_5577,N_5612);
nand U7623 (N_7623,N_5610,N_4297);
nor U7624 (N_7624,N_5062,N_5104);
and U7625 (N_7625,N_4335,N_4400);
nor U7626 (N_7626,N_4967,N_5046);
and U7627 (N_7627,N_4843,N_4456);
nor U7628 (N_7628,N_5750,N_5079);
or U7629 (N_7629,N_4950,N_5234);
and U7630 (N_7630,N_5443,N_4490);
nand U7631 (N_7631,N_4168,N_5498);
or U7632 (N_7632,N_5498,N_5360);
and U7633 (N_7633,N_4258,N_4819);
nor U7634 (N_7634,N_4489,N_5647);
and U7635 (N_7635,N_5593,N_5285);
and U7636 (N_7636,N_5787,N_4707);
nand U7637 (N_7637,N_4789,N_5928);
or U7638 (N_7638,N_5985,N_5649);
or U7639 (N_7639,N_5722,N_4455);
or U7640 (N_7640,N_5436,N_5409);
and U7641 (N_7641,N_4493,N_4565);
nand U7642 (N_7642,N_5440,N_5853);
nor U7643 (N_7643,N_5714,N_4557);
nand U7644 (N_7644,N_5608,N_5075);
nor U7645 (N_7645,N_5943,N_5443);
nand U7646 (N_7646,N_5788,N_4575);
nor U7647 (N_7647,N_5995,N_4327);
and U7648 (N_7648,N_4590,N_5871);
or U7649 (N_7649,N_5913,N_5712);
and U7650 (N_7650,N_5988,N_5806);
nor U7651 (N_7651,N_4404,N_4926);
nand U7652 (N_7652,N_4222,N_4748);
nand U7653 (N_7653,N_5025,N_5958);
nor U7654 (N_7654,N_5948,N_5403);
nor U7655 (N_7655,N_4122,N_4480);
and U7656 (N_7656,N_5191,N_5299);
nand U7657 (N_7657,N_5038,N_4668);
nor U7658 (N_7658,N_5509,N_5407);
nor U7659 (N_7659,N_4075,N_5524);
nor U7660 (N_7660,N_5501,N_5703);
nand U7661 (N_7661,N_5403,N_4042);
or U7662 (N_7662,N_5890,N_5396);
nand U7663 (N_7663,N_5959,N_4395);
nand U7664 (N_7664,N_5891,N_4800);
or U7665 (N_7665,N_4020,N_5880);
and U7666 (N_7666,N_5926,N_5214);
nand U7667 (N_7667,N_4573,N_5054);
nand U7668 (N_7668,N_5399,N_4414);
nor U7669 (N_7669,N_4527,N_4834);
and U7670 (N_7670,N_5320,N_5259);
nand U7671 (N_7671,N_4043,N_5357);
or U7672 (N_7672,N_4872,N_4463);
and U7673 (N_7673,N_5440,N_5654);
nand U7674 (N_7674,N_5794,N_5789);
or U7675 (N_7675,N_5564,N_4717);
nand U7676 (N_7676,N_5130,N_5521);
and U7677 (N_7677,N_4637,N_4921);
nand U7678 (N_7678,N_5574,N_5387);
nor U7679 (N_7679,N_5151,N_5853);
nand U7680 (N_7680,N_4932,N_5243);
or U7681 (N_7681,N_4481,N_4081);
nor U7682 (N_7682,N_4850,N_5733);
nor U7683 (N_7683,N_4102,N_4757);
nor U7684 (N_7684,N_5369,N_5197);
or U7685 (N_7685,N_4661,N_5121);
and U7686 (N_7686,N_4044,N_4865);
or U7687 (N_7687,N_5686,N_5998);
and U7688 (N_7688,N_5697,N_5058);
nand U7689 (N_7689,N_4614,N_4621);
or U7690 (N_7690,N_5765,N_4798);
nand U7691 (N_7691,N_5814,N_4517);
and U7692 (N_7692,N_4954,N_5804);
nand U7693 (N_7693,N_4001,N_4547);
nor U7694 (N_7694,N_5972,N_5673);
or U7695 (N_7695,N_4401,N_4635);
and U7696 (N_7696,N_5840,N_5297);
nand U7697 (N_7697,N_4402,N_4057);
and U7698 (N_7698,N_4692,N_4459);
and U7699 (N_7699,N_5811,N_4836);
or U7700 (N_7700,N_5246,N_4137);
nand U7701 (N_7701,N_4968,N_4502);
nand U7702 (N_7702,N_4192,N_4884);
nor U7703 (N_7703,N_5779,N_4340);
nor U7704 (N_7704,N_4201,N_4442);
or U7705 (N_7705,N_4106,N_4263);
or U7706 (N_7706,N_4520,N_4145);
nand U7707 (N_7707,N_4390,N_4551);
or U7708 (N_7708,N_5733,N_4924);
nor U7709 (N_7709,N_5816,N_5728);
and U7710 (N_7710,N_4098,N_4529);
or U7711 (N_7711,N_5400,N_5575);
nand U7712 (N_7712,N_4144,N_5155);
and U7713 (N_7713,N_4324,N_4894);
or U7714 (N_7714,N_5140,N_5225);
or U7715 (N_7715,N_4964,N_4671);
nor U7716 (N_7716,N_5613,N_4622);
or U7717 (N_7717,N_4037,N_5518);
nand U7718 (N_7718,N_5543,N_5804);
nand U7719 (N_7719,N_5843,N_5527);
or U7720 (N_7720,N_5867,N_4680);
and U7721 (N_7721,N_4245,N_5000);
nor U7722 (N_7722,N_4189,N_5685);
nand U7723 (N_7723,N_5168,N_5815);
nand U7724 (N_7724,N_5776,N_5867);
nand U7725 (N_7725,N_4727,N_5342);
nor U7726 (N_7726,N_5184,N_5155);
nand U7727 (N_7727,N_5078,N_4118);
or U7728 (N_7728,N_5608,N_5609);
or U7729 (N_7729,N_5623,N_4172);
nor U7730 (N_7730,N_5601,N_5613);
nor U7731 (N_7731,N_4739,N_4850);
and U7732 (N_7732,N_4907,N_4815);
nor U7733 (N_7733,N_5582,N_4810);
or U7734 (N_7734,N_4052,N_4707);
or U7735 (N_7735,N_5797,N_4582);
nor U7736 (N_7736,N_4322,N_5123);
nor U7737 (N_7737,N_4175,N_5833);
nor U7738 (N_7738,N_4269,N_5872);
or U7739 (N_7739,N_4756,N_4436);
nor U7740 (N_7740,N_4393,N_4467);
nor U7741 (N_7741,N_4129,N_5103);
nor U7742 (N_7742,N_4452,N_5426);
or U7743 (N_7743,N_5168,N_5321);
and U7744 (N_7744,N_5713,N_4646);
and U7745 (N_7745,N_4845,N_4549);
nor U7746 (N_7746,N_5223,N_5298);
or U7747 (N_7747,N_4689,N_5218);
nor U7748 (N_7748,N_5278,N_4335);
or U7749 (N_7749,N_4707,N_5852);
and U7750 (N_7750,N_4063,N_4707);
nand U7751 (N_7751,N_5329,N_4192);
nor U7752 (N_7752,N_4913,N_4427);
or U7753 (N_7753,N_5290,N_4787);
and U7754 (N_7754,N_4364,N_4635);
and U7755 (N_7755,N_5702,N_5419);
or U7756 (N_7756,N_5364,N_4468);
nor U7757 (N_7757,N_4138,N_4702);
nand U7758 (N_7758,N_5710,N_5781);
and U7759 (N_7759,N_4064,N_5963);
and U7760 (N_7760,N_4407,N_4853);
nor U7761 (N_7761,N_4813,N_4227);
nand U7762 (N_7762,N_5547,N_4670);
nand U7763 (N_7763,N_5400,N_5498);
nand U7764 (N_7764,N_4808,N_4729);
or U7765 (N_7765,N_5592,N_5330);
nor U7766 (N_7766,N_4191,N_4073);
and U7767 (N_7767,N_4224,N_4312);
and U7768 (N_7768,N_5994,N_4130);
or U7769 (N_7769,N_4852,N_4124);
nor U7770 (N_7770,N_4094,N_5870);
and U7771 (N_7771,N_5824,N_4417);
and U7772 (N_7772,N_5526,N_5511);
nor U7773 (N_7773,N_4456,N_4820);
or U7774 (N_7774,N_4412,N_4808);
and U7775 (N_7775,N_4736,N_4290);
or U7776 (N_7776,N_5957,N_5473);
nor U7777 (N_7777,N_5389,N_5078);
nor U7778 (N_7778,N_5159,N_4759);
or U7779 (N_7779,N_5861,N_5660);
nor U7780 (N_7780,N_4958,N_5172);
and U7781 (N_7781,N_5956,N_5311);
or U7782 (N_7782,N_4474,N_5981);
and U7783 (N_7783,N_5748,N_4925);
nand U7784 (N_7784,N_5143,N_4646);
nand U7785 (N_7785,N_4060,N_4872);
nand U7786 (N_7786,N_5476,N_4553);
nand U7787 (N_7787,N_5958,N_5956);
nand U7788 (N_7788,N_4173,N_4123);
nand U7789 (N_7789,N_4654,N_5426);
nand U7790 (N_7790,N_5760,N_5175);
nor U7791 (N_7791,N_4503,N_5689);
nand U7792 (N_7792,N_4951,N_4529);
nand U7793 (N_7793,N_5965,N_5563);
and U7794 (N_7794,N_5916,N_5246);
and U7795 (N_7795,N_5534,N_4190);
nor U7796 (N_7796,N_4377,N_4799);
or U7797 (N_7797,N_4532,N_5660);
or U7798 (N_7798,N_5678,N_5031);
and U7799 (N_7799,N_4382,N_5451);
nor U7800 (N_7800,N_4905,N_4986);
nor U7801 (N_7801,N_4509,N_5611);
nand U7802 (N_7802,N_5380,N_4603);
nor U7803 (N_7803,N_4163,N_4216);
or U7804 (N_7804,N_4265,N_5016);
or U7805 (N_7805,N_4624,N_5355);
and U7806 (N_7806,N_5107,N_5560);
nor U7807 (N_7807,N_5152,N_5511);
and U7808 (N_7808,N_5160,N_4213);
nand U7809 (N_7809,N_5083,N_5349);
nor U7810 (N_7810,N_4398,N_5439);
xnor U7811 (N_7811,N_5329,N_5018);
or U7812 (N_7812,N_4396,N_4230);
and U7813 (N_7813,N_4127,N_4631);
nand U7814 (N_7814,N_4874,N_5853);
nand U7815 (N_7815,N_5332,N_5983);
nor U7816 (N_7816,N_4562,N_5407);
or U7817 (N_7817,N_5261,N_4976);
nor U7818 (N_7818,N_4422,N_5096);
nor U7819 (N_7819,N_5130,N_5297);
and U7820 (N_7820,N_4006,N_4720);
nand U7821 (N_7821,N_4308,N_5053);
and U7822 (N_7822,N_5117,N_5042);
nor U7823 (N_7823,N_4269,N_4990);
and U7824 (N_7824,N_4416,N_5307);
and U7825 (N_7825,N_5374,N_4188);
and U7826 (N_7826,N_4041,N_5427);
nor U7827 (N_7827,N_4302,N_4188);
and U7828 (N_7828,N_4346,N_4612);
and U7829 (N_7829,N_5763,N_5845);
or U7830 (N_7830,N_4195,N_4791);
nand U7831 (N_7831,N_4096,N_5905);
nor U7832 (N_7832,N_5823,N_5409);
and U7833 (N_7833,N_5593,N_5595);
or U7834 (N_7834,N_4990,N_5950);
or U7835 (N_7835,N_5433,N_4460);
or U7836 (N_7836,N_4082,N_5565);
and U7837 (N_7837,N_5340,N_4877);
and U7838 (N_7838,N_5957,N_5441);
or U7839 (N_7839,N_4283,N_4371);
or U7840 (N_7840,N_5293,N_5640);
nand U7841 (N_7841,N_5788,N_4489);
and U7842 (N_7842,N_4558,N_5231);
or U7843 (N_7843,N_5898,N_5699);
xnor U7844 (N_7844,N_5585,N_5246);
and U7845 (N_7845,N_4433,N_5985);
nor U7846 (N_7846,N_5383,N_5673);
or U7847 (N_7847,N_4692,N_5342);
nand U7848 (N_7848,N_5299,N_4619);
nor U7849 (N_7849,N_4615,N_5773);
and U7850 (N_7850,N_5889,N_4526);
nor U7851 (N_7851,N_4483,N_4892);
or U7852 (N_7852,N_4403,N_4092);
nor U7853 (N_7853,N_5555,N_5922);
nand U7854 (N_7854,N_5005,N_5689);
or U7855 (N_7855,N_4395,N_4138);
nand U7856 (N_7856,N_5220,N_4563);
or U7857 (N_7857,N_4854,N_5224);
nand U7858 (N_7858,N_5301,N_5589);
nand U7859 (N_7859,N_5192,N_4473);
or U7860 (N_7860,N_5972,N_4941);
nand U7861 (N_7861,N_4188,N_5717);
and U7862 (N_7862,N_4360,N_4420);
or U7863 (N_7863,N_4476,N_4840);
and U7864 (N_7864,N_5033,N_5186);
and U7865 (N_7865,N_5252,N_4619);
or U7866 (N_7866,N_4377,N_5006);
or U7867 (N_7867,N_4341,N_5626);
and U7868 (N_7868,N_5003,N_4020);
or U7869 (N_7869,N_5619,N_4737);
nor U7870 (N_7870,N_5120,N_4291);
or U7871 (N_7871,N_4958,N_4636);
and U7872 (N_7872,N_4656,N_5133);
and U7873 (N_7873,N_4337,N_4400);
nor U7874 (N_7874,N_5842,N_5144);
and U7875 (N_7875,N_4927,N_5748);
nand U7876 (N_7876,N_5240,N_5067);
nand U7877 (N_7877,N_4995,N_4180);
or U7878 (N_7878,N_5122,N_4805);
nand U7879 (N_7879,N_4434,N_4455);
and U7880 (N_7880,N_4605,N_4335);
or U7881 (N_7881,N_5258,N_4590);
nor U7882 (N_7882,N_5200,N_5551);
or U7883 (N_7883,N_4502,N_5134);
or U7884 (N_7884,N_5384,N_5615);
nand U7885 (N_7885,N_4898,N_4048);
and U7886 (N_7886,N_5748,N_5647);
nand U7887 (N_7887,N_4099,N_5872);
nor U7888 (N_7888,N_5918,N_4439);
nor U7889 (N_7889,N_5463,N_4769);
nand U7890 (N_7890,N_5432,N_4521);
or U7891 (N_7891,N_4622,N_5175);
nor U7892 (N_7892,N_5102,N_4309);
and U7893 (N_7893,N_4098,N_4007);
or U7894 (N_7894,N_5412,N_4211);
or U7895 (N_7895,N_4314,N_5981);
and U7896 (N_7896,N_4415,N_5357);
nand U7897 (N_7897,N_5686,N_5094);
and U7898 (N_7898,N_4540,N_4479);
nor U7899 (N_7899,N_5009,N_5761);
nor U7900 (N_7900,N_5499,N_5595);
nand U7901 (N_7901,N_5713,N_5551);
nand U7902 (N_7902,N_5668,N_4824);
nand U7903 (N_7903,N_4221,N_4306);
nand U7904 (N_7904,N_4417,N_5515);
nand U7905 (N_7905,N_5741,N_4485);
and U7906 (N_7906,N_4050,N_5701);
and U7907 (N_7907,N_4312,N_4013);
and U7908 (N_7908,N_4062,N_5702);
or U7909 (N_7909,N_4716,N_5880);
nor U7910 (N_7910,N_4021,N_5167);
and U7911 (N_7911,N_4818,N_4807);
nand U7912 (N_7912,N_5912,N_5231);
or U7913 (N_7913,N_4121,N_5277);
and U7914 (N_7914,N_5369,N_5346);
and U7915 (N_7915,N_4785,N_5523);
nor U7916 (N_7916,N_5503,N_4609);
and U7917 (N_7917,N_4198,N_5737);
or U7918 (N_7918,N_5719,N_5010);
or U7919 (N_7919,N_4532,N_5292);
or U7920 (N_7920,N_5542,N_4464);
and U7921 (N_7921,N_5766,N_4995);
nor U7922 (N_7922,N_4633,N_4739);
or U7923 (N_7923,N_4728,N_5245);
and U7924 (N_7924,N_5832,N_4903);
or U7925 (N_7925,N_4791,N_5014);
nand U7926 (N_7926,N_4641,N_4661);
or U7927 (N_7927,N_5688,N_4591);
nand U7928 (N_7928,N_5308,N_5432);
nor U7929 (N_7929,N_4759,N_4293);
and U7930 (N_7930,N_5541,N_4393);
or U7931 (N_7931,N_5878,N_4997);
nand U7932 (N_7932,N_4885,N_4612);
nand U7933 (N_7933,N_5509,N_5252);
and U7934 (N_7934,N_5410,N_5633);
nand U7935 (N_7935,N_4709,N_4316);
xor U7936 (N_7936,N_5445,N_4831);
or U7937 (N_7937,N_5889,N_5580);
or U7938 (N_7938,N_4861,N_5388);
nand U7939 (N_7939,N_4137,N_4074);
and U7940 (N_7940,N_5280,N_4812);
and U7941 (N_7941,N_4717,N_4358);
xor U7942 (N_7942,N_5410,N_4760);
or U7943 (N_7943,N_4734,N_5701);
and U7944 (N_7944,N_4375,N_5805);
xnor U7945 (N_7945,N_5773,N_4826);
nand U7946 (N_7946,N_4992,N_5197);
nor U7947 (N_7947,N_4822,N_5473);
and U7948 (N_7948,N_4175,N_4672);
nor U7949 (N_7949,N_5350,N_5324);
nand U7950 (N_7950,N_5221,N_5262);
or U7951 (N_7951,N_4840,N_4680);
or U7952 (N_7952,N_4708,N_4432);
nand U7953 (N_7953,N_4492,N_4234);
or U7954 (N_7954,N_4248,N_5376);
nand U7955 (N_7955,N_4247,N_4466);
nand U7956 (N_7956,N_4296,N_4512);
and U7957 (N_7957,N_5253,N_4615);
or U7958 (N_7958,N_5209,N_5190);
nor U7959 (N_7959,N_4023,N_4848);
nand U7960 (N_7960,N_5974,N_5699);
xor U7961 (N_7961,N_5925,N_4633);
nand U7962 (N_7962,N_5015,N_5335);
nand U7963 (N_7963,N_4131,N_4423);
or U7964 (N_7964,N_5872,N_4104);
nand U7965 (N_7965,N_5149,N_4225);
or U7966 (N_7966,N_4314,N_5310);
or U7967 (N_7967,N_4778,N_5375);
nor U7968 (N_7968,N_4711,N_5910);
nor U7969 (N_7969,N_5851,N_4427);
nand U7970 (N_7970,N_4667,N_4509);
nor U7971 (N_7971,N_5611,N_5789);
nand U7972 (N_7972,N_4799,N_4393);
nand U7973 (N_7973,N_4567,N_5077);
and U7974 (N_7974,N_4651,N_4624);
and U7975 (N_7975,N_4096,N_4806);
or U7976 (N_7976,N_5295,N_5269);
and U7977 (N_7977,N_5023,N_5431);
or U7978 (N_7978,N_4719,N_4618);
or U7979 (N_7979,N_4883,N_4123);
nor U7980 (N_7980,N_5026,N_4487);
and U7981 (N_7981,N_5772,N_5009);
nand U7982 (N_7982,N_5679,N_5035);
and U7983 (N_7983,N_5570,N_4387);
or U7984 (N_7984,N_5080,N_4519);
and U7985 (N_7985,N_5296,N_4725);
or U7986 (N_7986,N_5808,N_4992);
nand U7987 (N_7987,N_4776,N_4627);
or U7988 (N_7988,N_4408,N_4137);
nor U7989 (N_7989,N_4155,N_5395);
nor U7990 (N_7990,N_4645,N_5346);
or U7991 (N_7991,N_4425,N_4086);
or U7992 (N_7992,N_5581,N_4200);
or U7993 (N_7993,N_5978,N_5582);
nor U7994 (N_7994,N_4689,N_4872);
or U7995 (N_7995,N_4240,N_5839);
and U7996 (N_7996,N_5996,N_5448);
nand U7997 (N_7997,N_4997,N_4487);
nor U7998 (N_7998,N_4867,N_5724);
nor U7999 (N_7999,N_4388,N_5815);
nor U8000 (N_8000,N_7669,N_7215);
and U8001 (N_8001,N_6211,N_6556);
nor U8002 (N_8002,N_6438,N_7498);
or U8003 (N_8003,N_6667,N_6068);
or U8004 (N_8004,N_6006,N_6803);
or U8005 (N_8005,N_7516,N_7470);
nor U8006 (N_8006,N_7693,N_7964);
nand U8007 (N_8007,N_6084,N_7011);
nand U8008 (N_8008,N_7762,N_7068);
nand U8009 (N_8009,N_6315,N_7243);
nand U8010 (N_8010,N_7449,N_6625);
and U8011 (N_8011,N_6745,N_7835);
nor U8012 (N_8012,N_7763,N_7357);
nand U8013 (N_8013,N_6053,N_6437);
nor U8014 (N_8014,N_6340,N_6615);
nand U8015 (N_8015,N_7335,N_6020);
and U8016 (N_8016,N_7887,N_7624);
and U8017 (N_8017,N_7833,N_7950);
or U8018 (N_8018,N_6689,N_7953);
and U8019 (N_8019,N_6930,N_6806);
nor U8020 (N_8020,N_7792,N_6546);
or U8021 (N_8021,N_7663,N_6077);
and U8022 (N_8022,N_7928,N_7736);
and U8023 (N_8023,N_7188,N_6558);
and U8024 (N_8024,N_7692,N_6732);
nor U8025 (N_8025,N_7151,N_6705);
nor U8026 (N_8026,N_7428,N_7227);
nand U8027 (N_8027,N_7001,N_7466);
or U8028 (N_8028,N_7678,N_6280);
nor U8029 (N_8029,N_6092,N_7668);
nand U8030 (N_8030,N_7542,N_6367);
nand U8031 (N_8031,N_6061,N_6722);
or U8032 (N_8032,N_6790,N_7787);
nand U8033 (N_8033,N_6958,N_7019);
nor U8034 (N_8034,N_7353,N_6633);
nor U8035 (N_8035,N_7195,N_7976);
and U8036 (N_8036,N_7558,N_6002);
or U8037 (N_8037,N_7281,N_6814);
and U8038 (N_8038,N_6196,N_7012);
and U8039 (N_8039,N_6690,N_6605);
nor U8040 (N_8040,N_7643,N_6992);
nor U8041 (N_8041,N_6099,N_6226);
and U8042 (N_8042,N_7153,N_7440);
and U8043 (N_8043,N_6236,N_7530);
and U8044 (N_8044,N_6279,N_7280);
and U8045 (N_8045,N_6425,N_7237);
nand U8046 (N_8046,N_6496,N_7163);
and U8047 (N_8047,N_6976,N_6116);
nand U8048 (N_8048,N_6140,N_7711);
nor U8049 (N_8049,N_7483,N_7347);
and U8050 (N_8050,N_6013,N_7911);
and U8051 (N_8051,N_7297,N_7829);
nor U8052 (N_8052,N_6662,N_7596);
and U8053 (N_8053,N_6602,N_6240);
nand U8054 (N_8054,N_6168,N_7584);
nor U8055 (N_8055,N_6833,N_7020);
and U8056 (N_8056,N_7408,N_7332);
nand U8057 (N_8057,N_6523,N_7699);
nand U8058 (N_8058,N_7644,N_7646);
nand U8059 (N_8059,N_7202,N_7629);
nor U8060 (N_8060,N_7476,N_6947);
or U8061 (N_8061,N_6305,N_6697);
nand U8062 (N_8062,N_6350,N_7654);
nor U8063 (N_8063,N_6940,N_6986);
nand U8064 (N_8064,N_7688,N_7588);
nand U8065 (N_8065,N_6977,N_7058);
nand U8066 (N_8066,N_7574,N_6054);
and U8067 (N_8067,N_7377,N_7304);
nor U8068 (N_8068,N_6498,N_7446);
xnor U8069 (N_8069,N_7217,N_6097);
or U8070 (N_8070,N_6862,N_7619);
or U8071 (N_8071,N_7898,N_7568);
and U8072 (N_8072,N_7289,N_6552);
nor U8073 (N_8073,N_7945,N_6674);
and U8074 (N_8074,N_7790,N_6098);
nand U8075 (N_8075,N_6287,N_6318);
or U8076 (N_8076,N_7176,N_7991);
and U8077 (N_8077,N_6677,N_6235);
and U8078 (N_8078,N_7370,N_7576);
and U8079 (N_8079,N_7747,N_6812);
nand U8080 (N_8080,N_7034,N_6826);
nand U8081 (N_8081,N_7623,N_7321);
and U8082 (N_8082,N_7415,N_6572);
and U8083 (N_8083,N_7456,N_7102);
or U8084 (N_8084,N_7830,N_7900);
nor U8085 (N_8085,N_7444,N_6752);
and U8086 (N_8086,N_7719,N_6816);
and U8087 (N_8087,N_7645,N_7988);
nand U8088 (N_8088,N_7252,N_7837);
and U8089 (N_8089,N_6829,N_7635);
nand U8090 (N_8090,N_7059,N_7655);
nand U8091 (N_8091,N_7512,N_6292);
and U8092 (N_8092,N_6458,N_6301);
or U8093 (N_8093,N_7130,N_6758);
or U8094 (N_8094,N_6881,N_7256);
or U8095 (N_8095,N_7480,N_7072);
and U8096 (N_8096,N_7735,N_7422);
and U8097 (N_8097,N_6048,N_7264);
nand U8098 (N_8098,N_6778,N_6701);
nor U8099 (N_8099,N_7031,N_6673);
nor U8100 (N_8100,N_7875,N_6743);
nand U8101 (N_8101,N_6581,N_6709);
or U8102 (N_8102,N_6921,N_6578);
xnor U8103 (N_8103,N_7608,N_7326);
nand U8104 (N_8104,N_6138,N_6510);
and U8105 (N_8105,N_6208,N_6057);
nor U8106 (N_8106,N_6165,N_7520);
or U8107 (N_8107,N_6285,N_7862);
nor U8108 (N_8108,N_6639,N_7865);
nand U8109 (N_8109,N_7184,N_7778);
nor U8110 (N_8110,N_6272,N_6832);
nor U8111 (N_8111,N_6353,N_7818);
and U8112 (N_8112,N_7975,N_6514);
nor U8113 (N_8113,N_7404,N_6435);
or U8114 (N_8114,N_6991,N_6485);
or U8115 (N_8115,N_6500,N_6649);
or U8116 (N_8116,N_7302,N_7433);
and U8117 (N_8117,N_7394,N_7391);
and U8118 (N_8118,N_7864,N_6617);
nand U8119 (N_8119,N_6336,N_6129);
nand U8120 (N_8120,N_7538,N_6174);
and U8121 (N_8121,N_6933,N_6804);
nand U8122 (N_8122,N_7544,N_6374);
nor U8123 (N_8123,N_7101,N_7495);
nor U8124 (N_8124,N_7567,N_7078);
or U8125 (N_8125,N_6936,N_6085);
nor U8126 (N_8126,N_6968,N_6499);
nand U8127 (N_8127,N_7192,N_6532);
nor U8128 (N_8128,N_7152,N_7856);
and U8129 (N_8129,N_6357,N_6014);
nand U8130 (N_8130,N_7791,N_7665);
and U8131 (N_8131,N_6724,N_7522);
and U8132 (N_8132,N_7859,N_6571);
nor U8133 (N_8133,N_7807,N_7994);
nand U8134 (N_8134,N_6952,N_7049);
or U8135 (N_8135,N_6463,N_7009);
nand U8136 (N_8136,N_6531,N_7587);
and U8137 (N_8137,N_6700,N_6985);
nand U8138 (N_8138,N_7380,N_6560);
and U8139 (N_8139,N_6345,N_7876);
nand U8140 (N_8140,N_7231,N_7943);
nor U8141 (N_8141,N_7491,N_6419);
nand U8142 (N_8142,N_7014,N_6923);
and U8143 (N_8143,N_7293,N_7944);
or U8144 (N_8144,N_6799,N_6711);
nor U8145 (N_8145,N_6997,N_6128);
nand U8146 (N_8146,N_7016,N_6426);
nand U8147 (N_8147,N_7201,N_6965);
and U8148 (N_8148,N_7882,N_7395);
or U8149 (N_8149,N_7499,N_7779);
nor U8150 (N_8150,N_6082,N_6993);
nand U8151 (N_8151,N_7378,N_6164);
or U8152 (N_8152,N_6884,N_6950);
nand U8153 (N_8153,N_7632,N_7717);
or U8154 (N_8154,N_6781,N_6202);
nand U8155 (N_8155,N_7165,N_7131);
or U8156 (N_8156,N_7559,N_7207);
nand U8157 (N_8157,N_7331,N_6948);
nor U8158 (N_8158,N_6584,N_7513);
or U8159 (N_8159,N_7927,N_7956);
nand U8160 (N_8160,N_7193,N_6576);
nand U8161 (N_8161,N_7505,N_6033);
nor U8162 (N_8162,N_6026,N_7222);
nor U8163 (N_8163,N_6623,N_6171);
or U8164 (N_8164,N_7006,N_6370);
or U8165 (N_8165,N_7661,N_6938);
nand U8166 (N_8166,N_6907,N_7569);
or U8167 (N_8167,N_6794,N_6113);
and U8168 (N_8168,N_6186,N_7066);
nand U8169 (N_8169,N_7734,N_7575);
or U8170 (N_8170,N_7253,N_7714);
nor U8171 (N_8171,N_7981,N_7371);
nand U8172 (N_8172,N_6870,N_7926);
nor U8173 (N_8173,N_7345,N_7314);
or U8174 (N_8174,N_6218,N_6133);
nand U8175 (N_8175,N_7294,N_7147);
and U8176 (N_8176,N_7720,N_6636);
and U8177 (N_8177,N_6646,N_6851);
and U8178 (N_8178,N_7552,N_6586);
nand U8179 (N_8179,N_7684,N_6343);
and U8180 (N_8180,N_7658,N_7946);
or U8181 (N_8181,N_6900,N_7182);
and U8182 (N_8182,N_7851,N_6232);
nor U8183 (N_8183,N_6720,N_7700);
nand U8184 (N_8184,N_6362,N_6856);
and U8185 (N_8185,N_6414,N_6598);
nor U8186 (N_8186,N_6502,N_6474);
nand U8187 (N_8187,N_7033,N_6431);
and U8188 (N_8188,N_7809,N_7703);
and U8189 (N_8189,N_7724,N_6775);
nor U8190 (N_8190,N_7250,N_6018);
nor U8191 (N_8191,N_7485,N_6738);
or U8192 (N_8192,N_7075,N_6595);
nor U8193 (N_8193,N_7113,N_7770);
nand U8194 (N_8194,N_7268,N_6820);
and U8195 (N_8195,N_6980,N_7450);
nor U8196 (N_8196,N_6213,N_7750);
xnor U8197 (N_8197,N_7417,N_7783);
nand U8198 (N_8198,N_7627,N_6616);
or U8199 (N_8199,N_6535,N_7581);
and U8200 (N_8200,N_7838,N_7155);
and U8201 (N_8201,N_7274,N_7196);
or U8202 (N_8202,N_7883,N_6102);
or U8203 (N_8203,N_7804,N_6131);
or U8204 (N_8204,N_7122,N_6878);
xor U8205 (N_8205,N_7521,N_7021);
or U8206 (N_8206,N_6508,N_6984);
or U8207 (N_8207,N_7285,N_6916);
or U8208 (N_8208,N_7174,N_7402);
or U8209 (N_8209,N_7346,N_6317);
nor U8210 (N_8210,N_6767,N_6073);
or U8211 (N_8211,N_6436,N_6117);
nor U8212 (N_8212,N_7503,N_7959);
nand U8213 (N_8213,N_6166,N_7537);
nand U8214 (N_8214,N_7482,N_6328);
or U8215 (N_8215,N_6488,N_6342);
nor U8216 (N_8216,N_6134,N_7247);
or U8217 (N_8217,N_7630,N_7112);
nand U8218 (N_8218,N_7897,N_7571);
nor U8219 (N_8219,N_6730,N_7808);
or U8220 (N_8220,N_6522,N_7842);
nand U8221 (N_8221,N_6119,N_6069);
and U8222 (N_8222,N_6599,N_6162);
and U8223 (N_8223,N_6086,N_7159);
nor U8224 (N_8224,N_6135,N_7213);
nor U8225 (N_8225,N_6258,N_6442);
nor U8226 (N_8226,N_6658,N_6528);
and U8227 (N_8227,N_7802,N_6902);
or U8228 (N_8228,N_6155,N_7874);
nor U8229 (N_8229,N_6214,N_7403);
or U8230 (N_8230,N_7270,N_7935);
nor U8231 (N_8231,N_6477,N_6380);
or U8232 (N_8232,N_7651,N_6101);
nand U8233 (N_8233,N_6717,N_7759);
nand U8234 (N_8234,N_7497,N_6580);
nand U8235 (N_8235,N_6934,N_6681);
or U8236 (N_8236,N_7190,N_7288);
nor U8237 (N_8237,N_6480,N_7179);
nor U8238 (N_8238,N_7570,N_7419);
nor U8239 (N_8239,N_6052,N_6517);
nand U8240 (N_8240,N_6899,N_6610);
and U8241 (N_8241,N_6282,N_6243);
or U8242 (N_8242,N_7824,N_6269);
nor U8243 (N_8243,N_7170,N_7834);
and U8244 (N_8244,N_7532,N_7080);
or U8245 (N_8245,N_7226,N_6579);
and U8246 (N_8246,N_7311,N_7696);
nand U8247 (N_8247,N_7600,N_7459);
and U8248 (N_8248,N_7464,N_6863);
nand U8249 (N_8249,N_6566,N_7869);
nand U8250 (N_8250,N_6462,N_7189);
and U8251 (N_8251,N_6904,N_6653);
nand U8252 (N_8252,N_7010,N_6180);
and U8253 (N_8253,N_6783,N_6755);
or U8254 (N_8254,N_6320,N_6453);
and U8255 (N_8255,N_6634,N_7847);
nand U8256 (N_8256,N_7076,N_7309);
or U8257 (N_8257,N_6945,N_7985);
and U8258 (N_8258,N_6307,N_7952);
nand U8259 (N_8259,N_6312,N_7702);
nor U8260 (N_8260,N_7392,N_6493);
and U8261 (N_8261,N_7091,N_6565);
or U8262 (N_8262,N_7306,N_6434);
nand U8263 (N_8263,N_6604,N_7566);
nor U8264 (N_8264,N_6967,N_6005);
nand U8265 (N_8265,N_6352,N_7723);
or U8266 (N_8266,N_6858,N_6927);
and U8267 (N_8267,N_7768,N_6664);
and U8268 (N_8268,N_7164,N_6702);
xor U8269 (N_8269,N_6205,N_6773);
or U8270 (N_8270,N_6928,N_6685);
nor U8271 (N_8271,N_7634,N_7168);
nand U8272 (N_8272,N_6257,N_7715);
or U8273 (N_8273,N_6228,N_7881);
nor U8274 (N_8274,N_7109,N_6311);
nand U8275 (N_8275,N_6375,N_7000);
nand U8276 (N_8276,N_7385,N_6201);
nand U8277 (N_8277,N_7732,N_6547);
and U8278 (N_8278,N_7259,N_7100);
and U8279 (N_8279,N_6156,N_6942);
nor U8280 (N_8280,N_7508,N_6088);
nor U8281 (N_8281,N_6562,N_7934);
nor U8282 (N_8282,N_7528,N_7209);
and U8283 (N_8283,N_7526,N_6430);
nand U8284 (N_8284,N_7695,N_6137);
nand U8285 (N_8285,N_7424,N_6151);
and U8286 (N_8286,N_6944,N_6268);
nand U8287 (N_8287,N_7782,N_7867);
nor U8288 (N_8288,N_7690,N_7580);
nand U8289 (N_8289,N_6420,N_7286);
nand U8290 (N_8290,N_6748,N_7187);
nor U8291 (N_8291,N_7341,N_7515);
nand U8292 (N_8292,N_7919,N_6076);
or U8293 (N_8293,N_7373,N_7043);
or U8294 (N_8294,N_7437,N_7666);
or U8295 (N_8295,N_6897,N_7050);
or U8296 (N_8296,N_6583,N_6801);
nor U8297 (N_8297,N_6678,N_7206);
and U8298 (N_8298,N_6010,N_6630);
nor U8299 (N_8299,N_6793,N_6682);
and U8300 (N_8300,N_7815,N_7997);
and U8301 (N_8301,N_6160,N_7716);
nand U8302 (N_8302,N_6015,N_7452);
nand U8303 (N_8303,N_6219,N_7936);
or U8304 (N_8304,N_6237,N_7148);
nor U8305 (N_8305,N_6982,N_6472);
nand U8306 (N_8306,N_6712,N_7477);
nor U8307 (N_8307,N_7040,N_6706);
nor U8308 (N_8308,N_7023,N_7729);
or U8309 (N_8309,N_6473,N_6210);
nand U8310 (N_8310,N_7605,N_6998);
and U8311 (N_8311,N_6729,N_6670);
nand U8312 (N_8312,N_7725,N_7914);
and U8313 (N_8313,N_7129,N_7501);
nor U8314 (N_8314,N_7032,N_7968);
or U8315 (N_8315,N_6512,N_6199);
or U8316 (N_8316,N_7622,N_6641);
or U8317 (N_8317,N_7510,N_7523);
and U8318 (N_8318,N_6910,N_6759);
nand U8319 (N_8319,N_7305,N_7942);
nor U8320 (N_8320,N_7890,N_6715);
nand U8321 (N_8321,N_7748,N_6760);
nand U8322 (N_8322,N_6153,N_7626);
and U8323 (N_8323,N_6632,N_6684);
nor U8324 (N_8324,N_6874,N_6503);
and U8325 (N_8325,N_6590,N_6635);
nor U8326 (N_8326,N_6003,N_6660);
nor U8327 (N_8327,N_7839,N_7296);
and U8328 (N_8328,N_6486,N_6421);
and U8329 (N_8329,N_7916,N_7099);
nand U8330 (N_8330,N_6567,N_6323);
or U8331 (N_8331,N_6959,N_7236);
nand U8332 (N_8332,N_6847,N_7721);
and U8333 (N_8333,N_6446,N_7784);
nand U8334 (N_8334,N_6726,N_7234);
nand U8335 (N_8335,N_6857,N_6839);
or U8336 (N_8336,N_7531,N_7899);
nor U8337 (N_8337,N_7962,N_6246);
and U8338 (N_8338,N_6450,N_7949);
nor U8339 (N_8339,N_6106,N_7667);
or U8340 (N_8340,N_7088,N_6441);
and U8341 (N_8341,N_7733,N_7816);
or U8342 (N_8342,N_7990,N_7396);
or U8343 (N_8343,N_7045,N_7984);
and U8344 (N_8344,N_7755,N_6638);
and U8345 (N_8345,N_7261,N_6284);
xnor U8346 (N_8346,N_7710,N_7880);
and U8347 (N_8347,N_7481,N_6957);
or U8348 (N_8348,N_6785,N_6611);
or U8349 (N_8349,N_6009,N_6538);
or U8350 (N_8350,N_6796,N_6169);
or U8351 (N_8351,N_7134,N_7740);
nand U8352 (N_8352,N_6850,N_7514);
nand U8353 (N_8353,N_6407,N_7966);
or U8354 (N_8354,N_7673,N_7359);
nand U8355 (N_8355,N_6574,N_6526);
or U8356 (N_8356,N_7056,N_7208);
and U8357 (N_8357,N_6844,N_6159);
nor U8358 (N_8358,N_6853,N_7469);
nand U8359 (N_8359,N_7300,N_6206);
nor U8360 (N_8360,N_7017,N_7219);
nor U8361 (N_8361,N_7682,N_7376);
nand U8362 (N_8362,N_6242,N_7519);
nor U8363 (N_8363,N_7382,N_6283);
nand U8364 (N_8364,N_6613,N_7850);
or U8365 (N_8365,N_7775,N_6838);
nand U8366 (N_8366,N_6824,N_6779);
or U8367 (N_8367,N_7255,N_7597);
or U8368 (N_8368,N_6805,N_6379);
nor U8369 (N_8369,N_6163,N_7751);
and U8370 (N_8370,N_6791,N_7960);
and U8371 (N_8371,N_7915,N_6046);
or U8372 (N_8372,N_7582,N_7212);
nor U8373 (N_8373,N_7015,N_6813);
nor U8374 (N_8374,N_7741,N_6591);
and U8375 (N_8375,N_6672,N_6527);
and U8376 (N_8376,N_6022,N_7381);
or U8377 (N_8377,N_7772,N_6596);
and U8378 (N_8378,N_7454,N_7194);
or U8379 (N_8379,N_7912,N_7098);
nor U8380 (N_8380,N_6593,N_6931);
nand U8381 (N_8381,N_6883,N_6244);
nand U8382 (N_8382,N_6797,N_6439);
nor U8383 (N_8383,N_7676,N_6573);
nor U8384 (N_8384,N_6247,N_7356);
nand U8385 (N_8385,N_6735,N_7607);
or U8386 (N_8386,N_6021,N_6569);
xor U8387 (N_8387,N_7731,N_6540);
nand U8388 (N_8388,N_7979,N_6229);
or U8389 (N_8389,N_6469,N_7551);
nor U8390 (N_8390,N_7149,N_6886);
nand U8391 (N_8391,N_7290,N_6424);
and U8392 (N_8392,N_7598,N_7205);
or U8393 (N_8393,N_6536,N_6185);
and U8394 (N_8394,N_7420,N_7572);
or U8395 (N_8395,N_7757,N_7465);
nor U8396 (N_8396,N_7200,N_6932);
nor U8397 (N_8397,N_7046,N_6975);
nand U8398 (N_8398,N_6124,N_6582);
or U8399 (N_8399,N_7117,N_6676);
and U8400 (N_8400,N_6918,N_6905);
or U8401 (N_8401,N_7048,N_7955);
and U8402 (N_8402,N_7279,N_6036);
and U8403 (N_8403,N_7333,N_7167);
or U8404 (N_8404,N_7978,N_7365);
nor U8405 (N_8405,N_7664,N_7947);
and U8406 (N_8406,N_6753,N_6093);
or U8407 (N_8407,N_6108,N_7819);
or U8408 (N_8408,N_7920,N_6062);
or U8409 (N_8409,N_7399,N_6941);
nor U8410 (N_8410,N_7108,N_7754);
or U8411 (N_8411,N_6999,N_6189);
and U8412 (N_8412,N_6704,N_7892);
nand U8413 (N_8413,N_7848,N_7478);
and U8414 (N_8414,N_6207,N_6460);
and U8415 (N_8415,N_6501,N_6482);
or U8416 (N_8416,N_7776,N_7178);
nor U8417 (N_8417,N_6392,N_6867);
and U8418 (N_8418,N_6683,N_7507);
nand U8419 (N_8419,N_7825,N_6860);
and U8420 (N_8420,N_6456,N_7933);
nor U8421 (N_8421,N_7362,N_6875);
and U8422 (N_8422,N_7271,N_6644);
or U8423 (N_8423,N_6648,N_6490);
and U8424 (N_8424,N_6074,N_7752);
and U8425 (N_8425,N_7931,N_6358);
nor U8426 (N_8426,N_6901,N_6507);
and U8427 (N_8427,N_7908,N_7562);
nor U8428 (N_8428,N_7832,N_7372);
and U8429 (N_8429,N_6551,N_7743);
nand U8430 (N_8430,N_6626,N_7447);
nor U8431 (N_8431,N_7327,N_6215);
nor U8432 (N_8432,N_7322,N_7092);
or U8433 (N_8433,N_6585,N_7342);
and U8434 (N_8434,N_7410,N_6198);
and U8435 (N_8435,N_7369,N_6448);
or U8436 (N_8436,N_6943,N_7060);
nand U8437 (N_8437,N_7873,N_6390);
or U8438 (N_8438,N_6680,N_7427);
nor U8439 (N_8439,N_6751,N_7007);
nand U8440 (N_8440,N_7987,N_7283);
or U8441 (N_8441,N_6286,N_6233);
nor U8442 (N_8442,N_6079,N_7885);
or U8443 (N_8443,N_6817,N_7840);
and U8444 (N_8444,N_7426,N_7612);
nor U8445 (N_8445,N_7907,N_6276);
and U8446 (N_8446,N_7652,N_7301);
and U8447 (N_8447,N_7786,N_7257);
and U8448 (N_8448,N_7339,N_7284);
nand U8449 (N_8449,N_6515,N_7282);
nor U8450 (N_8450,N_7706,N_7554);
nor U8451 (N_8451,N_6687,N_6483);
nand U8452 (N_8452,N_6854,N_6273);
or U8453 (N_8453,N_6831,N_6209);
nor U8454 (N_8454,N_6728,N_7039);
xnor U8455 (N_8455,N_6764,N_6607);
and U8456 (N_8456,N_7854,N_7533);
nor U8457 (N_8457,N_7621,N_7421);
nor U8458 (N_8458,N_7871,N_6810);
nor U8459 (N_8459,N_6840,N_6158);
and U8460 (N_8460,N_6447,N_6798);
nor U8461 (N_8461,N_6110,N_7648);
nand U8462 (N_8462,N_6471,N_6827);
nor U8463 (N_8463,N_7350,N_7064);
nor U8464 (N_8464,N_6339,N_6777);
nor U8465 (N_8465,N_7360,N_6511);
or U8466 (N_8466,N_6399,N_7313);
nand U8467 (N_8467,N_7161,N_6385);
nand U8468 (N_8468,N_6908,N_6714);
nand U8469 (N_8469,N_6418,N_6600);
or U8470 (N_8470,N_7577,N_6039);
nand U8471 (N_8471,N_7386,N_7096);
or U8472 (N_8472,N_7044,N_7689);
nand U8473 (N_8473,N_6698,N_6909);
or U8474 (N_8474,N_6139,N_7930);
or U8475 (N_8475,N_7351,N_6624);
or U8476 (N_8476,N_7005,N_7620);
nand U8477 (N_8477,N_7018,N_6464);
nand U8478 (N_8478,N_6346,N_6828);
or U8479 (N_8479,N_7269,N_6559);
or U8480 (N_8480,N_6167,N_7789);
nand U8481 (N_8481,N_7980,N_6087);
or U8482 (N_8482,N_6382,N_6443);
nand U8483 (N_8483,N_6761,N_6809);
or U8484 (N_8484,N_7698,N_7047);
or U8485 (N_8485,N_7003,N_6327);
nand U8486 (N_8486,N_6622,N_6182);
nand U8487 (N_8487,N_7249,N_6043);
nor U8488 (N_8488,N_6757,N_7860);
or U8489 (N_8489,N_6719,N_6296);
nand U8490 (N_8490,N_7974,N_7594);
nor U8491 (N_8491,N_6309,N_6360);
and U8492 (N_8492,N_7954,N_7375);
nand U8493 (N_8493,N_6710,N_7487);
nor U8494 (N_8494,N_7709,N_6772);
nand U8495 (N_8495,N_6412,N_6262);
xnor U8496 (N_8496,N_7463,N_6506);
nor U8497 (N_8497,N_7467,N_6529);
nand U8498 (N_8498,N_6118,N_6321);
or U8499 (N_8499,N_6238,N_7561);
and U8500 (N_8500,N_6946,N_7389);
or U8501 (N_8501,N_7133,N_6518);
and U8502 (N_8502,N_7251,N_6386);
nor U8503 (N_8503,N_7413,N_6603);
nand U8504 (N_8504,N_7121,N_6223);
nand U8505 (N_8505,N_6692,N_6568);
nand U8506 (N_8506,N_6197,N_6361);
and U8507 (N_8507,N_6173,N_6376);
and U8508 (N_8508,N_7822,N_7136);
or U8509 (N_8509,N_6668,N_6152);
nand U8510 (N_8510,N_7035,N_6645);
nor U8511 (N_8511,N_6554,N_6049);
and U8512 (N_8512,N_7811,N_6628);
or U8513 (N_8513,N_7453,N_7795);
nand U8514 (N_8514,N_6396,N_7343);
nor U8515 (N_8515,N_6981,N_6221);
or U8516 (N_8516,N_6121,N_6070);
or U8517 (N_8517,N_6170,N_7303);
and U8518 (N_8518,N_6267,N_6509);
and U8519 (N_8519,N_6191,N_7647);
and U8520 (N_8520,N_6024,N_7901);
and U8521 (N_8521,N_6837,N_7084);
nand U8522 (N_8522,N_6372,N_7705);
nand U8523 (N_8523,N_6561,N_7265);
nor U8524 (N_8524,N_6811,N_7166);
nand U8525 (N_8525,N_6393,N_6754);
nor U8526 (N_8526,N_7863,N_7337);
and U8527 (N_8527,N_6125,N_6356);
or U8528 (N_8528,N_6782,N_7810);
or U8529 (N_8529,N_7330,N_6808);
nor U8530 (N_8530,N_6181,N_6864);
and U8531 (N_8531,N_6721,N_6184);
or U8532 (N_8532,N_7083,N_7320);
and U8533 (N_8533,N_7145,N_6041);
and U8534 (N_8534,N_6802,N_6051);
nor U8535 (N_8535,N_6996,N_7686);
or U8536 (N_8536,N_7640,N_7140);
or U8537 (N_8537,N_7971,N_7504);
nor U8538 (N_8538,N_6731,N_7650);
nand U8539 (N_8539,N_7764,N_6872);
nand U8540 (N_8540,N_6222,N_7794);
nand U8541 (N_8541,N_6027,N_6744);
or U8542 (N_8542,N_6818,N_7107);
and U8543 (N_8543,N_6612,N_7126);
and U8544 (N_8544,N_6225,N_6890);
or U8545 (N_8545,N_6072,N_7799);
nor U8546 (N_8546,N_6019,N_6187);
and U8547 (N_8547,N_7115,N_7679);
or U8548 (N_8548,N_6478,N_6330);
and U8549 (N_8549,N_7739,N_7742);
nor U8550 (N_8550,N_7114,N_6953);
nor U8551 (N_8551,N_6115,N_7841);
or U8552 (N_8552,N_7336,N_7323);
nand U8553 (N_8553,N_7146,N_7073);
or U8554 (N_8554,N_6987,N_7820);
or U8555 (N_8555,N_7423,N_7937);
nand U8556 (N_8556,N_6629,N_7722);
nand U8557 (N_8557,N_6815,N_6428);
nand U8558 (N_8558,N_7004,N_6949);
and U8559 (N_8559,N_6251,N_6520);
or U8560 (N_8560,N_7905,N_6849);
and U8561 (N_8561,N_7616,N_6275);
and U8562 (N_8562,N_6234,N_7613);
nor U8563 (N_8563,N_6564,N_6368);
nor U8564 (N_8564,N_6132,N_7104);
nand U8565 (N_8565,N_6652,N_6302);
and U8566 (N_8566,N_6440,N_6391);
or U8567 (N_8567,N_6402,N_7767);
or U8568 (N_8568,N_7593,N_6707);
and U8569 (N_8569,N_6127,N_6869);
nor U8570 (N_8570,N_7097,N_7951);
or U8571 (N_8571,N_7547,N_6429);
and U8572 (N_8572,N_7081,N_7175);
and U8573 (N_8573,N_7473,N_7995);
nor U8574 (N_8574,N_7181,N_7529);
nand U8575 (N_8575,N_6025,N_7355);
nor U8576 (N_8576,N_6906,N_7683);
and U8577 (N_8577,N_7435,N_6696);
or U8578 (N_8578,N_7074,N_7534);
nor U8579 (N_8579,N_6979,N_7458);
and U8580 (N_8580,N_7614,N_7827);
and U8581 (N_8581,N_6614,N_7144);
or U8582 (N_8582,N_7254,N_6866);
nor U8583 (N_8583,N_6029,N_7334);
or U8584 (N_8584,N_6016,N_7555);
nand U8585 (N_8585,N_6675,N_6142);
nand U8586 (N_8586,N_6597,N_6589);
nand U8587 (N_8587,N_6444,N_7541);
nand U8588 (N_8588,N_6001,N_6300);
and U8589 (N_8589,N_7094,N_7055);
nand U8590 (N_8590,N_6415,N_6103);
and U8591 (N_8591,N_7586,N_7941);
or U8592 (N_8592,N_7340,N_6067);
and U8593 (N_8593,N_7638,N_6413);
nor U8594 (N_8594,N_6524,N_6042);
and U8595 (N_8595,N_7457,N_6969);
nand U8596 (N_8596,N_6786,N_7239);
nand U8597 (N_8597,N_7241,N_6823);
and U8598 (N_8598,N_7418,N_6270);
or U8599 (N_8599,N_7556,N_6335);
and U8600 (N_8600,N_6971,N_6298);
and U8601 (N_8601,N_7853,N_7712);
and U8602 (N_8602,N_6915,N_7354);
nor U8603 (N_8603,N_7298,N_6401);
nand U8604 (N_8604,N_7409,N_6742);
or U8605 (N_8605,N_7398,N_6746);
and U8606 (N_8606,N_7210,N_6373);
and U8607 (N_8607,N_6371,N_6245);
nor U8608 (N_8608,N_7494,N_7105);
or U8609 (N_8609,N_6126,N_7670);
or U8610 (N_8610,N_6461,N_7191);
or U8611 (N_8611,N_6876,N_6143);
nand U8612 (N_8612,N_7425,N_6819);
or U8613 (N_8613,N_6570,N_7656);
or U8614 (N_8614,N_6465,N_6792);
nand U8615 (N_8615,N_6954,N_6893);
nand U8616 (N_8616,N_7861,N_6065);
or U8617 (N_8617,N_6951,N_7983);
and U8618 (N_8618,N_7771,N_6964);
nor U8619 (N_8619,N_6459,N_6990);
nor U8620 (N_8620,N_6337,N_6530);
or U8621 (N_8621,N_7349,N_7030);
or U8622 (N_8622,N_7610,N_6080);
nor U8623 (N_8623,N_6050,N_6868);
or U8624 (N_8624,N_7744,N_7199);
or U8625 (N_8625,N_7002,N_7884);
nor U8626 (N_8626,N_7260,N_6333);
and U8627 (N_8627,N_6553,N_6903);
nand U8628 (N_8628,N_7774,N_7451);
nand U8629 (N_8629,N_6107,N_7583);
nor U8630 (N_8630,N_7028,N_7211);
nor U8631 (N_8631,N_6549,N_6120);
or U8632 (N_8632,N_6955,N_7625);
nand U8633 (N_8633,N_7545,N_7242);
and U8634 (N_8634,N_6594,N_6351);
nand U8635 (N_8635,N_6618,N_7492);
and U8636 (N_8636,N_6060,N_6193);
and U8637 (N_8637,N_6911,N_6995);
xor U8638 (N_8638,N_6663,N_6550);
nor U8639 (N_8639,N_7932,N_7218);
or U8640 (N_8640,N_7273,N_7070);
and U8641 (N_8641,N_6055,N_6063);
and U8642 (N_8642,N_7749,N_6313);
and U8643 (N_8643,N_6521,N_6771);
nor U8644 (N_8644,N_7866,N_7204);
or U8645 (N_8645,N_6718,N_6347);
or U8646 (N_8646,N_6306,N_6877);
and U8647 (N_8647,N_7266,N_7604);
and U8648 (N_8648,N_6334,N_6105);
and U8649 (N_8649,N_7393,N_7093);
or U8650 (N_8650,N_6261,N_6297);
nand U8651 (N_8651,N_7963,N_6822);
nor U8652 (N_8652,N_7071,N_7361);
nand U8653 (N_8653,N_7805,N_6555);
nor U8654 (N_8654,N_7069,N_7238);
or U8655 (N_8655,N_6889,N_6544);
and U8656 (N_8656,N_7244,N_7455);
or U8657 (N_8657,N_7036,N_7592);
and U8658 (N_8658,N_7352,N_6416);
or U8659 (N_8659,N_6481,N_7758);
nand U8660 (N_8660,N_6058,N_7405);
nor U8661 (N_8661,N_6427,N_6316);
nor U8662 (N_8662,N_7138,N_7917);
and U8663 (N_8663,N_7125,N_7893);
or U8664 (N_8664,N_6212,N_6491);
or U8665 (N_8665,N_7150,N_6484);
and U8666 (N_8666,N_6882,N_7157);
nor U8667 (N_8667,N_6030,N_7275);
nor U8668 (N_8668,N_6466,N_7183);
nor U8669 (N_8669,N_7139,N_6112);
or U8670 (N_8670,N_7468,N_6178);
or U8671 (N_8671,N_6651,N_6659);
or U8672 (N_8672,N_6256,N_7124);
or U8673 (N_8673,N_7379,N_7277);
or U8674 (N_8674,N_6825,N_7067);
or U8675 (N_8675,N_7760,N_6978);
or U8676 (N_8676,N_7407,N_6094);
nand U8677 (N_8677,N_7965,N_7564);
nor U8678 (N_8678,N_6935,N_6879);
xnor U8679 (N_8679,N_7814,N_7637);
nand U8680 (N_8680,N_7992,N_6621);
nor U8681 (N_8681,N_6354,N_6795);
nor U8682 (N_8682,N_6175,N_7158);
or U8683 (N_8683,N_6703,N_7697);
nand U8684 (N_8684,N_7718,N_6154);
and U8685 (N_8685,N_7141,N_7412);
nand U8686 (N_8686,N_6669,N_7090);
and U8687 (N_8687,N_6736,N_7162);
nor U8688 (N_8688,N_7922,N_7761);
and U8689 (N_8689,N_7524,N_6141);
nor U8690 (N_8690,N_6774,N_6545);
nor U8691 (N_8691,N_7546,N_6136);
or U8692 (N_8692,N_6387,N_6888);
and U8693 (N_8693,N_7278,N_6852);
nor U8694 (N_8694,N_7223,N_7110);
nor U8695 (N_8695,N_6433,N_7535);
or U8696 (N_8696,N_7599,N_6000);
nand U8697 (N_8697,N_7548,N_6150);
and U8698 (N_8698,N_7186,N_7845);
or U8699 (N_8699,N_7230,N_7258);
nor U8700 (N_8700,N_7633,N_7228);
nor U8701 (N_8701,N_7488,N_7411);
or U8702 (N_8702,N_7262,N_7287);
or U8703 (N_8703,N_6045,N_6800);
or U8704 (N_8704,N_7430,N_7479);
or U8705 (N_8705,N_7672,N_6411);
nand U8706 (N_8706,N_6973,N_6004);
and U8707 (N_8707,N_6331,N_6733);
and U8708 (N_8708,N_6255,N_6449);
and U8709 (N_8709,N_6765,N_6032);
nand U8710 (N_8710,N_6924,N_6608);
and U8711 (N_8711,N_7617,N_6661);
or U8712 (N_8712,N_6007,N_6383);
and U8713 (N_8713,N_6308,N_7496);
or U8714 (N_8714,N_7475,N_7601);
nand U8715 (N_8715,N_6044,N_7553);
or U8716 (N_8716,N_6939,N_7796);
nor U8717 (N_8717,N_6403,N_7106);
or U8718 (N_8718,N_7826,N_6972);
nor U8719 (N_8719,N_7628,N_7846);
nor U8720 (N_8720,N_7291,N_7728);
nand U8721 (N_8721,N_6203,N_7008);
nand U8722 (N_8722,N_6291,N_7961);
or U8723 (N_8723,N_7042,N_6912);
nor U8724 (N_8724,N_7197,N_7793);
and U8725 (N_8725,N_6542,N_7484);
nor U8726 (N_8726,N_6363,N_6470);
nor U8727 (N_8727,N_6533,N_6260);
nor U8728 (N_8728,N_6329,N_7416);
and U8729 (N_8729,N_7438,N_7143);
or U8730 (N_8730,N_7675,N_7660);
and U8731 (N_8731,N_6539,N_7989);
and U8732 (N_8732,N_6525,N_6492);
or U8733 (N_8733,N_6451,N_7474);
nand U8734 (N_8734,N_6395,N_7636);
nor U8735 (N_8735,N_6962,N_6655);
and U8736 (N_8736,N_7910,N_6926);
nand U8737 (N_8737,N_7649,N_7118);
nand U8738 (N_8738,N_7137,N_7431);
or U8739 (N_8739,N_7925,N_7086);
and U8740 (N_8740,N_7849,N_7879);
nand U8741 (N_8741,N_6494,N_6303);
and U8742 (N_8742,N_6548,N_7773);
xnor U8743 (N_8743,N_7730,N_6455);
or U8744 (N_8744,N_6384,N_6994);
nor U8745 (N_8745,N_7939,N_7891);
and U8746 (N_8746,N_6961,N_7315);
or U8747 (N_8747,N_6192,N_7123);
or U8748 (N_8748,N_7462,N_6937);
nor U8749 (N_8749,N_7310,N_6011);
or U8750 (N_8750,N_7065,N_7727);
and U8751 (N_8751,N_6468,N_7057);
and U8752 (N_8752,N_7358,N_7557);
nand U8753 (N_8753,N_6147,N_7324);
nor U8754 (N_8754,N_6650,N_6293);
nor U8755 (N_8755,N_7642,N_7214);
or U8756 (N_8756,N_7618,N_6322);
or U8757 (N_8757,N_7921,N_7135);
nand U8758 (N_8758,N_7517,N_6090);
nand U8759 (N_8759,N_7858,N_6619);
or U8760 (N_8760,N_7436,N_7051);
nand U8761 (N_8761,N_6325,N_7026);
nor U8762 (N_8762,N_6693,N_6278);
or U8763 (N_8763,N_6100,N_6842);
and U8764 (N_8764,N_7579,N_6871);
and U8765 (N_8765,N_6145,N_7240);
and U8766 (N_8766,N_6843,N_7077);
or U8767 (N_8767,N_6504,N_7606);
nor U8768 (N_8768,N_6266,N_7681);
or U8769 (N_8769,N_7061,N_6519);
nor U8770 (N_8770,N_6216,N_6104);
nor U8771 (N_8771,N_7235,N_6505);
nand U8772 (N_8772,N_7448,N_7590);
or U8773 (N_8773,N_7308,N_7777);
nand U8774 (N_8774,N_6059,N_7276);
nand U8775 (N_8775,N_6422,N_7857);
nand U8776 (N_8776,N_6040,N_7434);
nand U8777 (N_8777,N_7248,N_6111);
nand U8778 (N_8778,N_6177,N_6609);
and U8779 (N_8779,N_7868,N_6023);
nor U8780 (N_8780,N_7180,N_6423);
and U8781 (N_8781,N_6830,N_6516);
nor U8782 (N_8782,N_6400,N_6410);
nor U8783 (N_8783,N_7918,N_6627);
and U8784 (N_8784,N_6695,N_6254);
nor U8785 (N_8785,N_6359,N_7549);
nor U8786 (N_8786,N_6789,N_6475);
and U8787 (N_8787,N_7406,N_7662);
nor U8788 (N_8788,N_7785,N_6252);
nand U8789 (N_8789,N_7694,N_6885);
nand U8790 (N_8790,N_7027,N_7489);
or U8791 (N_8791,N_6035,N_7536);
nor U8792 (N_8792,N_7052,N_6841);
nand U8793 (N_8793,N_6096,N_6161);
nor U8794 (N_8794,N_7527,N_6366);
and U8795 (N_8795,N_7397,N_6089);
nor U8796 (N_8796,N_6265,N_7439);
and U8797 (N_8797,N_6541,N_6887);
nand U8798 (N_8798,N_7085,N_7390);
and U8799 (N_8799,N_6389,N_6845);
or U8800 (N_8800,N_6922,N_7609);
and U8801 (N_8801,N_6768,N_6304);
or U8802 (N_8802,N_6770,N_6960);
or U8803 (N_8803,N_7472,N_6204);
and U8804 (N_8804,N_7821,N_6388);
nor U8805 (N_8805,N_7299,N_7595);
nor U8806 (N_8806,N_7232,N_7511);
nor U8807 (N_8807,N_7550,N_7053);
or U8808 (N_8808,N_6457,N_6855);
and U8809 (N_8809,N_7025,N_7924);
nor U8810 (N_8810,N_6925,N_6378);
nor U8811 (N_8811,N_7788,N_7317);
nor U8812 (N_8812,N_6227,N_6271);
nand U8813 (N_8813,N_6149,N_7429);
or U8814 (N_8814,N_7461,N_6895);
nand U8815 (N_8815,N_7769,N_7903);
nor U8816 (N_8816,N_6694,N_6896);
nand U8817 (N_8817,N_6274,N_6708);
nand U8818 (N_8818,N_6643,N_7509);
and U8819 (N_8819,N_7539,N_7578);
or U8820 (N_8820,N_7338,N_6397);
and U8821 (N_8821,N_6723,N_7940);
and U8822 (N_8822,N_6679,N_6956);
and U8823 (N_8823,N_7127,N_7400);
or U8824 (N_8824,N_6691,N_6716);
nand U8825 (N_8825,N_6195,N_6821);
and U8826 (N_8826,N_7707,N_6489);
nor U8827 (N_8827,N_7704,N_6543);
and U8828 (N_8828,N_7348,N_7948);
nor U8829 (N_8829,N_6008,N_7801);
nand U8830 (N_8830,N_7224,N_7929);
nand U8831 (N_8831,N_7589,N_6966);
nor U8832 (N_8832,N_7318,N_7872);
or U8833 (N_8833,N_6666,N_7831);
and U8834 (N_8834,N_6537,N_7095);
or U8835 (N_8835,N_6750,N_7603);
and U8836 (N_8836,N_6788,N_7054);
xor U8837 (N_8837,N_6095,N_7708);
nand U8838 (N_8838,N_7038,N_7913);
nor U8839 (N_8839,N_6917,N_6846);
or U8840 (N_8840,N_6349,N_6575);
nand U8841 (N_8841,N_6355,N_7894);
or U8842 (N_8842,N_6642,N_7639);
and U8843 (N_8843,N_7969,N_6224);
nand U8844 (N_8844,N_7120,N_6487);
and U8845 (N_8845,N_7079,N_7982);
or U8846 (N_8846,N_6220,N_6637);
nor U8847 (N_8847,N_7677,N_6200);
nor U8848 (N_8848,N_6406,N_6495);
nand U8849 (N_8849,N_7471,N_7156);
nand U8850 (N_8850,N_6326,N_7221);
nor U8851 (N_8851,N_7756,N_6075);
nor U8852 (N_8852,N_7087,N_7828);
nand U8853 (N_8853,N_7737,N_7233);
or U8854 (N_8854,N_6408,N_7364);
nand U8855 (N_8855,N_7062,N_6740);
and U8856 (N_8856,N_7611,N_6563);
nand U8857 (N_8857,N_6038,N_7185);
nand U8858 (N_8858,N_6467,N_7388);
nand U8859 (N_8859,N_7726,N_6834);
and U8860 (N_8860,N_6078,N_7803);
and U8861 (N_8861,N_6289,N_7909);
xnor U8862 (N_8862,N_6176,N_7585);
nand U8863 (N_8863,N_7563,N_7367);
or U8864 (N_8864,N_7836,N_6310);
and U8865 (N_8865,N_7518,N_7765);
nor U8866 (N_8866,N_7432,N_6577);
nor U8867 (N_8867,N_7902,N_7923);
nor U8868 (N_8868,N_7877,N_6766);
or U8869 (N_8869,N_6749,N_7368);
nand U8870 (N_8870,N_7344,N_6557);
and U8871 (N_8871,N_6365,N_6012);
nand U8872 (N_8872,N_6264,N_7680);
or U8873 (N_8873,N_6314,N_7490);
nor U8874 (N_8874,N_6891,N_6476);
or U8875 (N_8875,N_7573,N_7312);
nand U8876 (N_8876,N_7797,N_6894);
nand U8877 (N_8877,N_7103,N_7906);
or U8878 (N_8878,N_6231,N_6737);
nand U8879 (N_8879,N_6281,N_7852);
nor U8880 (N_8880,N_7996,N_7560);
nand U8881 (N_8881,N_7986,N_7674);
or U8882 (N_8882,N_6123,N_7245);
and U8883 (N_8883,N_6807,N_7591);
nor U8884 (N_8884,N_6974,N_7817);
and U8885 (N_8885,N_7041,N_7753);
nand U8886 (N_8886,N_7295,N_6249);
nand U8887 (N_8887,N_7904,N_6377);
nor U8888 (N_8888,N_7082,N_6037);
and U8889 (N_8889,N_7895,N_7653);
and U8890 (N_8890,N_7374,N_7998);
or U8891 (N_8891,N_6686,N_6172);
nand U8892 (N_8892,N_7325,N_6725);
nor U8893 (N_8893,N_6873,N_6713);
and U8894 (N_8894,N_6341,N_7116);
and U8895 (N_8895,N_6109,N_6988);
nor U8896 (N_8896,N_7888,N_6091);
nand U8897 (N_8897,N_6865,N_6452);
nor U8898 (N_8898,N_6194,N_7844);
and U8899 (N_8899,N_7798,N_6534);
nand U8900 (N_8900,N_6157,N_6497);
nor U8901 (N_8901,N_6253,N_6130);
xnor U8902 (N_8902,N_6688,N_7691);
or U8903 (N_8903,N_6963,N_6381);
nand U8904 (N_8904,N_7999,N_7738);
nor U8905 (N_8905,N_6394,N_7855);
nor U8906 (N_8906,N_6028,N_7938);
or U8907 (N_8907,N_6248,N_6741);
nor U8908 (N_8908,N_6064,N_7387);
and U8909 (N_8909,N_7993,N_6409);
nand U8910 (N_8910,N_7812,N_6364);
nand U8911 (N_8911,N_6338,N_7870);
nand U8912 (N_8912,N_7177,N_7037);
and U8913 (N_8913,N_6190,N_6432);
nor U8914 (N_8914,N_7142,N_6620);
nor U8915 (N_8915,N_6230,N_7443);
nor U8916 (N_8916,N_6970,N_7363);
nor U8917 (N_8917,N_7384,N_6699);
and U8918 (N_8918,N_6989,N_6835);
nand U8919 (N_8919,N_7781,N_7022);
and U8920 (N_8920,N_6332,N_6259);
nand U8921 (N_8921,N_6183,N_7687);
nand U8922 (N_8922,N_6344,N_7813);
and U8923 (N_8923,N_6290,N_6739);
and U8924 (N_8924,N_7958,N_6513);
or U8925 (N_8925,N_7216,N_6241);
nor U8926 (N_8926,N_7229,N_7414);
and U8927 (N_8927,N_7957,N_6919);
or U8928 (N_8928,N_6288,N_7493);
nor U8929 (N_8929,N_6239,N_6914);
nor U8930 (N_8930,N_6769,N_6776);
or U8931 (N_8931,N_7225,N_7896);
or U8932 (N_8932,N_6295,N_7169);
or U8933 (N_8933,N_6348,N_7128);
xnor U8934 (N_8934,N_7442,N_7383);
and U8935 (N_8935,N_7502,N_7745);
or U8936 (N_8936,N_7063,N_6762);
nand U8937 (N_8937,N_7172,N_7713);
nor U8938 (N_8938,N_7886,N_7977);
or U8939 (N_8939,N_7171,N_6277);
or U8940 (N_8940,N_7460,N_7967);
nand U8941 (N_8941,N_6031,N_7970);
nor U8942 (N_8942,N_7685,N_7089);
nor U8943 (N_8943,N_6640,N_7203);
nor U8944 (N_8944,N_7319,N_7657);
nor U8945 (N_8945,N_6319,N_6324);
nand U8946 (N_8946,N_6250,N_6071);
and U8947 (N_8947,N_6836,N_6929);
nand U8948 (N_8948,N_7615,N_7973);
nand U8949 (N_8949,N_7659,N_7746);
nand U8950 (N_8950,N_7641,N_6445);
nand U8951 (N_8951,N_6479,N_6657);
nand U8952 (N_8952,N_7024,N_6654);
nand U8953 (N_8953,N_6034,N_7878);
and U8954 (N_8954,N_6144,N_6369);
or U8955 (N_8955,N_6665,N_7843);
and U8956 (N_8956,N_7307,N_6647);
or U8957 (N_8957,N_7500,N_7441);
and U8958 (N_8958,N_6587,N_6859);
and U8959 (N_8959,N_7671,N_7272);
nor U8960 (N_8960,N_6631,N_7486);
xor U8961 (N_8961,N_6756,N_6083);
and U8962 (N_8962,N_7160,N_6592);
nand U8963 (N_8963,N_6747,N_6148);
and U8964 (N_8964,N_7292,N_6263);
nor U8965 (N_8965,N_7800,N_6784);
nor U8966 (N_8966,N_6763,N_6454);
and U8967 (N_8967,N_6983,N_6920);
or U8968 (N_8968,N_7445,N_6217);
nor U8969 (N_8969,N_6066,N_7565);
nor U8970 (N_8970,N_7198,N_7766);
nor U8971 (N_8971,N_6179,N_7525);
or U8972 (N_8972,N_6601,N_7401);
and U8973 (N_8973,N_7602,N_6671);
nor U8974 (N_8974,N_6047,N_7246);
or U8975 (N_8975,N_7220,N_6892);
nor U8976 (N_8976,N_6146,N_7263);
or U8977 (N_8977,N_6056,N_6606);
nor U8978 (N_8978,N_7173,N_7823);
and U8979 (N_8979,N_6880,N_6780);
nor U8980 (N_8980,N_6913,N_6405);
or U8981 (N_8981,N_7154,N_6588);
xor U8982 (N_8982,N_6294,N_7119);
and U8983 (N_8983,N_6848,N_7029);
nand U8984 (N_8984,N_7631,N_7540);
and U8985 (N_8985,N_6787,N_7111);
and U8986 (N_8986,N_7506,N_7701);
or U8987 (N_8987,N_6404,N_6727);
nor U8988 (N_8988,N_6122,N_6417);
or U8989 (N_8989,N_6299,N_6898);
or U8990 (N_8990,N_7267,N_7132);
nand U8991 (N_8991,N_7780,N_6861);
or U8992 (N_8992,N_7329,N_6114);
and U8993 (N_8993,N_7806,N_7316);
or U8994 (N_8994,N_7543,N_6017);
nand U8995 (N_8995,N_7366,N_7889);
nand U8996 (N_8996,N_6734,N_6081);
or U8997 (N_8997,N_7972,N_7013);
and U8998 (N_8998,N_7328,N_6656);
nand U8999 (N_8999,N_6188,N_6398);
nor U9000 (N_9000,N_6466,N_7873);
nor U9001 (N_9001,N_6991,N_6828);
nor U9002 (N_9002,N_6190,N_7218);
and U9003 (N_9003,N_6388,N_6083);
or U9004 (N_9004,N_7809,N_7141);
nor U9005 (N_9005,N_7567,N_7752);
or U9006 (N_9006,N_7913,N_7004);
or U9007 (N_9007,N_7478,N_7180);
nand U9008 (N_9008,N_7654,N_7198);
nor U9009 (N_9009,N_6394,N_7149);
nand U9010 (N_9010,N_7749,N_6915);
nor U9011 (N_9011,N_6518,N_7177);
nor U9012 (N_9012,N_6195,N_7130);
nor U9013 (N_9013,N_7839,N_6159);
and U9014 (N_9014,N_7452,N_7451);
and U9015 (N_9015,N_7801,N_7457);
nand U9016 (N_9016,N_7928,N_6395);
nand U9017 (N_9017,N_6940,N_7481);
nand U9018 (N_9018,N_6146,N_7474);
or U9019 (N_9019,N_7252,N_7132);
or U9020 (N_9020,N_6582,N_6792);
nor U9021 (N_9021,N_6247,N_7432);
nand U9022 (N_9022,N_7414,N_6684);
nor U9023 (N_9023,N_6688,N_7839);
nand U9024 (N_9024,N_6187,N_7255);
nor U9025 (N_9025,N_7790,N_6181);
or U9026 (N_9026,N_7066,N_7221);
or U9027 (N_9027,N_6209,N_6420);
and U9028 (N_9028,N_7043,N_7200);
or U9029 (N_9029,N_6398,N_7664);
nor U9030 (N_9030,N_6332,N_6489);
nand U9031 (N_9031,N_6575,N_7329);
or U9032 (N_9032,N_6477,N_6625);
and U9033 (N_9033,N_7089,N_7317);
or U9034 (N_9034,N_6767,N_6698);
nor U9035 (N_9035,N_6941,N_6888);
nor U9036 (N_9036,N_7848,N_6688);
nor U9037 (N_9037,N_7723,N_6926);
nor U9038 (N_9038,N_7760,N_7676);
or U9039 (N_9039,N_7072,N_7890);
nor U9040 (N_9040,N_6988,N_7046);
nand U9041 (N_9041,N_6952,N_6147);
nor U9042 (N_9042,N_6711,N_6693);
nand U9043 (N_9043,N_7038,N_6003);
nor U9044 (N_9044,N_7455,N_6754);
and U9045 (N_9045,N_6827,N_7121);
or U9046 (N_9046,N_6967,N_7502);
or U9047 (N_9047,N_6887,N_6406);
nand U9048 (N_9048,N_7266,N_7477);
and U9049 (N_9049,N_7664,N_6831);
or U9050 (N_9050,N_6171,N_7309);
xor U9051 (N_9051,N_7064,N_6829);
nor U9052 (N_9052,N_7826,N_7989);
nor U9053 (N_9053,N_6175,N_6140);
nor U9054 (N_9054,N_6381,N_7819);
nand U9055 (N_9055,N_6255,N_6989);
and U9056 (N_9056,N_7556,N_6747);
nor U9057 (N_9057,N_7039,N_6458);
or U9058 (N_9058,N_7710,N_6382);
nand U9059 (N_9059,N_6555,N_7292);
nand U9060 (N_9060,N_7047,N_6962);
or U9061 (N_9061,N_6716,N_6860);
nand U9062 (N_9062,N_6601,N_7157);
and U9063 (N_9063,N_7777,N_6306);
and U9064 (N_9064,N_7138,N_7123);
and U9065 (N_9065,N_7005,N_6412);
nand U9066 (N_9066,N_6952,N_7513);
nor U9067 (N_9067,N_6893,N_6916);
nand U9068 (N_9068,N_6930,N_7290);
or U9069 (N_9069,N_6276,N_6399);
nand U9070 (N_9070,N_7333,N_7334);
nand U9071 (N_9071,N_7059,N_7562);
nor U9072 (N_9072,N_7508,N_6157);
and U9073 (N_9073,N_7673,N_6175);
and U9074 (N_9074,N_7198,N_7459);
nor U9075 (N_9075,N_7289,N_6235);
xor U9076 (N_9076,N_7915,N_7959);
nand U9077 (N_9077,N_6817,N_7877);
nand U9078 (N_9078,N_6653,N_7146);
nand U9079 (N_9079,N_7766,N_7778);
nor U9080 (N_9080,N_6597,N_7082);
and U9081 (N_9081,N_7154,N_6737);
and U9082 (N_9082,N_7372,N_7333);
nand U9083 (N_9083,N_7156,N_6551);
nand U9084 (N_9084,N_6215,N_6917);
and U9085 (N_9085,N_6406,N_7432);
nand U9086 (N_9086,N_7777,N_7222);
nand U9087 (N_9087,N_7675,N_7859);
nor U9088 (N_9088,N_6357,N_6447);
and U9089 (N_9089,N_6990,N_7372);
nor U9090 (N_9090,N_7366,N_6105);
nand U9091 (N_9091,N_7210,N_7810);
nor U9092 (N_9092,N_7389,N_6658);
nor U9093 (N_9093,N_7346,N_6636);
nand U9094 (N_9094,N_6029,N_6818);
or U9095 (N_9095,N_7827,N_7025);
nand U9096 (N_9096,N_7694,N_7055);
and U9097 (N_9097,N_6929,N_6170);
nor U9098 (N_9098,N_6921,N_7159);
or U9099 (N_9099,N_7559,N_6197);
nand U9100 (N_9100,N_7915,N_7656);
or U9101 (N_9101,N_7592,N_6768);
or U9102 (N_9102,N_6150,N_6985);
nand U9103 (N_9103,N_6048,N_7994);
nand U9104 (N_9104,N_7127,N_7741);
nand U9105 (N_9105,N_7721,N_7008);
nor U9106 (N_9106,N_6069,N_7611);
nand U9107 (N_9107,N_6337,N_6836);
and U9108 (N_9108,N_7056,N_6745);
and U9109 (N_9109,N_6271,N_6062);
xor U9110 (N_9110,N_7190,N_7103);
and U9111 (N_9111,N_7535,N_6886);
nand U9112 (N_9112,N_7954,N_6440);
or U9113 (N_9113,N_7057,N_7353);
nor U9114 (N_9114,N_6351,N_6256);
nand U9115 (N_9115,N_6397,N_6842);
nand U9116 (N_9116,N_7466,N_6968);
or U9117 (N_9117,N_6669,N_6379);
nor U9118 (N_9118,N_6809,N_6342);
or U9119 (N_9119,N_7199,N_7978);
nor U9120 (N_9120,N_7313,N_7430);
and U9121 (N_9121,N_6381,N_7381);
xor U9122 (N_9122,N_6623,N_7339);
and U9123 (N_9123,N_7911,N_6529);
and U9124 (N_9124,N_7966,N_7587);
and U9125 (N_9125,N_6016,N_7711);
or U9126 (N_9126,N_7057,N_7667);
nor U9127 (N_9127,N_6098,N_6859);
or U9128 (N_9128,N_6315,N_6560);
or U9129 (N_9129,N_7803,N_7531);
nand U9130 (N_9130,N_6134,N_7200);
and U9131 (N_9131,N_7840,N_6373);
or U9132 (N_9132,N_6169,N_6603);
and U9133 (N_9133,N_6613,N_6539);
and U9134 (N_9134,N_7068,N_7832);
nand U9135 (N_9135,N_6273,N_7862);
and U9136 (N_9136,N_6045,N_7496);
and U9137 (N_9137,N_6314,N_6899);
nor U9138 (N_9138,N_6492,N_6809);
nor U9139 (N_9139,N_7376,N_6267);
nor U9140 (N_9140,N_6599,N_6424);
or U9141 (N_9141,N_7895,N_6750);
nand U9142 (N_9142,N_6019,N_6035);
and U9143 (N_9143,N_7813,N_7584);
nor U9144 (N_9144,N_6081,N_7283);
nor U9145 (N_9145,N_7972,N_7340);
nand U9146 (N_9146,N_7303,N_6407);
or U9147 (N_9147,N_6832,N_6497);
or U9148 (N_9148,N_6386,N_7293);
nor U9149 (N_9149,N_7533,N_6848);
nand U9150 (N_9150,N_6468,N_6533);
nand U9151 (N_9151,N_7719,N_7131);
and U9152 (N_9152,N_7597,N_6035);
or U9153 (N_9153,N_7040,N_6940);
nor U9154 (N_9154,N_7552,N_6902);
or U9155 (N_9155,N_7344,N_7891);
or U9156 (N_9156,N_6072,N_6415);
nor U9157 (N_9157,N_6612,N_6465);
nor U9158 (N_9158,N_6024,N_6070);
nor U9159 (N_9159,N_6840,N_7175);
nand U9160 (N_9160,N_7138,N_7296);
nor U9161 (N_9161,N_6494,N_7041);
or U9162 (N_9162,N_7454,N_7589);
nand U9163 (N_9163,N_7219,N_7518);
and U9164 (N_9164,N_6997,N_7695);
nand U9165 (N_9165,N_6770,N_7958);
xnor U9166 (N_9166,N_7924,N_6077);
nand U9167 (N_9167,N_7801,N_7392);
nand U9168 (N_9168,N_7994,N_7321);
nor U9169 (N_9169,N_6219,N_7702);
or U9170 (N_9170,N_6752,N_7764);
or U9171 (N_9171,N_7311,N_7079);
nand U9172 (N_9172,N_7178,N_7306);
or U9173 (N_9173,N_7330,N_6396);
nor U9174 (N_9174,N_6996,N_7309);
or U9175 (N_9175,N_6030,N_7465);
nand U9176 (N_9176,N_7398,N_6868);
or U9177 (N_9177,N_7637,N_7941);
nor U9178 (N_9178,N_7531,N_6803);
or U9179 (N_9179,N_6458,N_7806);
nand U9180 (N_9180,N_6322,N_7373);
nand U9181 (N_9181,N_6930,N_7401);
or U9182 (N_9182,N_6913,N_6292);
and U9183 (N_9183,N_6598,N_6955);
and U9184 (N_9184,N_6678,N_7873);
nor U9185 (N_9185,N_7091,N_7854);
nand U9186 (N_9186,N_6579,N_7302);
and U9187 (N_9187,N_7059,N_6207);
nor U9188 (N_9188,N_7655,N_7379);
or U9189 (N_9189,N_6044,N_7679);
or U9190 (N_9190,N_7091,N_6784);
nand U9191 (N_9191,N_6240,N_7176);
or U9192 (N_9192,N_6488,N_7470);
and U9193 (N_9193,N_7922,N_6120);
or U9194 (N_9194,N_6664,N_7222);
or U9195 (N_9195,N_7629,N_7125);
and U9196 (N_9196,N_6092,N_6493);
and U9197 (N_9197,N_7541,N_6916);
or U9198 (N_9198,N_6095,N_6315);
nor U9199 (N_9199,N_7088,N_6053);
nand U9200 (N_9200,N_7092,N_6001);
and U9201 (N_9201,N_6218,N_7797);
nand U9202 (N_9202,N_7419,N_6612);
nor U9203 (N_9203,N_7359,N_6043);
nand U9204 (N_9204,N_7557,N_6495);
or U9205 (N_9205,N_7896,N_6621);
nor U9206 (N_9206,N_6254,N_6169);
or U9207 (N_9207,N_7587,N_6783);
and U9208 (N_9208,N_6065,N_7057);
or U9209 (N_9209,N_7847,N_7854);
nand U9210 (N_9210,N_7309,N_7598);
nand U9211 (N_9211,N_6359,N_6736);
nor U9212 (N_9212,N_7588,N_6121);
and U9213 (N_9213,N_6497,N_6840);
nor U9214 (N_9214,N_6081,N_6248);
nand U9215 (N_9215,N_6629,N_6669);
nor U9216 (N_9216,N_6332,N_6711);
or U9217 (N_9217,N_7968,N_7553);
and U9218 (N_9218,N_6294,N_7406);
nor U9219 (N_9219,N_6274,N_7516);
or U9220 (N_9220,N_6753,N_6080);
nor U9221 (N_9221,N_6578,N_7342);
nand U9222 (N_9222,N_6863,N_6349);
nor U9223 (N_9223,N_6217,N_6757);
or U9224 (N_9224,N_7367,N_6571);
and U9225 (N_9225,N_7370,N_7493);
nor U9226 (N_9226,N_6904,N_7084);
nand U9227 (N_9227,N_6075,N_7524);
or U9228 (N_9228,N_6434,N_7917);
nor U9229 (N_9229,N_6954,N_6076);
or U9230 (N_9230,N_7492,N_6080);
nor U9231 (N_9231,N_7998,N_7913);
or U9232 (N_9232,N_6090,N_7260);
nor U9233 (N_9233,N_6058,N_6168);
xor U9234 (N_9234,N_7404,N_7370);
nor U9235 (N_9235,N_6075,N_7715);
and U9236 (N_9236,N_6193,N_6399);
and U9237 (N_9237,N_6242,N_7334);
and U9238 (N_9238,N_6239,N_7121);
or U9239 (N_9239,N_6234,N_6213);
nor U9240 (N_9240,N_7206,N_6304);
and U9241 (N_9241,N_7137,N_7767);
and U9242 (N_9242,N_6458,N_6877);
and U9243 (N_9243,N_6135,N_6777);
or U9244 (N_9244,N_6597,N_6420);
nor U9245 (N_9245,N_6816,N_6448);
nor U9246 (N_9246,N_6326,N_6531);
nand U9247 (N_9247,N_7477,N_6857);
and U9248 (N_9248,N_7924,N_7298);
or U9249 (N_9249,N_7794,N_6354);
nor U9250 (N_9250,N_6327,N_7042);
nand U9251 (N_9251,N_7053,N_6201);
nand U9252 (N_9252,N_7220,N_7585);
nand U9253 (N_9253,N_6197,N_7584);
nor U9254 (N_9254,N_6985,N_6568);
and U9255 (N_9255,N_6653,N_7047);
nor U9256 (N_9256,N_6914,N_7652);
nand U9257 (N_9257,N_6044,N_7292);
or U9258 (N_9258,N_7591,N_6298);
nor U9259 (N_9259,N_7074,N_7776);
or U9260 (N_9260,N_7350,N_6615);
nor U9261 (N_9261,N_7219,N_6316);
and U9262 (N_9262,N_6459,N_7473);
nand U9263 (N_9263,N_6246,N_6415);
nand U9264 (N_9264,N_7412,N_6041);
nor U9265 (N_9265,N_6979,N_6676);
or U9266 (N_9266,N_6532,N_6497);
nor U9267 (N_9267,N_6992,N_7299);
nand U9268 (N_9268,N_7470,N_7445);
or U9269 (N_9269,N_6586,N_6920);
nor U9270 (N_9270,N_7284,N_7094);
or U9271 (N_9271,N_7481,N_7254);
nor U9272 (N_9272,N_6607,N_6797);
or U9273 (N_9273,N_6597,N_7366);
nor U9274 (N_9274,N_6882,N_6838);
or U9275 (N_9275,N_7593,N_6038);
nor U9276 (N_9276,N_7879,N_6658);
nand U9277 (N_9277,N_7492,N_7357);
and U9278 (N_9278,N_6605,N_7789);
and U9279 (N_9279,N_6821,N_6947);
or U9280 (N_9280,N_6449,N_7356);
xor U9281 (N_9281,N_7733,N_6854);
or U9282 (N_9282,N_7750,N_7508);
nand U9283 (N_9283,N_7852,N_7859);
nor U9284 (N_9284,N_7484,N_6678);
and U9285 (N_9285,N_6595,N_7399);
and U9286 (N_9286,N_6277,N_6757);
nand U9287 (N_9287,N_7950,N_6421);
nor U9288 (N_9288,N_7965,N_6178);
and U9289 (N_9289,N_6809,N_6505);
or U9290 (N_9290,N_6362,N_6018);
nor U9291 (N_9291,N_7582,N_7474);
nand U9292 (N_9292,N_7064,N_6693);
nor U9293 (N_9293,N_7442,N_6300);
or U9294 (N_9294,N_7365,N_7898);
nor U9295 (N_9295,N_7523,N_6289);
nor U9296 (N_9296,N_6353,N_7416);
and U9297 (N_9297,N_6589,N_7151);
and U9298 (N_9298,N_6068,N_6990);
nand U9299 (N_9299,N_7336,N_6760);
nand U9300 (N_9300,N_6040,N_7769);
or U9301 (N_9301,N_7686,N_7359);
or U9302 (N_9302,N_7114,N_7591);
nand U9303 (N_9303,N_7986,N_7895);
or U9304 (N_9304,N_6885,N_7324);
and U9305 (N_9305,N_7147,N_6527);
nor U9306 (N_9306,N_7353,N_7478);
and U9307 (N_9307,N_7531,N_6363);
nor U9308 (N_9308,N_7462,N_7609);
and U9309 (N_9309,N_6989,N_6710);
nand U9310 (N_9310,N_7011,N_6624);
nand U9311 (N_9311,N_7805,N_6599);
nor U9312 (N_9312,N_7715,N_6308);
nor U9313 (N_9313,N_6105,N_6197);
nor U9314 (N_9314,N_7581,N_7954);
and U9315 (N_9315,N_6067,N_7117);
or U9316 (N_9316,N_7471,N_6453);
or U9317 (N_9317,N_7593,N_6615);
nand U9318 (N_9318,N_7086,N_6106);
nor U9319 (N_9319,N_7986,N_7328);
or U9320 (N_9320,N_7504,N_7032);
and U9321 (N_9321,N_6072,N_6230);
nand U9322 (N_9322,N_7526,N_6411);
and U9323 (N_9323,N_7755,N_7279);
xnor U9324 (N_9324,N_6873,N_6862);
and U9325 (N_9325,N_7128,N_7821);
or U9326 (N_9326,N_7598,N_7006);
and U9327 (N_9327,N_7560,N_6410);
nand U9328 (N_9328,N_7409,N_6231);
and U9329 (N_9329,N_7343,N_7105);
and U9330 (N_9330,N_6205,N_6957);
or U9331 (N_9331,N_6744,N_7773);
and U9332 (N_9332,N_7237,N_6672);
nand U9333 (N_9333,N_6755,N_7842);
and U9334 (N_9334,N_7479,N_7090);
nor U9335 (N_9335,N_6449,N_7734);
nand U9336 (N_9336,N_7343,N_7237);
and U9337 (N_9337,N_6975,N_6804);
nand U9338 (N_9338,N_7864,N_7541);
and U9339 (N_9339,N_7024,N_7535);
or U9340 (N_9340,N_6806,N_6739);
nor U9341 (N_9341,N_6754,N_7381);
and U9342 (N_9342,N_7833,N_7670);
nand U9343 (N_9343,N_7239,N_6217);
nor U9344 (N_9344,N_7593,N_6226);
nand U9345 (N_9345,N_6054,N_7378);
and U9346 (N_9346,N_6543,N_7159);
or U9347 (N_9347,N_7591,N_6864);
nor U9348 (N_9348,N_7921,N_7607);
or U9349 (N_9349,N_7750,N_6513);
nand U9350 (N_9350,N_6886,N_7334);
nand U9351 (N_9351,N_6488,N_6331);
nand U9352 (N_9352,N_7354,N_7619);
or U9353 (N_9353,N_7155,N_6485);
or U9354 (N_9354,N_7444,N_7884);
and U9355 (N_9355,N_7772,N_7608);
and U9356 (N_9356,N_6582,N_7025);
and U9357 (N_9357,N_7473,N_7533);
and U9358 (N_9358,N_6062,N_7405);
or U9359 (N_9359,N_7470,N_7935);
nand U9360 (N_9360,N_7330,N_7519);
nand U9361 (N_9361,N_7838,N_7334);
and U9362 (N_9362,N_6411,N_7636);
nor U9363 (N_9363,N_7219,N_7621);
nor U9364 (N_9364,N_7414,N_7101);
nand U9365 (N_9365,N_7239,N_7154);
and U9366 (N_9366,N_6630,N_7551);
and U9367 (N_9367,N_6943,N_7516);
nor U9368 (N_9368,N_6157,N_6881);
and U9369 (N_9369,N_6294,N_7154);
or U9370 (N_9370,N_6505,N_6940);
and U9371 (N_9371,N_7258,N_6847);
nand U9372 (N_9372,N_6309,N_6611);
or U9373 (N_9373,N_6191,N_6938);
nor U9374 (N_9374,N_7606,N_7310);
nor U9375 (N_9375,N_7841,N_7978);
and U9376 (N_9376,N_7292,N_7279);
and U9377 (N_9377,N_6367,N_7999);
and U9378 (N_9378,N_7098,N_7640);
nor U9379 (N_9379,N_6236,N_6030);
nand U9380 (N_9380,N_7135,N_6441);
or U9381 (N_9381,N_7242,N_7485);
or U9382 (N_9382,N_7836,N_7084);
and U9383 (N_9383,N_7699,N_7384);
nor U9384 (N_9384,N_7968,N_7824);
and U9385 (N_9385,N_6506,N_7520);
nand U9386 (N_9386,N_6349,N_6037);
nand U9387 (N_9387,N_7626,N_6561);
nor U9388 (N_9388,N_7334,N_6380);
nand U9389 (N_9389,N_6219,N_6925);
nor U9390 (N_9390,N_6866,N_7340);
or U9391 (N_9391,N_6473,N_6585);
nor U9392 (N_9392,N_6554,N_7713);
and U9393 (N_9393,N_7242,N_6561);
and U9394 (N_9394,N_7257,N_6808);
or U9395 (N_9395,N_7821,N_7240);
or U9396 (N_9396,N_7929,N_6487);
and U9397 (N_9397,N_7897,N_7522);
nor U9398 (N_9398,N_6248,N_6886);
or U9399 (N_9399,N_6489,N_7778);
nor U9400 (N_9400,N_6899,N_7594);
nor U9401 (N_9401,N_7169,N_7319);
nand U9402 (N_9402,N_7762,N_7130);
and U9403 (N_9403,N_7470,N_6545);
nand U9404 (N_9404,N_6945,N_6529);
nand U9405 (N_9405,N_6166,N_6763);
nor U9406 (N_9406,N_6001,N_7298);
or U9407 (N_9407,N_6465,N_7040);
nor U9408 (N_9408,N_6367,N_6078);
nand U9409 (N_9409,N_7776,N_7738);
and U9410 (N_9410,N_6812,N_6013);
nor U9411 (N_9411,N_6687,N_6863);
nand U9412 (N_9412,N_6018,N_6853);
nor U9413 (N_9413,N_7210,N_6105);
nand U9414 (N_9414,N_7468,N_7270);
or U9415 (N_9415,N_6913,N_7776);
nor U9416 (N_9416,N_6939,N_7866);
and U9417 (N_9417,N_7831,N_6190);
nand U9418 (N_9418,N_7659,N_6728);
and U9419 (N_9419,N_7125,N_6492);
and U9420 (N_9420,N_6982,N_7971);
nand U9421 (N_9421,N_6775,N_6762);
and U9422 (N_9422,N_6073,N_6698);
nor U9423 (N_9423,N_7195,N_7656);
nor U9424 (N_9424,N_7993,N_7765);
or U9425 (N_9425,N_7287,N_7552);
nor U9426 (N_9426,N_6686,N_7611);
nor U9427 (N_9427,N_6810,N_6329);
nor U9428 (N_9428,N_7858,N_7772);
and U9429 (N_9429,N_7346,N_7301);
nand U9430 (N_9430,N_7257,N_7433);
nor U9431 (N_9431,N_7716,N_6743);
or U9432 (N_9432,N_6745,N_6960);
and U9433 (N_9433,N_7587,N_6464);
or U9434 (N_9434,N_6367,N_6229);
or U9435 (N_9435,N_7219,N_6840);
nor U9436 (N_9436,N_7778,N_7545);
nand U9437 (N_9437,N_7769,N_6275);
nor U9438 (N_9438,N_6444,N_7391);
nand U9439 (N_9439,N_7894,N_6738);
nor U9440 (N_9440,N_7566,N_6767);
or U9441 (N_9441,N_6617,N_7990);
and U9442 (N_9442,N_6887,N_7701);
or U9443 (N_9443,N_6902,N_7568);
nor U9444 (N_9444,N_7956,N_6688);
and U9445 (N_9445,N_7019,N_7605);
nand U9446 (N_9446,N_7320,N_6540);
nand U9447 (N_9447,N_6051,N_7144);
nor U9448 (N_9448,N_6429,N_7269);
nand U9449 (N_9449,N_6501,N_6728);
nor U9450 (N_9450,N_6277,N_6743);
or U9451 (N_9451,N_6977,N_6321);
or U9452 (N_9452,N_6251,N_6344);
or U9453 (N_9453,N_7531,N_7884);
nand U9454 (N_9454,N_6824,N_6176);
and U9455 (N_9455,N_7618,N_6194);
nand U9456 (N_9456,N_6334,N_6425);
nand U9457 (N_9457,N_7093,N_6915);
and U9458 (N_9458,N_6822,N_7880);
nand U9459 (N_9459,N_6051,N_7704);
nand U9460 (N_9460,N_6828,N_6120);
nor U9461 (N_9461,N_6523,N_7052);
and U9462 (N_9462,N_7925,N_6249);
or U9463 (N_9463,N_7121,N_7622);
and U9464 (N_9464,N_6526,N_6123);
nand U9465 (N_9465,N_6287,N_6929);
nor U9466 (N_9466,N_7726,N_6968);
nor U9467 (N_9467,N_6879,N_6823);
nand U9468 (N_9468,N_6719,N_6055);
or U9469 (N_9469,N_7963,N_6392);
nand U9470 (N_9470,N_7057,N_7159);
or U9471 (N_9471,N_6198,N_6031);
nor U9472 (N_9472,N_6814,N_7105);
or U9473 (N_9473,N_7458,N_6389);
nor U9474 (N_9474,N_7143,N_7782);
nor U9475 (N_9475,N_6572,N_6247);
nor U9476 (N_9476,N_7564,N_6521);
nand U9477 (N_9477,N_6542,N_6295);
or U9478 (N_9478,N_7767,N_6533);
xnor U9479 (N_9479,N_6449,N_7267);
nor U9480 (N_9480,N_6185,N_7144);
xor U9481 (N_9481,N_7508,N_6300);
nor U9482 (N_9482,N_7568,N_7519);
nor U9483 (N_9483,N_7402,N_6972);
nor U9484 (N_9484,N_7832,N_7301);
and U9485 (N_9485,N_7927,N_6958);
nand U9486 (N_9486,N_7624,N_6625);
nand U9487 (N_9487,N_6970,N_6088);
nor U9488 (N_9488,N_6125,N_6776);
nand U9489 (N_9489,N_7230,N_6247);
or U9490 (N_9490,N_7071,N_6158);
and U9491 (N_9491,N_6964,N_7001);
nand U9492 (N_9492,N_7615,N_6891);
nand U9493 (N_9493,N_7683,N_6486);
nor U9494 (N_9494,N_6350,N_7978);
or U9495 (N_9495,N_7447,N_7453);
nand U9496 (N_9496,N_7071,N_6329);
nand U9497 (N_9497,N_6356,N_7207);
or U9498 (N_9498,N_6604,N_7542);
and U9499 (N_9499,N_6161,N_7292);
and U9500 (N_9500,N_6655,N_6326);
and U9501 (N_9501,N_6247,N_6364);
nand U9502 (N_9502,N_7625,N_7584);
and U9503 (N_9503,N_6000,N_6511);
and U9504 (N_9504,N_7040,N_7813);
nor U9505 (N_9505,N_7271,N_7552);
nand U9506 (N_9506,N_7501,N_6131);
nand U9507 (N_9507,N_6546,N_7254);
nand U9508 (N_9508,N_6935,N_6666);
and U9509 (N_9509,N_6720,N_7202);
xor U9510 (N_9510,N_7435,N_7021);
nand U9511 (N_9511,N_6025,N_7526);
nand U9512 (N_9512,N_7930,N_6850);
nand U9513 (N_9513,N_6163,N_6415);
nor U9514 (N_9514,N_7352,N_6972);
or U9515 (N_9515,N_6346,N_6216);
nand U9516 (N_9516,N_6626,N_7564);
and U9517 (N_9517,N_6016,N_7708);
nor U9518 (N_9518,N_7651,N_7824);
nand U9519 (N_9519,N_7140,N_7399);
and U9520 (N_9520,N_7340,N_6351);
nand U9521 (N_9521,N_7133,N_7773);
and U9522 (N_9522,N_7760,N_6494);
nor U9523 (N_9523,N_7232,N_7553);
nand U9524 (N_9524,N_6772,N_6705);
or U9525 (N_9525,N_7356,N_7107);
or U9526 (N_9526,N_6336,N_7054);
or U9527 (N_9527,N_7563,N_6689);
and U9528 (N_9528,N_6341,N_6651);
nand U9529 (N_9529,N_6386,N_6738);
or U9530 (N_9530,N_7772,N_7142);
nand U9531 (N_9531,N_6058,N_6540);
nor U9532 (N_9532,N_6997,N_7963);
and U9533 (N_9533,N_7809,N_7666);
or U9534 (N_9534,N_7113,N_6546);
or U9535 (N_9535,N_7023,N_7405);
and U9536 (N_9536,N_7600,N_7631);
or U9537 (N_9537,N_7077,N_6855);
and U9538 (N_9538,N_7270,N_7229);
and U9539 (N_9539,N_7218,N_7752);
and U9540 (N_9540,N_7928,N_6594);
nor U9541 (N_9541,N_7545,N_6616);
nor U9542 (N_9542,N_6370,N_7148);
and U9543 (N_9543,N_7746,N_6516);
and U9544 (N_9544,N_6654,N_6678);
or U9545 (N_9545,N_6242,N_7718);
or U9546 (N_9546,N_6313,N_7669);
nand U9547 (N_9547,N_6427,N_7724);
nor U9548 (N_9548,N_6879,N_7542);
nor U9549 (N_9549,N_6705,N_7627);
and U9550 (N_9550,N_7148,N_7699);
nor U9551 (N_9551,N_6954,N_7343);
nand U9552 (N_9552,N_7068,N_7392);
nand U9553 (N_9553,N_6920,N_7945);
nand U9554 (N_9554,N_6485,N_7476);
or U9555 (N_9555,N_6307,N_7716);
or U9556 (N_9556,N_6548,N_6526);
or U9557 (N_9557,N_7826,N_7513);
and U9558 (N_9558,N_6013,N_7519);
nand U9559 (N_9559,N_6542,N_7144);
nand U9560 (N_9560,N_7713,N_7117);
or U9561 (N_9561,N_6347,N_6301);
and U9562 (N_9562,N_7677,N_7588);
or U9563 (N_9563,N_7260,N_6004);
nor U9564 (N_9564,N_6757,N_7125);
nand U9565 (N_9565,N_6482,N_7576);
nor U9566 (N_9566,N_7630,N_6860);
nand U9567 (N_9567,N_6145,N_7977);
and U9568 (N_9568,N_6489,N_7497);
and U9569 (N_9569,N_7579,N_7639);
nand U9570 (N_9570,N_7471,N_7665);
and U9571 (N_9571,N_6403,N_7933);
nor U9572 (N_9572,N_7416,N_6767);
and U9573 (N_9573,N_7108,N_6545);
and U9574 (N_9574,N_7640,N_6270);
or U9575 (N_9575,N_6505,N_6891);
nor U9576 (N_9576,N_7640,N_7774);
nor U9577 (N_9577,N_7628,N_7935);
nand U9578 (N_9578,N_6909,N_6371);
and U9579 (N_9579,N_7892,N_6847);
nor U9580 (N_9580,N_7163,N_6420);
and U9581 (N_9581,N_6911,N_6517);
or U9582 (N_9582,N_7017,N_6858);
and U9583 (N_9583,N_6851,N_7657);
nand U9584 (N_9584,N_7582,N_6172);
and U9585 (N_9585,N_6748,N_7579);
nand U9586 (N_9586,N_6057,N_6510);
or U9587 (N_9587,N_6642,N_7829);
nor U9588 (N_9588,N_6742,N_7283);
nand U9589 (N_9589,N_7448,N_6802);
nor U9590 (N_9590,N_6230,N_6922);
and U9591 (N_9591,N_6930,N_6899);
nor U9592 (N_9592,N_6222,N_6566);
or U9593 (N_9593,N_6861,N_6057);
nor U9594 (N_9594,N_7214,N_6604);
nor U9595 (N_9595,N_7569,N_6465);
nand U9596 (N_9596,N_7678,N_6384);
nand U9597 (N_9597,N_7409,N_7594);
nand U9598 (N_9598,N_6809,N_7889);
nor U9599 (N_9599,N_7155,N_7162);
nand U9600 (N_9600,N_6638,N_6519);
and U9601 (N_9601,N_6855,N_6366);
and U9602 (N_9602,N_7784,N_6880);
nand U9603 (N_9603,N_6475,N_6474);
and U9604 (N_9604,N_6708,N_6510);
or U9605 (N_9605,N_6461,N_7403);
nand U9606 (N_9606,N_6412,N_6758);
nand U9607 (N_9607,N_6960,N_6304);
nor U9608 (N_9608,N_7570,N_7728);
nor U9609 (N_9609,N_7212,N_7382);
or U9610 (N_9610,N_6328,N_7487);
and U9611 (N_9611,N_7124,N_7404);
and U9612 (N_9612,N_6322,N_6386);
or U9613 (N_9613,N_7999,N_7391);
nor U9614 (N_9614,N_7409,N_7345);
and U9615 (N_9615,N_7609,N_6712);
and U9616 (N_9616,N_7556,N_6684);
nand U9617 (N_9617,N_6567,N_7256);
and U9618 (N_9618,N_7033,N_6563);
nand U9619 (N_9619,N_7611,N_6459);
nand U9620 (N_9620,N_7022,N_6184);
or U9621 (N_9621,N_7331,N_7953);
and U9622 (N_9622,N_7951,N_7717);
and U9623 (N_9623,N_6555,N_6811);
or U9624 (N_9624,N_7945,N_6094);
nand U9625 (N_9625,N_7583,N_7026);
nand U9626 (N_9626,N_7658,N_7189);
and U9627 (N_9627,N_6282,N_7294);
xnor U9628 (N_9628,N_6933,N_7783);
nor U9629 (N_9629,N_6408,N_7942);
or U9630 (N_9630,N_6401,N_6942);
or U9631 (N_9631,N_6362,N_7736);
and U9632 (N_9632,N_7415,N_7178);
or U9633 (N_9633,N_6639,N_7766);
and U9634 (N_9634,N_6076,N_6989);
nor U9635 (N_9635,N_6618,N_7663);
and U9636 (N_9636,N_6371,N_7029);
and U9637 (N_9637,N_7040,N_7954);
and U9638 (N_9638,N_6689,N_7628);
nand U9639 (N_9639,N_6383,N_6863);
or U9640 (N_9640,N_7926,N_6368);
and U9641 (N_9641,N_6364,N_6842);
nand U9642 (N_9642,N_6365,N_7463);
nand U9643 (N_9643,N_6725,N_7811);
nand U9644 (N_9644,N_6315,N_6963);
nand U9645 (N_9645,N_6075,N_6755);
nor U9646 (N_9646,N_7994,N_6397);
nor U9647 (N_9647,N_7138,N_6322);
and U9648 (N_9648,N_7718,N_7532);
nor U9649 (N_9649,N_6883,N_6410);
and U9650 (N_9650,N_7926,N_6462);
nand U9651 (N_9651,N_7757,N_7439);
nand U9652 (N_9652,N_7279,N_7996);
nand U9653 (N_9653,N_6721,N_6368);
nor U9654 (N_9654,N_6425,N_6785);
or U9655 (N_9655,N_7293,N_7539);
and U9656 (N_9656,N_7520,N_7392);
and U9657 (N_9657,N_6587,N_7355);
and U9658 (N_9658,N_6688,N_7135);
nor U9659 (N_9659,N_7464,N_6697);
and U9660 (N_9660,N_7773,N_7073);
and U9661 (N_9661,N_6897,N_6282);
nor U9662 (N_9662,N_7944,N_6157);
nand U9663 (N_9663,N_7412,N_7945);
nor U9664 (N_9664,N_7871,N_6743);
nand U9665 (N_9665,N_7561,N_6551);
nor U9666 (N_9666,N_7468,N_6694);
nor U9667 (N_9667,N_7343,N_7124);
and U9668 (N_9668,N_6873,N_6108);
nand U9669 (N_9669,N_7413,N_6068);
and U9670 (N_9670,N_7942,N_6314);
and U9671 (N_9671,N_6286,N_7582);
or U9672 (N_9672,N_7879,N_7584);
nand U9673 (N_9673,N_6022,N_6497);
nor U9674 (N_9674,N_6883,N_7752);
nor U9675 (N_9675,N_6677,N_7579);
or U9676 (N_9676,N_7765,N_6778);
nand U9677 (N_9677,N_6779,N_6204);
nor U9678 (N_9678,N_6934,N_6160);
nand U9679 (N_9679,N_6745,N_6521);
or U9680 (N_9680,N_6143,N_7251);
nor U9681 (N_9681,N_7320,N_6032);
or U9682 (N_9682,N_7690,N_6037);
nor U9683 (N_9683,N_7350,N_7558);
or U9684 (N_9684,N_6222,N_6640);
nand U9685 (N_9685,N_6161,N_7975);
or U9686 (N_9686,N_7724,N_7518);
nand U9687 (N_9687,N_7729,N_7477);
nand U9688 (N_9688,N_7214,N_7713);
and U9689 (N_9689,N_6499,N_6288);
and U9690 (N_9690,N_6868,N_6904);
nand U9691 (N_9691,N_7907,N_6336);
nor U9692 (N_9692,N_7960,N_7610);
and U9693 (N_9693,N_6578,N_6506);
and U9694 (N_9694,N_6836,N_6018);
nor U9695 (N_9695,N_7458,N_6142);
and U9696 (N_9696,N_6503,N_7166);
nor U9697 (N_9697,N_7190,N_7395);
nand U9698 (N_9698,N_7313,N_7782);
or U9699 (N_9699,N_6912,N_6165);
or U9700 (N_9700,N_6926,N_7798);
or U9701 (N_9701,N_7417,N_7798);
or U9702 (N_9702,N_7570,N_7737);
nor U9703 (N_9703,N_6158,N_7162);
or U9704 (N_9704,N_7704,N_7899);
nand U9705 (N_9705,N_7037,N_7913);
and U9706 (N_9706,N_6351,N_6175);
or U9707 (N_9707,N_6009,N_6296);
nand U9708 (N_9708,N_6574,N_7354);
and U9709 (N_9709,N_7219,N_6648);
or U9710 (N_9710,N_7413,N_6412);
and U9711 (N_9711,N_6013,N_7646);
nor U9712 (N_9712,N_6324,N_6815);
nand U9713 (N_9713,N_6833,N_6916);
nor U9714 (N_9714,N_6078,N_7868);
nor U9715 (N_9715,N_6475,N_7927);
or U9716 (N_9716,N_6201,N_6594);
and U9717 (N_9717,N_7536,N_7621);
nand U9718 (N_9718,N_7862,N_6545);
nand U9719 (N_9719,N_7782,N_6785);
and U9720 (N_9720,N_7776,N_7134);
or U9721 (N_9721,N_6028,N_6526);
and U9722 (N_9722,N_6165,N_6155);
or U9723 (N_9723,N_7164,N_6552);
or U9724 (N_9724,N_6098,N_7602);
nor U9725 (N_9725,N_7043,N_7317);
nor U9726 (N_9726,N_6901,N_7244);
and U9727 (N_9727,N_6482,N_7133);
nand U9728 (N_9728,N_6856,N_6142);
nand U9729 (N_9729,N_7731,N_6456);
nand U9730 (N_9730,N_7053,N_7167);
or U9731 (N_9731,N_7439,N_7993);
and U9732 (N_9732,N_6021,N_6823);
nand U9733 (N_9733,N_6284,N_7342);
nand U9734 (N_9734,N_7008,N_6846);
and U9735 (N_9735,N_6490,N_6400);
nand U9736 (N_9736,N_6670,N_7635);
nand U9737 (N_9737,N_7832,N_6496);
and U9738 (N_9738,N_7914,N_6919);
nand U9739 (N_9739,N_7198,N_6986);
nand U9740 (N_9740,N_6753,N_6996);
nand U9741 (N_9741,N_7789,N_6358);
nand U9742 (N_9742,N_6598,N_7333);
and U9743 (N_9743,N_7408,N_6871);
nor U9744 (N_9744,N_7249,N_7276);
nand U9745 (N_9745,N_7423,N_7819);
and U9746 (N_9746,N_7241,N_6094);
nor U9747 (N_9747,N_6074,N_7274);
or U9748 (N_9748,N_7120,N_7881);
and U9749 (N_9749,N_7629,N_6644);
nor U9750 (N_9750,N_7354,N_7018);
nand U9751 (N_9751,N_7080,N_7688);
and U9752 (N_9752,N_6214,N_7707);
or U9753 (N_9753,N_6409,N_6305);
or U9754 (N_9754,N_6931,N_7353);
and U9755 (N_9755,N_6472,N_7553);
nor U9756 (N_9756,N_7482,N_6791);
nor U9757 (N_9757,N_7717,N_6773);
or U9758 (N_9758,N_7751,N_7789);
and U9759 (N_9759,N_7357,N_7976);
nor U9760 (N_9760,N_7703,N_6171);
nor U9761 (N_9761,N_7105,N_6079);
nand U9762 (N_9762,N_7088,N_6209);
nor U9763 (N_9763,N_6002,N_7325);
nor U9764 (N_9764,N_7036,N_6912);
nor U9765 (N_9765,N_7648,N_7790);
and U9766 (N_9766,N_7191,N_6183);
nand U9767 (N_9767,N_7221,N_6201);
or U9768 (N_9768,N_6196,N_7551);
and U9769 (N_9769,N_6040,N_6456);
nand U9770 (N_9770,N_6110,N_6703);
or U9771 (N_9771,N_7085,N_7715);
nand U9772 (N_9772,N_7819,N_6330);
and U9773 (N_9773,N_7066,N_7951);
or U9774 (N_9774,N_7274,N_7757);
or U9775 (N_9775,N_6552,N_7982);
nor U9776 (N_9776,N_6037,N_7080);
or U9777 (N_9777,N_6297,N_6153);
and U9778 (N_9778,N_6185,N_6372);
nand U9779 (N_9779,N_6566,N_6362);
nand U9780 (N_9780,N_7259,N_7243);
nor U9781 (N_9781,N_6867,N_7896);
and U9782 (N_9782,N_7116,N_6266);
nand U9783 (N_9783,N_6407,N_6468);
or U9784 (N_9784,N_7782,N_7322);
or U9785 (N_9785,N_7593,N_6739);
or U9786 (N_9786,N_7374,N_6654);
or U9787 (N_9787,N_6178,N_6877);
and U9788 (N_9788,N_7837,N_6712);
nand U9789 (N_9789,N_7902,N_7770);
nor U9790 (N_9790,N_7405,N_7524);
nor U9791 (N_9791,N_7320,N_7874);
or U9792 (N_9792,N_7858,N_7294);
and U9793 (N_9793,N_7744,N_7836);
nand U9794 (N_9794,N_7679,N_6198);
or U9795 (N_9795,N_6812,N_6071);
or U9796 (N_9796,N_7885,N_6736);
nor U9797 (N_9797,N_7019,N_7049);
and U9798 (N_9798,N_6876,N_6304);
nand U9799 (N_9799,N_7427,N_7850);
and U9800 (N_9800,N_6314,N_6822);
or U9801 (N_9801,N_7025,N_6623);
and U9802 (N_9802,N_6558,N_7874);
and U9803 (N_9803,N_6822,N_7437);
xor U9804 (N_9804,N_7799,N_6181);
nor U9805 (N_9805,N_7534,N_6896);
or U9806 (N_9806,N_6974,N_6957);
nor U9807 (N_9807,N_6997,N_7413);
and U9808 (N_9808,N_7563,N_7583);
nor U9809 (N_9809,N_6958,N_6810);
nand U9810 (N_9810,N_7390,N_6711);
and U9811 (N_9811,N_6140,N_6757);
and U9812 (N_9812,N_6667,N_6069);
nand U9813 (N_9813,N_7856,N_6444);
or U9814 (N_9814,N_6800,N_7532);
nor U9815 (N_9815,N_6976,N_6821);
and U9816 (N_9816,N_7675,N_6631);
nor U9817 (N_9817,N_7417,N_7586);
nor U9818 (N_9818,N_6570,N_7872);
and U9819 (N_9819,N_6552,N_7672);
or U9820 (N_9820,N_6623,N_6442);
or U9821 (N_9821,N_7202,N_7920);
nand U9822 (N_9822,N_7422,N_6255);
nor U9823 (N_9823,N_7112,N_6016);
or U9824 (N_9824,N_6827,N_6053);
nand U9825 (N_9825,N_6265,N_7249);
or U9826 (N_9826,N_6196,N_6844);
nand U9827 (N_9827,N_6958,N_6899);
or U9828 (N_9828,N_6649,N_7871);
nand U9829 (N_9829,N_6705,N_7096);
or U9830 (N_9830,N_6792,N_7757);
nand U9831 (N_9831,N_7030,N_6795);
nand U9832 (N_9832,N_6395,N_6630);
nor U9833 (N_9833,N_7599,N_7904);
and U9834 (N_9834,N_6408,N_7296);
or U9835 (N_9835,N_7971,N_6854);
nor U9836 (N_9836,N_6816,N_7519);
and U9837 (N_9837,N_7903,N_7307);
and U9838 (N_9838,N_7844,N_6429);
and U9839 (N_9839,N_6102,N_7892);
and U9840 (N_9840,N_7926,N_6745);
nand U9841 (N_9841,N_6994,N_6279);
nand U9842 (N_9842,N_7476,N_7221);
and U9843 (N_9843,N_7873,N_7005);
or U9844 (N_9844,N_7838,N_6054);
xnor U9845 (N_9845,N_6373,N_7628);
or U9846 (N_9846,N_6437,N_7925);
nand U9847 (N_9847,N_6624,N_6019);
nand U9848 (N_9848,N_6721,N_6554);
nand U9849 (N_9849,N_6946,N_6794);
nor U9850 (N_9850,N_6452,N_7803);
or U9851 (N_9851,N_6401,N_6887);
and U9852 (N_9852,N_6497,N_6611);
or U9853 (N_9853,N_6580,N_7294);
or U9854 (N_9854,N_6167,N_7932);
or U9855 (N_9855,N_6396,N_7648);
and U9856 (N_9856,N_6353,N_7297);
nand U9857 (N_9857,N_7390,N_7252);
or U9858 (N_9858,N_7731,N_7616);
and U9859 (N_9859,N_7100,N_7434);
or U9860 (N_9860,N_6453,N_7164);
nor U9861 (N_9861,N_6943,N_6244);
and U9862 (N_9862,N_7865,N_7553);
and U9863 (N_9863,N_7858,N_7769);
nor U9864 (N_9864,N_6421,N_6460);
or U9865 (N_9865,N_7766,N_7915);
nor U9866 (N_9866,N_6092,N_7546);
nand U9867 (N_9867,N_6857,N_7317);
or U9868 (N_9868,N_7625,N_6650);
or U9869 (N_9869,N_7300,N_7304);
nor U9870 (N_9870,N_7681,N_6184);
nand U9871 (N_9871,N_7885,N_6041);
and U9872 (N_9872,N_7650,N_7900);
nand U9873 (N_9873,N_7744,N_6579);
and U9874 (N_9874,N_6595,N_6979);
nand U9875 (N_9875,N_7496,N_6683);
and U9876 (N_9876,N_6635,N_6102);
nand U9877 (N_9877,N_6197,N_6163);
and U9878 (N_9878,N_7025,N_7290);
nor U9879 (N_9879,N_7874,N_7281);
or U9880 (N_9880,N_6322,N_6716);
nand U9881 (N_9881,N_6273,N_7572);
or U9882 (N_9882,N_6804,N_7646);
and U9883 (N_9883,N_6742,N_6060);
and U9884 (N_9884,N_7095,N_7380);
and U9885 (N_9885,N_6012,N_7427);
nand U9886 (N_9886,N_6863,N_6600);
xnor U9887 (N_9887,N_6519,N_6670);
and U9888 (N_9888,N_7910,N_7070);
nand U9889 (N_9889,N_7079,N_7328);
xor U9890 (N_9890,N_7562,N_6817);
nand U9891 (N_9891,N_7374,N_7410);
nand U9892 (N_9892,N_7959,N_6892);
nor U9893 (N_9893,N_6947,N_6138);
xor U9894 (N_9894,N_7048,N_6979);
or U9895 (N_9895,N_6870,N_6828);
or U9896 (N_9896,N_7609,N_6866);
nand U9897 (N_9897,N_6114,N_7054);
nor U9898 (N_9898,N_6114,N_7184);
and U9899 (N_9899,N_6557,N_7561);
or U9900 (N_9900,N_7624,N_7342);
and U9901 (N_9901,N_7478,N_7546);
and U9902 (N_9902,N_6755,N_7413);
nand U9903 (N_9903,N_7633,N_7169);
and U9904 (N_9904,N_6354,N_6098);
and U9905 (N_9905,N_7375,N_6419);
or U9906 (N_9906,N_6035,N_6323);
or U9907 (N_9907,N_6873,N_7921);
nand U9908 (N_9908,N_7531,N_6231);
nor U9909 (N_9909,N_6432,N_7451);
and U9910 (N_9910,N_6322,N_6478);
or U9911 (N_9911,N_7305,N_6639);
nand U9912 (N_9912,N_7218,N_7410);
nor U9913 (N_9913,N_7868,N_7458);
and U9914 (N_9914,N_6331,N_7591);
nor U9915 (N_9915,N_6074,N_7081);
nor U9916 (N_9916,N_6393,N_6308);
or U9917 (N_9917,N_7637,N_7373);
nor U9918 (N_9918,N_6714,N_7190);
or U9919 (N_9919,N_7119,N_7020);
or U9920 (N_9920,N_7577,N_6424);
and U9921 (N_9921,N_6738,N_6842);
nor U9922 (N_9922,N_6656,N_7578);
nor U9923 (N_9923,N_6020,N_7001);
nor U9924 (N_9924,N_7447,N_6653);
and U9925 (N_9925,N_7402,N_6351);
or U9926 (N_9926,N_6963,N_6078);
or U9927 (N_9927,N_7580,N_6690);
nor U9928 (N_9928,N_7560,N_6821);
and U9929 (N_9929,N_7802,N_7151);
and U9930 (N_9930,N_6903,N_6179);
or U9931 (N_9931,N_7654,N_6550);
or U9932 (N_9932,N_7848,N_6258);
nor U9933 (N_9933,N_7331,N_7654);
and U9934 (N_9934,N_7570,N_7323);
or U9935 (N_9935,N_7205,N_7860);
and U9936 (N_9936,N_7087,N_7886);
or U9937 (N_9937,N_7798,N_6986);
or U9938 (N_9938,N_7644,N_6847);
nand U9939 (N_9939,N_6150,N_7456);
nand U9940 (N_9940,N_6737,N_6671);
and U9941 (N_9941,N_6563,N_7668);
and U9942 (N_9942,N_6795,N_7881);
and U9943 (N_9943,N_6303,N_6259);
or U9944 (N_9944,N_6000,N_7155);
nor U9945 (N_9945,N_6685,N_6607);
nand U9946 (N_9946,N_6405,N_6719);
and U9947 (N_9947,N_6218,N_6591);
nand U9948 (N_9948,N_7618,N_6306);
and U9949 (N_9949,N_6696,N_6295);
nand U9950 (N_9950,N_7321,N_7173);
nor U9951 (N_9951,N_7865,N_6250);
or U9952 (N_9952,N_6127,N_7471);
nor U9953 (N_9953,N_7904,N_6950);
and U9954 (N_9954,N_6454,N_7114);
nor U9955 (N_9955,N_7876,N_7235);
nor U9956 (N_9956,N_6769,N_7388);
nand U9957 (N_9957,N_6731,N_6184);
and U9958 (N_9958,N_6301,N_6036);
and U9959 (N_9959,N_7660,N_7041);
nor U9960 (N_9960,N_6298,N_7230);
nor U9961 (N_9961,N_6111,N_6302);
or U9962 (N_9962,N_7437,N_7891);
nand U9963 (N_9963,N_7450,N_6849);
and U9964 (N_9964,N_7938,N_7820);
xor U9965 (N_9965,N_7885,N_7592);
nor U9966 (N_9966,N_7637,N_6097);
xnor U9967 (N_9967,N_6659,N_6928);
and U9968 (N_9968,N_7793,N_6906);
and U9969 (N_9969,N_6532,N_7763);
nand U9970 (N_9970,N_7605,N_6740);
and U9971 (N_9971,N_6810,N_7356);
and U9972 (N_9972,N_7496,N_6817);
nand U9973 (N_9973,N_7540,N_6727);
nand U9974 (N_9974,N_7192,N_6313);
nor U9975 (N_9975,N_7112,N_7782);
nor U9976 (N_9976,N_7257,N_6366);
or U9977 (N_9977,N_7883,N_6568);
nand U9978 (N_9978,N_6744,N_6601);
or U9979 (N_9979,N_7730,N_7281);
and U9980 (N_9980,N_7577,N_7193);
and U9981 (N_9981,N_7673,N_7362);
nor U9982 (N_9982,N_7087,N_6905);
and U9983 (N_9983,N_6283,N_7681);
nor U9984 (N_9984,N_6200,N_6529);
nand U9985 (N_9985,N_7592,N_6992);
nor U9986 (N_9986,N_6948,N_6438);
or U9987 (N_9987,N_6307,N_6222);
or U9988 (N_9988,N_7412,N_7313);
and U9989 (N_9989,N_7762,N_6143);
or U9990 (N_9990,N_7570,N_6083);
nand U9991 (N_9991,N_6943,N_6991);
nor U9992 (N_9992,N_7368,N_7480);
nor U9993 (N_9993,N_6529,N_6017);
nor U9994 (N_9994,N_7557,N_7629);
and U9995 (N_9995,N_6704,N_6004);
or U9996 (N_9996,N_7229,N_6961);
nand U9997 (N_9997,N_7853,N_6950);
nor U9998 (N_9998,N_6814,N_6681);
or U9999 (N_9999,N_6482,N_6955);
or UO_0 (O_0,N_8635,N_8043);
nor UO_1 (O_1,N_8880,N_8817);
nor UO_2 (O_2,N_8244,N_9513);
and UO_3 (O_3,N_8514,N_8254);
nand UO_4 (O_4,N_8386,N_8944);
or UO_5 (O_5,N_8310,N_8031);
nor UO_6 (O_6,N_9303,N_9692);
nor UO_7 (O_7,N_8882,N_8594);
or UO_8 (O_8,N_9994,N_8166);
and UO_9 (O_9,N_9419,N_8577);
xnor UO_10 (O_10,N_8107,N_9267);
and UO_11 (O_11,N_8558,N_8400);
or UO_12 (O_12,N_8858,N_9298);
nor UO_13 (O_13,N_8103,N_9817);
nor UO_14 (O_14,N_8768,N_8266);
nand UO_15 (O_15,N_8194,N_8988);
or UO_16 (O_16,N_8681,N_8280);
nor UO_17 (O_17,N_8460,N_8814);
and UO_18 (O_18,N_8971,N_8949);
or UO_19 (O_19,N_9159,N_9234);
or UO_20 (O_20,N_8890,N_9903);
nand UO_21 (O_21,N_8838,N_9579);
and UO_22 (O_22,N_9696,N_9237);
or UO_23 (O_23,N_8936,N_9001);
or UO_24 (O_24,N_8193,N_8160);
and UO_25 (O_25,N_9408,N_8220);
nor UO_26 (O_26,N_8791,N_9388);
nand UO_27 (O_27,N_9431,N_9614);
and UO_28 (O_28,N_8520,N_8128);
or UO_29 (O_29,N_9951,N_9199);
and UO_30 (O_30,N_9185,N_8983);
nand UO_31 (O_31,N_8684,N_8109);
nand UO_32 (O_32,N_8172,N_9908);
or UO_33 (O_33,N_8579,N_9942);
and UO_34 (O_34,N_8546,N_8354);
and UO_35 (O_35,N_9631,N_9134);
nor UO_36 (O_36,N_8132,N_9675);
and UO_37 (O_37,N_9057,N_9931);
or UO_38 (O_38,N_9041,N_8037);
nand UO_39 (O_39,N_8207,N_8086);
nand UO_40 (O_40,N_9430,N_8426);
nor UO_41 (O_41,N_8085,N_9182);
and UO_42 (O_42,N_9799,N_8126);
and UO_43 (O_43,N_8344,N_8063);
nor UO_44 (O_44,N_8407,N_9027);
nand UO_45 (O_45,N_9088,N_9280);
or UO_46 (O_46,N_8715,N_8932);
nand UO_47 (O_47,N_9583,N_9060);
nor UO_48 (O_48,N_8591,N_8134);
nand UO_49 (O_49,N_8404,N_8600);
and UO_50 (O_50,N_9301,N_9665);
nand UO_51 (O_51,N_9380,N_9978);
nor UO_52 (O_52,N_9873,N_8551);
nor UO_53 (O_53,N_8722,N_9745);
nor UO_54 (O_54,N_8141,N_9012);
or UO_55 (O_55,N_8054,N_9445);
nor UO_56 (O_56,N_8078,N_9868);
nand UO_57 (O_57,N_8067,N_8652);
nand UO_58 (O_58,N_8784,N_8545);
and UO_59 (O_59,N_9619,N_9819);
nor UO_60 (O_60,N_8281,N_9544);
nand UO_61 (O_61,N_9098,N_8330);
and UO_62 (O_62,N_8848,N_8780);
or UO_63 (O_63,N_8883,N_8997);
xnor UO_64 (O_64,N_9054,N_9527);
nand UO_65 (O_65,N_9487,N_8159);
or UO_66 (O_66,N_9018,N_9421);
and UO_67 (O_67,N_8110,N_8902);
or UO_68 (O_68,N_8973,N_8495);
nor UO_69 (O_69,N_8030,N_8154);
or UO_70 (O_70,N_8359,N_8236);
nor UO_71 (O_71,N_9105,N_8197);
and UO_72 (O_72,N_8967,N_9106);
nand UO_73 (O_73,N_9037,N_8291);
xnor UO_74 (O_74,N_8010,N_9078);
and UO_75 (O_75,N_8089,N_8341);
nor UO_76 (O_76,N_8405,N_8060);
nand UO_77 (O_77,N_8148,N_8438);
or UO_78 (O_78,N_9166,N_9202);
nand UO_79 (O_79,N_8124,N_9714);
and UO_80 (O_80,N_9687,N_8852);
nor UO_81 (O_81,N_9092,N_8501);
nand UO_82 (O_82,N_8621,N_9257);
nand UO_83 (O_83,N_9443,N_8705);
and UO_84 (O_84,N_8284,N_8928);
or UO_85 (O_85,N_8497,N_8674);
nor UO_86 (O_86,N_9005,N_8756);
nand UO_87 (O_87,N_9118,N_8427);
and UO_88 (O_88,N_8216,N_8387);
nand UO_89 (O_89,N_9703,N_8217);
nor UO_90 (O_90,N_8362,N_8155);
nand UO_91 (O_91,N_9925,N_9640);
nor UO_92 (O_92,N_9140,N_8805);
nor UO_93 (O_93,N_9712,N_8927);
xnor UO_94 (O_94,N_8275,N_9126);
and UO_95 (O_95,N_8508,N_8845);
nand UO_96 (O_96,N_9417,N_9693);
nor UO_97 (O_97,N_9839,N_9859);
nand UO_98 (O_98,N_9764,N_9706);
nor UO_99 (O_99,N_8071,N_9558);
nor UO_100 (O_100,N_9890,N_8419);
nor UO_101 (O_101,N_8531,N_9580);
nor UO_102 (O_102,N_8680,N_8799);
nor UO_103 (O_103,N_8486,N_9788);
and UO_104 (O_104,N_9676,N_8099);
or UO_105 (O_105,N_9644,N_8733);
nand UO_106 (O_106,N_9128,N_8249);
nor UO_107 (O_107,N_9715,N_8543);
and UO_108 (O_108,N_8530,N_9882);
nand UO_109 (O_109,N_9958,N_9353);
and UO_110 (O_110,N_8907,N_8730);
or UO_111 (O_111,N_8425,N_8646);
nor UO_112 (O_112,N_8802,N_9108);
and UO_113 (O_113,N_9989,N_9173);
xnor UO_114 (O_114,N_9139,N_9974);
or UO_115 (O_115,N_8662,N_9113);
and UO_116 (O_116,N_9773,N_9137);
nor UO_117 (O_117,N_9387,N_8410);
or UO_118 (O_118,N_9986,N_8296);
nor UO_119 (O_119,N_8349,N_9291);
nor UO_120 (O_120,N_8849,N_8627);
and UO_121 (O_121,N_8668,N_9322);
nor UO_122 (O_122,N_8653,N_8533);
or UO_123 (O_123,N_9339,N_9800);
nor UO_124 (O_124,N_9996,N_8637);
and UO_125 (O_125,N_8252,N_9411);
nand UO_126 (O_126,N_8396,N_9273);
or UO_127 (O_127,N_9645,N_9241);
and UO_128 (O_128,N_8956,N_9500);
nor UO_129 (O_129,N_9014,N_9300);
nor UO_130 (O_130,N_9420,N_9984);
nor UO_131 (O_131,N_8998,N_8070);
and UO_132 (O_132,N_9959,N_8716);
or UO_133 (O_133,N_9452,N_8611);
nand UO_134 (O_134,N_8383,N_8300);
nor UO_135 (O_135,N_8005,N_8747);
nand UO_136 (O_136,N_9953,N_9683);
or UO_137 (O_137,N_9306,N_9590);
and UO_138 (O_138,N_9471,N_8444);
and UO_139 (O_139,N_8875,N_8554);
and UO_140 (O_140,N_9501,N_8262);
nor UO_141 (O_141,N_8263,N_8368);
nand UO_142 (O_142,N_9837,N_9827);
or UO_143 (O_143,N_8638,N_9874);
nand UO_144 (O_144,N_8959,N_8226);
nand UO_145 (O_145,N_9393,N_8632);
nor UO_146 (O_146,N_8834,N_9547);
and UO_147 (O_147,N_9283,N_8815);
nor UO_148 (O_148,N_9065,N_8755);
or UO_149 (O_149,N_8870,N_9962);
or UO_150 (O_150,N_9497,N_8829);
or UO_151 (O_151,N_8553,N_9285);
nor UO_152 (O_152,N_8536,N_9743);
and UO_153 (O_153,N_9632,N_9224);
and UO_154 (O_154,N_9063,N_9600);
and UO_155 (O_155,N_8761,N_8395);
xnor UO_156 (O_156,N_9153,N_9794);
or UO_157 (O_157,N_9004,N_9344);
nand UO_158 (O_158,N_9635,N_9177);
nand UO_159 (O_159,N_8463,N_8446);
or UO_160 (O_160,N_8881,N_8261);
and UO_161 (O_161,N_8930,N_8174);
and UO_162 (O_162,N_8806,N_8229);
nor UO_163 (O_163,N_8872,N_9574);
nand UO_164 (O_164,N_8417,N_8447);
nor UO_165 (O_165,N_8735,N_9945);
or UO_166 (O_166,N_8087,N_8313);
or UO_167 (O_167,N_9368,N_8714);
or UO_168 (O_168,N_9403,N_9294);
nand UO_169 (O_169,N_8992,N_9789);
nand UO_170 (O_170,N_8813,N_8625);
nand UO_171 (O_171,N_8596,N_9010);
nor UO_172 (O_172,N_9246,N_8038);
nor UO_173 (O_173,N_8707,N_9311);
and UO_174 (O_174,N_9372,N_8989);
nor UO_175 (O_175,N_8879,N_9730);
or UO_176 (O_176,N_9491,N_8575);
nor UO_177 (O_177,N_8511,N_8527);
and UO_178 (O_178,N_8887,N_8481);
and UO_179 (O_179,N_9049,N_8108);
and UO_180 (O_180,N_8299,N_9489);
or UO_181 (O_181,N_8462,N_8473);
and UO_182 (O_182,N_9402,N_9056);
and UO_183 (O_183,N_8754,N_8620);
and UO_184 (O_184,N_8050,N_9720);
or UO_185 (O_185,N_8414,N_9766);
or UO_186 (O_186,N_9238,N_8841);
nor UO_187 (O_187,N_9970,N_9840);
or UO_188 (O_188,N_8374,N_9820);
nand UO_189 (O_189,N_8686,N_9499);
nor UO_190 (O_190,N_8149,N_8176);
and UO_191 (O_191,N_8051,N_9206);
nor UO_192 (O_192,N_8699,N_8454);
or UO_193 (O_193,N_8540,N_8146);
or UO_194 (O_194,N_9308,N_8597);
and UO_195 (O_195,N_9522,N_9472);
nor UO_196 (O_196,N_9039,N_8476);
nand UO_197 (O_197,N_9170,N_8616);
nand UO_198 (O_198,N_8117,N_9757);
nor UO_199 (O_199,N_8270,N_9553);
nor UO_200 (O_200,N_9504,N_9198);
nor UO_201 (O_201,N_8539,N_8029);
nand UO_202 (O_202,N_9214,N_9381);
or UO_203 (O_203,N_9576,N_8151);
and UO_204 (O_204,N_8505,N_9662);
nor UO_205 (O_205,N_9284,N_9923);
and UO_206 (O_206,N_9647,N_9243);
nor UO_207 (O_207,N_9950,N_8757);
nand UO_208 (O_208,N_9832,N_8198);
and UO_209 (O_209,N_8810,N_9966);
nor UO_210 (O_210,N_9319,N_9130);
or UO_211 (O_211,N_8415,N_9998);
or UO_212 (O_212,N_9935,N_9733);
or UO_213 (O_213,N_9876,N_8092);
or UO_214 (O_214,N_9537,N_8190);
and UO_215 (O_215,N_9685,N_8339);
and UO_216 (O_216,N_9272,N_9969);
nand UO_217 (O_217,N_9230,N_9806);
nand UO_218 (O_218,N_9535,N_8235);
nand UO_219 (O_219,N_9560,N_9588);
and UO_220 (O_220,N_9849,N_8599);
nand UO_221 (O_221,N_9091,N_9550);
nor UO_222 (O_222,N_8905,N_8948);
or UO_223 (O_223,N_9968,N_9707);
and UO_224 (O_224,N_8456,N_8474);
and UO_225 (O_225,N_9768,N_9035);
nand UO_226 (O_226,N_8990,N_8855);
nand UO_227 (O_227,N_8184,N_8677);
nand UO_228 (O_228,N_9119,N_8604);
nor UO_229 (O_229,N_9315,N_8630);
nor UO_230 (O_230,N_9864,N_8801);
or UO_231 (O_231,N_8534,N_8378);
or UO_232 (O_232,N_9666,N_8706);
nand UO_233 (O_233,N_8480,N_9236);
xor UO_234 (O_234,N_9440,N_9967);
nand UO_235 (O_235,N_8869,N_9628);
or UO_236 (O_236,N_9601,N_8464);
and UO_237 (O_237,N_8946,N_8168);
nand UO_238 (O_238,N_9436,N_9963);
or UO_239 (O_239,N_9716,N_9607);
nor UO_240 (O_240,N_9674,N_8352);
and UO_241 (O_241,N_8366,N_9798);
nor UO_242 (O_242,N_9019,N_9593);
or UO_243 (O_243,N_9016,N_8676);
nand UO_244 (O_244,N_8049,N_9911);
or UO_245 (O_245,N_9256,N_9176);
nand UO_246 (O_246,N_9532,N_9150);
and UO_247 (O_247,N_8242,N_9762);
or UO_248 (O_248,N_9023,N_9909);
and UO_249 (O_249,N_8022,N_9248);
and UO_250 (O_250,N_9055,N_9835);
and UO_251 (O_251,N_9725,N_9634);
or UO_252 (O_252,N_9852,N_9934);
nor UO_253 (O_253,N_9076,N_9684);
and UO_254 (O_254,N_9331,N_8718);
nand UO_255 (O_255,N_9573,N_9053);
nor UO_256 (O_256,N_9981,N_9554);
nor UO_257 (O_257,N_9575,N_9099);
and UO_258 (O_258,N_8698,N_9680);
or UO_259 (O_259,N_8958,N_8429);
or UO_260 (O_260,N_9069,N_9287);
nor UO_261 (O_261,N_8322,N_8072);
nor UO_262 (O_262,N_8820,N_9651);
or UO_263 (O_263,N_8265,N_9888);
or UO_264 (O_264,N_8547,N_8642);
nor UO_265 (O_265,N_8697,N_8048);
nor UO_266 (O_266,N_9578,N_9071);
and UO_267 (O_267,N_9704,N_8938);
and UO_268 (O_268,N_8450,N_9744);
and UO_269 (O_269,N_8683,N_8276);
nand UO_270 (O_270,N_9083,N_8101);
nand UO_271 (O_271,N_9734,N_9043);
and UO_272 (O_272,N_8131,N_9323);
and UO_273 (O_273,N_8304,N_9261);
nand UO_274 (O_274,N_9228,N_8376);
and UO_275 (O_275,N_8873,N_9771);
nor UO_276 (O_276,N_9865,N_9000);
nand UO_277 (O_277,N_9829,N_9936);
nand UO_278 (O_278,N_9048,N_8835);
nand UO_279 (O_279,N_8259,N_9210);
and UO_280 (O_280,N_8201,N_8622);
nor UO_281 (O_281,N_9979,N_9484);
and UO_282 (O_282,N_9358,N_8326);
and UO_283 (O_283,N_8423,N_8177);
and UO_284 (O_284,N_8443,N_8708);
nand UO_285 (O_285,N_8748,N_9017);
and UO_286 (O_286,N_9450,N_8644);
and UO_287 (O_287,N_9678,N_9517);
or UO_288 (O_288,N_9094,N_9758);
nand UO_289 (O_289,N_8267,N_9493);
nand UO_290 (O_290,N_8685,N_9955);
nor UO_291 (O_291,N_9562,N_9671);
nand UO_292 (O_292,N_8673,N_9127);
and UO_293 (O_293,N_8321,N_9643);
nand UO_294 (O_294,N_8777,N_8325);
or UO_295 (O_295,N_8592,N_9154);
nor UO_296 (O_296,N_8451,N_9565);
nor UO_297 (O_297,N_9917,N_8129);
or UO_298 (O_298,N_9196,N_9548);
nor UO_299 (O_299,N_9586,N_8439);
or UO_300 (O_300,N_9342,N_8239);
nor UO_301 (O_301,N_9459,N_9110);
and UO_302 (O_302,N_9157,N_9982);
and UO_303 (O_303,N_9494,N_9349);
or UO_304 (O_304,N_9506,N_8731);
nand UO_305 (O_305,N_8739,N_8911);
and UO_306 (O_306,N_9031,N_9040);
or UO_307 (O_307,N_8765,N_9193);
nand UO_308 (O_308,N_9061,N_8889);
or UO_309 (O_309,N_8336,N_9528);
nor UO_310 (O_310,N_9307,N_9728);
and UO_311 (O_311,N_8482,N_8348);
and UO_312 (O_312,N_9933,N_9605);
and UO_313 (O_313,N_8379,N_9072);
nand UO_314 (O_314,N_9032,N_9414);
nand UO_315 (O_315,N_8179,N_8100);
xor UO_316 (O_316,N_9581,N_9977);
nor UO_317 (O_317,N_8337,N_8691);
or UO_318 (O_318,N_9983,N_9441);
nand UO_319 (O_319,N_8695,N_8792);
and UO_320 (O_320,N_8953,N_8182);
and UO_321 (O_321,N_8830,N_8413);
or UO_322 (O_322,N_8024,N_9229);
nor UO_323 (O_323,N_8526,N_9318);
or UO_324 (O_324,N_8812,N_9812);
nand UO_325 (O_325,N_9514,N_8323);
nand UO_326 (O_326,N_8068,N_9412);
nand UO_327 (O_327,N_9880,N_9121);
and UO_328 (O_328,N_8130,N_8016);
or UO_329 (O_329,N_8893,N_8178);
and UO_330 (O_330,N_8789,N_9188);
or UO_331 (O_331,N_9737,N_8862);
nand UO_332 (O_332,N_8183,N_8328);
nand UO_333 (O_333,N_9862,N_8571);
and UO_334 (O_334,N_9218,N_8549);
and UO_335 (O_335,N_9821,N_9021);
and UO_336 (O_336,N_9906,N_8181);
nand UO_337 (O_337,N_9512,N_8645);
and UO_338 (O_338,N_8351,N_9075);
or UO_339 (O_339,N_8639,N_9603);
and UO_340 (O_340,N_8257,N_8827);
and UO_341 (O_341,N_9391,N_9013);
or UO_342 (O_342,N_9332,N_8047);
nand UO_343 (O_343,N_8279,N_9980);
and UO_344 (O_344,N_8657,N_9952);
and UO_345 (O_345,N_9597,N_9699);
nor UO_346 (O_346,N_8350,N_9723);
nand UO_347 (O_347,N_8826,N_9426);
nor UO_348 (O_348,N_8225,N_8459);
or UO_349 (O_349,N_9965,N_9244);
nand UO_350 (O_350,N_8568,N_9329);
and UO_351 (O_351,N_9572,N_9729);
nand UO_352 (O_352,N_9203,N_9801);
or UO_353 (O_353,N_8742,N_8924);
and UO_354 (O_354,N_8065,N_8819);
or UO_355 (O_355,N_8665,N_8836);
and UO_356 (O_356,N_8567,N_9112);
nor UO_357 (O_357,N_9446,N_8980);
or UO_358 (O_358,N_8560,N_8271);
or UO_359 (O_359,N_9618,N_9582);
or UO_360 (O_360,N_9926,N_8795);
and UO_361 (O_361,N_9370,N_8609);
or UO_362 (O_362,N_8895,N_8669);
nor UO_363 (O_363,N_8661,N_9397);
nor UO_364 (O_364,N_8926,N_9305);
or UO_365 (O_365,N_8306,N_9468);
nand UO_366 (O_366,N_9405,N_8420);
nor UO_367 (O_367,N_9813,N_8475);
and UO_368 (O_368,N_9330,N_8741);
and UO_369 (O_369,N_9668,N_9138);
nor UO_370 (O_370,N_8012,N_9416);
or UO_371 (O_371,N_8021,N_8861);
nand UO_372 (O_372,N_8593,N_8878);
nor UO_373 (O_373,N_9422,N_9557);
nor UO_374 (O_374,N_8433,N_8211);
or UO_375 (O_375,N_9184,N_8610);
nor UO_376 (O_376,N_9142,N_9149);
nand UO_377 (O_377,N_8228,N_9427);
nand UO_378 (O_378,N_8507,N_8607);
nor UO_379 (O_379,N_9165,N_9029);
nand UO_380 (O_380,N_9247,N_8504);
nor UO_381 (O_381,N_9144,N_8595);
and UO_382 (O_382,N_8187,N_8189);
and UO_383 (O_383,N_9760,N_9467);
or UO_384 (O_384,N_9062,N_8562);
nand UO_385 (O_385,N_8461,N_9136);
and UO_386 (O_386,N_8040,N_8251);
nand UO_387 (O_387,N_8289,N_9551);
nor UO_388 (O_388,N_8011,N_9396);
or UO_389 (O_389,N_9382,N_8724);
nor UO_390 (O_390,N_9924,N_9369);
nor UO_391 (O_391,N_8794,N_9498);
nor UO_392 (O_392,N_9304,N_9464);
or UO_393 (O_393,N_9477,N_8144);
nor UO_394 (O_394,N_9317,N_9104);
nand UO_395 (O_395,N_9204,N_9390);
nor UO_396 (O_396,N_8689,N_8112);
nand UO_397 (O_397,N_8122,N_8094);
and UO_398 (O_398,N_9089,N_8401);
and UO_399 (O_399,N_8723,N_9650);
and UO_400 (O_400,N_8363,N_8003);
or UO_401 (O_401,N_8796,N_9038);
nand UO_402 (O_402,N_8167,N_9178);
nor UO_403 (O_403,N_9846,N_8369);
nor UO_404 (O_404,N_9713,N_8576);
nor UO_405 (O_405,N_8598,N_8510);
or UO_406 (O_406,N_8985,N_8161);
xor UO_407 (O_407,N_9753,N_8904);
nor UO_408 (O_408,N_9781,N_9367);
nand UO_409 (O_409,N_9325,N_8648);
or UO_410 (O_410,N_8032,N_8965);
and UO_411 (O_411,N_8116,N_8240);
or UO_412 (O_412,N_9025,N_9920);
nor UO_413 (O_413,N_8305,N_9988);
or UO_414 (O_414,N_9592,N_9997);
or UO_415 (O_415,N_9691,N_9145);
nor UO_416 (O_416,N_8013,N_9266);
nor UO_417 (O_417,N_9598,N_8960);
or UO_418 (O_418,N_9406,N_8840);
nor UO_419 (O_419,N_9482,N_8237);
or UO_420 (O_420,N_8800,N_8452);
nand UO_421 (O_421,N_8014,N_9033);
nor UO_422 (O_422,N_8392,N_8329);
or UO_423 (O_423,N_8994,N_9886);
and UO_424 (O_424,N_9919,N_8628);
nor UO_425 (O_425,N_8290,N_9123);
or UO_426 (O_426,N_8783,N_8335);
nand UO_427 (O_427,N_8710,N_8017);
and UO_428 (O_428,N_9718,N_8937);
nor UO_429 (O_429,N_9878,N_9872);
or UO_430 (O_430,N_9156,N_8538);
or UO_431 (O_431,N_9541,N_9389);
nand UO_432 (O_432,N_9486,N_8143);
nand UO_433 (O_433,N_8298,N_8028);
nand UO_434 (O_434,N_8214,N_8727);
nand UO_435 (O_435,N_9463,N_9425);
nand UO_436 (O_436,N_8867,N_9480);
or UO_437 (O_437,N_9120,N_8565);
nor UO_438 (O_438,N_9451,N_9058);
nor UO_439 (O_439,N_9245,N_9205);
or UO_440 (O_440,N_9928,N_8209);
nor UO_441 (O_441,N_9885,N_9404);
and UO_442 (O_442,N_9802,N_8286);
nand UO_443 (O_443,N_9769,N_9594);
or UO_444 (O_444,N_9454,N_9456);
or UO_445 (O_445,N_9295,N_8618);
nand UO_446 (O_446,N_9804,N_8470);
nand UO_447 (O_447,N_9066,N_8499);
nor UO_448 (O_448,N_9843,N_8524);
nand UO_449 (O_449,N_9275,N_8671);
or UO_450 (O_450,N_8205,N_8023);
and UO_451 (O_451,N_9465,N_8375);
nor UO_452 (O_452,N_8918,N_8672);
nor UO_453 (O_453,N_8097,N_9070);
nor UO_454 (O_454,N_8496,N_9347);
nand UO_455 (O_455,N_8402,N_9770);
nand UO_456 (O_456,N_9792,N_9401);
and UO_457 (O_457,N_9314,N_9956);
or UO_458 (O_458,N_9507,N_8961);
and UO_459 (O_459,N_9719,N_8169);
and UO_460 (O_460,N_8165,N_9352);
nor UO_461 (O_461,N_9439,N_8516);
and UO_462 (O_462,N_8922,N_9937);
and UO_463 (O_463,N_8619,N_8479);
and UO_464 (O_464,N_9502,N_8912);
nand UO_465 (O_465,N_9972,N_9736);
nand UO_466 (O_466,N_9516,N_9476);
and UO_467 (O_467,N_8787,N_8026);
or UO_468 (O_468,N_9398,N_9350);
and UO_469 (O_469,N_9672,N_9235);
and UO_470 (O_470,N_9141,N_9115);
or UO_471 (O_471,N_8466,N_9194);
nor UO_472 (O_472,N_9378,N_9240);
or UO_473 (O_473,N_9346,N_9722);
and UO_474 (O_474,N_9050,N_8797);
nand UO_475 (O_475,N_8856,N_9732);
and UO_476 (O_476,N_9045,N_8809);
nand UO_477 (O_477,N_9225,N_9495);
and UO_478 (O_478,N_8589,N_8725);
nand UO_479 (O_479,N_8424,N_8258);
and UO_480 (O_480,N_8080,N_9570);
nand UO_481 (O_481,N_8139,N_9927);
nor UO_482 (O_482,N_8512,N_8968);
and UO_483 (O_483,N_9709,N_8572);
nand UO_484 (O_484,N_8403,N_8776);
and UO_485 (O_485,N_8309,N_9552);
nand UO_486 (O_486,N_8264,N_8745);
or UO_487 (O_487,N_8098,N_8519);
nor UO_488 (O_488,N_8036,N_8090);
and UO_489 (O_489,N_9641,N_8656);
nand UO_490 (O_490,N_9630,N_8432);
nor UO_491 (O_491,N_9667,N_8441);
or UO_492 (O_492,N_8253,N_9073);
nor UO_493 (O_493,N_8106,N_9615);
nand UO_494 (O_494,N_8314,N_9523);
and UO_495 (O_495,N_8191,N_8859);
nor UO_496 (O_496,N_8234,N_8940);
nand UO_497 (O_497,N_9189,N_9784);
nor UO_498 (O_498,N_8909,N_8521);
nor UO_499 (O_499,N_8153,N_9778);
nand UO_500 (O_500,N_8069,N_9783);
nor UO_501 (O_501,N_8839,N_8602);
xor UO_502 (O_502,N_8162,N_9701);
and UO_503 (O_503,N_9940,N_8157);
and UO_504 (O_504,N_8771,N_8525);
or UO_505 (O_505,N_9960,N_8303);
nor UO_506 (O_506,N_9964,N_8982);
or UO_507 (O_507,N_8891,N_9183);
nand UO_508 (O_508,N_8919,N_8453);
nor UO_509 (O_509,N_8978,N_8035);
nand UO_510 (O_510,N_8357,N_9084);
nand UO_511 (O_511,N_8573,N_9702);
nor UO_512 (O_512,N_9530,N_8623);
nor UO_513 (O_513,N_8736,N_8230);
and UO_514 (O_514,N_8898,N_8876);
nor UO_515 (O_515,N_9791,N_8758);
or UO_516 (O_516,N_9836,N_8766);
or UO_517 (O_517,N_9460,N_8709);
or UO_518 (O_518,N_8941,N_9221);
and UO_519 (O_519,N_8608,N_8634);
and UO_520 (O_520,N_9625,N_8260);
or UO_521 (O_521,N_9681,N_9661);
nand UO_522 (O_522,N_9216,N_9394);
nor UO_523 (O_523,N_9540,N_9677);
nand UO_524 (O_524,N_9793,N_8212);
nor UO_525 (O_525,N_8465,N_8914);
and UO_526 (O_526,N_8939,N_9360);
nand UO_527 (O_527,N_8615,N_8282);
nor UO_528 (O_528,N_8899,N_9051);
xnor UO_529 (O_529,N_8850,N_8002);
nor UO_530 (O_530,N_9556,N_9742);
or UO_531 (O_531,N_8808,N_8371);
or UO_532 (O_532,N_9220,N_9124);
nor UO_533 (O_533,N_8219,N_8206);
nor UO_534 (O_534,N_8788,N_9409);
and UO_535 (O_535,N_9143,N_9648);
or UO_536 (O_536,N_9201,N_8384);
nor UO_537 (O_537,N_8843,N_9587);
or UO_538 (O_538,N_8435,N_9690);
nand UO_539 (O_539,N_9449,N_8886);
nand UO_540 (O_540,N_9302,N_9081);
and UO_541 (O_541,N_9343,N_8987);
and UO_542 (O_542,N_8951,N_8255);
or UO_543 (O_543,N_8863,N_8045);
or UO_544 (O_544,N_9686,N_9250);
and UO_545 (O_545,N_8837,N_8059);
or UO_546 (O_546,N_8601,N_8185);
nor UO_547 (O_547,N_9496,N_8633);
or UO_548 (O_548,N_9262,N_8906);
and UO_549 (O_549,N_9584,N_9858);
and UO_550 (O_550,N_8612,N_9428);
and UO_551 (O_551,N_8666,N_8636);
or UO_552 (O_552,N_8113,N_9660);
nand UO_553 (O_553,N_9602,N_9096);
or UO_554 (O_554,N_9620,N_8690);
nand UO_555 (O_555,N_8584,N_8566);
nand UO_556 (O_556,N_9355,N_8390);
nor UO_557 (O_557,N_8581,N_9227);
nand UO_558 (O_558,N_8995,N_9990);
and UO_559 (O_559,N_9971,N_9524);
and UO_560 (O_560,N_9595,N_9341);
nor UO_561 (O_561,N_8273,N_9761);
nor UO_562 (O_562,N_8541,N_9871);
nor UO_563 (O_563,N_8897,N_9571);
nor UO_564 (O_564,N_8347,N_8587);
or UO_565 (O_565,N_9067,N_9538);
nand UO_566 (O_566,N_8256,N_8215);
and UO_567 (O_567,N_8900,N_9622);
and UO_568 (O_568,N_9192,N_8917);
and UO_569 (O_569,N_9656,N_8203);
and UO_570 (O_570,N_9828,N_9239);
nor UO_571 (O_571,N_9985,N_9488);
or UO_572 (O_572,N_8397,N_8247);
and UO_573 (O_573,N_8204,N_9077);
or UO_574 (O_574,N_8847,N_9161);
or UO_575 (O_575,N_9779,N_8311);
and UO_576 (O_576,N_8746,N_8871);
or UO_577 (O_577,N_8467,N_8079);
and UO_578 (O_578,N_8208,N_9252);
or UO_579 (O_579,N_8767,N_9585);
nor UO_580 (O_580,N_8066,N_9561);
nor UO_581 (O_581,N_9082,N_8186);
and UO_582 (O_582,N_8778,N_9433);
nand UO_583 (O_583,N_8233,N_9533);
nand UO_584 (O_584,N_9790,N_9209);
or UO_585 (O_585,N_8954,N_9442);
and UO_586 (O_586,N_9765,N_8523);
nand UO_587 (O_587,N_9900,N_9006);
nand UO_588 (O_588,N_8518,N_8854);
nor UO_589 (O_589,N_8073,N_9276);
nand UO_590 (O_590,N_9147,N_9902);
and UO_591 (O_591,N_8515,N_9299);
nand UO_592 (O_592,N_8908,N_9392);
nor UO_593 (O_593,N_9435,N_9898);
nand UO_594 (O_594,N_8316,N_8894);
or UO_595 (O_595,N_9608,N_8729);
nor UO_596 (O_596,N_9455,N_8020);
or UO_597 (O_597,N_9169,N_8578);
nor UO_598 (O_598,N_8111,N_9100);
or UO_599 (O_599,N_9337,N_8142);
or UO_600 (O_600,N_9132,N_9044);
and UO_601 (O_601,N_9362,N_9860);
nor UO_602 (O_602,N_9929,N_9938);
nand UO_603 (O_603,N_9152,N_8238);
nor UO_604 (O_604,N_9356,N_9755);
and UO_605 (O_605,N_8552,N_8093);
nand UO_606 (O_606,N_8704,N_8651);
and UO_607 (O_607,N_9599,N_9175);
or UO_608 (O_608,N_9825,N_9265);
or UO_609 (O_609,N_8312,N_8096);
and UO_610 (O_610,N_9374,N_8221);
nand UO_611 (O_611,N_9232,N_9429);
nor UO_612 (O_612,N_8811,N_8966);
nor UO_613 (O_613,N_8664,N_9424);
nor UO_614 (O_614,N_8004,N_8509);
nor UO_615 (O_615,N_8582,N_8295);
nor UO_616 (O_616,N_8963,N_8019);
nor UO_617 (O_617,N_9932,N_8667);
nor UO_618 (O_618,N_9505,N_8137);
or UO_619 (O_619,N_8317,N_9577);
nor UO_620 (O_620,N_8484,N_8232);
nand UO_621 (O_621,N_9866,N_8775);
and UO_622 (O_622,N_8896,N_9694);
or UO_623 (O_623,N_9795,N_8062);
or UO_624 (O_624,N_8687,N_8364);
nor UO_625 (O_625,N_9162,N_9695);
or UO_626 (O_626,N_9223,N_8377);
nor UO_627 (O_627,N_8743,N_8487);
nand UO_628 (O_628,N_8039,N_8535);
nor UO_629 (O_629,N_9642,N_9856);
and UO_630 (O_630,N_8857,N_8408);
nor UO_631 (O_631,N_8081,N_9282);
and UO_632 (O_632,N_8822,N_9320);
and UO_633 (O_633,N_9187,N_9453);
nor UO_634 (O_634,N_9700,N_8851);
nor UO_635 (O_635,N_8288,N_8133);
nand UO_636 (O_636,N_8913,N_9155);
and UO_637 (O_637,N_8196,N_9503);
nor UO_638 (O_638,N_8156,N_9782);
nor UO_639 (O_639,N_8200,N_9851);
or UO_640 (O_640,N_8389,N_9164);
nand UO_641 (O_641,N_9815,N_8824);
nand UO_642 (O_642,N_8701,N_9892);
or UO_643 (O_643,N_8485,N_8865);
or UO_644 (O_644,N_9669,N_9271);
nor UO_645 (O_645,N_9738,N_9407);
nand UO_646 (O_646,N_9167,N_9213);
and UO_647 (O_647,N_9270,N_8658);
and UO_648 (O_648,N_9327,N_9808);
nand UO_649 (O_649,N_8702,N_8864);
or UO_650 (O_650,N_9726,N_9186);
nor UO_651 (O_651,N_9448,N_8125);
nor UO_652 (O_652,N_8529,N_9749);
nand UO_653 (O_653,N_8431,N_9415);
nand UO_654 (O_654,N_8537,N_8660);
nor UO_655 (O_655,N_9434,N_9334);
nor UO_656 (O_656,N_9461,N_8287);
nor UO_657 (O_657,N_8975,N_9508);
or UO_658 (O_658,N_9546,N_9811);
and UO_659 (O_659,N_9881,N_8345);
and UO_660 (O_660,N_8564,N_8772);
nor UO_661 (O_661,N_8892,N_8355);
and UO_662 (O_662,N_9080,N_9174);
or UO_663 (O_663,N_9735,N_9479);
nand UO_664 (O_664,N_9525,N_9913);
nor UO_665 (O_665,N_9286,N_8749);
and UO_666 (O_666,N_9633,N_9148);
and UO_667 (O_667,N_8561,N_8763);
nand UO_668 (O_668,N_8947,N_9377);
and UO_669 (O_669,N_9810,N_8751);
or UO_670 (O_670,N_9559,N_8991);
nand UO_671 (O_671,N_9101,N_8970);
nand UO_672 (O_672,N_9172,N_8115);
and UO_673 (O_673,N_9754,N_8770);
nor UO_674 (O_674,N_9646,N_8779);
and UO_675 (O_675,N_8605,N_8006);
nand UO_676 (O_676,N_8436,N_8563);
nand UO_677 (O_677,N_8494,N_8150);
nand UO_678 (O_678,N_9258,N_9191);
nor UO_679 (O_679,N_9916,N_8356);
nor UO_680 (O_680,N_9568,N_9215);
or UO_681 (O_681,N_8825,N_9399);
nand UO_682 (O_682,N_9046,N_9002);
and UO_683 (O_683,N_8421,N_8367);
nand UO_684 (O_684,N_8910,N_9814);
nor UO_685 (O_685,N_8224,N_9831);
nand UO_686 (O_686,N_9896,N_9312);
nand UO_687 (O_687,N_9759,N_8365);
nand UO_688 (O_688,N_8744,N_8753);
nand UO_689 (O_689,N_8471,N_8781);
or UO_690 (O_690,N_9746,N_8500);
or UO_691 (O_691,N_9670,N_9263);
xor UO_692 (O_692,N_8964,N_8015);
nand UO_693 (O_693,N_9260,N_8726);
and UO_694 (O_694,N_8613,N_8569);
nor UO_695 (O_695,N_8301,N_9373);
nor UO_696 (O_696,N_9190,N_8626);
nand UO_697 (O_697,N_9365,N_9103);
nand UO_698 (O_698,N_8506,N_8380);
or UO_699 (O_699,N_9948,N_9673);
nand UO_700 (O_700,N_9922,N_8663);
or UO_701 (O_701,N_8807,N_9944);
nor UO_702 (O_702,N_8346,N_8574);
nand UO_703 (O_703,N_9775,N_9549);
nor UO_704 (O_704,N_9207,N_8332);
or UO_705 (O_705,N_8327,N_9122);
nor UO_706 (O_706,N_8957,N_8449);
nor UO_707 (O_707,N_8943,N_8550);
and UO_708 (O_708,N_9921,N_9529);
or UO_709 (O_709,N_8728,N_9975);
or UO_710 (O_710,N_9087,N_8361);
nand UO_711 (O_711,N_8095,N_9613);
and UO_712 (O_712,N_8489,N_8793);
and UO_713 (O_713,N_8557,N_9947);
or UO_714 (O_714,N_9129,N_9474);
and UO_715 (O_715,N_8675,N_8737);
or UO_716 (O_716,N_8996,N_9845);
and UO_717 (O_717,N_9316,N_8091);
nand UO_718 (O_718,N_8493,N_9796);
and UO_719 (O_719,N_9993,N_8659);
and UO_720 (O_720,N_9612,N_8720);
and UO_721 (O_721,N_8274,N_8041);
nand UO_722 (O_722,N_9991,N_9279);
nor UO_723 (O_723,N_8052,N_9109);
or UO_724 (O_724,N_8764,N_8853);
nand UO_725 (O_725,N_9563,N_9135);
nor UO_726 (O_726,N_9297,N_9509);
or UO_727 (O_727,N_9995,N_9750);
nor UO_728 (O_728,N_8418,N_8370);
nand UO_729 (O_729,N_9212,N_8246);
or UO_730 (O_730,N_8218,N_8163);
nand UO_731 (O_731,N_8542,N_8977);
or UO_732 (O_732,N_8445,N_8199);
or UO_733 (O_733,N_9269,N_9976);
nand UO_734 (O_734,N_9627,N_8170);
or UO_735 (O_735,N_9515,N_8703);
nor UO_736 (O_736,N_9357,N_9466);
and UO_737 (O_737,N_8434,N_8818);
and UO_738 (O_738,N_8785,N_9912);
nor UO_739 (O_739,N_8868,N_9180);
and UO_740 (O_740,N_9253,N_9114);
or UO_741 (O_741,N_8009,N_8333);
or UO_742 (O_742,N_8308,N_8409);
and UO_743 (O_743,N_9107,N_8606);
nand UO_744 (O_744,N_8738,N_8933);
nor UO_745 (O_745,N_9682,N_8307);
nand UO_746 (O_746,N_9961,N_9863);
or UO_747 (O_747,N_8654,N_8650);
nor UO_748 (O_748,N_8428,N_8319);
or UO_749 (O_749,N_8468,N_9534);
nand UO_750 (O_750,N_8821,N_8472);
nor UO_751 (O_751,N_9767,N_9366);
or UO_752 (O_752,N_9891,N_9288);
or UO_753 (O_753,N_9335,N_9785);
and UO_754 (O_754,N_9226,N_8734);
nand UO_755 (O_755,N_8885,N_8192);
and UO_756 (O_756,N_9086,N_9893);
and UO_757 (O_757,N_8888,N_9274);
or UO_758 (O_758,N_8076,N_8713);
nand UO_759 (O_759,N_9310,N_8334);
nor UO_760 (O_760,N_9249,N_8119);
nand UO_761 (O_761,N_9168,N_8057);
and UO_762 (O_762,N_9340,N_8935);
and UO_763 (O_763,N_9609,N_9987);
nor UO_764 (O_764,N_8340,N_9003);
or UO_765 (O_765,N_8860,N_9711);
nor UO_766 (O_766,N_8750,N_8469);
and UO_767 (O_767,N_9805,N_8590);
nand UO_768 (O_768,N_8498,N_9724);
and UO_769 (O_769,N_8679,N_9200);
nand UO_770 (O_770,N_9281,N_9823);
nand UO_771 (O_771,N_8969,N_9208);
and UO_772 (O_772,N_8832,N_9042);
or UO_773 (O_773,N_9847,N_9807);
nand UO_774 (O_774,N_9555,N_8585);
nor UO_775 (O_775,N_9364,N_9117);
and UO_776 (O_776,N_9657,N_8981);
nor UO_777 (O_777,N_9333,N_9649);
and UO_778 (O_778,N_8008,N_8786);
and UO_779 (O_779,N_9999,N_9567);
nor UO_780 (O_780,N_9776,N_9930);
or UO_781 (O_781,N_8044,N_9521);
nand UO_782 (O_782,N_8302,N_9697);
nor UO_783 (O_783,N_9949,N_9542);
nor UO_784 (O_784,N_8210,N_8001);
or UO_785 (O_785,N_8692,N_9376);
or UO_786 (O_786,N_9418,N_9473);
nand UO_787 (O_787,N_9395,N_8570);
or UO_788 (O_788,N_8682,N_8269);
nor UO_789 (O_789,N_8175,N_8528);
or UO_790 (O_790,N_8195,N_8158);
and UO_791 (O_791,N_8874,N_8488);
or UO_792 (O_792,N_9211,N_8643);
or UO_793 (O_793,N_9824,N_8945);
or UO_794 (O_794,N_8647,N_9102);
or UO_795 (O_795,N_8513,N_9163);
nand UO_796 (O_796,N_9731,N_8123);
or UO_797 (O_797,N_9095,N_9354);
and UO_798 (O_798,N_8171,N_9545);
or UO_799 (O_799,N_8816,N_9158);
and UO_800 (O_800,N_8382,N_9111);
and UO_801 (O_801,N_8136,N_9705);
or UO_802 (O_802,N_8490,N_9941);
nand UO_803 (O_803,N_9708,N_9313);
and UO_804 (O_804,N_9336,N_8719);
nand UO_805 (O_805,N_8394,N_8077);
and UO_806 (O_806,N_8614,N_8272);
nand UO_807 (O_807,N_8088,N_9659);
nor UO_808 (O_808,N_9492,N_9748);
or UO_809 (O_809,N_8053,N_9093);
or UO_810 (O_810,N_9052,N_9458);
or UO_811 (O_811,N_9777,N_9363);
nand UO_812 (O_812,N_8422,N_8972);
nand UO_813 (O_813,N_8188,N_9740);
and UO_814 (O_814,N_9375,N_8769);
nand UO_815 (O_815,N_9511,N_8920);
nor UO_816 (O_816,N_8752,N_9278);
or UO_817 (O_817,N_9531,N_9009);
nand UO_818 (O_818,N_8712,N_8398);
nor UO_819 (O_819,N_8759,N_9655);
or UO_820 (O_820,N_8058,N_9520);
or UO_821 (O_821,N_9809,N_9068);
nand UO_822 (O_822,N_9841,N_9899);
nand UO_823 (O_823,N_8104,N_9097);
nand UO_824 (O_824,N_8721,N_8268);
nand UO_825 (O_825,N_8711,N_8250);
nor UO_826 (O_826,N_8140,N_8603);
and UO_827 (O_827,N_8999,N_8952);
and UO_828 (O_828,N_8903,N_9030);
and UO_829 (O_829,N_8243,N_9015);
or UO_830 (O_830,N_9007,N_9384);
nor UO_831 (O_831,N_8491,N_8544);
nor UO_832 (O_832,N_9475,N_8866);
nor UO_833 (O_833,N_8717,N_9179);
nand UO_834 (O_834,N_8297,N_9992);
and UO_835 (O_835,N_8655,N_9803);
or UO_836 (O_836,N_9654,N_8804);
nand UO_837 (O_837,N_8694,N_9710);
nand UO_838 (O_838,N_9717,N_8477);
and UO_839 (O_839,N_9751,N_9910);
or UO_840 (O_840,N_9869,N_8976);
nor UO_841 (O_841,N_9623,N_8202);
and UO_842 (O_842,N_8277,N_9797);
xor UO_843 (O_843,N_8732,N_8145);
or UO_844 (O_844,N_8278,N_8292);
nand UO_845 (O_845,N_9739,N_9752);
and UO_846 (O_846,N_8555,N_8138);
nand UO_847 (O_847,N_9321,N_8147);
or UO_848 (O_848,N_8381,N_8458);
nor UO_849 (O_849,N_9470,N_8033);
or UO_850 (O_850,N_8556,N_8641);
or UO_851 (O_851,N_9639,N_9116);
and UO_852 (O_852,N_9059,N_8640);
nor UO_853 (O_853,N_8588,N_8846);
nor UO_854 (O_854,N_8986,N_9518);
nor UO_855 (O_855,N_8025,N_8828);
or UO_856 (O_856,N_8135,N_9231);
nor UO_857 (O_857,N_9151,N_9658);
or UO_858 (O_858,N_8248,N_8790);
nand UO_859 (O_859,N_9763,N_9008);
and UO_860 (O_860,N_8315,N_9589);
and UO_861 (O_861,N_9079,N_8118);
nor UO_862 (O_862,N_9219,N_8984);
and UO_863 (O_863,N_9217,N_8478);
nor UO_864 (O_864,N_8522,N_8055);
and UO_865 (O_865,N_8974,N_8338);
nor UO_866 (O_866,N_8121,N_9604);
nor UO_867 (O_867,N_8173,N_9359);
nand UO_868 (O_868,N_9386,N_9481);
or UO_869 (O_869,N_8283,N_8000);
nor UO_870 (O_870,N_9490,N_8979);
nor UO_871 (O_871,N_8844,N_9171);
nor UO_872 (O_872,N_8114,N_9787);
nor UO_873 (O_873,N_9462,N_9591);
nor UO_874 (O_874,N_9146,N_8503);
or UO_875 (O_875,N_9383,N_9020);
nor UO_876 (O_876,N_8700,N_9345);
nor UO_877 (O_877,N_9816,N_9652);
xnor UO_878 (O_878,N_9879,N_9914);
or UO_879 (O_879,N_9125,N_9251);
nand UO_880 (O_880,N_8061,N_8105);
or UO_881 (O_881,N_8760,N_8074);
and UO_882 (O_882,N_9638,N_9379);
and UO_883 (O_883,N_9432,N_9689);
nand UO_884 (O_884,N_9904,N_9606);
or UO_885 (O_885,N_9943,N_8688);
nor UO_886 (O_886,N_9850,N_8416);
nand UO_887 (O_887,N_9510,N_8084);
and UO_888 (O_888,N_8670,N_9255);
and UO_889 (O_889,N_8442,N_8950);
and UO_890 (O_890,N_8007,N_9973);
and UO_891 (O_891,N_9222,N_9889);
nand UO_892 (O_892,N_9698,N_9289);
and UO_893 (O_893,N_8884,N_9772);
nor UO_894 (O_894,N_8831,N_9064);
or UO_895 (O_895,N_8227,N_9822);
nand UO_896 (O_896,N_9022,N_9254);
and UO_897 (O_897,N_9653,N_9309);
nor UO_898 (O_898,N_9324,N_9478);
and UO_899 (O_899,N_8762,N_8027);
and UO_900 (O_900,N_8385,N_9611);
nor UO_901 (O_901,N_9688,N_8393);
or UO_902 (O_902,N_9861,N_8360);
nor UO_903 (O_903,N_8245,N_8532);
nand UO_904 (O_904,N_8457,N_8923);
nand UO_905 (O_905,N_9918,N_9907);
nand UO_906 (O_906,N_8921,N_9519);
or UO_907 (O_907,N_8223,N_9328);
and UO_908 (O_908,N_9526,N_9400);
or UO_909 (O_909,N_8152,N_9637);
or UO_910 (O_910,N_8222,N_8580);
and UO_911 (O_911,N_8075,N_8120);
nand UO_912 (O_912,N_8774,N_9085);
and UO_913 (O_913,N_8411,N_9833);
nor UO_914 (O_914,N_9894,N_8320);
nand UO_915 (O_915,N_9629,N_8931);
and UO_916 (O_916,N_8064,N_9897);
and UO_917 (O_917,N_9624,N_8833);
and UO_918 (O_918,N_9348,N_9915);
or UO_919 (O_919,N_8740,N_8372);
xor UO_920 (O_920,N_8180,N_8678);
or UO_921 (O_921,N_9756,N_9438);
or UO_922 (O_922,N_8213,N_8492);
nor UO_923 (O_923,N_9423,N_9011);
nand UO_924 (O_924,N_8929,N_9197);
nand UO_925 (O_925,N_8342,N_9293);
and UO_926 (O_926,N_8399,N_8548);
nand UO_927 (O_927,N_8915,N_8046);
and UO_928 (O_928,N_9371,N_9483);
nor UO_929 (O_929,N_9090,N_9569);
or UO_930 (O_930,N_9536,N_9596);
nor UO_931 (O_931,N_8293,N_9664);
and UO_932 (O_932,N_8082,N_9663);
nor UO_933 (O_933,N_9539,N_8586);
nand UO_934 (O_934,N_9844,N_9268);
nand UO_935 (O_935,N_9954,N_9447);
nand UO_936 (O_936,N_9290,N_9877);
nand UO_937 (O_937,N_8901,N_8437);
nor UO_938 (O_938,N_9131,N_9679);
and UO_939 (O_939,N_9727,N_8056);
nor UO_940 (O_940,N_9195,N_8916);
nand UO_941 (O_941,N_9946,N_8934);
nand UO_942 (O_942,N_8448,N_8034);
nand UO_943 (O_943,N_8993,N_9485);
and UO_944 (O_944,N_9883,N_9028);
nor UO_945 (O_945,N_9636,N_9242);
or UO_946 (O_946,N_9233,N_9361);
and UO_947 (O_947,N_8358,N_8583);
and UO_948 (O_948,N_8231,N_8517);
nand UO_949 (O_949,N_9838,N_8430);
nor UO_950 (O_950,N_8649,N_9543);
and UO_951 (O_951,N_9848,N_9855);
nor UO_952 (O_952,N_9895,N_9160);
nand UO_953 (O_953,N_9617,N_9957);
nand UO_954 (O_954,N_9410,N_8241);
and UO_955 (O_955,N_9626,N_9853);
nor UO_956 (O_956,N_8388,N_9444);
nand UO_957 (O_957,N_9351,N_9901);
and UO_958 (O_958,N_9905,N_8164);
or UO_959 (O_959,N_9566,N_8877);
and UO_960 (O_960,N_8842,N_9867);
or UO_961 (O_961,N_8773,N_9181);
or UO_962 (O_962,N_9780,N_9047);
or UO_963 (O_963,N_9610,N_9741);
nand UO_964 (O_964,N_9818,N_9875);
nor UO_965 (O_965,N_8502,N_8483);
nand UO_966 (O_966,N_9457,N_9259);
and UO_967 (O_967,N_8406,N_8294);
nor UO_968 (O_968,N_8925,N_8693);
nor UO_969 (O_969,N_9338,N_9437);
or UO_970 (O_970,N_9326,N_9292);
and UO_971 (O_971,N_9857,N_8559);
and UO_972 (O_972,N_9721,N_8696);
or UO_973 (O_973,N_9616,N_8955);
nand UO_974 (O_974,N_8318,N_8083);
and UO_975 (O_975,N_8440,N_9296);
or UO_976 (O_976,N_8617,N_8782);
nor UO_977 (O_977,N_9074,N_9747);
and UO_978 (O_978,N_9564,N_8455);
nor UO_979 (O_979,N_9034,N_8042);
nor UO_980 (O_980,N_8412,N_8018);
nor UO_981 (O_981,N_8373,N_8102);
and UO_982 (O_982,N_8343,N_9842);
and UO_983 (O_983,N_8962,N_8823);
and UO_984 (O_984,N_8803,N_8942);
nor UO_985 (O_985,N_9884,N_9826);
nor UO_986 (O_986,N_8324,N_8624);
nand UO_987 (O_987,N_9024,N_9036);
and UO_988 (O_988,N_9834,N_8331);
and UO_989 (O_989,N_9385,N_8629);
and UO_990 (O_990,N_8285,N_9469);
and UO_991 (O_991,N_8798,N_9854);
and UO_992 (O_992,N_8127,N_9786);
nand UO_993 (O_993,N_9774,N_9870);
and UO_994 (O_994,N_9887,N_9413);
nor UO_995 (O_995,N_9264,N_9133);
nand UO_996 (O_996,N_8391,N_9277);
and UO_997 (O_997,N_9939,N_9026);
and UO_998 (O_998,N_9830,N_8353);
nand UO_999 (O_999,N_8631,N_9621);
nand UO_1000 (O_1000,N_8719,N_8817);
nor UO_1001 (O_1001,N_8670,N_9229);
nand UO_1002 (O_1002,N_8131,N_8568);
nor UO_1003 (O_1003,N_9290,N_8485);
nand UO_1004 (O_1004,N_8798,N_8746);
and UO_1005 (O_1005,N_8433,N_9240);
and UO_1006 (O_1006,N_8832,N_9927);
or UO_1007 (O_1007,N_8874,N_9499);
nor UO_1008 (O_1008,N_8562,N_8230);
or UO_1009 (O_1009,N_9247,N_8654);
nor UO_1010 (O_1010,N_8467,N_8901);
nand UO_1011 (O_1011,N_9847,N_8335);
or UO_1012 (O_1012,N_9932,N_9413);
or UO_1013 (O_1013,N_9160,N_8835);
and UO_1014 (O_1014,N_8544,N_8148);
nor UO_1015 (O_1015,N_8884,N_8975);
nor UO_1016 (O_1016,N_9917,N_8544);
or UO_1017 (O_1017,N_9379,N_8762);
nor UO_1018 (O_1018,N_9056,N_9950);
and UO_1019 (O_1019,N_8982,N_8805);
or UO_1020 (O_1020,N_8094,N_9268);
xor UO_1021 (O_1021,N_9554,N_9208);
nand UO_1022 (O_1022,N_8718,N_9639);
or UO_1023 (O_1023,N_9952,N_8533);
nor UO_1024 (O_1024,N_9519,N_9001);
or UO_1025 (O_1025,N_9991,N_9930);
and UO_1026 (O_1026,N_8543,N_8360);
nor UO_1027 (O_1027,N_8710,N_8731);
or UO_1028 (O_1028,N_9445,N_9798);
nand UO_1029 (O_1029,N_9434,N_9198);
nor UO_1030 (O_1030,N_9862,N_9886);
and UO_1031 (O_1031,N_8088,N_8778);
and UO_1032 (O_1032,N_8036,N_9628);
nand UO_1033 (O_1033,N_8585,N_9116);
nand UO_1034 (O_1034,N_9241,N_8154);
or UO_1035 (O_1035,N_9782,N_9211);
and UO_1036 (O_1036,N_8419,N_9037);
nor UO_1037 (O_1037,N_8492,N_9119);
or UO_1038 (O_1038,N_8233,N_8939);
and UO_1039 (O_1039,N_8996,N_9685);
and UO_1040 (O_1040,N_8720,N_8825);
xor UO_1041 (O_1041,N_8079,N_8278);
or UO_1042 (O_1042,N_9825,N_8335);
or UO_1043 (O_1043,N_8892,N_8250);
nand UO_1044 (O_1044,N_9481,N_9103);
and UO_1045 (O_1045,N_8005,N_8173);
nor UO_1046 (O_1046,N_9728,N_9256);
and UO_1047 (O_1047,N_8280,N_9120);
or UO_1048 (O_1048,N_8234,N_9011);
and UO_1049 (O_1049,N_8406,N_8696);
nand UO_1050 (O_1050,N_9013,N_8401);
nand UO_1051 (O_1051,N_9729,N_8207);
nand UO_1052 (O_1052,N_8684,N_8745);
and UO_1053 (O_1053,N_9442,N_8949);
and UO_1054 (O_1054,N_9517,N_8081);
and UO_1055 (O_1055,N_9542,N_9361);
or UO_1056 (O_1056,N_9917,N_9844);
or UO_1057 (O_1057,N_8824,N_9969);
nand UO_1058 (O_1058,N_8178,N_8219);
or UO_1059 (O_1059,N_9124,N_8222);
or UO_1060 (O_1060,N_9617,N_8130);
nor UO_1061 (O_1061,N_9704,N_8531);
xor UO_1062 (O_1062,N_9498,N_9095);
or UO_1063 (O_1063,N_9359,N_9012);
or UO_1064 (O_1064,N_8977,N_8558);
nor UO_1065 (O_1065,N_8765,N_8869);
or UO_1066 (O_1066,N_9347,N_8940);
and UO_1067 (O_1067,N_9865,N_9963);
nand UO_1068 (O_1068,N_8280,N_8570);
nor UO_1069 (O_1069,N_9683,N_9120);
or UO_1070 (O_1070,N_9839,N_8377);
nor UO_1071 (O_1071,N_8052,N_9119);
or UO_1072 (O_1072,N_9887,N_9640);
and UO_1073 (O_1073,N_9761,N_9955);
and UO_1074 (O_1074,N_9874,N_9454);
or UO_1075 (O_1075,N_9037,N_9228);
nor UO_1076 (O_1076,N_8001,N_9819);
and UO_1077 (O_1077,N_8834,N_8145);
nand UO_1078 (O_1078,N_9592,N_9894);
nand UO_1079 (O_1079,N_8692,N_9231);
nor UO_1080 (O_1080,N_8051,N_9576);
nand UO_1081 (O_1081,N_9764,N_8828);
nor UO_1082 (O_1082,N_8972,N_9351);
and UO_1083 (O_1083,N_8828,N_8580);
nor UO_1084 (O_1084,N_9304,N_9540);
nor UO_1085 (O_1085,N_9571,N_9356);
nand UO_1086 (O_1086,N_8493,N_9523);
or UO_1087 (O_1087,N_8818,N_9879);
nand UO_1088 (O_1088,N_9136,N_8270);
or UO_1089 (O_1089,N_9995,N_9467);
and UO_1090 (O_1090,N_8319,N_8309);
or UO_1091 (O_1091,N_9887,N_8826);
nand UO_1092 (O_1092,N_9981,N_9855);
nand UO_1093 (O_1093,N_9145,N_9681);
and UO_1094 (O_1094,N_8536,N_9764);
or UO_1095 (O_1095,N_8755,N_9531);
and UO_1096 (O_1096,N_9647,N_8940);
nor UO_1097 (O_1097,N_8799,N_8248);
or UO_1098 (O_1098,N_9952,N_9283);
xnor UO_1099 (O_1099,N_9267,N_9780);
and UO_1100 (O_1100,N_8357,N_9552);
and UO_1101 (O_1101,N_9094,N_8293);
nor UO_1102 (O_1102,N_9177,N_8444);
or UO_1103 (O_1103,N_9922,N_8519);
nand UO_1104 (O_1104,N_9084,N_9374);
or UO_1105 (O_1105,N_8352,N_9896);
or UO_1106 (O_1106,N_9336,N_9606);
nor UO_1107 (O_1107,N_9825,N_9447);
nor UO_1108 (O_1108,N_9673,N_9469);
and UO_1109 (O_1109,N_8924,N_8941);
and UO_1110 (O_1110,N_9406,N_9150);
or UO_1111 (O_1111,N_8369,N_8441);
and UO_1112 (O_1112,N_8921,N_9970);
or UO_1113 (O_1113,N_8439,N_8676);
nand UO_1114 (O_1114,N_9432,N_9418);
and UO_1115 (O_1115,N_9332,N_9005);
nand UO_1116 (O_1116,N_9936,N_8472);
nand UO_1117 (O_1117,N_8924,N_9796);
nor UO_1118 (O_1118,N_8735,N_9112);
nor UO_1119 (O_1119,N_9914,N_9686);
xnor UO_1120 (O_1120,N_9698,N_8962);
or UO_1121 (O_1121,N_9824,N_8224);
nor UO_1122 (O_1122,N_9476,N_9385);
nand UO_1123 (O_1123,N_8736,N_9909);
nand UO_1124 (O_1124,N_9450,N_8957);
and UO_1125 (O_1125,N_8550,N_9812);
xnor UO_1126 (O_1126,N_9040,N_9670);
and UO_1127 (O_1127,N_8182,N_9339);
nand UO_1128 (O_1128,N_9652,N_9509);
or UO_1129 (O_1129,N_9196,N_8759);
nor UO_1130 (O_1130,N_8782,N_9427);
and UO_1131 (O_1131,N_9794,N_8565);
nand UO_1132 (O_1132,N_8416,N_9090);
or UO_1133 (O_1133,N_8711,N_8788);
and UO_1134 (O_1134,N_9621,N_9522);
and UO_1135 (O_1135,N_8604,N_8415);
or UO_1136 (O_1136,N_8789,N_9093);
nand UO_1137 (O_1137,N_8738,N_9314);
nand UO_1138 (O_1138,N_8806,N_9465);
or UO_1139 (O_1139,N_8971,N_9495);
and UO_1140 (O_1140,N_9460,N_8245);
nand UO_1141 (O_1141,N_8037,N_9148);
nand UO_1142 (O_1142,N_8421,N_8406);
or UO_1143 (O_1143,N_8280,N_9981);
nand UO_1144 (O_1144,N_8231,N_8284);
and UO_1145 (O_1145,N_9112,N_9844);
nand UO_1146 (O_1146,N_9496,N_9987);
and UO_1147 (O_1147,N_9277,N_9661);
or UO_1148 (O_1148,N_8137,N_9591);
and UO_1149 (O_1149,N_9373,N_9224);
nand UO_1150 (O_1150,N_9818,N_8214);
nor UO_1151 (O_1151,N_8946,N_8170);
nand UO_1152 (O_1152,N_8897,N_8211);
and UO_1153 (O_1153,N_8421,N_8559);
nor UO_1154 (O_1154,N_9414,N_9580);
nor UO_1155 (O_1155,N_9070,N_8601);
and UO_1156 (O_1156,N_8739,N_8957);
nand UO_1157 (O_1157,N_9716,N_9817);
nand UO_1158 (O_1158,N_8305,N_8547);
and UO_1159 (O_1159,N_9609,N_8495);
nand UO_1160 (O_1160,N_8762,N_8025);
and UO_1161 (O_1161,N_9845,N_8354);
and UO_1162 (O_1162,N_9554,N_8496);
or UO_1163 (O_1163,N_8810,N_8016);
nand UO_1164 (O_1164,N_9464,N_9852);
nor UO_1165 (O_1165,N_8459,N_9819);
and UO_1166 (O_1166,N_9611,N_8563);
and UO_1167 (O_1167,N_8571,N_9328);
and UO_1168 (O_1168,N_9033,N_8228);
nor UO_1169 (O_1169,N_9488,N_9581);
and UO_1170 (O_1170,N_8152,N_9748);
or UO_1171 (O_1171,N_8100,N_8567);
or UO_1172 (O_1172,N_8588,N_8915);
nor UO_1173 (O_1173,N_9717,N_8806);
nor UO_1174 (O_1174,N_9894,N_9406);
or UO_1175 (O_1175,N_9478,N_9958);
or UO_1176 (O_1176,N_9868,N_9324);
or UO_1177 (O_1177,N_8654,N_8835);
and UO_1178 (O_1178,N_9718,N_9249);
or UO_1179 (O_1179,N_8349,N_9792);
nand UO_1180 (O_1180,N_8396,N_8263);
nand UO_1181 (O_1181,N_8139,N_9658);
and UO_1182 (O_1182,N_8284,N_9840);
nand UO_1183 (O_1183,N_9750,N_8319);
and UO_1184 (O_1184,N_8838,N_9658);
or UO_1185 (O_1185,N_9136,N_9470);
or UO_1186 (O_1186,N_9578,N_9410);
and UO_1187 (O_1187,N_8020,N_8412);
and UO_1188 (O_1188,N_8199,N_8212);
nor UO_1189 (O_1189,N_8444,N_8270);
and UO_1190 (O_1190,N_8644,N_8758);
nand UO_1191 (O_1191,N_9024,N_8269);
and UO_1192 (O_1192,N_8316,N_8881);
or UO_1193 (O_1193,N_9200,N_8717);
nor UO_1194 (O_1194,N_8632,N_9822);
nand UO_1195 (O_1195,N_9015,N_8772);
nor UO_1196 (O_1196,N_8703,N_9561);
nand UO_1197 (O_1197,N_8663,N_8214);
or UO_1198 (O_1198,N_9619,N_8622);
or UO_1199 (O_1199,N_9115,N_8722);
nand UO_1200 (O_1200,N_8532,N_8229);
nor UO_1201 (O_1201,N_9769,N_8297);
and UO_1202 (O_1202,N_9486,N_9117);
nand UO_1203 (O_1203,N_8220,N_8161);
nand UO_1204 (O_1204,N_9301,N_8577);
nor UO_1205 (O_1205,N_8035,N_9471);
nand UO_1206 (O_1206,N_9144,N_9911);
nand UO_1207 (O_1207,N_8917,N_8542);
and UO_1208 (O_1208,N_9753,N_8216);
nor UO_1209 (O_1209,N_8461,N_9575);
nand UO_1210 (O_1210,N_9482,N_9028);
and UO_1211 (O_1211,N_9109,N_8435);
nand UO_1212 (O_1212,N_8411,N_8956);
or UO_1213 (O_1213,N_9994,N_8937);
nand UO_1214 (O_1214,N_9757,N_8975);
or UO_1215 (O_1215,N_8831,N_9355);
nand UO_1216 (O_1216,N_8488,N_9054);
nand UO_1217 (O_1217,N_9217,N_9501);
or UO_1218 (O_1218,N_8398,N_9887);
and UO_1219 (O_1219,N_9806,N_9575);
or UO_1220 (O_1220,N_9184,N_8286);
and UO_1221 (O_1221,N_9456,N_8580);
nor UO_1222 (O_1222,N_8286,N_9227);
nand UO_1223 (O_1223,N_8265,N_8987);
or UO_1224 (O_1224,N_9864,N_9000);
or UO_1225 (O_1225,N_9663,N_9948);
or UO_1226 (O_1226,N_8973,N_9381);
or UO_1227 (O_1227,N_9959,N_9396);
and UO_1228 (O_1228,N_9182,N_9310);
and UO_1229 (O_1229,N_9416,N_8372);
nand UO_1230 (O_1230,N_8201,N_8614);
nor UO_1231 (O_1231,N_9673,N_8654);
nand UO_1232 (O_1232,N_9885,N_9503);
or UO_1233 (O_1233,N_9835,N_8643);
nand UO_1234 (O_1234,N_8552,N_9277);
and UO_1235 (O_1235,N_8122,N_8509);
nor UO_1236 (O_1236,N_9773,N_8652);
nand UO_1237 (O_1237,N_8115,N_9858);
and UO_1238 (O_1238,N_9322,N_8219);
and UO_1239 (O_1239,N_9521,N_9169);
nand UO_1240 (O_1240,N_8490,N_8414);
and UO_1241 (O_1241,N_9557,N_9409);
nand UO_1242 (O_1242,N_8648,N_8386);
or UO_1243 (O_1243,N_9322,N_8291);
nor UO_1244 (O_1244,N_9495,N_8364);
nor UO_1245 (O_1245,N_9056,N_9381);
and UO_1246 (O_1246,N_9100,N_9623);
nand UO_1247 (O_1247,N_8563,N_8841);
and UO_1248 (O_1248,N_9797,N_9828);
or UO_1249 (O_1249,N_8355,N_9322);
and UO_1250 (O_1250,N_9923,N_8660);
nor UO_1251 (O_1251,N_9910,N_8170);
nor UO_1252 (O_1252,N_9027,N_8674);
or UO_1253 (O_1253,N_9669,N_8748);
nor UO_1254 (O_1254,N_8808,N_9557);
nor UO_1255 (O_1255,N_9316,N_8765);
nor UO_1256 (O_1256,N_8569,N_9321);
nor UO_1257 (O_1257,N_9295,N_8638);
or UO_1258 (O_1258,N_8667,N_8611);
nand UO_1259 (O_1259,N_8399,N_9435);
and UO_1260 (O_1260,N_8496,N_9028);
nor UO_1261 (O_1261,N_8000,N_8823);
nor UO_1262 (O_1262,N_8120,N_8552);
and UO_1263 (O_1263,N_9870,N_9886);
nand UO_1264 (O_1264,N_8042,N_9407);
nor UO_1265 (O_1265,N_8691,N_8715);
nand UO_1266 (O_1266,N_8636,N_9179);
and UO_1267 (O_1267,N_8256,N_8299);
nor UO_1268 (O_1268,N_9304,N_9181);
nor UO_1269 (O_1269,N_8073,N_9887);
nor UO_1270 (O_1270,N_8980,N_9556);
nand UO_1271 (O_1271,N_9317,N_9668);
and UO_1272 (O_1272,N_8364,N_9063);
or UO_1273 (O_1273,N_9354,N_8803);
or UO_1274 (O_1274,N_8288,N_8473);
nor UO_1275 (O_1275,N_9201,N_8866);
nand UO_1276 (O_1276,N_8573,N_9592);
or UO_1277 (O_1277,N_8093,N_9059);
nand UO_1278 (O_1278,N_9064,N_9003);
or UO_1279 (O_1279,N_8710,N_8879);
or UO_1280 (O_1280,N_8387,N_9531);
nand UO_1281 (O_1281,N_8256,N_8342);
and UO_1282 (O_1282,N_9296,N_8359);
and UO_1283 (O_1283,N_9739,N_9887);
or UO_1284 (O_1284,N_8435,N_8869);
nor UO_1285 (O_1285,N_9989,N_8549);
nor UO_1286 (O_1286,N_8521,N_8162);
nor UO_1287 (O_1287,N_8286,N_8256);
nor UO_1288 (O_1288,N_9206,N_8116);
and UO_1289 (O_1289,N_9708,N_8439);
nor UO_1290 (O_1290,N_9183,N_9013);
and UO_1291 (O_1291,N_8120,N_9518);
or UO_1292 (O_1292,N_9245,N_8014);
and UO_1293 (O_1293,N_9036,N_9087);
nor UO_1294 (O_1294,N_8408,N_9489);
and UO_1295 (O_1295,N_8657,N_8294);
or UO_1296 (O_1296,N_9422,N_9183);
nand UO_1297 (O_1297,N_8210,N_9295);
nand UO_1298 (O_1298,N_8337,N_9621);
or UO_1299 (O_1299,N_9930,N_8261);
nor UO_1300 (O_1300,N_9282,N_8781);
or UO_1301 (O_1301,N_8083,N_8834);
and UO_1302 (O_1302,N_8681,N_8778);
nand UO_1303 (O_1303,N_9413,N_8153);
nor UO_1304 (O_1304,N_9985,N_8722);
or UO_1305 (O_1305,N_9100,N_8491);
or UO_1306 (O_1306,N_9669,N_9910);
nor UO_1307 (O_1307,N_8381,N_8704);
or UO_1308 (O_1308,N_9467,N_9276);
nand UO_1309 (O_1309,N_8706,N_8363);
and UO_1310 (O_1310,N_9753,N_8942);
nor UO_1311 (O_1311,N_9751,N_9125);
and UO_1312 (O_1312,N_8838,N_9313);
nand UO_1313 (O_1313,N_8967,N_8831);
nand UO_1314 (O_1314,N_8095,N_9734);
or UO_1315 (O_1315,N_9635,N_8650);
nand UO_1316 (O_1316,N_8552,N_8756);
nand UO_1317 (O_1317,N_9504,N_8970);
and UO_1318 (O_1318,N_9409,N_9577);
or UO_1319 (O_1319,N_9311,N_8342);
nor UO_1320 (O_1320,N_9164,N_9260);
nor UO_1321 (O_1321,N_8103,N_8737);
nor UO_1322 (O_1322,N_8336,N_8842);
and UO_1323 (O_1323,N_8971,N_9218);
nand UO_1324 (O_1324,N_8555,N_9129);
nor UO_1325 (O_1325,N_8649,N_9736);
nand UO_1326 (O_1326,N_9406,N_8528);
and UO_1327 (O_1327,N_8550,N_8588);
and UO_1328 (O_1328,N_9455,N_9700);
and UO_1329 (O_1329,N_8288,N_9915);
or UO_1330 (O_1330,N_8845,N_9450);
or UO_1331 (O_1331,N_9156,N_9361);
nand UO_1332 (O_1332,N_9169,N_8816);
nor UO_1333 (O_1333,N_9109,N_9407);
nand UO_1334 (O_1334,N_8524,N_8663);
nand UO_1335 (O_1335,N_9059,N_8889);
and UO_1336 (O_1336,N_8340,N_8091);
nor UO_1337 (O_1337,N_8143,N_8737);
nand UO_1338 (O_1338,N_9314,N_8149);
or UO_1339 (O_1339,N_8223,N_9584);
nand UO_1340 (O_1340,N_9448,N_9538);
and UO_1341 (O_1341,N_8410,N_8435);
nand UO_1342 (O_1342,N_9147,N_9380);
or UO_1343 (O_1343,N_8445,N_8074);
nand UO_1344 (O_1344,N_9913,N_8828);
and UO_1345 (O_1345,N_9990,N_9211);
and UO_1346 (O_1346,N_8835,N_9800);
and UO_1347 (O_1347,N_8103,N_8741);
nor UO_1348 (O_1348,N_8760,N_9454);
nand UO_1349 (O_1349,N_9079,N_8549);
or UO_1350 (O_1350,N_9290,N_9073);
and UO_1351 (O_1351,N_8064,N_9021);
or UO_1352 (O_1352,N_8173,N_8074);
nand UO_1353 (O_1353,N_8442,N_8673);
nand UO_1354 (O_1354,N_8845,N_9334);
nor UO_1355 (O_1355,N_8532,N_9632);
or UO_1356 (O_1356,N_9734,N_9473);
nand UO_1357 (O_1357,N_8118,N_8448);
and UO_1358 (O_1358,N_8661,N_9425);
nand UO_1359 (O_1359,N_8459,N_9886);
xnor UO_1360 (O_1360,N_9910,N_8293);
nand UO_1361 (O_1361,N_9246,N_9488);
or UO_1362 (O_1362,N_8315,N_9856);
nor UO_1363 (O_1363,N_8595,N_8019);
nand UO_1364 (O_1364,N_9130,N_8258);
and UO_1365 (O_1365,N_9278,N_8220);
nand UO_1366 (O_1366,N_9131,N_8103);
and UO_1367 (O_1367,N_9615,N_8418);
nor UO_1368 (O_1368,N_8015,N_8461);
and UO_1369 (O_1369,N_8535,N_8252);
or UO_1370 (O_1370,N_8331,N_9461);
and UO_1371 (O_1371,N_8088,N_9998);
xnor UO_1372 (O_1372,N_8719,N_9796);
or UO_1373 (O_1373,N_8087,N_9270);
nand UO_1374 (O_1374,N_8985,N_8059);
nand UO_1375 (O_1375,N_9316,N_8050);
or UO_1376 (O_1376,N_8338,N_9161);
or UO_1377 (O_1377,N_9323,N_8711);
nor UO_1378 (O_1378,N_9566,N_8711);
nand UO_1379 (O_1379,N_9663,N_8219);
and UO_1380 (O_1380,N_8321,N_9754);
or UO_1381 (O_1381,N_8848,N_9724);
nor UO_1382 (O_1382,N_9335,N_9599);
nand UO_1383 (O_1383,N_9628,N_8963);
and UO_1384 (O_1384,N_9787,N_9402);
nor UO_1385 (O_1385,N_8833,N_8022);
nor UO_1386 (O_1386,N_9508,N_8464);
nor UO_1387 (O_1387,N_8950,N_8030);
nor UO_1388 (O_1388,N_8705,N_9831);
nor UO_1389 (O_1389,N_8710,N_9372);
nand UO_1390 (O_1390,N_8730,N_9024);
and UO_1391 (O_1391,N_8571,N_8311);
and UO_1392 (O_1392,N_8825,N_8682);
or UO_1393 (O_1393,N_8501,N_9994);
or UO_1394 (O_1394,N_8296,N_9979);
nand UO_1395 (O_1395,N_9571,N_9825);
nor UO_1396 (O_1396,N_9016,N_9084);
and UO_1397 (O_1397,N_8424,N_8365);
or UO_1398 (O_1398,N_9064,N_9174);
nand UO_1399 (O_1399,N_8237,N_9406);
or UO_1400 (O_1400,N_9392,N_9153);
nor UO_1401 (O_1401,N_8634,N_8968);
or UO_1402 (O_1402,N_9963,N_9634);
or UO_1403 (O_1403,N_9253,N_9276);
nand UO_1404 (O_1404,N_9484,N_9755);
or UO_1405 (O_1405,N_8993,N_9984);
nand UO_1406 (O_1406,N_8767,N_8318);
nor UO_1407 (O_1407,N_8530,N_9199);
or UO_1408 (O_1408,N_8626,N_8663);
nand UO_1409 (O_1409,N_9021,N_8564);
nor UO_1410 (O_1410,N_8580,N_8843);
or UO_1411 (O_1411,N_9133,N_8394);
or UO_1412 (O_1412,N_9464,N_9062);
or UO_1413 (O_1413,N_8010,N_9899);
nor UO_1414 (O_1414,N_9170,N_9045);
nor UO_1415 (O_1415,N_8876,N_9421);
nor UO_1416 (O_1416,N_9975,N_9385);
or UO_1417 (O_1417,N_9626,N_9126);
and UO_1418 (O_1418,N_9732,N_9371);
and UO_1419 (O_1419,N_8061,N_9648);
nand UO_1420 (O_1420,N_8051,N_9587);
nor UO_1421 (O_1421,N_8546,N_9393);
nand UO_1422 (O_1422,N_9729,N_8600);
nand UO_1423 (O_1423,N_8596,N_8841);
nand UO_1424 (O_1424,N_8121,N_9835);
nor UO_1425 (O_1425,N_8988,N_9927);
nand UO_1426 (O_1426,N_8604,N_8142);
or UO_1427 (O_1427,N_8878,N_9255);
nand UO_1428 (O_1428,N_9692,N_8543);
and UO_1429 (O_1429,N_9973,N_8755);
and UO_1430 (O_1430,N_9431,N_8224);
nor UO_1431 (O_1431,N_9076,N_8450);
or UO_1432 (O_1432,N_8674,N_9799);
or UO_1433 (O_1433,N_9156,N_9258);
nand UO_1434 (O_1434,N_8643,N_9070);
or UO_1435 (O_1435,N_9764,N_8564);
nand UO_1436 (O_1436,N_8521,N_8663);
nor UO_1437 (O_1437,N_9343,N_9009);
and UO_1438 (O_1438,N_8961,N_8637);
nor UO_1439 (O_1439,N_8929,N_9256);
or UO_1440 (O_1440,N_9499,N_9024);
nor UO_1441 (O_1441,N_9074,N_9929);
and UO_1442 (O_1442,N_8071,N_9063);
nand UO_1443 (O_1443,N_8670,N_9143);
and UO_1444 (O_1444,N_9726,N_9402);
or UO_1445 (O_1445,N_8748,N_8629);
or UO_1446 (O_1446,N_8758,N_9325);
and UO_1447 (O_1447,N_9346,N_8014);
and UO_1448 (O_1448,N_8424,N_9859);
nor UO_1449 (O_1449,N_8520,N_8095);
or UO_1450 (O_1450,N_9415,N_9267);
and UO_1451 (O_1451,N_9061,N_9964);
or UO_1452 (O_1452,N_9069,N_8674);
or UO_1453 (O_1453,N_9490,N_9984);
or UO_1454 (O_1454,N_8685,N_9864);
nand UO_1455 (O_1455,N_9122,N_9050);
xor UO_1456 (O_1456,N_9937,N_9555);
and UO_1457 (O_1457,N_9505,N_8993);
nor UO_1458 (O_1458,N_8593,N_9731);
and UO_1459 (O_1459,N_9243,N_9060);
xor UO_1460 (O_1460,N_8318,N_9391);
xor UO_1461 (O_1461,N_9556,N_8969);
nor UO_1462 (O_1462,N_8332,N_9101);
or UO_1463 (O_1463,N_9075,N_9533);
nor UO_1464 (O_1464,N_8637,N_8410);
xor UO_1465 (O_1465,N_9559,N_9106);
nor UO_1466 (O_1466,N_9574,N_9114);
or UO_1467 (O_1467,N_8098,N_8423);
nor UO_1468 (O_1468,N_8422,N_8575);
or UO_1469 (O_1469,N_8851,N_8353);
nor UO_1470 (O_1470,N_9818,N_8523);
xnor UO_1471 (O_1471,N_8575,N_9352);
or UO_1472 (O_1472,N_9598,N_8335);
nor UO_1473 (O_1473,N_9267,N_9325);
or UO_1474 (O_1474,N_8504,N_8626);
nand UO_1475 (O_1475,N_9018,N_9048);
or UO_1476 (O_1476,N_8309,N_9396);
nand UO_1477 (O_1477,N_9259,N_9252);
nand UO_1478 (O_1478,N_8659,N_9173);
and UO_1479 (O_1479,N_9106,N_8843);
nor UO_1480 (O_1480,N_8284,N_9529);
and UO_1481 (O_1481,N_9193,N_8504);
nand UO_1482 (O_1482,N_9901,N_8958);
and UO_1483 (O_1483,N_8525,N_8816);
and UO_1484 (O_1484,N_8941,N_8096);
and UO_1485 (O_1485,N_9227,N_9762);
and UO_1486 (O_1486,N_8959,N_9907);
and UO_1487 (O_1487,N_8700,N_8799);
and UO_1488 (O_1488,N_8635,N_9622);
nor UO_1489 (O_1489,N_9030,N_9208);
and UO_1490 (O_1490,N_9231,N_9239);
nor UO_1491 (O_1491,N_8876,N_9014);
or UO_1492 (O_1492,N_8464,N_8860);
or UO_1493 (O_1493,N_8563,N_8666);
nor UO_1494 (O_1494,N_9759,N_9817);
and UO_1495 (O_1495,N_8340,N_9236);
and UO_1496 (O_1496,N_8204,N_8901);
or UO_1497 (O_1497,N_8719,N_9203);
nand UO_1498 (O_1498,N_8327,N_9799);
nand UO_1499 (O_1499,N_9456,N_9666);
endmodule