module basic_2000_20000_2500_10_levels_5xor_3(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999;
or U0 (N_0,In_39,In_1273);
xnor U1 (N_1,In_893,In_1287);
nor U2 (N_2,In_600,In_1541);
and U3 (N_3,In_793,In_607);
nor U4 (N_4,In_1326,In_405);
nor U5 (N_5,In_330,In_1357);
xnor U6 (N_6,In_92,In_364);
xor U7 (N_7,In_1243,In_639);
nor U8 (N_8,In_316,In_574);
nand U9 (N_9,In_878,In_437);
nor U10 (N_10,In_1725,In_470);
and U11 (N_11,In_1871,In_1684);
nor U12 (N_12,In_219,In_519);
and U13 (N_13,In_848,In_1338);
nand U14 (N_14,In_1030,In_818);
nand U15 (N_15,In_962,In_1613);
nor U16 (N_16,In_1551,In_295);
nand U17 (N_17,In_11,In_1199);
xnor U18 (N_18,In_1997,In_1240);
xor U19 (N_19,In_1437,In_1635);
nor U20 (N_20,In_1227,In_1215);
xor U21 (N_21,In_732,In_551);
nand U22 (N_22,In_102,In_862);
nor U23 (N_23,In_823,In_185);
nand U24 (N_24,In_681,In_974);
nand U25 (N_25,In_897,In_1723);
nor U26 (N_26,In_716,In_441);
nor U27 (N_27,In_1773,In_56);
and U28 (N_28,In_356,In_1832);
or U29 (N_29,In_221,In_579);
or U30 (N_30,In_1789,In_237);
nor U31 (N_31,In_90,In_79);
or U32 (N_32,In_1519,In_1987);
nor U33 (N_33,In_1162,In_580);
and U34 (N_34,In_36,In_58);
nand U35 (N_35,In_1974,In_936);
and U36 (N_36,In_231,In_1529);
nand U37 (N_37,In_83,In_945);
nor U38 (N_38,In_1976,In_31);
nor U39 (N_39,In_747,In_1419);
nor U40 (N_40,In_876,In_1739);
or U41 (N_41,In_1523,In_224);
nor U42 (N_42,In_1284,In_1880);
xnor U43 (N_43,In_1319,In_808);
nand U44 (N_44,In_1986,In_1370);
and U45 (N_45,In_1194,In_1536);
nand U46 (N_46,In_1904,In_660);
xnor U47 (N_47,In_78,In_463);
nor U48 (N_48,In_1935,In_1810);
xnor U49 (N_49,In_326,In_1163);
and U50 (N_50,In_81,In_1881);
nor U51 (N_51,In_542,In_628);
or U52 (N_52,In_973,In_777);
nand U53 (N_53,In_1246,In_1957);
nor U54 (N_54,In_1527,In_120);
and U55 (N_55,In_63,In_835);
or U56 (N_56,In_544,In_697);
and U57 (N_57,In_1460,In_178);
and U58 (N_58,In_191,In_220);
and U59 (N_59,In_817,In_1205);
and U60 (N_60,In_863,In_443);
nor U61 (N_61,In_1663,In_1599);
nand U62 (N_62,In_243,In_57);
nor U63 (N_63,In_605,In_883);
nor U64 (N_64,In_869,In_1753);
or U65 (N_65,In_95,In_1433);
nor U66 (N_66,In_208,In_374);
nor U67 (N_67,In_1461,In_436);
and U68 (N_68,In_859,In_257);
nor U69 (N_69,In_711,In_718);
xor U70 (N_70,In_1265,In_957);
or U71 (N_71,In_748,In_1615);
and U72 (N_72,In_1320,In_928);
and U73 (N_73,In_961,In_1601);
nor U74 (N_74,In_563,In_595);
or U75 (N_75,In_1274,In_1127);
and U76 (N_76,In_1301,In_1268);
xnor U77 (N_77,In_1090,In_1920);
xor U78 (N_78,In_1761,In_1294);
nor U79 (N_79,In_907,In_1041);
or U80 (N_80,In_1256,In_1954);
nor U81 (N_81,In_1961,In_390);
or U82 (N_82,In_1702,In_810);
nand U83 (N_83,In_365,In_722);
or U84 (N_84,In_774,In_917);
and U85 (N_85,In_1557,In_392);
nor U86 (N_86,In_1735,In_1547);
xor U87 (N_87,In_1838,In_1740);
or U88 (N_88,In_1455,In_1799);
nand U89 (N_89,In_1448,In_753);
nand U90 (N_90,In_821,In_1905);
or U91 (N_91,In_1745,In_587);
and U92 (N_92,In_337,In_1015);
or U93 (N_93,In_223,In_1768);
and U94 (N_94,In_635,In_1754);
nor U95 (N_95,In_1766,In_1478);
nand U96 (N_96,In_880,In_1791);
or U97 (N_97,In_1975,In_1185);
or U98 (N_98,In_912,In_1836);
nor U99 (N_99,In_1874,In_241);
nand U100 (N_100,In_825,In_613);
nor U101 (N_101,In_1116,In_1355);
xor U102 (N_102,In_3,In_319);
nand U103 (N_103,In_1973,In_1129);
or U104 (N_104,In_1956,In_1432);
nor U105 (N_105,In_638,In_1701);
or U106 (N_106,In_686,In_1123);
nor U107 (N_107,In_834,In_116);
and U108 (N_108,In_664,In_976);
nor U109 (N_109,In_1902,In_278);
nor U110 (N_110,In_499,In_22);
nand U111 (N_111,In_1007,In_1855);
nand U112 (N_112,In_1397,In_1704);
and U113 (N_113,In_354,In_864);
nor U114 (N_114,In_1387,In_798);
nor U115 (N_115,In_643,In_1656);
nand U116 (N_116,In_949,In_302);
and U117 (N_117,In_577,In_355);
or U118 (N_118,In_1641,In_1606);
or U119 (N_119,In_1025,In_1984);
nand U120 (N_120,In_1180,In_1252);
and U121 (N_121,In_327,In_252);
xnor U122 (N_122,In_387,In_1339);
and U123 (N_123,In_73,In_1578);
or U124 (N_124,In_1166,In_1858);
and U125 (N_125,In_750,In_1164);
or U126 (N_126,In_1752,In_74);
and U127 (N_127,In_1781,In_1549);
or U128 (N_128,In_471,In_1833);
and U129 (N_129,In_778,In_626);
and U130 (N_130,In_474,In_135);
xor U131 (N_131,In_1762,In_1038);
and U132 (N_132,In_633,In_1614);
nor U133 (N_133,In_110,In_1383);
and U134 (N_134,In_46,In_1143);
or U135 (N_135,In_1085,In_476);
nand U136 (N_136,In_28,In_1012);
or U137 (N_137,In_1503,In_1457);
nand U138 (N_138,In_816,In_1934);
nor U139 (N_139,In_512,In_115);
nor U140 (N_140,In_588,In_1310);
and U141 (N_141,In_1089,In_145);
or U142 (N_142,In_1290,In_1170);
and U143 (N_143,In_1235,In_1378);
or U144 (N_144,In_561,In_1711);
nand U145 (N_145,In_304,In_1230);
or U146 (N_146,In_509,In_274);
xor U147 (N_147,In_153,In_589);
or U148 (N_148,In_382,In_1410);
and U149 (N_149,In_1347,In_867);
nand U150 (N_150,In_1024,In_738);
or U151 (N_151,In_1224,In_1767);
or U152 (N_152,In_1600,In_847);
xor U153 (N_153,In_282,In_1135);
xnor U154 (N_154,In_1292,In_204);
or U155 (N_155,In_1183,In_572);
nand U156 (N_156,In_363,In_797);
or U157 (N_157,In_35,In_1542);
or U158 (N_158,In_213,In_916);
or U159 (N_159,In_1354,In_1017);
or U160 (N_160,In_60,In_420);
nand U161 (N_161,In_473,In_1628);
or U162 (N_162,In_978,In_483);
nand U163 (N_163,In_1807,In_995);
nor U164 (N_164,In_1585,In_1271);
and U165 (N_165,In_743,In_306);
nand U166 (N_166,In_1996,In_1146);
and U167 (N_167,In_1122,In_1468);
or U168 (N_168,In_809,In_235);
and U169 (N_169,In_49,In_653);
and U170 (N_170,In_554,In_1169);
nand U171 (N_171,In_851,In_1808);
nand U172 (N_172,In_854,In_1106);
nor U173 (N_173,In_1534,In_1187);
or U174 (N_174,In_247,In_1982);
nand U175 (N_175,In_783,In_1848);
nor U176 (N_176,In_273,In_569);
and U177 (N_177,In_904,In_1298);
nor U178 (N_178,In_138,In_725);
or U179 (N_179,In_1335,In_1634);
nor U180 (N_180,In_1658,In_475);
xor U181 (N_181,In_1306,In_1342);
and U182 (N_182,In_1657,In_1411);
nand U183 (N_183,In_122,In_567);
xor U184 (N_184,In_1955,In_1396);
or U185 (N_185,In_1186,In_1640);
and U186 (N_186,In_581,In_1406);
and U187 (N_187,In_1108,In_837);
and U188 (N_188,In_421,In_1334);
nor U189 (N_189,In_1371,In_159);
and U190 (N_190,In_989,In_1720);
nor U191 (N_191,In_1321,In_1337);
or U192 (N_192,In_324,In_1039);
nor U193 (N_193,In_1184,In_1900);
and U194 (N_194,In_433,In_10);
nand U195 (N_195,In_256,In_1936);
and U196 (N_196,In_1716,In_173);
nor U197 (N_197,In_1736,In_1391);
nand U198 (N_198,In_1804,In_887);
or U199 (N_199,In_910,In_1824);
and U200 (N_200,In_1490,In_432);
nand U201 (N_201,In_998,In_712);
xnor U202 (N_202,In_1384,In_232);
or U203 (N_203,In_999,In_1167);
or U204 (N_204,In_1,In_1883);
or U205 (N_205,In_271,In_1266);
nor U206 (N_206,In_1071,In_1098);
and U207 (N_207,In_739,In_1176);
xor U208 (N_208,In_1400,In_152);
or U209 (N_209,In_180,In_1083);
nor U210 (N_210,In_647,In_1998);
nand U211 (N_211,In_1050,In_1653);
nor U212 (N_212,In_393,In_685);
xnor U213 (N_213,In_1423,In_1137);
xor U214 (N_214,In_856,In_77);
nor U215 (N_215,In_1308,In_766);
nand U216 (N_216,In_675,In_620);
nor U217 (N_217,In_1939,In_203);
xor U218 (N_218,In_983,In_118);
nand U219 (N_219,In_1282,In_866);
nor U220 (N_220,In_1075,In_1403);
and U221 (N_221,In_1792,In_1312);
and U222 (N_222,In_50,In_1811);
nor U223 (N_223,In_171,In_840);
and U224 (N_224,In_361,In_388);
or U225 (N_225,In_85,In_1897);
nor U226 (N_226,In_1210,In_611);
nor U227 (N_227,In_1722,In_320);
and U228 (N_228,In_1964,In_1124);
or U229 (N_229,In_1485,In_1788);
and U230 (N_230,In_1595,In_1484);
nand U231 (N_231,In_558,In_1237);
or U232 (N_232,In_1582,In_1719);
and U233 (N_233,In_591,In_762);
xnor U234 (N_234,In_1901,In_694);
nand U235 (N_235,In_871,In_309);
xnor U236 (N_236,In_651,In_264);
and U237 (N_237,In_1088,In_795);
or U238 (N_238,In_87,In_1348);
and U239 (N_239,In_98,In_1802);
nor U240 (N_240,In_1254,In_1577);
and U241 (N_241,In_24,In_1119);
and U242 (N_242,In_347,In_339);
and U243 (N_243,In_1280,In_710);
or U244 (N_244,In_955,In_625);
nand U245 (N_245,In_687,In_1200);
nand U246 (N_246,In_418,In_1607);
nand U247 (N_247,In_7,In_93);
or U248 (N_248,In_164,In_33);
nor U249 (N_249,In_258,In_1362);
nor U250 (N_250,In_1664,In_1061);
nand U251 (N_251,In_646,In_668);
xnor U252 (N_252,In_970,In_230);
nor U253 (N_253,In_202,In_1759);
nand U254 (N_254,In_670,In_1550);
or U255 (N_255,In_1456,In_953);
and U256 (N_256,In_1868,In_1506);
nor U257 (N_257,In_1450,In_458);
nand U258 (N_258,In_1245,In_62);
xor U259 (N_259,In_1795,In_715);
nor U260 (N_260,In_1856,In_1933);
and U261 (N_261,In_570,In_407);
and U262 (N_262,In_822,In_599);
or U263 (N_263,In_246,In_805);
nand U264 (N_264,In_1695,In_1544);
and U265 (N_265,In_1352,In_1692);
nand U266 (N_266,In_367,In_196);
xor U267 (N_267,In_129,In_398);
nand U268 (N_268,In_391,In_440);
and U269 (N_269,In_1144,In_1329);
nand U270 (N_270,In_394,In_858);
nor U271 (N_271,In_857,In_1053);
and U272 (N_272,In_467,In_1925);
nand U273 (N_273,In_915,In_1746);
and U274 (N_274,In_332,In_1912);
nand U275 (N_275,In_1676,In_1963);
and U276 (N_276,In_954,In_721);
nor U277 (N_277,In_526,In_336);
nor U278 (N_278,In_444,In_99);
nand U279 (N_279,In_1983,In_1511);
nor U280 (N_280,In_1580,In_490);
and U281 (N_281,In_67,In_1532);
nand U282 (N_282,In_1943,In_1046);
or U283 (N_283,In_669,In_1248);
or U284 (N_284,In_720,In_629);
xnor U285 (N_285,In_19,In_1890);
nor U286 (N_286,In_1474,In_585);
and U287 (N_287,In_1498,In_1875);
and U288 (N_288,In_16,In_1466);
nor U289 (N_289,In_992,In_201);
xnor U290 (N_290,In_91,In_1979);
and U291 (N_291,In_690,In_424);
and U292 (N_292,In_450,In_1140);
nand U293 (N_293,In_1251,In_142);
nand U294 (N_294,In_609,In_253);
nor U295 (N_295,In_225,In_1814);
nand U296 (N_296,In_1980,In_329);
and U297 (N_297,In_756,In_507);
or U298 (N_298,In_1576,In_1662);
or U299 (N_299,In_1299,In_1786);
and U300 (N_300,In_663,In_630);
nand U301 (N_301,In_301,In_791);
xor U302 (N_302,In_1022,In_1013);
nand U303 (N_303,In_283,In_1289);
nor U304 (N_304,In_1323,In_1927);
nand U305 (N_305,In_1878,In_1769);
or U306 (N_306,In_1545,In_537);
or U307 (N_307,In_1110,In_197);
and U308 (N_308,In_692,In_385);
nor U309 (N_309,In_839,In_1877);
and U310 (N_310,In_746,In_481);
xor U311 (N_311,In_598,In_1057);
nor U312 (N_312,In_1750,In_773);
xnor U313 (N_313,In_1340,In_898);
and U314 (N_314,In_117,In_265);
nor U315 (N_315,In_888,In_624);
nor U316 (N_316,In_1278,In_1211);
and U317 (N_317,In_27,In_133);
nand U318 (N_318,In_1392,In_34);
nor U319 (N_319,In_455,In_901);
nor U320 (N_320,In_1937,In_1004);
nand U321 (N_321,In_167,In_1675);
nand U322 (N_322,In_824,In_1018);
nor U323 (N_323,In_807,In_1771);
xnor U324 (N_324,In_1639,In_540);
nand U325 (N_325,In_1908,In_576);
nand U326 (N_326,In_788,In_993);
and U327 (N_327,In_759,In_211);
nand U328 (N_328,In_792,In_728);
nand U329 (N_329,In_1158,In_556);
nand U330 (N_330,In_395,In_1665);
xnor U331 (N_331,In_1581,In_1388);
nand U332 (N_332,In_1863,In_1680);
and U333 (N_333,In_1703,In_298);
or U334 (N_334,In_1648,In_1546);
nand U335 (N_335,In_518,In_632);
nand U336 (N_336,In_1142,In_113);
and U337 (N_337,In_1520,In_1277);
xor U338 (N_338,In_654,In_1168);
nor U339 (N_339,In_1304,In_1286);
or U340 (N_340,In_1531,In_442);
and U341 (N_341,In_1239,In_658);
or U342 (N_342,In_1058,In_166);
and U343 (N_343,In_1372,In_1650);
xnor U344 (N_344,In_144,In_1002);
nand U345 (N_345,In_1583,In_1341);
or U346 (N_346,In_496,In_1107);
nand U347 (N_347,In_1222,In_228);
or U348 (N_348,In_1941,In_1221);
and U349 (N_349,In_1827,In_353);
nor U350 (N_350,In_376,In_565);
xor U351 (N_351,In_1741,In_1867);
or U352 (N_352,In_1849,In_1862);
nand U353 (N_353,In_1196,In_761);
nand U354 (N_354,In_200,In_1263);
or U355 (N_355,In_1255,In_1717);
or U356 (N_356,In_381,In_943);
nor U357 (N_357,In_704,In_1285);
and U358 (N_358,In_1638,In_814);
or U359 (N_359,In_524,In_1491);
or U360 (N_360,In_338,In_841);
and U361 (N_361,In_1001,In_452);
and U362 (N_362,In_1622,In_1949);
and U363 (N_363,In_1825,In_1620);
nand U364 (N_364,In_1672,In_303);
and U365 (N_365,In_1147,In_165);
nand U366 (N_366,In_503,In_1830);
and U367 (N_367,In_935,In_603);
or U368 (N_368,In_1894,In_714);
or U369 (N_369,In_784,In_492);
nand U370 (N_370,In_621,In_1366);
and U371 (N_371,In_351,In_1189);
xor U372 (N_372,In_1059,In_1907);
and U373 (N_373,In_1842,In_1300);
and U374 (N_374,In_1178,In_1495);
or U375 (N_375,In_176,In_188);
nand U376 (N_376,In_1835,In_1886);
xor U377 (N_377,In_741,In_1358);
nor U378 (N_378,In_1005,In_297);
nor U379 (N_379,In_1625,In_1885);
or U380 (N_380,In_1928,In_1482);
or U381 (N_381,In_1344,In_1096);
and U382 (N_382,In_1062,In_97);
nand U383 (N_383,In_1356,In_1193);
nor U384 (N_384,In_1133,In_1483);
nor U385 (N_385,In_707,In_1777);
and U386 (N_386,In_1081,In_931);
xnor U387 (N_387,In_938,In_1154);
nand U388 (N_388,In_1439,In_1330);
and U389 (N_389,In_828,In_396);
nand U390 (N_390,In_48,In_1785);
nand U391 (N_391,In_465,In_1198);
nand U392 (N_392,In_59,In_1236);
nor U393 (N_393,In_1642,In_108);
and U394 (N_394,In_616,In_870);
or U395 (N_395,In_383,In_1379);
or U396 (N_396,In_1420,In_1365);
nand U397 (N_397,In_13,In_794);
xnor U398 (N_398,In_1353,In_1798);
and U399 (N_399,In_932,In_1393);
nand U400 (N_400,In_331,In_636);
nor U401 (N_401,In_960,In_990);
xor U402 (N_402,In_987,In_1034);
nand U403 (N_403,In_1010,In_1924);
nor U404 (N_404,In_1705,In_1568);
and U405 (N_405,In_1467,In_514);
or U406 (N_406,In_170,In_1846);
xor U407 (N_407,In_6,In_1592);
or U408 (N_408,In_343,In_838);
nand U409 (N_409,In_259,In_693);
and U410 (N_410,In_349,In_251);
or U411 (N_411,In_1203,In_1818);
or U412 (N_412,In_51,In_239);
and U413 (N_413,In_695,In_1295);
nor U414 (N_414,In_758,In_1594);
nor U415 (N_415,In_1117,In_1631);
and U416 (N_416,In_1202,In_422);
nor U417 (N_417,In_189,In_1524);
and U418 (N_418,In_754,In_765);
xor U419 (N_419,In_434,In_662);
nor U420 (N_420,In_547,In_1931);
or U421 (N_421,In_312,In_1819);
nor U422 (N_422,In_1749,In_1318);
and U423 (N_423,In_501,In_665);
or U424 (N_424,In_1471,In_1428);
or U425 (N_425,In_1624,In_1315);
xor U426 (N_426,In_341,In_1120);
and U427 (N_427,In_334,In_1048);
or U428 (N_428,In_377,In_30);
or U429 (N_429,In_1346,In_1293);
or U430 (N_430,In_911,In_84);
and U431 (N_431,In_1561,In_187);
or U432 (N_432,In_130,In_933);
or U433 (N_433,In_240,In_1952);
nand U434 (N_434,In_1730,In_1047);
nor U435 (N_435,In_157,In_1258);
nor U436 (N_436,In_1445,In_1510);
xor U437 (N_437,In_951,In_1829);
xor U438 (N_438,In_104,In_975);
nand U439 (N_439,In_448,In_850);
nand U440 (N_440,In_811,In_886);
xor U441 (N_441,In_656,In_435);
nand U442 (N_442,In_582,In_1386);
and U443 (N_443,In_604,In_1801);
nand U444 (N_444,In_1130,In_640);
nor U445 (N_445,In_666,In_1728);
nor U446 (N_446,In_803,In_1113);
xor U447 (N_447,In_1102,In_1247);
nor U448 (N_448,In_1674,In_1077);
nand U449 (N_449,In_275,In_1369);
nand U450 (N_450,In_1125,In_151);
nor U451 (N_451,In_1914,In_143);
xor U452 (N_452,In_702,In_642);
or U453 (N_453,In_1512,In_1233);
xnor U454 (N_454,In_1453,In_1724);
xnor U455 (N_455,In_318,In_1591);
and U456 (N_456,In_1302,In_1165);
nor U457 (N_457,In_269,In_597);
and U458 (N_458,In_1834,In_516);
nand U459 (N_459,In_1380,In_1569);
nor U460 (N_460,In_1500,In_1045);
and U461 (N_461,In_447,In_449);
nand U462 (N_462,In_719,In_984);
nor U463 (N_463,In_1884,In_1843);
nor U464 (N_464,In_689,In_1570);
nand U465 (N_465,In_266,In_477);
nor U466 (N_466,In_1898,In_775);
nand U467 (N_467,In_671,In_1345);
nand U468 (N_468,In_485,In_348);
nand U469 (N_469,In_1562,In_763);
xnor U470 (N_470,In_149,In_1528);
nand U471 (N_471,In_1422,In_1596);
xnor U472 (N_472,In_1000,In_1430);
nor U473 (N_473,In_1381,In_884);
xnor U474 (N_474,In_875,In_1942);
nor U475 (N_475,In_769,In_140);
and U476 (N_476,In_1099,In_1732);
or U477 (N_477,In_119,In_101);
or U478 (N_478,In_568,In_678);
nand U479 (N_479,In_513,In_1627);
nor U480 (N_480,In_64,In_1993);
xnor U481 (N_481,In_1840,In_1408);
nand U482 (N_482,In_1463,In_1054);
nor U483 (N_483,In_934,In_745);
nor U484 (N_484,In_293,In_1213);
nor U485 (N_485,In_1155,In_192);
nand U486 (N_486,In_534,In_688);
and U487 (N_487,In_1991,In_1401);
or U488 (N_488,In_431,In_487);
nand U489 (N_489,In_522,In_1131);
nand U490 (N_490,In_1906,In_305);
xnor U491 (N_491,In_849,In_186);
nor U492 (N_492,In_1037,In_1873);
nor U493 (N_493,In_1261,In_1114);
xnor U494 (N_494,In_1276,In_1610);
nand U495 (N_495,In_1064,In_172);
nand U496 (N_496,In_1360,In_986);
nor U497 (N_497,In_852,In_757);
nand U498 (N_498,In_1543,In_787);
nor U499 (N_499,In_1160,In_212);
or U500 (N_500,In_1593,In_400);
and U501 (N_501,In_845,In_1313);
nand U502 (N_502,In_1518,In_923);
or U503 (N_503,In_1152,In_1616);
and U504 (N_504,In_1260,In_123);
nor U505 (N_505,In_1267,In_139);
nor U506 (N_506,In_1844,In_25);
and U507 (N_507,In_535,In_1328);
nor U508 (N_508,In_372,In_287);
or U509 (N_509,In_284,In_0);
or U510 (N_510,In_1847,In_1307);
or U511 (N_511,In_198,In_1097);
nand U512 (N_512,In_1493,In_146);
xor U513 (N_513,In_667,In_826);
nand U514 (N_514,In_781,In_1481);
nand U515 (N_515,In_1686,In_752);
nor U516 (N_516,In_1159,In_1820);
nand U517 (N_517,In_1696,In_1563);
and U518 (N_518,In_193,In_958);
or U519 (N_519,In_1962,In_1872);
and U520 (N_520,In_829,In_459);
or U521 (N_521,In_125,In_1632);
xnor U522 (N_522,In_1476,In_1305);
nor U523 (N_523,In_1892,In_1604);
nor U524 (N_524,In_229,In_386);
xnor U525 (N_525,In_1816,In_1416);
and U526 (N_526,In_623,In_1115);
nor U527 (N_527,In_1179,In_109);
nor U528 (N_528,In_1783,In_292);
nor U529 (N_529,In_89,In_767);
or U530 (N_530,In_659,In_1153);
nor U531 (N_531,In_233,In_1522);
and U532 (N_532,In_414,In_1516);
and U533 (N_533,In_1434,In_1431);
or U534 (N_534,In_1575,In_1033);
nand U535 (N_535,In_1689,In_1316);
and U536 (N_536,In_61,In_183);
nand U537 (N_537,In_1659,In_896);
xor U538 (N_538,In_1218,In_627);
and U539 (N_539,In_956,In_1608);
or U540 (N_540,In_926,In_137);
and U541 (N_541,In_1076,In_1683);
nand U542 (N_542,In_1212,In_1707);
nor U543 (N_543,In_65,In_919);
and U544 (N_544,In_128,In_1737);
or U545 (N_545,In_163,In_371);
and U546 (N_546,In_150,In_1633);
nand U547 (N_547,In_285,In_1910);
or U548 (N_548,In_941,In_1139);
or U549 (N_549,In_1138,In_1073);
nand U550 (N_550,In_619,In_1778);
or U551 (N_551,In_1454,In_994);
or U552 (N_552,In_502,In_1241);
nor U553 (N_553,In_1609,In_158);
xor U554 (N_554,In_478,In_1182);
or U555 (N_555,In_1333,In_1879);
nor U556 (N_556,In_397,In_1782);
or U557 (N_557,In_902,In_1209);
nor U558 (N_558,In_242,In_357);
nor U559 (N_559,In_602,In_1363);
nor U560 (N_560,In_380,In_105);
nor U561 (N_561,In_412,In_344);
and U562 (N_562,In_952,In_453);
or U563 (N_563,In_724,In_1228);
xnor U564 (N_564,In_234,In_657);
nand U565 (N_565,In_1967,In_317);
and U566 (N_566,In_482,In_226);
xor U567 (N_567,In_1970,In_408);
xnor U568 (N_568,In_1364,In_723);
nor U569 (N_569,In_844,In_679);
and U570 (N_570,In_1784,In_1028);
nor U571 (N_571,In_610,In_445);
nand U572 (N_572,In_1191,In_1118);
nor U573 (N_573,In_982,In_855);
and U574 (N_574,In_593,In_1322);
and U575 (N_575,In_836,In_914);
and U576 (N_576,In_736,In_121);
nand U577 (N_577,In_804,In_1929);
or U578 (N_578,In_1262,In_43);
and U579 (N_579,In_1111,In_1190);
or U580 (N_580,In_819,In_942);
nor U581 (N_581,In_564,In_299);
or U582 (N_582,In_895,In_1923);
or U583 (N_583,In_1693,In_1042);
and U584 (N_584,In_1797,In_131);
nor U585 (N_585,In_1854,In_468);
nand U586 (N_586,In_126,In_1417);
nand U587 (N_587,In_1201,In_1713);
or U588 (N_588,In_559,In_346);
nand U589 (N_589,In_464,In_1223);
and U590 (N_590,In_1994,In_1035);
nand U591 (N_591,In_1779,In_45);
nor U592 (N_592,In_1501,In_112);
and U593 (N_593,In_573,In_776);
or U594 (N_594,In_1681,In_1803);
nor U595 (N_595,In_1776,In_182);
or U596 (N_596,In_1951,In_1586);
or U597 (N_597,In_1105,In_75);
and U598 (N_598,In_735,In_1853);
and U599 (N_599,In_44,In_517);
or U600 (N_600,In_1470,In_76);
or U601 (N_601,In_1208,In_322);
nor U602 (N_602,In_489,In_1444);
nand U603 (N_603,In_1459,In_833);
or U604 (N_604,In_500,In_1666);
or U605 (N_605,In_637,In_325);
xor U606 (N_606,In_411,In_429);
or U607 (N_607,In_1947,In_1612);
nand U608 (N_608,In_790,In_890);
xor U609 (N_609,In_260,In_1504);
or U610 (N_610,In_419,In_592);
or U611 (N_611,In_1385,In_682);
nor U612 (N_612,In_1815,In_154);
or U613 (N_613,In_1269,In_280);
or U614 (N_614,In_1181,In_1670);
nor U615 (N_615,In_562,In_1508);
nand U616 (N_616,In_9,In_583);
xnor U617 (N_617,In_103,In_296);
nor U618 (N_618,In_179,In_206);
nor U619 (N_619,In_1995,In_155);
or U620 (N_620,In_1172,In_345);
and U621 (N_621,In_1960,In_1515);
or U622 (N_622,In_1817,In_717);
and U623 (N_623,In_575,In_1579);
and U624 (N_624,In_1216,In_370);
or U625 (N_625,In_520,In_107);
or U626 (N_626,In_1109,In_882);
or U627 (N_627,In_972,In_1554);
xnor U628 (N_628,In_1336,In_831);
and U629 (N_629,In_1985,In_925);
nor U630 (N_630,In_1291,In_359);
nor U631 (N_631,In_1903,In_1831);
nor U632 (N_632,In_1311,In_785);
xor U633 (N_633,In_789,In_1394);
nor U634 (N_634,In_1051,In_1377);
nor U635 (N_635,In_796,In_1275);
nor U636 (N_636,In_1597,In_401);
nor U637 (N_637,In_15,In_308);
and U638 (N_638,In_1494,In_1479);
nand U639 (N_639,In_1671,In_53);
and U640 (N_640,In_1425,In_1916);
and U641 (N_641,In_190,In_699);
nand U642 (N_642,In_1100,In_800);
nand U643 (N_643,In_14,In_47);
nand U644 (N_644,In_1857,In_1649);
and U645 (N_645,In_1006,In_997);
or U646 (N_646,In_1171,In_261);
nand U647 (N_647,In_661,In_529);
nor U648 (N_648,In_42,In_272);
nor U649 (N_649,In_913,In_1464);
and U650 (N_650,In_1559,In_1514);
nor U651 (N_651,In_673,In_1414);
or U652 (N_652,In_927,In_1850);
nand U653 (N_653,In_533,In_438);
nand U654 (N_654,In_545,In_404);
xnor U655 (N_655,In_618,In_1940);
nor U656 (N_656,In_1132,In_1888);
and U657 (N_657,In_1134,In_1036);
nand U658 (N_658,In_1462,In_1760);
nand U659 (N_659,In_590,In_969);
or U660 (N_660,In_1564,In_1990);
xnor U661 (N_661,In_885,In_1327);
nand U662 (N_662,In_1584,In_1052);
nor U663 (N_663,In_1447,In_1751);
nand U664 (N_664,In_1661,In_1351);
or U665 (N_665,In_277,In_1104);
or U666 (N_666,In_768,In_649);
xor U667 (N_667,In_389,In_555);
nand U668 (N_668,In_1101,In_497);
or U669 (N_669,In_315,In_423);
and U670 (N_670,In_1558,In_1978);
or U671 (N_671,In_648,In_399);
and U672 (N_672,In_709,In_1436);
or U673 (N_673,In_1489,In_21);
and U674 (N_674,In_379,In_1404);
and U675 (N_675,In_1525,In_23);
and U676 (N_676,In_472,In_1350);
or U677 (N_677,In_1887,In_1572);
and U678 (N_678,In_968,In_1418);
nor U679 (N_679,In_1161,In_622);
or U680 (N_680,In_861,In_1647);
nand U681 (N_681,In_508,In_1136);
nor U682 (N_682,In_771,In_1623);
and U683 (N_683,In_124,In_1095);
nor U684 (N_684,In_906,In_1238);
nor U685 (N_685,In_55,In_446);
nor U686 (N_686,In_1965,In_413);
nor U687 (N_687,In_1992,In_1694);
and U688 (N_688,In_106,In_415);
xor U689 (N_689,In_1082,In_606);
nor U690 (N_690,In_674,In_1296);
nor U691 (N_691,In_696,In_1678);
nand U692 (N_692,In_734,In_250);
or U693 (N_693,In_1981,In_1281);
nand U694 (N_694,In_615,In_1552);
nand U695 (N_695,In_216,In_1743);
and U696 (N_696,In_1192,In_352);
and U697 (N_697,In_505,In_698);
nand U698 (N_698,In_532,In_32);
nand U699 (N_699,In_217,In_1477);
xnor U700 (N_700,In_779,In_1521);
and U701 (N_701,In_1809,In_1590);
or U702 (N_702,In_1253,In_1069);
and U703 (N_703,In_1283,In_209);
nand U704 (N_704,In_484,In_1225);
nand U705 (N_705,In_1698,In_740);
nand U706 (N_706,In_1813,In_162);
nor U707 (N_707,In_69,In_289);
and U708 (N_708,In_1079,In_12);
or U709 (N_709,In_335,In_966);
and U710 (N_710,In_236,In_1009);
and U711 (N_711,In_566,In_1325);
and U712 (N_712,In_1921,In_1950);
nand U713 (N_713,In_1063,In_1718);
nand U714 (N_714,In_1679,In_631);
xnor U715 (N_715,In_1895,In_215);
and U716 (N_716,In_523,In_944);
nor U717 (N_717,In_891,In_417);
nand U718 (N_718,In_286,In_1427);
or U719 (N_719,In_1851,In_1043);
or U720 (N_720,In_1712,In_1688);
nand U721 (N_721,In_1244,In_321);
nand U722 (N_722,In_38,In_1821);
and U723 (N_723,In_1398,In_1621);
or U724 (N_724,In_1072,In_1660);
and U725 (N_725,In_1645,In_780);
nor U726 (N_726,In_920,In_290);
or U727 (N_727,In_980,In_451);
nor U728 (N_728,In_1442,In_1669);
xnor U729 (N_729,In_922,In_1288);
and U730 (N_730,In_410,In_601);
or U731 (N_731,In_147,In_1926);
or U732 (N_732,In_1449,In_1421);
or U733 (N_733,In_672,In_1011);
xor U734 (N_734,In_358,In_708);
or U735 (N_735,In_1837,In_614);
nand U736 (N_736,In_1775,In_644);
xnor U737 (N_737,In_82,In_1026);
nor U738 (N_738,In_1770,In_426);
xor U739 (N_739,In_1440,In_868);
nor U740 (N_740,In_281,In_294);
nand U741 (N_741,In_1429,In_5);
or U742 (N_742,In_244,In_510);
or U743 (N_743,In_731,In_1708);
nor U744 (N_744,In_1763,In_1588);
nor U745 (N_745,In_222,In_1567);
or U746 (N_746,In_1044,In_937);
and U747 (N_747,In_1870,In_806);
or U748 (N_748,In_1988,In_1852);
nor U749 (N_749,In_136,In_1611);
or U750 (N_750,In_1744,In_918);
nand U751 (N_751,In_617,In_1822);
or U752 (N_752,In_1673,In_469);
nand U753 (N_753,In_1395,In_1016);
nor U754 (N_754,In_218,In_1891);
and U755 (N_755,In_1971,In_1413);
or U756 (N_756,In_964,In_655);
or U757 (N_757,In_1589,In_853);
and U758 (N_758,In_506,In_1861);
or U759 (N_759,In_1757,In_1019);
nor U760 (N_760,In_1726,In_1710);
or U761 (N_761,In_1845,In_584);
and U762 (N_762,In_291,In_1764);
or U763 (N_763,In_37,In_940);
xor U764 (N_764,In_457,In_1727);
or U765 (N_765,In_947,In_1571);
nand U766 (N_766,In_892,In_889);
nand U767 (N_767,In_1499,In_1959);
or U768 (N_768,In_307,In_1565);
and U769 (N_769,In_1794,In_1864);
nor U770 (N_770,In_860,In_729);
nand U771 (N_771,In_1505,In_403);
nand U772 (N_772,In_1204,In_1272);
or U773 (N_773,In_701,In_531);
or U774 (N_774,In_1324,In_1424);
nand U775 (N_775,In_1946,In_94);
nand U776 (N_776,In_946,In_1715);
nor U777 (N_777,In_1556,In_1574);
xor U778 (N_778,In_1128,In_1823);
xor U779 (N_779,In_1636,In_262);
or U780 (N_780,In_495,In_425);
nand U781 (N_781,In_1948,In_1112);
and U782 (N_782,In_705,In_786);
nand U783 (N_783,In_454,In_1748);
nor U784 (N_784,In_68,In_132);
nand U785 (N_785,In_1093,In_1008);
nand U786 (N_786,In_1317,In_1480);
nor U787 (N_787,In_586,In_1709);
nand U788 (N_788,In_249,In_894);
nor U789 (N_789,In_1538,In_1643);
xor U790 (N_790,In_596,In_1219);
nand U791 (N_791,In_427,In_751);
nand U792 (N_792,In_1332,In_1426);
nand U793 (N_793,In_406,In_504);
xor U794 (N_794,In_1188,In_1655);
and U795 (N_795,In_360,In_557);
xor U796 (N_796,In_548,In_1535);
nand U797 (N_797,In_530,In_461);
nor U798 (N_798,In_1359,In_921);
or U799 (N_799,In_1969,In_1668);
or U800 (N_800,In_700,In_1373);
or U801 (N_801,In_1932,In_1084);
or U802 (N_802,In_1882,In_1452);
and U803 (N_803,In_1899,In_813);
nand U804 (N_804,In_802,In_96);
nor U805 (N_805,In_1629,In_1530);
and U806 (N_806,In_378,In_801);
or U807 (N_807,In_1517,In_1772);
nand U808 (N_808,In_1415,In_194);
nor U809 (N_809,In_161,In_1331);
and U810 (N_810,In_210,In_1533);
nand U811 (N_811,In_991,In_214);
or U812 (N_812,In_1859,In_1573);
or U813 (N_813,In_1121,In_1297);
or U814 (N_814,In_1031,In_1896);
xnor U815 (N_815,In_1780,In_1021);
xor U816 (N_816,In_175,In_342);
nor U817 (N_817,In_830,In_881);
or U818 (N_818,In_981,In_1540);
nor U819 (N_819,In_549,In_1866);
or U820 (N_820,In_402,In_1930);
xnor U821 (N_821,In_900,In_1214);
nor U822 (N_822,In_842,In_428);
nor U823 (N_823,In_1443,In_1806);
nand U824 (N_824,In_1148,In_985);
and U825 (N_825,In_908,In_1587);
or U826 (N_826,In_1537,In_1721);
nand U827 (N_827,In_1697,In_1376);
or U828 (N_828,In_1826,In_1755);
and U829 (N_829,In_1279,In_1509);
nor U830 (N_830,In_552,In_141);
or U831 (N_831,In_1314,In_939);
or U832 (N_832,In_1465,In_1068);
nand U833 (N_833,In_1066,In_1958);
or U834 (N_834,In_1382,In_1092);
and U835 (N_835,In_1919,In_340);
or U836 (N_836,In_1409,In_877);
or U837 (N_837,In_310,In_493);
nor U838 (N_838,In_169,In_268);
and U839 (N_839,In_1526,In_1361);
or U840 (N_840,In_1685,In_1023);
nor U841 (N_841,In_1150,In_1488);
xor U842 (N_842,In_874,In_1756);
nand U843 (N_843,In_350,In_930);
and U844 (N_844,In_929,In_1682);
xnor U845 (N_845,In_1555,In_726);
or U846 (N_846,In_1687,In_1787);
nand U847 (N_847,In_174,In_706);
xnor U848 (N_848,In_267,In_770);
nand U849 (N_849,In_384,In_1513);
xor U850 (N_850,In_683,In_1175);
and U851 (N_851,In_1654,In_1617);
nor U852 (N_852,In_1765,In_100);
xor U853 (N_853,In_72,In_1618);
nand U854 (N_854,In_1677,In_373);
and U855 (N_855,In_1156,In_899);
or U856 (N_856,In_270,In_70);
nand U857 (N_857,In_703,In_1876);
or U858 (N_858,In_1691,In_1800);
nor U859 (N_859,In_1435,In_815);
nand U860 (N_860,In_1989,In_1539);
nand U861 (N_861,In_1630,In_80);
nand U862 (N_862,In_772,In_1177);
nor U863 (N_863,In_362,In_950);
nand U864 (N_864,In_634,In_1195);
nor U865 (N_865,In_608,In_460);
xnor U866 (N_866,In_300,In_1145);
nand U867 (N_867,In_1953,In_1738);
xnor U868 (N_868,In_820,In_71);
or U869 (N_869,In_1605,In_1734);
nor U870 (N_870,In_466,In_1094);
nor U871 (N_871,In_1487,In_1566);
xnor U872 (N_872,In_1226,In_480);
or U873 (N_873,In_1032,In_1103);
nor U874 (N_874,In_134,In_1412);
xnor U875 (N_875,In_948,In_311);
and U876 (N_876,In_1839,In_288);
nand U877 (N_877,In_650,In_684);
nor U878 (N_878,In_924,In_1472);
nor U879 (N_879,In_1259,In_313);
nor U880 (N_880,In_1560,In_1700);
and U881 (N_881,In_375,In_254);
or U882 (N_882,In_1173,In_546);
xor U883 (N_883,In_967,In_538);
nand U884 (N_884,In_1217,In_737);
nand U885 (N_885,In_1812,In_1074);
or U886 (N_886,In_368,In_1250);
or U887 (N_887,In_594,In_553);
or U888 (N_888,In_799,In_1492);
and U889 (N_889,In_872,In_1141);
xnor U890 (N_890,In_965,In_1231);
and U891 (N_891,In_1913,In_903);
nor U892 (N_892,In_1399,In_86);
or U893 (N_893,In_26,In_1309);
xor U894 (N_894,In_1229,In_54);
and U895 (N_895,In_1264,In_8);
nand U896 (N_896,In_29,In_111);
or U897 (N_897,In_1911,In_612);
nor U898 (N_898,In_1619,In_1603);
or U899 (N_899,In_525,In_1441);
and U900 (N_900,In_1349,In_521);
xnor U901 (N_901,In_645,In_527);
or U902 (N_902,In_430,In_1938);
nor U903 (N_903,In_1602,In_652);
or U904 (N_904,In_40,In_971);
nand U905 (N_905,In_491,In_641);
nor U906 (N_906,In_543,In_742);
nand U907 (N_907,In_279,In_1405);
nand U908 (N_908,In_199,In_1966);
or U909 (N_909,In_1507,In_511);
and U910 (N_910,In_1055,In_1014);
xnor U911 (N_911,In_541,In_1714);
or U912 (N_912,In_1805,In_1220);
nor U913 (N_913,In_1060,In_255);
and U914 (N_914,In_730,In_1027);
nor U915 (N_915,In_1473,In_2);
and U916 (N_916,In_160,In_205);
nor U917 (N_917,In_1496,In_1706);
or U918 (N_918,In_1869,In_1086);
or U919 (N_919,In_988,In_41);
and U920 (N_920,In_1157,In_148);
or U921 (N_921,In_238,In_227);
or U922 (N_922,In_846,In_1070);
nor U923 (N_923,In_996,In_1374);
nand U924 (N_924,In_416,In_1197);
xor U925 (N_925,In_1909,In_865);
nor U926 (N_926,In_764,In_1078);
nor U927 (N_927,In_1151,In_909);
nand U928 (N_928,In_1644,In_1368);
and U929 (N_929,In_1790,In_812);
nand U930 (N_930,In_979,In_1758);
nor U931 (N_931,In_1889,In_1375);
nor U932 (N_932,In_1548,In_1977);
nor U933 (N_933,In_733,In_1793);
nor U934 (N_934,In_713,In_749);
nor U935 (N_935,In_539,In_1091);
or U936 (N_936,In_1390,In_1065);
or U937 (N_937,In_1796,In_1020);
nor U938 (N_938,In_550,In_879);
or U939 (N_939,In_1865,In_52);
and U940 (N_940,In_1087,In_314);
or U941 (N_941,In_366,In_323);
or U942 (N_942,In_1841,In_680);
and U943 (N_943,In_1918,In_1497);
or U944 (N_944,In_832,In_1922);
and U945 (N_945,In_1402,In_1651);
nor U946 (N_946,In_177,In_536);
nand U947 (N_947,In_1207,In_1774);
nand U948 (N_948,In_486,In_156);
nor U949 (N_949,In_479,In_1206);
nand U950 (N_950,In_1652,In_1126);
xnor U951 (N_951,In_18,In_263);
or U952 (N_952,In_727,In_1174);
or U953 (N_953,In_494,In_456);
xor U954 (N_954,In_1598,In_333);
nand U955 (N_955,In_498,In_905);
and U956 (N_956,In_184,In_560);
and U957 (N_957,In_843,In_1944);
or U958 (N_958,In_1637,In_328);
nand U959 (N_959,In_127,In_1729);
nor U960 (N_960,In_977,In_181);
or U961 (N_961,In_1917,In_1747);
and U962 (N_962,In_760,In_1999);
or U963 (N_963,In_488,In_1343);
and U964 (N_964,In_1446,In_88);
or U965 (N_965,In_168,In_1080);
nand U966 (N_966,In_1733,In_114);
and U967 (N_967,In_1029,In_1486);
nor U968 (N_968,In_677,In_1270);
and U969 (N_969,In_1040,In_1003);
nor U970 (N_970,In_1438,In_1407);
or U971 (N_971,In_1731,In_1249);
and U972 (N_972,In_1232,In_17);
or U973 (N_973,In_248,In_571);
or U974 (N_974,In_959,In_1067);
nand U975 (N_975,In_827,In_755);
nand U976 (N_976,In_1667,In_1626);
xor U977 (N_977,In_1968,In_1234);
or U978 (N_978,In_20,In_515);
nand U979 (N_979,In_1646,In_1257);
nand U980 (N_980,In_1553,In_691);
xnor U981 (N_981,In_963,In_1367);
or U982 (N_982,In_462,In_1502);
nand U983 (N_983,In_744,In_1242);
and U984 (N_984,In_1149,In_1742);
nor U985 (N_985,In_1690,In_1303);
nand U986 (N_986,In_1893,In_409);
xor U987 (N_987,In_66,In_1458);
and U988 (N_988,In_1475,In_1945);
nor U989 (N_989,In_676,In_782);
nand U990 (N_990,In_1451,In_1049);
nor U991 (N_991,In_528,In_578);
or U992 (N_992,In_276,In_439);
nor U993 (N_993,In_1972,In_873);
nor U994 (N_994,In_4,In_207);
nand U995 (N_995,In_1056,In_1915);
xnor U996 (N_996,In_369,In_245);
nand U997 (N_997,In_1828,In_195);
and U998 (N_998,In_1860,In_1469);
nand U999 (N_999,In_1389,In_1699);
nand U1000 (N_1000,In_1124,In_973);
nor U1001 (N_1001,In_664,In_491);
and U1002 (N_1002,In_1573,In_1480);
or U1003 (N_1003,In_639,In_975);
or U1004 (N_1004,In_107,In_1442);
nor U1005 (N_1005,In_344,In_50);
and U1006 (N_1006,In_96,In_56);
and U1007 (N_1007,In_1777,In_386);
or U1008 (N_1008,In_807,In_963);
and U1009 (N_1009,In_1716,In_1451);
nor U1010 (N_1010,In_1762,In_986);
and U1011 (N_1011,In_768,In_511);
nand U1012 (N_1012,In_1893,In_1149);
or U1013 (N_1013,In_1052,In_726);
nand U1014 (N_1014,In_1475,In_1348);
nor U1015 (N_1015,In_1800,In_878);
and U1016 (N_1016,In_915,In_1045);
or U1017 (N_1017,In_169,In_456);
and U1018 (N_1018,In_371,In_1829);
nor U1019 (N_1019,In_1863,In_458);
nor U1020 (N_1020,In_130,In_1286);
and U1021 (N_1021,In_583,In_1469);
nor U1022 (N_1022,In_1935,In_800);
and U1023 (N_1023,In_1414,In_1553);
and U1024 (N_1024,In_51,In_1185);
nand U1025 (N_1025,In_1848,In_1425);
and U1026 (N_1026,In_699,In_1649);
and U1027 (N_1027,In_538,In_1446);
nand U1028 (N_1028,In_883,In_1273);
or U1029 (N_1029,In_408,In_1355);
xnor U1030 (N_1030,In_1630,In_1034);
nor U1031 (N_1031,In_1139,In_793);
nor U1032 (N_1032,In_749,In_545);
nor U1033 (N_1033,In_1975,In_524);
and U1034 (N_1034,In_176,In_1225);
nand U1035 (N_1035,In_669,In_1530);
and U1036 (N_1036,In_843,In_330);
or U1037 (N_1037,In_299,In_1550);
nand U1038 (N_1038,In_1035,In_1613);
nand U1039 (N_1039,In_564,In_1533);
nand U1040 (N_1040,In_189,In_979);
nand U1041 (N_1041,In_1573,In_1539);
and U1042 (N_1042,In_1409,In_141);
and U1043 (N_1043,In_1604,In_289);
nor U1044 (N_1044,In_1434,In_28);
nor U1045 (N_1045,In_1694,In_259);
nand U1046 (N_1046,In_1961,In_34);
nand U1047 (N_1047,In_303,In_1963);
nor U1048 (N_1048,In_529,In_1811);
and U1049 (N_1049,In_1317,In_833);
nand U1050 (N_1050,In_67,In_1976);
or U1051 (N_1051,In_18,In_1578);
and U1052 (N_1052,In_1543,In_1407);
nor U1053 (N_1053,In_1795,In_1777);
nor U1054 (N_1054,In_1722,In_222);
or U1055 (N_1055,In_601,In_1224);
xnor U1056 (N_1056,In_1291,In_556);
nor U1057 (N_1057,In_1794,In_1594);
nand U1058 (N_1058,In_1575,In_139);
nor U1059 (N_1059,In_1050,In_823);
or U1060 (N_1060,In_1364,In_231);
and U1061 (N_1061,In_1134,In_142);
xnor U1062 (N_1062,In_1457,In_1675);
xnor U1063 (N_1063,In_728,In_751);
nand U1064 (N_1064,In_1886,In_1731);
nor U1065 (N_1065,In_108,In_806);
and U1066 (N_1066,In_1951,In_1075);
or U1067 (N_1067,In_530,In_1318);
or U1068 (N_1068,In_1814,In_1751);
nand U1069 (N_1069,In_1738,In_1768);
and U1070 (N_1070,In_1724,In_515);
or U1071 (N_1071,In_1565,In_1838);
nand U1072 (N_1072,In_501,In_53);
and U1073 (N_1073,In_1059,In_1078);
nor U1074 (N_1074,In_641,In_860);
and U1075 (N_1075,In_85,In_1269);
and U1076 (N_1076,In_910,In_497);
and U1077 (N_1077,In_234,In_1384);
nor U1078 (N_1078,In_147,In_1707);
or U1079 (N_1079,In_1160,In_1354);
and U1080 (N_1080,In_250,In_1352);
xnor U1081 (N_1081,In_1920,In_431);
nand U1082 (N_1082,In_264,In_1828);
and U1083 (N_1083,In_98,In_1136);
and U1084 (N_1084,In_1710,In_816);
xnor U1085 (N_1085,In_1380,In_498);
nor U1086 (N_1086,In_1934,In_449);
xnor U1087 (N_1087,In_1813,In_940);
xnor U1088 (N_1088,In_1651,In_1469);
xor U1089 (N_1089,In_1487,In_394);
or U1090 (N_1090,In_1921,In_1926);
nor U1091 (N_1091,In_89,In_54);
nand U1092 (N_1092,In_1424,In_1618);
and U1093 (N_1093,In_1552,In_111);
nand U1094 (N_1094,In_608,In_1472);
xnor U1095 (N_1095,In_571,In_1797);
or U1096 (N_1096,In_822,In_1864);
nand U1097 (N_1097,In_1963,In_1514);
nor U1098 (N_1098,In_757,In_989);
or U1099 (N_1099,In_725,In_141);
or U1100 (N_1100,In_322,In_472);
nand U1101 (N_1101,In_1884,In_840);
nor U1102 (N_1102,In_849,In_958);
nand U1103 (N_1103,In_1376,In_322);
nand U1104 (N_1104,In_1845,In_1527);
and U1105 (N_1105,In_1839,In_1290);
and U1106 (N_1106,In_1175,In_1507);
xnor U1107 (N_1107,In_1829,In_1502);
xnor U1108 (N_1108,In_45,In_971);
or U1109 (N_1109,In_554,In_408);
nand U1110 (N_1110,In_398,In_693);
nor U1111 (N_1111,In_1810,In_1203);
and U1112 (N_1112,In_1763,In_57);
nor U1113 (N_1113,In_539,In_615);
or U1114 (N_1114,In_1118,In_775);
or U1115 (N_1115,In_1706,In_1605);
or U1116 (N_1116,In_901,In_1108);
nand U1117 (N_1117,In_345,In_577);
xnor U1118 (N_1118,In_794,In_510);
or U1119 (N_1119,In_1467,In_328);
and U1120 (N_1120,In_1384,In_648);
and U1121 (N_1121,In_1955,In_1599);
xor U1122 (N_1122,In_326,In_1860);
nor U1123 (N_1123,In_142,In_834);
nand U1124 (N_1124,In_1564,In_974);
nand U1125 (N_1125,In_626,In_928);
or U1126 (N_1126,In_1373,In_1931);
and U1127 (N_1127,In_999,In_1267);
and U1128 (N_1128,In_427,In_570);
nand U1129 (N_1129,In_1576,In_804);
xnor U1130 (N_1130,In_1752,In_317);
nand U1131 (N_1131,In_1182,In_813);
or U1132 (N_1132,In_1350,In_1559);
xnor U1133 (N_1133,In_1981,In_1319);
nor U1134 (N_1134,In_1957,In_1161);
nor U1135 (N_1135,In_856,In_443);
nand U1136 (N_1136,In_236,In_1964);
and U1137 (N_1137,In_459,In_1371);
nor U1138 (N_1138,In_107,In_1189);
or U1139 (N_1139,In_58,In_634);
nor U1140 (N_1140,In_744,In_876);
nor U1141 (N_1141,In_1694,In_1145);
nor U1142 (N_1142,In_1295,In_275);
and U1143 (N_1143,In_790,In_1388);
xnor U1144 (N_1144,In_676,In_1318);
and U1145 (N_1145,In_1242,In_1914);
nor U1146 (N_1146,In_422,In_1759);
nand U1147 (N_1147,In_304,In_576);
and U1148 (N_1148,In_724,In_935);
xnor U1149 (N_1149,In_633,In_218);
or U1150 (N_1150,In_350,In_74);
nor U1151 (N_1151,In_958,In_718);
and U1152 (N_1152,In_534,In_458);
or U1153 (N_1153,In_1336,In_1951);
or U1154 (N_1154,In_1738,In_1074);
and U1155 (N_1155,In_933,In_856);
nor U1156 (N_1156,In_470,In_331);
nand U1157 (N_1157,In_640,In_1151);
and U1158 (N_1158,In_1472,In_82);
nor U1159 (N_1159,In_651,In_1123);
nand U1160 (N_1160,In_915,In_882);
nand U1161 (N_1161,In_1171,In_367);
and U1162 (N_1162,In_1754,In_452);
nor U1163 (N_1163,In_1533,In_183);
and U1164 (N_1164,In_1994,In_226);
xor U1165 (N_1165,In_244,In_1494);
nor U1166 (N_1166,In_892,In_1861);
and U1167 (N_1167,In_743,In_1002);
nand U1168 (N_1168,In_462,In_181);
and U1169 (N_1169,In_309,In_936);
or U1170 (N_1170,In_148,In_777);
nor U1171 (N_1171,In_620,In_1231);
xor U1172 (N_1172,In_153,In_1428);
xor U1173 (N_1173,In_1952,In_517);
nor U1174 (N_1174,In_1148,In_878);
nand U1175 (N_1175,In_1390,In_1340);
nand U1176 (N_1176,In_538,In_1040);
and U1177 (N_1177,In_1424,In_841);
nand U1178 (N_1178,In_1921,In_1662);
xor U1179 (N_1179,In_1442,In_861);
or U1180 (N_1180,In_525,In_1108);
nand U1181 (N_1181,In_1824,In_439);
and U1182 (N_1182,In_1553,In_980);
or U1183 (N_1183,In_228,In_1564);
xnor U1184 (N_1184,In_1801,In_1417);
nand U1185 (N_1185,In_1425,In_2);
nor U1186 (N_1186,In_560,In_625);
or U1187 (N_1187,In_627,In_1908);
nor U1188 (N_1188,In_225,In_262);
and U1189 (N_1189,In_188,In_271);
nand U1190 (N_1190,In_1739,In_1400);
nand U1191 (N_1191,In_269,In_1394);
nor U1192 (N_1192,In_280,In_1349);
or U1193 (N_1193,In_299,In_16);
nand U1194 (N_1194,In_1133,In_716);
xnor U1195 (N_1195,In_839,In_602);
or U1196 (N_1196,In_1558,In_1926);
or U1197 (N_1197,In_827,In_1053);
nor U1198 (N_1198,In_1859,In_1913);
or U1199 (N_1199,In_301,In_1432);
nand U1200 (N_1200,In_1790,In_1571);
xor U1201 (N_1201,In_1295,In_1929);
nor U1202 (N_1202,In_1712,In_405);
nor U1203 (N_1203,In_1144,In_512);
nor U1204 (N_1204,In_339,In_1380);
or U1205 (N_1205,In_948,In_117);
or U1206 (N_1206,In_576,In_1680);
nand U1207 (N_1207,In_408,In_1625);
nand U1208 (N_1208,In_753,In_1980);
and U1209 (N_1209,In_1580,In_1250);
nand U1210 (N_1210,In_116,In_557);
nand U1211 (N_1211,In_1161,In_302);
and U1212 (N_1212,In_1544,In_201);
nor U1213 (N_1213,In_49,In_1900);
nor U1214 (N_1214,In_487,In_6);
and U1215 (N_1215,In_1988,In_1575);
nand U1216 (N_1216,In_378,In_234);
nor U1217 (N_1217,In_1400,In_1556);
or U1218 (N_1218,In_1982,In_46);
nor U1219 (N_1219,In_292,In_1023);
and U1220 (N_1220,In_1101,In_1308);
nand U1221 (N_1221,In_1994,In_656);
nand U1222 (N_1222,In_99,In_272);
nand U1223 (N_1223,In_1156,In_831);
nand U1224 (N_1224,In_1489,In_619);
nand U1225 (N_1225,In_1076,In_70);
and U1226 (N_1226,In_298,In_1968);
nand U1227 (N_1227,In_1509,In_633);
xor U1228 (N_1228,In_1668,In_326);
nor U1229 (N_1229,In_1575,In_757);
and U1230 (N_1230,In_1565,In_1164);
xnor U1231 (N_1231,In_1697,In_244);
nand U1232 (N_1232,In_1427,In_807);
and U1233 (N_1233,In_286,In_1787);
or U1234 (N_1234,In_1230,In_1505);
nor U1235 (N_1235,In_977,In_1406);
xnor U1236 (N_1236,In_599,In_349);
nand U1237 (N_1237,In_1160,In_932);
nor U1238 (N_1238,In_1039,In_873);
nand U1239 (N_1239,In_1172,In_1870);
and U1240 (N_1240,In_927,In_197);
nand U1241 (N_1241,In_1602,In_1101);
or U1242 (N_1242,In_126,In_756);
and U1243 (N_1243,In_1120,In_1730);
xor U1244 (N_1244,In_888,In_749);
and U1245 (N_1245,In_920,In_560);
nand U1246 (N_1246,In_69,In_1242);
and U1247 (N_1247,In_274,In_134);
nor U1248 (N_1248,In_1639,In_1311);
nor U1249 (N_1249,In_242,In_1544);
or U1250 (N_1250,In_1037,In_1088);
or U1251 (N_1251,In_1052,In_47);
and U1252 (N_1252,In_438,In_1892);
nor U1253 (N_1253,In_1586,In_1308);
nor U1254 (N_1254,In_502,In_1222);
and U1255 (N_1255,In_1128,In_1705);
and U1256 (N_1256,In_530,In_77);
nand U1257 (N_1257,In_1558,In_1856);
nand U1258 (N_1258,In_1460,In_17);
or U1259 (N_1259,In_190,In_205);
nor U1260 (N_1260,In_1503,In_1247);
and U1261 (N_1261,In_1038,In_1747);
or U1262 (N_1262,In_1649,In_429);
nor U1263 (N_1263,In_874,In_1139);
nor U1264 (N_1264,In_1480,In_130);
and U1265 (N_1265,In_1030,In_523);
nand U1266 (N_1266,In_1461,In_1342);
and U1267 (N_1267,In_1904,In_784);
nand U1268 (N_1268,In_1103,In_1316);
xor U1269 (N_1269,In_435,In_276);
nor U1270 (N_1270,In_1181,In_1024);
or U1271 (N_1271,In_996,In_357);
nor U1272 (N_1272,In_476,In_1113);
nand U1273 (N_1273,In_998,In_1014);
and U1274 (N_1274,In_464,In_929);
or U1275 (N_1275,In_1131,In_743);
nand U1276 (N_1276,In_1326,In_1138);
or U1277 (N_1277,In_161,In_863);
and U1278 (N_1278,In_232,In_1956);
xor U1279 (N_1279,In_1869,In_608);
and U1280 (N_1280,In_1037,In_1925);
or U1281 (N_1281,In_417,In_863);
nor U1282 (N_1282,In_360,In_1688);
xor U1283 (N_1283,In_1653,In_1961);
or U1284 (N_1284,In_980,In_1470);
nand U1285 (N_1285,In_998,In_1328);
nor U1286 (N_1286,In_1758,In_255);
and U1287 (N_1287,In_1798,In_1550);
nand U1288 (N_1288,In_532,In_726);
nand U1289 (N_1289,In_1791,In_647);
or U1290 (N_1290,In_1352,In_62);
nand U1291 (N_1291,In_294,In_905);
nor U1292 (N_1292,In_745,In_344);
and U1293 (N_1293,In_1679,In_1784);
nor U1294 (N_1294,In_1415,In_57);
or U1295 (N_1295,In_853,In_1751);
and U1296 (N_1296,In_1733,In_594);
or U1297 (N_1297,In_237,In_575);
and U1298 (N_1298,In_708,In_714);
nor U1299 (N_1299,In_674,In_877);
or U1300 (N_1300,In_1361,In_1694);
nor U1301 (N_1301,In_1355,In_767);
nand U1302 (N_1302,In_1750,In_1297);
nand U1303 (N_1303,In_1602,In_1583);
xnor U1304 (N_1304,In_791,In_1523);
nand U1305 (N_1305,In_1908,In_662);
nor U1306 (N_1306,In_104,In_408);
nor U1307 (N_1307,In_107,In_1678);
or U1308 (N_1308,In_630,In_885);
xor U1309 (N_1309,In_1647,In_1581);
nand U1310 (N_1310,In_1075,In_1083);
and U1311 (N_1311,In_275,In_849);
and U1312 (N_1312,In_284,In_1333);
and U1313 (N_1313,In_167,In_975);
nor U1314 (N_1314,In_178,In_849);
nor U1315 (N_1315,In_435,In_1772);
and U1316 (N_1316,In_401,In_305);
xor U1317 (N_1317,In_1575,In_518);
or U1318 (N_1318,In_1884,In_1463);
nand U1319 (N_1319,In_1606,In_249);
xor U1320 (N_1320,In_1340,In_1792);
and U1321 (N_1321,In_428,In_1606);
or U1322 (N_1322,In_1525,In_1363);
and U1323 (N_1323,In_90,In_1864);
nor U1324 (N_1324,In_1080,In_1523);
nor U1325 (N_1325,In_243,In_673);
xor U1326 (N_1326,In_735,In_1580);
xor U1327 (N_1327,In_43,In_1936);
and U1328 (N_1328,In_1080,In_603);
and U1329 (N_1329,In_1232,In_1539);
or U1330 (N_1330,In_1453,In_342);
or U1331 (N_1331,In_1462,In_430);
nor U1332 (N_1332,In_905,In_1401);
xor U1333 (N_1333,In_1271,In_1643);
and U1334 (N_1334,In_1168,In_109);
nand U1335 (N_1335,In_229,In_380);
nor U1336 (N_1336,In_1836,In_941);
or U1337 (N_1337,In_449,In_1035);
nand U1338 (N_1338,In_78,In_164);
nor U1339 (N_1339,In_631,In_1388);
or U1340 (N_1340,In_902,In_1929);
or U1341 (N_1341,In_1385,In_741);
nor U1342 (N_1342,In_1670,In_1085);
xnor U1343 (N_1343,In_1860,In_725);
nand U1344 (N_1344,In_1325,In_1836);
and U1345 (N_1345,In_1493,In_377);
or U1346 (N_1346,In_1602,In_1820);
and U1347 (N_1347,In_392,In_408);
nor U1348 (N_1348,In_607,In_1485);
xor U1349 (N_1349,In_1693,In_932);
and U1350 (N_1350,In_52,In_327);
xor U1351 (N_1351,In_588,In_1099);
nor U1352 (N_1352,In_20,In_543);
and U1353 (N_1353,In_744,In_1270);
nand U1354 (N_1354,In_1552,In_1722);
nor U1355 (N_1355,In_537,In_680);
and U1356 (N_1356,In_525,In_650);
nor U1357 (N_1357,In_441,In_839);
and U1358 (N_1358,In_1170,In_427);
and U1359 (N_1359,In_773,In_754);
and U1360 (N_1360,In_1785,In_356);
nor U1361 (N_1361,In_273,In_49);
or U1362 (N_1362,In_1157,In_758);
or U1363 (N_1363,In_229,In_991);
and U1364 (N_1364,In_994,In_1760);
or U1365 (N_1365,In_658,In_1231);
or U1366 (N_1366,In_1869,In_351);
or U1367 (N_1367,In_1531,In_976);
nor U1368 (N_1368,In_301,In_290);
and U1369 (N_1369,In_93,In_543);
or U1370 (N_1370,In_1262,In_1224);
nor U1371 (N_1371,In_1848,In_1339);
nor U1372 (N_1372,In_1248,In_1996);
nor U1373 (N_1373,In_1300,In_889);
and U1374 (N_1374,In_1095,In_1768);
and U1375 (N_1375,In_647,In_275);
nand U1376 (N_1376,In_777,In_963);
nor U1377 (N_1377,In_1146,In_1835);
nor U1378 (N_1378,In_389,In_1686);
or U1379 (N_1379,In_829,In_1842);
nor U1380 (N_1380,In_1576,In_476);
and U1381 (N_1381,In_83,In_1739);
xnor U1382 (N_1382,In_287,In_1670);
or U1383 (N_1383,In_1367,In_1295);
or U1384 (N_1384,In_1443,In_28);
nor U1385 (N_1385,In_1387,In_810);
or U1386 (N_1386,In_1490,In_1562);
nand U1387 (N_1387,In_341,In_703);
nor U1388 (N_1388,In_1597,In_1632);
nor U1389 (N_1389,In_66,In_557);
xnor U1390 (N_1390,In_364,In_36);
or U1391 (N_1391,In_1590,In_643);
nand U1392 (N_1392,In_784,In_1203);
nand U1393 (N_1393,In_1843,In_827);
or U1394 (N_1394,In_243,In_744);
nand U1395 (N_1395,In_457,In_1471);
nand U1396 (N_1396,In_198,In_1080);
nor U1397 (N_1397,In_1119,In_311);
nor U1398 (N_1398,In_1435,In_1455);
nor U1399 (N_1399,In_230,In_1712);
and U1400 (N_1400,In_742,In_1923);
xnor U1401 (N_1401,In_331,In_1467);
or U1402 (N_1402,In_1054,In_379);
nor U1403 (N_1403,In_1082,In_1861);
nand U1404 (N_1404,In_1850,In_1925);
or U1405 (N_1405,In_925,In_565);
and U1406 (N_1406,In_1748,In_1932);
and U1407 (N_1407,In_31,In_1624);
nor U1408 (N_1408,In_436,In_1571);
nand U1409 (N_1409,In_231,In_475);
or U1410 (N_1410,In_1809,In_1026);
xnor U1411 (N_1411,In_1478,In_1241);
or U1412 (N_1412,In_636,In_526);
nand U1413 (N_1413,In_429,In_1275);
nand U1414 (N_1414,In_1738,In_615);
xor U1415 (N_1415,In_1980,In_1172);
nor U1416 (N_1416,In_919,In_1641);
xnor U1417 (N_1417,In_1451,In_441);
nand U1418 (N_1418,In_821,In_1835);
or U1419 (N_1419,In_1785,In_1033);
and U1420 (N_1420,In_1541,In_617);
and U1421 (N_1421,In_1861,In_267);
and U1422 (N_1422,In_1562,In_1602);
xor U1423 (N_1423,In_177,In_1684);
or U1424 (N_1424,In_1724,In_1305);
or U1425 (N_1425,In_210,In_259);
or U1426 (N_1426,In_910,In_1340);
or U1427 (N_1427,In_61,In_1648);
nor U1428 (N_1428,In_400,In_1762);
and U1429 (N_1429,In_1564,In_835);
and U1430 (N_1430,In_848,In_1558);
or U1431 (N_1431,In_1455,In_267);
nand U1432 (N_1432,In_489,In_874);
xnor U1433 (N_1433,In_620,In_614);
nor U1434 (N_1434,In_1138,In_515);
or U1435 (N_1435,In_1142,In_74);
or U1436 (N_1436,In_653,In_720);
nand U1437 (N_1437,In_430,In_86);
xor U1438 (N_1438,In_424,In_267);
nand U1439 (N_1439,In_1844,In_1585);
xor U1440 (N_1440,In_1966,In_1542);
nand U1441 (N_1441,In_1257,In_1509);
and U1442 (N_1442,In_1477,In_644);
and U1443 (N_1443,In_59,In_1897);
nand U1444 (N_1444,In_1269,In_996);
or U1445 (N_1445,In_1710,In_323);
or U1446 (N_1446,In_118,In_1454);
or U1447 (N_1447,In_1979,In_460);
nand U1448 (N_1448,In_1438,In_428);
nand U1449 (N_1449,In_1897,In_1997);
xnor U1450 (N_1450,In_1766,In_788);
nand U1451 (N_1451,In_1347,In_1316);
nor U1452 (N_1452,In_748,In_705);
or U1453 (N_1453,In_66,In_1215);
and U1454 (N_1454,In_163,In_29);
xor U1455 (N_1455,In_447,In_1814);
or U1456 (N_1456,In_1238,In_1007);
nor U1457 (N_1457,In_1680,In_1521);
nand U1458 (N_1458,In_1414,In_285);
nand U1459 (N_1459,In_1231,In_1013);
or U1460 (N_1460,In_415,In_827);
nand U1461 (N_1461,In_696,In_1276);
or U1462 (N_1462,In_831,In_846);
nor U1463 (N_1463,In_995,In_872);
nand U1464 (N_1464,In_593,In_1258);
nand U1465 (N_1465,In_1333,In_215);
nor U1466 (N_1466,In_694,In_1127);
and U1467 (N_1467,In_1318,In_1305);
nand U1468 (N_1468,In_1332,In_1736);
xor U1469 (N_1469,In_606,In_251);
and U1470 (N_1470,In_1307,In_701);
and U1471 (N_1471,In_1464,In_1769);
nor U1472 (N_1472,In_1821,In_326);
and U1473 (N_1473,In_1660,In_1509);
and U1474 (N_1474,In_1262,In_1978);
or U1475 (N_1475,In_1741,In_345);
and U1476 (N_1476,In_1762,In_1313);
or U1477 (N_1477,In_1013,In_1241);
or U1478 (N_1478,In_1106,In_1067);
nand U1479 (N_1479,In_1385,In_1618);
xor U1480 (N_1480,In_289,In_1262);
or U1481 (N_1481,In_1581,In_1618);
nand U1482 (N_1482,In_258,In_83);
nand U1483 (N_1483,In_1345,In_1539);
or U1484 (N_1484,In_983,In_464);
or U1485 (N_1485,In_433,In_28);
and U1486 (N_1486,In_1582,In_1445);
xor U1487 (N_1487,In_1362,In_645);
nand U1488 (N_1488,In_1223,In_1709);
and U1489 (N_1489,In_1874,In_219);
or U1490 (N_1490,In_1285,In_625);
or U1491 (N_1491,In_1899,In_1303);
nand U1492 (N_1492,In_318,In_1472);
nor U1493 (N_1493,In_1517,In_1764);
nand U1494 (N_1494,In_162,In_630);
nand U1495 (N_1495,In_894,In_1852);
and U1496 (N_1496,In_131,In_134);
xor U1497 (N_1497,In_1376,In_724);
nor U1498 (N_1498,In_1861,In_1352);
or U1499 (N_1499,In_295,In_1308);
nand U1500 (N_1500,In_1057,In_1839);
nand U1501 (N_1501,In_462,In_1105);
and U1502 (N_1502,In_349,In_436);
nand U1503 (N_1503,In_897,In_1186);
nand U1504 (N_1504,In_1096,In_263);
or U1505 (N_1505,In_488,In_1002);
nor U1506 (N_1506,In_1062,In_1434);
xnor U1507 (N_1507,In_1706,In_607);
and U1508 (N_1508,In_876,In_605);
or U1509 (N_1509,In_1414,In_377);
nor U1510 (N_1510,In_31,In_365);
xor U1511 (N_1511,In_601,In_2);
nand U1512 (N_1512,In_485,In_1829);
and U1513 (N_1513,In_983,In_1860);
nor U1514 (N_1514,In_98,In_1652);
nand U1515 (N_1515,In_654,In_429);
and U1516 (N_1516,In_912,In_108);
nor U1517 (N_1517,In_1113,In_615);
and U1518 (N_1518,In_1241,In_51);
or U1519 (N_1519,In_614,In_1333);
and U1520 (N_1520,In_698,In_1142);
or U1521 (N_1521,In_1080,In_1878);
nor U1522 (N_1522,In_390,In_1742);
and U1523 (N_1523,In_1223,In_877);
nand U1524 (N_1524,In_1257,In_1012);
xor U1525 (N_1525,In_586,In_261);
nor U1526 (N_1526,In_1595,In_1945);
nand U1527 (N_1527,In_107,In_383);
and U1528 (N_1528,In_143,In_1097);
nor U1529 (N_1529,In_1114,In_1407);
and U1530 (N_1530,In_336,In_1899);
nand U1531 (N_1531,In_1780,In_399);
or U1532 (N_1532,In_742,In_26);
nand U1533 (N_1533,In_916,In_1806);
nand U1534 (N_1534,In_207,In_609);
xor U1535 (N_1535,In_177,In_104);
and U1536 (N_1536,In_1539,In_1572);
nor U1537 (N_1537,In_1190,In_1394);
and U1538 (N_1538,In_431,In_1037);
nand U1539 (N_1539,In_1203,In_794);
or U1540 (N_1540,In_683,In_69);
or U1541 (N_1541,In_1425,In_1179);
xnor U1542 (N_1542,In_1263,In_59);
nor U1543 (N_1543,In_1814,In_407);
nor U1544 (N_1544,In_608,In_837);
xor U1545 (N_1545,In_859,In_1617);
nand U1546 (N_1546,In_1652,In_1157);
and U1547 (N_1547,In_1419,In_848);
nor U1548 (N_1548,In_1732,In_1611);
nand U1549 (N_1549,In_1430,In_1278);
and U1550 (N_1550,In_1854,In_111);
nor U1551 (N_1551,In_260,In_837);
nor U1552 (N_1552,In_1773,In_179);
xor U1553 (N_1553,In_71,In_1715);
nand U1554 (N_1554,In_774,In_1415);
and U1555 (N_1555,In_1536,In_56);
or U1556 (N_1556,In_452,In_990);
nand U1557 (N_1557,In_1490,In_989);
xor U1558 (N_1558,In_632,In_309);
nor U1559 (N_1559,In_447,In_1599);
xnor U1560 (N_1560,In_1536,In_175);
nand U1561 (N_1561,In_1617,In_1180);
and U1562 (N_1562,In_1897,In_1718);
nor U1563 (N_1563,In_25,In_935);
nor U1564 (N_1564,In_1143,In_1508);
or U1565 (N_1565,In_404,In_184);
xor U1566 (N_1566,In_13,In_177);
xnor U1567 (N_1567,In_1400,In_30);
nand U1568 (N_1568,In_1705,In_1516);
nand U1569 (N_1569,In_1167,In_701);
nand U1570 (N_1570,In_1392,In_1608);
nand U1571 (N_1571,In_1041,In_1136);
or U1572 (N_1572,In_475,In_347);
nand U1573 (N_1573,In_777,In_1650);
or U1574 (N_1574,In_157,In_487);
and U1575 (N_1575,In_1763,In_770);
xor U1576 (N_1576,In_883,In_52);
nand U1577 (N_1577,In_1088,In_930);
nand U1578 (N_1578,In_1470,In_924);
and U1579 (N_1579,In_701,In_1654);
or U1580 (N_1580,In_959,In_737);
nand U1581 (N_1581,In_604,In_1286);
and U1582 (N_1582,In_1993,In_1091);
or U1583 (N_1583,In_767,In_618);
nand U1584 (N_1584,In_1630,In_1706);
or U1585 (N_1585,In_1856,In_766);
nor U1586 (N_1586,In_1718,In_1108);
nand U1587 (N_1587,In_735,In_591);
nor U1588 (N_1588,In_677,In_397);
or U1589 (N_1589,In_1773,In_787);
and U1590 (N_1590,In_423,In_1905);
or U1591 (N_1591,In_1599,In_1071);
and U1592 (N_1592,In_1195,In_561);
or U1593 (N_1593,In_394,In_724);
nand U1594 (N_1594,In_1601,In_464);
and U1595 (N_1595,In_1557,In_266);
or U1596 (N_1596,In_886,In_1964);
nand U1597 (N_1597,In_1688,In_1349);
xor U1598 (N_1598,In_969,In_1027);
nor U1599 (N_1599,In_1614,In_939);
or U1600 (N_1600,In_46,In_1156);
or U1601 (N_1601,In_1767,In_1577);
nor U1602 (N_1602,In_1935,In_405);
and U1603 (N_1603,In_1116,In_510);
nor U1604 (N_1604,In_1093,In_813);
nor U1605 (N_1605,In_905,In_146);
xor U1606 (N_1606,In_1051,In_1063);
nand U1607 (N_1607,In_704,In_777);
nand U1608 (N_1608,In_650,In_1608);
nand U1609 (N_1609,In_746,In_263);
xor U1610 (N_1610,In_1557,In_1198);
and U1611 (N_1611,In_1019,In_400);
nor U1612 (N_1612,In_1495,In_722);
or U1613 (N_1613,In_908,In_197);
nand U1614 (N_1614,In_492,In_589);
nand U1615 (N_1615,In_1920,In_314);
nand U1616 (N_1616,In_1885,In_412);
or U1617 (N_1617,In_171,In_1003);
nor U1618 (N_1618,In_1783,In_1202);
nand U1619 (N_1619,In_856,In_233);
and U1620 (N_1620,In_1753,In_1842);
nor U1621 (N_1621,In_1861,In_1875);
nor U1622 (N_1622,In_1209,In_611);
nand U1623 (N_1623,In_292,In_1290);
nand U1624 (N_1624,In_1794,In_1821);
nor U1625 (N_1625,In_1394,In_1884);
or U1626 (N_1626,In_1941,In_1176);
nor U1627 (N_1627,In_960,In_172);
xnor U1628 (N_1628,In_1732,In_885);
xor U1629 (N_1629,In_429,In_1540);
xnor U1630 (N_1630,In_1401,In_445);
and U1631 (N_1631,In_608,In_1768);
or U1632 (N_1632,In_410,In_1593);
nand U1633 (N_1633,In_877,In_915);
nand U1634 (N_1634,In_1327,In_1662);
or U1635 (N_1635,In_1428,In_462);
and U1636 (N_1636,In_1614,In_397);
nor U1637 (N_1637,In_666,In_1202);
and U1638 (N_1638,In_471,In_442);
nand U1639 (N_1639,In_1587,In_260);
nor U1640 (N_1640,In_181,In_210);
nand U1641 (N_1641,In_1624,In_1280);
nor U1642 (N_1642,In_561,In_942);
nor U1643 (N_1643,In_297,In_517);
and U1644 (N_1644,In_1110,In_1049);
nand U1645 (N_1645,In_955,In_241);
nand U1646 (N_1646,In_1577,In_328);
and U1647 (N_1647,In_231,In_208);
nor U1648 (N_1648,In_185,In_1471);
nand U1649 (N_1649,In_1293,In_1599);
or U1650 (N_1650,In_150,In_656);
nor U1651 (N_1651,In_1056,In_681);
nor U1652 (N_1652,In_587,In_1299);
or U1653 (N_1653,In_1207,In_1551);
and U1654 (N_1654,In_89,In_1596);
nand U1655 (N_1655,In_1776,In_107);
nand U1656 (N_1656,In_1726,In_1296);
nor U1657 (N_1657,In_978,In_1776);
nand U1658 (N_1658,In_1462,In_838);
nand U1659 (N_1659,In_1635,In_436);
nand U1660 (N_1660,In_1514,In_1768);
nor U1661 (N_1661,In_1173,In_1615);
and U1662 (N_1662,In_1302,In_186);
nand U1663 (N_1663,In_371,In_38);
nor U1664 (N_1664,In_892,In_958);
nand U1665 (N_1665,In_723,In_880);
nor U1666 (N_1666,In_420,In_1860);
nor U1667 (N_1667,In_445,In_1547);
or U1668 (N_1668,In_223,In_751);
nand U1669 (N_1669,In_1748,In_1492);
nor U1670 (N_1670,In_1095,In_520);
nor U1671 (N_1671,In_1731,In_1954);
nand U1672 (N_1672,In_483,In_229);
and U1673 (N_1673,In_1827,In_1758);
nand U1674 (N_1674,In_551,In_451);
or U1675 (N_1675,In_1267,In_72);
nor U1676 (N_1676,In_790,In_1751);
and U1677 (N_1677,In_316,In_1576);
nor U1678 (N_1678,In_565,In_1155);
xor U1679 (N_1679,In_357,In_1361);
and U1680 (N_1680,In_1134,In_67);
or U1681 (N_1681,In_291,In_1146);
nand U1682 (N_1682,In_321,In_1919);
and U1683 (N_1683,In_1490,In_1997);
or U1684 (N_1684,In_1652,In_1429);
or U1685 (N_1685,In_312,In_1406);
and U1686 (N_1686,In_102,In_1993);
and U1687 (N_1687,In_1926,In_1563);
nor U1688 (N_1688,In_1833,In_998);
xor U1689 (N_1689,In_114,In_791);
or U1690 (N_1690,In_1066,In_622);
nand U1691 (N_1691,In_905,In_487);
nand U1692 (N_1692,In_126,In_668);
nor U1693 (N_1693,In_1143,In_1662);
and U1694 (N_1694,In_1495,In_819);
and U1695 (N_1695,In_1242,In_189);
nor U1696 (N_1696,In_1946,In_924);
nand U1697 (N_1697,In_1375,In_1041);
nor U1698 (N_1698,In_1872,In_1098);
nor U1699 (N_1699,In_942,In_258);
xnor U1700 (N_1700,In_22,In_1570);
and U1701 (N_1701,In_1248,In_671);
xnor U1702 (N_1702,In_1650,In_348);
nand U1703 (N_1703,In_593,In_79);
or U1704 (N_1704,In_316,In_1118);
nand U1705 (N_1705,In_1209,In_224);
or U1706 (N_1706,In_136,In_1502);
nand U1707 (N_1707,In_215,In_291);
or U1708 (N_1708,In_1349,In_316);
nand U1709 (N_1709,In_1352,In_1378);
and U1710 (N_1710,In_800,In_481);
nor U1711 (N_1711,In_1030,In_598);
or U1712 (N_1712,In_1787,In_1989);
and U1713 (N_1713,In_209,In_1984);
or U1714 (N_1714,In_1102,In_626);
nand U1715 (N_1715,In_355,In_1234);
or U1716 (N_1716,In_1180,In_1683);
nor U1717 (N_1717,In_1089,In_1529);
nand U1718 (N_1718,In_746,In_749);
and U1719 (N_1719,In_716,In_1819);
nor U1720 (N_1720,In_1005,In_1339);
nand U1721 (N_1721,In_286,In_203);
nand U1722 (N_1722,In_1736,In_1756);
and U1723 (N_1723,In_509,In_1767);
nand U1724 (N_1724,In_660,In_748);
and U1725 (N_1725,In_1910,In_554);
nor U1726 (N_1726,In_1089,In_1266);
nand U1727 (N_1727,In_1541,In_337);
and U1728 (N_1728,In_493,In_463);
and U1729 (N_1729,In_150,In_1031);
nor U1730 (N_1730,In_1865,In_1042);
xnor U1731 (N_1731,In_709,In_1094);
and U1732 (N_1732,In_203,In_155);
or U1733 (N_1733,In_1977,In_444);
or U1734 (N_1734,In_438,In_1495);
nand U1735 (N_1735,In_971,In_1191);
and U1736 (N_1736,In_1908,In_10);
xnor U1737 (N_1737,In_862,In_1025);
nor U1738 (N_1738,In_431,In_1152);
xor U1739 (N_1739,In_1307,In_1128);
or U1740 (N_1740,In_1462,In_378);
and U1741 (N_1741,In_624,In_495);
nand U1742 (N_1742,In_1945,In_1662);
xnor U1743 (N_1743,In_1327,In_727);
xor U1744 (N_1744,In_225,In_1713);
nor U1745 (N_1745,In_355,In_1517);
nand U1746 (N_1746,In_196,In_562);
nand U1747 (N_1747,In_1753,In_470);
nor U1748 (N_1748,In_857,In_142);
and U1749 (N_1749,In_1859,In_1057);
nor U1750 (N_1750,In_1698,In_714);
and U1751 (N_1751,In_626,In_608);
nor U1752 (N_1752,In_1959,In_141);
nand U1753 (N_1753,In_1,In_624);
nand U1754 (N_1754,In_1637,In_1421);
nor U1755 (N_1755,In_479,In_1533);
or U1756 (N_1756,In_940,In_1871);
and U1757 (N_1757,In_868,In_147);
nand U1758 (N_1758,In_1441,In_1149);
or U1759 (N_1759,In_1897,In_603);
and U1760 (N_1760,In_1945,In_1593);
nand U1761 (N_1761,In_1065,In_1469);
xnor U1762 (N_1762,In_1308,In_182);
and U1763 (N_1763,In_932,In_1989);
and U1764 (N_1764,In_1694,In_482);
nor U1765 (N_1765,In_655,In_1918);
or U1766 (N_1766,In_1101,In_52);
or U1767 (N_1767,In_818,In_1811);
nor U1768 (N_1768,In_681,In_1548);
or U1769 (N_1769,In_1208,In_1364);
or U1770 (N_1770,In_1334,In_1782);
nand U1771 (N_1771,In_1947,In_274);
nor U1772 (N_1772,In_993,In_115);
and U1773 (N_1773,In_1388,In_1895);
nand U1774 (N_1774,In_1066,In_446);
xor U1775 (N_1775,In_892,In_1746);
nor U1776 (N_1776,In_149,In_855);
or U1777 (N_1777,In_1532,In_1715);
and U1778 (N_1778,In_654,In_800);
nor U1779 (N_1779,In_173,In_525);
nor U1780 (N_1780,In_1559,In_433);
or U1781 (N_1781,In_1722,In_822);
and U1782 (N_1782,In_329,In_949);
and U1783 (N_1783,In_548,In_1235);
or U1784 (N_1784,In_1245,In_1515);
nor U1785 (N_1785,In_647,In_987);
nor U1786 (N_1786,In_1190,In_399);
and U1787 (N_1787,In_1085,In_199);
nand U1788 (N_1788,In_394,In_1395);
nand U1789 (N_1789,In_1159,In_1104);
xor U1790 (N_1790,In_770,In_1610);
or U1791 (N_1791,In_316,In_906);
nand U1792 (N_1792,In_215,In_406);
nand U1793 (N_1793,In_1174,In_1380);
and U1794 (N_1794,In_1297,In_645);
nor U1795 (N_1795,In_902,In_1510);
xnor U1796 (N_1796,In_1408,In_1618);
nand U1797 (N_1797,In_167,In_1542);
or U1798 (N_1798,In_1307,In_273);
nor U1799 (N_1799,In_548,In_648);
or U1800 (N_1800,In_1945,In_1447);
nand U1801 (N_1801,In_340,In_482);
nand U1802 (N_1802,In_1118,In_697);
or U1803 (N_1803,In_310,In_974);
and U1804 (N_1804,In_1797,In_958);
nor U1805 (N_1805,In_716,In_1000);
nor U1806 (N_1806,In_1644,In_206);
nand U1807 (N_1807,In_622,In_527);
nor U1808 (N_1808,In_35,In_720);
nand U1809 (N_1809,In_617,In_533);
and U1810 (N_1810,In_1950,In_1375);
or U1811 (N_1811,In_1630,In_1123);
or U1812 (N_1812,In_894,In_1254);
or U1813 (N_1813,In_675,In_422);
nor U1814 (N_1814,In_205,In_1917);
or U1815 (N_1815,In_606,In_1345);
or U1816 (N_1816,In_1527,In_89);
nor U1817 (N_1817,In_310,In_1176);
nand U1818 (N_1818,In_394,In_1656);
and U1819 (N_1819,In_567,In_1333);
nor U1820 (N_1820,In_799,In_1092);
and U1821 (N_1821,In_677,In_1094);
nand U1822 (N_1822,In_845,In_408);
or U1823 (N_1823,In_1506,In_100);
and U1824 (N_1824,In_1490,In_869);
nand U1825 (N_1825,In_1890,In_1601);
and U1826 (N_1826,In_1033,In_1812);
xor U1827 (N_1827,In_1820,In_414);
or U1828 (N_1828,In_1925,In_1195);
nand U1829 (N_1829,In_1888,In_791);
or U1830 (N_1830,In_699,In_62);
or U1831 (N_1831,In_1654,In_1491);
and U1832 (N_1832,In_498,In_1437);
nor U1833 (N_1833,In_1427,In_94);
nand U1834 (N_1834,In_682,In_749);
or U1835 (N_1835,In_1203,In_246);
nor U1836 (N_1836,In_1862,In_1475);
xnor U1837 (N_1837,In_1112,In_1161);
and U1838 (N_1838,In_292,In_1693);
and U1839 (N_1839,In_535,In_623);
and U1840 (N_1840,In_875,In_245);
or U1841 (N_1841,In_117,In_1211);
nor U1842 (N_1842,In_543,In_685);
or U1843 (N_1843,In_1444,In_1689);
nand U1844 (N_1844,In_76,In_488);
xnor U1845 (N_1845,In_580,In_1289);
and U1846 (N_1846,In_482,In_945);
nand U1847 (N_1847,In_121,In_899);
nand U1848 (N_1848,In_1999,In_1837);
nand U1849 (N_1849,In_502,In_808);
or U1850 (N_1850,In_530,In_31);
nand U1851 (N_1851,In_813,In_1739);
and U1852 (N_1852,In_788,In_1948);
or U1853 (N_1853,In_472,In_1071);
nand U1854 (N_1854,In_356,In_1014);
nor U1855 (N_1855,In_1995,In_1635);
nand U1856 (N_1856,In_462,In_1202);
and U1857 (N_1857,In_227,In_1048);
nor U1858 (N_1858,In_22,In_470);
or U1859 (N_1859,In_1213,In_564);
or U1860 (N_1860,In_1655,In_856);
nor U1861 (N_1861,In_1467,In_561);
and U1862 (N_1862,In_21,In_1685);
or U1863 (N_1863,In_146,In_920);
or U1864 (N_1864,In_1481,In_323);
nand U1865 (N_1865,In_1563,In_413);
nand U1866 (N_1866,In_1669,In_215);
nor U1867 (N_1867,In_1457,In_1100);
and U1868 (N_1868,In_625,In_1649);
xor U1869 (N_1869,In_271,In_1918);
or U1870 (N_1870,In_1241,In_1069);
nand U1871 (N_1871,In_1022,In_801);
xor U1872 (N_1872,In_1015,In_449);
xor U1873 (N_1873,In_641,In_958);
or U1874 (N_1874,In_1560,In_746);
or U1875 (N_1875,In_661,In_1896);
and U1876 (N_1876,In_1909,In_1131);
xor U1877 (N_1877,In_306,In_259);
nor U1878 (N_1878,In_1161,In_432);
or U1879 (N_1879,In_1998,In_38);
xnor U1880 (N_1880,In_1501,In_574);
nand U1881 (N_1881,In_1756,In_299);
or U1882 (N_1882,In_521,In_345);
nor U1883 (N_1883,In_1780,In_895);
nand U1884 (N_1884,In_1177,In_1290);
nand U1885 (N_1885,In_15,In_1339);
and U1886 (N_1886,In_9,In_395);
and U1887 (N_1887,In_1984,In_262);
nand U1888 (N_1888,In_1677,In_1195);
or U1889 (N_1889,In_264,In_1024);
xnor U1890 (N_1890,In_1261,In_1634);
xor U1891 (N_1891,In_1531,In_617);
xnor U1892 (N_1892,In_610,In_1426);
or U1893 (N_1893,In_462,In_651);
or U1894 (N_1894,In_1274,In_1723);
nor U1895 (N_1895,In_1732,In_595);
or U1896 (N_1896,In_1340,In_647);
and U1897 (N_1897,In_1506,In_563);
and U1898 (N_1898,In_1554,In_614);
and U1899 (N_1899,In_1912,In_116);
or U1900 (N_1900,In_1862,In_431);
or U1901 (N_1901,In_339,In_1543);
or U1902 (N_1902,In_178,In_1619);
or U1903 (N_1903,In_913,In_1596);
nor U1904 (N_1904,In_196,In_91);
or U1905 (N_1905,In_1746,In_801);
and U1906 (N_1906,In_297,In_1867);
nor U1907 (N_1907,In_1405,In_550);
and U1908 (N_1908,In_1936,In_116);
nor U1909 (N_1909,In_1846,In_197);
nand U1910 (N_1910,In_1924,In_1650);
or U1911 (N_1911,In_118,In_1504);
nor U1912 (N_1912,In_619,In_594);
or U1913 (N_1913,In_1317,In_439);
nor U1914 (N_1914,In_653,In_794);
nand U1915 (N_1915,In_500,In_401);
nand U1916 (N_1916,In_795,In_1750);
nand U1917 (N_1917,In_913,In_43);
nand U1918 (N_1918,In_1291,In_1156);
nor U1919 (N_1919,In_55,In_561);
nand U1920 (N_1920,In_1536,In_368);
or U1921 (N_1921,In_1110,In_722);
nor U1922 (N_1922,In_109,In_778);
nand U1923 (N_1923,In_1640,In_1532);
xnor U1924 (N_1924,In_738,In_1289);
nor U1925 (N_1925,In_1001,In_75);
nand U1926 (N_1926,In_566,In_467);
nor U1927 (N_1927,In_61,In_6);
or U1928 (N_1928,In_1867,In_385);
xor U1929 (N_1929,In_1698,In_601);
nand U1930 (N_1930,In_1929,In_1133);
and U1931 (N_1931,In_1541,In_795);
nor U1932 (N_1932,In_1087,In_532);
or U1933 (N_1933,In_518,In_1209);
and U1934 (N_1934,In_321,In_978);
nor U1935 (N_1935,In_1770,In_721);
or U1936 (N_1936,In_1358,In_1068);
or U1937 (N_1937,In_1421,In_1994);
nor U1938 (N_1938,In_475,In_1461);
nand U1939 (N_1939,In_575,In_287);
and U1940 (N_1940,In_513,In_1708);
nand U1941 (N_1941,In_1331,In_491);
and U1942 (N_1942,In_338,In_297);
nand U1943 (N_1943,In_713,In_1202);
or U1944 (N_1944,In_234,In_1959);
or U1945 (N_1945,In_1529,In_1804);
and U1946 (N_1946,In_1090,In_1819);
or U1947 (N_1947,In_512,In_969);
and U1948 (N_1948,In_1407,In_1919);
or U1949 (N_1949,In_935,In_200);
and U1950 (N_1950,In_292,In_1352);
and U1951 (N_1951,In_64,In_1898);
or U1952 (N_1952,In_1907,In_991);
xnor U1953 (N_1953,In_469,In_302);
nand U1954 (N_1954,In_1954,In_1138);
nand U1955 (N_1955,In_387,In_528);
nor U1956 (N_1956,In_229,In_1010);
and U1957 (N_1957,In_1951,In_1938);
nor U1958 (N_1958,In_1341,In_1417);
nand U1959 (N_1959,In_1157,In_1821);
nand U1960 (N_1960,In_1820,In_522);
nand U1961 (N_1961,In_225,In_1343);
nand U1962 (N_1962,In_426,In_1578);
nor U1963 (N_1963,In_633,In_1519);
xnor U1964 (N_1964,In_1682,In_1462);
or U1965 (N_1965,In_134,In_1483);
or U1966 (N_1966,In_925,In_1348);
xnor U1967 (N_1967,In_472,In_722);
and U1968 (N_1968,In_1251,In_50);
and U1969 (N_1969,In_1183,In_1531);
or U1970 (N_1970,In_148,In_443);
nor U1971 (N_1971,In_1007,In_972);
nand U1972 (N_1972,In_966,In_317);
xnor U1973 (N_1973,In_1520,In_1742);
or U1974 (N_1974,In_1301,In_410);
xor U1975 (N_1975,In_1822,In_349);
and U1976 (N_1976,In_1493,In_826);
nand U1977 (N_1977,In_1429,In_481);
xor U1978 (N_1978,In_552,In_1504);
or U1979 (N_1979,In_402,In_1211);
or U1980 (N_1980,In_1562,In_1878);
or U1981 (N_1981,In_1105,In_1723);
and U1982 (N_1982,In_375,In_1949);
nor U1983 (N_1983,In_1156,In_1453);
or U1984 (N_1984,In_1974,In_479);
or U1985 (N_1985,In_1958,In_1210);
nor U1986 (N_1986,In_677,In_1095);
and U1987 (N_1987,In_186,In_81);
and U1988 (N_1988,In_1697,In_1574);
nand U1989 (N_1989,In_637,In_160);
and U1990 (N_1990,In_867,In_652);
nor U1991 (N_1991,In_1718,In_513);
or U1992 (N_1992,In_1720,In_1013);
and U1993 (N_1993,In_585,In_1227);
nand U1994 (N_1994,In_1997,In_268);
nand U1995 (N_1995,In_1146,In_1094);
nor U1996 (N_1996,In_925,In_1806);
or U1997 (N_1997,In_1491,In_1729);
nor U1998 (N_1998,In_1318,In_269);
nand U1999 (N_1999,In_1594,In_1147);
or U2000 (N_2000,N_862,N_426);
nor U2001 (N_2001,N_1783,N_94);
nand U2002 (N_2002,N_1807,N_617);
and U2003 (N_2003,N_638,N_7);
nor U2004 (N_2004,N_353,N_759);
nor U2005 (N_2005,N_1305,N_92);
nand U2006 (N_2006,N_471,N_871);
nand U2007 (N_2007,N_1086,N_229);
or U2008 (N_2008,N_937,N_1659);
nor U2009 (N_2009,N_1918,N_232);
and U2010 (N_2010,N_905,N_888);
nor U2011 (N_2011,N_309,N_974);
or U2012 (N_2012,N_1015,N_1324);
and U2013 (N_2013,N_554,N_855);
nor U2014 (N_2014,N_1106,N_58);
nand U2015 (N_2015,N_1625,N_843);
xnor U2016 (N_2016,N_169,N_1507);
and U2017 (N_2017,N_1632,N_957);
and U2018 (N_2018,N_1233,N_668);
nand U2019 (N_2019,N_1368,N_161);
nor U2020 (N_2020,N_1350,N_1841);
xnor U2021 (N_2021,N_462,N_603);
nand U2022 (N_2022,N_972,N_838);
nand U2023 (N_2023,N_40,N_1478);
or U2024 (N_2024,N_343,N_1953);
xor U2025 (N_2025,N_481,N_1873);
xnor U2026 (N_2026,N_1171,N_380);
and U2027 (N_2027,N_158,N_1662);
nor U2028 (N_2028,N_1422,N_126);
nor U2029 (N_2029,N_1517,N_1696);
nand U2030 (N_2030,N_1413,N_66);
xor U2031 (N_2031,N_990,N_1263);
and U2032 (N_2032,N_872,N_1765);
and U2033 (N_2033,N_1854,N_1874);
or U2034 (N_2034,N_1195,N_934);
and U2035 (N_2035,N_362,N_679);
nand U2036 (N_2036,N_1661,N_36);
or U2037 (N_2037,N_1099,N_732);
nor U2038 (N_2038,N_1815,N_541);
nor U2039 (N_2039,N_195,N_1675);
nand U2040 (N_2040,N_1347,N_1101);
nor U2041 (N_2041,N_1083,N_1361);
xor U2042 (N_2042,N_1363,N_1870);
nor U2043 (N_2043,N_1446,N_363);
nor U2044 (N_2044,N_1141,N_1743);
and U2045 (N_2045,N_1029,N_516);
or U2046 (N_2046,N_1964,N_42);
nand U2047 (N_2047,N_1572,N_1767);
nor U2048 (N_2048,N_1828,N_544);
xor U2049 (N_2049,N_144,N_1489);
nor U2050 (N_2050,N_1822,N_1608);
or U2051 (N_2051,N_631,N_1339);
and U2052 (N_2052,N_228,N_1555);
and U2053 (N_2053,N_1417,N_249);
and U2054 (N_2054,N_491,N_289);
or U2055 (N_2055,N_1510,N_1485);
nand U2056 (N_2056,N_523,N_904);
and U2057 (N_2057,N_1343,N_63);
nand U2058 (N_2058,N_739,N_649);
or U2059 (N_2059,N_468,N_1120);
nor U2060 (N_2060,N_373,N_1913);
and U2061 (N_2061,N_355,N_1096);
or U2062 (N_2062,N_203,N_884);
nor U2063 (N_2063,N_1118,N_671);
nand U2064 (N_2064,N_1938,N_1455);
xnor U2065 (N_2065,N_883,N_1809);
and U2066 (N_2066,N_548,N_1470);
or U2067 (N_2067,N_1338,N_552);
nor U2068 (N_2068,N_1234,N_1158);
and U2069 (N_2069,N_1944,N_712);
or U2070 (N_2070,N_1900,N_1628);
and U2071 (N_2071,N_3,N_160);
nand U2072 (N_2072,N_1191,N_263);
or U2073 (N_2073,N_931,N_1871);
or U2074 (N_2074,N_1087,N_607);
nand U2075 (N_2075,N_51,N_1502);
or U2076 (N_2076,N_291,N_1883);
and U2077 (N_2077,N_1432,N_1845);
or U2078 (N_2078,N_135,N_261);
and U2079 (N_2079,N_1812,N_1801);
and U2080 (N_2080,N_1619,N_857);
and U2081 (N_2081,N_1356,N_1786);
nand U2082 (N_2082,N_181,N_207);
nand U2083 (N_2083,N_1253,N_245);
nor U2084 (N_2084,N_1258,N_948);
nor U2085 (N_2085,N_1906,N_1513);
nand U2086 (N_2086,N_1853,N_1535);
xnor U2087 (N_2087,N_547,N_1551);
or U2088 (N_2088,N_1341,N_1890);
and U2089 (N_2089,N_1344,N_1462);
and U2090 (N_2090,N_1621,N_1303);
or U2091 (N_2091,N_1333,N_1986);
nand U2092 (N_2092,N_1125,N_6);
nand U2093 (N_2093,N_204,N_1686);
nor U2094 (N_2094,N_1114,N_1017);
nand U2095 (N_2095,N_1075,N_216);
nor U2096 (N_2096,N_728,N_856);
nand U2097 (N_2097,N_236,N_1553);
nor U2098 (N_2098,N_432,N_15);
xor U2099 (N_2099,N_1394,N_164);
nor U2100 (N_2100,N_74,N_535);
nand U2101 (N_2101,N_1868,N_1227);
or U2102 (N_2102,N_9,N_1746);
and U2103 (N_2103,N_1062,N_286);
or U2104 (N_2104,N_533,N_773);
and U2105 (N_2105,N_955,N_1730);
or U2106 (N_2106,N_750,N_325);
and U2107 (N_2107,N_1219,N_848);
or U2108 (N_2108,N_434,N_1840);
and U2109 (N_2109,N_796,N_1838);
or U2110 (N_2110,N_1349,N_519);
and U2111 (N_2111,N_1724,N_1928);
nand U2112 (N_2112,N_1032,N_1025);
xor U2113 (N_2113,N_29,N_1579);
xor U2114 (N_2114,N_1805,N_882);
nand U2115 (N_2115,N_558,N_1117);
nand U2116 (N_2116,N_1629,N_1051);
and U2117 (N_2117,N_635,N_449);
nor U2118 (N_2118,N_267,N_1179);
and U2119 (N_2119,N_460,N_394);
nand U2120 (N_2120,N_107,N_425);
nand U2121 (N_2121,N_1833,N_944);
nor U2122 (N_2122,N_738,N_1583);
nor U2123 (N_2123,N_1149,N_310);
and U2124 (N_2124,N_1708,N_718);
nor U2125 (N_2125,N_482,N_526);
nand U2126 (N_2126,N_69,N_317);
nand U2127 (N_2127,N_1399,N_1990);
or U2128 (N_2128,N_876,N_1323);
xor U2129 (N_2129,N_304,N_803);
nand U2130 (N_2130,N_445,N_1565);
or U2131 (N_2131,N_1274,N_1915);
or U2132 (N_2132,N_1818,N_1395);
or U2133 (N_2133,N_1346,N_487);
xnor U2134 (N_2134,N_1795,N_1894);
nand U2135 (N_2135,N_663,N_1917);
or U2136 (N_2136,N_290,N_1558);
or U2137 (N_2137,N_1302,N_32);
or U2138 (N_2138,N_1111,N_1855);
xor U2139 (N_2139,N_262,N_298);
or U2140 (N_2140,N_1452,N_702);
and U2141 (N_2141,N_441,N_1459);
nor U2142 (N_2142,N_1524,N_350);
and U2143 (N_2143,N_1610,N_1451);
or U2144 (N_2144,N_1332,N_420);
nand U2145 (N_2145,N_1094,N_1095);
and U2146 (N_2146,N_1788,N_14);
and U2147 (N_2147,N_1359,N_1653);
xnor U2148 (N_2148,N_1823,N_597);
and U2149 (N_2149,N_1292,N_1007);
or U2150 (N_2150,N_1284,N_25);
nand U2151 (N_2151,N_1705,N_1951);
nand U2152 (N_2152,N_969,N_1634);
or U2153 (N_2153,N_191,N_1576);
nand U2154 (N_2154,N_1693,N_706);
or U2155 (N_2155,N_522,N_1445);
or U2156 (N_2156,N_637,N_1942);
nand U2157 (N_2157,N_1711,N_11);
nor U2158 (N_2158,N_1568,N_1666);
or U2159 (N_2159,N_19,N_247);
or U2160 (N_2160,N_602,N_1476);
nand U2161 (N_2161,N_949,N_1642);
and U2162 (N_2162,N_1378,N_143);
nand U2163 (N_2163,N_1116,N_314);
nor U2164 (N_2164,N_1646,N_1071);
nor U2165 (N_2165,N_1027,N_1479);
nor U2166 (N_2166,N_1793,N_1406);
nand U2167 (N_2167,N_1415,N_1469);
nand U2168 (N_2168,N_810,N_469);
nand U2169 (N_2169,N_1612,N_1720);
and U2170 (N_2170,N_456,N_1772);
nand U2171 (N_2171,N_1384,N_584);
and U2172 (N_2172,N_1506,N_703);
nor U2173 (N_2173,N_225,N_214);
nor U2174 (N_2174,N_556,N_1971);
xor U2175 (N_2175,N_696,N_1442);
nand U2176 (N_2176,N_772,N_1790);
nand U2177 (N_2177,N_1600,N_1174);
nand U2178 (N_2178,N_1526,N_1992);
nand U2179 (N_2179,N_1620,N_1758);
nor U2180 (N_2180,N_954,N_1367);
and U2181 (N_2181,N_758,N_172);
or U2182 (N_2182,N_1474,N_623);
and U2183 (N_2183,N_134,N_1220);
or U2184 (N_2184,N_1533,N_559);
nor U2185 (N_2185,N_963,N_1963);
or U2186 (N_2186,N_643,N_681);
and U2187 (N_2187,N_430,N_754);
and U2188 (N_2188,N_1969,N_1611);
nor U2189 (N_2189,N_1391,N_1617);
or U2190 (N_2190,N_374,N_335);
nand U2191 (N_2191,N_1026,N_1799);
nand U2192 (N_2192,N_964,N_958);
nand U2193 (N_2193,N_13,N_776);
nand U2194 (N_2194,N_813,N_1050);
or U2195 (N_2195,N_893,N_1092);
nand U2196 (N_2196,N_1176,N_114);
nor U2197 (N_2197,N_785,N_1755);
nand U2198 (N_2198,N_672,N_439);
xnor U2199 (N_2199,N_266,N_486);
nand U2200 (N_2200,N_1736,N_1960);
or U2201 (N_2201,N_1945,N_1335);
and U2202 (N_2202,N_1864,N_945);
nor U2203 (N_2203,N_338,N_1392);
nor U2204 (N_2204,N_724,N_765);
nor U2205 (N_2205,N_1570,N_527);
nand U2206 (N_2206,N_709,N_716);
and U2207 (N_2207,N_61,N_270);
nor U2208 (N_2208,N_1259,N_1269);
or U2209 (N_2209,N_532,N_1345);
nor U2210 (N_2210,N_847,N_720);
nand U2211 (N_2211,N_766,N_1172);
and U2212 (N_2212,N_1924,N_1678);
xor U2213 (N_2213,N_762,N_1537);
or U2214 (N_2214,N_780,N_1859);
nand U2215 (N_2215,N_1782,N_1364);
nand U2216 (N_2216,N_682,N_248);
or U2217 (N_2217,N_1658,N_1567);
nand U2218 (N_2218,N_666,N_387);
nor U2219 (N_2219,N_825,N_288);
nand U2220 (N_2220,N_722,N_665);
nand U2221 (N_2221,N_585,N_524);
and U2222 (N_2222,N_1067,N_379);
nand U2223 (N_2223,N_1377,N_1268);
and U2224 (N_2224,N_253,N_727);
nor U2225 (N_2225,N_879,N_1714);
xor U2226 (N_2226,N_1140,N_339);
or U2227 (N_2227,N_1456,N_81);
and U2228 (N_2228,N_113,N_795);
and U2229 (N_2229,N_1858,N_485);
nand U2230 (N_2230,N_1307,N_1491);
nor U2231 (N_2231,N_1273,N_564);
or U2232 (N_2232,N_1203,N_992);
and U2233 (N_2233,N_1310,N_612);
nor U2234 (N_2234,N_145,N_837);
xnor U2235 (N_2235,N_1909,N_0);
nand U2236 (N_2236,N_1631,N_833);
and U2237 (N_2237,N_1719,N_269);
nor U2238 (N_2238,N_112,N_165);
xnor U2239 (N_2239,N_587,N_802);
nor U2240 (N_2240,N_102,N_1301);
nor U2241 (N_2241,N_595,N_1309);
xor U2242 (N_2242,N_755,N_293);
and U2243 (N_2243,N_659,N_977);
and U2244 (N_2244,N_278,N_390);
and U2245 (N_2245,N_133,N_1433);
or U2246 (N_2246,N_1242,N_793);
nand U2247 (N_2247,N_4,N_1523);
or U2248 (N_2248,N_1463,N_226);
or U2249 (N_2249,N_705,N_1319);
and U2250 (N_2250,N_389,N_534);
nor U2251 (N_2251,N_1006,N_1069);
or U2252 (N_2252,N_407,N_1129);
and U2253 (N_2253,N_1369,N_1519);
nor U2254 (N_2254,N_1295,N_1293);
nand U2255 (N_2255,N_1768,N_1283);
nor U2256 (N_2256,N_279,N_1213);
nor U2257 (N_2257,N_892,N_208);
and U2258 (N_2258,N_1712,N_1595);
or U2259 (N_2259,N_422,N_323);
nand U2260 (N_2260,N_930,N_1903);
nand U2261 (N_2261,N_503,N_952);
nand U2262 (N_2262,N_334,N_345);
xor U2263 (N_2263,N_369,N_1824);
nor U2264 (N_2264,N_1396,N_1122);
or U2265 (N_2265,N_1898,N_546);
xnor U2266 (N_2266,N_178,N_606);
nor U2267 (N_2267,N_1144,N_543);
and U2268 (N_2268,N_27,N_790);
and U2269 (N_2269,N_517,N_1441);
or U2270 (N_2270,N_187,N_302);
nand U2271 (N_2271,N_72,N_109);
or U2272 (N_2272,N_84,N_988);
xnor U2273 (N_2273,N_1892,N_213);
and U2274 (N_2274,N_1905,N_1460);
nor U2275 (N_2275,N_1707,N_1152);
or U2276 (N_2276,N_1573,N_1146);
or U2277 (N_2277,N_1166,N_128);
nand U2278 (N_2278,N_1254,N_1353);
xor U2279 (N_2279,N_563,N_271);
and U2280 (N_2280,N_139,N_1260);
nor U2281 (N_2281,N_987,N_798);
xor U2282 (N_2282,N_922,N_80);
or U2283 (N_2283,N_1819,N_1252);
nor U2284 (N_2284,N_1958,N_1054);
or U2285 (N_2285,N_717,N_925);
or U2286 (N_2286,N_1225,N_382);
and U2287 (N_2287,N_807,N_1649);
nor U2288 (N_2288,N_1635,N_736);
nor U2289 (N_2289,N_472,N_1287);
nand U2290 (N_2290,N_1516,N_52);
nand U2291 (N_2291,N_1919,N_1729);
nor U2292 (N_2292,N_497,N_1577);
nand U2293 (N_2293,N_1676,N_513);
or U2294 (N_2294,N_695,N_1170);
and U2295 (N_2295,N_936,N_56);
or U2296 (N_2296,N_1546,N_1820);
nor U2297 (N_2297,N_1499,N_1785);
or U2298 (N_2298,N_572,N_1668);
or U2299 (N_2299,N_31,N_348);
and U2300 (N_2300,N_316,N_147);
nor U2301 (N_2301,N_1531,N_1251);
nand U2302 (N_2302,N_1817,N_1030);
or U2303 (N_2303,N_1811,N_1186);
nand U2304 (N_2304,N_62,N_836);
nand U2305 (N_2305,N_1457,N_1185);
nor U2306 (N_2306,N_1246,N_1052);
or U2307 (N_2307,N_48,N_1340);
and U2308 (N_2308,N_393,N_633);
nand U2309 (N_2309,N_285,N_1754);
xnor U2310 (N_2310,N_189,N_182);
nor U2311 (N_2311,N_902,N_520);
nand U2312 (N_2312,N_1154,N_1464);
nand U2313 (N_2313,N_116,N_1737);
and U2314 (N_2314,N_1382,N_1580);
nor U2315 (N_2315,N_846,N_1749);
nor U2316 (N_2316,N_723,N_971);
nand U2317 (N_2317,N_530,N_866);
nand U2318 (N_2318,N_1379,N_1650);
and U2319 (N_2319,N_8,N_1780);
or U2320 (N_2320,N_235,N_742);
nor U2321 (N_2321,N_447,N_18);
nor U2322 (N_2322,N_1001,N_488);
and U2323 (N_2323,N_540,N_1312);
and U2324 (N_2324,N_894,N_1436);
or U2325 (N_2325,N_734,N_1270);
or U2326 (N_2326,N_1437,N_1016);
nor U2327 (N_2327,N_700,N_142);
and U2328 (N_2328,N_1839,N_1372);
nor U2329 (N_2329,N_1426,N_1849);
nand U2330 (N_2330,N_419,N_1726);
nor U2331 (N_2331,N_1881,N_1060);
nand U2332 (N_2332,N_1723,N_489);
nor U2333 (N_2333,N_315,N_1012);
nor U2334 (N_2334,N_746,N_1561);
nor U2335 (N_2335,N_805,N_454);
nor U2336 (N_2336,N_1728,N_1362);
nor U2337 (N_2337,N_1398,N_664);
xor U2338 (N_2338,N_1511,N_392);
and U2339 (N_2339,N_781,N_1420);
or U2340 (N_2340,N_1068,N_1753);
nand U2341 (N_2341,N_1689,N_1641);
nand U2342 (N_2342,N_886,N_771);
and U2343 (N_2343,N_1500,N_1503);
nor U2344 (N_2344,N_1132,N_436);
and U2345 (N_2345,N_1107,N_1961);
nor U2346 (N_2346,N_573,N_1177);
nand U2347 (N_2347,N_965,N_512);
nor U2348 (N_2348,N_1827,N_763);
nor U2349 (N_2349,N_550,N_1688);
and U2350 (N_2350,N_277,N_313);
nand U2351 (N_2351,N_1893,N_1342);
nor U2352 (N_2352,N_1355,N_791);
xor U2353 (N_2353,N_737,N_93);
xnor U2354 (N_2354,N_411,N_50);
nor U2355 (N_2355,N_1334,N_769);
nor U2356 (N_2356,N_811,N_673);
and U2357 (N_2357,N_1532,N_1745);
or U2358 (N_2358,N_1552,N_683);
nor U2359 (N_2359,N_16,N_1256);
nor U2360 (N_2360,N_364,N_1695);
or U2361 (N_2361,N_779,N_667);
and U2362 (N_2362,N_1080,N_1127);
or U2363 (N_2363,N_1846,N_721);
or U2364 (N_2364,N_1314,N_1280);
or U2365 (N_2365,N_1447,N_613);
nand U2366 (N_2366,N_870,N_1907);
and U2367 (N_2367,N_175,N_1444);
or U2368 (N_2368,N_1867,N_1761);
nor U2369 (N_2369,N_311,N_525);
xnor U2370 (N_2370,N_414,N_1575);
and U2371 (N_2371,N_1212,N_320);
xnor U2372 (N_2372,N_443,N_1237);
and U2373 (N_2373,N_1727,N_1589);
and U2374 (N_2374,N_1574,N_138);
and U2375 (N_2375,N_1188,N_661);
or U2376 (N_2376,N_1286,N_829);
nor U2377 (N_2377,N_828,N_1710);
or U2378 (N_2378,N_1781,N_1181);
or U2379 (N_2379,N_1687,N_90);
or U2380 (N_2380,N_1241,N_598);
nor U2381 (N_2381,N_73,N_1070);
and U2382 (N_2382,N_1607,N_1716);
nor U2383 (N_2383,N_1104,N_376);
or U2384 (N_2384,N_37,N_747);
or U2385 (N_2385,N_1036,N_1003);
nand U2386 (N_2386,N_1412,N_704);
nor U2387 (N_2387,N_1606,N_939);
nor U2388 (N_2388,N_1315,N_1147);
nand U2389 (N_2389,N_1074,N_1091);
xnor U2390 (N_2390,N_366,N_1979);
nand U2391 (N_2391,N_1105,N_538);
and U2392 (N_2392,N_1515,N_507);
xor U2393 (N_2393,N_151,N_475);
or U2394 (N_2394,N_1311,N_280);
and U2395 (N_2395,N_642,N_1908);
and U2396 (N_2396,N_670,N_1317);
nor U2397 (N_2397,N_1848,N_1798);
nor U2398 (N_2398,N_1124,N_636);
nor U2399 (N_2399,N_242,N_692);
or U2400 (N_2400,N_730,N_574);
or U2401 (N_2401,N_615,N_179);
nor U2402 (N_2402,N_79,N_596);
or U2403 (N_2403,N_577,N_921);
nand U2404 (N_2404,N_17,N_45);
or U2405 (N_2405,N_627,N_675);
nor U2406 (N_2406,N_130,N_197);
nor U2407 (N_2407,N_1747,N_609);
and U2408 (N_2408,N_1508,N_864);
nand U2409 (N_2409,N_252,N_405);
nand U2410 (N_2410,N_1983,N_167);
or U2411 (N_2411,N_1085,N_254);
nor U2412 (N_2412,N_1701,N_1081);
and U2413 (N_2413,N_1151,N_186);
or U2414 (N_2414,N_1352,N_1477);
and U2415 (N_2415,N_129,N_1571);
nand U2416 (N_2416,N_435,N_1159);
xor U2417 (N_2417,N_1955,N_312);
nand U2418 (N_2418,N_131,N_624);
xnor U2419 (N_2419,N_1680,N_647);
nor U2420 (N_2420,N_86,N_352);
nand U2421 (N_2421,N_1133,N_132);
and U2422 (N_2422,N_192,N_853);
nand U2423 (N_2423,N_782,N_1775);
nor U2424 (N_2424,N_1198,N_1157);
nor U2425 (N_2425,N_1999,N_174);
or U2426 (N_2426,N_457,N_804);
nor U2427 (N_2427,N_555,N_938);
or U2428 (N_2428,N_1637,N_222);
and U2429 (N_2429,N_841,N_1648);
nand U2430 (N_2430,N_1058,N_1238);
and U2431 (N_2431,N_827,N_137);
and U2432 (N_2432,N_1763,N_1214);
nand U2433 (N_2433,N_1078,N_1542);
and U2434 (N_2434,N_1590,N_1393);
xor U2435 (N_2435,N_1977,N_1375);
or U2436 (N_2436,N_1946,N_1496);
nand U2437 (N_2437,N_1088,N_993);
or U2438 (N_2438,N_234,N_1313);
nor U2439 (N_2439,N_108,N_1173);
nand U2440 (N_2440,N_588,N_404);
or U2441 (N_2441,N_1897,N_1414);
or U2442 (N_2442,N_375,N_241);
nor U2443 (N_2443,N_1483,N_684);
nor U2444 (N_2444,N_1102,N_1509);
nor U2445 (N_2445,N_823,N_1562);
nor U2446 (N_2446,N_1126,N_946);
or U2447 (N_2447,N_982,N_1825);
nor U2448 (N_2448,N_561,N_177);
nand U2449 (N_2449,N_1019,N_428);
and U2450 (N_2450,N_714,N_321);
nor U2451 (N_2451,N_579,N_85);
nand U2452 (N_2452,N_1539,N_1584);
and U2453 (N_2453,N_940,N_402);
xnor U2454 (N_2454,N_97,N_551);
or U2455 (N_2455,N_1331,N_1501);
xnor U2456 (N_2456,N_1427,N_1388);
and U2457 (N_2457,N_578,N_1262);
nor U2458 (N_2458,N_1813,N_357);
xnor U2459 (N_2459,N_1547,N_1722);
and U2460 (N_2460,N_386,N_421);
nor U2461 (N_2461,N_1912,N_975);
nand U2462 (N_2462,N_240,N_725);
nor U2463 (N_2463,N_506,N_715);
nor U2464 (N_2464,N_1266,N_1581);
or U2465 (N_2465,N_162,N_1700);
nand U2466 (N_2466,N_246,N_1592);
or U2467 (N_2467,N_877,N_652);
nor U2468 (N_2468,N_110,N_125);
nand U2469 (N_2469,N_1880,N_365);
nand U2470 (N_2470,N_1821,N_580);
nor U2471 (N_2471,N_1564,N_1156);
or U2472 (N_2472,N_1850,N_184);
nand U2473 (N_2473,N_986,N_528);
nand U2474 (N_2474,N_869,N_1076);
nand U2475 (N_2475,N_1370,N_1598);
and U2476 (N_2476,N_619,N_1603);
and U2477 (N_2477,N_1288,N_38);
xor U2478 (N_2478,N_1504,N_660);
and U2479 (N_2479,N_1633,N_1425);
or U2480 (N_2480,N_205,N_1486);
or U2481 (N_2481,N_983,N_361);
and U2482 (N_2482,N_1837,N_1599);
xnor U2483 (N_2483,N_576,N_53);
nor U2484 (N_2484,N_171,N_1285);
xnor U2485 (N_2485,N_1109,N_383);
and U2486 (N_2486,N_654,N_1713);
nor U2487 (N_2487,N_494,N_748);
or U2488 (N_2488,N_1236,N_1520);
or U2489 (N_2489,N_1950,N_1299);
and U2490 (N_2490,N_1694,N_1040);
and U2491 (N_2491,N_634,N_1984);
and U2492 (N_2492,N_1965,N_450);
or U2493 (N_2493,N_1941,N_970);
or U2494 (N_2494,N_1932,N_1929);
nand U2495 (N_2495,N_1647,N_1901);
or U2496 (N_2496,N_1430,N_1360);
nor U2497 (N_2497,N_1265,N_622);
nor U2498 (N_2498,N_816,N_1998);
nand U2499 (N_2499,N_985,N_1328);
nor U2500 (N_2500,N_764,N_1702);
or U2501 (N_2501,N_1865,N_644);
nand U2502 (N_2502,N_1401,N_1381);
nor U2503 (N_2503,N_1139,N_508);
nor U2504 (N_2504,N_1993,N_981);
nor U2505 (N_2505,N_1204,N_223);
nand U2506 (N_2506,N_371,N_1803);
nand U2507 (N_2507,N_283,N_1431);
xnor U2508 (N_2508,N_844,N_1578);
nand U2509 (N_2509,N_356,N_1232);
and U2510 (N_2510,N_935,N_1059);
nor U2511 (N_2511,N_1044,N_1624);
or U2512 (N_2512,N_401,N_865);
and U2513 (N_2513,N_1229,N_687);
nand U2514 (N_2514,N_768,N_1327);
xor U2515 (N_2515,N_1856,N_1777);
nor U2516 (N_2516,N_1836,N_370);
nand U2517 (N_2517,N_1056,N_95);
xnor U2518 (N_2518,N_1512,N_1654);
and U2519 (N_2519,N_947,N_1153);
nor U2520 (N_2520,N_306,N_347);
nand U2521 (N_2521,N_1863,N_185);
nor U2522 (N_2522,N_1216,N_1494);
xor U2523 (N_2523,N_111,N_307);
nand U2524 (N_2524,N_1326,N_1100);
xor U2525 (N_2525,N_997,N_1636);
nand U2526 (N_2526,N_333,N_54);
and U2527 (N_2527,N_1771,N_1530);
or U2528 (N_2528,N_1609,N_331);
xnor U2529 (N_2529,N_873,N_65);
and U2530 (N_2530,N_1454,N_710);
nor U2531 (N_2531,N_1759,N_1691);
xnor U2532 (N_2532,N_1748,N_156);
and U2533 (N_2533,N_1742,N_1936);
nor U2534 (N_2534,N_1887,N_806);
or U2535 (N_2535,N_1740,N_1222);
and U2536 (N_2536,N_1980,N_359);
or U2537 (N_2537,N_1731,N_1554);
and U2538 (N_2538,N_1482,N_1134);
xor U2539 (N_2539,N_605,N_163);
nand U2540 (N_2540,N_655,N_224);
and U2541 (N_2541,N_238,N_1484);
nand U2542 (N_2542,N_1769,N_817);
and U2543 (N_2543,N_809,N_994);
nor U2544 (N_2544,N_368,N_438);
and U2545 (N_2545,N_509,N_914);
xnor U2546 (N_2546,N_403,N_1738);
and U2547 (N_2547,N_850,N_1308);
nor U2548 (N_2548,N_1304,N_1434);
or U2549 (N_2549,N_698,N_593);
nand U2550 (N_2550,N_951,N_927);
nand U2551 (N_2551,N_1291,N_1792);
or U2552 (N_2552,N_1065,N_35);
or U2553 (N_2553,N_1429,N_341);
or U2554 (N_2554,N_96,N_452);
or U2555 (N_2555,N_1910,N_1271);
nor U2556 (N_2556,N_217,N_821);
nand U2557 (N_2557,N_568,N_1536);
xnor U2558 (N_2558,N_1498,N_300);
or U2559 (N_2559,N_1832,N_1587);
nor U2560 (N_2560,N_91,N_1113);
and U2561 (N_2561,N_1760,N_943);
nand U2562 (N_2562,N_451,N_41);
and U2563 (N_2563,N_1490,N_1468);
nand U2564 (N_2564,N_1289,N_1390);
and U2565 (N_2565,N_244,N_693);
nand U2566 (N_2566,N_1373,N_1014);
xnor U2567 (N_2567,N_1387,N_950);
and U2568 (N_2568,N_1593,N_1073);
and U2569 (N_2569,N_1325,N_1002);
nand U2570 (N_2570,N_777,N_1704);
nand U2571 (N_2571,N_1320,N_453);
nand U2572 (N_2572,N_1208,N_694);
or U2573 (N_2573,N_395,N_1756);
and U2574 (N_2574,N_1168,N_1869);
and U2575 (N_2575,N_1739,N_1994);
and U2576 (N_2576,N_657,N_1779);
nor U2577 (N_2577,N_1911,N_1187);
or U2578 (N_2578,N_196,N_1940);
and U2579 (N_2579,N_416,N_1752);
nor U2580 (N_2580,N_1055,N_188);
and U2581 (N_2581,N_1959,N_1541);
nand U2582 (N_2582,N_1321,N_868);
nor U2583 (N_2583,N_575,N_961);
nor U2584 (N_2584,N_230,N_466);
or U2585 (N_2585,N_1221,N_20);
and U2586 (N_2586,N_43,N_1904);
nand U2587 (N_2587,N_1358,N_1560);
and U2588 (N_2588,N_923,N_1136);
nor U2589 (N_2589,N_1569,N_1119);
nand U2590 (N_2590,N_1732,N_1879);
or U2591 (N_2591,N_431,N_388);
and U2592 (N_2592,N_1656,N_1559);
or U2593 (N_2593,N_1215,N_1810);
nand U2594 (N_2594,N_148,N_1639);
nor U2595 (N_2595,N_1644,N_168);
nand U2596 (N_2596,N_1645,N_1896);
xor U2597 (N_2597,N_1538,N_326);
nand U2598 (N_2598,N_1371,N_676);
or U2599 (N_2599,N_909,N_1178);
or U2600 (N_2600,N_998,N_822);
nor U2601 (N_2601,N_913,N_688);
or U2602 (N_2602,N_1926,N_470);
or U2603 (N_2603,N_294,N_743);
or U2604 (N_2604,N_860,N_529);
or U2605 (N_2605,N_1115,N_980);
nor U2606 (N_2606,N_645,N_1857);
xnor U2607 (N_2607,N_1690,N_1090);
or U2608 (N_2608,N_1834,N_212);
nand U2609 (N_2609,N_272,N_840);
or U2610 (N_2610,N_149,N_1605);
nand U2611 (N_2611,N_1615,N_358);
and U2612 (N_2612,N_59,N_1318);
nor U2613 (N_2613,N_1962,N_372);
or U2614 (N_2614,N_23,N_1439);
and U2615 (N_2615,N_1218,N_1021);
and U2616 (N_2616,N_719,N_1038);
nand U2617 (N_2617,N_221,N_788);
or U2618 (N_2618,N_851,N_1013);
nor U2619 (N_2619,N_1135,N_378);
xor U2620 (N_2620,N_1063,N_1243);
nor U2621 (N_2621,N_1161,N_1630);
nor U2622 (N_2622,N_708,N_1316);
and U2623 (N_2623,N_33,N_1480);
nor U2624 (N_2624,N_408,N_942);
nand U2625 (N_2625,N_1843,N_87);
xnor U2626 (N_2626,N_194,N_303);
or U2627 (N_2627,N_908,N_1039);
xnor U2628 (N_2628,N_819,N_1791);
nor U2629 (N_2629,N_504,N_1250);
and U2630 (N_2630,N_1949,N_1473);
nor U2631 (N_2631,N_258,N_1891);
and U2632 (N_2632,N_502,N_193);
and U2633 (N_2633,N_808,N_960);
nor U2634 (N_2634,N_1000,N_1209);
nand U2635 (N_2635,N_117,N_180);
nor U2636 (N_2636,N_233,N_1112);
nand U2637 (N_2637,N_60,N_1438);
or U2638 (N_2638,N_1272,N_1297);
and U2639 (N_2639,N_424,N_480);
xor U2640 (N_2640,N_219,N_490);
nand U2641 (N_2641,N_1721,N_1996);
and U2642 (N_2642,N_745,N_1416);
nand U2643 (N_2643,N_75,N_691);
and U2644 (N_2644,N_1652,N_1145);
nand U2645 (N_2645,N_630,N_1466);
xnor U2646 (N_2646,N_199,N_381);
and U2647 (N_2647,N_1336,N_646);
and U2648 (N_2648,N_891,N_1981);
or U2649 (N_2649,N_1108,N_1471);
and U2650 (N_2650,N_1023,N_464);
and U2651 (N_2651,N_1860,N_966);
nand U2652 (N_2652,N_1084,N_920);
or U2653 (N_2653,N_295,N_28);
nand U2654 (N_2654,N_418,N_500);
nor U2655 (N_2655,N_478,N_582);
or U2656 (N_2656,N_880,N_55);
nand U2657 (N_2657,N_824,N_726);
and U2658 (N_2658,N_792,N_662);
and U2659 (N_2659,N_1397,N_775);
or U2660 (N_2660,N_653,N_1987);
xnor U2661 (N_2661,N_391,N_608);
nor U2662 (N_2662,N_354,N_299);
or U2663 (N_2663,N_1549,N_1276);
xnor U2664 (N_2664,N_268,N_427);
or U2665 (N_2665,N_1672,N_1180);
nand U2666 (N_2666,N_209,N_1638);
nor U2667 (N_2667,N_282,N_173);
xnor U2668 (N_2668,N_978,N_1762);
xnor U2669 (N_2669,N_99,N_1385);
and U2670 (N_2670,N_1525,N_1366);
xnor U2671 (N_2671,N_1235,N_996);
nor U2672 (N_2672,N_1231,N_1585);
and U2673 (N_2673,N_360,N_1923);
nand U2674 (N_2674,N_1402,N_1684);
xnor U2675 (N_2675,N_1475,N_783);
nand U2676 (N_2676,N_1957,N_458);
xnor U2677 (N_2677,N_999,N_677);
or U2678 (N_2678,N_628,N_1814);
nor U2679 (N_2679,N_1028,N_1935);
and U2680 (N_2680,N_397,N_484);
xor U2681 (N_2681,N_1202,N_104);
nand U2682 (N_2682,N_1718,N_1383);
nor U2683 (N_2683,N_284,N_874);
nor U2684 (N_2684,N_835,N_678);
nand U2685 (N_2685,N_1540,N_124);
and U2686 (N_2686,N_136,N_919);
xnor U2687 (N_2687,N_505,N_1764);
nor U2688 (N_2688,N_1279,N_1403);
and U2689 (N_2689,N_592,N_260);
nor U2690 (N_2690,N_928,N_281);
nand U2691 (N_2691,N_800,N_761);
and U2692 (N_2692,N_1757,N_859);
and U2693 (N_2693,N_1064,N_959);
and U2694 (N_2694,N_152,N_1275);
nand U2695 (N_2695,N_995,N_1844);
or U2696 (N_2696,N_256,N_176);
nor U2697 (N_2697,N_962,N_1223);
or U2698 (N_2698,N_308,N_1199);
nand U2699 (N_2699,N_483,N_926);
and U2700 (N_2700,N_398,N_1045);
nor U2701 (N_2701,N_1985,N_586);
nand U2702 (N_2702,N_1481,N_1183);
and U2703 (N_2703,N_967,N_814);
or U2704 (N_2704,N_1925,N_1528);
nand U2705 (N_2705,N_202,N_429);
and U2706 (N_2706,N_1920,N_616);
and U2707 (N_2707,N_1563,N_1037);
and U2708 (N_2708,N_1206,N_1626);
nor U2709 (N_2709,N_1797,N_685);
or U2710 (N_2710,N_1937,N_68);
xnor U2711 (N_2711,N_1947,N_477);
nand U2712 (N_2712,N_1493,N_157);
and U2713 (N_2713,N_887,N_1966);
and U2714 (N_2714,N_898,N_77);
nand U2715 (N_2715,N_1142,N_1751);
nand U2716 (N_2716,N_1008,N_47);
or U2717 (N_2717,N_1667,N_567);
and U2718 (N_2718,N_583,N_437);
xnor U2719 (N_2719,N_70,N_328);
or U2720 (N_2720,N_1205,N_44);
or U2721 (N_2721,N_337,N_377);
nand U2722 (N_2722,N_1692,N_501);
xor U2723 (N_2723,N_257,N_1882);
nand U2724 (N_2724,N_1098,N_863);
or U2725 (N_2725,N_498,N_118);
or U2726 (N_2726,N_1899,N_1294);
xor U2727 (N_2727,N_442,N_1952);
nand U2728 (N_2728,N_30,N_1123);
nand U2729 (N_2729,N_570,N_1072);
nor U2730 (N_2730,N_1972,N_911);
nor U2731 (N_2731,N_1669,N_701);
nor U2732 (N_2732,N_1357,N_467);
xnor U2733 (N_2733,N_1982,N_1024);
nand U2734 (N_2734,N_1582,N_697);
xor U2735 (N_2735,N_433,N_1956);
or U2736 (N_2736,N_1789,N_915);
and U2737 (N_2737,N_1365,N_198);
nor U2738 (N_2738,N_1192,N_1794);
nand U2739 (N_2739,N_1835,N_1703);
nor U2740 (N_2740,N_1277,N_1622);
xor U2741 (N_2741,N_818,N_273);
nor U2742 (N_2742,N_367,N_1773);
nand U2743 (N_2743,N_1,N_1495);
or U2744 (N_2744,N_330,N_329);
or U2745 (N_2745,N_49,N_1348);
nand U2746 (N_2746,N_1010,N_1831);
xor U2747 (N_2747,N_1043,N_1405);
or U2748 (N_2748,N_1804,N_1664);
nor U2749 (N_2749,N_1954,N_711);
nand U2750 (N_2750,N_1933,N_64);
nor U2751 (N_2751,N_1137,N_1009);
xor U2752 (N_2752,N_1706,N_1829);
or U2753 (N_2753,N_82,N_1774);
nor U2754 (N_2754,N_155,N_384);
or U2755 (N_2755,N_1047,N_1097);
and U2756 (N_2756,N_658,N_1715);
and U2757 (N_2757,N_140,N_318);
or U2758 (N_2758,N_342,N_889);
nand U2759 (N_2759,N_1110,N_542);
xnor U2760 (N_2760,N_744,N_1851);
or U2761 (N_2761,N_1766,N_1614);
xor U2762 (N_2762,N_21,N_1816);
nand U2763 (N_2763,N_5,N_201);
and U2764 (N_2764,N_1643,N_1698);
xnor U2765 (N_2765,N_417,N_515);
and U2766 (N_2766,N_680,N_590);
or U2767 (N_2767,N_1862,N_918);
and U2768 (N_2768,N_1679,N_621);
nand U2769 (N_2769,N_1921,N_292);
nand U2770 (N_2770,N_1613,N_444);
xor U2771 (N_2771,N_569,N_1974);
nand U2772 (N_2772,N_1386,N_220);
nor U2773 (N_2773,N_1601,N_1784);
and U2774 (N_2774,N_1261,N_115);
nand U2775 (N_2775,N_154,N_752);
nand U2776 (N_2776,N_1267,N_1847);
xor U2777 (N_2777,N_396,N_903);
or U2778 (N_2778,N_1443,N_1995);
and U2779 (N_2779,N_1699,N_346);
and U2780 (N_2780,N_473,N_1300);
xor U2781 (N_2781,N_1093,N_406);
or U2782 (N_2782,N_1458,N_581);
or U2783 (N_2783,N_103,N_1975);
and U2784 (N_2784,N_1492,N_531);
nand U2785 (N_2785,N_753,N_1872);
or U2786 (N_2786,N_976,N_1596);
or U2787 (N_2787,N_1042,N_1020);
nor U2788 (N_2788,N_1602,N_1389);
and U2789 (N_2789,N_912,N_324);
nor U2790 (N_2790,N_907,N_24);
or U2791 (N_2791,N_1226,N_1197);
or U2792 (N_2792,N_571,N_1591);
or U2793 (N_2793,N_1978,N_1683);
nand U2794 (N_2794,N_1281,N_106);
and U2795 (N_2795,N_1376,N_1770);
and U2796 (N_2796,N_231,N_618);
nor U2797 (N_2797,N_200,N_297);
nor U2798 (N_2798,N_275,N_1682);
nor U2799 (N_2799,N_1976,N_39);
and U2800 (N_2800,N_699,N_797);
xor U2801 (N_2801,N_1895,N_1296);
nand U2802 (N_2802,N_1733,N_1351);
and U2803 (N_2803,N_881,N_1717);
and U2804 (N_2804,N_924,N_1467);
nand U2805 (N_2805,N_190,N_1597);
nand U2806 (N_2806,N_239,N_22);
and U2807 (N_2807,N_1194,N_1306);
or U2808 (N_2808,N_1184,N_1130);
nor U2809 (N_2809,N_153,N_170);
and U2810 (N_2810,N_34,N_1927);
xor U2811 (N_2811,N_1527,N_1207);
or U2812 (N_2812,N_929,N_1550);
or U2813 (N_2813,N_896,N_159);
and U2814 (N_2814,N_499,N_991);
or U2815 (N_2815,N_932,N_956);
or U2816 (N_2816,N_474,N_1830);
nor U2817 (N_2817,N_562,N_1160);
and U2818 (N_2818,N_749,N_1245);
and U2819 (N_2819,N_119,N_1380);
nor U2820 (N_2820,N_1004,N_1247);
or U2821 (N_2821,N_251,N_1408);
nor U2822 (N_2822,N_514,N_674);
and U2823 (N_2823,N_1970,N_1228);
or U2824 (N_2824,N_1670,N_250);
or U2825 (N_2825,N_121,N_10);
nor U2826 (N_2826,N_789,N_614);
xnor U2827 (N_2827,N_1034,N_495);
or U2828 (N_2828,N_1278,N_265);
nor U2829 (N_2829,N_1143,N_1167);
nand U2830 (N_2830,N_1175,N_150);
xnor U2831 (N_2831,N_296,N_1889);
and U2832 (N_2832,N_1488,N_274);
and U2833 (N_2833,N_1423,N_1543);
or U2834 (N_2834,N_1505,N_496);
and U2835 (N_2835,N_1866,N_650);
nand U2836 (N_2836,N_1709,N_799);
xnor U2837 (N_2837,N_1224,N_767);
nor U2838 (N_2838,N_933,N_2);
or U2839 (N_2839,N_1660,N_536);
or U2840 (N_2840,N_1046,N_1244);
xnor U2841 (N_2841,N_842,N_861);
nor U2842 (N_2842,N_1618,N_778);
xor U2843 (N_2843,N_78,N_101);
nand U2844 (N_2844,N_910,N_812);
or U2845 (N_2845,N_461,N_1930);
nand U2846 (N_2846,N_67,N_1131);
or U2847 (N_2847,N_1997,N_410);
xor U2848 (N_2848,N_901,N_629);
nand U2849 (N_2849,N_565,N_218);
nor U2850 (N_2850,N_1035,N_1031);
and U2851 (N_2851,N_1461,N_895);
and U2852 (N_2852,N_423,N_1735);
xnor U2853 (N_2853,N_1162,N_770);
nand U2854 (N_2854,N_1796,N_399);
and U2855 (N_2855,N_1264,N_1787);
nand U2856 (N_2856,N_1651,N_801);
and U2857 (N_2857,N_412,N_71);
or U2858 (N_2858,N_120,N_1193);
nor U2859 (N_2859,N_786,N_1778);
and U2860 (N_2860,N_1424,N_953);
nand U2861 (N_2861,N_1239,N_1079);
or U2862 (N_2862,N_1472,N_1967);
nor U2863 (N_2863,N_141,N_757);
and U2864 (N_2864,N_105,N_1230);
xor U2865 (N_2865,N_1189,N_557);
or U2866 (N_2866,N_1586,N_760);
nand U2867 (N_2867,N_1041,N_1518);
or U2868 (N_2868,N_1257,N_1196);
xor U2869 (N_2869,N_641,N_834);
or U2870 (N_2870,N_1240,N_322);
or U2871 (N_2871,N_1182,N_875);
and U2872 (N_2872,N_845,N_1411);
nor U2873 (N_2873,N_707,N_1066);
nor U2874 (N_2874,N_413,N_211);
or U2875 (N_2875,N_123,N_1077);
and U2876 (N_2876,N_849,N_1671);
and U2877 (N_2877,N_1627,N_1148);
or U2878 (N_2878,N_351,N_1663);
nor U2879 (N_2879,N_1556,N_463);
xor U2880 (N_2880,N_1640,N_1165);
and U2881 (N_2881,N_259,N_1011);
xnor U2882 (N_2882,N_917,N_1407);
and U2883 (N_2883,N_1487,N_301);
nor U2884 (N_2884,N_89,N_1916);
nand U2885 (N_2885,N_1623,N_510);
or U2886 (N_2886,N_591,N_1409);
and U2887 (N_2887,N_858,N_820);
xnor U2888 (N_2888,N_1018,N_98);
nor U2889 (N_2889,N_968,N_686);
nand U2890 (N_2890,N_88,N_1852);
nand U2891 (N_2891,N_46,N_831);
and U2892 (N_2892,N_83,N_1808);
nor U2893 (N_2893,N_12,N_264);
or U2894 (N_2894,N_740,N_1544);
or U2895 (N_2895,N_479,N_1534);
or U2896 (N_2896,N_287,N_989);
or U2897 (N_2897,N_319,N_465);
or U2898 (N_2898,N_1604,N_1685);
and U2899 (N_2899,N_166,N_545);
nor U2900 (N_2900,N_839,N_854);
or U2901 (N_2901,N_566,N_1750);
and U2902 (N_2902,N_852,N_1322);
nand U2903 (N_2903,N_560,N_332);
and U2904 (N_2904,N_1201,N_890);
nand U2905 (N_2905,N_1128,N_651);
or U2906 (N_2906,N_1082,N_1138);
or U2907 (N_2907,N_620,N_1057);
and U2908 (N_2908,N_832,N_1989);
nor U2909 (N_2909,N_1448,N_1665);
nor U2910 (N_2910,N_794,N_146);
and U2911 (N_2911,N_787,N_1876);
or U2912 (N_2912,N_1005,N_1404);
or U2913 (N_2913,N_589,N_1988);
nand U2914 (N_2914,N_518,N_648);
or U2915 (N_2915,N_1410,N_1169);
xnor U2916 (N_2916,N_327,N_57);
xnor U2917 (N_2917,N_984,N_1673);
xor U2918 (N_2918,N_1545,N_1330);
and U2919 (N_2919,N_215,N_1155);
or U2920 (N_2920,N_1053,N_741);
or U2921 (N_2921,N_1655,N_210);
nand U2922 (N_2922,N_610,N_897);
nor U2923 (N_2923,N_1826,N_1744);
and U2924 (N_2924,N_1973,N_899);
and U2925 (N_2925,N_1048,N_1697);
nand U2926 (N_2926,N_1806,N_1211);
nand U2927 (N_2927,N_1374,N_973);
xnor U2928 (N_2928,N_1725,N_867);
or U2929 (N_2929,N_1150,N_340);
and U2930 (N_2930,N_511,N_1914);
nor U2931 (N_2931,N_1877,N_900);
nor U2932 (N_2932,N_601,N_243);
nor U2933 (N_2933,N_1800,N_1674);
nand U2934 (N_2934,N_476,N_916);
nand U2935 (N_2935,N_1418,N_1657);
xnor U2936 (N_2936,N_594,N_826);
nor U2937 (N_2937,N_1450,N_1934);
or U2938 (N_2938,N_227,N_1419);
nand U2939 (N_2939,N_1061,N_1548);
or U2940 (N_2940,N_1400,N_122);
nor U2941 (N_2941,N_1566,N_830);
or U2942 (N_2942,N_1522,N_1354);
xnor U2943 (N_2943,N_349,N_1428);
nand U2944 (N_2944,N_885,N_446);
and U2945 (N_2945,N_100,N_689);
or U2946 (N_2946,N_731,N_415);
nor U2947 (N_2947,N_255,N_1337);
or U2948 (N_2948,N_1435,N_237);
nor U2949 (N_2949,N_183,N_1677);
nand U2950 (N_2950,N_521,N_1884);
nor U2951 (N_2951,N_1948,N_729);
nor U2952 (N_2952,N_553,N_537);
nand U2953 (N_2953,N_26,N_625);
nor U2954 (N_2954,N_1298,N_1885);
and U2955 (N_2955,N_400,N_336);
and U2956 (N_2956,N_1248,N_276);
and U2957 (N_2957,N_1875,N_1842);
and U2958 (N_2958,N_1255,N_206);
nor U2959 (N_2959,N_1103,N_600);
or U2960 (N_2960,N_385,N_1931);
nand U2961 (N_2961,N_1449,N_639);
or U2962 (N_2962,N_1164,N_1249);
nand U2963 (N_2963,N_878,N_1943);
nand U2964 (N_2964,N_815,N_713);
or U2965 (N_2965,N_1616,N_784);
nor U2966 (N_2966,N_493,N_1290);
nand U2967 (N_2967,N_1163,N_690);
xor U2968 (N_2968,N_1200,N_76);
or U2969 (N_2969,N_1594,N_1902);
nand U2970 (N_2970,N_1741,N_459);
or U2971 (N_2971,N_979,N_599);
or U2972 (N_2972,N_604,N_626);
and U2973 (N_2973,N_1497,N_735);
nor U2974 (N_2974,N_669,N_1878);
nor U2975 (N_2975,N_1968,N_344);
or U2976 (N_2976,N_1421,N_1465);
and U2977 (N_2977,N_1861,N_941);
or U2978 (N_2978,N_127,N_1529);
nand U2979 (N_2979,N_1588,N_632);
nor U2980 (N_2980,N_1210,N_774);
or U2981 (N_2981,N_1802,N_756);
xnor U2982 (N_2982,N_906,N_1922);
or U2983 (N_2983,N_1022,N_455);
nand U2984 (N_2984,N_1121,N_305);
nand U2985 (N_2985,N_1991,N_1514);
nand U2986 (N_2986,N_1521,N_1888);
nand U2987 (N_2987,N_1190,N_1329);
and U2988 (N_2988,N_1886,N_1282);
nand U2989 (N_2989,N_440,N_1440);
and U2990 (N_2990,N_1089,N_492);
or U2991 (N_2991,N_656,N_611);
and U2992 (N_2992,N_1557,N_539);
and U2993 (N_2993,N_1734,N_1049);
nor U2994 (N_2994,N_1453,N_751);
or U2995 (N_2995,N_1033,N_1681);
or U2996 (N_2996,N_549,N_1217);
or U2997 (N_2997,N_640,N_733);
and U2998 (N_2998,N_1939,N_448);
or U2999 (N_2999,N_409,N_1776);
xor U3000 (N_3000,N_833,N_1675);
nor U3001 (N_3001,N_1986,N_395);
or U3002 (N_3002,N_1660,N_1395);
and U3003 (N_3003,N_470,N_992);
nor U3004 (N_3004,N_268,N_317);
nor U3005 (N_3005,N_1306,N_1920);
nand U3006 (N_3006,N_349,N_1978);
nand U3007 (N_3007,N_1463,N_797);
nor U3008 (N_3008,N_112,N_1467);
nor U3009 (N_3009,N_1545,N_1167);
or U3010 (N_3010,N_299,N_1653);
nand U3011 (N_3011,N_1829,N_1069);
nand U3012 (N_3012,N_105,N_1015);
and U3013 (N_3013,N_1257,N_623);
and U3014 (N_3014,N_1057,N_1760);
and U3015 (N_3015,N_1235,N_1328);
nor U3016 (N_3016,N_1255,N_1802);
nor U3017 (N_3017,N_1434,N_132);
or U3018 (N_3018,N_1897,N_455);
nand U3019 (N_3019,N_1509,N_1285);
or U3020 (N_3020,N_1266,N_537);
or U3021 (N_3021,N_796,N_171);
nand U3022 (N_3022,N_494,N_1664);
nand U3023 (N_3023,N_544,N_253);
nor U3024 (N_3024,N_169,N_921);
nand U3025 (N_3025,N_203,N_491);
or U3026 (N_3026,N_283,N_1330);
and U3027 (N_3027,N_1184,N_1784);
xor U3028 (N_3028,N_797,N_5);
or U3029 (N_3029,N_1538,N_61);
and U3030 (N_3030,N_1201,N_806);
xnor U3031 (N_3031,N_1622,N_1553);
or U3032 (N_3032,N_1250,N_1887);
xor U3033 (N_3033,N_1869,N_949);
or U3034 (N_3034,N_1013,N_101);
nand U3035 (N_3035,N_1406,N_241);
and U3036 (N_3036,N_1337,N_830);
nor U3037 (N_3037,N_503,N_1614);
nor U3038 (N_3038,N_1662,N_1674);
or U3039 (N_3039,N_1955,N_1611);
and U3040 (N_3040,N_1530,N_1477);
or U3041 (N_3041,N_531,N_697);
nor U3042 (N_3042,N_1113,N_1356);
nor U3043 (N_3043,N_492,N_1948);
nand U3044 (N_3044,N_993,N_1345);
or U3045 (N_3045,N_122,N_1701);
or U3046 (N_3046,N_758,N_985);
xor U3047 (N_3047,N_747,N_717);
nand U3048 (N_3048,N_872,N_951);
nand U3049 (N_3049,N_211,N_1811);
nor U3050 (N_3050,N_413,N_1811);
nor U3051 (N_3051,N_1030,N_1186);
nor U3052 (N_3052,N_1537,N_1767);
and U3053 (N_3053,N_891,N_1257);
nor U3054 (N_3054,N_248,N_1519);
nand U3055 (N_3055,N_419,N_524);
nand U3056 (N_3056,N_217,N_323);
and U3057 (N_3057,N_633,N_842);
nor U3058 (N_3058,N_1059,N_957);
and U3059 (N_3059,N_1377,N_911);
nor U3060 (N_3060,N_1924,N_1257);
and U3061 (N_3061,N_364,N_1046);
and U3062 (N_3062,N_1822,N_1740);
xor U3063 (N_3063,N_1786,N_1476);
or U3064 (N_3064,N_437,N_436);
or U3065 (N_3065,N_193,N_1326);
and U3066 (N_3066,N_303,N_731);
and U3067 (N_3067,N_1283,N_728);
or U3068 (N_3068,N_1484,N_362);
and U3069 (N_3069,N_209,N_1455);
nor U3070 (N_3070,N_1391,N_1466);
nand U3071 (N_3071,N_4,N_1006);
and U3072 (N_3072,N_444,N_999);
nand U3073 (N_3073,N_198,N_1163);
nor U3074 (N_3074,N_1222,N_275);
xor U3075 (N_3075,N_120,N_1814);
nor U3076 (N_3076,N_1963,N_588);
nand U3077 (N_3077,N_679,N_1109);
nor U3078 (N_3078,N_1153,N_346);
nor U3079 (N_3079,N_138,N_944);
or U3080 (N_3080,N_1210,N_1845);
nand U3081 (N_3081,N_900,N_1897);
xnor U3082 (N_3082,N_1341,N_1698);
and U3083 (N_3083,N_1078,N_377);
nor U3084 (N_3084,N_1900,N_1027);
xnor U3085 (N_3085,N_107,N_1051);
nand U3086 (N_3086,N_1878,N_1674);
nand U3087 (N_3087,N_1121,N_1796);
xor U3088 (N_3088,N_1762,N_944);
and U3089 (N_3089,N_1585,N_842);
or U3090 (N_3090,N_787,N_1145);
or U3091 (N_3091,N_1368,N_566);
nor U3092 (N_3092,N_986,N_767);
nand U3093 (N_3093,N_240,N_1449);
and U3094 (N_3094,N_1135,N_21);
and U3095 (N_3095,N_316,N_1599);
nand U3096 (N_3096,N_1157,N_1423);
nor U3097 (N_3097,N_1367,N_255);
or U3098 (N_3098,N_347,N_1336);
or U3099 (N_3099,N_287,N_1351);
nor U3100 (N_3100,N_337,N_1599);
or U3101 (N_3101,N_1307,N_1604);
or U3102 (N_3102,N_177,N_1323);
or U3103 (N_3103,N_1054,N_30);
or U3104 (N_3104,N_1475,N_440);
nor U3105 (N_3105,N_354,N_364);
nor U3106 (N_3106,N_102,N_1142);
or U3107 (N_3107,N_259,N_692);
and U3108 (N_3108,N_1726,N_1519);
nor U3109 (N_3109,N_1345,N_1701);
nor U3110 (N_3110,N_50,N_1350);
nor U3111 (N_3111,N_1365,N_852);
xnor U3112 (N_3112,N_91,N_1923);
nor U3113 (N_3113,N_280,N_289);
nand U3114 (N_3114,N_415,N_1899);
xnor U3115 (N_3115,N_1331,N_1237);
and U3116 (N_3116,N_1426,N_372);
nand U3117 (N_3117,N_1874,N_910);
or U3118 (N_3118,N_350,N_877);
xor U3119 (N_3119,N_701,N_1457);
nor U3120 (N_3120,N_929,N_769);
and U3121 (N_3121,N_1090,N_1330);
nor U3122 (N_3122,N_500,N_1976);
and U3123 (N_3123,N_970,N_1437);
nor U3124 (N_3124,N_1567,N_937);
and U3125 (N_3125,N_247,N_1404);
and U3126 (N_3126,N_363,N_1699);
and U3127 (N_3127,N_74,N_1903);
nor U3128 (N_3128,N_1344,N_1501);
xor U3129 (N_3129,N_1964,N_1888);
nand U3130 (N_3130,N_666,N_1689);
and U3131 (N_3131,N_926,N_473);
nor U3132 (N_3132,N_271,N_1758);
nand U3133 (N_3133,N_811,N_1361);
nand U3134 (N_3134,N_487,N_1415);
nand U3135 (N_3135,N_1826,N_80);
xnor U3136 (N_3136,N_1499,N_499);
nor U3137 (N_3137,N_695,N_1683);
and U3138 (N_3138,N_727,N_1311);
xor U3139 (N_3139,N_421,N_1610);
xor U3140 (N_3140,N_1883,N_1520);
and U3141 (N_3141,N_1603,N_545);
nor U3142 (N_3142,N_551,N_1383);
and U3143 (N_3143,N_93,N_988);
nand U3144 (N_3144,N_638,N_130);
nand U3145 (N_3145,N_1301,N_1096);
and U3146 (N_3146,N_1180,N_658);
and U3147 (N_3147,N_145,N_1381);
nand U3148 (N_3148,N_1336,N_1759);
nor U3149 (N_3149,N_451,N_1127);
and U3150 (N_3150,N_463,N_44);
or U3151 (N_3151,N_243,N_1837);
or U3152 (N_3152,N_1010,N_1839);
nand U3153 (N_3153,N_1919,N_663);
nand U3154 (N_3154,N_1522,N_1180);
nand U3155 (N_3155,N_1597,N_440);
or U3156 (N_3156,N_865,N_542);
nand U3157 (N_3157,N_543,N_1920);
or U3158 (N_3158,N_1405,N_1916);
or U3159 (N_3159,N_420,N_1706);
nor U3160 (N_3160,N_961,N_1365);
nor U3161 (N_3161,N_889,N_641);
nand U3162 (N_3162,N_1913,N_1825);
nor U3163 (N_3163,N_284,N_1680);
or U3164 (N_3164,N_125,N_1674);
nand U3165 (N_3165,N_1207,N_866);
nand U3166 (N_3166,N_75,N_796);
or U3167 (N_3167,N_1368,N_279);
xnor U3168 (N_3168,N_186,N_262);
nand U3169 (N_3169,N_501,N_1838);
nor U3170 (N_3170,N_766,N_1399);
nand U3171 (N_3171,N_468,N_934);
xor U3172 (N_3172,N_1212,N_1262);
nand U3173 (N_3173,N_1730,N_459);
nand U3174 (N_3174,N_723,N_591);
or U3175 (N_3175,N_1565,N_1267);
nor U3176 (N_3176,N_1998,N_920);
nor U3177 (N_3177,N_984,N_641);
nand U3178 (N_3178,N_1079,N_864);
and U3179 (N_3179,N_190,N_1600);
or U3180 (N_3180,N_1589,N_1502);
nand U3181 (N_3181,N_9,N_654);
or U3182 (N_3182,N_17,N_1042);
xnor U3183 (N_3183,N_107,N_1129);
nor U3184 (N_3184,N_1853,N_935);
nand U3185 (N_3185,N_741,N_1017);
nor U3186 (N_3186,N_1748,N_1182);
or U3187 (N_3187,N_1815,N_1765);
xor U3188 (N_3188,N_1954,N_824);
nor U3189 (N_3189,N_328,N_280);
nand U3190 (N_3190,N_684,N_577);
or U3191 (N_3191,N_265,N_82);
nand U3192 (N_3192,N_185,N_1059);
nor U3193 (N_3193,N_1589,N_1781);
nor U3194 (N_3194,N_731,N_1012);
nor U3195 (N_3195,N_111,N_1036);
or U3196 (N_3196,N_406,N_1931);
nor U3197 (N_3197,N_1034,N_1380);
nand U3198 (N_3198,N_1793,N_1598);
nand U3199 (N_3199,N_504,N_256);
nand U3200 (N_3200,N_1448,N_19);
nand U3201 (N_3201,N_1925,N_679);
and U3202 (N_3202,N_1343,N_1534);
nor U3203 (N_3203,N_464,N_1746);
nor U3204 (N_3204,N_584,N_552);
nor U3205 (N_3205,N_1442,N_1026);
and U3206 (N_3206,N_227,N_1431);
and U3207 (N_3207,N_1808,N_659);
or U3208 (N_3208,N_562,N_1362);
nor U3209 (N_3209,N_1694,N_1747);
and U3210 (N_3210,N_348,N_25);
or U3211 (N_3211,N_318,N_1379);
nor U3212 (N_3212,N_1426,N_132);
nand U3213 (N_3213,N_166,N_289);
and U3214 (N_3214,N_714,N_461);
xor U3215 (N_3215,N_595,N_1125);
or U3216 (N_3216,N_437,N_1267);
xor U3217 (N_3217,N_1134,N_1291);
nor U3218 (N_3218,N_36,N_243);
and U3219 (N_3219,N_1059,N_751);
nor U3220 (N_3220,N_499,N_1151);
xnor U3221 (N_3221,N_261,N_486);
xnor U3222 (N_3222,N_77,N_1880);
or U3223 (N_3223,N_1242,N_786);
xor U3224 (N_3224,N_184,N_1950);
nand U3225 (N_3225,N_32,N_1130);
nor U3226 (N_3226,N_153,N_459);
and U3227 (N_3227,N_1679,N_1793);
or U3228 (N_3228,N_1357,N_351);
nand U3229 (N_3229,N_1690,N_1519);
nor U3230 (N_3230,N_783,N_1587);
nand U3231 (N_3231,N_893,N_761);
nand U3232 (N_3232,N_616,N_683);
and U3233 (N_3233,N_1135,N_1117);
or U3234 (N_3234,N_1994,N_984);
and U3235 (N_3235,N_912,N_1638);
xor U3236 (N_3236,N_38,N_1786);
nand U3237 (N_3237,N_1872,N_645);
and U3238 (N_3238,N_345,N_178);
or U3239 (N_3239,N_1429,N_515);
or U3240 (N_3240,N_1519,N_1746);
and U3241 (N_3241,N_1278,N_1374);
nor U3242 (N_3242,N_1329,N_978);
and U3243 (N_3243,N_410,N_417);
nand U3244 (N_3244,N_370,N_1056);
xnor U3245 (N_3245,N_1760,N_1331);
nor U3246 (N_3246,N_982,N_616);
or U3247 (N_3247,N_448,N_286);
and U3248 (N_3248,N_1500,N_70);
and U3249 (N_3249,N_1512,N_1182);
xor U3250 (N_3250,N_1854,N_1488);
or U3251 (N_3251,N_476,N_1584);
and U3252 (N_3252,N_1228,N_1222);
xor U3253 (N_3253,N_731,N_1830);
or U3254 (N_3254,N_929,N_427);
or U3255 (N_3255,N_1892,N_1630);
or U3256 (N_3256,N_620,N_1696);
xor U3257 (N_3257,N_66,N_1699);
or U3258 (N_3258,N_1993,N_1445);
nor U3259 (N_3259,N_1762,N_1676);
nor U3260 (N_3260,N_149,N_1983);
and U3261 (N_3261,N_1071,N_1224);
xnor U3262 (N_3262,N_202,N_1928);
nor U3263 (N_3263,N_1797,N_844);
xnor U3264 (N_3264,N_141,N_1302);
xnor U3265 (N_3265,N_1021,N_535);
nor U3266 (N_3266,N_1637,N_559);
nor U3267 (N_3267,N_1741,N_1521);
nand U3268 (N_3268,N_919,N_1152);
nand U3269 (N_3269,N_452,N_1537);
xor U3270 (N_3270,N_1082,N_1442);
or U3271 (N_3271,N_1185,N_964);
and U3272 (N_3272,N_1052,N_831);
or U3273 (N_3273,N_1566,N_1497);
nand U3274 (N_3274,N_275,N_1622);
or U3275 (N_3275,N_234,N_1469);
and U3276 (N_3276,N_672,N_276);
nand U3277 (N_3277,N_1345,N_1977);
nor U3278 (N_3278,N_256,N_1441);
nor U3279 (N_3279,N_1773,N_1699);
nand U3280 (N_3280,N_83,N_1034);
nor U3281 (N_3281,N_460,N_1250);
nand U3282 (N_3282,N_643,N_1942);
and U3283 (N_3283,N_1325,N_1406);
nor U3284 (N_3284,N_934,N_60);
nor U3285 (N_3285,N_1591,N_1193);
nand U3286 (N_3286,N_1534,N_1794);
nor U3287 (N_3287,N_646,N_1750);
nor U3288 (N_3288,N_59,N_522);
nor U3289 (N_3289,N_1369,N_1681);
xnor U3290 (N_3290,N_499,N_692);
and U3291 (N_3291,N_1866,N_86);
or U3292 (N_3292,N_167,N_1048);
and U3293 (N_3293,N_273,N_1787);
or U3294 (N_3294,N_1653,N_995);
or U3295 (N_3295,N_938,N_509);
and U3296 (N_3296,N_1073,N_1618);
xnor U3297 (N_3297,N_1406,N_815);
and U3298 (N_3298,N_829,N_1460);
nand U3299 (N_3299,N_84,N_1893);
and U3300 (N_3300,N_1063,N_753);
xnor U3301 (N_3301,N_1821,N_104);
or U3302 (N_3302,N_1786,N_143);
and U3303 (N_3303,N_790,N_219);
and U3304 (N_3304,N_1331,N_878);
and U3305 (N_3305,N_626,N_1038);
nand U3306 (N_3306,N_634,N_272);
and U3307 (N_3307,N_1670,N_630);
xnor U3308 (N_3308,N_962,N_333);
or U3309 (N_3309,N_399,N_838);
and U3310 (N_3310,N_1881,N_316);
nor U3311 (N_3311,N_1536,N_1721);
nand U3312 (N_3312,N_1571,N_348);
or U3313 (N_3313,N_994,N_537);
and U3314 (N_3314,N_1668,N_677);
nor U3315 (N_3315,N_839,N_1537);
and U3316 (N_3316,N_872,N_1543);
nor U3317 (N_3317,N_796,N_886);
nand U3318 (N_3318,N_971,N_1079);
nor U3319 (N_3319,N_606,N_1648);
xnor U3320 (N_3320,N_1131,N_1441);
nand U3321 (N_3321,N_569,N_1477);
or U3322 (N_3322,N_1263,N_1203);
or U3323 (N_3323,N_803,N_876);
xor U3324 (N_3324,N_1254,N_1907);
and U3325 (N_3325,N_931,N_517);
or U3326 (N_3326,N_792,N_532);
nor U3327 (N_3327,N_663,N_44);
nor U3328 (N_3328,N_231,N_1385);
nand U3329 (N_3329,N_1743,N_861);
nand U3330 (N_3330,N_1609,N_549);
nand U3331 (N_3331,N_1280,N_574);
and U3332 (N_3332,N_144,N_727);
nand U3333 (N_3333,N_1601,N_1016);
or U3334 (N_3334,N_1395,N_83);
or U3335 (N_3335,N_847,N_1621);
nor U3336 (N_3336,N_1654,N_787);
nor U3337 (N_3337,N_96,N_1185);
and U3338 (N_3338,N_59,N_1929);
or U3339 (N_3339,N_505,N_1855);
xor U3340 (N_3340,N_796,N_92);
xnor U3341 (N_3341,N_246,N_1139);
xnor U3342 (N_3342,N_66,N_914);
or U3343 (N_3343,N_909,N_1055);
or U3344 (N_3344,N_305,N_90);
nor U3345 (N_3345,N_1955,N_1074);
nand U3346 (N_3346,N_783,N_616);
and U3347 (N_3347,N_974,N_1962);
xor U3348 (N_3348,N_521,N_610);
nand U3349 (N_3349,N_1643,N_1186);
nand U3350 (N_3350,N_370,N_703);
or U3351 (N_3351,N_214,N_515);
xnor U3352 (N_3352,N_178,N_1653);
nand U3353 (N_3353,N_320,N_106);
nor U3354 (N_3354,N_1848,N_1790);
nor U3355 (N_3355,N_1078,N_517);
nand U3356 (N_3356,N_696,N_364);
and U3357 (N_3357,N_675,N_1027);
and U3358 (N_3358,N_1599,N_1208);
nor U3359 (N_3359,N_564,N_1931);
and U3360 (N_3360,N_1462,N_1656);
nand U3361 (N_3361,N_527,N_1906);
nor U3362 (N_3362,N_1764,N_567);
or U3363 (N_3363,N_179,N_728);
and U3364 (N_3364,N_645,N_526);
nand U3365 (N_3365,N_532,N_1480);
nand U3366 (N_3366,N_423,N_1539);
xnor U3367 (N_3367,N_1306,N_1059);
or U3368 (N_3368,N_1153,N_844);
nor U3369 (N_3369,N_1562,N_1511);
and U3370 (N_3370,N_1151,N_1613);
xnor U3371 (N_3371,N_1480,N_1103);
nand U3372 (N_3372,N_795,N_172);
nor U3373 (N_3373,N_948,N_1918);
and U3374 (N_3374,N_1431,N_338);
nand U3375 (N_3375,N_1027,N_222);
xnor U3376 (N_3376,N_1675,N_468);
nor U3377 (N_3377,N_543,N_465);
nand U3378 (N_3378,N_1869,N_1486);
nand U3379 (N_3379,N_1784,N_1664);
nand U3380 (N_3380,N_1343,N_1949);
and U3381 (N_3381,N_1728,N_1384);
xnor U3382 (N_3382,N_658,N_322);
and U3383 (N_3383,N_927,N_308);
and U3384 (N_3384,N_1156,N_788);
nor U3385 (N_3385,N_470,N_654);
nand U3386 (N_3386,N_1497,N_1828);
nor U3387 (N_3387,N_1581,N_68);
nor U3388 (N_3388,N_1451,N_48);
xor U3389 (N_3389,N_1881,N_1985);
or U3390 (N_3390,N_1227,N_1092);
xor U3391 (N_3391,N_897,N_1836);
and U3392 (N_3392,N_82,N_553);
nand U3393 (N_3393,N_1427,N_881);
and U3394 (N_3394,N_127,N_421);
and U3395 (N_3395,N_1633,N_1689);
and U3396 (N_3396,N_1067,N_7);
nor U3397 (N_3397,N_508,N_276);
nor U3398 (N_3398,N_531,N_146);
and U3399 (N_3399,N_756,N_463);
or U3400 (N_3400,N_1701,N_396);
nand U3401 (N_3401,N_371,N_1542);
nand U3402 (N_3402,N_107,N_1982);
or U3403 (N_3403,N_365,N_1528);
and U3404 (N_3404,N_1129,N_305);
xnor U3405 (N_3405,N_532,N_1107);
nand U3406 (N_3406,N_1298,N_1665);
nor U3407 (N_3407,N_1666,N_996);
and U3408 (N_3408,N_1399,N_591);
and U3409 (N_3409,N_1014,N_1591);
or U3410 (N_3410,N_561,N_862);
nand U3411 (N_3411,N_1417,N_365);
and U3412 (N_3412,N_53,N_1661);
nor U3413 (N_3413,N_393,N_70);
and U3414 (N_3414,N_1212,N_158);
nor U3415 (N_3415,N_1668,N_4);
and U3416 (N_3416,N_728,N_731);
xnor U3417 (N_3417,N_1310,N_116);
nand U3418 (N_3418,N_1929,N_71);
nand U3419 (N_3419,N_513,N_1450);
nor U3420 (N_3420,N_168,N_1365);
and U3421 (N_3421,N_1413,N_1127);
or U3422 (N_3422,N_799,N_1674);
or U3423 (N_3423,N_700,N_920);
or U3424 (N_3424,N_1331,N_1103);
and U3425 (N_3425,N_1028,N_748);
nor U3426 (N_3426,N_1605,N_716);
nor U3427 (N_3427,N_0,N_1260);
or U3428 (N_3428,N_58,N_1492);
or U3429 (N_3429,N_162,N_335);
xor U3430 (N_3430,N_1793,N_419);
xor U3431 (N_3431,N_1864,N_827);
nor U3432 (N_3432,N_1993,N_408);
nor U3433 (N_3433,N_186,N_960);
nand U3434 (N_3434,N_1023,N_931);
nor U3435 (N_3435,N_650,N_642);
nor U3436 (N_3436,N_21,N_1434);
nor U3437 (N_3437,N_894,N_1113);
xor U3438 (N_3438,N_755,N_433);
nor U3439 (N_3439,N_695,N_21);
xnor U3440 (N_3440,N_229,N_1640);
nand U3441 (N_3441,N_1320,N_1967);
nor U3442 (N_3442,N_1432,N_1192);
nand U3443 (N_3443,N_158,N_750);
and U3444 (N_3444,N_159,N_1073);
or U3445 (N_3445,N_1070,N_1385);
nand U3446 (N_3446,N_1429,N_135);
nor U3447 (N_3447,N_99,N_138);
nand U3448 (N_3448,N_1317,N_397);
nand U3449 (N_3449,N_1816,N_7);
nand U3450 (N_3450,N_476,N_1335);
or U3451 (N_3451,N_1614,N_530);
and U3452 (N_3452,N_118,N_1272);
or U3453 (N_3453,N_1620,N_1958);
nor U3454 (N_3454,N_441,N_1352);
nand U3455 (N_3455,N_144,N_1605);
and U3456 (N_3456,N_1963,N_1147);
nand U3457 (N_3457,N_432,N_768);
xor U3458 (N_3458,N_1093,N_476);
or U3459 (N_3459,N_1843,N_1260);
nor U3460 (N_3460,N_1346,N_1457);
nor U3461 (N_3461,N_1678,N_944);
or U3462 (N_3462,N_911,N_1164);
nor U3463 (N_3463,N_803,N_607);
or U3464 (N_3464,N_514,N_1475);
nand U3465 (N_3465,N_1935,N_1832);
nor U3466 (N_3466,N_1581,N_306);
xnor U3467 (N_3467,N_1424,N_1914);
nor U3468 (N_3468,N_1202,N_1809);
or U3469 (N_3469,N_162,N_548);
xor U3470 (N_3470,N_1464,N_749);
and U3471 (N_3471,N_1470,N_258);
nand U3472 (N_3472,N_477,N_862);
nand U3473 (N_3473,N_1447,N_1129);
nand U3474 (N_3474,N_937,N_1901);
nand U3475 (N_3475,N_813,N_1693);
nand U3476 (N_3476,N_494,N_479);
nand U3477 (N_3477,N_799,N_210);
xor U3478 (N_3478,N_1200,N_724);
nor U3479 (N_3479,N_1165,N_925);
nand U3480 (N_3480,N_1385,N_206);
xnor U3481 (N_3481,N_1517,N_1092);
nor U3482 (N_3482,N_1206,N_94);
or U3483 (N_3483,N_1750,N_19);
and U3484 (N_3484,N_1812,N_475);
and U3485 (N_3485,N_407,N_466);
and U3486 (N_3486,N_1775,N_671);
or U3487 (N_3487,N_1085,N_1700);
nor U3488 (N_3488,N_1301,N_1348);
or U3489 (N_3489,N_1731,N_770);
and U3490 (N_3490,N_178,N_547);
and U3491 (N_3491,N_363,N_108);
and U3492 (N_3492,N_1523,N_781);
nand U3493 (N_3493,N_1826,N_1282);
nor U3494 (N_3494,N_1758,N_391);
nor U3495 (N_3495,N_668,N_729);
nand U3496 (N_3496,N_1549,N_1902);
and U3497 (N_3497,N_719,N_1549);
xor U3498 (N_3498,N_938,N_905);
nand U3499 (N_3499,N_746,N_193);
and U3500 (N_3500,N_401,N_994);
nor U3501 (N_3501,N_356,N_65);
nand U3502 (N_3502,N_1267,N_1668);
and U3503 (N_3503,N_1634,N_656);
nand U3504 (N_3504,N_1809,N_993);
and U3505 (N_3505,N_1682,N_1360);
or U3506 (N_3506,N_1135,N_1377);
and U3507 (N_3507,N_610,N_1215);
or U3508 (N_3508,N_458,N_435);
or U3509 (N_3509,N_1307,N_1204);
or U3510 (N_3510,N_166,N_900);
nand U3511 (N_3511,N_1341,N_335);
nor U3512 (N_3512,N_776,N_867);
nand U3513 (N_3513,N_71,N_488);
or U3514 (N_3514,N_1495,N_1803);
and U3515 (N_3515,N_1270,N_1736);
nor U3516 (N_3516,N_1436,N_294);
or U3517 (N_3517,N_1389,N_1524);
nand U3518 (N_3518,N_635,N_1818);
nand U3519 (N_3519,N_517,N_801);
nand U3520 (N_3520,N_473,N_1415);
nor U3521 (N_3521,N_783,N_66);
and U3522 (N_3522,N_1541,N_1868);
and U3523 (N_3523,N_1020,N_936);
nor U3524 (N_3524,N_639,N_730);
and U3525 (N_3525,N_1610,N_617);
or U3526 (N_3526,N_201,N_1991);
nor U3527 (N_3527,N_1551,N_185);
or U3528 (N_3528,N_773,N_1825);
and U3529 (N_3529,N_1075,N_605);
or U3530 (N_3530,N_291,N_107);
nand U3531 (N_3531,N_160,N_207);
xnor U3532 (N_3532,N_1940,N_1261);
or U3533 (N_3533,N_491,N_853);
nand U3534 (N_3534,N_1461,N_929);
nand U3535 (N_3535,N_1792,N_1165);
xnor U3536 (N_3536,N_1917,N_798);
nor U3537 (N_3537,N_528,N_701);
nand U3538 (N_3538,N_1970,N_1595);
nand U3539 (N_3539,N_423,N_1960);
nor U3540 (N_3540,N_1424,N_1258);
xnor U3541 (N_3541,N_460,N_1048);
xor U3542 (N_3542,N_819,N_1753);
or U3543 (N_3543,N_842,N_509);
and U3544 (N_3544,N_983,N_560);
nand U3545 (N_3545,N_907,N_1312);
nand U3546 (N_3546,N_1086,N_1349);
and U3547 (N_3547,N_148,N_526);
or U3548 (N_3548,N_777,N_77);
or U3549 (N_3549,N_1396,N_1294);
and U3550 (N_3550,N_1776,N_871);
nor U3551 (N_3551,N_1826,N_512);
or U3552 (N_3552,N_350,N_1747);
xor U3553 (N_3553,N_1940,N_188);
xnor U3554 (N_3554,N_493,N_1164);
and U3555 (N_3555,N_1763,N_1109);
or U3556 (N_3556,N_817,N_165);
or U3557 (N_3557,N_1749,N_1017);
and U3558 (N_3558,N_1020,N_183);
nand U3559 (N_3559,N_348,N_104);
and U3560 (N_3560,N_1719,N_1883);
xnor U3561 (N_3561,N_781,N_18);
nor U3562 (N_3562,N_1036,N_258);
xnor U3563 (N_3563,N_89,N_452);
and U3564 (N_3564,N_194,N_830);
nor U3565 (N_3565,N_1028,N_40);
xor U3566 (N_3566,N_589,N_145);
nor U3567 (N_3567,N_884,N_1190);
nor U3568 (N_3568,N_1121,N_969);
xnor U3569 (N_3569,N_962,N_792);
and U3570 (N_3570,N_1368,N_330);
or U3571 (N_3571,N_1780,N_491);
nor U3572 (N_3572,N_735,N_1351);
or U3573 (N_3573,N_1748,N_1839);
xor U3574 (N_3574,N_922,N_1838);
nor U3575 (N_3575,N_1278,N_674);
or U3576 (N_3576,N_1441,N_1673);
or U3577 (N_3577,N_917,N_983);
or U3578 (N_3578,N_675,N_944);
and U3579 (N_3579,N_1057,N_989);
and U3580 (N_3580,N_560,N_1840);
or U3581 (N_3581,N_1166,N_520);
and U3582 (N_3582,N_1732,N_1473);
or U3583 (N_3583,N_725,N_1322);
nor U3584 (N_3584,N_1620,N_481);
nor U3585 (N_3585,N_521,N_1001);
or U3586 (N_3586,N_1390,N_1510);
or U3587 (N_3587,N_179,N_1764);
nand U3588 (N_3588,N_202,N_1763);
nor U3589 (N_3589,N_629,N_584);
or U3590 (N_3590,N_1665,N_334);
or U3591 (N_3591,N_72,N_738);
nor U3592 (N_3592,N_1858,N_1025);
and U3593 (N_3593,N_1748,N_1034);
nor U3594 (N_3594,N_1770,N_1700);
or U3595 (N_3595,N_648,N_852);
xor U3596 (N_3596,N_1310,N_0);
and U3597 (N_3597,N_1290,N_1776);
and U3598 (N_3598,N_700,N_952);
and U3599 (N_3599,N_537,N_1048);
and U3600 (N_3600,N_295,N_560);
nand U3601 (N_3601,N_65,N_1653);
or U3602 (N_3602,N_1990,N_379);
and U3603 (N_3603,N_476,N_1386);
nand U3604 (N_3604,N_221,N_601);
nand U3605 (N_3605,N_891,N_614);
nor U3606 (N_3606,N_502,N_1010);
nand U3607 (N_3607,N_1875,N_511);
and U3608 (N_3608,N_1531,N_1467);
and U3609 (N_3609,N_1066,N_278);
nand U3610 (N_3610,N_1605,N_1672);
xnor U3611 (N_3611,N_1984,N_1627);
or U3612 (N_3612,N_368,N_1978);
nor U3613 (N_3613,N_58,N_1979);
and U3614 (N_3614,N_707,N_1068);
xor U3615 (N_3615,N_575,N_436);
nor U3616 (N_3616,N_880,N_497);
or U3617 (N_3617,N_1714,N_209);
xnor U3618 (N_3618,N_127,N_394);
and U3619 (N_3619,N_659,N_1652);
nand U3620 (N_3620,N_742,N_1419);
nor U3621 (N_3621,N_1382,N_42);
nor U3622 (N_3622,N_160,N_753);
or U3623 (N_3623,N_1947,N_1293);
or U3624 (N_3624,N_850,N_1095);
and U3625 (N_3625,N_918,N_1099);
or U3626 (N_3626,N_1467,N_349);
nor U3627 (N_3627,N_1583,N_1373);
nand U3628 (N_3628,N_1553,N_92);
and U3629 (N_3629,N_1641,N_1102);
nand U3630 (N_3630,N_1624,N_727);
nor U3631 (N_3631,N_1038,N_1075);
and U3632 (N_3632,N_61,N_52);
and U3633 (N_3633,N_1376,N_585);
nor U3634 (N_3634,N_1139,N_1511);
and U3635 (N_3635,N_1992,N_649);
nand U3636 (N_3636,N_140,N_271);
or U3637 (N_3637,N_31,N_879);
nor U3638 (N_3638,N_365,N_34);
or U3639 (N_3639,N_1858,N_1386);
nand U3640 (N_3640,N_98,N_497);
and U3641 (N_3641,N_254,N_1256);
or U3642 (N_3642,N_1039,N_1103);
nor U3643 (N_3643,N_1973,N_989);
and U3644 (N_3644,N_798,N_905);
xnor U3645 (N_3645,N_1629,N_7);
nor U3646 (N_3646,N_1449,N_1134);
nand U3647 (N_3647,N_1345,N_1097);
xor U3648 (N_3648,N_407,N_1125);
and U3649 (N_3649,N_1498,N_78);
or U3650 (N_3650,N_1229,N_575);
nor U3651 (N_3651,N_1369,N_702);
nor U3652 (N_3652,N_191,N_433);
xor U3653 (N_3653,N_933,N_35);
nor U3654 (N_3654,N_561,N_1753);
xnor U3655 (N_3655,N_394,N_1201);
and U3656 (N_3656,N_380,N_1540);
and U3657 (N_3657,N_1118,N_1567);
nand U3658 (N_3658,N_578,N_224);
nand U3659 (N_3659,N_1941,N_983);
or U3660 (N_3660,N_1582,N_646);
nor U3661 (N_3661,N_145,N_1501);
nor U3662 (N_3662,N_933,N_731);
nand U3663 (N_3663,N_806,N_1267);
and U3664 (N_3664,N_219,N_592);
and U3665 (N_3665,N_1413,N_1581);
nor U3666 (N_3666,N_440,N_926);
xor U3667 (N_3667,N_10,N_1672);
nor U3668 (N_3668,N_720,N_108);
xor U3669 (N_3669,N_793,N_1124);
or U3670 (N_3670,N_872,N_1759);
xnor U3671 (N_3671,N_1866,N_1197);
and U3672 (N_3672,N_1074,N_236);
and U3673 (N_3673,N_143,N_795);
and U3674 (N_3674,N_588,N_28);
nand U3675 (N_3675,N_1553,N_1274);
nand U3676 (N_3676,N_1148,N_1757);
nor U3677 (N_3677,N_1409,N_543);
nand U3678 (N_3678,N_1940,N_1633);
nand U3679 (N_3679,N_1740,N_1877);
nor U3680 (N_3680,N_411,N_817);
and U3681 (N_3681,N_49,N_1442);
and U3682 (N_3682,N_811,N_1038);
or U3683 (N_3683,N_1866,N_1719);
or U3684 (N_3684,N_930,N_4);
nor U3685 (N_3685,N_843,N_707);
nor U3686 (N_3686,N_1997,N_782);
or U3687 (N_3687,N_1900,N_888);
nand U3688 (N_3688,N_660,N_1327);
nand U3689 (N_3689,N_1266,N_463);
or U3690 (N_3690,N_1928,N_671);
nand U3691 (N_3691,N_1959,N_370);
nand U3692 (N_3692,N_1642,N_1612);
nor U3693 (N_3693,N_1886,N_648);
xnor U3694 (N_3694,N_1859,N_1253);
xor U3695 (N_3695,N_1383,N_1566);
or U3696 (N_3696,N_1343,N_227);
or U3697 (N_3697,N_262,N_555);
nor U3698 (N_3698,N_1609,N_575);
or U3699 (N_3699,N_916,N_1151);
or U3700 (N_3700,N_107,N_363);
or U3701 (N_3701,N_257,N_427);
xor U3702 (N_3702,N_993,N_1108);
or U3703 (N_3703,N_537,N_807);
and U3704 (N_3704,N_1640,N_834);
nor U3705 (N_3705,N_109,N_796);
and U3706 (N_3706,N_1444,N_1163);
nor U3707 (N_3707,N_176,N_1909);
nand U3708 (N_3708,N_414,N_622);
nand U3709 (N_3709,N_383,N_507);
or U3710 (N_3710,N_303,N_720);
nand U3711 (N_3711,N_1852,N_374);
nor U3712 (N_3712,N_578,N_1032);
or U3713 (N_3713,N_1046,N_961);
nor U3714 (N_3714,N_1127,N_1446);
nor U3715 (N_3715,N_1061,N_940);
and U3716 (N_3716,N_5,N_594);
or U3717 (N_3717,N_586,N_1679);
nor U3718 (N_3718,N_879,N_1105);
and U3719 (N_3719,N_637,N_1344);
or U3720 (N_3720,N_200,N_1099);
nand U3721 (N_3721,N_177,N_280);
nor U3722 (N_3722,N_1526,N_1378);
nor U3723 (N_3723,N_327,N_66);
nand U3724 (N_3724,N_195,N_467);
nor U3725 (N_3725,N_1348,N_1514);
and U3726 (N_3726,N_1135,N_1993);
and U3727 (N_3727,N_818,N_1523);
or U3728 (N_3728,N_815,N_402);
xor U3729 (N_3729,N_1196,N_62);
or U3730 (N_3730,N_1449,N_1182);
nand U3731 (N_3731,N_1458,N_1408);
nor U3732 (N_3732,N_559,N_1775);
and U3733 (N_3733,N_327,N_531);
or U3734 (N_3734,N_219,N_526);
nand U3735 (N_3735,N_1555,N_637);
or U3736 (N_3736,N_201,N_1030);
or U3737 (N_3737,N_1096,N_1893);
nor U3738 (N_3738,N_493,N_1581);
nor U3739 (N_3739,N_278,N_49);
and U3740 (N_3740,N_9,N_599);
nand U3741 (N_3741,N_1562,N_573);
nand U3742 (N_3742,N_793,N_1262);
and U3743 (N_3743,N_1241,N_978);
and U3744 (N_3744,N_655,N_1072);
nand U3745 (N_3745,N_499,N_489);
nand U3746 (N_3746,N_1485,N_1534);
nand U3747 (N_3747,N_1215,N_841);
nand U3748 (N_3748,N_871,N_1823);
nor U3749 (N_3749,N_1742,N_1573);
nand U3750 (N_3750,N_250,N_1795);
nor U3751 (N_3751,N_1133,N_231);
and U3752 (N_3752,N_452,N_408);
nor U3753 (N_3753,N_482,N_838);
or U3754 (N_3754,N_1204,N_1100);
or U3755 (N_3755,N_980,N_1744);
nor U3756 (N_3756,N_1386,N_1785);
or U3757 (N_3757,N_71,N_530);
nor U3758 (N_3758,N_1942,N_1264);
nand U3759 (N_3759,N_653,N_1038);
and U3760 (N_3760,N_520,N_597);
and U3761 (N_3761,N_1136,N_1217);
nand U3762 (N_3762,N_1682,N_1950);
nor U3763 (N_3763,N_1311,N_21);
or U3764 (N_3764,N_420,N_1201);
nor U3765 (N_3765,N_713,N_435);
or U3766 (N_3766,N_1811,N_67);
nand U3767 (N_3767,N_774,N_549);
nor U3768 (N_3768,N_958,N_192);
nor U3769 (N_3769,N_300,N_1625);
nand U3770 (N_3770,N_648,N_967);
and U3771 (N_3771,N_608,N_769);
nand U3772 (N_3772,N_1363,N_1494);
xnor U3773 (N_3773,N_1279,N_1513);
nand U3774 (N_3774,N_1848,N_94);
or U3775 (N_3775,N_501,N_1387);
xor U3776 (N_3776,N_1858,N_1317);
nor U3777 (N_3777,N_1929,N_1309);
or U3778 (N_3778,N_378,N_838);
xor U3779 (N_3779,N_1067,N_1481);
or U3780 (N_3780,N_1000,N_1921);
nor U3781 (N_3781,N_1850,N_1040);
or U3782 (N_3782,N_260,N_792);
nand U3783 (N_3783,N_353,N_1138);
or U3784 (N_3784,N_282,N_1994);
nand U3785 (N_3785,N_700,N_1194);
or U3786 (N_3786,N_342,N_157);
nand U3787 (N_3787,N_1138,N_875);
nand U3788 (N_3788,N_866,N_12);
and U3789 (N_3789,N_339,N_912);
xnor U3790 (N_3790,N_442,N_1282);
xor U3791 (N_3791,N_1924,N_1287);
nor U3792 (N_3792,N_424,N_1476);
nor U3793 (N_3793,N_961,N_1425);
nor U3794 (N_3794,N_31,N_501);
nand U3795 (N_3795,N_174,N_733);
nor U3796 (N_3796,N_1041,N_1667);
or U3797 (N_3797,N_31,N_1786);
nand U3798 (N_3798,N_178,N_236);
or U3799 (N_3799,N_429,N_1812);
xor U3800 (N_3800,N_526,N_1314);
xnor U3801 (N_3801,N_241,N_1681);
nor U3802 (N_3802,N_338,N_343);
or U3803 (N_3803,N_550,N_1718);
nor U3804 (N_3804,N_1564,N_1263);
nor U3805 (N_3805,N_1035,N_624);
and U3806 (N_3806,N_715,N_1506);
nor U3807 (N_3807,N_1154,N_995);
and U3808 (N_3808,N_1222,N_1829);
xor U3809 (N_3809,N_1415,N_1338);
and U3810 (N_3810,N_309,N_555);
and U3811 (N_3811,N_806,N_1729);
nor U3812 (N_3812,N_1924,N_962);
nand U3813 (N_3813,N_941,N_582);
nor U3814 (N_3814,N_1592,N_762);
and U3815 (N_3815,N_1980,N_1960);
or U3816 (N_3816,N_1949,N_699);
nand U3817 (N_3817,N_1992,N_555);
and U3818 (N_3818,N_749,N_562);
and U3819 (N_3819,N_1179,N_90);
and U3820 (N_3820,N_1798,N_1300);
nand U3821 (N_3821,N_648,N_800);
or U3822 (N_3822,N_374,N_1773);
or U3823 (N_3823,N_1361,N_1864);
nor U3824 (N_3824,N_820,N_486);
or U3825 (N_3825,N_1900,N_132);
nand U3826 (N_3826,N_729,N_97);
nor U3827 (N_3827,N_1132,N_1852);
nand U3828 (N_3828,N_747,N_398);
nand U3829 (N_3829,N_1482,N_945);
and U3830 (N_3830,N_1980,N_1436);
nand U3831 (N_3831,N_179,N_1472);
xnor U3832 (N_3832,N_1204,N_120);
and U3833 (N_3833,N_1973,N_1822);
nand U3834 (N_3834,N_1002,N_1154);
nor U3835 (N_3835,N_778,N_1525);
nand U3836 (N_3836,N_1937,N_1883);
or U3837 (N_3837,N_1237,N_1950);
xor U3838 (N_3838,N_1800,N_1421);
nor U3839 (N_3839,N_1140,N_1778);
and U3840 (N_3840,N_616,N_1230);
nand U3841 (N_3841,N_1383,N_89);
nor U3842 (N_3842,N_364,N_1754);
nand U3843 (N_3843,N_1633,N_562);
nand U3844 (N_3844,N_1787,N_449);
xnor U3845 (N_3845,N_1965,N_1872);
nand U3846 (N_3846,N_1946,N_510);
nand U3847 (N_3847,N_1295,N_624);
and U3848 (N_3848,N_1649,N_770);
nor U3849 (N_3849,N_190,N_903);
nand U3850 (N_3850,N_606,N_250);
and U3851 (N_3851,N_1633,N_150);
nand U3852 (N_3852,N_945,N_1933);
nor U3853 (N_3853,N_156,N_21);
or U3854 (N_3854,N_1264,N_402);
nand U3855 (N_3855,N_1999,N_569);
nand U3856 (N_3856,N_1042,N_1615);
nand U3857 (N_3857,N_786,N_1186);
xnor U3858 (N_3858,N_588,N_543);
and U3859 (N_3859,N_1031,N_1402);
and U3860 (N_3860,N_1391,N_1164);
nor U3861 (N_3861,N_1021,N_582);
nand U3862 (N_3862,N_1651,N_1060);
and U3863 (N_3863,N_442,N_729);
or U3864 (N_3864,N_957,N_1248);
nor U3865 (N_3865,N_1641,N_267);
or U3866 (N_3866,N_1417,N_44);
nand U3867 (N_3867,N_1458,N_874);
or U3868 (N_3868,N_513,N_999);
and U3869 (N_3869,N_333,N_1236);
nand U3870 (N_3870,N_1410,N_470);
nor U3871 (N_3871,N_1387,N_1426);
or U3872 (N_3872,N_449,N_71);
xnor U3873 (N_3873,N_1207,N_34);
xor U3874 (N_3874,N_1855,N_1843);
nor U3875 (N_3875,N_513,N_1652);
or U3876 (N_3876,N_1003,N_1735);
and U3877 (N_3877,N_1701,N_894);
and U3878 (N_3878,N_1568,N_803);
or U3879 (N_3879,N_1760,N_917);
nor U3880 (N_3880,N_799,N_1614);
nand U3881 (N_3881,N_1739,N_549);
and U3882 (N_3882,N_1497,N_1887);
nor U3883 (N_3883,N_1532,N_1356);
and U3884 (N_3884,N_1301,N_647);
xnor U3885 (N_3885,N_300,N_740);
nand U3886 (N_3886,N_784,N_1549);
and U3887 (N_3887,N_304,N_1373);
nor U3888 (N_3888,N_273,N_34);
xor U3889 (N_3889,N_1973,N_1387);
nand U3890 (N_3890,N_1947,N_510);
or U3891 (N_3891,N_1154,N_328);
or U3892 (N_3892,N_43,N_227);
and U3893 (N_3893,N_1855,N_962);
or U3894 (N_3894,N_1943,N_1010);
and U3895 (N_3895,N_1047,N_596);
nor U3896 (N_3896,N_1714,N_547);
nand U3897 (N_3897,N_1725,N_1908);
nand U3898 (N_3898,N_719,N_1789);
nand U3899 (N_3899,N_723,N_1647);
and U3900 (N_3900,N_1045,N_838);
and U3901 (N_3901,N_1333,N_1603);
xor U3902 (N_3902,N_1196,N_1061);
xor U3903 (N_3903,N_1821,N_220);
nand U3904 (N_3904,N_574,N_482);
and U3905 (N_3905,N_441,N_636);
and U3906 (N_3906,N_818,N_1960);
nand U3907 (N_3907,N_1563,N_1081);
and U3908 (N_3908,N_431,N_1044);
and U3909 (N_3909,N_1927,N_107);
nor U3910 (N_3910,N_37,N_570);
nor U3911 (N_3911,N_1866,N_1814);
or U3912 (N_3912,N_1720,N_1410);
and U3913 (N_3913,N_78,N_1018);
nor U3914 (N_3914,N_1880,N_1546);
nor U3915 (N_3915,N_1327,N_578);
or U3916 (N_3916,N_464,N_729);
xnor U3917 (N_3917,N_1094,N_1035);
nor U3918 (N_3918,N_1522,N_1469);
or U3919 (N_3919,N_1303,N_1148);
and U3920 (N_3920,N_1837,N_1140);
or U3921 (N_3921,N_1696,N_851);
nand U3922 (N_3922,N_1370,N_44);
nor U3923 (N_3923,N_1092,N_902);
nand U3924 (N_3924,N_779,N_1640);
nor U3925 (N_3925,N_1473,N_606);
nand U3926 (N_3926,N_1662,N_720);
nand U3927 (N_3927,N_1345,N_280);
or U3928 (N_3928,N_312,N_328);
and U3929 (N_3929,N_125,N_258);
or U3930 (N_3930,N_1083,N_288);
nor U3931 (N_3931,N_1442,N_1931);
nor U3932 (N_3932,N_1793,N_1555);
or U3933 (N_3933,N_1225,N_1658);
nand U3934 (N_3934,N_1639,N_472);
and U3935 (N_3935,N_874,N_1510);
and U3936 (N_3936,N_1625,N_1998);
and U3937 (N_3937,N_30,N_726);
nand U3938 (N_3938,N_1434,N_1413);
and U3939 (N_3939,N_898,N_1908);
nor U3940 (N_3940,N_581,N_1918);
or U3941 (N_3941,N_791,N_721);
xnor U3942 (N_3942,N_195,N_88);
or U3943 (N_3943,N_936,N_1235);
or U3944 (N_3944,N_757,N_1064);
nand U3945 (N_3945,N_942,N_1835);
and U3946 (N_3946,N_1094,N_61);
nand U3947 (N_3947,N_689,N_1412);
nand U3948 (N_3948,N_336,N_90);
nor U3949 (N_3949,N_1607,N_1754);
nor U3950 (N_3950,N_1853,N_1344);
xor U3951 (N_3951,N_402,N_537);
nand U3952 (N_3952,N_34,N_1481);
and U3953 (N_3953,N_653,N_1816);
and U3954 (N_3954,N_1205,N_912);
nor U3955 (N_3955,N_786,N_960);
and U3956 (N_3956,N_1279,N_542);
or U3957 (N_3957,N_246,N_1376);
nand U3958 (N_3958,N_1330,N_1051);
xnor U3959 (N_3959,N_1768,N_162);
and U3960 (N_3960,N_1466,N_1093);
nor U3961 (N_3961,N_478,N_611);
nor U3962 (N_3962,N_1535,N_1496);
and U3963 (N_3963,N_980,N_353);
or U3964 (N_3964,N_644,N_926);
and U3965 (N_3965,N_240,N_1749);
or U3966 (N_3966,N_1872,N_1047);
and U3967 (N_3967,N_2,N_788);
xor U3968 (N_3968,N_1238,N_266);
xor U3969 (N_3969,N_1000,N_1349);
nor U3970 (N_3970,N_1252,N_993);
and U3971 (N_3971,N_82,N_1058);
and U3972 (N_3972,N_1499,N_1563);
or U3973 (N_3973,N_1583,N_1386);
and U3974 (N_3974,N_1616,N_770);
and U3975 (N_3975,N_459,N_411);
nand U3976 (N_3976,N_498,N_1953);
or U3977 (N_3977,N_65,N_412);
or U3978 (N_3978,N_588,N_834);
or U3979 (N_3979,N_1644,N_552);
nor U3980 (N_3980,N_1220,N_1908);
xnor U3981 (N_3981,N_585,N_1882);
nand U3982 (N_3982,N_1412,N_750);
nand U3983 (N_3983,N_1518,N_362);
nand U3984 (N_3984,N_127,N_1480);
and U3985 (N_3985,N_845,N_718);
and U3986 (N_3986,N_1044,N_68);
nor U3987 (N_3987,N_1400,N_829);
or U3988 (N_3988,N_75,N_1756);
nor U3989 (N_3989,N_743,N_1532);
or U3990 (N_3990,N_910,N_936);
nor U3991 (N_3991,N_1238,N_823);
nor U3992 (N_3992,N_220,N_399);
xnor U3993 (N_3993,N_783,N_1152);
nand U3994 (N_3994,N_1510,N_475);
and U3995 (N_3995,N_1945,N_1445);
nor U3996 (N_3996,N_50,N_1876);
nor U3997 (N_3997,N_1043,N_1601);
and U3998 (N_3998,N_1103,N_880);
or U3999 (N_3999,N_195,N_588);
nor U4000 (N_4000,N_2673,N_3938);
and U4001 (N_4001,N_3270,N_3563);
nand U4002 (N_4002,N_2834,N_2622);
nand U4003 (N_4003,N_2844,N_2062);
nand U4004 (N_4004,N_2193,N_2083);
nor U4005 (N_4005,N_3792,N_3004);
nor U4006 (N_4006,N_2442,N_2361);
or U4007 (N_4007,N_2082,N_2323);
nor U4008 (N_4008,N_2359,N_3067);
and U4009 (N_4009,N_3000,N_2146);
nand U4010 (N_4010,N_2043,N_2642);
and U4011 (N_4011,N_3888,N_2240);
or U4012 (N_4012,N_2746,N_3984);
xnor U4013 (N_4013,N_3690,N_2572);
and U4014 (N_4014,N_2813,N_3552);
nand U4015 (N_4015,N_2392,N_2461);
nor U4016 (N_4016,N_3358,N_3264);
nor U4017 (N_4017,N_2898,N_3853);
and U4018 (N_4018,N_3080,N_2071);
nor U4019 (N_4019,N_3583,N_3720);
and U4020 (N_4020,N_3254,N_2923);
or U4021 (N_4021,N_3497,N_3472);
nand U4022 (N_4022,N_3926,N_2244);
nand U4023 (N_4023,N_3279,N_3842);
and U4024 (N_4024,N_3307,N_2591);
and U4025 (N_4025,N_3907,N_2942);
nand U4026 (N_4026,N_3285,N_3900);
nand U4027 (N_4027,N_3483,N_2383);
and U4028 (N_4028,N_3560,N_2829);
nor U4029 (N_4029,N_3868,N_3796);
or U4030 (N_4030,N_2706,N_3007);
nand U4031 (N_4031,N_2034,N_2724);
and U4032 (N_4032,N_2238,N_3337);
or U4033 (N_4033,N_3241,N_2830);
or U4034 (N_4034,N_2200,N_2938);
nor U4035 (N_4035,N_3089,N_2725);
and U4036 (N_4036,N_2550,N_3245);
or U4037 (N_4037,N_3533,N_2876);
nand U4038 (N_4038,N_2395,N_2935);
or U4039 (N_4039,N_2079,N_3315);
or U4040 (N_4040,N_2552,N_3079);
nor U4041 (N_4041,N_2266,N_3460);
and U4042 (N_4042,N_3828,N_3542);
and U4043 (N_4043,N_3649,N_3357);
xnor U4044 (N_4044,N_3503,N_2901);
nor U4045 (N_4045,N_3744,N_2566);
xor U4046 (N_4046,N_3424,N_2772);
xor U4047 (N_4047,N_2320,N_3210);
and U4048 (N_4048,N_3688,N_2979);
or U4049 (N_4049,N_2421,N_2908);
nand U4050 (N_4050,N_2149,N_3887);
xnor U4051 (N_4051,N_2311,N_2729);
or U4052 (N_4052,N_3031,N_2096);
or U4053 (N_4053,N_3819,N_2865);
nand U4054 (N_4054,N_2807,N_2986);
or U4055 (N_4055,N_2771,N_2191);
or U4056 (N_4056,N_3738,N_2815);
or U4057 (N_4057,N_3145,N_3893);
and U4058 (N_4058,N_3641,N_3223);
or U4059 (N_4059,N_2267,N_3468);
or U4060 (N_4060,N_2039,N_2620);
nor U4061 (N_4061,N_2067,N_2786);
or U4062 (N_4062,N_3675,N_2855);
or U4063 (N_4063,N_2489,N_2093);
and U4064 (N_4064,N_2188,N_2895);
nor U4065 (N_4065,N_2674,N_2055);
nand U4066 (N_4066,N_3843,N_2549);
nor U4067 (N_4067,N_2580,N_2977);
and U4068 (N_4068,N_2298,N_3695);
or U4069 (N_4069,N_3822,N_2070);
or U4070 (N_4070,N_3184,N_3767);
nand U4071 (N_4071,N_2946,N_2514);
nor U4072 (N_4072,N_3415,N_2627);
or U4073 (N_4073,N_3502,N_3345);
or U4074 (N_4074,N_2475,N_2181);
nand U4075 (N_4075,N_2235,N_3491);
and U4076 (N_4076,N_2886,N_2808);
or U4077 (N_4077,N_3433,N_2177);
or U4078 (N_4078,N_2542,N_2709);
nor U4079 (N_4079,N_2215,N_3188);
nand U4080 (N_4080,N_2887,N_2218);
and U4081 (N_4081,N_2948,N_2293);
xor U4082 (N_4082,N_3495,N_2018);
nand U4083 (N_4083,N_2125,N_2049);
nand U4084 (N_4084,N_2516,N_3258);
nor U4085 (N_4085,N_2372,N_3230);
nand U4086 (N_4086,N_3289,N_3655);
or U4087 (N_4087,N_2905,N_2890);
or U4088 (N_4088,N_3643,N_3795);
nor U4089 (N_4089,N_3911,N_2641);
nand U4090 (N_4090,N_2152,N_3021);
and U4091 (N_4091,N_2233,N_3086);
nor U4092 (N_4092,N_2732,N_3523);
and U4093 (N_4093,N_3557,N_3074);
and U4094 (N_4094,N_2755,N_3359);
or U4095 (N_4095,N_2336,N_3136);
nor U4096 (N_4096,N_2026,N_2332);
nand U4097 (N_4097,N_3319,N_3908);
or U4098 (N_4098,N_3311,N_3799);
nor U4099 (N_4099,N_2427,N_2458);
xor U4100 (N_4100,N_3801,N_2992);
nor U4101 (N_4101,N_3905,N_2775);
nor U4102 (N_4102,N_3158,N_2749);
or U4103 (N_4103,N_3239,N_2434);
and U4104 (N_4104,N_3252,N_2646);
or U4105 (N_4105,N_3480,N_3628);
and U4106 (N_4106,N_2403,N_2751);
nor U4107 (N_4107,N_3185,N_2249);
or U4108 (N_4108,N_2230,N_2636);
or U4109 (N_4109,N_2241,N_3212);
and U4110 (N_4110,N_2389,N_2608);
nand U4111 (N_4111,N_2217,N_3963);
xor U4112 (N_4112,N_2902,N_2020);
nor U4113 (N_4113,N_2237,N_2957);
nor U4114 (N_4114,N_3193,N_3127);
nor U4115 (N_4115,N_3394,N_3321);
nand U4116 (N_4116,N_2577,N_2394);
nor U4117 (N_4117,N_2573,N_2987);
nand U4118 (N_4118,N_3789,N_2816);
nor U4119 (N_4119,N_3006,N_3214);
nor U4120 (N_4120,N_2207,N_2927);
nand U4121 (N_4121,N_2285,N_2019);
nor U4122 (N_4122,N_3618,N_2998);
and U4123 (N_4123,N_3488,N_2765);
and U4124 (N_4124,N_3626,N_2214);
xnor U4125 (N_4125,N_3847,N_3861);
or U4126 (N_4126,N_3949,N_3869);
nand U4127 (N_4127,N_2360,N_2316);
nor U4128 (N_4128,N_3120,N_2046);
or U4129 (N_4129,N_2909,N_2907);
nor U4130 (N_4130,N_2113,N_3066);
or U4131 (N_4131,N_3175,N_3780);
nor U4132 (N_4132,N_3035,N_2970);
nand U4133 (N_4133,N_3482,N_3050);
nor U4134 (N_4134,N_3501,N_3186);
or U4135 (N_4135,N_3419,N_3904);
nor U4136 (N_4136,N_3437,N_3440);
nor U4137 (N_4137,N_2199,N_2187);
nand U4138 (N_4138,N_2462,N_3397);
and U4139 (N_4139,N_2420,N_2006);
and U4140 (N_4140,N_2645,N_3221);
nor U4141 (N_4141,N_2415,N_2994);
or U4142 (N_4142,N_2715,N_2474);
or U4143 (N_4143,N_2969,N_2952);
or U4144 (N_4144,N_3978,N_3678);
nand U4145 (N_4145,N_2799,N_2033);
or U4146 (N_4146,N_3585,N_3640);
and U4147 (N_4147,N_3972,N_2499);
nand U4148 (N_4148,N_2762,N_2433);
and U4149 (N_4149,N_2903,N_3263);
and U4150 (N_4150,N_3469,N_3739);
nand U4151 (N_4151,N_3920,N_3566);
and U4152 (N_4152,N_3444,N_3361);
or U4153 (N_4153,N_3377,N_3676);
or U4154 (N_4154,N_3934,N_2115);
or U4155 (N_4155,N_3055,N_3854);
or U4156 (N_4156,N_3764,N_3191);
or U4157 (N_4157,N_2047,N_2364);
nand U4158 (N_4158,N_3148,N_2091);
xnor U4159 (N_4159,N_3290,N_2600);
nand U4160 (N_4160,N_2576,N_2617);
nor U4161 (N_4161,N_3748,N_3840);
or U4162 (N_4162,N_3753,N_2839);
nand U4163 (N_4163,N_3068,N_3862);
nor U4164 (N_4164,N_2124,N_2208);
xor U4165 (N_4165,N_2041,N_2077);
nand U4166 (N_4166,N_2086,N_2468);
nand U4167 (N_4167,N_2509,N_2679);
nand U4168 (N_4168,N_3492,N_2716);
xnor U4169 (N_4169,N_2411,N_2105);
nor U4170 (N_4170,N_3332,N_3395);
nor U4171 (N_4171,N_3236,N_2512);
and U4172 (N_4172,N_2660,N_3546);
nand U4173 (N_4173,N_2268,N_3613);
or U4174 (N_4174,N_3831,N_2692);
and U4175 (N_4175,N_2060,N_2261);
xor U4176 (N_4176,N_3825,N_2104);
or U4177 (N_4177,N_2707,N_2401);
nor U4178 (N_4178,N_3126,N_3692);
nand U4179 (N_4179,N_2423,N_3844);
nand U4180 (N_4180,N_2974,N_3088);
or U4181 (N_4181,N_3924,N_2459);
and U4182 (N_4182,N_2581,N_3138);
nand U4183 (N_4183,N_2232,N_2934);
or U4184 (N_4184,N_3986,N_2156);
nand U4185 (N_4185,N_2085,N_2900);
xnor U4186 (N_4186,N_3671,N_2335);
nand U4187 (N_4187,N_2805,N_2963);
or U4188 (N_4188,N_2857,N_3448);
nor U4189 (N_4189,N_2988,N_3165);
or U4190 (N_4190,N_2697,N_2072);
nor U4191 (N_4191,N_3180,N_2426);
xnor U4192 (N_4192,N_3561,N_3500);
or U4193 (N_4193,N_3063,N_3071);
nor U4194 (N_4194,N_3346,N_2226);
or U4195 (N_4195,N_2625,N_3473);
or U4196 (N_4196,N_3755,N_2297);
nor U4197 (N_4197,N_2453,N_3586);
nand U4198 (N_4198,N_2176,N_2483);
nand U4199 (N_4199,N_3256,N_2363);
nand U4200 (N_4200,N_2947,N_3855);
xor U4201 (N_4201,N_3711,N_3867);
or U4202 (N_4202,N_3942,N_2075);
nand U4203 (N_4203,N_2711,N_2161);
nand U4204 (N_4204,N_2467,N_2092);
or U4205 (N_4205,N_3336,N_2384);
nand U4206 (N_4206,N_3324,N_2779);
nand U4207 (N_4207,N_3879,N_3749);
nand U4208 (N_4208,N_2720,N_2357);
xor U4209 (N_4209,N_3016,N_3570);
xor U4210 (N_4210,N_2430,N_3807);
and U4211 (N_4211,N_2398,N_3135);
xnor U4212 (N_4212,N_3830,N_2252);
nor U4213 (N_4213,N_2614,N_2893);
and U4214 (N_4214,N_2140,N_2410);
nor U4215 (N_4215,N_3567,N_2400);
or U4216 (N_4216,N_3093,N_3343);
xor U4217 (N_4217,N_3642,N_3334);
or U4218 (N_4218,N_2350,N_3808);
nor U4219 (N_4219,N_3190,N_3846);
nand U4220 (N_4220,N_2980,N_3446);
or U4221 (N_4221,N_2570,N_3562);
or U4222 (N_4222,N_3342,N_2823);
nor U4223 (N_4223,N_3330,N_3697);
nand U4224 (N_4224,N_3967,N_3030);
nand U4225 (N_4225,N_3875,N_3723);
or U4226 (N_4226,N_2160,N_2319);
or U4227 (N_4227,N_3454,N_3709);
or U4228 (N_4228,N_3237,N_2011);
nor U4229 (N_4229,N_2012,N_3824);
or U4230 (N_4230,N_2469,N_2277);
and U4231 (N_4231,N_3891,N_2223);
or U4232 (N_4232,N_2874,N_2151);
or U4233 (N_4233,N_2741,N_2279);
and U4234 (N_4234,N_3047,N_2849);
or U4235 (N_4235,N_3681,N_3961);
xnor U4236 (N_4236,N_3860,N_3203);
or U4237 (N_4237,N_3464,N_3215);
nor U4238 (N_4238,N_3043,N_2528);
nor U4239 (N_4239,N_3968,N_2730);
or U4240 (N_4240,N_2127,N_3354);
and U4241 (N_4241,N_3710,N_2953);
nand U4242 (N_4242,N_3880,N_2449);
xor U4243 (N_4243,N_3405,N_2429);
nand U4244 (N_4244,N_3020,N_3945);
nand U4245 (N_4245,N_3970,N_3196);
and U4246 (N_4246,N_2144,N_3033);
or U4247 (N_4247,N_2317,N_3216);
or U4248 (N_4248,N_2183,N_3933);
xor U4249 (N_4249,N_3130,N_3353);
and U4250 (N_4250,N_2851,N_3046);
nor U4251 (N_4251,N_2048,N_3244);
nor U4252 (N_4252,N_2287,N_2435);
nand U4253 (N_4253,N_2776,N_3247);
nand U4254 (N_4254,N_3775,N_3573);
nand U4255 (N_4255,N_2037,N_2780);
and U4256 (N_4256,N_2413,N_3356);
nand U4257 (N_4257,N_3917,N_2123);
or U4258 (N_4258,N_3721,N_3713);
nand U4259 (N_4259,N_2295,N_2676);
and U4260 (N_4260,N_3699,N_3457);
nor U4261 (N_4261,N_3943,N_3877);
nand U4262 (N_4262,N_2508,N_2662);
or U4263 (N_4263,N_2141,N_3788);
nand U4264 (N_4264,N_2533,N_2283);
or U4265 (N_4265,N_2002,N_2655);
nand U4266 (N_4266,N_3049,N_2321);
nor U4267 (N_4267,N_2536,N_3105);
or U4268 (N_4268,N_2278,N_2866);
nand U4269 (N_4269,N_2584,N_3073);
nor U4270 (N_4270,N_3725,N_2425);
nand U4271 (N_4271,N_2112,N_2366);
and U4272 (N_4272,N_2349,N_2594);
or U4273 (N_4273,N_2993,N_2589);
nand U4274 (N_4274,N_3112,N_2373);
and U4275 (N_4275,N_3429,N_2723);
nor U4276 (N_4276,N_2678,N_3117);
nand U4277 (N_4277,N_3179,N_2685);
xnor U4278 (N_4278,N_2066,N_2675);
and U4279 (N_4279,N_2431,N_3296);
nand U4280 (N_4280,N_2888,N_2030);
nor U4281 (N_4281,N_3009,N_2510);
xnor U4282 (N_4282,N_2009,N_3392);
nand U4283 (N_4283,N_2719,N_2159);
nor U4284 (N_4284,N_3134,N_2473);
nor U4285 (N_4285,N_3144,N_3601);
nor U4286 (N_4286,N_3224,N_3227);
xnor U4287 (N_4287,N_2001,N_2978);
nand U4288 (N_4288,N_3981,N_2480);
and U4289 (N_4289,N_2440,N_3450);
or U4290 (N_4290,N_3376,N_2562);
or U4291 (N_4291,N_3008,N_2209);
and U4292 (N_4292,N_2007,N_2472);
nand U4293 (N_4293,N_2748,N_3839);
nand U4294 (N_4294,N_3040,N_3584);
nand U4295 (N_4295,N_2212,N_3019);
nor U4296 (N_4296,N_3017,N_3368);
xor U4297 (N_4297,N_3889,N_2554);
nor U4298 (N_4298,N_2479,N_3052);
nand U4299 (N_4299,N_2683,N_3520);
xnor U4300 (N_4300,N_2455,N_3139);
or U4301 (N_4301,N_2116,N_3261);
and U4302 (N_4302,N_3260,N_3275);
or U4303 (N_4303,N_2882,N_3703);
or U4304 (N_4304,N_3110,N_2052);
and U4305 (N_4305,N_3374,N_3565);
and U4306 (N_4306,N_3335,N_2179);
or U4307 (N_4307,N_3229,N_2061);
xnor U4308 (N_4308,N_2471,N_3619);
and U4309 (N_4309,N_2281,N_2170);
nand U4310 (N_4310,N_2586,N_2595);
xor U4311 (N_4311,N_3282,N_3650);
and U4312 (N_4312,N_3892,N_3527);
or U4313 (N_4313,N_2537,N_3832);
or U4314 (N_4314,N_2497,N_2407);
or U4315 (N_4315,N_2688,N_3208);
and U4316 (N_4316,N_2728,N_2899);
nand U4317 (N_4317,N_3129,N_2733);
or U4318 (N_4318,N_3577,N_3028);
or U4319 (N_4319,N_2255,N_3137);
nor U4320 (N_4320,N_3508,N_2211);
and U4321 (N_4321,N_3351,N_2657);
nand U4322 (N_4322,N_3271,N_2910);
nand U4323 (N_4323,N_2204,N_3418);
or U4324 (N_4324,N_2968,N_3559);
and U4325 (N_4325,N_2122,N_3779);
or U4326 (N_4326,N_3059,N_2131);
nor U4327 (N_4327,N_3550,N_2257);
nand U4328 (N_4328,N_3689,N_2387);
nand U4329 (N_4329,N_3802,N_2153);
nor U4330 (N_4330,N_2515,N_3940);
nor U4331 (N_4331,N_2326,N_2973);
nand U4332 (N_4332,N_2520,N_2290);
nand U4333 (N_4333,N_2504,N_3316);
xor U4334 (N_4334,N_2492,N_3107);
nand U4335 (N_4335,N_2376,N_3806);
nor U4336 (N_4336,N_3011,N_3598);
nand U4337 (N_4337,N_3202,N_3528);
nand U4338 (N_4338,N_2758,N_2526);
and U4339 (N_4339,N_2681,N_2135);
and U4340 (N_4340,N_2792,N_3811);
or U4341 (N_4341,N_3916,N_3848);
and U4342 (N_4342,N_2169,N_2243);
nor U4343 (N_4343,N_3250,N_3896);
nor U4344 (N_4344,N_2721,N_3338);
and U4345 (N_4345,N_3147,N_2548);
nor U4346 (N_4346,N_2864,N_3034);
nand U4347 (N_4347,N_2932,N_3672);
and U4348 (N_4348,N_3538,N_2643);
nor U4349 (N_4349,N_3360,N_3515);
and U4350 (N_4350,N_2590,N_3280);
or U4351 (N_4351,N_3143,N_3679);
and U4352 (N_4352,N_3114,N_3918);
and U4353 (N_4353,N_3461,N_3155);
nor U4354 (N_4354,N_3576,N_2754);
xnor U4355 (N_4355,N_3750,N_2056);
and U4356 (N_4356,N_3101,N_2097);
nor U4357 (N_4357,N_2598,N_3646);
nand U4358 (N_4358,N_2975,N_3727);
and U4359 (N_4359,N_2929,N_2791);
nand U4360 (N_4360,N_2774,N_2111);
nand U4361 (N_4361,N_3425,N_2972);
xor U4362 (N_4362,N_2155,N_2736);
nor U4363 (N_4363,N_2951,N_3947);
and U4364 (N_4364,N_3232,N_2546);
nor U4365 (N_4365,N_2309,N_3973);
nand U4366 (N_4366,N_3836,N_3732);
xor U4367 (N_4367,N_2377,N_2846);
xnor U4368 (N_4368,N_2023,N_2302);
nor U4369 (N_4369,N_3841,N_2119);
or U4370 (N_4370,N_3962,N_3288);
nor U4371 (N_4371,N_2369,N_2228);
and U4372 (N_4372,N_3677,N_3187);
nor U4373 (N_4373,N_2853,N_3680);
nand U4374 (N_4374,N_2303,N_3730);
nand U4375 (N_4375,N_2305,N_3434);
or U4376 (N_4376,N_2275,N_3674);
or U4377 (N_4377,N_2069,N_2880);
nor U4378 (N_4378,N_3410,N_3507);
nor U4379 (N_4379,N_2166,N_3170);
and U4380 (N_4380,N_2253,N_2700);
nor U4381 (N_4381,N_2206,N_3589);
and U4382 (N_4382,N_3371,N_2753);
nor U4383 (N_4383,N_2647,N_3421);
and U4384 (N_4384,N_3234,N_3382);
nor U4385 (N_4385,N_2102,N_3005);
or U4386 (N_4386,N_2618,N_3463);
or U4387 (N_4387,N_3015,N_2213);
or U4388 (N_4388,N_2565,N_2470);
or U4389 (N_4389,N_2322,N_2405);
xor U4390 (N_4390,N_2227,N_2971);
or U4391 (N_4391,N_2539,N_2606);
nand U4392 (N_4392,N_3192,N_3724);
and U4393 (N_4393,N_2856,N_3818);
xor U4394 (N_4394,N_2448,N_3517);
nor U4395 (N_4395,N_2517,N_3754);
xor U4396 (N_4396,N_2623,N_2068);
or U4397 (N_4397,N_2958,N_3793);
and U4398 (N_4398,N_3763,N_2802);
nand U4399 (N_4399,N_3535,N_3594);
nand U4400 (N_4400,N_2250,N_2010);
or U4401 (N_4401,N_3274,N_2763);
xnor U4402 (N_4402,N_3298,N_2718);
and U4403 (N_4403,N_3662,N_3514);
or U4404 (N_4404,N_2672,N_3606);
nand U4405 (N_4405,N_2547,N_3458);
or U4406 (N_4406,N_3639,N_3572);
nor U4407 (N_4407,N_3142,N_2693);
nor U4408 (N_4408,N_3693,N_3845);
nor U4409 (N_4409,N_3791,N_3310);
nand U4410 (N_4410,N_3803,N_3849);
or U4411 (N_4411,N_2928,N_3901);
and U4412 (N_4412,N_2234,N_2342);
nor U4413 (N_4413,N_2652,N_2095);
and U4414 (N_4414,N_2976,N_3122);
or U4415 (N_4415,N_3442,N_2045);
and U4416 (N_4416,N_3785,N_2502);
nor U4417 (N_4417,N_3574,N_3156);
and U4418 (N_4418,N_2684,N_3992);
nor U4419 (N_4419,N_3631,N_3554);
nand U4420 (N_4420,N_2878,N_3997);
and U4421 (N_4421,N_2158,N_3431);
nand U4422 (N_4422,N_3519,N_2478);
or U4423 (N_4423,N_2996,N_2629);
and U4424 (N_4424,N_2417,N_2698);
and U4425 (N_4425,N_2621,N_2966);
and U4426 (N_4426,N_3183,N_2128);
nor U4427 (N_4427,N_2640,N_2631);
or U4428 (N_4428,N_2883,N_3391);
nand U4429 (N_4429,N_3199,N_2983);
or U4430 (N_4430,N_3581,N_2852);
and U4431 (N_4431,N_3506,N_3441);
or U4432 (N_4432,N_3609,N_3131);
xnor U4433 (N_4433,N_3612,N_3665);
and U4434 (N_4434,N_2087,N_3102);
nor U4435 (N_4435,N_2059,N_3115);
and U4436 (N_4436,N_3633,N_2954);
or U4437 (N_4437,N_2867,N_2490);
nand U4438 (N_4438,N_3540,N_2186);
nand U4439 (N_4439,N_3766,N_3453);
or U4440 (N_4440,N_3349,N_2889);
nor U4441 (N_4441,N_3160,N_3683);
and U4442 (N_4442,N_2619,N_3477);
nor U4443 (N_4443,N_2103,N_3883);
and U4444 (N_4444,N_3702,N_2906);
or U4445 (N_4445,N_3995,N_2378);
and U4446 (N_4446,N_2612,N_3784);
nand U4447 (N_4447,N_3691,N_3976);
and U4448 (N_4448,N_2269,N_2670);
or U4449 (N_4449,N_3365,N_3804);
and U4450 (N_4450,N_2569,N_2875);
xnor U4451 (N_4451,N_2789,N_3176);
nor U4452 (N_4452,N_3707,N_2588);
xor U4453 (N_4453,N_3012,N_3608);
nand U4454 (N_4454,N_3189,N_3985);
or U4455 (N_4455,N_2262,N_3948);
nand U4456 (N_4456,N_3061,N_3859);
nor U4457 (N_4457,N_2477,N_2167);
nor U4458 (N_4458,N_2328,N_2860);
nor U4459 (N_4459,N_3718,N_2424);
nor U4460 (N_4460,N_3659,N_3714);
and U4461 (N_4461,N_2696,N_3060);
and U4462 (N_4462,N_3588,N_3816);
nand U4463 (N_4463,N_2739,N_3914);
xor U4464 (N_4464,N_3094,N_3308);
xor U4465 (N_4465,N_3874,N_3657);
nand U4466 (N_4466,N_2216,N_2922);
nor U4467 (N_4467,N_2560,N_3253);
and U4468 (N_4468,N_3910,N_3163);
and U4469 (N_4469,N_3872,N_3977);
nor U4470 (N_4470,N_2282,N_3380);
and U4471 (N_4471,N_2375,N_2745);
nor U4472 (N_4472,N_2837,N_3002);
nand U4473 (N_4473,N_2343,N_3745);
and U4474 (N_4474,N_3291,N_2961);
or U4475 (N_4475,N_2985,N_3476);
nand U4476 (N_4476,N_2251,N_3706);
nor U4477 (N_4477,N_2759,N_3790);
or U4478 (N_4478,N_2769,N_3760);
nand U4479 (N_4479,N_2120,N_3529);
and U4480 (N_4480,N_3870,N_3304);
or U4481 (N_4481,N_2171,N_2933);
nor U4482 (N_4482,N_3420,N_3571);
nand U4483 (N_4483,N_2339,N_2106);
nor U4484 (N_4484,N_2511,N_3827);
nand U4485 (N_4485,N_3003,N_3599);
or U4486 (N_4486,N_2936,N_2556);
or U4487 (N_4487,N_3341,N_3098);
xnor U4488 (N_4488,N_2638,N_3352);
nor U4489 (N_4489,N_3965,N_3704);
nand U4490 (N_4490,N_2659,N_2991);
or U4491 (N_4491,N_2944,N_2025);
nand U4492 (N_4492,N_2630,N_3301);
nor U4493 (N_4493,N_3851,N_3373);
and U4494 (N_4494,N_3462,N_3820);
nor U4495 (N_4495,N_2585,N_3240);
nand U4496 (N_4496,N_2545,N_3580);
nor U4497 (N_4497,N_2794,N_3980);
and U4498 (N_4498,N_2165,N_3235);
or U4499 (N_4499,N_3556,N_2286);
or U4500 (N_4500,N_3758,N_3095);
and U4501 (N_4501,N_2017,N_2635);
or U4502 (N_4502,N_2873,N_3379);
or U4503 (N_4503,N_3076,N_2826);
and U4504 (N_4504,N_3927,N_3960);
nor U4505 (N_4505,N_2368,N_3666);
xnor U4506 (N_4506,N_2337,N_3975);
nor U4507 (N_4507,N_2354,N_2132);
or U4508 (N_4508,N_3438,N_2661);
nor U4509 (N_4509,N_3414,N_2254);
nand U4510 (N_4510,N_2098,N_2414);
nand U4511 (N_4511,N_3484,N_2452);
nand U4512 (N_4512,N_2174,N_2422);
or U4513 (N_4513,N_2381,N_2203);
nor U4514 (N_4514,N_2854,N_2727);
nor U4515 (N_4515,N_3591,N_2456);
or U4516 (N_4516,N_2788,N_2157);
and U4517 (N_4517,N_3057,N_2245);
nor U4518 (N_4518,N_3164,N_2327);
xnor U4519 (N_4519,N_2574,N_3181);
and U4520 (N_4520,N_2710,N_3177);
nor U4521 (N_4521,N_2787,N_2582);
nand U4522 (N_4522,N_2032,N_3884);
or U4523 (N_4523,N_3166,N_3375);
nor U4524 (N_4524,N_3347,N_3326);
nand U4525 (N_4525,N_2821,N_2564);
or U4526 (N_4526,N_2583,N_2783);
and U4527 (N_4527,N_2668,N_2500);
and U4528 (N_4528,N_3249,N_2221);
nand U4529 (N_4529,N_3182,N_3146);
nand U4530 (N_4530,N_3637,N_2760);
or U4531 (N_4531,N_3838,N_3762);
xor U4532 (N_4532,N_3099,N_3548);
or U4533 (N_4533,N_2879,N_3422);
or U4534 (N_4534,N_2699,N_3238);
and U4535 (N_4535,N_3297,N_2129);
nand U4536 (N_4536,N_3387,N_2943);
and U4537 (N_4537,N_3850,N_2438);
nor U4538 (N_4538,N_2142,N_2040);
or U4539 (N_4539,N_2063,N_2201);
nor U4540 (N_4540,N_2248,N_3834);
and U4541 (N_4541,N_3823,N_3814);
nand U4542 (N_4542,N_2133,N_3154);
nand U4543 (N_4543,N_3416,N_3964);
and U4544 (N_4544,N_2735,N_3773);
nand U4545 (N_4545,N_2107,N_2027);
nand U4546 (N_4546,N_2990,N_2604);
xnor U4547 (N_4547,N_3037,N_2371);
and U4548 (N_4548,N_3969,N_3881);
nor U4549 (N_4549,N_2108,N_2524);
or U4550 (N_4550,N_3794,N_3829);
nand U4551 (N_4551,N_3096,N_3409);
and U4552 (N_4552,N_2385,N_2355);
or U4553 (N_4553,N_3417,N_3797);
or U4554 (N_4554,N_2386,N_2825);
nor U4555 (N_4555,N_2145,N_2460);
and U4556 (N_4556,N_2189,N_2173);
nand U4557 (N_4557,N_2352,N_3530);
or U4558 (N_4558,N_3620,N_3010);
or U4559 (N_4559,N_3592,N_3698);
nand U4560 (N_4560,N_3747,N_2778);
nor U4561 (N_4561,N_2518,N_2481);
nor U4562 (N_4562,N_2818,N_2114);
xor U4563 (N_4563,N_2353,N_2258);
xor U4564 (N_4564,N_2088,N_2225);
nand U4565 (N_4565,N_2379,N_2797);
and U4566 (N_4566,N_2054,N_2703);
xor U4567 (N_4567,N_2348,N_3075);
xor U4568 (N_4568,N_2781,N_2965);
nor U4569 (N_4569,N_2304,N_3284);
or U4570 (N_4570,N_3157,N_3197);
nand U4571 (N_4571,N_3490,N_3663);
nor U4572 (N_4572,N_3299,N_2862);
and U4573 (N_4573,N_3622,N_3056);
xor U4574 (N_4574,N_3344,N_3950);
xor U4575 (N_4575,N_2832,N_2651);
and U4576 (N_4576,N_2219,N_3553);
and U4577 (N_4577,N_2796,N_2742);
and U4578 (N_4578,N_3231,N_3092);
or U4579 (N_4579,N_3498,N_3087);
nand U4580 (N_4580,N_3396,N_3604);
nand U4581 (N_4581,N_3809,N_2761);
and U4582 (N_4582,N_3988,N_3314);
xor U4583 (N_4583,N_2205,N_2222);
nor U4584 (N_4584,N_3487,N_2911);
nand U4585 (N_4585,N_2744,N_3257);
or U4586 (N_4586,N_2418,N_3505);
or U4587 (N_4587,N_3638,N_2168);
and U4588 (N_4588,N_2447,N_3894);
xor U4589 (N_4589,N_2446,N_2809);
and U4590 (N_4590,N_3778,N_3812);
nor U4591 (N_4591,N_2004,N_2464);
and U4592 (N_4592,N_3267,N_2344);
or U4593 (N_4593,N_3798,N_3813);
nor U4594 (N_4594,N_2610,N_2308);
nor U4595 (N_4595,N_2812,N_2432);
and U4596 (N_4596,N_2292,N_2465);
nor U4597 (N_4597,N_3233,N_3367);
or U4598 (N_4598,N_2559,N_2817);
nor U4599 (N_4599,N_2571,N_3761);
nand U4600 (N_4600,N_2615,N_2486);
nand U4601 (N_4601,N_3857,N_2443);
nor U4602 (N_4602,N_3939,N_2894);
and U4603 (N_4603,N_2726,N_3069);
and U4604 (N_4604,N_3123,N_2592);
nand U4605 (N_4605,N_3481,N_2731);
nor U4606 (N_4606,N_3958,N_3277);
and U4607 (N_4607,N_3768,N_2325);
or U4608 (N_4608,N_2596,N_2466);
xor U4609 (N_4609,N_3384,N_3485);
and U4610 (N_4610,N_3954,N_3524);
nand U4611 (N_4611,N_2734,N_2544);
and U4612 (N_4612,N_2210,N_3652);
nor U4613 (N_4613,N_3333,N_2441);
or U4614 (N_4614,N_3630,N_3023);
nand U4615 (N_4615,N_3171,N_3350);
nand U4616 (N_4616,N_3941,N_2090);
and U4617 (N_4617,N_2892,N_2450);
nand U4618 (N_4618,N_2828,N_2757);
nor U4619 (N_4619,N_3178,N_2263);
nand U4620 (N_4620,N_2811,N_3478);
nor U4621 (N_4621,N_2930,N_2195);
xor U4622 (N_4622,N_2708,N_2270);
xor U4623 (N_4623,N_3558,N_3971);
xor U4624 (N_4624,N_2801,N_3815);
and U4625 (N_4625,N_3856,N_2785);
nor U4626 (N_4626,N_2412,N_3246);
nand U4627 (N_4627,N_2599,N_2329);
nor U4628 (N_4628,N_2324,N_2436);
xnor U4629 (N_4629,N_3774,N_3474);
or U4630 (N_4630,N_3653,N_3078);
xnor U4631 (N_4631,N_2242,N_3516);
or U4632 (N_4632,N_3886,N_2265);
or U4633 (N_4633,N_2836,N_2995);
or U4634 (N_4634,N_2840,N_3328);
nor U4635 (N_4635,N_3198,N_3610);
or U4636 (N_4636,N_2005,N_2220);
xor U4637 (N_4637,N_3451,N_2172);
or U4638 (N_4638,N_3644,N_3355);
nor U4639 (N_4639,N_2613,N_2897);
nor U4640 (N_4640,N_2841,N_3300);
or U4641 (N_4641,N_2872,N_2605);
nand U4642 (N_4642,N_3624,N_3787);
or U4643 (N_4643,N_3259,N_3537);
and U4644 (N_4644,N_2338,N_2937);
nand U4645 (N_4645,N_3489,N_3617);
and U4646 (N_4646,N_3090,N_2848);
nor U4647 (N_4647,N_2689,N_2722);
or U4648 (N_4648,N_3106,N_3081);
and U4649 (N_4649,N_2137,N_3636);
and U4650 (N_4650,N_2845,N_3922);
nor U4651 (N_4651,N_2859,N_2686);
and U4652 (N_4652,N_2182,N_3024);
or U4653 (N_4653,N_2451,N_2404);
nor U4654 (N_4654,N_2967,N_2756);
or U4655 (N_4655,N_2521,N_3897);
nor U4656 (N_4656,N_3408,N_2498);
and U4657 (N_4657,N_3996,N_3756);
nand U4658 (N_4658,N_3161,N_3670);
or U4659 (N_4659,N_2568,N_2925);
and U4660 (N_4660,N_3782,N_3479);
or U4661 (N_4661,N_3045,N_3737);
and U4662 (N_4662,N_2924,N_2197);
nand U4663 (N_4663,N_2491,N_2038);
nand U4664 (N_4664,N_3470,N_3590);
or U4665 (N_4665,N_3740,N_3293);
nor U4666 (N_4666,N_2671,N_3759);
and U4667 (N_4667,N_3281,N_2989);
and U4668 (N_4668,N_2399,N_2868);
nor U4669 (N_4669,N_3032,N_2587);
nand U4670 (N_4670,N_2869,N_3781);
nor U4671 (N_4671,N_3925,N_2022);
nand U4672 (N_4672,N_3213,N_2192);
nor U4673 (N_4673,N_3518,N_3393);
xor U4674 (N_4674,N_2346,N_2532);
and U4675 (N_4675,N_2143,N_3705);
or U4676 (N_4676,N_3575,N_3522);
or U4677 (N_4677,N_3909,N_2044);
nand U4678 (N_4678,N_3313,N_3268);
nand U4679 (N_4679,N_2984,N_3826);
xnor U4680 (N_4680,N_2624,N_3401);
nand U4681 (N_4681,N_3614,N_2496);
or U4682 (N_4682,N_2691,N_2154);
and U4683 (N_4683,N_3684,N_3772);
or U4684 (N_4684,N_2959,N_2150);
nand U4685 (N_4685,N_2820,N_2777);
xnor U4686 (N_4686,N_2340,N_2485);
xnor U4687 (N_4687,N_3648,N_3716);
nor U4688 (N_4688,N_3635,N_3615);
or U4689 (N_4689,N_2028,N_2029);
and U4690 (N_4690,N_3225,N_2551);
or U4691 (N_4691,N_3051,N_2312);
nor U4692 (N_4692,N_2861,N_3915);
and U4693 (N_4693,N_3456,N_3991);
nand U4694 (N_4694,N_2917,N_2136);
or U4695 (N_4695,N_3194,N_3306);
xor U4696 (N_4696,N_2331,N_2365);
xor U4697 (N_4697,N_3436,N_3776);
or U4698 (N_4698,N_3952,N_2053);
nand U4699 (N_4699,N_3001,N_2704);
nand U4700 (N_4700,N_2273,N_2738);
or U4701 (N_4701,N_2926,N_2015);
and U4702 (N_4702,N_3510,N_2330);
nor U4703 (N_4703,N_3097,N_2714);
xnor U4704 (N_4704,N_3731,N_2522);
nor U4705 (N_4705,N_2842,N_2259);
and U4706 (N_4706,N_2541,N_3070);
nor U4707 (N_4707,N_2717,N_2705);
and U4708 (N_4708,N_2784,N_2891);
nand U4709 (N_4709,N_3153,N_3475);
and U4710 (N_4710,N_2945,N_3833);
and U4711 (N_4711,N_3656,N_2519);
nand U4712 (N_4712,N_2603,N_2918);
nand U4713 (N_4713,N_3603,N_3890);
xnor U4714 (N_4714,N_2740,N_2870);
xor U4715 (N_4715,N_3471,N_2941);
nand U4716 (N_4716,N_2164,N_2850);
nand U4717 (N_4717,N_3701,N_3103);
or U4718 (N_4718,N_2543,N_2099);
and U4719 (N_4719,N_3255,N_3651);
nand U4720 (N_4720,N_3878,N_3228);
nor U4721 (N_4721,N_3531,N_3312);
or U4722 (N_4722,N_2094,N_3302);
nand U4723 (N_4723,N_3226,N_2402);
and U4724 (N_4724,N_2677,N_2914);
nor U4725 (N_4725,N_2667,N_2607);
nand U4726 (N_4726,N_2637,N_3443);
xor U4727 (N_4727,N_3174,N_3309);
nand U4728 (N_4728,N_3018,N_3769);
or U4729 (N_4729,N_2003,N_3218);
nand U4730 (N_4730,N_3751,N_3389);
and U4731 (N_4731,N_2493,N_2089);
nor U4732 (N_4732,N_3536,N_3276);
nor U4733 (N_4733,N_3953,N_3132);
nor U4734 (N_4734,N_3430,N_2148);
nand U4735 (N_4735,N_3661,N_2682);
or U4736 (N_4736,N_3800,N_2921);
or U4737 (N_4737,N_3083,N_2318);
or U4738 (N_4738,N_3569,N_2663);
or U4739 (N_4739,N_3195,N_3549);
or U4740 (N_4740,N_2351,N_3647);
nor U4741 (N_4741,N_2743,N_2904);
xor U4742 (N_4742,N_2484,N_3383);
and U4743 (N_4743,N_2081,N_2482);
nand U4744 (N_4744,N_2827,N_2271);
nand U4745 (N_4745,N_3741,N_2306);
or U4746 (N_4746,N_3168,N_2358);
nand U4747 (N_4747,N_2408,N_3983);
xor U4748 (N_4748,N_2824,N_3363);
and U4749 (N_4749,N_3398,N_2912);
nand U4750 (N_4750,N_2628,N_3404);
nand U4751 (N_4751,N_2505,N_2073);
nand U4752 (N_4752,N_2076,N_3882);
xnor U4753 (N_4753,N_2180,N_3390);
or U4754 (N_4754,N_2184,N_3634);
xnor U4755 (N_4755,N_2031,N_2014);
or U4756 (N_4756,N_2231,N_2611);
or U4757 (N_4757,N_3269,N_2557);
nor U4758 (N_4758,N_3109,N_3728);
xnor U4759 (N_4759,N_2766,N_3771);
and U4760 (N_4760,N_3700,N_2260);
and U4761 (N_4761,N_3765,N_2503);
and U4762 (N_4762,N_3091,N_3370);
xor U4763 (N_4763,N_3124,N_3876);
nand U4764 (N_4764,N_3685,N_2050);
or U4765 (N_4765,N_3459,N_2695);
nor U4766 (N_4766,N_3381,N_3956);
or U4767 (N_4767,N_2649,N_2831);
and U4768 (N_4768,N_2527,N_3817);
nand U4769 (N_4769,N_3402,N_2896);
nand U4770 (N_4770,N_3865,N_3935);
and U4771 (N_4771,N_2178,N_2563);
and U4772 (N_4772,N_3042,N_2530);
and U4773 (N_4773,N_3629,N_3979);
or U4774 (N_4774,N_2822,N_3466);
nand U4775 (N_4775,N_3064,N_2008);
nor U4776 (N_4776,N_3810,N_3757);
nand U4777 (N_4777,N_3898,N_3329);
nor U4778 (N_4778,N_3399,N_3578);
xnor U4779 (N_4779,N_2881,N_2202);
nand U4780 (N_4780,N_3128,N_3864);
and U4781 (N_4781,N_2185,N_2110);
nand U4782 (N_4782,N_2000,N_3512);
or U4783 (N_4783,N_2313,N_2654);
nor U4784 (N_4784,N_2939,N_2701);
nand U4785 (N_4785,N_2289,N_3726);
and U4786 (N_4786,N_3770,N_2163);
nor U4787 (N_4787,N_2393,N_2370);
nor U4788 (N_4788,N_2669,N_2666);
nand U4789 (N_4789,N_3172,N_3222);
xor U4790 (N_4790,N_2314,N_3366);
nor U4791 (N_4791,N_2013,N_2871);
or U4792 (N_4792,N_2065,N_2838);
xor U4793 (N_4793,N_3786,N_3292);
nand U4794 (N_4794,N_3509,N_3272);
nand U4795 (N_4795,N_2397,N_3946);
nand U4796 (N_4796,N_3932,N_2632);
or U4797 (N_4797,N_2885,N_2531);
nand U4798 (N_4798,N_3339,N_3989);
and U4799 (N_4799,N_2074,N_2256);
and U4800 (N_4800,N_2877,N_3694);
or U4801 (N_4801,N_3207,N_2656);
and U4802 (N_4802,N_3428,N_3085);
or U4803 (N_4803,N_3895,N_2162);
and U4804 (N_4804,N_3435,N_3752);
nor U4805 (N_4805,N_3587,N_2488);
or U4806 (N_4806,N_3348,N_2997);
nand U4807 (N_4807,N_2428,N_2962);
and U4808 (N_4808,N_3525,N_2795);
nor U4809 (N_4809,N_3959,N_3493);
nor U4810 (N_4810,N_3201,N_3219);
nor U4811 (N_4811,N_2529,N_3113);
or U4812 (N_4812,N_3044,N_2367);
nand U4813 (N_4813,N_2476,N_2333);
nand U4814 (N_4814,N_2567,N_3735);
and U4815 (N_4815,N_2042,N_3217);
and U4816 (N_4816,N_2858,N_3455);
and U4817 (N_4817,N_2694,N_3320);
or U4818 (N_4818,N_2236,N_3957);
or U4819 (N_4819,N_3852,N_3805);
nand U4820 (N_4820,N_2345,N_2558);
nor U4821 (N_4821,N_3526,N_3499);
nor U4822 (N_4822,N_2382,N_2535);
xnor U4823 (N_4823,N_3159,N_2296);
or U4824 (N_4824,N_2109,N_2284);
and U4825 (N_4825,N_2534,N_2080);
and U4826 (N_4826,N_3607,N_3209);
or U4827 (N_4827,N_2602,N_3951);
or U4828 (N_4828,N_3048,N_2847);
nand U4829 (N_4829,N_2138,N_2956);
xor U4830 (N_4830,N_3658,N_3746);
nor U4831 (N_4831,N_3777,N_3167);
or U4832 (N_4832,N_2117,N_3140);
nand U4833 (N_4833,N_3303,N_3717);
nor U4834 (N_4834,N_2513,N_2523);
nand U4835 (N_4835,N_3467,N_3885);
and U4836 (N_4836,N_3990,N_3664);
and U4837 (N_4837,N_3955,N_3072);
nand U4838 (N_4838,N_3062,N_3982);
xor U4839 (N_4839,N_3162,N_2687);
and U4840 (N_4840,N_2773,N_3273);
nand U4841 (N_4841,N_2747,N_3669);
or U4842 (N_4842,N_3149,N_2445);
and U4843 (N_4843,N_3821,N_3539);
nor U4844 (N_4844,N_2380,N_2920);
nor U4845 (N_4845,N_3734,N_3863);
nor U4846 (N_4846,N_3866,N_2833);
nor U4847 (N_4847,N_3084,N_2121);
nand U4848 (N_4848,N_2793,N_3385);
nand U4849 (N_4849,N_3719,N_2021);
or U4850 (N_4850,N_2916,N_2919);
nor U4851 (N_4851,N_2100,N_2648);
nand U4852 (N_4852,N_3205,N_3906);
or U4853 (N_4853,N_2288,N_3151);
nand U4854 (N_4854,N_2819,N_2981);
nand U4855 (N_4855,N_3119,N_2374);
or U4856 (N_4856,N_3595,N_3715);
xor U4857 (N_4857,N_3654,N_3447);
nor U4858 (N_4858,N_2501,N_2982);
or U4859 (N_4859,N_2506,N_2639);
xor U4860 (N_4860,N_2634,N_2764);
nand U4861 (N_4861,N_2419,N_3597);
or U4862 (N_4862,N_2356,N_2579);
nand U4863 (N_4863,N_3627,N_3611);
or U4864 (N_4864,N_3364,N_3682);
nand U4865 (N_4865,N_3993,N_2101);
xor U4866 (N_4866,N_2915,N_3504);
or U4867 (N_4867,N_3736,N_3036);
nand U4868 (N_4868,N_2416,N_3513);
nand U4869 (N_4869,N_2495,N_3369);
xor U4870 (N_4870,N_2064,N_2036);
xnor U4871 (N_4871,N_2561,N_2609);
or U4872 (N_4872,N_2454,N_3555);
nand U4873 (N_4873,N_2884,N_2391);
or U4874 (N_4874,N_2690,N_2814);
nand U4875 (N_4875,N_3331,N_3200);
nand U4876 (N_4876,N_3027,N_3362);
nand U4877 (N_4877,N_3026,N_3937);
nor U4878 (N_4878,N_3921,N_3660);
or U4879 (N_4879,N_3465,N_3108);
nand U4880 (N_4880,N_3014,N_3593);
xnor U4881 (N_4881,N_3278,N_3041);
nor U4882 (N_4882,N_2175,N_3407);
nand U4883 (N_4883,N_2626,N_3411);
or U4884 (N_4884,N_2960,N_3742);
or U4885 (N_4885,N_2964,N_2084);
nor U4886 (N_4886,N_3403,N_3251);
and U4887 (N_4887,N_3903,N_3564);
nor U4888 (N_4888,N_2650,N_3025);
or U4889 (N_4889,N_3323,N_2553);
and U4890 (N_4890,N_3141,N_3013);
xor U4891 (N_4891,N_2931,N_2307);
nor U4892 (N_4892,N_3708,N_3150);
or U4893 (N_4893,N_2198,N_3733);
and U4894 (N_4894,N_3998,N_3449);
and U4895 (N_4895,N_2134,N_3966);
or U4896 (N_4896,N_2347,N_2437);
and U4897 (N_4897,N_3388,N_3835);
or U4898 (N_4898,N_2294,N_2835);
and U4899 (N_4899,N_3065,N_2291);
or U4900 (N_4900,N_3220,N_3243);
nor U4901 (N_4901,N_3211,N_3133);
nor U4902 (N_4902,N_3545,N_2601);
nor U4903 (N_4903,N_3722,N_2664);
or U4904 (N_4904,N_2130,N_3712);
nand U4905 (N_4905,N_3022,N_2439);
nor U4906 (N_4906,N_2750,N_2444);
nand U4907 (N_4907,N_2247,N_3305);
xnor U4908 (N_4908,N_3286,N_2658);
nor U4909 (N_4909,N_3265,N_3543);
xnor U4910 (N_4910,N_3111,N_3605);
nand U4911 (N_4911,N_2790,N_2940);
nor U4912 (N_4912,N_2224,N_3317);
nand U4913 (N_4913,N_3521,N_3936);
nor U4914 (N_4914,N_3994,N_3039);
nor U4915 (N_4915,N_3930,N_2024);
xor U4916 (N_4916,N_3547,N_3100);
nor U4917 (N_4917,N_3928,N_2999);
nand U4918 (N_4918,N_2806,N_2315);
or U4919 (N_4919,N_3423,N_2194);
nand U4920 (N_4920,N_2388,N_3668);
nand U4921 (N_4921,N_3929,N_2644);
or U4922 (N_4922,N_2680,N_2955);
or U4923 (N_4923,N_3412,N_2078);
or U4924 (N_4924,N_2406,N_3206);
and U4925 (N_4925,N_3262,N_3426);
or U4926 (N_4926,N_3783,N_3999);
nor U4927 (N_4927,N_3919,N_3053);
nand U4928 (N_4928,N_3173,N_3118);
nor U4929 (N_4929,N_3534,N_3686);
and U4930 (N_4930,N_2300,N_2390);
xor U4931 (N_4931,N_3318,N_3445);
nor U4932 (N_4932,N_3873,N_3406);
and U4933 (N_4933,N_2139,N_2737);
nor U4934 (N_4934,N_2276,N_3532);
and U4935 (N_4935,N_2767,N_2341);
and U4936 (N_4936,N_3322,N_3541);
nor U4937 (N_4937,N_3544,N_3837);
nand U4938 (N_4938,N_3511,N_2616);
xor U4939 (N_4939,N_3623,N_3413);
nor U4940 (N_4940,N_2665,N_3029);
nand U4941 (N_4941,N_3579,N_3729);
nor U4942 (N_4942,N_3616,N_3987);
nand U4943 (N_4943,N_3294,N_2494);
or U4944 (N_4944,N_3551,N_3116);
nand U4945 (N_4945,N_2239,N_2310);
nand U4946 (N_4946,N_2713,N_3944);
and U4947 (N_4947,N_3913,N_3568);
or U4948 (N_4948,N_3340,N_2538);
nand U4949 (N_4949,N_3287,N_3327);
and U4950 (N_4950,N_3600,N_3902);
nand U4951 (N_4951,N_3204,N_3452);
nor U4952 (N_4952,N_3054,N_3378);
and U4953 (N_4953,N_3283,N_3687);
xor U4954 (N_4954,N_3439,N_3602);
nand U4955 (N_4955,N_3121,N_2487);
or U4956 (N_4956,N_3432,N_2301);
and U4957 (N_4957,N_3743,N_3242);
nand U4958 (N_4958,N_2299,N_3596);
nor U4959 (N_4959,N_2147,N_2810);
and U4960 (N_4960,N_3931,N_3386);
xor U4961 (N_4961,N_2507,N_2575);
nor U4962 (N_4962,N_2653,N_2246);
or U4963 (N_4963,N_3082,N_3871);
or U4964 (N_4964,N_2051,N_2396);
or U4965 (N_4965,N_2633,N_3169);
xnor U4966 (N_4966,N_3486,N_3248);
and U4967 (N_4967,N_2770,N_2035);
or U4968 (N_4968,N_2058,N_2949);
or U4969 (N_4969,N_2752,N_3266);
or U4970 (N_4970,N_3899,N_2229);
nand U4971 (N_4971,N_3494,N_2463);
nand U4972 (N_4972,N_2803,N_2578);
nor U4973 (N_4973,N_2798,N_3400);
and U4974 (N_4974,N_2950,N_3625);
or U4975 (N_4975,N_3667,N_2782);
or U4976 (N_4976,N_2118,N_3372);
and U4977 (N_4977,N_2525,N_3427);
or U4978 (N_4978,N_2362,N_3673);
xnor U4979 (N_4979,N_2768,N_3582);
or U4980 (N_4980,N_3325,N_2409);
or U4981 (N_4981,N_2196,N_3912);
nor U4982 (N_4982,N_2804,N_2274);
nor U4983 (N_4983,N_2555,N_2863);
nor U4984 (N_4984,N_2016,N_2593);
or U4985 (N_4985,N_3125,N_3632);
nor U4986 (N_4986,N_3038,N_2800);
nand U4987 (N_4987,N_2843,N_3858);
xor U4988 (N_4988,N_3645,N_2712);
or U4989 (N_4989,N_2597,N_2540);
nand U4990 (N_4990,N_2457,N_2264);
and U4991 (N_4991,N_2280,N_3058);
or U4992 (N_4992,N_3923,N_3974);
nor U4993 (N_4993,N_3696,N_3621);
or U4994 (N_4994,N_3104,N_2334);
or U4995 (N_4995,N_2913,N_3077);
and U4996 (N_4996,N_3496,N_2057);
xnor U4997 (N_4997,N_3152,N_2190);
or U4998 (N_4998,N_2702,N_2126);
xor U4999 (N_4999,N_3295,N_2272);
or U5000 (N_5000,N_2953,N_2830);
or U5001 (N_5001,N_2267,N_3391);
nor U5002 (N_5002,N_2880,N_2925);
nor U5003 (N_5003,N_2330,N_3331);
or U5004 (N_5004,N_2132,N_2781);
or U5005 (N_5005,N_3955,N_2358);
and U5006 (N_5006,N_3280,N_2346);
and U5007 (N_5007,N_2965,N_2930);
or U5008 (N_5008,N_3513,N_2683);
or U5009 (N_5009,N_2410,N_3633);
nor U5010 (N_5010,N_2485,N_3456);
nand U5011 (N_5011,N_3202,N_2957);
or U5012 (N_5012,N_3562,N_3175);
nor U5013 (N_5013,N_3645,N_3065);
and U5014 (N_5014,N_2093,N_3609);
nor U5015 (N_5015,N_2503,N_3722);
and U5016 (N_5016,N_2188,N_3256);
and U5017 (N_5017,N_2019,N_2978);
nand U5018 (N_5018,N_3232,N_2146);
nand U5019 (N_5019,N_2511,N_2452);
or U5020 (N_5020,N_3434,N_3281);
or U5021 (N_5021,N_2875,N_3395);
and U5022 (N_5022,N_2506,N_2129);
nor U5023 (N_5023,N_2930,N_2841);
and U5024 (N_5024,N_3455,N_2364);
nor U5025 (N_5025,N_2539,N_2570);
nand U5026 (N_5026,N_2467,N_3829);
or U5027 (N_5027,N_2949,N_3062);
xor U5028 (N_5028,N_2192,N_3677);
nand U5029 (N_5029,N_3295,N_3419);
nand U5030 (N_5030,N_2738,N_3826);
and U5031 (N_5031,N_2177,N_2184);
and U5032 (N_5032,N_2494,N_2311);
nor U5033 (N_5033,N_2122,N_3627);
or U5034 (N_5034,N_2010,N_3012);
and U5035 (N_5035,N_3804,N_2333);
nand U5036 (N_5036,N_2993,N_2027);
nand U5037 (N_5037,N_3326,N_2701);
or U5038 (N_5038,N_3547,N_2363);
or U5039 (N_5039,N_2399,N_3985);
or U5040 (N_5040,N_3702,N_3298);
nor U5041 (N_5041,N_3074,N_3308);
or U5042 (N_5042,N_3816,N_2065);
nor U5043 (N_5043,N_3351,N_3684);
and U5044 (N_5044,N_3251,N_3677);
or U5045 (N_5045,N_3001,N_2541);
and U5046 (N_5046,N_2106,N_3915);
nor U5047 (N_5047,N_3567,N_2614);
xnor U5048 (N_5048,N_2664,N_3026);
nand U5049 (N_5049,N_3940,N_2714);
and U5050 (N_5050,N_3740,N_3176);
xnor U5051 (N_5051,N_3928,N_3500);
and U5052 (N_5052,N_3962,N_3179);
or U5053 (N_5053,N_3788,N_2437);
and U5054 (N_5054,N_3010,N_3884);
or U5055 (N_5055,N_3277,N_2947);
and U5056 (N_5056,N_2249,N_3738);
nand U5057 (N_5057,N_2531,N_3483);
nor U5058 (N_5058,N_3497,N_3489);
nor U5059 (N_5059,N_3435,N_3992);
nand U5060 (N_5060,N_2608,N_3495);
nand U5061 (N_5061,N_3724,N_2547);
or U5062 (N_5062,N_2372,N_2473);
nand U5063 (N_5063,N_2530,N_2328);
nor U5064 (N_5064,N_2374,N_3190);
or U5065 (N_5065,N_2065,N_2204);
xnor U5066 (N_5066,N_3041,N_2750);
nand U5067 (N_5067,N_2625,N_2440);
nor U5068 (N_5068,N_2868,N_2584);
or U5069 (N_5069,N_3456,N_2774);
nand U5070 (N_5070,N_3477,N_2707);
or U5071 (N_5071,N_2807,N_3570);
nand U5072 (N_5072,N_3027,N_2448);
nor U5073 (N_5073,N_2092,N_2327);
and U5074 (N_5074,N_3737,N_3273);
nor U5075 (N_5075,N_2955,N_3434);
or U5076 (N_5076,N_3788,N_2644);
and U5077 (N_5077,N_2740,N_2501);
nand U5078 (N_5078,N_2483,N_3561);
nand U5079 (N_5079,N_3547,N_3159);
and U5080 (N_5080,N_3389,N_2181);
or U5081 (N_5081,N_3594,N_3385);
nor U5082 (N_5082,N_3762,N_2665);
nand U5083 (N_5083,N_3467,N_3432);
nor U5084 (N_5084,N_3743,N_3381);
nand U5085 (N_5085,N_3194,N_3211);
or U5086 (N_5086,N_2844,N_3714);
or U5087 (N_5087,N_2302,N_3512);
nand U5088 (N_5088,N_3375,N_3807);
nor U5089 (N_5089,N_2704,N_2886);
nor U5090 (N_5090,N_2121,N_2925);
and U5091 (N_5091,N_2484,N_3175);
or U5092 (N_5092,N_2110,N_3573);
or U5093 (N_5093,N_2679,N_2139);
nor U5094 (N_5094,N_2723,N_2819);
and U5095 (N_5095,N_2556,N_3109);
nor U5096 (N_5096,N_3301,N_2597);
or U5097 (N_5097,N_3529,N_2806);
or U5098 (N_5098,N_2373,N_2829);
xnor U5099 (N_5099,N_2833,N_3037);
and U5100 (N_5100,N_3609,N_2619);
xor U5101 (N_5101,N_3205,N_3420);
nand U5102 (N_5102,N_3384,N_2451);
or U5103 (N_5103,N_2880,N_2160);
and U5104 (N_5104,N_3542,N_2765);
and U5105 (N_5105,N_3121,N_3722);
xnor U5106 (N_5106,N_3213,N_3732);
and U5107 (N_5107,N_2374,N_3278);
or U5108 (N_5108,N_2795,N_3678);
or U5109 (N_5109,N_3085,N_3533);
xnor U5110 (N_5110,N_3680,N_2920);
and U5111 (N_5111,N_2485,N_2676);
or U5112 (N_5112,N_2805,N_3296);
nand U5113 (N_5113,N_2270,N_2151);
nand U5114 (N_5114,N_2431,N_3330);
nand U5115 (N_5115,N_3924,N_3321);
or U5116 (N_5116,N_3137,N_3690);
or U5117 (N_5117,N_3450,N_3566);
nor U5118 (N_5118,N_3512,N_3011);
and U5119 (N_5119,N_3062,N_2307);
or U5120 (N_5120,N_2804,N_2857);
nand U5121 (N_5121,N_2438,N_2179);
or U5122 (N_5122,N_2303,N_2503);
nor U5123 (N_5123,N_3159,N_2281);
nor U5124 (N_5124,N_2260,N_3749);
nor U5125 (N_5125,N_3606,N_3052);
or U5126 (N_5126,N_2054,N_2707);
or U5127 (N_5127,N_3543,N_2394);
nor U5128 (N_5128,N_2219,N_2603);
or U5129 (N_5129,N_3159,N_2431);
nand U5130 (N_5130,N_2088,N_2360);
nand U5131 (N_5131,N_3313,N_3685);
nand U5132 (N_5132,N_2517,N_2671);
nand U5133 (N_5133,N_2416,N_3960);
xnor U5134 (N_5134,N_3526,N_3763);
or U5135 (N_5135,N_3029,N_2439);
or U5136 (N_5136,N_3595,N_2740);
or U5137 (N_5137,N_3422,N_3818);
nand U5138 (N_5138,N_3589,N_2541);
or U5139 (N_5139,N_2853,N_2502);
and U5140 (N_5140,N_2788,N_3160);
nor U5141 (N_5141,N_2907,N_2633);
and U5142 (N_5142,N_3186,N_2594);
or U5143 (N_5143,N_3954,N_3860);
or U5144 (N_5144,N_2214,N_3473);
nor U5145 (N_5145,N_2183,N_2424);
xnor U5146 (N_5146,N_3328,N_2230);
nor U5147 (N_5147,N_3807,N_2667);
or U5148 (N_5148,N_3749,N_2254);
or U5149 (N_5149,N_2357,N_2437);
xor U5150 (N_5150,N_3153,N_3297);
nor U5151 (N_5151,N_2383,N_2177);
xnor U5152 (N_5152,N_3979,N_2202);
and U5153 (N_5153,N_3776,N_3598);
or U5154 (N_5154,N_2868,N_3904);
nor U5155 (N_5155,N_2206,N_2345);
nand U5156 (N_5156,N_2885,N_3619);
or U5157 (N_5157,N_3271,N_2928);
nand U5158 (N_5158,N_3632,N_2800);
nand U5159 (N_5159,N_2547,N_3479);
or U5160 (N_5160,N_3193,N_3106);
and U5161 (N_5161,N_2718,N_3060);
nor U5162 (N_5162,N_3880,N_3738);
xnor U5163 (N_5163,N_2105,N_2290);
and U5164 (N_5164,N_3721,N_2927);
nor U5165 (N_5165,N_2558,N_3486);
nor U5166 (N_5166,N_2753,N_3728);
and U5167 (N_5167,N_2937,N_2846);
nor U5168 (N_5168,N_3075,N_3542);
nor U5169 (N_5169,N_2953,N_3241);
nor U5170 (N_5170,N_2003,N_2883);
or U5171 (N_5171,N_3457,N_3020);
nor U5172 (N_5172,N_3452,N_2632);
nor U5173 (N_5173,N_3334,N_3699);
and U5174 (N_5174,N_3138,N_2950);
nand U5175 (N_5175,N_2969,N_3314);
and U5176 (N_5176,N_3617,N_2173);
and U5177 (N_5177,N_2862,N_2613);
nor U5178 (N_5178,N_3345,N_3512);
and U5179 (N_5179,N_2335,N_2453);
nor U5180 (N_5180,N_3205,N_2654);
nand U5181 (N_5181,N_2823,N_2550);
nor U5182 (N_5182,N_3461,N_2485);
nor U5183 (N_5183,N_2436,N_2840);
nand U5184 (N_5184,N_3228,N_3197);
xnor U5185 (N_5185,N_2537,N_3547);
or U5186 (N_5186,N_2279,N_3852);
or U5187 (N_5187,N_3135,N_3184);
or U5188 (N_5188,N_2808,N_2006);
or U5189 (N_5189,N_3334,N_2287);
and U5190 (N_5190,N_2184,N_3161);
nor U5191 (N_5191,N_3371,N_3735);
and U5192 (N_5192,N_2270,N_3614);
or U5193 (N_5193,N_3049,N_3989);
and U5194 (N_5194,N_2707,N_2109);
nor U5195 (N_5195,N_3119,N_3941);
nand U5196 (N_5196,N_2078,N_3834);
or U5197 (N_5197,N_3408,N_3766);
xnor U5198 (N_5198,N_2478,N_3889);
nor U5199 (N_5199,N_3145,N_3926);
xor U5200 (N_5200,N_2835,N_3241);
and U5201 (N_5201,N_3681,N_2995);
and U5202 (N_5202,N_3520,N_3951);
and U5203 (N_5203,N_2954,N_2973);
or U5204 (N_5204,N_3076,N_2269);
or U5205 (N_5205,N_3632,N_3043);
nand U5206 (N_5206,N_3454,N_3771);
or U5207 (N_5207,N_2232,N_2464);
xnor U5208 (N_5208,N_2397,N_3531);
or U5209 (N_5209,N_3159,N_3956);
and U5210 (N_5210,N_2885,N_2075);
nor U5211 (N_5211,N_3191,N_3109);
and U5212 (N_5212,N_2606,N_3539);
nor U5213 (N_5213,N_3894,N_2794);
nand U5214 (N_5214,N_2662,N_3317);
or U5215 (N_5215,N_2952,N_3824);
nor U5216 (N_5216,N_3927,N_2318);
nand U5217 (N_5217,N_3123,N_2336);
xnor U5218 (N_5218,N_2549,N_3271);
nand U5219 (N_5219,N_3677,N_3276);
or U5220 (N_5220,N_2054,N_3021);
nor U5221 (N_5221,N_3164,N_3885);
or U5222 (N_5222,N_2088,N_3840);
nand U5223 (N_5223,N_2673,N_2579);
and U5224 (N_5224,N_2780,N_3776);
or U5225 (N_5225,N_3104,N_2598);
or U5226 (N_5226,N_2213,N_2712);
or U5227 (N_5227,N_2298,N_2787);
nor U5228 (N_5228,N_3301,N_3135);
and U5229 (N_5229,N_2311,N_2593);
and U5230 (N_5230,N_2974,N_2477);
and U5231 (N_5231,N_3455,N_2532);
nand U5232 (N_5232,N_2019,N_3574);
and U5233 (N_5233,N_3043,N_3771);
and U5234 (N_5234,N_3028,N_2609);
xor U5235 (N_5235,N_3446,N_3036);
nor U5236 (N_5236,N_2735,N_3030);
and U5237 (N_5237,N_2739,N_2267);
nor U5238 (N_5238,N_2128,N_2734);
or U5239 (N_5239,N_3619,N_2110);
or U5240 (N_5240,N_2002,N_2816);
or U5241 (N_5241,N_3371,N_2767);
and U5242 (N_5242,N_2692,N_3941);
nor U5243 (N_5243,N_2818,N_2797);
or U5244 (N_5244,N_2609,N_3161);
or U5245 (N_5245,N_3331,N_3375);
or U5246 (N_5246,N_3665,N_2668);
nor U5247 (N_5247,N_2269,N_3546);
nand U5248 (N_5248,N_3555,N_2394);
xnor U5249 (N_5249,N_3915,N_2344);
nor U5250 (N_5250,N_3040,N_2953);
nor U5251 (N_5251,N_2303,N_3869);
nand U5252 (N_5252,N_2782,N_3732);
and U5253 (N_5253,N_2179,N_2431);
and U5254 (N_5254,N_3452,N_2815);
nand U5255 (N_5255,N_2945,N_2866);
or U5256 (N_5256,N_3382,N_3406);
nand U5257 (N_5257,N_2633,N_2582);
xor U5258 (N_5258,N_3601,N_2761);
nor U5259 (N_5259,N_2262,N_3354);
xor U5260 (N_5260,N_3213,N_3236);
nand U5261 (N_5261,N_2106,N_2760);
or U5262 (N_5262,N_2439,N_2299);
and U5263 (N_5263,N_2114,N_3944);
or U5264 (N_5264,N_2333,N_2817);
and U5265 (N_5265,N_3421,N_3372);
and U5266 (N_5266,N_3475,N_2157);
or U5267 (N_5267,N_2584,N_3836);
or U5268 (N_5268,N_3476,N_3304);
nor U5269 (N_5269,N_3086,N_2327);
nor U5270 (N_5270,N_3235,N_3111);
or U5271 (N_5271,N_2404,N_2093);
xor U5272 (N_5272,N_3846,N_3602);
nand U5273 (N_5273,N_3856,N_2512);
nor U5274 (N_5274,N_3314,N_3293);
or U5275 (N_5275,N_3136,N_2297);
nand U5276 (N_5276,N_3627,N_2337);
nand U5277 (N_5277,N_3429,N_3295);
and U5278 (N_5278,N_3783,N_3422);
xor U5279 (N_5279,N_2461,N_2400);
nor U5280 (N_5280,N_2680,N_2246);
nand U5281 (N_5281,N_3725,N_3421);
nand U5282 (N_5282,N_3346,N_2795);
xnor U5283 (N_5283,N_3822,N_3813);
nor U5284 (N_5284,N_2280,N_3314);
nor U5285 (N_5285,N_2374,N_3481);
or U5286 (N_5286,N_2866,N_3770);
and U5287 (N_5287,N_2240,N_2003);
or U5288 (N_5288,N_3103,N_3154);
or U5289 (N_5289,N_2873,N_3311);
or U5290 (N_5290,N_3287,N_2305);
and U5291 (N_5291,N_3180,N_3333);
xor U5292 (N_5292,N_3926,N_3049);
and U5293 (N_5293,N_2830,N_3130);
nand U5294 (N_5294,N_3651,N_2766);
nand U5295 (N_5295,N_3239,N_3000);
nor U5296 (N_5296,N_2123,N_2586);
or U5297 (N_5297,N_3367,N_2920);
nor U5298 (N_5298,N_2605,N_3709);
nor U5299 (N_5299,N_2067,N_3090);
and U5300 (N_5300,N_3169,N_2176);
nor U5301 (N_5301,N_2268,N_3283);
xor U5302 (N_5302,N_2867,N_2037);
nor U5303 (N_5303,N_3471,N_3046);
and U5304 (N_5304,N_2540,N_2545);
xnor U5305 (N_5305,N_2782,N_3957);
nand U5306 (N_5306,N_3380,N_2337);
nand U5307 (N_5307,N_3133,N_3855);
and U5308 (N_5308,N_2296,N_3768);
and U5309 (N_5309,N_3481,N_3117);
or U5310 (N_5310,N_3687,N_2514);
and U5311 (N_5311,N_3830,N_3019);
or U5312 (N_5312,N_2216,N_2927);
xnor U5313 (N_5313,N_2662,N_2888);
nand U5314 (N_5314,N_3520,N_2636);
or U5315 (N_5315,N_3446,N_2826);
nor U5316 (N_5316,N_2581,N_2153);
and U5317 (N_5317,N_3716,N_2403);
or U5318 (N_5318,N_2134,N_3429);
nor U5319 (N_5319,N_3620,N_3738);
nor U5320 (N_5320,N_3957,N_3555);
and U5321 (N_5321,N_2333,N_3182);
nand U5322 (N_5322,N_2321,N_2350);
xor U5323 (N_5323,N_3996,N_2607);
or U5324 (N_5324,N_2438,N_3468);
or U5325 (N_5325,N_2381,N_2302);
nor U5326 (N_5326,N_3174,N_2713);
or U5327 (N_5327,N_2488,N_3001);
or U5328 (N_5328,N_3847,N_2205);
nor U5329 (N_5329,N_2963,N_3815);
xor U5330 (N_5330,N_2826,N_3541);
nor U5331 (N_5331,N_3438,N_3267);
or U5332 (N_5332,N_3719,N_3965);
or U5333 (N_5333,N_3987,N_3082);
nand U5334 (N_5334,N_2946,N_2314);
or U5335 (N_5335,N_2298,N_3161);
and U5336 (N_5336,N_2883,N_3184);
nor U5337 (N_5337,N_3528,N_3826);
nor U5338 (N_5338,N_2024,N_2678);
nand U5339 (N_5339,N_2698,N_3539);
xor U5340 (N_5340,N_3904,N_2550);
or U5341 (N_5341,N_2359,N_2411);
and U5342 (N_5342,N_3179,N_2842);
nand U5343 (N_5343,N_3298,N_3198);
and U5344 (N_5344,N_2080,N_2290);
nand U5345 (N_5345,N_2896,N_3467);
and U5346 (N_5346,N_2980,N_2059);
and U5347 (N_5347,N_2922,N_3884);
nor U5348 (N_5348,N_3060,N_3430);
nor U5349 (N_5349,N_3622,N_3854);
or U5350 (N_5350,N_2382,N_3352);
nand U5351 (N_5351,N_2009,N_2312);
or U5352 (N_5352,N_2451,N_2017);
or U5353 (N_5353,N_2603,N_3317);
or U5354 (N_5354,N_2543,N_2805);
and U5355 (N_5355,N_3615,N_2494);
or U5356 (N_5356,N_3538,N_3650);
and U5357 (N_5357,N_3649,N_2250);
nand U5358 (N_5358,N_2842,N_3189);
nor U5359 (N_5359,N_2949,N_3118);
and U5360 (N_5360,N_3010,N_3571);
or U5361 (N_5361,N_3312,N_3900);
nand U5362 (N_5362,N_2986,N_3390);
and U5363 (N_5363,N_3537,N_3812);
nand U5364 (N_5364,N_3398,N_3186);
nand U5365 (N_5365,N_2646,N_2761);
nand U5366 (N_5366,N_3844,N_2861);
nand U5367 (N_5367,N_3890,N_3860);
nor U5368 (N_5368,N_3586,N_2122);
and U5369 (N_5369,N_2269,N_2571);
nor U5370 (N_5370,N_3099,N_2209);
xor U5371 (N_5371,N_3268,N_3029);
or U5372 (N_5372,N_2183,N_2688);
and U5373 (N_5373,N_3286,N_2292);
or U5374 (N_5374,N_2329,N_2718);
and U5375 (N_5375,N_2648,N_3467);
nand U5376 (N_5376,N_2803,N_2259);
nand U5377 (N_5377,N_3083,N_2775);
nor U5378 (N_5378,N_2629,N_2223);
nand U5379 (N_5379,N_2879,N_3575);
xor U5380 (N_5380,N_2896,N_2209);
or U5381 (N_5381,N_2470,N_3953);
xnor U5382 (N_5382,N_3589,N_2577);
nand U5383 (N_5383,N_2752,N_2268);
and U5384 (N_5384,N_2568,N_3423);
and U5385 (N_5385,N_3908,N_3274);
nand U5386 (N_5386,N_3009,N_3798);
and U5387 (N_5387,N_2509,N_3589);
nor U5388 (N_5388,N_3364,N_3769);
or U5389 (N_5389,N_3135,N_2584);
or U5390 (N_5390,N_3138,N_2740);
or U5391 (N_5391,N_2022,N_3280);
and U5392 (N_5392,N_3150,N_3827);
or U5393 (N_5393,N_2774,N_3357);
and U5394 (N_5394,N_3033,N_2086);
nand U5395 (N_5395,N_2499,N_2385);
and U5396 (N_5396,N_3110,N_3423);
and U5397 (N_5397,N_3091,N_3265);
or U5398 (N_5398,N_2941,N_2600);
nand U5399 (N_5399,N_3440,N_3206);
nand U5400 (N_5400,N_3909,N_2535);
nor U5401 (N_5401,N_3614,N_2758);
and U5402 (N_5402,N_3073,N_3089);
or U5403 (N_5403,N_2753,N_3686);
nor U5404 (N_5404,N_2888,N_3382);
and U5405 (N_5405,N_2318,N_3066);
xor U5406 (N_5406,N_2312,N_2933);
or U5407 (N_5407,N_3956,N_3445);
nor U5408 (N_5408,N_3633,N_3184);
xor U5409 (N_5409,N_3745,N_2009);
nand U5410 (N_5410,N_3152,N_2333);
nor U5411 (N_5411,N_3281,N_3508);
and U5412 (N_5412,N_3993,N_3655);
and U5413 (N_5413,N_2473,N_3341);
and U5414 (N_5414,N_2855,N_3265);
and U5415 (N_5415,N_3510,N_3204);
nor U5416 (N_5416,N_3872,N_3765);
xor U5417 (N_5417,N_3145,N_3777);
nand U5418 (N_5418,N_3288,N_2438);
and U5419 (N_5419,N_3884,N_3387);
or U5420 (N_5420,N_3944,N_3895);
nor U5421 (N_5421,N_3332,N_3199);
nand U5422 (N_5422,N_3861,N_3116);
nand U5423 (N_5423,N_3628,N_2229);
nor U5424 (N_5424,N_2142,N_3465);
nand U5425 (N_5425,N_3136,N_2985);
nor U5426 (N_5426,N_3287,N_3972);
or U5427 (N_5427,N_2356,N_3732);
nor U5428 (N_5428,N_2676,N_2918);
and U5429 (N_5429,N_3225,N_3651);
and U5430 (N_5430,N_2101,N_3102);
nor U5431 (N_5431,N_3176,N_3571);
and U5432 (N_5432,N_2721,N_2957);
or U5433 (N_5433,N_3362,N_2792);
and U5434 (N_5434,N_2058,N_3307);
nor U5435 (N_5435,N_2969,N_3170);
nand U5436 (N_5436,N_3905,N_3032);
nor U5437 (N_5437,N_2197,N_2274);
nand U5438 (N_5438,N_2561,N_3289);
nor U5439 (N_5439,N_2053,N_3433);
nor U5440 (N_5440,N_3114,N_2801);
or U5441 (N_5441,N_3828,N_2458);
nand U5442 (N_5442,N_3665,N_3232);
nand U5443 (N_5443,N_2851,N_2567);
xnor U5444 (N_5444,N_3849,N_3785);
nor U5445 (N_5445,N_3644,N_3011);
nand U5446 (N_5446,N_2683,N_2840);
nand U5447 (N_5447,N_3813,N_2471);
nor U5448 (N_5448,N_3337,N_2264);
and U5449 (N_5449,N_2101,N_2162);
nand U5450 (N_5450,N_2116,N_3928);
nand U5451 (N_5451,N_3659,N_3647);
or U5452 (N_5452,N_2529,N_2201);
or U5453 (N_5453,N_2706,N_2426);
and U5454 (N_5454,N_3074,N_2707);
xor U5455 (N_5455,N_3044,N_2495);
and U5456 (N_5456,N_2440,N_3913);
nor U5457 (N_5457,N_2489,N_3148);
and U5458 (N_5458,N_3738,N_2905);
and U5459 (N_5459,N_3424,N_3705);
or U5460 (N_5460,N_2196,N_3875);
nor U5461 (N_5461,N_2175,N_2252);
nand U5462 (N_5462,N_2899,N_3669);
xnor U5463 (N_5463,N_2316,N_3382);
nor U5464 (N_5464,N_3942,N_3175);
or U5465 (N_5465,N_2385,N_2447);
xor U5466 (N_5466,N_3789,N_2676);
and U5467 (N_5467,N_2118,N_3682);
and U5468 (N_5468,N_3361,N_3721);
and U5469 (N_5469,N_2528,N_3521);
and U5470 (N_5470,N_3489,N_2971);
or U5471 (N_5471,N_2580,N_2075);
nand U5472 (N_5472,N_3024,N_3678);
and U5473 (N_5473,N_2191,N_3076);
and U5474 (N_5474,N_2184,N_3775);
or U5475 (N_5475,N_2084,N_2771);
nand U5476 (N_5476,N_3130,N_3543);
nand U5477 (N_5477,N_2336,N_3240);
or U5478 (N_5478,N_2696,N_3830);
nand U5479 (N_5479,N_2843,N_2277);
xor U5480 (N_5480,N_3747,N_2159);
nand U5481 (N_5481,N_3884,N_2422);
xnor U5482 (N_5482,N_2267,N_2831);
and U5483 (N_5483,N_2412,N_3989);
or U5484 (N_5484,N_3762,N_3848);
or U5485 (N_5485,N_3521,N_2150);
or U5486 (N_5486,N_2065,N_2303);
nor U5487 (N_5487,N_2325,N_3219);
nor U5488 (N_5488,N_3980,N_2582);
and U5489 (N_5489,N_2207,N_2144);
and U5490 (N_5490,N_3558,N_2038);
and U5491 (N_5491,N_3059,N_3556);
or U5492 (N_5492,N_3428,N_2696);
or U5493 (N_5493,N_2414,N_3141);
nor U5494 (N_5494,N_2196,N_3290);
xor U5495 (N_5495,N_2901,N_3423);
nand U5496 (N_5496,N_3282,N_3318);
xor U5497 (N_5497,N_2071,N_3692);
nor U5498 (N_5498,N_2783,N_2053);
and U5499 (N_5499,N_2250,N_2825);
nor U5500 (N_5500,N_3048,N_3959);
or U5501 (N_5501,N_2905,N_3244);
or U5502 (N_5502,N_2284,N_3524);
nand U5503 (N_5503,N_3208,N_3257);
or U5504 (N_5504,N_2626,N_3683);
or U5505 (N_5505,N_2934,N_2240);
nand U5506 (N_5506,N_3166,N_3411);
or U5507 (N_5507,N_2946,N_3256);
or U5508 (N_5508,N_3397,N_3273);
nor U5509 (N_5509,N_2420,N_3291);
or U5510 (N_5510,N_2692,N_2795);
or U5511 (N_5511,N_3405,N_3706);
or U5512 (N_5512,N_3229,N_2661);
and U5513 (N_5513,N_3794,N_2406);
and U5514 (N_5514,N_3622,N_2604);
nand U5515 (N_5515,N_2700,N_3691);
nand U5516 (N_5516,N_3527,N_2817);
or U5517 (N_5517,N_2280,N_2165);
or U5518 (N_5518,N_3229,N_2448);
nand U5519 (N_5519,N_2150,N_2600);
or U5520 (N_5520,N_3624,N_3420);
and U5521 (N_5521,N_3729,N_3423);
and U5522 (N_5522,N_3220,N_2798);
nand U5523 (N_5523,N_2497,N_2957);
or U5524 (N_5524,N_2815,N_3253);
nor U5525 (N_5525,N_3857,N_2751);
nor U5526 (N_5526,N_2680,N_3664);
or U5527 (N_5527,N_2045,N_3420);
xor U5528 (N_5528,N_3666,N_2113);
nor U5529 (N_5529,N_3922,N_3411);
nand U5530 (N_5530,N_3280,N_2546);
nand U5531 (N_5531,N_2681,N_3179);
nand U5532 (N_5532,N_2760,N_3284);
or U5533 (N_5533,N_2110,N_2213);
nand U5534 (N_5534,N_2633,N_3293);
nor U5535 (N_5535,N_3577,N_3234);
or U5536 (N_5536,N_2753,N_3048);
nor U5537 (N_5537,N_2241,N_2553);
xnor U5538 (N_5538,N_3613,N_2577);
xnor U5539 (N_5539,N_3077,N_2808);
nor U5540 (N_5540,N_3714,N_3049);
nor U5541 (N_5541,N_3116,N_2773);
or U5542 (N_5542,N_2401,N_3615);
nor U5543 (N_5543,N_2262,N_2738);
nor U5544 (N_5544,N_3917,N_2063);
xor U5545 (N_5545,N_2837,N_2533);
or U5546 (N_5546,N_3883,N_3855);
and U5547 (N_5547,N_2023,N_2925);
or U5548 (N_5548,N_3823,N_3391);
and U5549 (N_5549,N_2989,N_3001);
nand U5550 (N_5550,N_2006,N_3320);
and U5551 (N_5551,N_2689,N_2163);
and U5552 (N_5552,N_2087,N_2546);
and U5553 (N_5553,N_3271,N_3599);
xnor U5554 (N_5554,N_3649,N_3647);
or U5555 (N_5555,N_2266,N_2751);
xnor U5556 (N_5556,N_2450,N_2815);
nor U5557 (N_5557,N_2943,N_3732);
or U5558 (N_5558,N_2174,N_3665);
or U5559 (N_5559,N_2486,N_3332);
nand U5560 (N_5560,N_3135,N_2504);
nand U5561 (N_5561,N_3406,N_3154);
or U5562 (N_5562,N_2690,N_3489);
xor U5563 (N_5563,N_2682,N_3010);
and U5564 (N_5564,N_2631,N_3453);
nor U5565 (N_5565,N_2558,N_3962);
or U5566 (N_5566,N_2432,N_2949);
and U5567 (N_5567,N_3053,N_2689);
nand U5568 (N_5568,N_3431,N_3754);
nand U5569 (N_5569,N_2598,N_3870);
or U5570 (N_5570,N_2111,N_2026);
xnor U5571 (N_5571,N_2906,N_3283);
nand U5572 (N_5572,N_3751,N_2507);
and U5573 (N_5573,N_3340,N_2830);
nor U5574 (N_5574,N_3754,N_2085);
nand U5575 (N_5575,N_3294,N_2216);
nand U5576 (N_5576,N_2149,N_2108);
nand U5577 (N_5577,N_2461,N_2901);
and U5578 (N_5578,N_3102,N_2040);
and U5579 (N_5579,N_3746,N_2909);
or U5580 (N_5580,N_3220,N_3354);
nand U5581 (N_5581,N_2187,N_3950);
or U5582 (N_5582,N_3672,N_2419);
nand U5583 (N_5583,N_2547,N_3525);
nor U5584 (N_5584,N_3245,N_2697);
nand U5585 (N_5585,N_3038,N_2725);
nand U5586 (N_5586,N_3081,N_3966);
or U5587 (N_5587,N_3240,N_3573);
or U5588 (N_5588,N_2221,N_3070);
and U5589 (N_5589,N_3995,N_3548);
nand U5590 (N_5590,N_2170,N_3990);
or U5591 (N_5591,N_3351,N_3476);
nor U5592 (N_5592,N_2023,N_3263);
nand U5593 (N_5593,N_2443,N_3503);
and U5594 (N_5594,N_3861,N_3155);
nor U5595 (N_5595,N_2537,N_3708);
or U5596 (N_5596,N_3016,N_3159);
nand U5597 (N_5597,N_3390,N_3212);
nand U5598 (N_5598,N_3447,N_2758);
xor U5599 (N_5599,N_2018,N_2213);
xnor U5600 (N_5600,N_2720,N_2563);
nand U5601 (N_5601,N_2974,N_2883);
or U5602 (N_5602,N_3172,N_3428);
and U5603 (N_5603,N_2316,N_3872);
nand U5604 (N_5604,N_2353,N_3770);
nand U5605 (N_5605,N_2041,N_3718);
xor U5606 (N_5606,N_3468,N_2414);
nand U5607 (N_5607,N_2378,N_2435);
or U5608 (N_5608,N_3413,N_3952);
and U5609 (N_5609,N_3005,N_2124);
xor U5610 (N_5610,N_3516,N_3464);
and U5611 (N_5611,N_2268,N_2365);
nor U5612 (N_5612,N_2074,N_3460);
and U5613 (N_5613,N_3094,N_2927);
nor U5614 (N_5614,N_3891,N_2942);
or U5615 (N_5615,N_3695,N_3503);
nand U5616 (N_5616,N_2397,N_2458);
or U5617 (N_5617,N_3694,N_3190);
xor U5618 (N_5618,N_2194,N_2462);
nand U5619 (N_5619,N_3576,N_2037);
nor U5620 (N_5620,N_3993,N_3649);
and U5621 (N_5621,N_3131,N_2646);
and U5622 (N_5622,N_3124,N_2405);
xor U5623 (N_5623,N_2245,N_2225);
and U5624 (N_5624,N_2275,N_3315);
or U5625 (N_5625,N_2585,N_2142);
and U5626 (N_5626,N_2546,N_2170);
or U5627 (N_5627,N_3122,N_3651);
nor U5628 (N_5628,N_3546,N_3739);
and U5629 (N_5629,N_2904,N_2648);
xor U5630 (N_5630,N_3546,N_3616);
and U5631 (N_5631,N_3490,N_3395);
and U5632 (N_5632,N_3524,N_3465);
or U5633 (N_5633,N_3583,N_2107);
nor U5634 (N_5634,N_3414,N_3276);
and U5635 (N_5635,N_2576,N_2447);
or U5636 (N_5636,N_3129,N_3509);
nand U5637 (N_5637,N_2476,N_2877);
nor U5638 (N_5638,N_3593,N_3223);
nand U5639 (N_5639,N_3957,N_3135);
nand U5640 (N_5640,N_2477,N_3712);
and U5641 (N_5641,N_2646,N_2145);
nand U5642 (N_5642,N_2818,N_2236);
nor U5643 (N_5643,N_2451,N_2698);
and U5644 (N_5644,N_2675,N_3130);
or U5645 (N_5645,N_2107,N_2045);
nand U5646 (N_5646,N_3968,N_2941);
or U5647 (N_5647,N_2324,N_3679);
nor U5648 (N_5648,N_2785,N_3977);
nor U5649 (N_5649,N_2003,N_3452);
nor U5650 (N_5650,N_2326,N_3893);
nor U5651 (N_5651,N_2341,N_2005);
nor U5652 (N_5652,N_3239,N_3401);
or U5653 (N_5653,N_3029,N_2748);
and U5654 (N_5654,N_2464,N_3095);
or U5655 (N_5655,N_2234,N_3945);
or U5656 (N_5656,N_3163,N_2901);
and U5657 (N_5657,N_3146,N_2993);
nand U5658 (N_5658,N_3485,N_3034);
and U5659 (N_5659,N_2763,N_2281);
or U5660 (N_5660,N_2108,N_3147);
xor U5661 (N_5661,N_2898,N_3824);
or U5662 (N_5662,N_3092,N_3175);
or U5663 (N_5663,N_2569,N_3623);
nor U5664 (N_5664,N_3382,N_2029);
or U5665 (N_5665,N_2810,N_3824);
or U5666 (N_5666,N_3186,N_3102);
or U5667 (N_5667,N_3768,N_3587);
nand U5668 (N_5668,N_3156,N_3796);
or U5669 (N_5669,N_3103,N_2428);
nand U5670 (N_5670,N_2092,N_2133);
and U5671 (N_5671,N_2903,N_2901);
nand U5672 (N_5672,N_3307,N_3280);
nand U5673 (N_5673,N_2644,N_3824);
nand U5674 (N_5674,N_3613,N_3776);
or U5675 (N_5675,N_2049,N_3656);
or U5676 (N_5676,N_3057,N_2184);
or U5677 (N_5677,N_2900,N_3927);
and U5678 (N_5678,N_3944,N_2368);
and U5679 (N_5679,N_2445,N_2973);
nand U5680 (N_5680,N_3588,N_2110);
nor U5681 (N_5681,N_3036,N_3624);
nor U5682 (N_5682,N_3885,N_3757);
or U5683 (N_5683,N_3503,N_3476);
nand U5684 (N_5684,N_3958,N_3408);
nor U5685 (N_5685,N_3170,N_3083);
or U5686 (N_5686,N_2059,N_3039);
and U5687 (N_5687,N_3490,N_3180);
or U5688 (N_5688,N_2592,N_2383);
and U5689 (N_5689,N_2946,N_2071);
or U5690 (N_5690,N_3248,N_3255);
nand U5691 (N_5691,N_2050,N_2497);
nand U5692 (N_5692,N_3192,N_3688);
and U5693 (N_5693,N_2205,N_2754);
or U5694 (N_5694,N_3050,N_3537);
and U5695 (N_5695,N_3801,N_2935);
or U5696 (N_5696,N_2465,N_3680);
nand U5697 (N_5697,N_2231,N_3086);
xor U5698 (N_5698,N_3752,N_3485);
nand U5699 (N_5699,N_2776,N_3073);
and U5700 (N_5700,N_3994,N_2333);
nor U5701 (N_5701,N_3467,N_2515);
and U5702 (N_5702,N_3604,N_2432);
xor U5703 (N_5703,N_2816,N_3464);
nor U5704 (N_5704,N_3863,N_2625);
nor U5705 (N_5705,N_3844,N_2930);
nor U5706 (N_5706,N_3602,N_2563);
or U5707 (N_5707,N_2101,N_3116);
or U5708 (N_5708,N_3613,N_2849);
nor U5709 (N_5709,N_2583,N_3415);
and U5710 (N_5710,N_2139,N_2918);
xor U5711 (N_5711,N_2343,N_2667);
xor U5712 (N_5712,N_3240,N_3166);
nand U5713 (N_5713,N_3370,N_2214);
and U5714 (N_5714,N_2083,N_2437);
or U5715 (N_5715,N_2093,N_2984);
nor U5716 (N_5716,N_2215,N_3612);
xnor U5717 (N_5717,N_3792,N_3074);
nor U5718 (N_5718,N_2007,N_2021);
nand U5719 (N_5719,N_2861,N_2386);
nor U5720 (N_5720,N_3741,N_2575);
and U5721 (N_5721,N_2960,N_3489);
or U5722 (N_5722,N_2316,N_2169);
nand U5723 (N_5723,N_3659,N_2658);
or U5724 (N_5724,N_3281,N_3954);
nor U5725 (N_5725,N_2961,N_2491);
and U5726 (N_5726,N_3460,N_2802);
nand U5727 (N_5727,N_3849,N_3482);
nand U5728 (N_5728,N_3406,N_2095);
and U5729 (N_5729,N_2706,N_2776);
nor U5730 (N_5730,N_3656,N_3247);
or U5731 (N_5731,N_2616,N_3209);
or U5732 (N_5732,N_3542,N_3552);
nand U5733 (N_5733,N_3261,N_2534);
nor U5734 (N_5734,N_2570,N_2714);
nand U5735 (N_5735,N_3331,N_3870);
or U5736 (N_5736,N_2001,N_3251);
or U5737 (N_5737,N_2929,N_3413);
nand U5738 (N_5738,N_3766,N_3853);
nor U5739 (N_5739,N_2042,N_2566);
or U5740 (N_5740,N_2421,N_3405);
and U5741 (N_5741,N_2247,N_3451);
nor U5742 (N_5742,N_3770,N_2775);
nand U5743 (N_5743,N_2343,N_2972);
and U5744 (N_5744,N_2753,N_3384);
nor U5745 (N_5745,N_2300,N_3024);
nand U5746 (N_5746,N_2963,N_2087);
or U5747 (N_5747,N_2539,N_2832);
or U5748 (N_5748,N_3785,N_2204);
or U5749 (N_5749,N_2872,N_3881);
xor U5750 (N_5750,N_2264,N_2390);
nand U5751 (N_5751,N_3060,N_2250);
nor U5752 (N_5752,N_2435,N_2710);
nor U5753 (N_5753,N_3007,N_2625);
and U5754 (N_5754,N_3436,N_2505);
and U5755 (N_5755,N_2835,N_3808);
nor U5756 (N_5756,N_3515,N_2055);
xor U5757 (N_5757,N_3295,N_3838);
nor U5758 (N_5758,N_3578,N_2865);
nand U5759 (N_5759,N_2125,N_2877);
and U5760 (N_5760,N_2303,N_3160);
or U5761 (N_5761,N_3543,N_3608);
nor U5762 (N_5762,N_2876,N_2677);
or U5763 (N_5763,N_2447,N_2894);
nand U5764 (N_5764,N_2576,N_2584);
or U5765 (N_5765,N_3720,N_2751);
or U5766 (N_5766,N_3375,N_2312);
and U5767 (N_5767,N_2537,N_2517);
nand U5768 (N_5768,N_3146,N_3118);
xnor U5769 (N_5769,N_3372,N_3415);
and U5770 (N_5770,N_2251,N_3414);
nand U5771 (N_5771,N_2603,N_3596);
xor U5772 (N_5772,N_3542,N_2996);
nand U5773 (N_5773,N_2121,N_3935);
and U5774 (N_5774,N_3356,N_3884);
or U5775 (N_5775,N_3646,N_3108);
or U5776 (N_5776,N_3625,N_3486);
nand U5777 (N_5777,N_3626,N_2313);
nand U5778 (N_5778,N_3916,N_2914);
or U5779 (N_5779,N_3037,N_3947);
or U5780 (N_5780,N_2130,N_2930);
nand U5781 (N_5781,N_2991,N_2762);
and U5782 (N_5782,N_3770,N_2852);
nand U5783 (N_5783,N_2248,N_2157);
nand U5784 (N_5784,N_3798,N_3953);
nor U5785 (N_5785,N_2476,N_3653);
nand U5786 (N_5786,N_3316,N_2315);
nor U5787 (N_5787,N_3049,N_2247);
or U5788 (N_5788,N_3349,N_2115);
or U5789 (N_5789,N_3839,N_2653);
or U5790 (N_5790,N_2299,N_2643);
or U5791 (N_5791,N_3684,N_3884);
or U5792 (N_5792,N_3029,N_3003);
nor U5793 (N_5793,N_3085,N_2502);
or U5794 (N_5794,N_3003,N_2771);
and U5795 (N_5795,N_3163,N_2625);
nand U5796 (N_5796,N_2370,N_3592);
or U5797 (N_5797,N_2377,N_3591);
and U5798 (N_5798,N_3530,N_3482);
nand U5799 (N_5799,N_3885,N_2459);
or U5800 (N_5800,N_2145,N_3010);
nor U5801 (N_5801,N_3619,N_2252);
nand U5802 (N_5802,N_3021,N_3533);
nand U5803 (N_5803,N_3037,N_2113);
and U5804 (N_5804,N_3918,N_3714);
nor U5805 (N_5805,N_3242,N_3690);
or U5806 (N_5806,N_3484,N_3337);
nor U5807 (N_5807,N_3660,N_2961);
nor U5808 (N_5808,N_2562,N_3885);
and U5809 (N_5809,N_3232,N_3173);
or U5810 (N_5810,N_3022,N_3055);
and U5811 (N_5811,N_2448,N_2422);
nand U5812 (N_5812,N_3548,N_3009);
nand U5813 (N_5813,N_3892,N_3775);
nor U5814 (N_5814,N_3220,N_2997);
nand U5815 (N_5815,N_2383,N_3030);
and U5816 (N_5816,N_3961,N_2158);
and U5817 (N_5817,N_2843,N_2362);
nor U5818 (N_5818,N_2128,N_3448);
or U5819 (N_5819,N_3564,N_3170);
or U5820 (N_5820,N_2405,N_2067);
xor U5821 (N_5821,N_2883,N_2593);
and U5822 (N_5822,N_2994,N_3498);
or U5823 (N_5823,N_3317,N_2945);
or U5824 (N_5824,N_3354,N_3486);
xor U5825 (N_5825,N_2374,N_2110);
or U5826 (N_5826,N_3761,N_3391);
xnor U5827 (N_5827,N_2688,N_2786);
nor U5828 (N_5828,N_3049,N_2049);
nand U5829 (N_5829,N_2059,N_3922);
nand U5830 (N_5830,N_3974,N_2519);
nor U5831 (N_5831,N_2656,N_3621);
xnor U5832 (N_5832,N_2487,N_2172);
or U5833 (N_5833,N_3087,N_2627);
nand U5834 (N_5834,N_2817,N_2481);
or U5835 (N_5835,N_2501,N_3662);
or U5836 (N_5836,N_3348,N_2726);
or U5837 (N_5837,N_3699,N_2088);
and U5838 (N_5838,N_3384,N_3330);
and U5839 (N_5839,N_2338,N_2429);
nor U5840 (N_5840,N_3901,N_2249);
and U5841 (N_5841,N_2121,N_3419);
nor U5842 (N_5842,N_2815,N_2566);
nor U5843 (N_5843,N_2445,N_2071);
nor U5844 (N_5844,N_3546,N_3963);
nand U5845 (N_5845,N_3629,N_3811);
nand U5846 (N_5846,N_2761,N_2580);
and U5847 (N_5847,N_3312,N_3931);
nor U5848 (N_5848,N_3234,N_2659);
nand U5849 (N_5849,N_2207,N_3686);
nor U5850 (N_5850,N_2225,N_3840);
nand U5851 (N_5851,N_2914,N_3880);
nand U5852 (N_5852,N_2069,N_3357);
xnor U5853 (N_5853,N_3026,N_2609);
nand U5854 (N_5854,N_3976,N_3526);
nor U5855 (N_5855,N_3786,N_3079);
xnor U5856 (N_5856,N_2138,N_3400);
nor U5857 (N_5857,N_3954,N_3537);
nor U5858 (N_5858,N_2432,N_2752);
nand U5859 (N_5859,N_3710,N_2060);
and U5860 (N_5860,N_2611,N_3463);
nor U5861 (N_5861,N_3562,N_2168);
nand U5862 (N_5862,N_3611,N_3417);
nor U5863 (N_5863,N_2015,N_3506);
nor U5864 (N_5864,N_3065,N_3816);
or U5865 (N_5865,N_3760,N_3813);
xnor U5866 (N_5866,N_2374,N_3874);
and U5867 (N_5867,N_2591,N_3843);
and U5868 (N_5868,N_2544,N_3979);
xor U5869 (N_5869,N_2124,N_3552);
or U5870 (N_5870,N_2529,N_3105);
or U5871 (N_5871,N_2781,N_2549);
nor U5872 (N_5872,N_3345,N_2200);
nor U5873 (N_5873,N_2189,N_3639);
nor U5874 (N_5874,N_2868,N_3080);
nand U5875 (N_5875,N_3825,N_3308);
or U5876 (N_5876,N_3660,N_3968);
or U5877 (N_5877,N_3608,N_3601);
nor U5878 (N_5878,N_2174,N_3732);
and U5879 (N_5879,N_2883,N_3407);
nand U5880 (N_5880,N_2960,N_2683);
or U5881 (N_5881,N_2566,N_2531);
nand U5882 (N_5882,N_2275,N_2692);
xnor U5883 (N_5883,N_3742,N_3490);
nand U5884 (N_5884,N_2425,N_3795);
and U5885 (N_5885,N_2215,N_2859);
nor U5886 (N_5886,N_3238,N_2431);
nand U5887 (N_5887,N_2939,N_3407);
nor U5888 (N_5888,N_3297,N_2453);
nand U5889 (N_5889,N_2725,N_2100);
nand U5890 (N_5890,N_3542,N_2309);
and U5891 (N_5891,N_3883,N_3448);
and U5892 (N_5892,N_3030,N_3490);
and U5893 (N_5893,N_3518,N_2062);
and U5894 (N_5894,N_3859,N_2869);
nand U5895 (N_5895,N_2935,N_2734);
nor U5896 (N_5896,N_2182,N_2903);
or U5897 (N_5897,N_3935,N_2133);
or U5898 (N_5898,N_2515,N_3128);
or U5899 (N_5899,N_2977,N_3179);
and U5900 (N_5900,N_2941,N_2918);
and U5901 (N_5901,N_2587,N_3613);
nor U5902 (N_5902,N_3133,N_2698);
and U5903 (N_5903,N_3602,N_3504);
nand U5904 (N_5904,N_2172,N_3682);
and U5905 (N_5905,N_2475,N_3742);
nor U5906 (N_5906,N_3416,N_3648);
and U5907 (N_5907,N_2749,N_3166);
and U5908 (N_5908,N_2025,N_3504);
and U5909 (N_5909,N_3971,N_2190);
and U5910 (N_5910,N_3025,N_2847);
nor U5911 (N_5911,N_2894,N_3982);
nand U5912 (N_5912,N_2504,N_3157);
and U5913 (N_5913,N_3010,N_3314);
or U5914 (N_5914,N_3346,N_3849);
or U5915 (N_5915,N_3445,N_3594);
or U5916 (N_5916,N_3175,N_3842);
nor U5917 (N_5917,N_2392,N_2989);
xor U5918 (N_5918,N_2661,N_3775);
or U5919 (N_5919,N_3164,N_3631);
and U5920 (N_5920,N_3877,N_2515);
xor U5921 (N_5921,N_2344,N_3394);
and U5922 (N_5922,N_2169,N_2744);
and U5923 (N_5923,N_2667,N_2214);
and U5924 (N_5924,N_3949,N_3271);
nand U5925 (N_5925,N_3247,N_3104);
or U5926 (N_5926,N_2408,N_3517);
and U5927 (N_5927,N_3858,N_3996);
nor U5928 (N_5928,N_2999,N_2056);
nand U5929 (N_5929,N_3303,N_3506);
or U5930 (N_5930,N_3333,N_3484);
nor U5931 (N_5931,N_3758,N_2432);
nor U5932 (N_5932,N_2056,N_2476);
or U5933 (N_5933,N_2749,N_2316);
nand U5934 (N_5934,N_3185,N_3184);
and U5935 (N_5935,N_2276,N_3758);
nor U5936 (N_5936,N_3089,N_2501);
or U5937 (N_5937,N_3940,N_2700);
xor U5938 (N_5938,N_2202,N_3858);
xor U5939 (N_5939,N_3190,N_3838);
or U5940 (N_5940,N_2207,N_3412);
nand U5941 (N_5941,N_3367,N_3532);
nor U5942 (N_5942,N_3168,N_2994);
nand U5943 (N_5943,N_2996,N_3637);
nor U5944 (N_5944,N_2315,N_3742);
and U5945 (N_5945,N_3404,N_2020);
nand U5946 (N_5946,N_3560,N_2431);
xor U5947 (N_5947,N_2553,N_3520);
nor U5948 (N_5948,N_2297,N_2430);
and U5949 (N_5949,N_3295,N_3817);
nand U5950 (N_5950,N_3839,N_2076);
nor U5951 (N_5951,N_2658,N_3462);
nor U5952 (N_5952,N_3536,N_3215);
nor U5953 (N_5953,N_3401,N_2116);
and U5954 (N_5954,N_3616,N_3910);
nand U5955 (N_5955,N_3428,N_3475);
nand U5956 (N_5956,N_2091,N_3866);
or U5957 (N_5957,N_3906,N_3498);
nor U5958 (N_5958,N_3969,N_2761);
or U5959 (N_5959,N_2387,N_3637);
nand U5960 (N_5960,N_3735,N_3800);
nand U5961 (N_5961,N_3538,N_2822);
nor U5962 (N_5962,N_3744,N_2527);
nor U5963 (N_5963,N_3882,N_3549);
nor U5964 (N_5964,N_2663,N_2100);
nand U5965 (N_5965,N_3903,N_3624);
nor U5966 (N_5966,N_2978,N_3159);
nand U5967 (N_5967,N_2504,N_3545);
or U5968 (N_5968,N_3538,N_3888);
or U5969 (N_5969,N_2256,N_2285);
xnor U5970 (N_5970,N_3540,N_2705);
and U5971 (N_5971,N_2830,N_2401);
or U5972 (N_5972,N_3797,N_2436);
or U5973 (N_5973,N_3362,N_3677);
nand U5974 (N_5974,N_2120,N_2902);
and U5975 (N_5975,N_2138,N_2786);
or U5976 (N_5976,N_3308,N_2444);
nand U5977 (N_5977,N_2314,N_3083);
and U5978 (N_5978,N_2742,N_2469);
nor U5979 (N_5979,N_3146,N_2070);
nor U5980 (N_5980,N_3692,N_3494);
nand U5981 (N_5981,N_2346,N_3595);
nand U5982 (N_5982,N_3128,N_2887);
nor U5983 (N_5983,N_2399,N_3416);
nor U5984 (N_5984,N_2222,N_3084);
and U5985 (N_5985,N_3664,N_2160);
xor U5986 (N_5986,N_2635,N_3895);
nand U5987 (N_5987,N_2332,N_3597);
nand U5988 (N_5988,N_2895,N_2803);
and U5989 (N_5989,N_3838,N_2984);
nand U5990 (N_5990,N_2014,N_3294);
xor U5991 (N_5991,N_3194,N_3721);
nand U5992 (N_5992,N_3746,N_2720);
nor U5993 (N_5993,N_3813,N_3397);
nor U5994 (N_5994,N_3221,N_2939);
nand U5995 (N_5995,N_2150,N_3371);
and U5996 (N_5996,N_2365,N_2834);
nand U5997 (N_5997,N_2348,N_3379);
xnor U5998 (N_5998,N_2274,N_2093);
and U5999 (N_5999,N_3350,N_3184);
and U6000 (N_6000,N_4692,N_4973);
or U6001 (N_6001,N_4102,N_4621);
xor U6002 (N_6002,N_4785,N_4775);
or U6003 (N_6003,N_4222,N_4461);
nor U6004 (N_6004,N_4831,N_5290);
nor U6005 (N_6005,N_4752,N_5280);
nand U6006 (N_6006,N_5439,N_5814);
xnor U6007 (N_6007,N_4818,N_4781);
nand U6008 (N_6008,N_4708,N_5821);
xor U6009 (N_6009,N_5637,N_5760);
or U6010 (N_6010,N_5223,N_4980);
and U6011 (N_6011,N_4177,N_5119);
or U6012 (N_6012,N_4024,N_5277);
or U6013 (N_6013,N_4599,N_4936);
nand U6014 (N_6014,N_5213,N_4852);
and U6015 (N_6015,N_4881,N_4487);
xnor U6016 (N_6016,N_5710,N_5150);
nand U6017 (N_6017,N_5692,N_5998);
and U6018 (N_6018,N_4760,N_4679);
nand U6019 (N_6019,N_5406,N_5047);
and U6020 (N_6020,N_4310,N_4424);
and U6021 (N_6021,N_4464,N_5698);
or U6022 (N_6022,N_4105,N_4815);
and U6023 (N_6023,N_5454,N_4218);
nor U6024 (N_6024,N_5167,N_5105);
and U6025 (N_6025,N_5164,N_4624);
xor U6026 (N_6026,N_4472,N_4788);
nand U6027 (N_6027,N_4646,N_5563);
nor U6028 (N_6028,N_4062,N_5743);
nor U6029 (N_6029,N_5070,N_5524);
nand U6030 (N_6030,N_4003,N_4063);
or U6031 (N_6031,N_4871,N_5324);
and U6032 (N_6032,N_4888,N_5308);
and U6033 (N_6033,N_4299,N_4408);
and U6034 (N_6034,N_4690,N_4608);
nand U6035 (N_6035,N_4638,N_5428);
xnor U6036 (N_6036,N_5441,N_5611);
nand U6037 (N_6037,N_5986,N_5048);
nand U6038 (N_6038,N_5688,N_5538);
or U6039 (N_6039,N_5146,N_5776);
nand U6040 (N_6040,N_5209,N_5615);
nor U6041 (N_6041,N_4449,N_5486);
and U6042 (N_6042,N_4026,N_5915);
or U6043 (N_6043,N_4877,N_4450);
nand U6044 (N_6044,N_5478,N_5786);
and U6045 (N_6045,N_4720,N_5234);
or U6046 (N_6046,N_4071,N_4804);
and U6047 (N_6047,N_5154,N_5497);
nor U6048 (N_6048,N_4987,N_4600);
xor U6049 (N_6049,N_4274,N_5465);
nor U6050 (N_6050,N_4511,N_4578);
and U6051 (N_6051,N_5459,N_4210);
and U6052 (N_6052,N_4830,N_4069);
nand U6053 (N_6053,N_5340,N_4339);
nand U6054 (N_6054,N_4750,N_4158);
nor U6055 (N_6055,N_4746,N_4510);
xor U6056 (N_6056,N_4494,N_5550);
and U6057 (N_6057,N_5176,N_4983);
nand U6058 (N_6058,N_4576,N_4090);
nand U6059 (N_6059,N_4759,N_5616);
nand U6060 (N_6060,N_5542,N_4451);
nor U6061 (N_6061,N_5668,N_5415);
or U6062 (N_6062,N_4168,N_5118);
nand U6063 (N_6063,N_5633,N_4557);
nand U6064 (N_6064,N_4758,N_4525);
and U6065 (N_6065,N_4731,N_4364);
nand U6066 (N_6066,N_5943,N_4550);
nand U6067 (N_6067,N_5457,N_5355);
nand U6068 (N_6068,N_4796,N_4154);
and U6069 (N_6069,N_5212,N_5723);
and U6070 (N_6070,N_5980,N_5206);
nand U6071 (N_6071,N_4944,N_5326);
or U6072 (N_6072,N_4139,N_4734);
nor U6073 (N_6073,N_4659,N_5354);
nand U6074 (N_6074,N_4545,N_4801);
and U6075 (N_6075,N_5867,N_4187);
and U6076 (N_6076,N_4933,N_4379);
or U6077 (N_6077,N_4219,N_5500);
or U6078 (N_6078,N_5064,N_4531);
nor U6079 (N_6079,N_4955,N_5417);
nor U6080 (N_6080,N_5197,N_5282);
and U6081 (N_6081,N_5519,N_4146);
or U6082 (N_6082,N_4671,N_5382);
nand U6083 (N_6083,N_4763,N_5215);
nand U6084 (N_6084,N_4841,N_5475);
nand U6085 (N_6085,N_5818,N_4403);
or U6086 (N_6086,N_5174,N_4940);
nand U6087 (N_6087,N_5046,N_4360);
nand U6088 (N_6088,N_5963,N_5676);
and U6089 (N_6089,N_5796,N_5893);
nand U6090 (N_6090,N_5313,N_4025);
and U6091 (N_6091,N_4225,N_4833);
nand U6092 (N_6092,N_5879,N_4631);
or U6093 (N_6093,N_5485,N_5396);
xor U6094 (N_6094,N_5987,N_4514);
nor U6095 (N_6095,N_4686,N_5896);
xor U6096 (N_6096,N_5014,N_5230);
nor U6097 (N_6097,N_5504,N_4007);
and U6098 (N_6098,N_4911,N_4534);
and U6099 (N_6099,N_5464,N_5139);
nor U6100 (N_6100,N_4967,N_5175);
xor U6101 (N_6101,N_4323,N_5788);
and U6102 (N_6102,N_4335,N_5012);
nand U6103 (N_6103,N_5029,N_5674);
and U6104 (N_6104,N_5067,N_5283);
xnor U6105 (N_6105,N_4918,N_4952);
nand U6106 (N_6106,N_5192,N_4390);
or U6107 (N_6107,N_5799,N_5222);
and U6108 (N_6108,N_4513,N_5721);
and U6109 (N_6109,N_4491,N_5775);
or U6110 (N_6110,N_5286,N_4991);
or U6111 (N_6111,N_5708,N_4280);
and U6112 (N_6112,N_4753,N_5703);
nor U6113 (N_6113,N_5096,N_5138);
nand U6114 (N_6114,N_4418,N_5106);
xnor U6115 (N_6115,N_4048,N_5148);
or U6116 (N_6116,N_5999,N_5009);
and U6117 (N_6117,N_5112,N_4668);
xor U6118 (N_6118,N_5476,N_4421);
and U6119 (N_6119,N_5431,N_5673);
and U6120 (N_6120,N_4727,N_5503);
xor U6121 (N_6121,N_4340,N_4460);
xor U6122 (N_6122,N_4257,N_5489);
or U6123 (N_6123,N_5309,N_5199);
or U6124 (N_6124,N_5375,N_4712);
and U6125 (N_6125,N_4214,N_4713);
nor U6126 (N_6126,N_4295,N_4732);
and U6127 (N_6127,N_5002,N_4142);
nand U6128 (N_6128,N_4145,N_5071);
nor U6129 (N_6129,N_4837,N_4542);
or U6130 (N_6130,N_5907,N_5751);
and U6131 (N_6131,N_4341,N_5380);
nand U6132 (N_6132,N_5813,N_5677);
nor U6133 (N_6133,N_5525,N_4328);
or U6134 (N_6134,N_4838,N_5532);
xor U6135 (N_6135,N_5143,N_5360);
or U6136 (N_6136,N_5044,N_5684);
nor U6137 (N_6137,N_5809,N_4046);
xor U6138 (N_6138,N_4721,N_4194);
or U6139 (N_6139,N_4907,N_5975);
nor U6140 (N_6140,N_4163,N_4296);
or U6141 (N_6141,N_4478,N_4636);
nand U6142 (N_6142,N_5032,N_5017);
nand U6143 (N_6143,N_5667,N_4508);
xnor U6144 (N_6144,N_5471,N_5574);
nor U6145 (N_6145,N_5381,N_4014);
and U6146 (N_6146,N_4902,N_4311);
xnor U6147 (N_6147,N_5491,N_4320);
nand U6148 (N_6148,N_5837,N_4835);
nor U6149 (N_6149,N_4124,N_4604);
and U6150 (N_6150,N_5188,N_4544);
or U6151 (N_6151,N_4172,N_4935);
nand U6152 (N_6152,N_4148,N_4362);
nor U6153 (N_6153,N_5262,N_5801);
nor U6154 (N_6154,N_5742,N_4894);
nor U6155 (N_6155,N_4258,N_5718);
nand U6156 (N_6156,N_4656,N_4221);
xor U6157 (N_6157,N_5707,N_4495);
nand U6158 (N_6158,N_5217,N_5460);
xnor U6159 (N_6159,N_5603,N_4680);
nor U6160 (N_6160,N_4255,N_4052);
and U6161 (N_6161,N_5618,N_5870);
and U6162 (N_6162,N_4794,N_5635);
nor U6163 (N_6163,N_4038,N_5482);
nor U6164 (N_6164,N_5768,N_4467);
nor U6165 (N_6165,N_5091,N_4689);
and U6166 (N_6166,N_5534,N_4614);
nand U6167 (N_6167,N_5652,N_4256);
nor U6168 (N_6168,N_4057,N_5035);
nor U6169 (N_6169,N_4463,N_5462);
or U6170 (N_6170,N_5777,N_5432);
nor U6171 (N_6171,N_5369,N_4343);
or U6172 (N_6172,N_5235,N_5828);
or U6173 (N_6173,N_5614,N_4622);
and U6174 (N_6174,N_5990,N_5502);
or U6175 (N_6175,N_5256,N_4251);
and U6176 (N_6176,N_4675,N_5874);
nand U6177 (N_6177,N_4290,N_4681);
nor U6178 (N_6178,N_4928,N_5292);
nor U6179 (N_6179,N_4620,N_4329);
and U6180 (N_6180,N_5040,N_5229);
or U6181 (N_6181,N_5935,N_5304);
and U6182 (N_6182,N_5254,N_4009);
nor U6183 (N_6183,N_5897,N_4774);
or U6184 (N_6184,N_4874,N_4301);
and U6185 (N_6185,N_5551,N_4365);
nor U6186 (N_6186,N_5808,N_5772);
or U6187 (N_6187,N_4388,N_4363);
or U6188 (N_6188,N_5994,N_5631);
nor U6189 (N_6189,N_4372,N_4591);
xor U6190 (N_6190,N_4593,N_4792);
and U6191 (N_6191,N_4040,N_5820);
or U6192 (N_6192,N_5069,N_5038);
or U6193 (N_6193,N_5345,N_4305);
or U6194 (N_6194,N_4609,N_4131);
nand U6195 (N_6195,N_5509,N_4238);
nor U6196 (N_6196,N_4440,N_5608);
nand U6197 (N_6197,N_5974,N_5658);
and U6198 (N_6198,N_4411,N_4786);
or U6199 (N_6199,N_5545,N_5807);
nor U6200 (N_6200,N_5898,N_5361);
nand U6201 (N_6201,N_5007,N_4227);
nand U6202 (N_6202,N_4828,N_5285);
or U6203 (N_6203,N_5116,N_5425);
and U6204 (N_6204,N_5852,N_4095);
nand U6205 (N_6205,N_5765,N_5448);
and U6206 (N_6206,N_5936,N_4143);
and U6207 (N_6207,N_4699,N_4672);
nand U6208 (N_6208,N_5594,N_4137);
or U6209 (N_6209,N_5013,N_5085);
and U6210 (N_6210,N_5761,N_5356);
nand U6211 (N_6211,N_4824,N_4897);
nor U6212 (N_6212,N_4486,N_5279);
and U6213 (N_6213,N_4387,N_4455);
nand U6214 (N_6214,N_5607,N_5258);
nand U6215 (N_6215,N_5805,N_5930);
and U6216 (N_6216,N_5001,N_4559);
nand U6217 (N_6217,N_5605,N_4917);
or U6218 (N_6218,N_5712,N_5783);
or U6219 (N_6219,N_4027,N_4433);
or U6220 (N_6220,N_5853,N_5988);
or U6221 (N_6221,N_4572,N_4873);
nand U6222 (N_6222,N_5172,N_4442);
nor U6223 (N_6223,N_4673,N_5544);
and U6224 (N_6224,N_4106,N_5626);
xnor U6225 (N_6225,N_5627,N_4755);
and U6226 (N_6226,N_5394,N_4964);
nor U6227 (N_6227,N_4931,N_4651);
nand U6228 (N_6228,N_5245,N_5274);
xnor U6229 (N_6229,N_5317,N_4549);
and U6230 (N_6230,N_5592,N_4068);
nor U6231 (N_6231,N_4524,N_4556);
or U6232 (N_6232,N_5762,N_4189);
nor U6233 (N_6233,N_5622,N_5985);
nor U6234 (N_6234,N_5984,N_4400);
xor U6235 (N_6235,N_5132,N_4884);
or U6236 (N_6236,N_5060,N_4036);
or U6237 (N_6237,N_4919,N_5977);
or U6238 (N_6238,N_5490,N_4470);
xnor U6239 (N_6239,N_4739,N_5477);
xor U6240 (N_6240,N_5310,N_5125);
nor U6241 (N_6241,N_4317,N_4985);
xor U6242 (N_6242,N_5555,N_4822);
nand U6243 (N_6243,N_4506,N_4259);
or U6244 (N_6244,N_4322,N_4780);
nor U6245 (N_6245,N_5077,N_5514);
nor U6246 (N_6246,N_5399,N_5606);
nand U6247 (N_6247,N_5716,N_5833);
and U6248 (N_6248,N_4401,N_4910);
xnor U6249 (N_6249,N_4308,N_4192);
nor U6250 (N_6250,N_5653,N_5543);
or U6251 (N_6251,N_4722,N_5857);
nor U6252 (N_6252,N_5320,N_5421);
or U6253 (N_6253,N_4004,N_4565);
or U6254 (N_6254,N_4862,N_5347);
nand U6255 (N_6255,N_5709,N_4444);
and U6256 (N_6256,N_5691,N_4598);
and U6257 (N_6257,N_4055,N_4112);
and U6258 (N_6258,N_4635,N_4744);
or U6259 (N_6259,N_5034,N_4882);
nor U6260 (N_6260,N_5225,N_4517);
nand U6261 (N_6261,N_5208,N_5409);
nor U6262 (N_6262,N_4733,N_4089);
nor U6263 (N_6263,N_5377,N_5863);
nand U6264 (N_6264,N_4051,N_5925);
or U6265 (N_6265,N_5352,N_5104);
or U6266 (N_6266,N_4784,N_4325);
or U6267 (N_6267,N_4594,N_4080);
and U6268 (N_6268,N_5960,N_5025);
nand U6269 (N_6269,N_5507,N_4235);
or U6270 (N_6270,N_4880,N_5200);
xnor U6271 (N_6271,N_4682,N_4698);
or U6272 (N_6272,N_4596,N_5794);
or U6273 (N_6273,N_5171,N_4246);
nand U6274 (N_6274,N_4954,N_5445);
nor U6275 (N_6275,N_4416,N_5939);
nand U6276 (N_6276,N_5184,N_4767);
and U6277 (N_6277,N_4567,N_4745);
nor U6278 (N_6278,N_4371,N_4962);
or U6279 (N_6279,N_4773,N_4454);
or U6280 (N_6280,N_5388,N_5533);
nor U6281 (N_6281,N_5798,N_4606);
nor U6282 (N_6282,N_5068,N_5926);
nor U6283 (N_6283,N_5889,N_5868);
or U6284 (N_6284,N_4459,N_4707);
nor U6285 (N_6285,N_4414,N_4943);
nand U6286 (N_6286,N_5523,N_5259);
and U6287 (N_6287,N_5881,N_4044);
and U6288 (N_6288,N_5236,N_5321);
nor U6289 (N_6289,N_4382,N_4913);
nor U6290 (N_6290,N_5458,N_4509);
nand U6291 (N_6291,N_4426,N_5110);
and U6292 (N_6292,N_5284,N_4876);
nand U6293 (N_6293,N_4564,N_5900);
nor U6294 (N_6294,N_5797,N_4123);
nor U6295 (N_6295,N_5314,N_5216);
nand U6296 (N_6296,N_5095,N_4021);
and U6297 (N_6297,N_5792,N_4554);
or U6298 (N_6298,N_4735,N_4428);
xnor U6299 (N_6299,N_5549,N_5403);
or U6300 (N_6300,N_5662,N_4061);
nand U6301 (N_6301,N_5528,N_4272);
xor U6302 (N_6302,N_4330,N_5251);
nand U6303 (N_6303,N_4354,N_5186);
nor U6304 (N_6304,N_4005,N_4499);
or U6305 (N_6305,N_5581,N_5480);
or U6306 (N_6306,N_4979,N_4237);
nand U6307 (N_6307,N_4754,N_5090);
or U6308 (N_6308,N_5978,N_4657);
nand U6309 (N_6309,N_5590,N_5553);
nand U6310 (N_6310,N_4547,N_4164);
xnor U6311 (N_6311,N_5329,N_5364);
nor U6312 (N_6312,N_5122,N_4688);
or U6313 (N_6313,N_5263,N_5588);
or U6314 (N_6314,N_4676,N_5938);
nor U6315 (N_6315,N_5782,N_4429);
nor U6316 (N_6316,N_5207,N_5312);
nor U6317 (N_6317,N_5273,N_4017);
nand U6318 (N_6318,N_4167,N_5479);
or U6319 (N_6319,N_4160,N_4856);
nand U6320 (N_6320,N_5335,N_5815);
and U6321 (N_6321,N_5363,N_5949);
xnor U6322 (N_6322,N_4846,N_4015);
nor U6323 (N_6323,N_4705,N_5024);
nor U6324 (N_6324,N_4171,N_5404);
nand U6325 (N_6325,N_4060,N_5149);
and U6326 (N_6326,N_5976,N_5883);
nor U6327 (N_6327,N_4205,N_4002);
and U6328 (N_6328,N_4479,N_4355);
and U6329 (N_6329,N_4976,N_5057);
nand U6330 (N_6330,N_5840,N_4262);
and U6331 (N_6331,N_5089,N_5932);
xnor U6332 (N_6332,N_4798,N_4268);
nand U6333 (N_6333,N_4766,N_5842);
nand U6334 (N_6334,N_5730,N_5447);
nor U6335 (N_6335,N_5851,N_4905);
or U6336 (N_6336,N_5075,N_4224);
nor U6337 (N_6337,N_4729,N_5967);
xor U6338 (N_6338,N_4077,N_4764);
nand U6339 (N_6339,N_4423,N_5401);
or U6340 (N_6340,N_5027,N_4847);
or U6341 (N_6341,N_4503,N_4446);
or U6342 (N_6342,N_4972,N_5166);
or U6343 (N_6343,N_4075,N_4213);
or U6344 (N_6344,N_5028,N_4351);
or U6345 (N_6345,N_5650,N_4445);
nor U6346 (N_6346,N_5934,N_5194);
nor U6347 (N_6347,N_5584,N_5130);
nand U6348 (N_6348,N_5706,N_5580);
xor U6349 (N_6349,N_5501,N_5604);
xor U6350 (N_6350,N_5496,N_4126);
or U6351 (N_6351,N_4946,N_4723);
nor U6352 (N_6352,N_4054,N_5437);
nand U6353 (N_6353,N_4751,N_4253);
nand U6354 (N_6354,N_4903,N_4336);
nor U6355 (N_6355,N_5512,N_4949);
xnor U6356 (N_6356,N_5625,N_4821);
nand U6357 (N_6357,N_4230,N_4169);
nor U6358 (N_6358,N_5714,N_5111);
or U6359 (N_6359,N_5526,N_4728);
nand U6360 (N_6360,N_4776,N_5136);
xor U6361 (N_6361,N_4097,N_5657);
nand U6362 (N_6362,N_4706,N_5056);
nand U6363 (N_6363,N_4399,N_5291);
or U6364 (N_6364,N_5386,N_4197);
nor U6365 (N_6365,N_5656,N_5036);
nor U6366 (N_6366,N_4165,N_4493);
nand U6367 (N_6367,N_4179,N_5892);
and U6368 (N_6368,N_5917,N_4020);
or U6369 (N_6369,N_4816,N_5573);
or U6370 (N_6370,N_5031,N_5233);
and U6371 (N_6371,N_5271,N_4701);
and U6372 (N_6372,N_4033,N_5011);
or U6373 (N_6373,N_4278,N_5747);
and U6374 (N_6374,N_4857,N_4074);
or U6375 (N_6375,N_5331,N_4883);
and U6376 (N_6376,N_5871,N_4181);
and U6377 (N_6377,N_5670,N_5391);
and U6378 (N_6378,N_5785,N_5763);
or U6379 (N_6379,N_5153,N_4997);
nand U6380 (N_6380,N_4050,N_4220);
and U6381 (N_6381,N_5520,N_4358);
nor U6382 (N_6382,N_4867,N_4670);
nor U6383 (N_6383,N_5498,N_5080);
nand U6384 (N_6384,N_4802,N_4412);
nor U6385 (N_6385,N_4432,N_4281);
or U6386 (N_6386,N_4349,N_5373);
xnor U6387 (N_6387,N_5952,N_5882);
nor U6388 (N_6388,N_4836,N_4346);
nor U6389 (N_6389,N_4666,N_5749);
xnor U6390 (N_6390,N_4331,N_5483);
or U6391 (N_6391,N_4231,N_4045);
nor U6392 (N_6392,N_5481,N_5327);
nand U6393 (N_6393,N_5076,N_4629);
nand U6394 (N_6394,N_4085,N_4865);
xor U6395 (N_6395,N_4756,N_4826);
nor U6396 (N_6396,N_5756,N_5643);
nand U6397 (N_6397,N_5365,N_5913);
and U6398 (N_6398,N_4992,N_4497);
and U6399 (N_6399,N_5341,N_5346);
nand U6400 (N_6400,N_4120,N_4647);
nor U6401 (N_6401,N_5244,N_5648);
and U6402 (N_6402,N_4201,N_5073);
nand U6403 (N_6403,N_5738,N_5623);
or U6404 (N_6404,N_5472,N_4208);
and U6405 (N_6405,N_5231,N_4893);
and U6406 (N_6406,N_4583,N_4639);
or U6407 (N_6407,N_5033,N_4695);
nor U6408 (N_6408,N_5145,N_4602);
nand U6409 (N_6409,N_5645,N_5342);
nand U6410 (N_6410,N_4855,N_5996);
xor U6411 (N_6411,N_5536,N_5120);
nand U6412 (N_6412,N_4866,N_4298);
nand U6413 (N_6413,N_5646,N_5433);
nand U6414 (N_6414,N_4327,N_5727);
or U6415 (N_6415,N_5412,N_4239);
nor U6416 (N_6416,N_4284,N_5052);
or U6417 (N_6417,N_5750,N_5152);
xnor U6418 (N_6418,N_4086,N_4191);
or U6419 (N_6419,N_5293,N_4842);
or U6420 (N_6420,N_4162,N_5741);
xor U6421 (N_6421,N_5400,N_5711);
nor U6422 (N_6422,N_5933,N_5795);
nand U6423 (N_6423,N_4155,N_4084);
or U6424 (N_6424,N_4117,N_4561);
nor U6425 (N_6425,N_5944,N_5793);
nor U6426 (N_6426,N_4338,N_5571);
or U6427 (N_6427,N_5300,N_5005);
xor U6428 (N_6428,N_4711,N_5018);
nor U6429 (N_6429,N_4104,N_5701);
or U6430 (N_6430,N_4999,N_5098);
and U6431 (N_6431,N_5950,N_5671);
nand U6432 (N_6432,N_4190,N_4757);
or U6433 (N_6433,N_4013,N_4736);
nor U6434 (N_6434,N_4245,N_5367);
and U6435 (N_6435,N_5844,N_5566);
xnor U6436 (N_6436,N_4114,N_5804);
or U6437 (N_6437,N_4501,N_4070);
xor U6438 (N_6438,N_5374,N_4490);
nand U6439 (N_6439,N_4693,N_4570);
or U6440 (N_6440,N_4378,N_4324);
and U6441 (N_6441,N_5759,N_5189);
nand U6442 (N_6442,N_4996,N_5610);
and U6443 (N_6443,N_5264,N_4587);
and U6444 (N_6444,N_4533,N_4207);
nor U6445 (N_6445,N_5126,N_4648);
xnor U6446 (N_6446,N_5778,N_5318);
or U6447 (N_6447,N_5198,N_4420);
nand U6448 (N_6448,N_4306,N_5461);
nand U6449 (N_6449,N_4006,N_4153);
nor U6450 (N_6450,N_4138,N_4603);
nand U6451 (N_6451,N_5557,N_5983);
nand U6452 (N_6452,N_5856,N_4369);
and U6453 (N_6453,N_5695,N_4717);
nor U6454 (N_6454,N_5886,N_4872);
nor U6455 (N_6455,N_5904,N_4998);
or U6456 (N_6456,N_4481,N_5920);
or U6457 (N_6457,N_5436,N_5736);
or U6458 (N_6458,N_5651,N_5468);
nand U6459 (N_6459,N_4768,N_4209);
and U6460 (N_6460,N_5484,N_5488);
or U6461 (N_6461,N_5659,N_5953);
nor U6462 (N_6462,N_4610,N_5181);
nand U6463 (N_6463,N_4924,N_4252);
nor U6464 (N_6464,N_4617,N_5168);
nand U6465 (N_6465,N_4391,N_4396);
nand U6466 (N_6466,N_4260,N_4537);
nor U6467 (N_6467,N_4129,N_4042);
nand U6468 (N_6468,N_5826,N_4226);
nor U6469 (N_6469,N_4849,N_4034);
or U6470 (N_6470,N_5921,N_4083);
nand U6471 (N_6471,N_5101,N_5784);
and U6472 (N_6472,N_5989,N_4417);
nor U6473 (N_6473,N_4730,N_5587);
nor U6474 (N_6474,N_4615,N_4439);
nand U6475 (N_6475,N_4474,N_4184);
or U6476 (N_6476,N_5929,N_5315);
nor U6477 (N_6477,N_5003,N_4202);
or U6478 (N_6478,N_5855,N_5474);
and U6479 (N_6479,N_4186,N_5687);
nand U6480 (N_6480,N_4392,N_5865);
or U6481 (N_6481,N_5613,N_4568);
nand U6482 (N_6482,N_4366,N_5829);
nand U6483 (N_6483,N_4977,N_5846);
nor U6484 (N_6484,N_4410,N_4318);
nand U6485 (N_6485,N_5252,N_4951);
or U6486 (N_6486,N_4834,N_5713);
nor U6487 (N_6487,N_4500,N_4538);
xor U6488 (N_6488,N_5601,N_5426);
and U6489 (N_6489,N_5914,N_4694);
and U6490 (N_6490,N_4523,N_4916);
nand U6491 (N_6491,N_4580,N_5694);
nand U6492 (N_6492,N_5466,N_5059);
nand U6493 (N_6493,N_5912,N_4627);
and U6494 (N_6494,N_5583,N_5140);
nor U6495 (N_6495,N_4067,N_5850);
nand U6496 (N_6496,N_5732,N_4654);
xnor U6497 (N_6497,N_5169,N_5115);
nor U6498 (N_6498,N_5201,N_4887);
xnor U6499 (N_6499,N_5268,N_4658);
or U6500 (N_6500,N_4397,N_4476);
and U6501 (N_6501,N_4283,N_4637);
or U6502 (N_6502,N_5411,N_5299);
nand U6503 (N_6503,N_4304,N_4546);
and U6504 (N_6504,N_4183,N_4669);
or U6505 (N_6505,N_4718,N_5022);
or U6506 (N_6506,N_4813,N_4458);
nand U6507 (N_6507,N_4619,N_5816);
nor U6508 (N_6508,N_5430,N_4035);
nand U6509 (N_6509,N_4741,N_5596);
and U6510 (N_6510,N_5649,N_4640);
and U6511 (N_6511,N_5243,N_4912);
nor U6512 (N_6512,N_5734,N_5958);
xnor U6513 (N_6513,N_4303,N_4150);
or U6514 (N_6514,N_4661,N_4116);
or U6515 (N_6515,N_4193,N_5379);
nor U6516 (N_6516,N_5773,N_4316);
and U6517 (N_6517,N_5887,N_5281);
nor U6518 (N_6518,N_4103,N_4823);
xnor U6519 (N_6519,N_4447,N_4772);
nor U6520 (N_6520,N_5724,N_4858);
or U6521 (N_6521,N_4832,N_5505);
xor U6522 (N_6522,N_5770,N_4456);
or U6523 (N_6523,N_5961,N_5739);
or U6524 (N_6524,N_5839,N_4969);
nor U6525 (N_6525,N_4477,N_5752);
xor U6526 (N_6526,N_4286,N_4018);
and U6527 (N_6527,N_4496,N_4065);
and U6528 (N_6528,N_4093,N_4267);
nor U6529 (N_6529,N_4203,N_4443);
nor U6530 (N_6530,N_4294,N_5906);
or U6531 (N_6531,N_4927,N_5858);
nand U6532 (N_6532,N_4938,N_4118);
and U6533 (N_6533,N_5924,N_4377);
xor U6534 (N_6534,N_5306,N_4725);
and U6535 (N_6535,N_5141,N_5822);
or U6536 (N_6536,N_4982,N_5416);
or U6537 (N_6537,N_4498,N_4504);
nand U6538 (N_6538,N_4469,N_5419);
xor U6539 (N_6539,N_5636,N_4385);
xnor U6540 (N_6540,N_4829,N_4353);
and U6541 (N_6541,N_4863,N_5540);
nor U6542 (N_6542,N_4770,N_5753);
nor U6543 (N_6543,N_4404,N_4749);
nor U6544 (N_6544,N_5518,N_5812);
nor U6545 (N_6545,N_4240,N_4288);
nand U6546 (N_6546,N_5307,N_4660);
and U6547 (N_6547,N_5726,N_4914);
nor U6548 (N_6548,N_4195,N_4814);
and U6549 (N_6549,N_4645,N_5825);
nand U6550 (N_6550,N_4652,N_4783);
nor U6551 (N_6551,N_4200,N_5050);
and U6552 (N_6552,N_4762,N_5358);
xnor U6553 (N_6553,N_5000,N_4710);
xor U6554 (N_6554,N_4127,N_4709);
or U6555 (N_6555,N_4386,N_5910);
or U6556 (N_6556,N_4769,N_4958);
and U6557 (N_6557,N_4047,N_4532);
nand U6558 (N_6558,N_5848,N_4361);
nand U6559 (N_6559,N_5398,N_5434);
and U6560 (N_6560,N_4072,N_5560);
nor U6561 (N_6561,N_4087,N_5248);
nand U6562 (N_6562,N_5239,N_4277);
xnor U6563 (N_6563,N_4023,N_5418);
or U6564 (N_6564,N_4700,N_5004);
or U6565 (N_6565,N_5384,N_5074);
or U6566 (N_6566,N_5162,N_4223);
or U6567 (N_6567,N_5100,N_5087);
nor U6568 (N_6568,N_4049,N_4348);
or U6569 (N_6569,N_4875,N_4696);
and U6570 (N_6570,N_5578,N_4597);
nor U6571 (N_6571,N_5982,N_5144);
xnor U6572 (N_6572,N_4334,N_4374);
xor U6573 (N_6573,N_5699,N_4276);
or U6574 (N_6574,N_5552,N_4805);
nand U6575 (N_6575,N_5289,N_5927);
and U6576 (N_6576,N_4791,N_5991);
or U6577 (N_6577,N_5187,N_5683);
or U6578 (N_6578,N_5269,N_4765);
nor U6579 (N_6579,N_5303,N_5219);
or U6580 (N_6580,N_4000,N_4878);
xor U6581 (N_6581,N_4552,N_5541);
and U6582 (N_6582,N_5294,N_5026);
nor U6583 (N_6583,N_5227,N_4098);
and U6584 (N_6584,N_5877,N_5302);
nor U6585 (N_6585,N_5966,N_5278);
nand U6586 (N_6586,N_5393,N_5947);
and U6587 (N_6587,N_5655,N_5506);
nand U6588 (N_6588,N_5903,N_5021);
and U6589 (N_6589,N_4409,N_4056);
nand U6590 (N_6590,N_5338,N_4108);
nor U6591 (N_6591,N_4817,N_4683);
nor U6592 (N_6592,N_4585,N_5962);
nor U6593 (N_6593,N_4948,N_5901);
and U6594 (N_6594,N_5564,N_5971);
nand U6595 (N_6595,N_5134,N_4466);
xor U6596 (N_6596,N_4206,N_5895);
xnor U6597 (N_6597,N_5452,N_5769);
xor U6598 (N_6598,N_4144,N_5835);
nor U6599 (N_6599,N_4900,N_4512);
and U6600 (N_6600,N_4437,N_5495);
nand U6601 (N_6601,N_5093,N_5385);
and U6602 (N_6602,N_5053,N_4932);
nand U6603 (N_6603,N_5487,N_4521);
nor U6604 (N_6604,N_4929,N_4844);
nand U6605 (N_6605,N_5218,N_5876);
nor U6606 (N_6606,N_4215,N_5697);
or U6607 (N_6607,N_5371,N_5629);
and U6608 (N_6608,N_4623,N_5348);
nor U6609 (N_6609,N_5582,N_4820);
nand U6610 (N_6610,N_5530,N_4860);
xnor U6611 (N_6611,N_4111,N_5737);
or U6612 (N_6612,N_4465,N_4152);
nand U6613 (N_6613,N_4357,N_4975);
xnor U6614 (N_6614,N_5728,N_4265);
nor U6615 (N_6615,N_5493,N_5873);
and U6616 (N_6616,N_4406,N_5672);
or U6617 (N_6617,N_5276,N_4347);
and U6618 (N_6618,N_5993,N_5602);
nand U6619 (N_6619,N_4122,N_4551);
nand U6620 (N_6620,N_4642,N_4438);
and U6621 (N_6621,N_4321,N_5968);
nor U6622 (N_6622,N_4425,N_4242);
and U6623 (N_6623,N_5665,N_4810);
and U6624 (N_6624,N_4966,N_4119);
nor U6625 (N_6625,N_5275,N_4853);
and U6626 (N_6626,N_5869,N_5124);
xor U6627 (N_6627,N_4182,N_4279);
nor U6628 (N_6628,N_4422,N_5664);
and U6629 (N_6629,N_5539,N_4300);
nor U6630 (N_6630,N_5979,N_5435);
and U6631 (N_6631,N_4984,N_5802);
nor U6632 (N_6632,N_5647,N_5083);
nand U6633 (N_6633,N_5058,N_4058);
or U6634 (N_6634,N_5595,N_4703);
nand U6635 (N_6635,N_5810,N_5499);
and U6636 (N_6636,N_5621,N_4384);
and U6637 (N_6637,N_4275,N_4527);
nor U6638 (N_6638,N_5395,N_5767);
and U6639 (N_6639,N_5827,N_5689);
nand U6640 (N_6640,N_4199,N_4157);
xnor U6641 (N_6641,N_4263,N_4107);
nand U6642 (N_6642,N_4314,N_5715);
and U6643 (N_6643,N_4522,N_5155);
nor U6644 (N_6644,N_5620,N_5948);
and U6645 (N_6645,N_5193,N_5638);
and U6646 (N_6646,N_4502,N_4248);
nand U6647 (N_6647,N_5758,N_4315);
or U6648 (N_6648,N_5681,N_5531);
or U6649 (N_6649,N_4886,N_4665);
nor U6650 (N_6650,N_4861,N_5015);
and U6651 (N_6651,N_4266,N_5861);
nand U6652 (N_6652,N_5598,N_5558);
xnor U6653 (N_6653,N_4309,N_5147);
nor U6654 (N_6654,N_5562,N_5241);
nor U6655 (N_6655,N_5654,N_4678);
nor U6656 (N_6656,N_4247,N_4435);
or U6657 (N_6657,N_5135,N_5088);
nand U6658 (N_6658,N_5177,N_4930);
and U6659 (N_6659,N_5267,N_5287);
or U6660 (N_6660,N_5467,N_4742);
nand U6661 (N_6661,N_4302,N_5817);
or U6662 (N_6662,N_5911,N_5051);
xnor U6663 (N_6663,N_4649,N_5942);
or U6664 (N_6664,N_4848,N_5909);
nand U6665 (N_6665,N_4904,N_5639);
nor U6666 (N_6666,N_5224,N_5295);
or U6667 (N_6667,N_5065,N_4441);
or U6668 (N_6668,N_4475,N_5030);
and U6669 (N_6669,N_4779,N_5232);
nor U6670 (N_6670,N_5663,N_5246);
nand U6671 (N_6671,N_4342,N_4563);
nor U6672 (N_6672,N_4211,N_5450);
nor U6673 (N_6673,N_4628,N_5325);
xnor U6674 (N_6674,N_4462,N_4581);
or U6675 (N_6675,N_4737,N_4241);
nor U6676 (N_6676,N_5204,N_5546);
nand U6677 (N_6677,N_4516,N_4891);
or U6678 (N_6678,N_4413,N_4771);
or U6679 (N_6679,N_5859,N_4039);
or U6680 (N_6680,N_5023,N_5513);
nor U6681 (N_6681,N_4961,N_5781);
and U6682 (N_6682,N_4249,N_5344);
and U6683 (N_6683,N_5729,N_5661);
xnor U6684 (N_6684,N_4555,N_4797);
nor U6685 (N_6685,N_4393,N_5160);
and U6686 (N_6686,N_4541,N_5221);
nand U6687 (N_6687,N_5054,N_4337);
xor U6688 (N_6688,N_4088,N_5641);
or U6689 (N_6689,N_5946,N_5323);
or U6690 (N_6690,N_5353,N_5332);
nand U6691 (N_6691,N_4079,N_5261);
and U6692 (N_6692,N_5806,N_4133);
nor U6693 (N_6693,N_5366,N_4471);
nor U6694 (N_6694,N_4136,N_4250);
and U6695 (N_6695,N_4663,N_4643);
xnor U6696 (N_6696,N_5916,N_5045);
nand U6697 (N_6697,N_4845,N_5954);
nand U6698 (N_6698,N_5066,N_5675);
nor U6699 (N_6699,N_4092,N_4174);
nand U6700 (N_6700,N_5755,N_4799);
or U6701 (N_6701,N_5158,N_4715);
and U6702 (N_6702,N_4008,N_4217);
and U6703 (N_6703,N_4868,N_4626);
and U6704 (N_6704,N_5884,N_5630);
or U6705 (N_6705,N_4198,N_4677);
nand U6706 (N_6706,N_4515,N_5311);
nand U6707 (N_6707,N_5473,N_5109);
nand U6708 (N_6708,N_5780,N_4151);
or U6709 (N_6709,N_5529,N_5748);
nor U6710 (N_6710,N_4332,N_5919);
and U6711 (N_6711,N_4282,N_5569);
or U6712 (N_6712,N_5790,N_4968);
nor U6713 (N_6713,N_4398,N_5191);
and U6714 (N_6714,N_5576,N_5129);
or U6715 (N_6715,N_4584,N_4519);
and U6716 (N_6716,N_5628,N_4970);
and U6717 (N_6717,N_5547,N_5951);
or U6718 (N_6718,N_5238,N_4032);
nor U6719 (N_6719,N_5845,N_4540);
or U6720 (N_6720,N_4028,N_5740);
and U6721 (N_6721,N_5612,N_5362);
nand U6722 (N_6722,N_4380,N_4457);
nor U6723 (N_6723,N_5567,N_4287);
or U6724 (N_6724,N_5572,N_5376);
nor U6725 (N_6725,N_5413,N_5890);
nor U6726 (N_6726,N_5682,N_4633);
and U6727 (N_6727,N_4001,N_4548);
nand U6728 (N_6728,N_5429,N_5800);
or U6729 (N_6729,N_5020,N_4945);
nor U6730 (N_6730,N_4528,N_5764);
nand U6731 (N_6731,N_5255,N_4543);
or U6732 (N_6732,N_5240,N_4261);
and U6733 (N_6733,N_5337,N_5854);
nand U6734 (N_6734,N_5992,N_5832);
and U6735 (N_6735,N_4381,N_4934);
xnor U6736 (N_6736,N_5062,N_4787);
xnor U6737 (N_6737,N_5719,N_5632);
and U6738 (N_6738,N_4234,N_5266);
and U6739 (N_6739,N_4895,N_5872);
or U6740 (N_6740,N_5745,N_5226);
or U6741 (N_6741,N_4589,N_4373);
or U6742 (N_6742,N_5257,N_4839);
nand U6743 (N_6743,N_5669,N_4653);
nand U6744 (N_6744,N_5301,N_5237);
or U6745 (N_6745,N_5619,N_5438);
and U6746 (N_6746,N_4579,N_4031);
or U6747 (N_6747,N_5972,N_4293);
or U6748 (N_6748,N_5908,N_4269);
and U6749 (N_6749,N_4535,N_4960);
nand U6750 (N_6750,N_5843,N_5744);
or U6751 (N_6751,N_5296,N_5754);
nor U6752 (N_6752,N_4704,N_5420);
and U6753 (N_6753,N_4134,N_4577);
or U6754 (N_6754,N_5082,N_4778);
and U6755 (N_6755,N_5679,N_4782);
nor U6756 (N_6756,N_4906,N_4890);
nor U6757 (N_6757,N_4662,N_4161);
nor U6758 (N_6758,N_4612,N_4022);
nor U6759 (N_6759,N_4843,N_4993);
and U6760 (N_6760,N_5789,N_4790);
and U6761 (N_6761,N_5746,N_4947);
and U6762 (N_6762,N_5527,N_4613);
nand U6763 (N_6763,N_4923,N_5956);
nor U6764 (N_6764,N_5092,N_5157);
nor U6765 (N_6765,N_4344,N_5161);
and U6766 (N_6766,N_5774,N_5771);
xor U6767 (N_6767,N_4965,N_4244);
nor U6768 (N_6768,N_5589,N_5617);
or U6769 (N_6769,N_5705,N_5508);
nor U6770 (N_6770,N_5586,N_5179);
xnor U6771 (N_6771,N_4942,N_5019);
nor U6772 (N_6772,N_5862,N_4212);
and U6773 (N_6773,N_5591,N_4402);
or U6774 (N_6774,N_5405,N_4529);
and U6775 (N_6775,N_5137,N_5521);
nand U6776 (N_6776,N_4920,N_4819);
and U6777 (N_6777,N_4452,N_4803);
and U6778 (N_6778,N_4574,N_4175);
nor U6779 (N_6779,N_4530,N_5195);
nand U6780 (N_6780,N_4896,N_4076);
nor U6781 (N_6781,N_4825,N_4655);
nand U6782 (N_6782,N_4959,N_5957);
or U6783 (N_6783,N_4430,N_4053);
xnor U6784 (N_6784,N_5556,N_5173);
nor U6785 (N_6785,N_5378,N_4011);
nand U6786 (N_6786,N_4562,N_5880);
nand U6787 (N_6787,N_4395,N_4702);
and U6788 (N_6788,N_5453,N_5593);
and U6789 (N_6789,N_4073,N_5841);
and U6790 (N_6790,N_5336,N_5725);
and U6791 (N_6791,N_4204,N_4125);
nand U6792 (N_6792,N_5559,N_5733);
nor U6793 (N_6793,N_5039,N_5178);
and U6794 (N_6794,N_4569,N_5128);
nand U6795 (N_6795,N_4808,N_5372);
or U6796 (N_6796,N_5108,N_5931);
nand U6797 (N_6797,N_5228,N_4536);
and U6798 (N_6798,N_4870,N_5196);
nor U6799 (N_6799,N_4128,N_4064);
xor U6800 (N_6800,N_4939,N_4611);
nor U6801 (N_6801,N_4854,N_4526);
and U6802 (N_6802,N_5940,N_4473);
and U6803 (N_6803,N_5443,N_5702);
and U6804 (N_6804,N_5402,N_5242);
nand U6805 (N_6805,N_5392,N_4312);
or U6806 (N_6806,N_4812,N_5265);
or U6807 (N_6807,N_4030,N_5634);
or U6808 (N_6808,N_4571,N_4687);
nand U6809 (N_6809,N_5316,N_5247);
nor U6810 (N_6810,N_5370,N_4010);
xnor U6811 (N_6811,N_4505,N_5010);
nor U6812 (N_6812,N_4096,N_4586);
and U6813 (N_6813,N_4178,N_5410);
or U6814 (N_6814,N_5599,N_5390);
nor U6815 (N_6815,N_4356,N_4156);
and U6816 (N_6816,N_5114,N_5678);
or U6817 (N_6817,N_5511,N_5693);
or U6818 (N_6818,N_4507,N_4313);
nor U6819 (N_6819,N_4394,N_5298);
and U6820 (N_6820,N_5981,N_4921);
xor U6821 (N_6821,N_5644,N_5343);
or U6822 (N_6822,N_4885,N_5959);
nor U6823 (N_6823,N_4407,N_4141);
nand U6824 (N_6824,N_5600,N_5440);
or U6825 (N_6825,N_4431,N_4480);
and U6826 (N_6826,N_4468,N_4099);
nand U6827 (N_6827,N_5535,N_5554);
nor U6828 (N_6828,N_4216,N_4898);
xnor U6829 (N_6829,N_5055,N_4807);
nor U6830 (N_6830,N_5834,N_4685);
nor U6831 (N_6831,N_5609,N_5170);
or U6832 (N_6832,N_4484,N_4101);
or U6833 (N_6833,N_4777,N_5270);
and U6834 (N_6834,N_5891,N_5455);
and U6835 (N_6835,N_4029,N_4909);
nand U6836 (N_6836,N_5214,N_5334);
nor U6837 (N_6837,N_4869,N_4616);
or U6838 (N_6838,N_4297,N_4560);
or U6839 (N_6839,N_5185,N_4345);
and U6840 (N_6840,N_4100,N_4436);
or U6841 (N_6841,N_5642,N_4595);
or U6842 (N_6842,N_5250,N_4482);
or U6843 (N_6843,N_5819,N_4974);
and U6844 (N_6844,N_5875,N_5333);
nor U6845 (N_6845,N_4605,N_4684);
and U6846 (N_6846,N_4795,N_5941);
nand U6847 (N_6847,N_5685,N_5078);
xor U6848 (N_6848,N_4448,N_5690);
nor U6849 (N_6849,N_5061,N_4434);
and U6850 (N_6850,N_5937,N_5322);
and U6851 (N_6851,N_5575,N_4389);
xnor U6852 (N_6852,N_5383,N_4809);
or U6853 (N_6853,N_4634,N_5803);
or U6854 (N_6854,N_4566,N_5585);
nand U6855 (N_6855,N_4851,N_5717);
nand U6856 (N_6856,N_5902,N_5203);
and U6857 (N_6857,N_4520,N_5463);
nor U6858 (N_6858,N_4691,N_4582);
and U6859 (N_6859,N_5253,N_5183);
or U6860 (N_6860,N_4188,N_5042);
or U6861 (N_6861,N_5423,N_5494);
or U6862 (N_6862,N_5894,N_5123);
nor U6863 (N_6863,N_4243,N_5131);
and U6864 (N_6864,N_5117,N_5964);
or U6865 (N_6865,N_4950,N_5107);
or U6866 (N_6866,N_4453,N_4081);
nor U6867 (N_6867,N_4254,N_5446);
nor U6868 (N_6868,N_5757,N_4196);
and U6869 (N_6869,N_4724,N_4415);
nor U6870 (N_6870,N_4740,N_4630);
and U6871 (N_6871,N_4850,N_5451);
nor U6872 (N_6872,N_4738,N_5885);
or U6873 (N_6873,N_4588,N_4273);
nand U6874 (N_6874,N_5305,N_5151);
nor U6875 (N_6875,N_4915,N_5389);
nor U6876 (N_6876,N_5522,N_5923);
nor U6877 (N_6877,N_5368,N_5099);
nor U6878 (N_6878,N_5680,N_4326);
xnor U6879 (N_6879,N_5079,N_5696);
and U6880 (N_6880,N_4019,N_4995);
nand U6881 (N_6881,N_5735,N_4370);
nor U6882 (N_6882,N_5387,N_5811);
and U6883 (N_6883,N_4925,N_5260);
and U6884 (N_6884,N_4664,N_5142);
and U6885 (N_6885,N_4644,N_5577);
xnor U6886 (N_6886,N_4285,N_4059);
or U6887 (N_6887,N_5444,N_5163);
and U6888 (N_6888,N_5469,N_5548);
and U6889 (N_6889,N_4228,N_4988);
nor U6890 (N_6890,N_4233,N_4132);
and U6891 (N_6891,N_5704,N_5202);
or U6892 (N_6892,N_4185,N_4989);
nor U6893 (N_6893,N_5165,N_5133);
and U6894 (N_6894,N_4159,N_4289);
and U6895 (N_6895,N_5288,N_5830);
or U6896 (N_6896,N_4697,N_4899);
xor U6897 (N_6897,N_4864,N_5973);
nor U6898 (N_6898,N_4264,N_4016);
or U6899 (N_6899,N_5249,N_4978);
nor U6900 (N_6900,N_5836,N_4590);
xor U6901 (N_6901,N_5359,N_4789);
nor U6902 (N_6902,N_5182,N_4082);
nor U6903 (N_6903,N_4483,N_4292);
nor U6904 (N_6904,N_4492,N_4518);
nand U6905 (N_6905,N_4650,N_4922);
and U6906 (N_6906,N_4376,N_4859);
nor U6907 (N_6907,N_4990,N_5849);
and U6908 (N_6908,N_5510,N_5686);
nand U6909 (N_6909,N_4641,N_5449);
nor U6910 (N_6910,N_5397,N_5492);
nor U6911 (N_6911,N_5103,N_4840);
nor U6912 (N_6912,N_4575,N_4173);
nor U6913 (N_6913,N_4043,N_5081);
nor U6914 (N_6914,N_4236,N_4714);
xor U6915 (N_6915,N_5722,N_5905);
nor U6916 (N_6916,N_5847,N_5720);
and U6917 (N_6917,N_4012,N_5121);
xnor U6918 (N_6918,N_4037,N_4066);
or U6919 (N_6919,N_5350,N_4180);
or U6920 (N_6920,N_5995,N_5211);
nand U6921 (N_6921,N_4553,N_5407);
nor U6922 (N_6922,N_5700,N_5330);
or U6923 (N_6923,N_4375,N_5955);
xor U6924 (N_6924,N_4170,N_4941);
or U6925 (N_6925,N_5470,N_5180);
or U6926 (N_6926,N_5823,N_4091);
or U6927 (N_6927,N_4926,N_5190);
nand U6928 (N_6928,N_4761,N_5220);
nand U6929 (N_6929,N_4994,N_5094);
or U6930 (N_6930,N_5408,N_5970);
nand U6931 (N_6931,N_5888,N_4889);
and U6932 (N_6932,N_5640,N_4908);
or U6933 (N_6933,N_5666,N_4485);
nand U6934 (N_6934,N_5339,N_4405);
nand U6935 (N_6935,N_4726,N_4953);
and U6936 (N_6936,N_5016,N_4957);
nor U6937 (N_6937,N_5561,N_4719);
or U6938 (N_6938,N_4140,N_5965);
or U6939 (N_6939,N_5624,N_5899);
nor U6940 (N_6940,N_4121,N_4110);
nor U6941 (N_6941,N_5831,N_5041);
and U6942 (N_6942,N_5787,N_5210);
and U6943 (N_6943,N_4419,N_4539);
nand U6944 (N_6944,N_5766,N_4094);
or U6945 (N_6945,N_5427,N_4800);
nor U6946 (N_6946,N_4319,N_4618);
nor U6947 (N_6947,N_5072,N_5866);
nor U6948 (N_6948,N_4901,N_5049);
and U6949 (N_6949,N_5037,N_5864);
or U6950 (N_6950,N_5928,N_4359);
nand U6951 (N_6951,N_4963,N_5517);
nand U6952 (N_6952,N_4176,N_4149);
and U6953 (N_6953,N_5779,N_4981);
or U6954 (N_6954,N_5006,N_5918);
xor U6955 (N_6955,N_5456,N_5860);
and U6956 (N_6956,N_4793,N_5424);
nor U6957 (N_6957,N_5731,N_4748);
nand U6958 (N_6958,N_5414,N_4307);
xor U6959 (N_6959,N_5945,N_4352);
xor U6960 (N_6960,N_4333,N_5127);
and U6961 (N_6961,N_4113,N_4607);
nand U6962 (N_6962,N_4573,N_5008);
or U6963 (N_6963,N_5328,N_5922);
nand U6964 (N_6964,N_5084,N_5097);
and U6965 (N_6965,N_4427,N_4489);
or U6966 (N_6966,N_4806,N_4350);
nand U6967 (N_6967,N_4625,N_4747);
nor U6968 (N_6968,N_5205,N_4632);
and U6969 (N_6969,N_4270,N_5319);
nand U6970 (N_6970,N_4271,N_4601);
or U6971 (N_6971,N_4956,N_4130);
nand U6972 (N_6972,N_5102,N_4667);
xnor U6973 (N_6973,N_5878,N_4367);
or U6974 (N_6974,N_5156,N_4674);
xnor U6975 (N_6975,N_4879,N_5086);
and U6976 (N_6976,N_4488,N_5997);
nor U6977 (N_6977,N_4147,N_4971);
nor U6978 (N_6978,N_4558,N_5824);
and U6979 (N_6979,N_4892,N_5565);
nand U6980 (N_6980,N_5297,N_5043);
or U6981 (N_6981,N_4811,N_4109);
nor U6982 (N_6982,N_5272,N_5515);
or U6983 (N_6983,N_5579,N_5357);
nand U6984 (N_6984,N_4368,N_4229);
or U6985 (N_6985,N_5660,N_5568);
and U6986 (N_6986,N_5422,N_5113);
nor U6987 (N_6987,N_5159,N_5597);
xnor U6988 (N_6988,N_4986,N_4115);
nand U6989 (N_6989,N_5838,N_4291);
nand U6990 (N_6990,N_5351,N_4827);
nand U6991 (N_6991,N_4592,N_5791);
and U6992 (N_6992,N_5516,N_4041);
nand U6993 (N_6993,N_5537,N_4716);
nor U6994 (N_6994,N_4166,N_4383);
xor U6995 (N_6995,N_5570,N_5969);
xnor U6996 (N_6996,N_4232,N_5349);
xor U6997 (N_6997,N_5442,N_5063);
or U6998 (N_6998,N_4078,N_4937);
and U6999 (N_6999,N_4743,N_4135);
xnor U7000 (N_7000,N_5597,N_5886);
and U7001 (N_7001,N_5769,N_5587);
nor U7002 (N_7002,N_4137,N_4830);
nand U7003 (N_7003,N_4442,N_5938);
or U7004 (N_7004,N_5171,N_4469);
nand U7005 (N_7005,N_4361,N_5008);
nand U7006 (N_7006,N_4329,N_4837);
nand U7007 (N_7007,N_5223,N_5259);
nand U7008 (N_7008,N_5032,N_5040);
or U7009 (N_7009,N_4492,N_5906);
nor U7010 (N_7010,N_5695,N_4041);
and U7011 (N_7011,N_4558,N_4868);
or U7012 (N_7012,N_5286,N_4198);
and U7013 (N_7013,N_4687,N_5525);
or U7014 (N_7014,N_5089,N_5496);
and U7015 (N_7015,N_4218,N_5001);
or U7016 (N_7016,N_5054,N_4687);
or U7017 (N_7017,N_4203,N_5765);
nand U7018 (N_7018,N_5076,N_5521);
nor U7019 (N_7019,N_4824,N_4541);
nor U7020 (N_7020,N_4319,N_5142);
and U7021 (N_7021,N_4338,N_5623);
or U7022 (N_7022,N_5506,N_4103);
and U7023 (N_7023,N_5967,N_5219);
nand U7024 (N_7024,N_5073,N_5730);
and U7025 (N_7025,N_4626,N_4960);
and U7026 (N_7026,N_4472,N_4851);
and U7027 (N_7027,N_5400,N_4565);
xnor U7028 (N_7028,N_5263,N_5039);
or U7029 (N_7029,N_4276,N_4850);
nor U7030 (N_7030,N_4392,N_4944);
nand U7031 (N_7031,N_4577,N_4014);
nand U7032 (N_7032,N_5792,N_5953);
and U7033 (N_7033,N_5280,N_4351);
nor U7034 (N_7034,N_5915,N_5579);
or U7035 (N_7035,N_5625,N_5831);
nor U7036 (N_7036,N_4174,N_5496);
or U7037 (N_7037,N_4885,N_5251);
nand U7038 (N_7038,N_5858,N_5012);
xnor U7039 (N_7039,N_4607,N_5172);
xor U7040 (N_7040,N_5873,N_5249);
and U7041 (N_7041,N_4722,N_5829);
or U7042 (N_7042,N_4064,N_5140);
or U7043 (N_7043,N_5083,N_5033);
nand U7044 (N_7044,N_4202,N_4411);
xor U7045 (N_7045,N_4953,N_4712);
and U7046 (N_7046,N_5769,N_5131);
and U7047 (N_7047,N_5677,N_5434);
and U7048 (N_7048,N_5428,N_5908);
nand U7049 (N_7049,N_4459,N_4065);
or U7050 (N_7050,N_4939,N_5897);
nor U7051 (N_7051,N_5101,N_5218);
nand U7052 (N_7052,N_4033,N_4525);
or U7053 (N_7053,N_4026,N_5373);
nor U7054 (N_7054,N_5890,N_4052);
and U7055 (N_7055,N_4627,N_4609);
or U7056 (N_7056,N_4671,N_4878);
and U7057 (N_7057,N_4660,N_5076);
or U7058 (N_7058,N_4441,N_4984);
or U7059 (N_7059,N_5002,N_5448);
and U7060 (N_7060,N_4528,N_5345);
xor U7061 (N_7061,N_4378,N_5932);
xor U7062 (N_7062,N_4597,N_5534);
and U7063 (N_7063,N_4126,N_5156);
nand U7064 (N_7064,N_5196,N_4032);
nor U7065 (N_7065,N_4804,N_4777);
nand U7066 (N_7066,N_5478,N_4046);
nor U7067 (N_7067,N_4003,N_4603);
and U7068 (N_7068,N_4402,N_4508);
nand U7069 (N_7069,N_4211,N_4006);
nor U7070 (N_7070,N_5458,N_5171);
nand U7071 (N_7071,N_5954,N_4706);
nor U7072 (N_7072,N_5092,N_5623);
or U7073 (N_7073,N_4671,N_4928);
nor U7074 (N_7074,N_5035,N_5688);
nand U7075 (N_7075,N_4142,N_4243);
nand U7076 (N_7076,N_5878,N_4238);
xnor U7077 (N_7077,N_5301,N_5273);
xor U7078 (N_7078,N_5916,N_5618);
nand U7079 (N_7079,N_5852,N_4466);
and U7080 (N_7080,N_4714,N_5688);
xor U7081 (N_7081,N_4617,N_4889);
or U7082 (N_7082,N_5444,N_5286);
nor U7083 (N_7083,N_5710,N_4319);
and U7084 (N_7084,N_5284,N_4456);
or U7085 (N_7085,N_5066,N_5038);
nor U7086 (N_7086,N_5680,N_5234);
and U7087 (N_7087,N_4801,N_5266);
nor U7088 (N_7088,N_5566,N_4150);
nand U7089 (N_7089,N_4621,N_5138);
nor U7090 (N_7090,N_5836,N_5261);
or U7091 (N_7091,N_4168,N_5049);
or U7092 (N_7092,N_4376,N_5076);
nand U7093 (N_7093,N_4281,N_4418);
nand U7094 (N_7094,N_4568,N_5001);
nor U7095 (N_7095,N_4754,N_5248);
nor U7096 (N_7096,N_4601,N_5479);
nor U7097 (N_7097,N_4918,N_5384);
nor U7098 (N_7098,N_5920,N_5963);
or U7099 (N_7099,N_4608,N_5023);
nand U7100 (N_7100,N_5100,N_4424);
nor U7101 (N_7101,N_5458,N_5497);
and U7102 (N_7102,N_4156,N_4146);
nand U7103 (N_7103,N_5638,N_4670);
nand U7104 (N_7104,N_4598,N_5689);
nor U7105 (N_7105,N_5551,N_5804);
nand U7106 (N_7106,N_4568,N_4273);
and U7107 (N_7107,N_4185,N_4625);
nand U7108 (N_7108,N_5247,N_4681);
nand U7109 (N_7109,N_5634,N_5417);
and U7110 (N_7110,N_4677,N_4361);
and U7111 (N_7111,N_5313,N_5338);
xnor U7112 (N_7112,N_5441,N_4787);
nand U7113 (N_7113,N_4721,N_5074);
xnor U7114 (N_7114,N_4127,N_4115);
nor U7115 (N_7115,N_5237,N_4100);
nor U7116 (N_7116,N_4086,N_5374);
nor U7117 (N_7117,N_5006,N_5158);
or U7118 (N_7118,N_5318,N_5103);
and U7119 (N_7119,N_4801,N_4852);
or U7120 (N_7120,N_4837,N_4973);
or U7121 (N_7121,N_4835,N_5714);
or U7122 (N_7122,N_5413,N_5338);
nand U7123 (N_7123,N_4710,N_5705);
nor U7124 (N_7124,N_5812,N_4085);
nor U7125 (N_7125,N_5639,N_4190);
xnor U7126 (N_7126,N_4809,N_4137);
and U7127 (N_7127,N_5177,N_4376);
and U7128 (N_7128,N_5883,N_5927);
nor U7129 (N_7129,N_5937,N_4747);
nor U7130 (N_7130,N_5956,N_4442);
nor U7131 (N_7131,N_5148,N_5843);
nand U7132 (N_7132,N_4331,N_4811);
nor U7133 (N_7133,N_4044,N_5052);
nand U7134 (N_7134,N_5341,N_4769);
xor U7135 (N_7135,N_5373,N_5672);
nor U7136 (N_7136,N_4771,N_5491);
nor U7137 (N_7137,N_4067,N_4834);
nor U7138 (N_7138,N_5161,N_5605);
nor U7139 (N_7139,N_4233,N_4942);
nor U7140 (N_7140,N_5569,N_5679);
and U7141 (N_7141,N_4754,N_5946);
nor U7142 (N_7142,N_4174,N_4984);
and U7143 (N_7143,N_4216,N_5950);
nor U7144 (N_7144,N_4146,N_5346);
nand U7145 (N_7145,N_4265,N_5088);
or U7146 (N_7146,N_4001,N_4135);
nand U7147 (N_7147,N_5754,N_4012);
and U7148 (N_7148,N_4512,N_5519);
nand U7149 (N_7149,N_5828,N_4189);
and U7150 (N_7150,N_5819,N_5769);
and U7151 (N_7151,N_4747,N_5430);
and U7152 (N_7152,N_4224,N_5814);
and U7153 (N_7153,N_5637,N_5733);
nor U7154 (N_7154,N_5580,N_5337);
nand U7155 (N_7155,N_4241,N_5865);
and U7156 (N_7156,N_5022,N_4901);
nor U7157 (N_7157,N_5383,N_5621);
xor U7158 (N_7158,N_5049,N_4362);
nand U7159 (N_7159,N_4534,N_5725);
nor U7160 (N_7160,N_5233,N_5425);
xor U7161 (N_7161,N_4164,N_5121);
or U7162 (N_7162,N_4904,N_4021);
nand U7163 (N_7163,N_4273,N_5670);
and U7164 (N_7164,N_4458,N_5741);
or U7165 (N_7165,N_4462,N_5008);
nand U7166 (N_7166,N_4690,N_5630);
nor U7167 (N_7167,N_4085,N_5429);
nor U7168 (N_7168,N_5292,N_4002);
or U7169 (N_7169,N_4006,N_5650);
and U7170 (N_7170,N_4497,N_4713);
or U7171 (N_7171,N_4401,N_5302);
nand U7172 (N_7172,N_4438,N_5572);
nand U7173 (N_7173,N_4292,N_4861);
and U7174 (N_7174,N_4762,N_4791);
and U7175 (N_7175,N_5026,N_5447);
nand U7176 (N_7176,N_4401,N_4537);
or U7177 (N_7177,N_4340,N_5666);
or U7178 (N_7178,N_4460,N_4318);
nand U7179 (N_7179,N_4108,N_4622);
nor U7180 (N_7180,N_4939,N_5245);
nor U7181 (N_7181,N_5570,N_4033);
nand U7182 (N_7182,N_4977,N_5128);
nor U7183 (N_7183,N_5965,N_5064);
or U7184 (N_7184,N_5796,N_5064);
or U7185 (N_7185,N_4478,N_5525);
nor U7186 (N_7186,N_5392,N_5076);
or U7187 (N_7187,N_4863,N_4064);
and U7188 (N_7188,N_5685,N_5671);
nor U7189 (N_7189,N_5503,N_5826);
nor U7190 (N_7190,N_5646,N_4304);
xnor U7191 (N_7191,N_5842,N_4614);
or U7192 (N_7192,N_4370,N_5936);
nand U7193 (N_7193,N_4319,N_4304);
nor U7194 (N_7194,N_5450,N_4429);
or U7195 (N_7195,N_4364,N_4352);
or U7196 (N_7196,N_4490,N_5689);
nor U7197 (N_7197,N_5162,N_5247);
nor U7198 (N_7198,N_4855,N_4633);
xor U7199 (N_7199,N_4092,N_5458);
and U7200 (N_7200,N_5258,N_5370);
nor U7201 (N_7201,N_4868,N_5951);
nor U7202 (N_7202,N_5080,N_4373);
and U7203 (N_7203,N_4030,N_5549);
and U7204 (N_7204,N_5301,N_4180);
nor U7205 (N_7205,N_5513,N_4633);
or U7206 (N_7206,N_4764,N_4891);
nor U7207 (N_7207,N_4276,N_4427);
nor U7208 (N_7208,N_5976,N_4657);
nor U7209 (N_7209,N_5190,N_4985);
xnor U7210 (N_7210,N_5447,N_4863);
nand U7211 (N_7211,N_4153,N_5171);
nor U7212 (N_7212,N_4071,N_5636);
or U7213 (N_7213,N_4782,N_4943);
and U7214 (N_7214,N_4032,N_4899);
or U7215 (N_7215,N_5621,N_4561);
and U7216 (N_7216,N_5952,N_4052);
nor U7217 (N_7217,N_4921,N_5305);
xor U7218 (N_7218,N_5454,N_5452);
and U7219 (N_7219,N_5489,N_4370);
nor U7220 (N_7220,N_4713,N_4597);
nor U7221 (N_7221,N_5479,N_5890);
nand U7222 (N_7222,N_4408,N_4861);
and U7223 (N_7223,N_4435,N_4510);
and U7224 (N_7224,N_4616,N_4993);
and U7225 (N_7225,N_5952,N_4324);
nand U7226 (N_7226,N_4975,N_5934);
nor U7227 (N_7227,N_5394,N_5947);
nand U7228 (N_7228,N_5928,N_5861);
nor U7229 (N_7229,N_4078,N_4322);
nand U7230 (N_7230,N_5318,N_5581);
nand U7231 (N_7231,N_4528,N_4478);
or U7232 (N_7232,N_5909,N_5772);
and U7233 (N_7233,N_4554,N_5044);
or U7234 (N_7234,N_5783,N_5354);
nand U7235 (N_7235,N_5461,N_5878);
nand U7236 (N_7236,N_4852,N_5987);
and U7237 (N_7237,N_4228,N_5515);
and U7238 (N_7238,N_5664,N_4250);
or U7239 (N_7239,N_4740,N_5588);
nor U7240 (N_7240,N_5523,N_4641);
and U7241 (N_7241,N_4292,N_5286);
and U7242 (N_7242,N_4329,N_4407);
and U7243 (N_7243,N_4627,N_5864);
and U7244 (N_7244,N_5475,N_4308);
nand U7245 (N_7245,N_4305,N_4277);
and U7246 (N_7246,N_4124,N_4378);
or U7247 (N_7247,N_4931,N_5198);
or U7248 (N_7248,N_4625,N_5236);
and U7249 (N_7249,N_5139,N_5495);
nand U7250 (N_7250,N_4587,N_4728);
nand U7251 (N_7251,N_5696,N_5083);
or U7252 (N_7252,N_4610,N_5355);
nor U7253 (N_7253,N_4823,N_5369);
or U7254 (N_7254,N_4183,N_4493);
nand U7255 (N_7255,N_5081,N_5401);
nor U7256 (N_7256,N_5367,N_4165);
and U7257 (N_7257,N_4735,N_5513);
xor U7258 (N_7258,N_4622,N_4506);
xor U7259 (N_7259,N_5032,N_4036);
nor U7260 (N_7260,N_5483,N_5563);
xnor U7261 (N_7261,N_5371,N_4249);
xor U7262 (N_7262,N_5743,N_4760);
and U7263 (N_7263,N_5306,N_4803);
nand U7264 (N_7264,N_4238,N_5070);
nor U7265 (N_7265,N_5604,N_5542);
nor U7266 (N_7266,N_5565,N_4351);
nand U7267 (N_7267,N_5136,N_4811);
and U7268 (N_7268,N_5781,N_5947);
or U7269 (N_7269,N_4162,N_4424);
or U7270 (N_7270,N_5821,N_4392);
and U7271 (N_7271,N_4300,N_5674);
nand U7272 (N_7272,N_5979,N_5260);
and U7273 (N_7273,N_5786,N_4322);
nand U7274 (N_7274,N_4104,N_4355);
nand U7275 (N_7275,N_4886,N_5871);
and U7276 (N_7276,N_5374,N_4733);
or U7277 (N_7277,N_5556,N_4562);
nand U7278 (N_7278,N_4241,N_4693);
and U7279 (N_7279,N_5382,N_4182);
or U7280 (N_7280,N_5960,N_5556);
and U7281 (N_7281,N_4517,N_4532);
nor U7282 (N_7282,N_5563,N_4552);
nand U7283 (N_7283,N_5195,N_5172);
and U7284 (N_7284,N_4244,N_4889);
nand U7285 (N_7285,N_4821,N_5314);
nand U7286 (N_7286,N_5730,N_5801);
xnor U7287 (N_7287,N_4765,N_4618);
xor U7288 (N_7288,N_5282,N_5638);
or U7289 (N_7289,N_5766,N_4945);
or U7290 (N_7290,N_4179,N_4654);
nand U7291 (N_7291,N_5755,N_4285);
or U7292 (N_7292,N_5878,N_5339);
nor U7293 (N_7293,N_5547,N_4175);
and U7294 (N_7294,N_4149,N_5949);
and U7295 (N_7295,N_4488,N_4811);
nor U7296 (N_7296,N_5842,N_5228);
xnor U7297 (N_7297,N_4212,N_4470);
xnor U7298 (N_7298,N_5392,N_5120);
or U7299 (N_7299,N_4098,N_4174);
and U7300 (N_7300,N_5623,N_4540);
or U7301 (N_7301,N_5635,N_4184);
xor U7302 (N_7302,N_5778,N_5156);
nor U7303 (N_7303,N_4992,N_4114);
nand U7304 (N_7304,N_4845,N_5923);
nor U7305 (N_7305,N_4796,N_5945);
xor U7306 (N_7306,N_5818,N_5943);
or U7307 (N_7307,N_4693,N_4576);
nand U7308 (N_7308,N_5745,N_4886);
xor U7309 (N_7309,N_4575,N_5153);
and U7310 (N_7310,N_5488,N_5825);
or U7311 (N_7311,N_4886,N_4735);
nor U7312 (N_7312,N_5341,N_4885);
nor U7313 (N_7313,N_4250,N_4380);
nor U7314 (N_7314,N_5806,N_5869);
and U7315 (N_7315,N_4136,N_4030);
or U7316 (N_7316,N_5466,N_4823);
nand U7317 (N_7317,N_4254,N_5964);
or U7318 (N_7318,N_5517,N_4956);
or U7319 (N_7319,N_4407,N_4116);
or U7320 (N_7320,N_4642,N_5505);
or U7321 (N_7321,N_4115,N_4686);
nor U7322 (N_7322,N_4390,N_4970);
and U7323 (N_7323,N_4069,N_5440);
xor U7324 (N_7324,N_5188,N_5633);
or U7325 (N_7325,N_5327,N_5775);
or U7326 (N_7326,N_4507,N_5380);
or U7327 (N_7327,N_4502,N_5321);
or U7328 (N_7328,N_5725,N_4993);
nand U7329 (N_7329,N_4642,N_4801);
and U7330 (N_7330,N_4456,N_5765);
or U7331 (N_7331,N_5654,N_4111);
or U7332 (N_7332,N_5855,N_5212);
nor U7333 (N_7333,N_5960,N_5559);
xnor U7334 (N_7334,N_4861,N_4278);
and U7335 (N_7335,N_4349,N_4206);
or U7336 (N_7336,N_5787,N_5686);
or U7337 (N_7337,N_4194,N_5993);
and U7338 (N_7338,N_5259,N_4570);
and U7339 (N_7339,N_5999,N_4725);
nand U7340 (N_7340,N_4972,N_4459);
nand U7341 (N_7341,N_4139,N_4157);
nand U7342 (N_7342,N_4815,N_5376);
nor U7343 (N_7343,N_5911,N_5719);
nand U7344 (N_7344,N_5152,N_5900);
nor U7345 (N_7345,N_5683,N_5987);
nor U7346 (N_7346,N_5085,N_5209);
xnor U7347 (N_7347,N_5187,N_5713);
nor U7348 (N_7348,N_5589,N_4177);
or U7349 (N_7349,N_4392,N_5309);
nand U7350 (N_7350,N_5469,N_5146);
or U7351 (N_7351,N_4494,N_5266);
and U7352 (N_7352,N_4224,N_5009);
nor U7353 (N_7353,N_4230,N_4283);
nand U7354 (N_7354,N_4132,N_4551);
and U7355 (N_7355,N_5919,N_4302);
nor U7356 (N_7356,N_5149,N_4452);
or U7357 (N_7357,N_4788,N_4266);
nand U7358 (N_7358,N_5941,N_5490);
and U7359 (N_7359,N_5080,N_4620);
and U7360 (N_7360,N_4286,N_4565);
and U7361 (N_7361,N_4148,N_4004);
nor U7362 (N_7362,N_5912,N_5202);
or U7363 (N_7363,N_4484,N_4592);
nand U7364 (N_7364,N_5996,N_5053);
nand U7365 (N_7365,N_4407,N_4224);
nand U7366 (N_7366,N_4034,N_4427);
or U7367 (N_7367,N_5926,N_5845);
and U7368 (N_7368,N_4888,N_5047);
or U7369 (N_7369,N_4016,N_4754);
and U7370 (N_7370,N_5029,N_5003);
nand U7371 (N_7371,N_5113,N_4766);
nand U7372 (N_7372,N_4953,N_5525);
or U7373 (N_7373,N_4828,N_5989);
and U7374 (N_7374,N_4090,N_4720);
or U7375 (N_7375,N_4821,N_5892);
and U7376 (N_7376,N_5216,N_5217);
nor U7377 (N_7377,N_4258,N_4540);
nor U7378 (N_7378,N_4559,N_5240);
and U7379 (N_7379,N_4328,N_5725);
and U7380 (N_7380,N_5866,N_4654);
nor U7381 (N_7381,N_4797,N_4810);
nor U7382 (N_7382,N_4200,N_5571);
nor U7383 (N_7383,N_5980,N_5615);
nor U7384 (N_7384,N_5718,N_4414);
and U7385 (N_7385,N_5939,N_5535);
nand U7386 (N_7386,N_5779,N_5264);
or U7387 (N_7387,N_4563,N_4925);
nand U7388 (N_7388,N_5102,N_4370);
or U7389 (N_7389,N_4144,N_5574);
or U7390 (N_7390,N_5056,N_4194);
nor U7391 (N_7391,N_4784,N_4925);
nand U7392 (N_7392,N_4885,N_4379);
or U7393 (N_7393,N_4613,N_5388);
and U7394 (N_7394,N_4736,N_5347);
nor U7395 (N_7395,N_4750,N_5878);
xor U7396 (N_7396,N_5089,N_4485);
nor U7397 (N_7397,N_5464,N_5697);
and U7398 (N_7398,N_5937,N_5379);
and U7399 (N_7399,N_4447,N_5003);
xor U7400 (N_7400,N_5292,N_5878);
nor U7401 (N_7401,N_4386,N_5072);
nand U7402 (N_7402,N_4976,N_5121);
nor U7403 (N_7403,N_4415,N_4169);
or U7404 (N_7404,N_4461,N_4748);
nand U7405 (N_7405,N_5668,N_5717);
nand U7406 (N_7406,N_5344,N_4231);
nor U7407 (N_7407,N_5580,N_4618);
xnor U7408 (N_7408,N_5049,N_5979);
and U7409 (N_7409,N_4577,N_5583);
nor U7410 (N_7410,N_4934,N_5044);
xor U7411 (N_7411,N_4822,N_5686);
or U7412 (N_7412,N_4480,N_5953);
xnor U7413 (N_7413,N_4542,N_4681);
nand U7414 (N_7414,N_5083,N_5404);
nand U7415 (N_7415,N_5066,N_4395);
or U7416 (N_7416,N_4739,N_4871);
xnor U7417 (N_7417,N_5890,N_5802);
nand U7418 (N_7418,N_5869,N_5364);
xnor U7419 (N_7419,N_5385,N_4623);
nand U7420 (N_7420,N_5326,N_4315);
xor U7421 (N_7421,N_4767,N_5052);
or U7422 (N_7422,N_5785,N_4110);
nand U7423 (N_7423,N_5767,N_5430);
and U7424 (N_7424,N_5936,N_4499);
nand U7425 (N_7425,N_4669,N_4951);
xor U7426 (N_7426,N_4986,N_4322);
and U7427 (N_7427,N_4880,N_5346);
or U7428 (N_7428,N_4492,N_5506);
nor U7429 (N_7429,N_4333,N_5227);
or U7430 (N_7430,N_4929,N_4618);
and U7431 (N_7431,N_4492,N_5916);
nor U7432 (N_7432,N_5326,N_4739);
or U7433 (N_7433,N_4944,N_5544);
and U7434 (N_7434,N_5720,N_5637);
nor U7435 (N_7435,N_5598,N_4061);
and U7436 (N_7436,N_5472,N_4324);
xnor U7437 (N_7437,N_5133,N_5054);
and U7438 (N_7438,N_4564,N_5870);
nand U7439 (N_7439,N_5445,N_4228);
nor U7440 (N_7440,N_4464,N_5062);
nor U7441 (N_7441,N_5167,N_5854);
or U7442 (N_7442,N_5773,N_4438);
and U7443 (N_7443,N_4858,N_4003);
or U7444 (N_7444,N_4765,N_4260);
or U7445 (N_7445,N_4887,N_4902);
nor U7446 (N_7446,N_4317,N_4622);
and U7447 (N_7447,N_4433,N_4643);
or U7448 (N_7448,N_5537,N_4243);
nor U7449 (N_7449,N_5782,N_4946);
and U7450 (N_7450,N_5174,N_5857);
xnor U7451 (N_7451,N_5176,N_5454);
or U7452 (N_7452,N_4282,N_4792);
nor U7453 (N_7453,N_4621,N_5464);
and U7454 (N_7454,N_5309,N_4922);
or U7455 (N_7455,N_5799,N_4070);
nand U7456 (N_7456,N_5091,N_4203);
xor U7457 (N_7457,N_5463,N_5994);
nand U7458 (N_7458,N_5965,N_4102);
or U7459 (N_7459,N_5886,N_4196);
nand U7460 (N_7460,N_4160,N_4799);
and U7461 (N_7461,N_5759,N_4611);
nand U7462 (N_7462,N_5267,N_4549);
or U7463 (N_7463,N_4594,N_5518);
xor U7464 (N_7464,N_5049,N_4116);
and U7465 (N_7465,N_4686,N_5452);
nand U7466 (N_7466,N_4828,N_5044);
or U7467 (N_7467,N_5644,N_5989);
or U7468 (N_7468,N_5575,N_5076);
nor U7469 (N_7469,N_4725,N_4167);
nor U7470 (N_7470,N_4147,N_5233);
and U7471 (N_7471,N_5547,N_5295);
and U7472 (N_7472,N_5622,N_4112);
or U7473 (N_7473,N_4269,N_5261);
and U7474 (N_7474,N_5324,N_5321);
nor U7475 (N_7475,N_4403,N_5443);
and U7476 (N_7476,N_4905,N_4486);
and U7477 (N_7477,N_4415,N_5584);
nor U7478 (N_7478,N_5671,N_4789);
or U7479 (N_7479,N_5854,N_4964);
nand U7480 (N_7480,N_5807,N_5926);
nor U7481 (N_7481,N_4135,N_4714);
and U7482 (N_7482,N_5698,N_5519);
nand U7483 (N_7483,N_4188,N_4365);
and U7484 (N_7484,N_4454,N_5960);
nor U7485 (N_7485,N_5202,N_4900);
or U7486 (N_7486,N_5806,N_5964);
or U7487 (N_7487,N_4255,N_4745);
and U7488 (N_7488,N_5491,N_5772);
and U7489 (N_7489,N_5518,N_4212);
xor U7490 (N_7490,N_4721,N_4356);
and U7491 (N_7491,N_4490,N_4083);
nor U7492 (N_7492,N_4312,N_5149);
nand U7493 (N_7493,N_4127,N_4917);
nand U7494 (N_7494,N_5613,N_4124);
nand U7495 (N_7495,N_5480,N_5221);
or U7496 (N_7496,N_4448,N_4927);
nand U7497 (N_7497,N_5187,N_5388);
nor U7498 (N_7498,N_4224,N_5375);
nor U7499 (N_7499,N_5949,N_4348);
or U7500 (N_7500,N_5135,N_5625);
nor U7501 (N_7501,N_5757,N_4785);
nand U7502 (N_7502,N_4485,N_5584);
and U7503 (N_7503,N_4921,N_4137);
nor U7504 (N_7504,N_5319,N_4407);
xnor U7505 (N_7505,N_4837,N_4906);
xnor U7506 (N_7506,N_5976,N_5219);
and U7507 (N_7507,N_4629,N_4139);
and U7508 (N_7508,N_5111,N_5554);
nor U7509 (N_7509,N_5595,N_5990);
nand U7510 (N_7510,N_5252,N_4629);
nand U7511 (N_7511,N_4265,N_4764);
nand U7512 (N_7512,N_4220,N_5692);
nor U7513 (N_7513,N_4092,N_5596);
nor U7514 (N_7514,N_4618,N_5301);
xor U7515 (N_7515,N_4425,N_4481);
and U7516 (N_7516,N_5661,N_4206);
nor U7517 (N_7517,N_5392,N_4701);
and U7518 (N_7518,N_4202,N_4320);
nor U7519 (N_7519,N_5948,N_4923);
nor U7520 (N_7520,N_5129,N_5804);
xor U7521 (N_7521,N_5234,N_5745);
and U7522 (N_7522,N_5293,N_4530);
xor U7523 (N_7523,N_4397,N_4935);
nor U7524 (N_7524,N_5365,N_5900);
or U7525 (N_7525,N_4138,N_5180);
nand U7526 (N_7526,N_5620,N_4884);
xnor U7527 (N_7527,N_5347,N_4226);
or U7528 (N_7528,N_5644,N_5598);
or U7529 (N_7529,N_5470,N_5904);
nand U7530 (N_7530,N_5456,N_5909);
nor U7531 (N_7531,N_5061,N_5691);
or U7532 (N_7532,N_5070,N_5001);
nand U7533 (N_7533,N_5749,N_5517);
nor U7534 (N_7534,N_4925,N_4183);
nand U7535 (N_7535,N_5511,N_5331);
or U7536 (N_7536,N_4183,N_5474);
and U7537 (N_7537,N_5260,N_5484);
nor U7538 (N_7538,N_4422,N_5111);
or U7539 (N_7539,N_4324,N_5769);
nand U7540 (N_7540,N_4403,N_4996);
and U7541 (N_7541,N_4286,N_4032);
or U7542 (N_7542,N_4408,N_4723);
xnor U7543 (N_7543,N_5115,N_5942);
xor U7544 (N_7544,N_5127,N_5424);
nand U7545 (N_7545,N_5262,N_4795);
and U7546 (N_7546,N_4254,N_5115);
nand U7547 (N_7547,N_4592,N_4002);
nor U7548 (N_7548,N_5173,N_5110);
or U7549 (N_7549,N_4701,N_5407);
nand U7550 (N_7550,N_5690,N_4840);
nor U7551 (N_7551,N_4517,N_5591);
or U7552 (N_7552,N_5463,N_5308);
xor U7553 (N_7553,N_4414,N_4355);
or U7554 (N_7554,N_4811,N_4525);
or U7555 (N_7555,N_5716,N_5572);
nor U7556 (N_7556,N_4492,N_4391);
nor U7557 (N_7557,N_4643,N_4609);
nor U7558 (N_7558,N_4859,N_4579);
nand U7559 (N_7559,N_4458,N_5481);
nor U7560 (N_7560,N_4482,N_5905);
nor U7561 (N_7561,N_4225,N_5008);
nor U7562 (N_7562,N_4669,N_4919);
or U7563 (N_7563,N_4553,N_5612);
and U7564 (N_7564,N_5493,N_4561);
nand U7565 (N_7565,N_4791,N_4413);
nor U7566 (N_7566,N_5595,N_4031);
nor U7567 (N_7567,N_5160,N_4994);
and U7568 (N_7568,N_4078,N_4042);
nor U7569 (N_7569,N_4604,N_4894);
nand U7570 (N_7570,N_4385,N_4956);
nand U7571 (N_7571,N_5822,N_5773);
nand U7572 (N_7572,N_4102,N_5691);
xor U7573 (N_7573,N_4723,N_4664);
nand U7574 (N_7574,N_4164,N_4628);
nor U7575 (N_7575,N_4827,N_4250);
and U7576 (N_7576,N_4597,N_5797);
nand U7577 (N_7577,N_4343,N_4124);
nand U7578 (N_7578,N_5493,N_4763);
nor U7579 (N_7579,N_4039,N_4583);
or U7580 (N_7580,N_5376,N_4658);
and U7581 (N_7581,N_4388,N_5973);
nand U7582 (N_7582,N_5612,N_5371);
nand U7583 (N_7583,N_5556,N_5933);
nor U7584 (N_7584,N_4373,N_5238);
and U7585 (N_7585,N_5374,N_5329);
nand U7586 (N_7586,N_4083,N_5982);
nor U7587 (N_7587,N_4462,N_5551);
xnor U7588 (N_7588,N_4911,N_5167);
nor U7589 (N_7589,N_4055,N_5199);
or U7590 (N_7590,N_5930,N_5376);
nor U7591 (N_7591,N_5594,N_4688);
xor U7592 (N_7592,N_4507,N_5118);
and U7593 (N_7593,N_4030,N_4380);
nor U7594 (N_7594,N_4607,N_4423);
or U7595 (N_7595,N_5406,N_4623);
or U7596 (N_7596,N_4326,N_4959);
and U7597 (N_7597,N_4879,N_5124);
nand U7598 (N_7598,N_5583,N_5648);
nor U7599 (N_7599,N_4903,N_5486);
or U7600 (N_7600,N_4353,N_4800);
and U7601 (N_7601,N_4997,N_5945);
nor U7602 (N_7602,N_4193,N_5773);
nand U7603 (N_7603,N_4045,N_5810);
xnor U7604 (N_7604,N_4599,N_4396);
and U7605 (N_7605,N_4547,N_5201);
and U7606 (N_7606,N_4936,N_4969);
nor U7607 (N_7607,N_4432,N_4148);
nand U7608 (N_7608,N_5978,N_4000);
nor U7609 (N_7609,N_5993,N_4008);
nor U7610 (N_7610,N_5820,N_5254);
and U7611 (N_7611,N_4971,N_4766);
nor U7612 (N_7612,N_5845,N_5468);
or U7613 (N_7613,N_5424,N_5155);
or U7614 (N_7614,N_4342,N_5147);
nand U7615 (N_7615,N_5098,N_5632);
and U7616 (N_7616,N_5588,N_4428);
and U7617 (N_7617,N_4098,N_5471);
and U7618 (N_7618,N_5401,N_5671);
nor U7619 (N_7619,N_5414,N_5027);
and U7620 (N_7620,N_5950,N_5744);
nand U7621 (N_7621,N_5578,N_5739);
or U7622 (N_7622,N_4447,N_5802);
nand U7623 (N_7623,N_4985,N_4461);
nor U7624 (N_7624,N_4167,N_4178);
nand U7625 (N_7625,N_4289,N_4128);
and U7626 (N_7626,N_5050,N_5243);
or U7627 (N_7627,N_4985,N_5670);
xor U7628 (N_7628,N_4058,N_4792);
nor U7629 (N_7629,N_5168,N_5447);
and U7630 (N_7630,N_4052,N_4743);
or U7631 (N_7631,N_4350,N_4381);
or U7632 (N_7632,N_4459,N_4946);
nand U7633 (N_7633,N_5013,N_4957);
or U7634 (N_7634,N_4291,N_5751);
or U7635 (N_7635,N_5547,N_4401);
and U7636 (N_7636,N_4478,N_5106);
nand U7637 (N_7637,N_5030,N_5469);
or U7638 (N_7638,N_4948,N_4454);
nand U7639 (N_7639,N_5686,N_4410);
nor U7640 (N_7640,N_5694,N_4733);
nand U7641 (N_7641,N_5579,N_4462);
and U7642 (N_7642,N_5330,N_4076);
xnor U7643 (N_7643,N_5608,N_4358);
nand U7644 (N_7644,N_4528,N_5881);
or U7645 (N_7645,N_5823,N_5767);
and U7646 (N_7646,N_5135,N_4434);
and U7647 (N_7647,N_5788,N_5740);
and U7648 (N_7648,N_4900,N_5662);
nor U7649 (N_7649,N_4033,N_4310);
or U7650 (N_7650,N_4026,N_5158);
and U7651 (N_7651,N_5813,N_5468);
xor U7652 (N_7652,N_4374,N_5132);
nand U7653 (N_7653,N_4735,N_4608);
xor U7654 (N_7654,N_4569,N_4900);
nand U7655 (N_7655,N_5912,N_5006);
nor U7656 (N_7656,N_4167,N_4995);
and U7657 (N_7657,N_4355,N_5144);
nand U7658 (N_7658,N_4879,N_5920);
or U7659 (N_7659,N_4660,N_5526);
nor U7660 (N_7660,N_4474,N_4018);
nand U7661 (N_7661,N_4683,N_4927);
nand U7662 (N_7662,N_5645,N_5859);
nor U7663 (N_7663,N_4487,N_4460);
nand U7664 (N_7664,N_5293,N_4832);
nand U7665 (N_7665,N_4730,N_5717);
and U7666 (N_7666,N_5123,N_5871);
nor U7667 (N_7667,N_5597,N_4697);
nand U7668 (N_7668,N_4413,N_4132);
or U7669 (N_7669,N_4260,N_4805);
and U7670 (N_7670,N_5620,N_5053);
or U7671 (N_7671,N_5557,N_4428);
nand U7672 (N_7672,N_5057,N_4959);
nand U7673 (N_7673,N_5532,N_4845);
nand U7674 (N_7674,N_4522,N_5603);
nand U7675 (N_7675,N_5184,N_4478);
xnor U7676 (N_7676,N_4775,N_5176);
nor U7677 (N_7677,N_4129,N_5714);
nand U7678 (N_7678,N_5217,N_4114);
and U7679 (N_7679,N_5163,N_4051);
xnor U7680 (N_7680,N_5349,N_5816);
xnor U7681 (N_7681,N_4920,N_5902);
nand U7682 (N_7682,N_4688,N_4065);
or U7683 (N_7683,N_4988,N_4978);
and U7684 (N_7684,N_5940,N_5464);
or U7685 (N_7685,N_4386,N_4972);
nor U7686 (N_7686,N_4687,N_4019);
or U7687 (N_7687,N_5625,N_5852);
nor U7688 (N_7688,N_5221,N_4895);
xor U7689 (N_7689,N_4201,N_5062);
nor U7690 (N_7690,N_4945,N_5976);
and U7691 (N_7691,N_5906,N_5490);
nand U7692 (N_7692,N_5947,N_5534);
or U7693 (N_7693,N_5470,N_4017);
nor U7694 (N_7694,N_4284,N_5721);
xnor U7695 (N_7695,N_5570,N_4544);
and U7696 (N_7696,N_5051,N_5100);
nand U7697 (N_7697,N_5275,N_4397);
and U7698 (N_7698,N_5068,N_5211);
or U7699 (N_7699,N_4212,N_4096);
and U7700 (N_7700,N_5576,N_4586);
or U7701 (N_7701,N_4394,N_4857);
nor U7702 (N_7702,N_4268,N_5249);
or U7703 (N_7703,N_5575,N_5191);
xnor U7704 (N_7704,N_4048,N_4399);
and U7705 (N_7705,N_4411,N_5969);
nor U7706 (N_7706,N_4561,N_5747);
and U7707 (N_7707,N_5521,N_4160);
or U7708 (N_7708,N_5915,N_5839);
nand U7709 (N_7709,N_4443,N_4104);
nor U7710 (N_7710,N_4102,N_4285);
nor U7711 (N_7711,N_4808,N_5009);
and U7712 (N_7712,N_5677,N_5638);
and U7713 (N_7713,N_5437,N_4256);
and U7714 (N_7714,N_5833,N_5401);
or U7715 (N_7715,N_4439,N_5533);
nor U7716 (N_7716,N_4484,N_5507);
nand U7717 (N_7717,N_5987,N_5754);
nor U7718 (N_7718,N_4900,N_5474);
or U7719 (N_7719,N_4584,N_5574);
and U7720 (N_7720,N_4587,N_4858);
nand U7721 (N_7721,N_5069,N_5099);
or U7722 (N_7722,N_5797,N_4481);
nor U7723 (N_7723,N_4946,N_4504);
and U7724 (N_7724,N_4959,N_5489);
or U7725 (N_7725,N_4546,N_5102);
or U7726 (N_7726,N_5850,N_4373);
nand U7727 (N_7727,N_4032,N_4931);
and U7728 (N_7728,N_5257,N_4121);
nand U7729 (N_7729,N_4834,N_4315);
and U7730 (N_7730,N_5001,N_4741);
nand U7731 (N_7731,N_4942,N_4929);
or U7732 (N_7732,N_4991,N_5132);
or U7733 (N_7733,N_5293,N_4328);
nand U7734 (N_7734,N_5776,N_4492);
nand U7735 (N_7735,N_5038,N_5919);
or U7736 (N_7736,N_4201,N_5496);
nand U7737 (N_7737,N_4662,N_4305);
and U7738 (N_7738,N_5506,N_4110);
xor U7739 (N_7739,N_5371,N_5985);
nor U7740 (N_7740,N_5866,N_4028);
or U7741 (N_7741,N_5517,N_4867);
xor U7742 (N_7742,N_4007,N_4182);
nor U7743 (N_7743,N_4903,N_4607);
and U7744 (N_7744,N_4559,N_4962);
or U7745 (N_7745,N_5234,N_4102);
nor U7746 (N_7746,N_5179,N_5761);
nor U7747 (N_7747,N_5949,N_4343);
nand U7748 (N_7748,N_5638,N_5245);
or U7749 (N_7749,N_5334,N_5851);
or U7750 (N_7750,N_5356,N_4956);
nand U7751 (N_7751,N_5084,N_4222);
or U7752 (N_7752,N_5379,N_4755);
or U7753 (N_7753,N_5712,N_4079);
nor U7754 (N_7754,N_4803,N_5730);
and U7755 (N_7755,N_4602,N_4770);
or U7756 (N_7756,N_4625,N_5234);
nor U7757 (N_7757,N_5672,N_5709);
nand U7758 (N_7758,N_4333,N_5735);
nand U7759 (N_7759,N_4758,N_4428);
nand U7760 (N_7760,N_5534,N_5189);
or U7761 (N_7761,N_5989,N_5144);
and U7762 (N_7762,N_4315,N_5975);
nand U7763 (N_7763,N_5246,N_4323);
nand U7764 (N_7764,N_4449,N_5079);
nand U7765 (N_7765,N_4413,N_4943);
or U7766 (N_7766,N_4622,N_5386);
and U7767 (N_7767,N_4316,N_4566);
nor U7768 (N_7768,N_5572,N_5089);
and U7769 (N_7769,N_5589,N_4956);
xnor U7770 (N_7770,N_5154,N_5892);
nand U7771 (N_7771,N_4672,N_4363);
or U7772 (N_7772,N_4363,N_5531);
and U7773 (N_7773,N_5054,N_5425);
and U7774 (N_7774,N_5705,N_5483);
or U7775 (N_7775,N_5218,N_5875);
xnor U7776 (N_7776,N_4564,N_4771);
nor U7777 (N_7777,N_5720,N_4062);
and U7778 (N_7778,N_5639,N_5460);
or U7779 (N_7779,N_4431,N_4651);
nand U7780 (N_7780,N_5045,N_5845);
xnor U7781 (N_7781,N_4855,N_4225);
xor U7782 (N_7782,N_4582,N_4507);
nand U7783 (N_7783,N_5264,N_5166);
and U7784 (N_7784,N_4408,N_4902);
and U7785 (N_7785,N_5557,N_4272);
nor U7786 (N_7786,N_5000,N_5001);
and U7787 (N_7787,N_5383,N_5572);
and U7788 (N_7788,N_4638,N_5747);
nor U7789 (N_7789,N_4102,N_5919);
and U7790 (N_7790,N_4907,N_5667);
and U7791 (N_7791,N_4117,N_5074);
nand U7792 (N_7792,N_5377,N_4843);
and U7793 (N_7793,N_4633,N_4050);
nand U7794 (N_7794,N_4124,N_5799);
and U7795 (N_7795,N_4954,N_4247);
nor U7796 (N_7796,N_4410,N_4480);
or U7797 (N_7797,N_4141,N_4618);
nand U7798 (N_7798,N_5215,N_5219);
or U7799 (N_7799,N_5127,N_4847);
nor U7800 (N_7800,N_4016,N_5936);
nand U7801 (N_7801,N_5989,N_4138);
nand U7802 (N_7802,N_5456,N_5718);
nor U7803 (N_7803,N_4845,N_4184);
nand U7804 (N_7804,N_5374,N_4489);
nor U7805 (N_7805,N_4936,N_5215);
nand U7806 (N_7806,N_4372,N_4949);
nor U7807 (N_7807,N_4828,N_5976);
nor U7808 (N_7808,N_4020,N_5866);
nor U7809 (N_7809,N_5809,N_5203);
or U7810 (N_7810,N_5034,N_5048);
and U7811 (N_7811,N_4676,N_5660);
nor U7812 (N_7812,N_5970,N_4919);
nand U7813 (N_7813,N_5170,N_4749);
nor U7814 (N_7814,N_4730,N_5876);
and U7815 (N_7815,N_5230,N_4887);
nor U7816 (N_7816,N_4212,N_4581);
nand U7817 (N_7817,N_5066,N_5435);
and U7818 (N_7818,N_5575,N_5408);
nand U7819 (N_7819,N_5601,N_5411);
nand U7820 (N_7820,N_5336,N_5903);
nand U7821 (N_7821,N_5054,N_5154);
and U7822 (N_7822,N_4817,N_5811);
nand U7823 (N_7823,N_4149,N_5208);
and U7824 (N_7824,N_4298,N_5555);
nor U7825 (N_7825,N_5931,N_4012);
nor U7826 (N_7826,N_5988,N_5819);
nor U7827 (N_7827,N_4025,N_5329);
nand U7828 (N_7828,N_4204,N_5748);
or U7829 (N_7829,N_4137,N_4986);
or U7830 (N_7830,N_4268,N_4195);
and U7831 (N_7831,N_4722,N_5092);
nand U7832 (N_7832,N_5151,N_5313);
and U7833 (N_7833,N_5287,N_5491);
or U7834 (N_7834,N_5076,N_5013);
nor U7835 (N_7835,N_4029,N_4066);
xnor U7836 (N_7836,N_5358,N_4416);
xor U7837 (N_7837,N_5678,N_4190);
nor U7838 (N_7838,N_4636,N_4640);
or U7839 (N_7839,N_5718,N_4755);
xnor U7840 (N_7840,N_5353,N_4556);
nand U7841 (N_7841,N_5300,N_4032);
and U7842 (N_7842,N_4285,N_4519);
or U7843 (N_7843,N_5814,N_4066);
nor U7844 (N_7844,N_4312,N_4146);
nand U7845 (N_7845,N_4025,N_5844);
nor U7846 (N_7846,N_5879,N_5785);
nand U7847 (N_7847,N_5023,N_5922);
nor U7848 (N_7848,N_5580,N_4828);
nand U7849 (N_7849,N_4645,N_5140);
nand U7850 (N_7850,N_5335,N_5920);
nand U7851 (N_7851,N_4621,N_5152);
xnor U7852 (N_7852,N_5804,N_5677);
nor U7853 (N_7853,N_5184,N_4143);
or U7854 (N_7854,N_5614,N_4086);
or U7855 (N_7855,N_5275,N_4894);
and U7856 (N_7856,N_5487,N_5177);
or U7857 (N_7857,N_5290,N_4382);
nor U7858 (N_7858,N_4720,N_4463);
or U7859 (N_7859,N_4206,N_4375);
and U7860 (N_7860,N_4649,N_5705);
xor U7861 (N_7861,N_5149,N_5053);
nand U7862 (N_7862,N_5670,N_4035);
nand U7863 (N_7863,N_4915,N_5460);
nor U7864 (N_7864,N_5149,N_4565);
nand U7865 (N_7865,N_4651,N_5782);
nand U7866 (N_7866,N_5267,N_4613);
nand U7867 (N_7867,N_4536,N_4944);
or U7868 (N_7868,N_4967,N_5061);
nor U7869 (N_7869,N_5836,N_5716);
or U7870 (N_7870,N_4999,N_5602);
nor U7871 (N_7871,N_4069,N_4817);
and U7872 (N_7872,N_4724,N_4882);
xor U7873 (N_7873,N_4417,N_5918);
and U7874 (N_7874,N_4553,N_5389);
nor U7875 (N_7875,N_4794,N_5632);
and U7876 (N_7876,N_4743,N_4091);
xor U7877 (N_7877,N_4422,N_5775);
xor U7878 (N_7878,N_5781,N_5123);
nand U7879 (N_7879,N_5694,N_5355);
nor U7880 (N_7880,N_5598,N_4541);
or U7881 (N_7881,N_5972,N_5896);
or U7882 (N_7882,N_5409,N_5553);
or U7883 (N_7883,N_4980,N_5129);
nand U7884 (N_7884,N_4697,N_4365);
nor U7885 (N_7885,N_4732,N_5025);
and U7886 (N_7886,N_5365,N_4511);
and U7887 (N_7887,N_4584,N_4386);
or U7888 (N_7888,N_4524,N_4643);
nand U7889 (N_7889,N_4509,N_5634);
nand U7890 (N_7890,N_5406,N_4274);
nor U7891 (N_7891,N_5089,N_4513);
and U7892 (N_7892,N_4901,N_5913);
nand U7893 (N_7893,N_5827,N_4533);
nand U7894 (N_7894,N_4905,N_5526);
nand U7895 (N_7895,N_5270,N_5812);
or U7896 (N_7896,N_4565,N_5199);
nand U7897 (N_7897,N_5119,N_4621);
or U7898 (N_7898,N_4296,N_4241);
nand U7899 (N_7899,N_5130,N_4878);
and U7900 (N_7900,N_4442,N_5110);
xor U7901 (N_7901,N_4856,N_5767);
nor U7902 (N_7902,N_4622,N_5200);
or U7903 (N_7903,N_4562,N_4707);
and U7904 (N_7904,N_5765,N_4523);
nand U7905 (N_7905,N_4500,N_4752);
xor U7906 (N_7906,N_4191,N_4662);
xnor U7907 (N_7907,N_5032,N_4006);
nand U7908 (N_7908,N_5783,N_4985);
nand U7909 (N_7909,N_5879,N_5542);
nand U7910 (N_7910,N_4217,N_5587);
and U7911 (N_7911,N_5945,N_4827);
and U7912 (N_7912,N_5209,N_4229);
nand U7913 (N_7913,N_5908,N_5837);
nand U7914 (N_7914,N_4442,N_4670);
and U7915 (N_7915,N_4217,N_4450);
nand U7916 (N_7916,N_4465,N_4685);
or U7917 (N_7917,N_4828,N_4810);
xor U7918 (N_7918,N_4493,N_5789);
nor U7919 (N_7919,N_4931,N_4841);
nor U7920 (N_7920,N_5363,N_4344);
nand U7921 (N_7921,N_4159,N_4866);
and U7922 (N_7922,N_4422,N_4753);
and U7923 (N_7923,N_4459,N_5557);
nor U7924 (N_7924,N_4536,N_5464);
or U7925 (N_7925,N_5418,N_5793);
xnor U7926 (N_7926,N_5811,N_4877);
xnor U7927 (N_7927,N_5640,N_4814);
or U7928 (N_7928,N_4860,N_4584);
and U7929 (N_7929,N_4657,N_5016);
nor U7930 (N_7930,N_5037,N_4478);
and U7931 (N_7931,N_4912,N_4120);
nor U7932 (N_7932,N_4209,N_4766);
or U7933 (N_7933,N_5652,N_5732);
and U7934 (N_7934,N_5900,N_5291);
nor U7935 (N_7935,N_5617,N_4956);
and U7936 (N_7936,N_5153,N_5247);
nor U7937 (N_7937,N_5078,N_4425);
nor U7938 (N_7938,N_5139,N_4593);
nand U7939 (N_7939,N_4609,N_4529);
and U7940 (N_7940,N_4722,N_5599);
and U7941 (N_7941,N_4176,N_5949);
nand U7942 (N_7942,N_4097,N_5689);
nor U7943 (N_7943,N_5984,N_5622);
nor U7944 (N_7944,N_4365,N_5814);
and U7945 (N_7945,N_4903,N_4732);
nor U7946 (N_7946,N_5254,N_5767);
nand U7947 (N_7947,N_5308,N_4757);
nand U7948 (N_7948,N_5562,N_4735);
or U7949 (N_7949,N_4141,N_4466);
xor U7950 (N_7950,N_5293,N_5925);
xor U7951 (N_7951,N_4694,N_5124);
nor U7952 (N_7952,N_4207,N_5357);
xor U7953 (N_7953,N_4985,N_5222);
nor U7954 (N_7954,N_4158,N_5189);
nand U7955 (N_7955,N_5636,N_4714);
nand U7956 (N_7956,N_5082,N_5156);
and U7957 (N_7957,N_5020,N_5313);
and U7958 (N_7958,N_4390,N_4191);
nand U7959 (N_7959,N_4222,N_4366);
or U7960 (N_7960,N_4258,N_5697);
or U7961 (N_7961,N_4604,N_5156);
and U7962 (N_7962,N_5296,N_5769);
nor U7963 (N_7963,N_4638,N_5687);
nor U7964 (N_7964,N_4998,N_5054);
nor U7965 (N_7965,N_4424,N_4548);
xor U7966 (N_7966,N_5414,N_4047);
and U7967 (N_7967,N_5950,N_5864);
nor U7968 (N_7968,N_5365,N_5978);
nor U7969 (N_7969,N_5079,N_5527);
and U7970 (N_7970,N_4554,N_5806);
nand U7971 (N_7971,N_4996,N_4622);
nand U7972 (N_7972,N_5976,N_5457);
and U7973 (N_7973,N_5505,N_4510);
and U7974 (N_7974,N_4385,N_4423);
or U7975 (N_7975,N_4102,N_5586);
or U7976 (N_7976,N_4429,N_5923);
nand U7977 (N_7977,N_4971,N_4226);
and U7978 (N_7978,N_5817,N_5761);
and U7979 (N_7979,N_4900,N_5149);
and U7980 (N_7980,N_5551,N_4747);
nor U7981 (N_7981,N_4857,N_5880);
xnor U7982 (N_7982,N_4732,N_4691);
and U7983 (N_7983,N_4734,N_5252);
nor U7984 (N_7984,N_4337,N_5814);
nand U7985 (N_7985,N_5643,N_4696);
nand U7986 (N_7986,N_5239,N_5416);
and U7987 (N_7987,N_5248,N_4876);
and U7988 (N_7988,N_5899,N_4751);
and U7989 (N_7989,N_4338,N_4404);
and U7990 (N_7990,N_5043,N_5253);
nor U7991 (N_7991,N_4328,N_5566);
or U7992 (N_7992,N_4909,N_4431);
nor U7993 (N_7993,N_4502,N_5044);
nor U7994 (N_7994,N_4001,N_5334);
and U7995 (N_7995,N_5848,N_5126);
xor U7996 (N_7996,N_4372,N_4529);
nand U7997 (N_7997,N_5727,N_5146);
nor U7998 (N_7998,N_5725,N_5973);
nand U7999 (N_7999,N_4265,N_4813);
and U8000 (N_8000,N_6015,N_6188);
or U8001 (N_8001,N_7220,N_7881);
nor U8002 (N_8002,N_7356,N_6416);
nand U8003 (N_8003,N_7239,N_6685);
nand U8004 (N_8004,N_6641,N_6036);
or U8005 (N_8005,N_6670,N_6940);
or U8006 (N_8006,N_6239,N_7707);
nand U8007 (N_8007,N_7882,N_7498);
nor U8008 (N_8008,N_6403,N_7493);
or U8009 (N_8009,N_7227,N_6843);
and U8010 (N_8010,N_6819,N_6147);
and U8011 (N_8011,N_7742,N_6005);
nand U8012 (N_8012,N_7645,N_6802);
or U8013 (N_8013,N_6155,N_7791);
or U8014 (N_8014,N_6750,N_6320);
or U8015 (N_8015,N_7515,N_7388);
xnor U8016 (N_8016,N_6718,N_6253);
nor U8017 (N_8017,N_6775,N_7991);
nand U8018 (N_8018,N_7318,N_6247);
xnor U8019 (N_8019,N_6343,N_6182);
and U8020 (N_8020,N_6699,N_7661);
and U8021 (N_8021,N_6591,N_7215);
or U8022 (N_8022,N_7244,N_7408);
and U8023 (N_8023,N_7848,N_7091);
nor U8024 (N_8024,N_6812,N_7856);
xnor U8025 (N_8025,N_6352,N_7424);
nor U8026 (N_8026,N_7474,N_7787);
nor U8027 (N_8027,N_6118,N_6071);
nand U8028 (N_8028,N_6527,N_6866);
nor U8029 (N_8029,N_6386,N_6728);
nand U8030 (N_8030,N_7681,N_7055);
nor U8031 (N_8031,N_7549,N_6515);
nand U8032 (N_8032,N_6538,N_6771);
nor U8033 (N_8033,N_7970,N_7092);
nor U8034 (N_8034,N_6855,N_6469);
nand U8035 (N_8035,N_7930,N_7536);
and U8036 (N_8036,N_7421,N_6902);
or U8037 (N_8037,N_6034,N_7067);
or U8038 (N_8038,N_7072,N_7964);
nor U8039 (N_8039,N_6686,N_6969);
nand U8040 (N_8040,N_6178,N_6755);
nand U8041 (N_8041,N_6257,N_6391);
nand U8042 (N_8042,N_7500,N_6568);
nor U8043 (N_8043,N_6964,N_7073);
nor U8044 (N_8044,N_6776,N_7156);
nor U8045 (N_8045,N_7088,N_6097);
or U8046 (N_8046,N_6479,N_7189);
or U8047 (N_8047,N_7838,N_6704);
and U8048 (N_8048,N_6768,N_7444);
and U8049 (N_8049,N_6872,N_7404);
and U8050 (N_8050,N_7130,N_6306);
or U8051 (N_8051,N_7766,N_6384);
nor U8052 (N_8052,N_6206,N_6581);
or U8053 (N_8053,N_7668,N_6448);
and U8054 (N_8054,N_6026,N_6122);
or U8055 (N_8055,N_7869,N_6100);
nor U8056 (N_8056,N_7828,N_6562);
nor U8057 (N_8057,N_7658,N_7858);
and U8058 (N_8058,N_7103,N_7855);
nand U8059 (N_8059,N_6689,N_7935);
nor U8060 (N_8060,N_7062,N_6839);
nand U8061 (N_8061,N_6040,N_7816);
and U8062 (N_8062,N_6613,N_7927);
and U8063 (N_8063,N_7949,N_7354);
and U8064 (N_8064,N_6633,N_7265);
xor U8065 (N_8065,N_7229,N_7298);
and U8066 (N_8066,N_7011,N_6914);
nand U8067 (N_8067,N_6042,N_7983);
or U8068 (N_8068,N_6460,N_7851);
nor U8069 (N_8069,N_6319,N_6455);
or U8070 (N_8070,N_6476,N_7303);
and U8071 (N_8071,N_7995,N_7590);
nand U8072 (N_8072,N_7208,N_6463);
or U8073 (N_8073,N_7050,N_7247);
nand U8074 (N_8074,N_6123,N_6105);
or U8075 (N_8075,N_6961,N_7035);
and U8076 (N_8076,N_6959,N_6081);
nor U8077 (N_8077,N_7107,N_6294);
nand U8078 (N_8078,N_7235,N_7642);
and U8079 (N_8079,N_7297,N_6186);
or U8080 (N_8080,N_7916,N_7662);
nor U8081 (N_8081,N_6804,N_6066);
or U8082 (N_8082,N_7114,N_7326);
or U8083 (N_8083,N_7528,N_6321);
or U8084 (N_8084,N_7431,N_6258);
nor U8085 (N_8085,N_7969,N_7041);
and U8086 (N_8086,N_7894,N_6871);
xnor U8087 (N_8087,N_6430,N_7192);
nand U8088 (N_8088,N_6607,N_6989);
nand U8089 (N_8089,N_6052,N_7384);
and U8090 (N_8090,N_6124,N_7144);
or U8091 (N_8091,N_7441,N_7559);
or U8092 (N_8092,N_6903,N_7012);
nand U8093 (N_8093,N_7802,N_6133);
xor U8094 (N_8094,N_6811,N_6762);
and U8095 (N_8095,N_7826,N_6471);
or U8096 (N_8096,N_7100,N_6786);
and U8097 (N_8097,N_6393,N_6078);
nor U8098 (N_8098,N_6588,N_6963);
and U8099 (N_8099,N_7467,N_7213);
or U8100 (N_8100,N_7275,N_7255);
nand U8101 (N_8101,N_7320,N_6721);
or U8102 (N_8102,N_7601,N_7204);
nor U8103 (N_8103,N_6723,N_7005);
and U8104 (N_8104,N_6380,N_7730);
xnor U8105 (N_8105,N_6698,N_7439);
or U8106 (N_8106,N_6473,N_7110);
xnor U8107 (N_8107,N_7793,N_7806);
nor U8108 (N_8108,N_6706,N_7425);
and U8109 (N_8109,N_6162,N_6332);
nor U8110 (N_8110,N_6060,N_7322);
or U8111 (N_8111,N_7462,N_7734);
or U8112 (N_8112,N_6494,N_7284);
nand U8113 (N_8113,N_7785,N_6399);
nor U8114 (N_8114,N_6315,N_7455);
nand U8115 (N_8115,N_6763,N_7176);
or U8116 (N_8116,N_6345,N_6892);
nor U8117 (N_8117,N_6807,N_7951);
nand U8118 (N_8118,N_7080,N_6908);
and U8119 (N_8119,N_7909,N_6682);
and U8120 (N_8120,N_7934,N_6838);
nand U8121 (N_8121,N_6367,N_7922);
and U8122 (N_8122,N_7401,N_7154);
or U8123 (N_8123,N_6518,N_7723);
nor U8124 (N_8124,N_6278,N_7403);
or U8125 (N_8125,N_7956,N_7483);
and U8126 (N_8126,N_6957,N_6697);
nor U8127 (N_8127,N_7013,N_6372);
or U8128 (N_8128,N_7884,N_6475);
and U8129 (N_8129,N_6406,N_7953);
or U8130 (N_8130,N_7988,N_7621);
and U8131 (N_8131,N_6353,N_7537);
and U8132 (N_8132,N_6945,N_7046);
and U8133 (N_8133,N_7538,N_7256);
nor U8134 (N_8134,N_7150,N_6396);
and U8135 (N_8135,N_6067,N_6068);
nor U8136 (N_8136,N_7691,N_7727);
xnor U8137 (N_8137,N_7832,N_6255);
and U8138 (N_8138,N_7686,N_6464);
nand U8139 (N_8139,N_7967,N_7327);
nor U8140 (N_8140,N_6260,N_7885);
or U8141 (N_8141,N_6334,N_6268);
nand U8142 (N_8142,N_6116,N_6438);
nand U8143 (N_8143,N_7409,N_6417);
nor U8144 (N_8144,N_6285,N_7418);
or U8145 (N_8145,N_6314,N_6251);
nor U8146 (N_8146,N_7671,N_6595);
nand U8147 (N_8147,N_7544,N_7288);
nand U8148 (N_8148,N_7776,N_7034);
and U8149 (N_8149,N_7127,N_6004);
and U8150 (N_8150,N_7736,N_6262);
xnor U8151 (N_8151,N_7852,N_7739);
xor U8152 (N_8152,N_7593,N_7513);
nand U8153 (N_8153,N_6062,N_6057);
or U8154 (N_8154,N_7757,N_7812);
nand U8155 (N_8155,N_6120,N_7083);
nor U8156 (N_8156,N_7866,N_7992);
nand U8157 (N_8157,N_7854,N_6664);
nand U8158 (N_8158,N_6139,N_6210);
or U8159 (N_8159,N_7711,N_6385);
and U8160 (N_8160,N_6690,N_6934);
or U8161 (N_8161,N_7960,N_7698);
nand U8162 (N_8162,N_7664,N_7744);
nand U8163 (N_8163,N_7132,N_6678);
and U8164 (N_8164,N_6240,N_7160);
nor U8165 (N_8165,N_7924,N_7546);
and U8166 (N_8166,N_6025,N_6408);
or U8167 (N_8167,N_7429,N_7372);
or U8168 (N_8168,N_6414,N_7638);
nor U8169 (N_8169,N_6860,N_7604);
or U8170 (N_8170,N_6759,N_7184);
xnor U8171 (N_8171,N_6366,N_7936);
nand U8172 (N_8172,N_7302,N_7112);
nand U8173 (N_8173,N_7603,N_7774);
and U8174 (N_8174,N_7482,N_6712);
nor U8175 (N_8175,N_7231,N_7847);
and U8176 (N_8176,N_6900,N_7889);
nor U8177 (N_8177,N_7501,N_7068);
nand U8178 (N_8178,N_6044,N_6700);
and U8179 (N_8179,N_7299,N_7625);
nor U8180 (N_8180,N_7348,N_6939);
nor U8181 (N_8181,N_6970,N_7314);
or U8182 (N_8182,N_6286,N_7491);
nand U8183 (N_8183,N_7428,N_7173);
or U8184 (N_8184,N_6342,N_6952);
nand U8185 (N_8185,N_6785,N_6249);
nor U8186 (N_8186,N_7933,N_6427);
nor U8187 (N_8187,N_6478,N_6917);
nor U8188 (N_8188,N_7135,N_7081);
xor U8189 (N_8189,N_6128,N_7290);
or U8190 (N_8190,N_7412,N_7534);
xnor U8191 (N_8191,N_6039,N_7249);
and U8192 (N_8192,N_7839,N_6996);
and U8193 (N_8193,N_7560,N_6445);
or U8194 (N_8194,N_7712,N_6567);
or U8195 (N_8195,N_7400,N_7416);
nor U8196 (N_8196,N_7531,N_7841);
nand U8197 (N_8197,N_7989,N_6500);
or U8198 (N_8198,N_6852,N_7520);
or U8199 (N_8199,N_6295,N_6933);
xnor U8200 (N_8200,N_6291,N_6263);
nand U8201 (N_8201,N_7892,N_6671);
and U8202 (N_8202,N_7190,N_7883);
xnor U8203 (N_8203,N_6307,N_7516);
nand U8204 (N_8204,N_7362,N_7913);
nor U8205 (N_8205,N_6730,N_7719);
or U8206 (N_8206,N_6508,N_7872);
nand U8207 (N_8207,N_7366,N_7825);
xnor U8208 (N_8208,N_7651,N_6809);
nor U8209 (N_8209,N_7598,N_6511);
nor U8210 (N_8210,N_6442,N_6389);
nand U8211 (N_8211,N_6313,N_7556);
xnor U8212 (N_8212,N_7219,N_6956);
and U8213 (N_8213,N_6447,N_7104);
and U8214 (N_8214,N_6873,N_6101);
or U8215 (N_8215,N_6737,N_6805);
nand U8216 (N_8216,N_6371,N_7809);
and U8217 (N_8217,N_6622,N_6724);
or U8218 (N_8218,N_7485,N_7174);
xor U8219 (N_8219,N_7900,N_7319);
nor U8220 (N_8220,N_6790,N_7126);
nand U8221 (N_8221,N_6381,N_7074);
nor U8222 (N_8222,N_6646,N_6126);
nand U8223 (N_8223,N_7371,N_7612);
nand U8224 (N_8224,N_7078,N_6987);
or U8225 (N_8225,N_7543,N_7289);
nand U8226 (N_8226,N_6201,N_6615);
xnor U8227 (N_8227,N_6221,N_7955);
or U8228 (N_8228,N_6745,N_7783);
and U8229 (N_8229,N_6121,N_6844);
or U8230 (N_8230,N_7810,N_6894);
or U8231 (N_8231,N_6450,N_7307);
nand U8232 (N_8232,N_6451,N_6605);
xnor U8233 (N_8233,N_7937,N_7709);
nor U8234 (N_8234,N_6711,N_7242);
nor U8235 (N_8235,N_7205,N_6165);
xnor U8236 (N_8236,N_6864,N_7216);
and U8237 (N_8237,N_6621,N_6619);
nor U8238 (N_8238,N_6108,N_7963);
nand U8239 (N_8239,N_6275,N_7393);
nand U8240 (N_8240,N_6573,N_6254);
nand U8241 (N_8241,N_7910,N_7918);
or U8242 (N_8242,N_7607,N_6146);
and U8243 (N_8243,N_6041,N_6196);
nand U8244 (N_8244,N_7273,N_7039);
or U8245 (N_8245,N_6536,N_6069);
nand U8246 (N_8246,N_7495,N_7565);
nor U8247 (N_8247,N_7925,N_6997);
and U8248 (N_8248,N_7557,N_7340);
xnor U8249 (N_8249,N_7767,N_7310);
nand U8250 (N_8250,N_6610,N_6404);
nor U8251 (N_8251,N_6720,N_6218);
nor U8252 (N_8252,N_7090,N_6548);
nor U8253 (N_8253,N_7442,N_6922);
nor U8254 (N_8254,N_7695,N_7419);
nand U8255 (N_8255,N_7702,N_6364);
nand U8256 (N_8256,N_6842,N_6231);
nand U8257 (N_8257,N_7504,N_6798);
and U8258 (N_8258,N_6318,N_7923);
and U8259 (N_8259,N_7952,N_6800);
nor U8260 (N_8260,N_6620,N_7053);
or U8261 (N_8261,N_7102,N_7579);
nor U8262 (N_8262,N_7061,N_7669);
or U8263 (N_8263,N_6335,N_6533);
or U8264 (N_8264,N_6604,N_6377);
and U8265 (N_8265,N_6795,N_6836);
and U8266 (N_8266,N_6824,N_7486);
or U8267 (N_8267,N_6356,N_7152);
nand U8268 (N_8268,N_7186,N_7168);
or U8269 (N_8269,N_7182,N_6177);
and U8270 (N_8270,N_6891,N_7300);
nor U8271 (N_8271,N_7274,N_6074);
or U8272 (N_8272,N_6975,N_7007);
nand U8273 (N_8273,N_7064,N_7262);
or U8274 (N_8274,N_6109,N_7143);
and U8275 (N_8275,N_6297,N_6426);
nand U8276 (N_8276,N_6955,N_6830);
nor U8277 (N_8277,N_7606,N_7292);
nand U8278 (N_8278,N_7232,N_6898);
and U8279 (N_8279,N_7140,N_7682);
nand U8280 (N_8280,N_7045,N_7201);
and U8281 (N_8281,N_7870,N_6135);
and U8282 (N_8282,N_6183,N_6281);
or U8283 (N_8283,N_6715,N_6707);
and U8284 (N_8284,N_7361,N_6991);
and U8285 (N_8285,N_7058,N_7093);
and U8286 (N_8286,N_6951,N_7451);
or U8287 (N_8287,N_7646,N_6259);
and U8288 (N_8288,N_6194,N_6974);
or U8289 (N_8289,N_7465,N_7990);
or U8290 (N_8290,N_7976,N_6184);
nor U8291 (N_8291,N_7212,N_6046);
or U8292 (N_8292,N_6137,N_7908);
nand U8293 (N_8293,N_7700,N_7749);
or U8294 (N_8294,N_7394,N_7505);
nand U8295 (N_8295,N_6093,N_6953);
xor U8296 (N_8296,N_6098,N_7263);
nand U8297 (N_8297,N_6023,N_6777);
xnor U8298 (N_8298,N_6107,N_6629);
or U8299 (N_8299,N_7115,N_6136);
or U8300 (N_8300,N_7972,N_7094);
nor U8301 (N_8301,N_7611,N_7281);
and U8302 (N_8302,N_6048,N_6801);
and U8303 (N_8303,N_6211,N_6157);
nor U8304 (N_8304,N_6420,N_7716);
and U8305 (N_8305,N_7740,N_6783);
nand U8306 (N_8306,N_6490,N_6609);
xor U8307 (N_8307,N_7022,N_6761);
or U8308 (N_8308,N_6327,N_6654);
nand U8309 (N_8309,N_6672,N_7773);
or U8310 (N_8310,N_7240,N_7512);
nor U8311 (N_8311,N_7591,N_7510);
and U8312 (N_8312,N_7199,N_6459);
xor U8313 (N_8313,N_6960,N_6350);
xor U8314 (N_8314,N_6113,N_7808);
and U8315 (N_8315,N_6153,N_6973);
and U8316 (N_8316,N_7835,N_7985);
nand U8317 (N_8317,N_7617,N_6962);
nor U8318 (N_8318,N_6365,N_6637);
nand U8319 (N_8319,N_6106,N_6862);
nor U8320 (N_8320,N_6190,N_6596);
nand U8321 (N_8321,N_7487,N_6375);
and U8322 (N_8322,N_7118,N_7675);
or U8323 (N_8323,N_7121,N_6912);
nor U8324 (N_8324,N_6592,N_6289);
nand U8325 (N_8325,N_7001,N_6002);
or U8326 (N_8326,N_7296,N_6336);
xor U8327 (N_8327,N_7316,N_6944);
or U8328 (N_8328,N_6090,N_7162);
or U8329 (N_8329,N_7010,N_7640);
xor U8330 (N_8330,N_6053,N_7206);
nor U8331 (N_8331,N_7197,N_7301);
and U8332 (N_8332,N_7803,N_7123);
or U8333 (N_8333,N_7929,N_7021);
or U8334 (N_8334,N_7586,N_6663);
nor U8335 (N_8335,N_6822,N_7194);
and U8336 (N_8336,N_6560,N_6741);
nor U8337 (N_8337,N_6156,N_7752);
or U8338 (N_8338,N_7243,N_6616);
or U8339 (N_8339,N_6674,N_6911);
nor U8340 (N_8340,N_6631,N_6729);
nand U8341 (N_8341,N_7432,N_7622);
nor U8342 (N_8342,N_6432,N_6506);
nor U8343 (N_8343,N_7202,N_7195);
nand U8344 (N_8344,N_7333,N_6214);
or U8345 (N_8345,N_7113,N_6667);
and U8346 (N_8346,N_6612,N_7398);
and U8347 (N_8347,N_6696,N_7876);
nand U8348 (N_8348,N_7506,N_7759);
xnor U8349 (N_8349,N_6215,N_6213);
nand U8350 (N_8350,N_7368,N_7177);
or U8351 (N_8351,N_6859,N_6544);
and U8352 (N_8352,N_7098,N_6643);
nor U8353 (N_8353,N_6764,N_6409);
or U8354 (N_8354,N_7821,N_6941);
or U8355 (N_8355,N_7193,N_6732);
nand U8356 (N_8356,N_7595,N_7230);
and U8357 (N_8357,N_6825,N_6150);
nand U8358 (N_8358,N_6791,N_7373);
nand U8359 (N_8359,N_7427,N_7754);
and U8360 (N_8360,N_6228,N_7188);
and U8361 (N_8361,N_6833,N_6347);
and U8362 (N_8362,N_7345,N_6096);
and U8363 (N_8363,N_6936,N_6865);
nand U8364 (N_8364,N_7452,N_7349);
or U8365 (N_8365,N_7765,N_7629);
and U8366 (N_8366,N_7679,N_7508);
and U8367 (N_8367,N_6570,N_7788);
xnor U8368 (N_8368,N_6413,N_6129);
or U8369 (N_8369,N_7674,N_6179);
or U8370 (N_8370,N_7655,N_6276);
and U8371 (N_8371,N_7258,N_6738);
or U8372 (N_8372,N_6339,N_6423);
and U8373 (N_8373,N_7066,N_7893);
and U8374 (N_8374,N_7797,N_7308);
nand U8375 (N_8375,N_7267,N_7836);
nand U8376 (N_8376,N_7279,N_6920);
xnor U8377 (N_8377,N_6803,N_7632);
nand U8378 (N_8378,N_6348,N_7799);
nand U8379 (N_8379,N_7502,N_6823);
nor U8380 (N_8380,N_7597,N_6195);
or U8381 (N_8381,N_6001,N_7221);
nand U8382 (N_8382,N_6007,N_6870);
nor U8383 (N_8383,N_6895,N_6608);
nand U8384 (N_8384,N_7397,N_7693);
and U8385 (N_8385,N_7417,N_6694);
or U8386 (N_8386,N_7097,N_7943);
and U8387 (N_8387,N_6145,N_7831);
nor U8388 (N_8388,N_6958,N_7850);
nor U8389 (N_8389,N_7618,N_6378);
or U8390 (N_8390,N_6283,N_7450);
nand U8391 (N_8391,N_6131,N_6896);
and U8392 (N_8392,N_7911,N_6983);
xor U8393 (N_8393,N_6027,N_6466);
nand U8394 (N_8394,N_7903,N_7178);
or U8395 (N_8395,N_6235,N_7818);
nand U8396 (N_8396,N_7975,N_7353);
or U8397 (N_8397,N_6014,N_6174);
nor U8398 (N_8398,N_6837,N_7561);
or U8399 (N_8399,N_7382,N_6808);
nand U8400 (N_8400,N_6248,N_7004);
or U8401 (N_8401,N_7337,N_6424);
or U8402 (N_8402,N_6209,N_7214);
nor U8403 (N_8403,N_7552,N_7426);
or U8404 (N_8404,N_7666,N_7743);
nor U8405 (N_8405,N_7763,N_7370);
or U8406 (N_8406,N_6454,N_7492);
nand U8407 (N_8407,N_7840,N_7489);
and U8408 (N_8408,N_6861,N_7111);
and U8409 (N_8409,N_6232,N_7445);
nand U8410 (N_8410,N_7181,N_6887);
nor U8411 (N_8411,N_7522,N_7237);
nand U8412 (N_8412,N_6882,N_7673);
and U8413 (N_8413,N_7696,N_7470);
xnor U8414 (N_8414,N_6993,N_7280);
or U8415 (N_8415,N_7476,N_6635);
or U8416 (N_8416,N_7772,N_6489);
xor U8417 (N_8417,N_6496,N_7456);
or U8418 (N_8418,N_6185,N_7864);
nor U8419 (N_8419,N_7507,N_6360);
nor U8420 (N_8420,N_6269,N_7436);
and U8421 (N_8421,N_7987,N_7430);
nor U8422 (N_8422,N_7191,N_7804);
nor U8423 (N_8423,N_7962,N_7844);
and U8424 (N_8424,N_6598,N_6574);
nor U8425 (N_8425,N_6901,N_7926);
and U8426 (N_8426,N_6769,N_6191);
nand U8427 (N_8427,N_7351,N_7805);
nor U8428 (N_8428,N_7849,N_7217);
and U8429 (N_8429,N_6847,N_6867);
and U8430 (N_8430,N_7873,N_6487);
or U8431 (N_8431,N_6749,N_7095);
nand U8432 (N_8432,N_7086,N_6751);
and U8433 (N_8433,N_7583,N_7338);
and U8434 (N_8434,N_6256,N_6154);
nor U8435 (N_8435,N_6030,N_7391);
nor U8436 (N_8436,N_6316,N_6415);
nor U8437 (N_8437,N_7762,N_6111);
or U8438 (N_8438,N_6173,N_6532);
or U8439 (N_8439,N_7768,N_6784);
nor U8440 (N_8440,N_6242,N_6552);
and U8441 (N_8441,N_7139,N_6687);
and U8442 (N_8442,N_7136,N_7820);
nand U8443 (N_8443,N_6429,N_7721);
and U8444 (N_8444,N_7724,N_6169);
or U8445 (N_8445,N_7656,N_6502);
and U8446 (N_8446,N_7017,N_7570);
or U8447 (N_8447,N_6726,N_7713);
and U8448 (N_8448,N_7683,N_6766);
nand U8449 (N_8449,N_6468,N_7203);
and U8450 (N_8450,N_7484,N_7875);
or U8451 (N_8451,N_6421,N_6639);
nor U8452 (N_8452,N_7670,N_6024);
and U8453 (N_8453,N_7582,N_7547);
and U8454 (N_8454,N_7633,N_7920);
and U8455 (N_8455,N_7331,N_6590);
and U8456 (N_8456,N_7697,N_6757);
or U8457 (N_8457,N_6501,N_7580);
nor U8458 (N_8458,N_6885,N_6398);
nand U8459 (N_8459,N_7837,N_6405);
nor U8460 (N_8460,N_6159,N_7717);
nand U8461 (N_8461,N_7099,N_7518);
or U8462 (N_8462,N_6158,N_7703);
nand U8463 (N_8463,N_6788,N_6792);
nor U8464 (N_8464,N_7994,N_7545);
and U8465 (N_8465,N_7792,N_7735);
nor U8466 (N_8466,N_6302,N_6743);
nor U8467 (N_8467,N_7120,N_7690);
nand U8468 (N_8468,N_7172,N_6828);
nor U8469 (N_8469,N_6237,N_6680);
nand U8470 (N_8470,N_6714,N_7986);
or U8471 (N_8471,N_7525,N_7868);
nor U8472 (N_8472,N_7116,N_6702);
or U8473 (N_8473,N_7532,N_7974);
and U8474 (N_8474,N_7018,N_6488);
or U8475 (N_8475,N_7813,N_6264);
and U8476 (N_8476,N_6119,N_6238);
nor U8477 (N_8477,N_7392,N_7888);
and U8478 (N_8478,N_6580,N_7663);
and U8479 (N_8479,N_7755,N_7228);
xnor U8480 (N_8480,N_7905,N_6437);
and U8481 (N_8481,N_7965,N_6008);
and U8482 (N_8482,N_7261,N_7238);
nand U8483 (N_8483,N_7211,N_7339);
nand U8484 (N_8484,N_6559,N_6772);
nor U8485 (N_8485,N_7822,N_6328);
or U8486 (N_8486,N_6733,N_7834);
and U8487 (N_8487,N_7902,N_7644);
nor U8488 (N_8488,N_6834,N_6651);
and U8489 (N_8489,N_6362,N_6781);
nand U8490 (N_8490,N_7605,N_6695);
nand U8491 (N_8491,N_6298,N_7464);
xor U8492 (N_8492,N_7945,N_6461);
or U8493 (N_8493,N_7169,N_7183);
nand U8494 (N_8494,N_7344,N_7321);
xnor U8495 (N_8495,N_6103,N_7260);
nor U8496 (N_8496,N_7628,N_6207);
nand U8497 (N_8497,N_6486,N_7448);
xor U8498 (N_8498,N_6849,N_7355);
or U8499 (N_8499,N_6234,N_6428);
or U8500 (N_8500,N_6018,N_7946);
or U8501 (N_8501,N_7044,N_6199);
nor U8502 (N_8502,N_6815,N_6166);
nor U8503 (N_8503,N_6602,N_6065);
and U8504 (N_8504,N_6374,N_6086);
nand U8505 (N_8505,N_6152,N_6634);
or U8506 (N_8506,N_6725,N_6087);
xor U8507 (N_8507,N_6497,N_6739);
nor U8508 (N_8508,N_7131,N_6530);
xor U8509 (N_8509,N_6753,N_7798);
nor U8510 (N_8510,N_6623,N_6467);
or U8511 (N_8511,N_7015,N_7659);
or U8512 (N_8512,N_6831,N_7019);
xnor U8513 (N_8513,N_6170,N_6701);
and U8514 (N_8514,N_7896,N_6351);
or U8515 (N_8515,N_6440,N_7459);
nand U8516 (N_8516,N_6904,N_7016);
or U8517 (N_8517,N_7306,N_7751);
nor U8518 (N_8518,N_7179,N_6884);
and U8519 (N_8519,N_7931,N_7689);
nand U8520 (N_8520,N_6913,N_6181);
nand U8521 (N_8521,N_6063,N_6752);
nand U8522 (N_8522,N_7282,N_6329);
nand U8523 (N_8523,N_7732,N_6075);
xnor U8524 (N_8524,N_7047,N_6407);
nor U8525 (N_8525,N_6611,N_7399);
or U8526 (N_8526,N_7886,N_6740);
nand U8527 (N_8527,N_6094,N_6540);
nand U8528 (N_8528,N_6011,N_6341);
xor U8529 (N_8529,N_6326,N_7954);
or U8530 (N_8530,N_7814,N_6000);
nor U8531 (N_8531,N_6304,N_6789);
and U8532 (N_8532,N_6986,N_6927);
xnor U8533 (N_8533,N_7657,N_7328);
and U8534 (N_8534,N_6683,N_6303);
or U8535 (N_8535,N_6675,N_6600);
nor U8536 (N_8536,N_6309,N_7584);
and U8537 (N_8537,N_7225,N_6400);
or U8538 (N_8538,N_6110,N_6735);
nor U8539 (N_8539,N_6431,N_6528);
or U8540 (N_8540,N_7846,N_7207);
and U8541 (N_8541,N_7277,N_7890);
nor U8542 (N_8542,N_6484,N_7517);
or U8543 (N_8543,N_6879,N_7006);
nand U8544 (N_8544,N_6979,N_6453);
nand U8545 (N_8545,N_6549,N_7291);
nor U8546 (N_8546,N_6806,N_7057);
and U8547 (N_8547,N_6322,N_6187);
nor U8548 (N_8548,N_7271,N_6197);
and U8549 (N_8549,N_7999,N_6925);
and U8550 (N_8550,N_6551,N_7141);
or U8551 (N_8551,N_7396,N_6893);
and U8552 (N_8552,N_6708,N_6624);
or U8553 (N_8553,N_7947,N_7575);
and U8554 (N_8554,N_7159,N_6102);
nand U8555 (N_8555,N_7295,N_6797);
nor U8556 (N_8556,N_6731,N_7959);
xor U8557 (N_8557,N_7082,N_6693);
and U8558 (N_8558,N_6433,N_6446);
xor U8559 (N_8559,N_6292,N_7599);
or U8560 (N_8560,N_7973,N_6924);
nand U8561 (N_8561,N_7312,N_7198);
nor U8562 (N_8562,N_7653,N_6587);
or U8563 (N_8563,N_7478,N_7259);
and U8564 (N_8564,N_6205,N_6003);
or U8565 (N_8565,N_7978,N_6401);
nand U8566 (N_8566,N_7823,N_7581);
nor U8567 (N_8567,N_6033,N_7551);
xor U8568 (N_8568,N_6009,N_7175);
and U8569 (N_8569,N_6584,N_6627);
and U8570 (N_8570,N_7819,N_7684);
xnor U8571 (N_8571,N_6954,N_7027);
or U8572 (N_8572,N_6035,N_6586);
and U8573 (N_8573,N_7054,N_6436);
or U8574 (N_8574,N_7944,N_6223);
xnor U8575 (N_8575,N_6642,N_6492);
nand U8576 (N_8576,N_6225,N_6507);
and U8577 (N_8577,N_6832,N_6636);
or U8578 (N_8578,N_6813,N_7899);
nor U8579 (N_8579,N_7789,N_6688);
nor U8580 (N_8580,N_6899,N_6638);
or U8581 (N_8581,N_7402,N_6338);
xnor U8582 (N_8582,N_7075,N_7037);
nand U8583 (N_8583,N_7056,N_6216);
and U8584 (N_8584,N_7079,N_6976);
and U8585 (N_8585,N_6045,N_7438);
nor U8586 (N_8586,N_6013,N_7033);
xnor U8587 (N_8587,N_7148,N_6299);
and U8588 (N_8588,N_6038,N_7639);
nand U8589 (N_8589,N_7449,N_7494);
or U8590 (N_8590,N_7790,N_7272);
or U8591 (N_8591,N_7435,N_6668);
nand U8592 (N_8592,N_7647,N_6346);
nor U8593 (N_8593,N_6555,N_7842);
nand U8594 (N_8594,N_7223,N_7725);
or U8595 (N_8595,N_6114,N_7966);
and U8596 (N_8596,N_6918,N_7076);
or U8597 (N_8597,N_7738,N_6212);
or U8598 (N_8598,N_7264,N_7481);
nand U8599 (N_8599,N_7541,N_6868);
nor U8600 (N_8600,N_6370,N_7921);
xnor U8601 (N_8601,N_6845,N_6856);
or U8602 (N_8602,N_7151,N_6665);
nand U8603 (N_8603,N_6512,N_7251);
nor U8604 (N_8604,N_7968,N_7912);
and U8605 (N_8605,N_7002,N_7539);
nand U8606 (N_8606,N_6876,N_7209);
or U8607 (N_8607,N_6577,N_6773);
and U8608 (N_8608,N_7248,N_6545);
and U8609 (N_8609,N_6966,N_7938);
nor U8610 (N_8610,N_6521,N_6452);
nand U8611 (N_8611,N_6470,N_7125);
or U8612 (N_8612,N_6357,N_7294);
and U8613 (N_8613,N_6394,N_7817);
nor U8614 (N_8614,N_6583,N_7065);
or U8615 (N_8615,N_6282,N_7038);
xnor U8616 (N_8616,N_7710,N_7957);
or U8617 (N_8617,N_7626,N_6349);
and U8618 (N_8618,N_7466,N_6647);
nor U8619 (N_8619,N_6143,N_6043);
xnor U8620 (N_8620,N_6513,N_6531);
or U8621 (N_8621,N_7950,N_6499);
nand U8622 (N_8622,N_7210,N_6099);
xor U8623 (N_8623,N_7026,N_7915);
nor U8624 (N_8624,N_6519,N_7422);
and U8625 (N_8625,N_6198,N_7149);
nand U8626 (N_8626,N_6368,N_7024);
or U8627 (N_8627,N_7117,N_7602);
or U8628 (N_8628,N_6514,N_7252);
or U8629 (N_8629,N_6907,N_7677);
nand U8630 (N_8630,N_7286,N_7218);
nor U8631 (N_8631,N_6382,N_6919);
and U8632 (N_8632,N_6713,N_6984);
nor U8633 (N_8633,N_7753,N_6246);
and U8634 (N_8634,N_7998,N_6760);
and U8635 (N_8635,N_6888,N_6458);
xor U8636 (N_8636,N_6245,N_6656);
nor U8637 (N_8637,N_6589,N_6571);
or U8638 (N_8638,N_7387,N_7276);
or U8639 (N_8639,N_6241,N_6625);
or U8640 (N_8640,N_7323,N_6333);
xnor U8641 (N_8641,N_7760,N_7468);
or U8642 (N_8642,N_6265,N_7853);
nand U8643 (N_8643,N_6799,N_7680);
and U8644 (N_8644,N_6504,N_6710);
nand U8645 (N_8645,N_6778,N_7378);
nor U8646 (N_8646,N_7443,N_7919);
and U8647 (N_8647,N_6193,N_7728);
xnor U8648 (N_8648,N_7096,N_6267);
nand U8649 (N_8649,N_6599,N_7857);
nand U8650 (N_8650,N_6456,N_6937);
xnor U8651 (N_8651,N_7385,N_6534);
nand U8652 (N_8652,N_6767,N_6076);
xor U8653 (N_8653,N_7420,N_6554);
nor U8654 (N_8654,N_7860,N_7796);
nor U8655 (N_8655,N_6363,N_7981);
nand U8656 (N_8656,N_7324,N_6857);
xnor U8657 (N_8657,N_7627,N_6387);
and U8658 (N_8658,N_7386,N_6817);
nand U8659 (N_8659,N_6425,N_7161);
or U8660 (N_8660,N_6271,N_7257);
or U8661 (N_8661,N_7624,N_6716);
and U8662 (N_8662,N_7558,N_6863);
or U8663 (N_8663,N_7437,N_6061);
nor U8664 (N_8664,N_6943,N_7524);
nand U8665 (N_8665,N_6085,N_7133);
or U8666 (N_8666,N_6161,N_7003);
or U8667 (N_8667,N_6946,N_6709);
nand U8668 (N_8668,N_6127,N_7706);
nor U8669 (N_8669,N_7077,N_6200);
or U8670 (N_8670,N_7167,N_7600);
or U8671 (N_8671,N_7845,N_6331);
and U8672 (N_8672,N_6084,N_7554);
nor U8673 (N_8673,N_7589,N_7374);
nor U8674 (N_8674,N_7070,N_7778);
or U8675 (N_8675,N_7527,N_7358);
nand U8676 (N_8676,N_7233,N_7381);
nand U8677 (N_8677,N_7843,N_6383);
and U8678 (N_8678,N_7577,N_6485);
nand U8679 (N_8679,N_6029,N_6858);
nand U8680 (N_8680,N_7770,N_6498);
or U8681 (N_8681,N_7619,N_7285);
nand U8682 (N_8682,N_6869,N_7071);
nand U8683 (N_8683,N_7729,N_6539);
nor U8684 (N_8684,N_6132,N_6719);
and U8685 (N_8685,N_6657,N_6585);
or U8686 (N_8686,N_6915,N_6529);
xor U8687 (N_8687,N_6104,N_6296);
nor U8688 (N_8688,N_7676,N_7897);
or U8689 (N_8689,N_6546,N_7971);
and U8690 (N_8690,N_7824,N_7472);
nand U8691 (N_8691,N_6483,N_7996);
nand U8692 (N_8692,N_6050,N_6340);
nand U8693 (N_8693,N_7028,N_6968);
or U8694 (N_8694,N_6854,N_6717);
and U8695 (N_8695,N_6779,N_7490);
and U8696 (N_8696,N_7410,N_6826);
nand U8697 (N_8697,N_6658,N_6480);
nand U8698 (N_8698,N_6140,N_7250);
and U8699 (N_8699,N_7380,N_7153);
nand U8700 (N_8700,N_6503,N_6395);
or U8701 (N_8701,N_6361,N_7708);
or U8702 (N_8702,N_7369,N_6410);
and U8703 (N_8703,N_7948,N_7771);
or U8704 (N_8704,N_7571,N_6203);
and U8705 (N_8705,N_6443,N_6222);
and U8706 (N_8706,N_7119,N_7043);
or U8707 (N_8707,N_6640,N_6525);
xor U8708 (N_8708,N_6681,N_7059);
and U8709 (N_8709,N_7051,N_6523);
and U8710 (N_8710,N_6550,N_7413);
or U8711 (N_8711,N_7980,N_6305);
nand U8712 (N_8712,N_6653,N_6593);
or U8713 (N_8713,N_6142,N_7158);
or U8714 (N_8714,N_7961,N_6542);
and U8715 (N_8715,N_6233,N_6853);
and U8716 (N_8716,N_7463,N_6020);
nor U8717 (N_8717,N_6827,N_6850);
nand U8718 (N_8718,N_7383,N_6279);
and U8719 (N_8719,N_7025,N_6557);
or U8720 (N_8720,N_7283,N_7171);
nor U8721 (N_8721,N_7830,N_7042);
or U8722 (N_8722,N_7036,N_7128);
nand U8723 (N_8723,N_7958,N_6816);
nor U8724 (N_8724,N_6669,N_7807);
nor U8725 (N_8725,N_7715,N_7758);
nor U8726 (N_8726,N_7040,N_7613);
nand U8727 (N_8727,N_7069,N_7731);
nand U8728 (N_8728,N_6821,N_7609);
or U8729 (N_8729,N_6079,N_7365);
and U8730 (N_8730,N_7566,N_7245);
nand U8731 (N_8731,N_7722,N_6558);
nor U8732 (N_8732,N_7779,N_6301);
nand U8733 (N_8733,N_7769,N_7704);
nand U8734 (N_8734,N_7811,N_6547);
xnor U8735 (N_8735,N_7335,N_6117);
nor U8736 (N_8736,N_6505,N_6509);
nor U8737 (N_8737,N_7196,N_7052);
or U8738 (N_8738,N_6661,N_6402);
nand U8739 (N_8739,N_6561,N_7637);
nand U8740 (N_8740,N_7756,N_6780);
nand U8741 (N_8741,N_6935,N_6566);
nand U8742 (N_8742,N_6376,N_7750);
xnor U8743 (N_8743,N_6359,N_7129);
nor U8744 (N_8744,N_6810,N_6787);
nand U8745 (N_8745,N_7932,N_7170);
and U8746 (N_8746,N_7761,N_7530);
nor U8747 (N_8747,N_6392,N_7906);
or U8748 (N_8748,N_6614,N_6878);
or U8749 (N_8749,N_6618,N_6481);
and U8750 (N_8750,N_6054,N_7106);
nand U8751 (N_8751,N_7907,N_6411);
xnor U8752 (N_8752,N_7406,N_7939);
and U8753 (N_8753,N_7342,N_7615);
nand U8754 (N_8754,N_7737,N_6578);
nor U8755 (N_8755,N_7877,N_6388);
xnor U8756 (N_8756,N_6910,N_6626);
and U8757 (N_8757,N_6971,N_6051);
or U8758 (N_8758,N_6835,N_7748);
nor U8759 (N_8759,N_6736,N_6535);
nand U8760 (N_8760,N_6441,N_7146);
and U8761 (N_8761,N_7269,N_7145);
nor U8762 (N_8762,N_7649,N_7315);
xor U8763 (N_8763,N_6765,N_7993);
nand U8764 (N_8764,N_6217,N_6981);
or U8765 (N_8765,N_7720,N_7157);
or U8766 (N_8766,N_7784,N_6125);
nor U8767 (N_8767,N_7726,N_6064);
or U8768 (N_8768,N_7781,N_6358);
or U8769 (N_8769,N_6543,N_7166);
nor U8770 (N_8770,N_6921,N_7891);
or U8771 (N_8771,N_6418,N_7519);
nand U8772 (N_8772,N_6684,N_6164);
and U8773 (N_8773,N_7567,N_6644);
or U8774 (N_8774,N_7705,N_7375);
nand U8775 (N_8775,N_7741,N_6660);
or U8776 (N_8776,N_7667,N_6666);
and U8777 (N_8777,N_7089,N_7304);
and U8778 (N_8778,N_6070,N_6541);
nor U8779 (N_8779,N_7029,N_7977);
nor U8780 (N_8780,N_7648,N_6923);
nand U8781 (N_8781,N_6758,N_6355);
nor U8782 (N_8782,N_6679,N_6877);
and U8783 (N_8783,N_6010,N_7347);
or U8784 (N_8784,N_7576,N_6273);
nor U8785 (N_8785,N_7147,N_7568);
and U8786 (N_8786,N_6457,N_6597);
and U8787 (N_8787,N_7030,N_7352);
and U8788 (N_8788,N_7454,N_7569);
or U8789 (N_8789,N_6982,N_6649);
and U8790 (N_8790,N_7614,N_7236);
nor U8791 (N_8791,N_7268,N_6949);
nor U8792 (N_8792,N_6293,N_6226);
and U8793 (N_8793,N_7032,N_7650);
nand U8794 (N_8794,N_7278,N_7733);
nor U8795 (N_8795,N_6229,N_6266);
nand U8796 (N_8796,N_7101,N_7475);
nand U8797 (N_8797,N_7469,N_7473);
nand U8798 (N_8798,N_6703,N_7880);
xor U8799 (N_8799,N_6080,N_7620);
nand U8800 (N_8800,N_6323,N_7660);
and U8801 (N_8801,N_7997,N_6677);
and U8802 (N_8802,N_7747,N_7138);
nor U8803 (N_8803,N_7574,N_6890);
and U8804 (N_8804,N_7578,N_6280);
or U8805 (N_8805,N_7254,N_6491);
and U8806 (N_8806,N_7867,N_6330);
nand U8807 (N_8807,N_7241,N_6373);
nand U8808 (N_8808,N_7270,N_7982);
xor U8809 (N_8809,N_7477,N_6676);
and U8810 (N_8810,N_6994,N_7453);
or U8811 (N_8811,N_7457,N_6883);
nand U8812 (N_8812,N_7555,N_6603);
or U8813 (N_8813,N_6390,N_7782);
and U8814 (N_8814,N_7222,N_7496);
nand U8815 (N_8815,N_7940,N_6379);
or U8816 (N_8816,N_6148,N_6012);
xnor U8817 (N_8817,N_7874,N_6909);
nor U8818 (N_8818,N_6300,N_7395);
or U8819 (N_8819,N_6047,N_6524);
and U8820 (N_8820,N_6575,N_6742);
or U8821 (N_8821,N_6517,N_6916);
nand U8822 (N_8822,N_6645,N_7941);
and U8823 (N_8823,N_6482,N_6134);
nand U8824 (N_8824,N_6522,N_7415);
or U8825 (N_8825,N_6932,N_7446);
nor U8826 (N_8826,N_7572,N_7631);
or U8827 (N_8827,N_7137,N_7325);
or U8828 (N_8828,N_6722,N_7009);
xor U8829 (N_8829,N_7878,N_6705);
xor U8830 (N_8830,N_6848,N_7596);
nor U8831 (N_8831,N_6841,N_7616);
or U8832 (N_8832,N_6261,N_7652);
xnor U8833 (N_8833,N_7000,N_6889);
nor U8834 (N_8834,N_7862,N_7563);
xnor U8835 (N_8835,N_7357,N_7346);
nand U8836 (N_8836,N_6988,N_6756);
or U8837 (N_8837,N_7887,N_7562);
nor U8838 (N_8838,N_6144,N_6493);
nand U8839 (N_8839,N_6092,N_6734);
xor U8840 (N_8840,N_7861,N_7688);
nand U8841 (N_8841,N_6202,N_7234);
nor U8842 (N_8842,N_7360,N_6980);
and U8843 (N_8843,N_6310,N_7122);
xnor U8844 (N_8844,N_7461,N_6397);
nand U8845 (N_8845,N_6032,N_6115);
and U8846 (N_8846,N_6272,N_6252);
xnor U8847 (N_8847,N_7311,N_6938);
or U8848 (N_8848,N_7521,N_6840);
and U8849 (N_8849,N_7390,N_7641);
xnor U8850 (N_8850,N_7458,N_6477);
nor U8851 (N_8851,N_7685,N_7984);
nor U8852 (N_8852,N_6942,N_6091);
or U8853 (N_8853,N_6793,N_7564);
or U8854 (N_8854,N_7594,N_6176);
or U8855 (N_8855,N_7503,N_6526);
or U8856 (N_8856,N_6985,N_7165);
nor U8857 (N_8857,N_6163,N_7087);
nor U8858 (N_8858,N_7509,N_7440);
nor U8859 (N_8859,N_6926,N_6650);
nor U8860 (N_8860,N_7678,N_7060);
nor U8861 (N_8861,N_6881,N_7701);
and U8862 (N_8862,N_6814,N_6874);
nor U8863 (N_8863,N_7049,N_7367);
nor U8864 (N_8864,N_7636,N_7411);
or U8865 (N_8865,N_6628,N_7334);
nor U8866 (N_8866,N_7665,N_6149);
and U8867 (N_8867,N_7800,N_6794);
and U8868 (N_8868,N_7898,N_7672);
and U8869 (N_8869,N_6058,N_6175);
nor U8870 (N_8870,N_6244,N_7871);
or U8871 (N_8871,N_6906,N_6172);
nor U8872 (N_8872,N_6462,N_7692);
or U8873 (N_8873,N_6171,N_7200);
nand U8874 (N_8874,N_6947,N_7533);
nand U8875 (N_8875,N_6082,N_6556);
or U8876 (N_8876,N_6141,N_7497);
xor U8877 (N_8877,N_7745,N_6439);
and U8878 (N_8878,N_7433,N_6754);
nor U8879 (N_8879,N_7350,N_7185);
or U8880 (N_8880,N_6230,N_6516);
nand U8881 (N_8881,N_6049,N_6782);
or U8882 (N_8882,N_6449,N_7901);
or U8883 (N_8883,N_7407,N_6325);
or U8884 (N_8884,N_6659,N_7488);
nor U8885 (N_8885,N_6056,N_6929);
or U8886 (N_8886,N_6208,N_7630);
and U8887 (N_8887,N_6059,N_6072);
nor U8888 (N_8888,N_6990,N_6016);
and U8889 (N_8889,N_7329,N_6189);
nor U8890 (N_8890,N_6655,N_7699);
nor U8891 (N_8891,N_7859,N_7542);
and U8892 (N_8892,N_7548,N_6652);
or U8893 (N_8893,N_6579,N_6998);
or U8894 (N_8894,N_6112,N_7460);
and U8895 (N_8895,N_7163,N_6875);
and U8896 (N_8896,N_7588,N_7523);
nor U8897 (N_8897,N_7511,N_6948);
and U8898 (N_8898,N_7928,N_7592);
and U8899 (N_8899,N_6250,N_7363);
nand U8900 (N_8900,N_7317,N_6277);
nand U8901 (N_8901,N_6021,N_7020);
xnor U8902 (N_8902,N_6077,N_6422);
and U8903 (N_8903,N_6083,N_6565);
and U8904 (N_8904,N_7942,N_7226);
xnor U8905 (N_8905,N_7377,N_6576);
and U8906 (N_8906,N_6317,N_7780);
nor U8907 (N_8907,N_6192,N_6287);
nand U8908 (N_8908,N_6037,N_6288);
nor U8909 (N_8909,N_7794,N_7332);
or U8910 (N_8910,N_7610,N_6846);
nand U8911 (N_8911,N_6474,N_7359);
nand U8912 (N_8912,N_7031,N_7313);
or U8913 (N_8913,N_6569,N_6829);
nor U8914 (N_8914,N_7376,N_7687);
nor U8915 (N_8915,N_6006,N_6662);
nor U8916 (N_8916,N_7305,N_6130);
nand U8917 (N_8917,N_7786,N_7405);
nand U8918 (N_8918,N_6897,N_6167);
xor U8919 (N_8919,N_6928,N_7635);
nor U8920 (N_8920,N_6747,N_7777);
or U8921 (N_8921,N_7573,N_7108);
nand U8922 (N_8922,N_6151,N_6630);
nand U8923 (N_8923,N_7587,N_6270);
xor U8924 (N_8924,N_7084,N_6180);
and U8925 (N_8925,N_6673,N_7471);
nand U8926 (N_8926,N_7085,N_7535);
nor U8927 (N_8927,N_7142,N_7801);
or U8928 (N_8928,N_7389,N_7364);
or U8929 (N_8929,N_6692,N_6369);
nor U8930 (N_8930,N_7643,N_6601);
nand U8931 (N_8931,N_6465,N_6274);
nand U8932 (N_8932,N_6617,N_7063);
nand U8933 (N_8933,N_7336,N_7879);
nor U8934 (N_8934,N_6243,N_6606);
nand U8935 (N_8935,N_6017,N_6999);
or U8936 (N_8936,N_6028,N_6648);
nand U8937 (N_8937,N_7134,N_7914);
or U8938 (N_8938,N_7827,N_6324);
and U8939 (N_8939,N_7865,N_6886);
nand U8940 (N_8940,N_6160,N_7917);
xor U8941 (N_8941,N_6419,N_7795);
nand U8942 (N_8942,N_6095,N_6972);
or U8943 (N_8943,N_6344,N_7023);
or U8944 (N_8944,N_7815,N_6227);
xor U8945 (N_8945,N_6995,N_6434);
or U8946 (N_8946,N_6290,N_6744);
or U8947 (N_8947,N_7124,N_7623);
nand U8948 (N_8948,N_7293,N_7694);
nor U8949 (N_8949,N_6880,N_7048);
and U8950 (N_8950,N_6691,N_7379);
nor U8951 (N_8951,N_6746,N_7224);
and U8952 (N_8952,N_6337,N_6851);
xor U8953 (N_8953,N_7187,N_6472);
or U8954 (N_8954,N_6495,N_6818);
or U8955 (N_8955,N_6594,N_6965);
nor U8956 (N_8956,N_6168,N_6931);
nand U8957 (N_8957,N_7634,N_6905);
and U8958 (N_8958,N_7529,N_7608);
and U8959 (N_8959,N_7266,N_7479);
nand U8960 (N_8960,N_6770,N_6219);
and U8961 (N_8961,N_6224,N_7434);
and U8962 (N_8962,N_6992,N_7341);
or U8963 (N_8963,N_6563,N_7423);
and U8964 (N_8964,N_6950,N_7109);
nand U8965 (N_8965,N_6930,N_7008);
nand U8966 (N_8966,N_7499,N_6796);
and U8967 (N_8967,N_6977,N_6236);
nor U8968 (N_8968,N_7904,N_6354);
or U8969 (N_8969,N_7654,N_7414);
xnor U8970 (N_8970,N_6727,N_7540);
or U8971 (N_8971,N_6073,N_6774);
nand U8972 (N_8972,N_6412,N_6022);
nand U8973 (N_8973,N_7829,N_6055);
xnor U8974 (N_8974,N_6572,N_6582);
nand U8975 (N_8975,N_7447,N_7164);
and U8976 (N_8976,N_7514,N_7895);
nand U8977 (N_8977,N_7526,N_6031);
and U8978 (N_8978,N_6510,N_6444);
nor U8979 (N_8979,N_7253,N_6632);
or U8980 (N_8980,N_7155,N_6138);
or U8981 (N_8981,N_7246,N_6748);
or U8982 (N_8982,N_7330,N_7833);
or U8983 (N_8983,N_7105,N_6820);
or U8984 (N_8984,N_6089,N_7718);
nor U8985 (N_8985,N_6978,N_7746);
xor U8986 (N_8986,N_7863,N_7979);
nand U8987 (N_8987,N_6019,N_7550);
and U8988 (N_8988,N_7764,N_6312);
xor U8989 (N_8989,N_6520,N_6088);
xor U8990 (N_8990,N_6308,N_7287);
nand U8991 (N_8991,N_7553,N_6284);
and U8992 (N_8992,N_6204,N_6553);
and U8993 (N_8993,N_6967,N_6220);
nor U8994 (N_8994,N_7014,N_7343);
nor U8995 (N_8995,N_7309,N_6311);
nor U8996 (N_8996,N_6537,N_6435);
or U8997 (N_8997,N_7775,N_7180);
nand U8998 (N_8998,N_7714,N_7585);
or U8999 (N_8999,N_7480,N_6564);
and U9000 (N_9000,N_7583,N_7108);
nand U9001 (N_9001,N_7323,N_6383);
nand U9002 (N_9002,N_7035,N_6995);
nand U9003 (N_9003,N_7694,N_6118);
xnor U9004 (N_9004,N_7241,N_6607);
nand U9005 (N_9005,N_7850,N_6331);
nand U9006 (N_9006,N_6840,N_7873);
nor U9007 (N_9007,N_6907,N_7525);
nand U9008 (N_9008,N_6874,N_7175);
nor U9009 (N_9009,N_7681,N_7820);
or U9010 (N_9010,N_7957,N_6765);
and U9011 (N_9011,N_7609,N_6902);
and U9012 (N_9012,N_7965,N_6622);
nor U9013 (N_9013,N_6749,N_7753);
nand U9014 (N_9014,N_6301,N_7046);
nor U9015 (N_9015,N_7160,N_7846);
and U9016 (N_9016,N_6581,N_7094);
nor U9017 (N_9017,N_7414,N_7524);
or U9018 (N_9018,N_7946,N_6472);
or U9019 (N_9019,N_7653,N_7782);
and U9020 (N_9020,N_6310,N_6727);
nand U9021 (N_9021,N_6112,N_6251);
or U9022 (N_9022,N_6672,N_6531);
nand U9023 (N_9023,N_7830,N_6729);
nand U9024 (N_9024,N_6688,N_6827);
xor U9025 (N_9025,N_6174,N_6239);
and U9026 (N_9026,N_6487,N_7558);
or U9027 (N_9027,N_7719,N_6811);
and U9028 (N_9028,N_6189,N_7441);
nor U9029 (N_9029,N_6316,N_7570);
or U9030 (N_9030,N_6723,N_7576);
or U9031 (N_9031,N_7564,N_6062);
nor U9032 (N_9032,N_6187,N_7171);
and U9033 (N_9033,N_7222,N_7880);
or U9034 (N_9034,N_7236,N_6402);
or U9035 (N_9035,N_7270,N_7459);
and U9036 (N_9036,N_6437,N_7608);
or U9037 (N_9037,N_7865,N_7733);
nand U9038 (N_9038,N_7439,N_7968);
nand U9039 (N_9039,N_6990,N_7229);
and U9040 (N_9040,N_7149,N_6244);
and U9041 (N_9041,N_6992,N_6624);
nor U9042 (N_9042,N_7565,N_7876);
or U9043 (N_9043,N_7388,N_6699);
nor U9044 (N_9044,N_6608,N_6992);
nor U9045 (N_9045,N_7305,N_7800);
nor U9046 (N_9046,N_6220,N_6342);
nand U9047 (N_9047,N_6647,N_7765);
and U9048 (N_9048,N_6473,N_7709);
and U9049 (N_9049,N_7560,N_7566);
nand U9050 (N_9050,N_6438,N_6203);
nor U9051 (N_9051,N_6954,N_6820);
nand U9052 (N_9052,N_6394,N_6633);
nand U9053 (N_9053,N_7322,N_6944);
and U9054 (N_9054,N_7038,N_6542);
nor U9055 (N_9055,N_7988,N_7005);
or U9056 (N_9056,N_6381,N_6530);
or U9057 (N_9057,N_7147,N_6382);
or U9058 (N_9058,N_7581,N_6790);
nor U9059 (N_9059,N_6416,N_7265);
or U9060 (N_9060,N_7385,N_7064);
and U9061 (N_9061,N_7934,N_7057);
and U9062 (N_9062,N_7878,N_6579);
nand U9063 (N_9063,N_7884,N_6107);
or U9064 (N_9064,N_7337,N_6325);
or U9065 (N_9065,N_7087,N_6803);
or U9066 (N_9066,N_6124,N_7120);
nand U9067 (N_9067,N_7749,N_7202);
or U9068 (N_9068,N_7781,N_6692);
or U9069 (N_9069,N_6909,N_7550);
or U9070 (N_9070,N_6531,N_7511);
and U9071 (N_9071,N_7057,N_7033);
and U9072 (N_9072,N_6549,N_7398);
nor U9073 (N_9073,N_6577,N_7509);
nand U9074 (N_9074,N_6102,N_7038);
nand U9075 (N_9075,N_7253,N_7038);
nor U9076 (N_9076,N_7328,N_7182);
or U9077 (N_9077,N_6322,N_6148);
nand U9078 (N_9078,N_6076,N_7883);
xnor U9079 (N_9079,N_7248,N_7619);
nand U9080 (N_9080,N_6262,N_6086);
nor U9081 (N_9081,N_7475,N_6295);
and U9082 (N_9082,N_7559,N_6430);
xor U9083 (N_9083,N_6834,N_7104);
or U9084 (N_9084,N_7639,N_6137);
and U9085 (N_9085,N_6795,N_6129);
or U9086 (N_9086,N_7841,N_7615);
and U9087 (N_9087,N_7959,N_6276);
and U9088 (N_9088,N_7559,N_6385);
xor U9089 (N_9089,N_7111,N_7729);
nor U9090 (N_9090,N_7604,N_6629);
xor U9091 (N_9091,N_6924,N_6147);
and U9092 (N_9092,N_7019,N_7581);
and U9093 (N_9093,N_7116,N_6808);
and U9094 (N_9094,N_6061,N_7170);
and U9095 (N_9095,N_6816,N_6863);
and U9096 (N_9096,N_7026,N_7433);
xor U9097 (N_9097,N_7381,N_6236);
or U9098 (N_9098,N_6163,N_6671);
nor U9099 (N_9099,N_6922,N_7949);
nand U9100 (N_9100,N_7175,N_7760);
or U9101 (N_9101,N_6423,N_7653);
or U9102 (N_9102,N_7037,N_6176);
or U9103 (N_9103,N_7219,N_7920);
or U9104 (N_9104,N_6553,N_6587);
or U9105 (N_9105,N_6507,N_7691);
xor U9106 (N_9106,N_7241,N_7571);
or U9107 (N_9107,N_6775,N_6737);
and U9108 (N_9108,N_6808,N_7574);
and U9109 (N_9109,N_6490,N_6797);
and U9110 (N_9110,N_6018,N_7486);
nand U9111 (N_9111,N_7069,N_6334);
or U9112 (N_9112,N_6590,N_6856);
nor U9113 (N_9113,N_7816,N_7988);
xnor U9114 (N_9114,N_7613,N_6876);
nand U9115 (N_9115,N_6697,N_7567);
nor U9116 (N_9116,N_6417,N_6847);
and U9117 (N_9117,N_6707,N_7635);
and U9118 (N_9118,N_7558,N_7867);
nand U9119 (N_9119,N_7800,N_6044);
nand U9120 (N_9120,N_7789,N_6123);
or U9121 (N_9121,N_6889,N_7974);
nand U9122 (N_9122,N_6866,N_7900);
nor U9123 (N_9123,N_7022,N_6146);
nand U9124 (N_9124,N_6856,N_6931);
nor U9125 (N_9125,N_6579,N_7063);
nor U9126 (N_9126,N_6605,N_7793);
xnor U9127 (N_9127,N_7623,N_7780);
or U9128 (N_9128,N_6964,N_6665);
nand U9129 (N_9129,N_6843,N_7668);
nand U9130 (N_9130,N_6324,N_7006);
nand U9131 (N_9131,N_6849,N_6338);
nor U9132 (N_9132,N_7926,N_7036);
nand U9133 (N_9133,N_6498,N_6654);
or U9134 (N_9134,N_7527,N_6707);
nor U9135 (N_9135,N_6307,N_6353);
nand U9136 (N_9136,N_6538,N_7558);
and U9137 (N_9137,N_6683,N_7922);
nor U9138 (N_9138,N_6868,N_6060);
xor U9139 (N_9139,N_6645,N_6291);
xnor U9140 (N_9140,N_7104,N_6176);
and U9141 (N_9141,N_6684,N_6901);
or U9142 (N_9142,N_7759,N_7075);
nor U9143 (N_9143,N_7408,N_6580);
or U9144 (N_9144,N_7306,N_6255);
nand U9145 (N_9145,N_7931,N_6226);
nand U9146 (N_9146,N_7005,N_6305);
nor U9147 (N_9147,N_6884,N_7144);
nand U9148 (N_9148,N_7036,N_7572);
and U9149 (N_9149,N_6392,N_6185);
xor U9150 (N_9150,N_6160,N_7941);
nand U9151 (N_9151,N_7143,N_6501);
nor U9152 (N_9152,N_6961,N_7402);
nor U9153 (N_9153,N_6907,N_6789);
nand U9154 (N_9154,N_6268,N_7833);
or U9155 (N_9155,N_7818,N_6297);
nand U9156 (N_9156,N_7924,N_6713);
nand U9157 (N_9157,N_7609,N_6422);
xor U9158 (N_9158,N_7211,N_6887);
nand U9159 (N_9159,N_6252,N_7784);
xor U9160 (N_9160,N_6095,N_6649);
nor U9161 (N_9161,N_6218,N_6157);
nand U9162 (N_9162,N_6674,N_7765);
xor U9163 (N_9163,N_7677,N_6415);
nand U9164 (N_9164,N_7604,N_6581);
and U9165 (N_9165,N_7891,N_6172);
or U9166 (N_9166,N_7180,N_7732);
nand U9167 (N_9167,N_6973,N_7401);
or U9168 (N_9168,N_7771,N_6113);
nor U9169 (N_9169,N_7978,N_6209);
nor U9170 (N_9170,N_6619,N_7192);
xor U9171 (N_9171,N_6355,N_6273);
and U9172 (N_9172,N_7051,N_7312);
xor U9173 (N_9173,N_6430,N_6078);
nand U9174 (N_9174,N_7853,N_6165);
xnor U9175 (N_9175,N_7484,N_6054);
nand U9176 (N_9176,N_6443,N_7504);
nor U9177 (N_9177,N_6810,N_6930);
and U9178 (N_9178,N_7980,N_7567);
and U9179 (N_9179,N_6974,N_7942);
or U9180 (N_9180,N_6672,N_7858);
xor U9181 (N_9181,N_6009,N_6048);
or U9182 (N_9182,N_6809,N_6981);
or U9183 (N_9183,N_6928,N_7386);
nand U9184 (N_9184,N_7245,N_7876);
or U9185 (N_9185,N_6479,N_6572);
xnor U9186 (N_9186,N_6046,N_7744);
or U9187 (N_9187,N_7178,N_7758);
nand U9188 (N_9188,N_6234,N_6921);
nand U9189 (N_9189,N_6254,N_7346);
nor U9190 (N_9190,N_6501,N_7851);
nand U9191 (N_9191,N_7027,N_7219);
nand U9192 (N_9192,N_7754,N_7932);
and U9193 (N_9193,N_7417,N_6834);
nor U9194 (N_9194,N_6393,N_6532);
or U9195 (N_9195,N_7787,N_7078);
nor U9196 (N_9196,N_6752,N_6257);
and U9197 (N_9197,N_7098,N_6762);
nand U9198 (N_9198,N_7831,N_7972);
nor U9199 (N_9199,N_6485,N_7952);
or U9200 (N_9200,N_6472,N_7697);
nor U9201 (N_9201,N_7767,N_6537);
and U9202 (N_9202,N_6051,N_6351);
or U9203 (N_9203,N_7926,N_6042);
or U9204 (N_9204,N_6108,N_7783);
and U9205 (N_9205,N_7021,N_6483);
and U9206 (N_9206,N_7028,N_7223);
and U9207 (N_9207,N_7169,N_7060);
xnor U9208 (N_9208,N_7730,N_7595);
or U9209 (N_9209,N_7430,N_6482);
and U9210 (N_9210,N_7969,N_7805);
nor U9211 (N_9211,N_6067,N_7883);
xor U9212 (N_9212,N_6892,N_7052);
or U9213 (N_9213,N_7944,N_7269);
nand U9214 (N_9214,N_6994,N_7741);
or U9215 (N_9215,N_7186,N_6791);
or U9216 (N_9216,N_6205,N_7758);
or U9217 (N_9217,N_7229,N_7559);
xor U9218 (N_9218,N_7061,N_6306);
nand U9219 (N_9219,N_6780,N_7800);
or U9220 (N_9220,N_7191,N_7846);
or U9221 (N_9221,N_6818,N_6115);
xnor U9222 (N_9222,N_6499,N_6045);
and U9223 (N_9223,N_6859,N_7828);
or U9224 (N_9224,N_6017,N_6575);
xor U9225 (N_9225,N_6728,N_7702);
nor U9226 (N_9226,N_7693,N_7644);
and U9227 (N_9227,N_7702,N_6615);
nor U9228 (N_9228,N_6825,N_7091);
or U9229 (N_9229,N_6869,N_6659);
and U9230 (N_9230,N_7009,N_7815);
or U9231 (N_9231,N_7776,N_6298);
and U9232 (N_9232,N_6912,N_7119);
nor U9233 (N_9233,N_6567,N_7518);
and U9234 (N_9234,N_7751,N_7728);
nand U9235 (N_9235,N_6738,N_6244);
nand U9236 (N_9236,N_6910,N_6717);
and U9237 (N_9237,N_6598,N_7399);
nand U9238 (N_9238,N_7962,N_7477);
and U9239 (N_9239,N_7832,N_7169);
xnor U9240 (N_9240,N_7752,N_6131);
xnor U9241 (N_9241,N_6761,N_6161);
xnor U9242 (N_9242,N_6320,N_6511);
nand U9243 (N_9243,N_7777,N_6365);
nor U9244 (N_9244,N_7220,N_6073);
xor U9245 (N_9245,N_6091,N_7362);
and U9246 (N_9246,N_6409,N_7994);
or U9247 (N_9247,N_6777,N_7852);
or U9248 (N_9248,N_7747,N_7473);
and U9249 (N_9249,N_6373,N_6193);
or U9250 (N_9250,N_7100,N_6606);
and U9251 (N_9251,N_6246,N_7607);
or U9252 (N_9252,N_7338,N_7198);
and U9253 (N_9253,N_7752,N_6475);
and U9254 (N_9254,N_7879,N_7106);
and U9255 (N_9255,N_6550,N_6227);
or U9256 (N_9256,N_6021,N_7290);
or U9257 (N_9257,N_6837,N_6464);
nor U9258 (N_9258,N_6135,N_6992);
nor U9259 (N_9259,N_6637,N_7838);
nor U9260 (N_9260,N_7251,N_7401);
nand U9261 (N_9261,N_7537,N_7746);
or U9262 (N_9262,N_7783,N_6762);
and U9263 (N_9263,N_7884,N_7109);
xnor U9264 (N_9264,N_6343,N_6846);
nand U9265 (N_9265,N_7779,N_6431);
nor U9266 (N_9266,N_7248,N_6098);
nand U9267 (N_9267,N_7529,N_6671);
and U9268 (N_9268,N_6987,N_6876);
and U9269 (N_9269,N_6173,N_7697);
nand U9270 (N_9270,N_7839,N_6317);
nor U9271 (N_9271,N_7810,N_6061);
nand U9272 (N_9272,N_6818,N_6286);
nand U9273 (N_9273,N_6500,N_6753);
and U9274 (N_9274,N_7974,N_7676);
and U9275 (N_9275,N_7674,N_7798);
or U9276 (N_9276,N_6035,N_7791);
or U9277 (N_9277,N_6147,N_6105);
or U9278 (N_9278,N_6164,N_7975);
nor U9279 (N_9279,N_7507,N_7060);
nor U9280 (N_9280,N_6761,N_7780);
nor U9281 (N_9281,N_6948,N_7979);
nor U9282 (N_9282,N_7623,N_6405);
and U9283 (N_9283,N_7704,N_7429);
nand U9284 (N_9284,N_6083,N_7756);
nor U9285 (N_9285,N_6950,N_6079);
or U9286 (N_9286,N_6779,N_6789);
nor U9287 (N_9287,N_7521,N_7106);
nor U9288 (N_9288,N_6671,N_6320);
xnor U9289 (N_9289,N_6230,N_7840);
nor U9290 (N_9290,N_6841,N_7221);
nor U9291 (N_9291,N_7746,N_6371);
and U9292 (N_9292,N_6378,N_7298);
and U9293 (N_9293,N_7695,N_7158);
nand U9294 (N_9294,N_6351,N_6843);
or U9295 (N_9295,N_7202,N_7514);
or U9296 (N_9296,N_6401,N_7322);
nand U9297 (N_9297,N_6494,N_7830);
nand U9298 (N_9298,N_6056,N_6286);
and U9299 (N_9299,N_6155,N_6975);
and U9300 (N_9300,N_6081,N_6771);
nand U9301 (N_9301,N_7361,N_6895);
nand U9302 (N_9302,N_6887,N_7111);
nor U9303 (N_9303,N_7361,N_7493);
xnor U9304 (N_9304,N_7075,N_7804);
nor U9305 (N_9305,N_6496,N_7416);
and U9306 (N_9306,N_7819,N_7614);
or U9307 (N_9307,N_6754,N_7971);
nand U9308 (N_9308,N_7411,N_6877);
and U9309 (N_9309,N_7651,N_7797);
xnor U9310 (N_9310,N_6527,N_7918);
nand U9311 (N_9311,N_7470,N_7638);
and U9312 (N_9312,N_7917,N_6759);
nor U9313 (N_9313,N_6877,N_7754);
and U9314 (N_9314,N_6856,N_6400);
nand U9315 (N_9315,N_6706,N_7337);
nor U9316 (N_9316,N_7271,N_7999);
xnor U9317 (N_9317,N_6703,N_7869);
xor U9318 (N_9318,N_7996,N_7750);
nor U9319 (N_9319,N_7633,N_6381);
nor U9320 (N_9320,N_7017,N_7078);
nand U9321 (N_9321,N_6323,N_6540);
or U9322 (N_9322,N_7774,N_6608);
nor U9323 (N_9323,N_6994,N_6862);
or U9324 (N_9324,N_6438,N_7367);
xnor U9325 (N_9325,N_7208,N_6882);
and U9326 (N_9326,N_6305,N_6173);
or U9327 (N_9327,N_7898,N_6483);
or U9328 (N_9328,N_7794,N_6678);
or U9329 (N_9329,N_6412,N_7919);
and U9330 (N_9330,N_7310,N_7872);
nand U9331 (N_9331,N_7227,N_7490);
nor U9332 (N_9332,N_7988,N_7265);
nand U9333 (N_9333,N_6553,N_6471);
or U9334 (N_9334,N_6897,N_6222);
nor U9335 (N_9335,N_6728,N_7261);
or U9336 (N_9336,N_7373,N_7828);
xnor U9337 (N_9337,N_6675,N_6389);
nand U9338 (N_9338,N_6746,N_7166);
nand U9339 (N_9339,N_6663,N_6842);
and U9340 (N_9340,N_7859,N_7905);
nor U9341 (N_9341,N_6938,N_7739);
nor U9342 (N_9342,N_6269,N_6354);
or U9343 (N_9343,N_7590,N_7412);
nand U9344 (N_9344,N_7328,N_6018);
nand U9345 (N_9345,N_6193,N_6677);
nand U9346 (N_9346,N_7913,N_6084);
and U9347 (N_9347,N_7324,N_6966);
nor U9348 (N_9348,N_7971,N_6783);
or U9349 (N_9349,N_7716,N_7416);
xor U9350 (N_9350,N_7316,N_7767);
nor U9351 (N_9351,N_6654,N_7203);
and U9352 (N_9352,N_7903,N_7376);
and U9353 (N_9353,N_6957,N_6380);
and U9354 (N_9354,N_6159,N_6773);
nor U9355 (N_9355,N_7145,N_7955);
and U9356 (N_9356,N_7545,N_7052);
or U9357 (N_9357,N_7715,N_7309);
nor U9358 (N_9358,N_7124,N_6545);
and U9359 (N_9359,N_6065,N_7481);
xor U9360 (N_9360,N_7625,N_7050);
nor U9361 (N_9361,N_7100,N_7966);
or U9362 (N_9362,N_6261,N_6196);
nand U9363 (N_9363,N_7740,N_7385);
nor U9364 (N_9364,N_6825,N_7794);
and U9365 (N_9365,N_7555,N_7752);
or U9366 (N_9366,N_6037,N_6147);
or U9367 (N_9367,N_7289,N_6110);
nor U9368 (N_9368,N_6607,N_7457);
nor U9369 (N_9369,N_7129,N_7531);
nand U9370 (N_9370,N_7466,N_6847);
or U9371 (N_9371,N_6685,N_6160);
nor U9372 (N_9372,N_7889,N_7060);
or U9373 (N_9373,N_7669,N_6570);
and U9374 (N_9374,N_7952,N_6776);
and U9375 (N_9375,N_7327,N_7111);
or U9376 (N_9376,N_6249,N_6770);
nand U9377 (N_9377,N_7030,N_7100);
and U9378 (N_9378,N_6332,N_6824);
and U9379 (N_9379,N_7730,N_7093);
or U9380 (N_9380,N_7152,N_7393);
and U9381 (N_9381,N_6395,N_6193);
or U9382 (N_9382,N_6032,N_6696);
and U9383 (N_9383,N_7777,N_6378);
nor U9384 (N_9384,N_7445,N_6265);
or U9385 (N_9385,N_7675,N_7635);
xnor U9386 (N_9386,N_7676,N_6090);
xnor U9387 (N_9387,N_6114,N_7575);
or U9388 (N_9388,N_7172,N_7176);
or U9389 (N_9389,N_6677,N_7885);
and U9390 (N_9390,N_6961,N_7539);
nor U9391 (N_9391,N_6746,N_6654);
nor U9392 (N_9392,N_7982,N_6281);
xnor U9393 (N_9393,N_6242,N_7430);
and U9394 (N_9394,N_6816,N_7051);
nor U9395 (N_9395,N_6835,N_6149);
nor U9396 (N_9396,N_7558,N_6789);
nand U9397 (N_9397,N_7188,N_7102);
and U9398 (N_9398,N_6794,N_6393);
nand U9399 (N_9399,N_6360,N_7001);
and U9400 (N_9400,N_6605,N_6325);
nor U9401 (N_9401,N_6074,N_6081);
xor U9402 (N_9402,N_7581,N_7701);
and U9403 (N_9403,N_7739,N_6568);
and U9404 (N_9404,N_7880,N_6964);
nand U9405 (N_9405,N_6012,N_6128);
nor U9406 (N_9406,N_6125,N_6168);
or U9407 (N_9407,N_6314,N_6627);
nand U9408 (N_9408,N_7664,N_7962);
xnor U9409 (N_9409,N_7518,N_6470);
nand U9410 (N_9410,N_7837,N_6034);
nand U9411 (N_9411,N_7091,N_6711);
or U9412 (N_9412,N_7510,N_6486);
xnor U9413 (N_9413,N_7381,N_6185);
and U9414 (N_9414,N_6841,N_7293);
nor U9415 (N_9415,N_7028,N_6128);
nand U9416 (N_9416,N_7254,N_6062);
and U9417 (N_9417,N_6522,N_6445);
and U9418 (N_9418,N_6231,N_6310);
and U9419 (N_9419,N_6101,N_7058);
and U9420 (N_9420,N_7797,N_7667);
nor U9421 (N_9421,N_6988,N_7523);
xnor U9422 (N_9422,N_7035,N_7039);
or U9423 (N_9423,N_6504,N_7877);
nor U9424 (N_9424,N_6806,N_7602);
or U9425 (N_9425,N_6076,N_7962);
nor U9426 (N_9426,N_6145,N_7964);
nand U9427 (N_9427,N_7972,N_7292);
and U9428 (N_9428,N_6767,N_7513);
nor U9429 (N_9429,N_7880,N_6601);
nor U9430 (N_9430,N_6792,N_7841);
and U9431 (N_9431,N_7237,N_7533);
and U9432 (N_9432,N_6445,N_7102);
or U9433 (N_9433,N_7364,N_6268);
or U9434 (N_9434,N_7628,N_6624);
nand U9435 (N_9435,N_7702,N_7029);
nand U9436 (N_9436,N_7535,N_6894);
nor U9437 (N_9437,N_7595,N_6939);
xnor U9438 (N_9438,N_7963,N_6516);
nor U9439 (N_9439,N_7240,N_6089);
xnor U9440 (N_9440,N_6615,N_7321);
and U9441 (N_9441,N_6839,N_7897);
and U9442 (N_9442,N_7289,N_6406);
nor U9443 (N_9443,N_7055,N_6774);
nand U9444 (N_9444,N_7094,N_6449);
nand U9445 (N_9445,N_6019,N_6601);
and U9446 (N_9446,N_7636,N_7660);
or U9447 (N_9447,N_6644,N_7196);
nor U9448 (N_9448,N_6143,N_6056);
or U9449 (N_9449,N_6177,N_6491);
or U9450 (N_9450,N_6547,N_6002);
and U9451 (N_9451,N_7129,N_7505);
nor U9452 (N_9452,N_6063,N_7966);
nand U9453 (N_9453,N_6190,N_7791);
nor U9454 (N_9454,N_6191,N_7930);
and U9455 (N_9455,N_6712,N_7149);
nor U9456 (N_9456,N_7519,N_6583);
nand U9457 (N_9457,N_7849,N_6881);
or U9458 (N_9458,N_7023,N_6955);
nand U9459 (N_9459,N_7293,N_6228);
and U9460 (N_9460,N_6855,N_6672);
or U9461 (N_9461,N_6155,N_6789);
or U9462 (N_9462,N_6711,N_6250);
nor U9463 (N_9463,N_7690,N_6340);
and U9464 (N_9464,N_6869,N_7201);
nor U9465 (N_9465,N_6191,N_6533);
and U9466 (N_9466,N_7847,N_7254);
or U9467 (N_9467,N_7547,N_7456);
nor U9468 (N_9468,N_6193,N_7789);
nor U9469 (N_9469,N_6898,N_7610);
and U9470 (N_9470,N_6685,N_6311);
and U9471 (N_9471,N_7532,N_6924);
or U9472 (N_9472,N_6972,N_7594);
nor U9473 (N_9473,N_6610,N_7399);
or U9474 (N_9474,N_7831,N_7044);
nor U9475 (N_9475,N_6871,N_6069);
or U9476 (N_9476,N_7354,N_6926);
and U9477 (N_9477,N_6138,N_7940);
nand U9478 (N_9478,N_6931,N_6854);
nand U9479 (N_9479,N_7111,N_7264);
or U9480 (N_9480,N_6832,N_6008);
nor U9481 (N_9481,N_7345,N_6964);
nor U9482 (N_9482,N_7645,N_6944);
xnor U9483 (N_9483,N_7571,N_7405);
and U9484 (N_9484,N_7778,N_6245);
and U9485 (N_9485,N_6075,N_6535);
nand U9486 (N_9486,N_7936,N_7190);
or U9487 (N_9487,N_7789,N_6276);
nand U9488 (N_9488,N_6664,N_6384);
nor U9489 (N_9489,N_6598,N_6769);
and U9490 (N_9490,N_6969,N_6540);
xor U9491 (N_9491,N_7328,N_6384);
nand U9492 (N_9492,N_6626,N_7382);
nand U9493 (N_9493,N_6958,N_6372);
or U9494 (N_9494,N_7207,N_7987);
or U9495 (N_9495,N_6521,N_7094);
nor U9496 (N_9496,N_6140,N_7320);
nand U9497 (N_9497,N_7232,N_6938);
and U9498 (N_9498,N_6827,N_6532);
nand U9499 (N_9499,N_6185,N_7136);
nand U9500 (N_9500,N_7077,N_7574);
nand U9501 (N_9501,N_7306,N_6857);
nand U9502 (N_9502,N_7382,N_6753);
nor U9503 (N_9503,N_7510,N_7604);
and U9504 (N_9504,N_6925,N_6037);
and U9505 (N_9505,N_7317,N_7711);
nor U9506 (N_9506,N_7844,N_6931);
nor U9507 (N_9507,N_7150,N_7279);
nand U9508 (N_9508,N_6527,N_6336);
or U9509 (N_9509,N_6031,N_6333);
and U9510 (N_9510,N_6855,N_6800);
or U9511 (N_9511,N_7853,N_6065);
and U9512 (N_9512,N_6057,N_6907);
or U9513 (N_9513,N_6626,N_6322);
or U9514 (N_9514,N_7875,N_6248);
nand U9515 (N_9515,N_6592,N_6380);
and U9516 (N_9516,N_7854,N_7422);
nand U9517 (N_9517,N_7618,N_7882);
and U9518 (N_9518,N_7753,N_7143);
and U9519 (N_9519,N_7079,N_6649);
nor U9520 (N_9520,N_7822,N_6397);
and U9521 (N_9521,N_6912,N_7701);
or U9522 (N_9522,N_7952,N_6803);
or U9523 (N_9523,N_7255,N_7368);
nand U9524 (N_9524,N_6738,N_7109);
or U9525 (N_9525,N_6897,N_7377);
nand U9526 (N_9526,N_7574,N_6119);
or U9527 (N_9527,N_7214,N_7621);
nor U9528 (N_9528,N_6797,N_6347);
or U9529 (N_9529,N_7558,N_6837);
or U9530 (N_9530,N_6640,N_7577);
and U9531 (N_9531,N_6603,N_6353);
nand U9532 (N_9532,N_6662,N_7584);
nand U9533 (N_9533,N_6330,N_7377);
nor U9534 (N_9534,N_7435,N_6022);
or U9535 (N_9535,N_6269,N_6248);
nand U9536 (N_9536,N_7397,N_7196);
or U9537 (N_9537,N_7137,N_6703);
xnor U9538 (N_9538,N_6719,N_7820);
nor U9539 (N_9539,N_6640,N_6128);
nand U9540 (N_9540,N_7108,N_7821);
nand U9541 (N_9541,N_6813,N_7786);
nor U9542 (N_9542,N_7907,N_7569);
or U9543 (N_9543,N_7150,N_7135);
and U9544 (N_9544,N_7800,N_7602);
nor U9545 (N_9545,N_7063,N_6074);
or U9546 (N_9546,N_7947,N_7346);
or U9547 (N_9547,N_7539,N_6398);
xor U9548 (N_9548,N_7343,N_6416);
xor U9549 (N_9549,N_6898,N_6540);
or U9550 (N_9550,N_6830,N_6137);
nand U9551 (N_9551,N_7434,N_6052);
nor U9552 (N_9552,N_6108,N_7000);
or U9553 (N_9553,N_7600,N_6421);
nor U9554 (N_9554,N_6498,N_7900);
nor U9555 (N_9555,N_7882,N_7935);
or U9556 (N_9556,N_6685,N_6222);
or U9557 (N_9557,N_6741,N_6984);
and U9558 (N_9558,N_6443,N_6089);
nand U9559 (N_9559,N_6888,N_7329);
or U9560 (N_9560,N_7497,N_6362);
nor U9561 (N_9561,N_6479,N_6658);
and U9562 (N_9562,N_7364,N_7271);
and U9563 (N_9563,N_6305,N_7643);
or U9564 (N_9564,N_7673,N_6236);
and U9565 (N_9565,N_7358,N_7586);
xor U9566 (N_9566,N_6244,N_7669);
and U9567 (N_9567,N_6089,N_7973);
nand U9568 (N_9568,N_7934,N_7278);
and U9569 (N_9569,N_6120,N_6700);
nand U9570 (N_9570,N_7717,N_6164);
xor U9571 (N_9571,N_6750,N_6305);
nor U9572 (N_9572,N_6086,N_7859);
xor U9573 (N_9573,N_6042,N_7468);
or U9574 (N_9574,N_7509,N_7156);
and U9575 (N_9575,N_6722,N_7366);
nand U9576 (N_9576,N_6716,N_7587);
or U9577 (N_9577,N_6039,N_7026);
and U9578 (N_9578,N_7997,N_7363);
and U9579 (N_9579,N_6639,N_7775);
nor U9580 (N_9580,N_7104,N_6886);
nor U9581 (N_9581,N_7090,N_7909);
xnor U9582 (N_9582,N_6205,N_7104);
nor U9583 (N_9583,N_7223,N_6188);
nand U9584 (N_9584,N_7327,N_6359);
nor U9585 (N_9585,N_7534,N_7489);
nor U9586 (N_9586,N_7605,N_7168);
and U9587 (N_9587,N_7558,N_6560);
nor U9588 (N_9588,N_7470,N_6356);
and U9589 (N_9589,N_7567,N_6105);
and U9590 (N_9590,N_7733,N_7657);
or U9591 (N_9591,N_7750,N_6400);
nor U9592 (N_9592,N_7674,N_7131);
and U9593 (N_9593,N_6152,N_6923);
nand U9594 (N_9594,N_6200,N_7582);
nand U9595 (N_9595,N_6898,N_6999);
and U9596 (N_9596,N_7796,N_6956);
nor U9597 (N_9597,N_7067,N_7096);
xor U9598 (N_9598,N_6476,N_7294);
nor U9599 (N_9599,N_7087,N_7207);
or U9600 (N_9600,N_6451,N_6809);
or U9601 (N_9601,N_6815,N_7402);
xor U9602 (N_9602,N_6612,N_7205);
nor U9603 (N_9603,N_6366,N_7648);
or U9604 (N_9604,N_6132,N_7609);
or U9605 (N_9605,N_6322,N_7597);
or U9606 (N_9606,N_6338,N_7050);
xor U9607 (N_9607,N_6954,N_7686);
nor U9608 (N_9608,N_7994,N_6560);
xnor U9609 (N_9609,N_7783,N_6761);
nand U9610 (N_9610,N_7464,N_7071);
nor U9611 (N_9611,N_7394,N_6595);
or U9612 (N_9612,N_7176,N_7068);
nor U9613 (N_9613,N_6125,N_7776);
and U9614 (N_9614,N_7443,N_7514);
and U9615 (N_9615,N_6823,N_7191);
or U9616 (N_9616,N_7533,N_6104);
nor U9617 (N_9617,N_6780,N_6760);
nor U9618 (N_9618,N_6721,N_7111);
nor U9619 (N_9619,N_6832,N_6502);
nor U9620 (N_9620,N_6885,N_6382);
nand U9621 (N_9621,N_6394,N_6098);
nand U9622 (N_9622,N_6711,N_6217);
nor U9623 (N_9623,N_7345,N_7245);
nor U9624 (N_9624,N_7531,N_7662);
nor U9625 (N_9625,N_7876,N_7196);
and U9626 (N_9626,N_6265,N_7549);
nand U9627 (N_9627,N_6425,N_6841);
nand U9628 (N_9628,N_7574,N_7320);
xnor U9629 (N_9629,N_7014,N_6922);
and U9630 (N_9630,N_7880,N_6834);
nor U9631 (N_9631,N_6531,N_6806);
and U9632 (N_9632,N_7696,N_7023);
or U9633 (N_9633,N_7050,N_7524);
nand U9634 (N_9634,N_6657,N_6426);
nor U9635 (N_9635,N_6714,N_6472);
nand U9636 (N_9636,N_7440,N_7371);
nor U9637 (N_9637,N_6146,N_6123);
or U9638 (N_9638,N_6675,N_6222);
and U9639 (N_9639,N_6847,N_7026);
or U9640 (N_9640,N_6167,N_7878);
or U9641 (N_9641,N_7052,N_7711);
nand U9642 (N_9642,N_7883,N_7695);
and U9643 (N_9643,N_7329,N_7970);
nor U9644 (N_9644,N_6186,N_7696);
nand U9645 (N_9645,N_6117,N_7071);
nor U9646 (N_9646,N_6431,N_6380);
and U9647 (N_9647,N_6861,N_7277);
nor U9648 (N_9648,N_7398,N_7331);
and U9649 (N_9649,N_7463,N_7551);
and U9650 (N_9650,N_6673,N_7842);
nor U9651 (N_9651,N_6119,N_7882);
or U9652 (N_9652,N_7717,N_6964);
nand U9653 (N_9653,N_7468,N_7391);
and U9654 (N_9654,N_6363,N_6722);
or U9655 (N_9655,N_7085,N_7364);
nand U9656 (N_9656,N_7612,N_7863);
nor U9657 (N_9657,N_6472,N_6697);
nand U9658 (N_9658,N_6048,N_7000);
and U9659 (N_9659,N_6628,N_6150);
and U9660 (N_9660,N_6062,N_6735);
xor U9661 (N_9661,N_7675,N_6551);
nand U9662 (N_9662,N_6558,N_7447);
nand U9663 (N_9663,N_7980,N_6056);
and U9664 (N_9664,N_6268,N_7284);
nor U9665 (N_9665,N_7457,N_6322);
nor U9666 (N_9666,N_6472,N_7588);
and U9667 (N_9667,N_6486,N_7767);
or U9668 (N_9668,N_7171,N_7199);
or U9669 (N_9669,N_6401,N_6929);
or U9670 (N_9670,N_7527,N_7946);
nand U9671 (N_9671,N_6021,N_7218);
and U9672 (N_9672,N_7415,N_7595);
and U9673 (N_9673,N_7133,N_6406);
or U9674 (N_9674,N_7721,N_6651);
nor U9675 (N_9675,N_6963,N_6725);
nand U9676 (N_9676,N_7963,N_6318);
nand U9677 (N_9677,N_7996,N_7709);
or U9678 (N_9678,N_6513,N_6637);
or U9679 (N_9679,N_7804,N_6473);
nand U9680 (N_9680,N_7558,N_6232);
and U9681 (N_9681,N_7017,N_7254);
nand U9682 (N_9682,N_7212,N_6594);
and U9683 (N_9683,N_7764,N_7822);
nor U9684 (N_9684,N_7094,N_7829);
and U9685 (N_9685,N_7209,N_7645);
nand U9686 (N_9686,N_7848,N_6555);
nor U9687 (N_9687,N_7685,N_6862);
nor U9688 (N_9688,N_6543,N_7893);
nand U9689 (N_9689,N_7922,N_7076);
or U9690 (N_9690,N_7616,N_6982);
nor U9691 (N_9691,N_6637,N_6491);
nor U9692 (N_9692,N_6280,N_6772);
xnor U9693 (N_9693,N_7351,N_7797);
and U9694 (N_9694,N_6546,N_6184);
nor U9695 (N_9695,N_7171,N_7838);
or U9696 (N_9696,N_6096,N_6430);
nand U9697 (N_9697,N_7595,N_7631);
xnor U9698 (N_9698,N_7771,N_6140);
or U9699 (N_9699,N_6326,N_6909);
or U9700 (N_9700,N_6966,N_7907);
and U9701 (N_9701,N_6624,N_7180);
and U9702 (N_9702,N_7540,N_6464);
and U9703 (N_9703,N_7262,N_7213);
and U9704 (N_9704,N_6429,N_6927);
nor U9705 (N_9705,N_6697,N_7393);
nor U9706 (N_9706,N_7727,N_6558);
and U9707 (N_9707,N_6059,N_6619);
and U9708 (N_9708,N_6947,N_7608);
nor U9709 (N_9709,N_6649,N_7072);
or U9710 (N_9710,N_7049,N_7411);
nand U9711 (N_9711,N_6718,N_7017);
and U9712 (N_9712,N_7429,N_7872);
nand U9713 (N_9713,N_7606,N_6054);
and U9714 (N_9714,N_6127,N_7081);
or U9715 (N_9715,N_7469,N_7132);
nand U9716 (N_9716,N_7729,N_7885);
and U9717 (N_9717,N_7208,N_6806);
and U9718 (N_9718,N_6112,N_7789);
or U9719 (N_9719,N_6405,N_6336);
and U9720 (N_9720,N_6001,N_6339);
or U9721 (N_9721,N_7608,N_6978);
xnor U9722 (N_9722,N_6750,N_6287);
nand U9723 (N_9723,N_6329,N_7753);
xnor U9724 (N_9724,N_6558,N_6705);
and U9725 (N_9725,N_6295,N_6032);
xor U9726 (N_9726,N_6850,N_7199);
nand U9727 (N_9727,N_7156,N_7296);
or U9728 (N_9728,N_6334,N_7015);
nor U9729 (N_9729,N_7744,N_6486);
nand U9730 (N_9730,N_7493,N_6098);
or U9731 (N_9731,N_7594,N_7194);
or U9732 (N_9732,N_6304,N_7847);
or U9733 (N_9733,N_7706,N_6511);
nand U9734 (N_9734,N_7764,N_6788);
or U9735 (N_9735,N_6403,N_7176);
and U9736 (N_9736,N_6207,N_7723);
and U9737 (N_9737,N_7377,N_6157);
nand U9738 (N_9738,N_6235,N_6447);
or U9739 (N_9739,N_6985,N_7628);
xnor U9740 (N_9740,N_7234,N_7920);
and U9741 (N_9741,N_6816,N_7512);
nand U9742 (N_9742,N_7540,N_7674);
nor U9743 (N_9743,N_7030,N_6298);
nand U9744 (N_9744,N_6589,N_6963);
xor U9745 (N_9745,N_6280,N_7221);
and U9746 (N_9746,N_6102,N_7868);
and U9747 (N_9747,N_7326,N_7518);
nor U9748 (N_9748,N_7421,N_7114);
and U9749 (N_9749,N_6911,N_6270);
xor U9750 (N_9750,N_7890,N_6521);
or U9751 (N_9751,N_6083,N_6698);
or U9752 (N_9752,N_7615,N_7591);
and U9753 (N_9753,N_7014,N_7914);
nor U9754 (N_9754,N_6245,N_7376);
nand U9755 (N_9755,N_6372,N_7189);
xor U9756 (N_9756,N_7066,N_6751);
nor U9757 (N_9757,N_6523,N_6431);
or U9758 (N_9758,N_7541,N_6846);
nor U9759 (N_9759,N_6947,N_7017);
and U9760 (N_9760,N_7260,N_6653);
and U9761 (N_9761,N_6013,N_6634);
or U9762 (N_9762,N_6958,N_6129);
nand U9763 (N_9763,N_7711,N_6323);
nor U9764 (N_9764,N_6417,N_7779);
nor U9765 (N_9765,N_7917,N_6822);
nor U9766 (N_9766,N_6708,N_7255);
and U9767 (N_9767,N_7509,N_6928);
nand U9768 (N_9768,N_7962,N_7983);
and U9769 (N_9769,N_6198,N_6958);
and U9770 (N_9770,N_7577,N_7442);
nor U9771 (N_9771,N_6709,N_7500);
and U9772 (N_9772,N_7699,N_7782);
and U9773 (N_9773,N_6523,N_7099);
nand U9774 (N_9774,N_7755,N_6749);
nor U9775 (N_9775,N_7876,N_7657);
or U9776 (N_9776,N_7266,N_6991);
nor U9777 (N_9777,N_7590,N_7078);
or U9778 (N_9778,N_7599,N_6906);
and U9779 (N_9779,N_7117,N_7596);
nand U9780 (N_9780,N_7339,N_6203);
nor U9781 (N_9781,N_7637,N_7070);
nand U9782 (N_9782,N_6509,N_7278);
and U9783 (N_9783,N_6533,N_6056);
nor U9784 (N_9784,N_6738,N_6800);
nand U9785 (N_9785,N_6645,N_7199);
or U9786 (N_9786,N_6886,N_6700);
xor U9787 (N_9787,N_7150,N_6216);
nor U9788 (N_9788,N_7163,N_6984);
and U9789 (N_9789,N_6682,N_7648);
nand U9790 (N_9790,N_6717,N_6209);
and U9791 (N_9791,N_6507,N_7754);
and U9792 (N_9792,N_7601,N_6356);
and U9793 (N_9793,N_6781,N_7617);
nand U9794 (N_9794,N_7101,N_6620);
nand U9795 (N_9795,N_6979,N_6291);
nor U9796 (N_9796,N_6181,N_6421);
and U9797 (N_9797,N_7926,N_6049);
nand U9798 (N_9798,N_6621,N_6271);
or U9799 (N_9799,N_6198,N_6996);
nor U9800 (N_9800,N_7192,N_6600);
xnor U9801 (N_9801,N_7831,N_7870);
and U9802 (N_9802,N_6381,N_7377);
and U9803 (N_9803,N_6977,N_7343);
nor U9804 (N_9804,N_6529,N_6628);
nand U9805 (N_9805,N_7524,N_7658);
nand U9806 (N_9806,N_6775,N_7183);
nand U9807 (N_9807,N_7654,N_7946);
nor U9808 (N_9808,N_7848,N_6131);
and U9809 (N_9809,N_6785,N_7542);
nor U9810 (N_9810,N_6474,N_6721);
nand U9811 (N_9811,N_6412,N_6096);
xor U9812 (N_9812,N_7104,N_6012);
nor U9813 (N_9813,N_6136,N_7801);
nor U9814 (N_9814,N_7349,N_6609);
and U9815 (N_9815,N_6011,N_6022);
or U9816 (N_9816,N_7167,N_7661);
and U9817 (N_9817,N_6187,N_7291);
and U9818 (N_9818,N_7487,N_6134);
or U9819 (N_9819,N_7027,N_7923);
nand U9820 (N_9820,N_6031,N_6392);
nand U9821 (N_9821,N_6034,N_6397);
or U9822 (N_9822,N_7889,N_7428);
and U9823 (N_9823,N_6443,N_6477);
and U9824 (N_9824,N_7490,N_6581);
or U9825 (N_9825,N_6828,N_7098);
nor U9826 (N_9826,N_7529,N_7471);
and U9827 (N_9827,N_6760,N_6705);
and U9828 (N_9828,N_7921,N_7302);
or U9829 (N_9829,N_6388,N_7499);
and U9830 (N_9830,N_6233,N_7455);
nand U9831 (N_9831,N_7508,N_7485);
nor U9832 (N_9832,N_7626,N_7820);
or U9833 (N_9833,N_7014,N_6016);
nor U9834 (N_9834,N_6636,N_6190);
or U9835 (N_9835,N_7064,N_7186);
nor U9836 (N_9836,N_6173,N_6573);
nand U9837 (N_9837,N_7671,N_6985);
or U9838 (N_9838,N_7880,N_6940);
or U9839 (N_9839,N_7150,N_7463);
nand U9840 (N_9840,N_6697,N_7987);
nor U9841 (N_9841,N_6969,N_7536);
nor U9842 (N_9842,N_6225,N_6158);
nor U9843 (N_9843,N_6573,N_7132);
or U9844 (N_9844,N_6597,N_7797);
and U9845 (N_9845,N_6173,N_6695);
nand U9846 (N_9846,N_6240,N_6777);
and U9847 (N_9847,N_6039,N_6134);
and U9848 (N_9848,N_6920,N_7602);
or U9849 (N_9849,N_7417,N_7426);
xor U9850 (N_9850,N_7726,N_6953);
nand U9851 (N_9851,N_7227,N_6276);
and U9852 (N_9852,N_6819,N_6983);
and U9853 (N_9853,N_7861,N_6153);
nand U9854 (N_9854,N_7525,N_7367);
xnor U9855 (N_9855,N_7987,N_6829);
xnor U9856 (N_9856,N_6680,N_6337);
or U9857 (N_9857,N_7765,N_6088);
or U9858 (N_9858,N_7051,N_6192);
nand U9859 (N_9859,N_7471,N_6239);
nand U9860 (N_9860,N_6630,N_6633);
and U9861 (N_9861,N_6284,N_7238);
or U9862 (N_9862,N_6317,N_6554);
and U9863 (N_9863,N_6591,N_6303);
nand U9864 (N_9864,N_6406,N_7560);
nand U9865 (N_9865,N_6825,N_6282);
nor U9866 (N_9866,N_7570,N_6699);
or U9867 (N_9867,N_6184,N_6485);
nor U9868 (N_9868,N_6018,N_7473);
and U9869 (N_9869,N_7678,N_7399);
nor U9870 (N_9870,N_7450,N_7920);
nor U9871 (N_9871,N_6153,N_6290);
nor U9872 (N_9872,N_6191,N_6621);
nor U9873 (N_9873,N_7514,N_6502);
nand U9874 (N_9874,N_6509,N_7861);
nand U9875 (N_9875,N_6754,N_7229);
or U9876 (N_9876,N_6877,N_7089);
nand U9877 (N_9877,N_6286,N_7461);
or U9878 (N_9878,N_7796,N_6960);
nand U9879 (N_9879,N_6863,N_7531);
and U9880 (N_9880,N_6704,N_6282);
xnor U9881 (N_9881,N_6923,N_6813);
and U9882 (N_9882,N_7963,N_7339);
xnor U9883 (N_9883,N_7296,N_7553);
nand U9884 (N_9884,N_6175,N_7042);
nor U9885 (N_9885,N_6057,N_7976);
nand U9886 (N_9886,N_7299,N_6509);
or U9887 (N_9887,N_6846,N_6761);
nor U9888 (N_9888,N_7818,N_7293);
and U9889 (N_9889,N_6166,N_6192);
nand U9890 (N_9890,N_7138,N_6297);
nand U9891 (N_9891,N_7167,N_6077);
or U9892 (N_9892,N_7167,N_7357);
or U9893 (N_9893,N_6981,N_6540);
nor U9894 (N_9894,N_6242,N_7056);
or U9895 (N_9895,N_6624,N_7674);
or U9896 (N_9896,N_7965,N_6500);
nor U9897 (N_9897,N_7485,N_7091);
xnor U9898 (N_9898,N_6837,N_6636);
or U9899 (N_9899,N_7714,N_6814);
nand U9900 (N_9900,N_6681,N_7999);
or U9901 (N_9901,N_6331,N_6056);
and U9902 (N_9902,N_7230,N_6569);
or U9903 (N_9903,N_7327,N_7504);
and U9904 (N_9904,N_6640,N_7287);
and U9905 (N_9905,N_6179,N_6419);
or U9906 (N_9906,N_7992,N_6509);
nor U9907 (N_9907,N_6417,N_6285);
xnor U9908 (N_9908,N_7336,N_7013);
nand U9909 (N_9909,N_6650,N_7095);
xnor U9910 (N_9910,N_7498,N_7765);
or U9911 (N_9911,N_7943,N_6631);
xor U9912 (N_9912,N_7430,N_6969);
xor U9913 (N_9913,N_6469,N_6126);
or U9914 (N_9914,N_7193,N_6393);
nor U9915 (N_9915,N_6984,N_6514);
or U9916 (N_9916,N_7488,N_6233);
nor U9917 (N_9917,N_6507,N_6815);
nor U9918 (N_9918,N_7421,N_6265);
and U9919 (N_9919,N_6563,N_7275);
nand U9920 (N_9920,N_7161,N_7819);
and U9921 (N_9921,N_7187,N_6125);
nor U9922 (N_9922,N_6419,N_7479);
nor U9923 (N_9923,N_7024,N_7430);
nor U9924 (N_9924,N_6582,N_7926);
and U9925 (N_9925,N_7984,N_7504);
and U9926 (N_9926,N_7660,N_6335);
nand U9927 (N_9927,N_6066,N_6751);
nor U9928 (N_9928,N_7699,N_6827);
or U9929 (N_9929,N_7171,N_7373);
or U9930 (N_9930,N_6101,N_6342);
nand U9931 (N_9931,N_7292,N_6871);
nor U9932 (N_9932,N_6030,N_6987);
nor U9933 (N_9933,N_7977,N_7464);
or U9934 (N_9934,N_6456,N_6537);
xor U9935 (N_9935,N_7378,N_6995);
xor U9936 (N_9936,N_7392,N_6159);
and U9937 (N_9937,N_7477,N_6091);
xnor U9938 (N_9938,N_6714,N_6796);
nor U9939 (N_9939,N_6486,N_7216);
nand U9940 (N_9940,N_7928,N_6788);
nand U9941 (N_9941,N_7657,N_6952);
nor U9942 (N_9942,N_6440,N_7009);
xnor U9943 (N_9943,N_6398,N_7153);
and U9944 (N_9944,N_7774,N_7265);
or U9945 (N_9945,N_6708,N_6429);
nor U9946 (N_9946,N_7301,N_7946);
nand U9947 (N_9947,N_7118,N_6733);
or U9948 (N_9948,N_7356,N_7811);
and U9949 (N_9949,N_7282,N_6085);
and U9950 (N_9950,N_6725,N_7210);
or U9951 (N_9951,N_6400,N_6531);
or U9952 (N_9952,N_7603,N_6262);
nand U9953 (N_9953,N_7776,N_6350);
nor U9954 (N_9954,N_6366,N_6342);
or U9955 (N_9955,N_7710,N_7497);
nand U9956 (N_9956,N_6603,N_6857);
nor U9957 (N_9957,N_6636,N_6618);
nor U9958 (N_9958,N_6814,N_7713);
xnor U9959 (N_9959,N_6088,N_6113);
or U9960 (N_9960,N_6417,N_6963);
nand U9961 (N_9961,N_6620,N_7060);
or U9962 (N_9962,N_7841,N_7118);
or U9963 (N_9963,N_7031,N_7849);
and U9964 (N_9964,N_7337,N_6168);
and U9965 (N_9965,N_6144,N_6283);
nand U9966 (N_9966,N_7696,N_6249);
nor U9967 (N_9967,N_6401,N_7509);
nand U9968 (N_9968,N_7734,N_6104);
or U9969 (N_9969,N_7707,N_6025);
nor U9970 (N_9970,N_6765,N_7484);
or U9971 (N_9971,N_6212,N_7177);
or U9972 (N_9972,N_6413,N_6352);
nand U9973 (N_9973,N_7323,N_7236);
nor U9974 (N_9974,N_7023,N_6887);
nand U9975 (N_9975,N_7635,N_7302);
or U9976 (N_9976,N_6214,N_6640);
nor U9977 (N_9977,N_6652,N_6854);
and U9978 (N_9978,N_6178,N_6601);
nand U9979 (N_9979,N_7182,N_7333);
xnor U9980 (N_9980,N_6724,N_7699);
nor U9981 (N_9981,N_7549,N_6011);
and U9982 (N_9982,N_7045,N_7162);
or U9983 (N_9983,N_7080,N_7573);
nor U9984 (N_9984,N_7756,N_6025);
xnor U9985 (N_9985,N_7598,N_6491);
and U9986 (N_9986,N_6415,N_6582);
and U9987 (N_9987,N_7998,N_6219);
or U9988 (N_9988,N_7626,N_7679);
nor U9989 (N_9989,N_6721,N_7535);
or U9990 (N_9990,N_7823,N_6091);
and U9991 (N_9991,N_6393,N_7874);
or U9992 (N_9992,N_7554,N_7751);
and U9993 (N_9993,N_7788,N_7236);
and U9994 (N_9994,N_7385,N_7857);
xor U9995 (N_9995,N_6431,N_6444);
nor U9996 (N_9996,N_7660,N_7391);
nand U9997 (N_9997,N_6113,N_7281);
or U9998 (N_9998,N_6007,N_6188);
nor U9999 (N_9999,N_6850,N_6164);
or U10000 (N_10000,N_8466,N_9333);
and U10001 (N_10001,N_8914,N_9005);
or U10002 (N_10002,N_9352,N_8637);
or U10003 (N_10003,N_9674,N_9868);
and U10004 (N_10004,N_9736,N_9617);
nor U10005 (N_10005,N_8190,N_8895);
or U10006 (N_10006,N_8715,N_8530);
nor U10007 (N_10007,N_8857,N_8900);
xor U10008 (N_10008,N_9864,N_9412);
nand U10009 (N_10009,N_8350,N_9320);
nand U10010 (N_10010,N_9407,N_8633);
nor U10011 (N_10011,N_8226,N_8000);
and U10012 (N_10012,N_8956,N_9162);
nand U10013 (N_10013,N_9874,N_8219);
or U10014 (N_10014,N_8120,N_9022);
xor U10015 (N_10015,N_8459,N_9664);
nor U10016 (N_10016,N_9002,N_8709);
or U10017 (N_10017,N_9156,N_8811);
and U10018 (N_10018,N_8400,N_9512);
nor U10019 (N_10019,N_9823,N_9479);
nand U10020 (N_10020,N_8996,N_8052);
or U10021 (N_10021,N_8985,N_8882);
or U10022 (N_10022,N_8818,N_9188);
and U10023 (N_10023,N_9871,N_8273);
and U10024 (N_10024,N_8886,N_8305);
or U10025 (N_10025,N_9701,N_9645);
nor U10026 (N_10026,N_9178,N_9014);
nor U10027 (N_10027,N_8366,N_9458);
or U10028 (N_10028,N_9265,N_9679);
or U10029 (N_10029,N_9263,N_9249);
nor U10030 (N_10030,N_9023,N_8789);
nor U10031 (N_10031,N_9060,N_9754);
nand U10032 (N_10032,N_8940,N_9238);
nand U10033 (N_10033,N_8370,N_9579);
and U10034 (N_10034,N_9834,N_9116);
and U10035 (N_10035,N_9291,N_9201);
nand U10036 (N_10036,N_8583,N_8840);
nand U10037 (N_10037,N_8127,N_8581);
and U10038 (N_10038,N_8729,N_8511);
and U10039 (N_10039,N_9184,N_8240);
nor U10040 (N_10040,N_8638,N_8510);
nor U10041 (N_10041,N_9809,N_8907);
or U10042 (N_10042,N_9563,N_9132);
and U10043 (N_10043,N_8184,N_8780);
nor U10044 (N_10044,N_9386,N_9801);
nand U10045 (N_10045,N_8391,N_8905);
and U10046 (N_10046,N_9878,N_9015);
nand U10047 (N_10047,N_8666,N_9665);
nand U10048 (N_10048,N_8041,N_8734);
xor U10049 (N_10049,N_9362,N_8997);
or U10050 (N_10050,N_8721,N_9280);
or U10051 (N_10051,N_9897,N_8233);
or U10052 (N_10052,N_8185,N_8093);
nor U10053 (N_10053,N_9328,N_9727);
or U10054 (N_10054,N_9428,N_8106);
or U10055 (N_10055,N_9444,N_9947);
nand U10056 (N_10056,N_8627,N_8977);
nor U10057 (N_10057,N_8222,N_9271);
nor U10058 (N_10058,N_8536,N_9840);
xnor U10059 (N_10059,N_9237,N_9297);
nor U10060 (N_10060,N_9854,N_9551);
xor U10061 (N_10061,N_9507,N_8778);
nor U10062 (N_10062,N_8471,N_8213);
nand U10063 (N_10063,N_8469,N_9949);
nand U10064 (N_10064,N_8053,N_9142);
nand U10065 (N_10065,N_8606,N_9626);
or U10066 (N_10066,N_9472,N_9715);
nor U10067 (N_10067,N_8991,N_8097);
and U10068 (N_10068,N_8896,N_9267);
or U10069 (N_10069,N_9991,N_8681);
nand U10070 (N_10070,N_9114,N_9985);
nor U10071 (N_10071,N_8232,N_8569);
xor U10072 (N_10072,N_8557,N_8060);
nor U10073 (N_10073,N_8340,N_9518);
and U10074 (N_10074,N_9079,N_8790);
xnor U10075 (N_10075,N_8989,N_9601);
or U10076 (N_10076,N_8570,N_9627);
and U10077 (N_10077,N_8188,N_8292);
and U10078 (N_10078,N_8519,N_8328);
or U10079 (N_10079,N_8777,N_8533);
nand U10080 (N_10080,N_9516,N_9223);
and U10081 (N_10081,N_9374,N_8373);
or U10082 (N_10082,N_8458,N_9403);
or U10083 (N_10083,N_8864,N_8480);
nand U10084 (N_10084,N_9668,N_9343);
or U10085 (N_10085,N_9911,N_9028);
and U10086 (N_10086,N_9347,N_9281);
and U10087 (N_10087,N_9851,N_8057);
and U10088 (N_10088,N_8877,N_8664);
nand U10089 (N_10089,N_9102,N_8594);
nor U10090 (N_10090,N_9568,N_9196);
or U10091 (N_10091,N_8786,N_8412);
xnor U10092 (N_10092,N_9647,N_8943);
and U10093 (N_10093,N_8794,N_9167);
nor U10094 (N_10094,N_9490,N_8971);
nand U10095 (N_10095,N_8700,N_9545);
nor U10096 (N_10096,N_8033,N_9327);
nor U10097 (N_10097,N_8140,N_9717);
or U10098 (N_10098,N_9232,N_8279);
nor U10099 (N_10099,N_8839,N_9597);
nor U10100 (N_10100,N_9211,N_9027);
nor U10101 (N_10101,N_8083,N_8548);
and U10102 (N_10102,N_9073,N_9961);
or U10103 (N_10103,N_9445,N_9559);
nor U10104 (N_10104,N_8830,N_8084);
nand U10105 (N_10105,N_8532,N_8356);
nand U10106 (N_10106,N_8756,N_9103);
or U10107 (N_10107,N_8441,N_9847);
or U10108 (N_10108,N_8755,N_8555);
and U10109 (N_10109,N_9222,N_8516);
or U10110 (N_10110,N_8175,N_8523);
or U10111 (N_10111,N_9760,N_9973);
and U10112 (N_10112,N_8159,N_9824);
xnor U10113 (N_10113,N_9540,N_8887);
xor U10114 (N_10114,N_9471,N_8793);
xnor U10115 (N_10115,N_8652,N_8976);
nor U10116 (N_10116,N_8559,N_8449);
nor U10117 (N_10117,N_8211,N_8810);
or U10118 (N_10118,N_8298,N_8157);
and U10119 (N_10119,N_9951,N_8270);
nor U10120 (N_10120,N_8168,N_9025);
nand U10121 (N_10121,N_8113,N_9181);
nand U10122 (N_10122,N_9318,N_9159);
nand U10123 (N_10123,N_8856,N_8595);
or U10124 (N_10124,N_8092,N_8915);
nor U10125 (N_10125,N_8932,N_8126);
or U10126 (N_10126,N_9887,N_8263);
nor U10127 (N_10127,N_9999,N_8284);
and U10128 (N_10128,N_8043,N_8472);
nor U10129 (N_10129,N_8927,N_8164);
nor U10130 (N_10130,N_8309,N_9606);
xor U10131 (N_10131,N_9534,N_9240);
nor U10132 (N_10132,N_9530,N_9946);
and U10133 (N_10133,N_9192,N_9261);
nor U10134 (N_10134,N_9622,N_9278);
nand U10135 (N_10135,N_8754,N_8901);
and U10136 (N_10136,N_9963,N_8906);
or U10137 (N_10137,N_9870,N_9165);
nor U10138 (N_10138,N_9144,N_8607);
and U10139 (N_10139,N_9976,N_9933);
nand U10140 (N_10140,N_9554,N_8771);
or U10141 (N_10141,N_9221,N_8100);
or U10142 (N_10142,N_8401,N_8359);
or U10143 (N_10143,N_8911,N_9924);
and U10144 (N_10144,N_9570,N_8908);
nand U10145 (N_10145,N_9058,N_9348);
xnor U10146 (N_10146,N_8040,N_8386);
nor U10147 (N_10147,N_9774,N_9344);
nor U10148 (N_10148,N_8757,N_8275);
and U10149 (N_10149,N_9312,N_9276);
nand U10150 (N_10150,N_8880,N_9409);
or U10151 (N_10151,N_9244,N_8266);
or U10152 (N_10152,N_8621,N_8416);
nand U10153 (N_10153,N_9171,N_8702);
or U10154 (N_10154,N_8950,N_9743);
and U10155 (N_10155,N_9372,N_9885);
and U10156 (N_10156,N_8728,N_8134);
nor U10157 (N_10157,N_9105,N_9186);
xnor U10158 (N_10158,N_9879,N_9842);
nor U10159 (N_10159,N_9299,N_9898);
nor U10160 (N_10160,N_8828,N_9705);
nor U10161 (N_10161,N_9069,N_9431);
and U10162 (N_10162,N_8545,N_8525);
or U10163 (N_10163,N_9293,N_9164);
or U10164 (N_10164,N_8264,N_9163);
or U10165 (N_10165,N_8885,N_9836);
nor U10166 (N_10166,N_8236,N_8220);
and U10167 (N_10167,N_8520,N_9972);
and U10168 (N_10168,N_8925,N_9654);
and U10169 (N_10169,N_9245,N_9199);
or U10170 (N_10170,N_8325,N_9535);
nor U10171 (N_10171,N_8930,N_9363);
or U10172 (N_10172,N_8549,N_9389);
or U10173 (N_10173,N_9179,N_9618);
nand U10174 (N_10174,N_8749,N_8751);
nor U10175 (N_10175,N_8972,N_8128);
nor U10176 (N_10176,N_9086,N_8640);
xnor U10177 (N_10177,N_9867,N_8390);
and U10178 (N_10178,N_8645,N_8868);
nand U10179 (N_10179,N_8936,N_8389);
and U10180 (N_10180,N_9738,N_8858);
or U10181 (N_10181,N_8020,N_9382);
nand U10182 (N_10182,N_8217,N_9331);
xnor U10183 (N_10183,N_9751,N_8429);
nor U10184 (N_10184,N_9942,N_8542);
nand U10185 (N_10185,N_8941,N_8180);
or U10186 (N_10186,N_9302,N_8518);
or U10187 (N_10187,N_8091,N_9752);
and U10188 (N_10188,N_8393,N_9408);
nand U10189 (N_10189,N_9477,N_8149);
nor U10190 (N_10190,N_9578,N_8626);
xor U10191 (N_10191,N_8625,N_8740);
or U10192 (N_10192,N_9140,N_8723);
and U10193 (N_10193,N_8503,N_8738);
and U10194 (N_10194,N_8920,N_9706);
and U10195 (N_10195,N_9430,N_9604);
xor U10196 (N_10196,N_9649,N_9906);
nor U10197 (N_10197,N_9848,N_9543);
nand U10198 (N_10198,N_8028,N_8307);
nor U10199 (N_10199,N_9149,N_8618);
nand U10200 (N_10200,N_9643,N_9183);
xor U10201 (N_10201,N_8602,N_9709);
nand U10202 (N_10202,N_8296,N_9741);
nor U10203 (N_10203,N_9029,N_9794);
xnor U10204 (N_10204,N_9776,N_8587);
or U10205 (N_10205,N_9173,N_9236);
nand U10206 (N_10206,N_8812,N_9620);
or U10207 (N_10207,N_9459,N_8584);
nand U10208 (N_10208,N_9599,N_9100);
and U10209 (N_10209,N_9255,N_9273);
and U10210 (N_10210,N_8062,N_8726);
or U10211 (N_10211,N_9960,N_8506);
nor U10212 (N_10212,N_9035,N_8687);
nor U10213 (N_10213,N_9903,N_8805);
nor U10214 (N_10214,N_9080,N_9537);
xor U10215 (N_10215,N_9126,N_8775);
nand U10216 (N_10216,N_8342,N_8639);
nor U10217 (N_10217,N_8833,N_8330);
or U10218 (N_10218,N_8678,N_8246);
xnor U10219 (N_10219,N_8365,N_9585);
nand U10220 (N_10220,N_9084,N_9763);
and U10221 (N_10221,N_8172,N_8966);
and U10222 (N_10222,N_9364,N_8817);
nor U10223 (N_10223,N_9541,N_9737);
nand U10224 (N_10224,N_8538,N_8317);
or U10225 (N_10225,N_9764,N_9688);
xnor U10226 (N_10226,N_9502,N_9909);
nor U10227 (N_10227,N_9912,N_8438);
or U10228 (N_10228,N_8135,N_8277);
nor U10229 (N_10229,N_8013,N_9595);
or U10230 (N_10230,N_9120,N_8623);
xor U10231 (N_10231,N_9673,N_9215);
or U10232 (N_10232,N_9111,N_9556);
nor U10233 (N_10233,N_9650,N_8029);
and U10234 (N_10234,N_8380,N_9208);
or U10235 (N_10235,N_9136,N_9243);
or U10236 (N_10236,N_8144,N_8482);
and U10237 (N_10237,N_9756,N_8661);
or U10238 (N_10238,N_9254,N_9075);
nor U10239 (N_10239,N_9460,N_8066);
and U10240 (N_10240,N_8762,N_9234);
or U10241 (N_10241,N_8884,N_9155);
and U10242 (N_10242,N_8448,N_9509);
nor U10243 (N_10243,N_9708,N_8613);
xnor U10244 (N_10244,N_8192,N_8614);
nand U10245 (N_10245,N_9786,N_8069);
xor U10246 (N_10246,N_8216,N_9306);
nand U10247 (N_10247,N_8862,N_9804);
nand U10248 (N_10248,N_9761,N_9695);
and U10249 (N_10249,N_8674,N_9499);
nand U10250 (N_10250,N_9603,N_8826);
and U10251 (N_10251,N_8848,N_8362);
or U10252 (N_10252,N_9390,N_9839);
nand U10253 (N_10253,N_8081,N_9217);
or U10254 (N_10254,N_8321,N_8339);
or U10255 (N_10255,N_8924,N_9807);
and U10256 (N_10256,N_9505,N_8115);
nand U10257 (N_10257,N_9910,N_9613);
nand U10258 (N_10258,N_9825,N_9977);
or U10259 (N_10259,N_9154,N_8680);
and U10260 (N_10260,N_8513,N_9307);
and U10261 (N_10261,N_8122,N_9124);
xnor U10262 (N_10262,N_9553,N_8038);
and U10263 (N_10263,N_8508,N_8892);
nor U10264 (N_10264,N_9623,N_9883);
and U10265 (N_10265,N_8163,N_8108);
nand U10266 (N_10266,N_8688,N_9091);
xor U10267 (N_10267,N_8061,N_9335);
nor U10268 (N_10268,N_8938,N_9896);
nand U10269 (N_10269,N_8692,N_9135);
nor U10270 (N_10270,N_9815,N_9197);
nand U10271 (N_10271,N_8801,N_9571);
xnor U10272 (N_10272,N_9264,N_8564);
nor U10273 (N_10273,N_8679,N_9796);
nor U10274 (N_10274,N_9956,N_8011);
or U10275 (N_10275,N_9117,N_8620);
nor U10276 (N_10276,N_9224,N_9104);
nor U10277 (N_10277,N_8733,N_9852);
and U10278 (N_10278,N_9855,N_8944);
or U10279 (N_10279,N_9078,N_9448);
and U10280 (N_10280,N_8854,N_8758);
nand U10281 (N_10281,N_8629,N_8921);
nor U10282 (N_10282,N_9063,N_8411);
or U10283 (N_10283,N_9675,N_8369);
nand U10284 (N_10284,N_9365,N_8478);
and U10285 (N_10285,N_8334,N_9371);
nand U10286 (N_10286,N_9097,N_9151);
and U10287 (N_10287,N_8306,N_8834);
and U10288 (N_10288,N_9630,N_9475);
or U10289 (N_10289,N_9316,N_8962);
xor U10290 (N_10290,N_9369,N_8059);
xnor U10291 (N_10291,N_9575,N_9228);
or U10292 (N_10292,N_8894,N_8204);
or U10293 (N_10293,N_8257,N_9997);
or U10294 (N_10294,N_9833,N_8909);
nand U10295 (N_10295,N_8417,N_8435);
nor U10296 (N_10296,N_9742,N_8054);
nor U10297 (N_10297,N_8912,N_9773);
nor U10298 (N_10298,N_8860,N_8430);
or U10299 (N_10299,N_9993,N_9076);
nand U10300 (N_10300,N_8974,N_9146);
or U10301 (N_10301,N_8312,N_8413);
nor U10302 (N_10302,N_9957,N_8443);
nor U10303 (N_10303,N_8580,N_9054);
nor U10304 (N_10304,N_9783,N_8212);
or U10305 (N_10305,N_9268,N_9336);
or U10306 (N_10306,N_8014,N_8933);
or U10307 (N_10307,N_8781,N_8016);
and U10308 (N_10308,N_9515,N_8524);
nand U10309 (N_10309,N_8194,N_9123);
nand U10310 (N_10310,N_8803,N_8546);
or U10311 (N_10311,N_9533,N_9048);
and U10312 (N_10312,N_9806,N_9158);
nand U10313 (N_10313,N_9095,N_8474);
nor U10314 (N_10314,N_8836,N_9388);
and U10315 (N_10315,N_8104,N_9990);
nand U10316 (N_10316,N_8865,N_8765);
or U10317 (N_10317,N_9770,N_9766);
xnor U10318 (N_10318,N_8540,N_8590);
or U10319 (N_10319,N_9865,N_8039);
and U10320 (N_10320,N_8197,N_8782);
nor U10321 (N_10321,N_9006,N_8165);
nand U10322 (N_10322,N_9681,N_9353);
nand U10323 (N_10323,N_9857,N_8156);
nor U10324 (N_10324,N_8406,N_8318);
nand U10325 (N_10325,N_8913,N_8042);
nand U10326 (N_10326,N_8534,N_9041);
nand U10327 (N_10327,N_9932,N_8207);
nand U10328 (N_10328,N_8005,N_9676);
nor U10329 (N_10329,N_8155,N_8179);
xnor U10330 (N_10330,N_8761,N_9303);
nor U10331 (N_10331,N_9292,N_9648);
and U10332 (N_10332,N_8671,N_8783);
and U10333 (N_10333,N_8125,N_9713);
or U10334 (N_10334,N_8931,N_8667);
nor U10335 (N_10335,N_8703,N_8599);
nand U10336 (N_10336,N_9587,N_9661);
nand U10337 (N_10337,N_8415,N_9133);
nor U10338 (N_10338,N_8952,N_8988);
or U10339 (N_10339,N_8842,N_8252);
nand U10340 (N_10340,N_9446,N_8034);
xnor U10341 (N_10341,N_9888,N_9295);
or U10342 (N_10342,N_8121,N_9394);
nand U10343 (N_10343,N_8048,N_9907);
nand U10344 (N_10344,N_9231,N_8716);
or U10345 (N_10345,N_8310,N_9050);
or U10346 (N_10346,N_9889,N_9979);
nor U10347 (N_10347,N_9758,N_8665);
and U10348 (N_10348,N_9747,N_8566);
nand U10349 (N_10349,N_8816,N_8874);
nor U10350 (N_10350,N_8424,N_9734);
nand U10351 (N_10351,N_9227,N_8183);
and U10352 (N_10352,N_8451,N_8012);
nand U10353 (N_10353,N_9939,N_8923);
and U10354 (N_10354,N_8653,N_8947);
and U10355 (N_10355,N_8145,N_9663);
nand U10356 (N_10356,N_8684,N_9844);
nor U10357 (N_10357,N_8300,N_9434);
xor U10358 (N_10358,N_9229,N_8278);
and U10359 (N_10359,N_9187,N_8398);
and U10360 (N_10360,N_8436,N_8281);
nand U10361 (N_10361,N_9427,N_8837);
nor U10362 (N_10362,N_9150,N_8396);
and U10363 (N_10363,N_8597,N_9121);
or U10364 (N_10364,N_9449,N_9829);
nor U10365 (N_10365,N_8831,N_8133);
nand U10366 (N_10366,N_9966,N_9762);
xnor U10367 (N_10367,N_9077,N_9241);
or U10368 (N_10368,N_9089,N_9677);
nand U10369 (N_10369,N_8249,N_9826);
nand U10370 (N_10370,N_8870,N_8274);
xnor U10371 (N_10371,N_8654,N_9740);
nor U10372 (N_10372,N_8426,N_9748);
nor U10373 (N_10373,N_9367,N_8644);
nand U10374 (N_10374,N_8158,N_9658);
and U10375 (N_10375,N_9420,N_8802);
and U10376 (N_10376,N_9088,N_8067);
and U10377 (N_10377,N_8089,N_9811);
or U10378 (N_10378,N_9441,N_9433);
and U10379 (N_10379,N_9191,N_9672);
nand U10380 (N_10380,N_8182,N_8804);
nand U10381 (N_10381,N_9242,N_9180);
nor U10382 (N_10382,N_8036,N_9719);
and U10383 (N_10383,N_8821,N_8313);
nand U10384 (N_10384,N_8747,N_8576);
nor U10385 (N_10385,N_8918,N_9656);
and U10386 (N_10386,N_8418,N_9980);
and U10387 (N_10387,N_9329,N_9732);
nand U10388 (N_10388,N_8772,N_8187);
nand U10389 (N_10389,N_9691,N_9454);
nand U10390 (N_10390,N_8460,N_8431);
nand U10391 (N_10391,N_8551,N_9784);
nor U10392 (N_10392,N_9426,N_9489);
nand U10393 (N_10393,N_9964,N_8405);
nor U10394 (N_10394,N_9219,N_8586);
nand U10395 (N_10395,N_9657,N_9629);
and U10396 (N_10396,N_9926,N_9612);
or U10397 (N_10397,N_8302,N_9061);
and U10398 (N_10398,N_8792,N_8208);
or U10399 (N_10399,N_8229,N_9831);
and U10400 (N_10400,N_8191,N_8642);
or U10401 (N_10401,N_8319,N_9724);
nor U10402 (N_10402,N_8254,N_8528);
nor U10403 (N_10403,N_9381,N_9652);
nor U10404 (N_10404,N_8676,N_9845);
nor U10405 (N_10405,N_9262,N_9904);
or U10406 (N_10406,N_9875,N_8922);
or U10407 (N_10407,N_9712,N_9166);
nand U10408 (N_10408,N_9416,N_8628);
and U10409 (N_10409,N_8859,N_8883);
and U10410 (N_10410,N_8779,N_9510);
nand U10411 (N_10411,N_8507,N_8027);
nand U10412 (N_10412,N_8078,N_9799);
nor U10413 (N_10413,N_8727,N_9493);
nor U10414 (N_10414,N_9821,N_8718);
and U10415 (N_10415,N_9378,N_9049);
and U10416 (N_10416,N_9203,N_8707);
or U10417 (N_10417,N_9918,N_8492);
nor U10418 (N_10418,N_8759,N_9660);
and U10419 (N_10419,N_9600,N_9813);
or U10420 (N_10420,N_9418,N_8673);
nor U10421 (N_10421,N_8588,N_8730);
xor U10422 (N_10422,N_9860,N_8440);
nor U10423 (N_10423,N_9682,N_8221);
and U10424 (N_10424,N_9018,N_9375);
xnor U10425 (N_10425,N_9368,N_9250);
and U10426 (N_10426,N_9891,N_8314);
and U10427 (N_10427,N_9992,N_9480);
and U10428 (N_10428,N_9359,N_9198);
nor U10429 (N_10429,N_8953,N_9702);
or U10430 (N_10430,N_8617,N_9220);
xnor U10431 (N_10431,N_9781,N_8351);
or U10432 (N_10432,N_8049,N_9283);
nand U10433 (N_10433,N_8682,N_9611);
nor U10434 (N_10434,N_8669,N_9465);
or U10435 (N_10435,N_8420,N_9300);
nor U10436 (N_10436,N_9859,N_8631);
nor U10437 (N_10437,N_8297,N_9286);
xor U10438 (N_10438,N_8161,N_9846);
and U10439 (N_10439,N_9216,N_9632);
or U10440 (N_10440,N_9012,N_9436);
nor U10441 (N_10441,N_8820,N_8376);
nand U10442 (N_10442,N_9131,N_8479);
or U10443 (N_10443,N_8237,N_8711);
nand U10444 (N_10444,N_9108,N_9772);
nand U10445 (N_10445,N_8822,N_8946);
xnor U10446 (N_10446,N_8979,N_8465);
nor U10447 (N_10447,N_9731,N_8395);
nor U10448 (N_10448,N_9404,N_9659);
nand U10449 (N_10449,N_9750,N_9323);
and U10450 (N_10450,N_8009,N_8798);
nand U10451 (N_10451,N_8129,N_8486);
or U10452 (N_10452,N_9621,N_9550);
nor U10453 (N_10453,N_9536,N_8539);
or U10454 (N_10454,N_9145,N_8589);
and U10455 (N_10455,N_9042,N_8869);
or U10456 (N_10456,N_9009,N_8402);
nor U10457 (N_10457,N_8535,N_8928);
or U10458 (N_10458,N_8142,N_8970);
nor U10459 (N_10459,N_8659,N_9795);
and U10460 (N_10460,N_8898,N_9596);
and U10461 (N_10461,N_9487,N_9152);
nor U10462 (N_10462,N_8147,N_9099);
and U10463 (N_10463,N_9314,N_8743);
and U10464 (N_10464,N_9143,N_8693);
and U10465 (N_10465,N_8999,N_9780);
nand U10466 (N_10466,N_9342,N_9213);
nor U10467 (N_10467,N_9256,N_9539);
nand U10468 (N_10468,N_9561,N_9608);
and U10469 (N_10469,N_9437,N_9830);
nand U10470 (N_10470,N_9130,N_9351);
nand U10471 (N_10471,N_9863,N_9856);
nand U10472 (N_10472,N_8295,N_9771);
nor U10473 (N_10473,N_8578,N_8713);
nor U10474 (N_10474,N_8732,N_9483);
nor U10475 (N_10475,N_9415,N_9233);
nand U10476 (N_10476,N_8209,N_8648);
nor U10477 (N_10477,N_9319,N_8967);
nand U10478 (N_10478,N_8919,N_9440);
nand U10479 (N_10479,N_9443,N_9817);
and U10480 (N_10480,N_8283,N_8004);
nand U10481 (N_10481,N_8099,N_8769);
xor U10482 (N_10482,N_8082,N_8017);
nand U10483 (N_10483,N_8259,N_8235);
or U10484 (N_10484,N_8572,N_9514);
nor U10485 (N_10485,N_9744,N_8643);
nand U10486 (N_10486,N_8591,N_8178);
and U10487 (N_10487,N_8473,N_9670);
nor U10488 (N_10488,N_8672,N_8464);
nand U10489 (N_10489,N_9628,N_9040);
nand U10490 (N_10490,N_8035,N_8963);
nand U10491 (N_10491,N_9619,N_8177);
or U10492 (N_10492,N_8090,N_8799);
nand U10493 (N_10493,N_8752,N_8800);
or U10494 (N_10494,N_9200,N_8787);
and U10495 (N_10495,N_9631,N_8095);
nand U10496 (N_10496,N_9730,N_8360);
and U10497 (N_10497,N_9853,N_9838);
nand U10498 (N_10498,N_8897,N_9927);
nand U10499 (N_10499,N_9697,N_8748);
nor U10500 (N_10500,N_9112,N_9759);
xor U10501 (N_10501,N_8600,N_9728);
or U10502 (N_10502,N_9057,N_9066);
or U10503 (N_10503,N_8153,N_9392);
or U10504 (N_10504,N_9513,N_9189);
or U10505 (N_10505,N_8024,N_9739);
and U10506 (N_10506,N_8452,N_9204);
xnor U10507 (N_10507,N_8047,N_8851);
and U10508 (N_10508,N_8556,N_9016);
nor U10509 (N_10509,N_8073,N_8008);
and U10510 (N_10510,N_9916,N_9610);
or U10511 (N_10511,N_8454,N_8916);
nand U10512 (N_10512,N_8150,N_8705);
nand U10513 (N_10513,N_9110,N_8526);
and U10514 (N_10514,N_8074,N_9549);
nor U10515 (N_10515,N_8541,N_9937);
xor U10516 (N_10516,N_8294,N_9988);
and U10517 (N_10517,N_9350,N_9634);
nand U10518 (N_10518,N_9068,N_9081);
nand U10519 (N_10519,N_9699,N_9936);
xor U10520 (N_10520,N_9030,N_9153);
nor U10521 (N_10521,N_8565,N_9257);
nor U10522 (N_10522,N_9573,N_8774);
nor U10523 (N_10523,N_9609,N_8875);
or U10524 (N_10524,N_9455,N_8993);
nor U10525 (N_10525,N_8481,N_9194);
or U10526 (N_10526,N_9405,N_8814);
nand U10527 (N_10527,N_9849,N_8987);
nand U10528 (N_10528,N_9055,N_8937);
nand U10529 (N_10529,N_8195,N_8462);
and U10530 (N_10530,N_9729,N_8291);
or U10531 (N_10531,N_8500,N_9792);
or U10532 (N_10532,N_8453,N_9464);
nor U10533 (N_10533,N_9401,N_9651);
nand U10534 (N_10534,N_8341,N_8215);
or U10535 (N_10535,N_9987,N_8439);
or U10536 (N_10536,N_8813,N_8861);
nor U10537 (N_10537,N_9562,N_8026);
xor U10538 (N_10538,N_9971,N_8745);
nor U10539 (N_10539,N_9583,N_8338);
or U10540 (N_10540,N_8132,N_9039);
or U10541 (N_10541,N_8367,N_8722);
or U10542 (N_10542,N_8845,N_9497);
nor U10543 (N_10543,N_9442,N_9995);
or U10544 (N_10544,N_8063,N_9065);
nor U10545 (N_10545,N_8611,N_8152);
nand U10546 (N_10546,N_9230,N_8505);
nor U10547 (N_10547,N_8990,N_8051);
nand U10548 (N_10548,N_8343,N_9172);
xnor U10549 (N_10549,N_9137,N_8873);
and U10550 (N_10550,N_9036,N_8382);
nand U10551 (N_10551,N_9716,N_8258);
and U10552 (N_10552,N_9572,N_8741);
nor U10553 (N_10553,N_8624,N_9519);
or U10554 (N_10554,N_8286,N_9067);
or U10555 (N_10555,N_9182,N_9814);
nor U10556 (N_10556,N_8675,N_8446);
and U10557 (N_10557,N_9866,N_8571);
nand U10558 (N_10558,N_8954,N_8574);
nand U10559 (N_10559,N_9438,N_9373);
and U10560 (N_10560,N_8414,N_9584);
xnor U10561 (N_10561,N_9638,N_9899);
nor U10562 (N_10562,N_9930,N_8998);
nor U10563 (N_10563,N_9998,N_8634);
nor U10564 (N_10564,N_9703,N_8983);
and U10565 (N_10565,N_8337,N_9026);
nand U10566 (N_10566,N_8495,N_9071);
nor U10567 (N_10567,N_9383,N_9582);
or U10568 (N_10568,N_9157,N_8585);
or U10569 (N_10569,N_9900,N_9338);
nand U10570 (N_10570,N_8841,N_8148);
and U10571 (N_10571,N_9462,N_9950);
nand U10572 (N_10572,N_9981,N_9476);
and U10573 (N_10573,N_9975,N_8227);
and U10574 (N_10574,N_9481,N_9835);
or U10575 (N_10575,N_9148,N_8846);
and U10576 (N_10576,N_8819,N_8223);
nor U10577 (N_10577,N_9484,N_8214);
and U10578 (N_10578,N_8683,N_9755);
nor U10579 (N_10579,N_8457,N_9892);
nand U10580 (N_10580,N_9246,N_8193);
or U10581 (N_10581,N_8903,N_9138);
and U10582 (N_10582,N_8656,N_9193);
nand U10583 (N_10583,N_9542,N_8691);
and U10584 (N_10584,N_9789,N_8714);
nor U10585 (N_10585,N_8102,N_8784);
nor U10586 (N_10586,N_8490,N_9447);
xor U10587 (N_10587,N_9978,N_9810);
nor U10588 (N_10588,N_9376,N_9053);
and U10589 (N_10589,N_9468,N_9315);
and U10590 (N_10590,N_8143,N_8456);
nor U10591 (N_10591,N_8668,N_8124);
or U10592 (N_10592,N_9642,N_9185);
nand U10593 (N_10593,N_8256,N_9546);
or U10594 (N_10594,N_8255,N_9798);
and U10595 (N_10595,N_9045,N_8136);
nand U10596 (N_10596,N_8975,N_9841);
or U10597 (N_10597,N_8348,N_9013);
and U10598 (N_10598,N_9565,N_9037);
or U10599 (N_10599,N_9925,N_9965);
nor U10600 (N_10600,N_8737,N_9285);
nand U10601 (N_10601,N_9345,N_8332);
nor U10602 (N_10602,N_8323,N_9317);
or U10603 (N_10603,N_8234,N_8387);
nand U10604 (N_10604,N_8336,N_8427);
and U10605 (N_10605,N_8001,N_9970);
nor U10606 (N_10606,N_8612,N_9461);
or U10607 (N_10607,N_8251,N_8166);
or U10608 (N_10608,N_9711,N_9305);
nand U10609 (N_10609,N_8630,N_8742);
nand U10610 (N_10610,N_9332,N_8850);
and U10611 (N_10611,N_9726,N_9790);
and U10612 (N_10612,N_8768,N_9996);
xnor U10613 (N_10613,N_8445,N_8697);
and U10614 (N_10614,N_8509,N_8304);
nand U10615 (N_10615,N_8434,N_8023);
and U10616 (N_10616,N_8037,N_9890);
nand U10617 (N_10617,N_9452,N_8550);
nand U10618 (N_10618,N_8425,N_9886);
nand U10619 (N_10619,N_9787,N_9310);
nand U10620 (N_10620,N_8635,N_8694);
nand U10621 (N_10621,N_8619,N_9355);
xor U10622 (N_10622,N_8824,N_8725);
and U10623 (N_10623,N_8392,N_8361);
nand U10624 (N_10624,N_9195,N_8889);
xor U10625 (N_10625,N_8695,N_8394);
xnor U10626 (N_10626,N_9881,N_8079);
nand U10627 (N_10627,N_9555,N_8450);
nor U10628 (N_10628,N_9683,N_8942);
or U10629 (N_10629,N_9425,N_8596);
nand U10630 (N_10630,N_9637,N_8493);
and U10631 (N_10631,N_9669,N_9858);
xor U10632 (N_10632,N_8267,N_9644);
nor U10633 (N_10633,N_9379,N_9785);
and U10634 (N_10634,N_9646,N_8357);
nor U10635 (N_10635,N_9033,N_9723);
nand U10636 (N_10636,N_9837,N_8046);
or U10637 (N_10637,N_8706,N_8731);
and U10638 (N_10638,N_8050,N_8379);
and U10639 (N_10639,N_9775,N_9284);
and U10640 (N_10640,N_8189,N_8174);
xnor U10641 (N_10641,N_9640,N_9377);
nor U10642 (N_10642,N_8065,N_8245);
and U10643 (N_10643,N_8577,N_9494);
or U10644 (N_10644,N_9004,N_9820);
xnor U10645 (N_10645,N_8965,N_9020);
and U10646 (N_10646,N_8146,N_8308);
or U10647 (N_10647,N_8111,N_9209);
and U10648 (N_10648,N_9520,N_9370);
nor U10649 (N_10649,N_8663,N_8250);
nand U10650 (N_10650,N_9843,N_9207);
nand U10651 (N_10651,N_9524,N_9056);
xnor U10652 (N_10652,N_8554,N_9805);
nand U10653 (N_10653,N_9928,N_8795);
nor U10654 (N_10654,N_9880,N_9832);
nand U10655 (N_10655,N_9361,N_9419);
nand U10656 (N_10656,N_8699,N_9722);
nand U10657 (N_10657,N_9083,N_9337);
nor U10658 (N_10658,N_8899,N_9357);
nor U10659 (N_10659,N_8437,N_8806);
and U10660 (N_10660,N_8973,N_8410);
nor U10661 (N_10661,N_8262,N_9788);
or U10662 (N_10662,N_8374,N_9349);
and U10663 (N_10663,N_9210,N_8173);
nand U10664 (N_10664,N_9552,N_8736);
xnor U10665 (N_10665,N_8660,N_8397);
and U10666 (N_10666,N_9096,N_9894);
nor U10667 (N_10667,N_9326,N_9704);
or U10668 (N_10668,N_9745,N_9294);
or U10669 (N_10669,N_9984,N_8658);
nor U10670 (N_10670,N_8579,N_8902);
or U10671 (N_10671,N_8763,N_8766);
nor U10672 (N_10672,N_9279,N_9531);
or U10673 (N_10673,N_9411,N_9134);
nor U10674 (N_10674,N_8767,N_9324);
xnor U10675 (N_10675,N_8499,N_8203);
nor U10676 (N_10676,N_9884,N_9414);
or U10677 (N_10677,N_9239,N_9001);
nor U10678 (N_10678,N_8244,N_9955);
and U10679 (N_10679,N_8206,N_9122);
nor U10680 (N_10680,N_9827,N_9687);
and U10681 (N_10681,N_9696,N_9962);
and U10682 (N_10682,N_9498,N_9693);
nor U10683 (N_10683,N_9517,N_9298);
xor U10684 (N_10684,N_8385,N_8844);
and U10685 (N_10685,N_8568,N_9607);
nand U10686 (N_10686,N_9269,N_8562);
and U10687 (N_10687,N_8018,N_9125);
xnor U10688 (N_10688,N_8218,N_9915);
xnor U10689 (N_10689,N_8949,N_9160);
nand U10690 (N_10690,N_9511,N_8750);
nor U10691 (N_10691,N_9340,N_8467);
xor U10692 (N_10692,N_8521,N_9119);
and U10693 (N_10693,N_9247,N_9003);
xnor U10694 (N_10694,N_9474,N_9862);
and U10695 (N_10695,N_9311,N_8904);
nor U10696 (N_10696,N_8285,N_8056);
nand U10697 (N_10697,N_8582,N_9958);
or U10698 (N_10698,N_9304,N_8558);
nor U10699 (N_10699,N_8388,N_8228);
nor U10700 (N_10700,N_8690,N_9588);
nand U10701 (N_10701,N_9923,N_8085);
and U10702 (N_10702,N_8335,N_8655);
nor U10703 (N_10703,N_9735,N_9589);
nor U10704 (N_10704,N_8331,N_9046);
xor U10705 (N_10705,N_8423,N_9346);
xor U10706 (N_10706,N_8269,N_8031);
or U10707 (N_10707,N_9322,N_8847);
nor U10708 (N_10708,N_9469,N_8287);
or U10709 (N_10709,N_8377,N_8485);
nand U10710 (N_10710,N_9574,N_8632);
and U10711 (N_10711,N_9274,N_8447);
and U10712 (N_10712,N_8372,N_9506);
nor U10713 (N_10713,N_8381,N_9707);
nor U10714 (N_10714,N_9793,N_9206);
or U10715 (N_10715,N_8890,N_9275);
nor U10716 (N_10716,N_9953,N_8968);
and U10717 (N_10717,N_9503,N_8708);
nand U10718 (N_10718,N_9308,N_8368);
and U10719 (N_10719,N_8021,N_9259);
and U10720 (N_10720,N_9396,N_8110);
or U10721 (N_10721,N_8247,N_8959);
or U10722 (N_10722,N_8151,N_9920);
nand U10723 (N_10723,N_8076,N_9500);
nor U10724 (N_10724,N_8230,N_9902);
nand U10725 (N_10725,N_8468,N_8408);
nor U10726 (N_10726,N_9684,N_8210);
nand U10727 (N_10727,N_9818,N_8419);
or U10728 (N_10728,N_8879,N_9385);
nor U10729 (N_10729,N_9115,N_8934);
nand U10730 (N_10730,N_8007,N_8112);
nor U10731 (N_10731,N_8958,N_9177);
and U10732 (N_10732,N_8487,N_8515);
nand U10733 (N_10733,N_9492,N_8253);
and U10734 (N_10734,N_8199,N_9616);
nand U10735 (N_10735,N_8383,N_9098);
and U10736 (N_10736,N_8717,N_8948);
nor U10737 (N_10737,N_8838,N_9641);
nand U10738 (N_10738,N_9901,N_9952);
and U10739 (N_10739,N_9129,N_9802);
nor U10740 (N_10740,N_9101,N_8871);
nor U10741 (N_10741,N_8231,N_8598);
xor U10742 (N_10742,N_9118,N_8677);
or U10743 (N_10743,N_8992,N_8271);
and U10744 (N_10744,N_9913,N_9463);
or U10745 (N_10745,N_8068,N_9994);
nor U10746 (N_10746,N_8225,N_8224);
nand U10747 (N_10747,N_9289,N_8261);
or U10748 (N_10748,N_8290,N_8239);
xor U10749 (N_10749,N_8724,N_9538);
nor U10750 (N_10750,N_8088,N_8827);
and U10751 (N_10751,N_8926,N_8288);
and U10752 (N_10752,N_8176,N_9598);
nor U10753 (N_10753,N_9218,N_9812);
nor U10754 (N_10754,N_9872,N_9592);
nand U10755 (N_10755,N_9380,N_8087);
and U10756 (N_10756,N_9034,N_9397);
nor U10757 (N_10757,N_8130,N_9749);
or U10758 (N_10758,N_8616,N_8399);
or U10759 (N_10759,N_8404,N_8552);
nand U10760 (N_10760,N_8375,N_9943);
xor U10761 (N_10761,N_8154,N_8403);
nor U10762 (N_10762,N_9021,N_8315);
and U10763 (N_10763,N_9453,N_8248);
nor U10764 (N_10764,N_9439,N_8641);
nor U10765 (N_10765,N_9334,N_9168);
or U10766 (N_10766,N_8696,N_9214);
or U10767 (N_10767,N_8333,N_9917);
and U10768 (N_10768,N_8592,N_9753);
and U10769 (N_10769,N_9175,N_8686);
and U10770 (N_10770,N_8422,N_8025);
nand U10771 (N_10771,N_8358,N_8719);
nand U10772 (N_10772,N_8103,N_8137);
and U10773 (N_10773,N_9782,N_8260);
and U10774 (N_10774,N_8646,N_8609);
nor U10775 (N_10775,N_9816,N_8407);
and U10776 (N_10776,N_9251,N_9085);
nand U10777 (N_10777,N_9486,N_9128);
and U10778 (N_10778,N_9147,N_8843);
nor U10779 (N_10779,N_9746,N_8608);
or U10780 (N_10780,N_9653,N_9698);
nand U10781 (N_10781,N_8537,N_9625);
nor U10782 (N_10782,N_9914,N_8796);
xor U10783 (N_10783,N_9877,N_8202);
or U10784 (N_10784,N_8689,N_9694);
nand U10785 (N_10785,N_8553,N_9576);
and U10786 (N_10786,N_8344,N_8575);
or U10787 (N_10787,N_8517,N_9127);
and U10788 (N_10788,N_9718,N_9290);
nor U10789 (N_10789,N_9495,N_9779);
or U10790 (N_10790,N_8010,N_9339);
nand U10791 (N_10791,N_9043,N_9417);
and U10792 (N_10792,N_8470,N_8371);
nand U10793 (N_10793,N_8957,N_8355);
and U10794 (N_10794,N_9800,N_8345);
and U10795 (N_10795,N_9934,N_8442);
nor U10796 (N_10796,N_9107,N_8935);
nor U10797 (N_10797,N_9680,N_8268);
nand U10798 (N_10798,N_8428,N_9919);
or U10799 (N_10799,N_9212,N_8986);
xnor U10800 (N_10800,N_9567,N_8863);
nand U10801 (N_10801,N_9488,N_9882);
and U10802 (N_10802,N_8893,N_8605);
or U10803 (N_10803,N_8077,N_8201);
and U10804 (N_10804,N_9090,N_8969);
nor U10805 (N_10805,N_9174,N_8476);
nor U10806 (N_10806,N_8704,N_8720);
nand U10807 (N_10807,N_9282,N_8980);
nand U10808 (N_10808,N_8698,N_8096);
or U10809 (N_10809,N_8735,N_8808);
and U10810 (N_10810,N_8186,N_9908);
and U10811 (N_10811,N_9508,N_9667);
or U10812 (N_10812,N_9501,N_9258);
nand U10813 (N_10813,N_8601,N_9202);
and U10814 (N_10814,N_8196,N_8662);
and U10815 (N_10815,N_9007,N_9496);
or U10816 (N_10816,N_8852,N_8138);
nand U10817 (N_10817,N_8563,N_9528);
and U10818 (N_10818,N_9525,N_8101);
xor U10819 (N_10819,N_8994,N_9032);
nand U10820 (N_10820,N_9000,N_9725);
or U10821 (N_10821,N_9569,N_9190);
nand U10822 (N_10822,N_8064,N_9959);
or U10823 (N_10823,N_8118,N_8501);
nor U10824 (N_10824,N_9354,N_9402);
and U10825 (N_10825,N_8354,N_8170);
and U10826 (N_10826,N_9954,N_8809);
or U10827 (N_10827,N_9624,N_8773);
xor U10828 (N_10828,N_8951,N_8105);
nand U10829 (N_10829,N_8477,N_8080);
and U10830 (N_10830,N_8561,N_8849);
nand U10831 (N_10831,N_9819,N_9767);
and U10832 (N_10832,N_9808,N_8316);
nor U10833 (N_10833,N_9047,N_8299);
and U10834 (N_10834,N_8324,N_8116);
nor U10835 (N_10835,N_9757,N_8109);
nor U10836 (N_10836,N_8701,N_8123);
nor U10837 (N_10837,N_8529,N_9633);
nor U10838 (N_10838,N_9491,N_8070);
or U10839 (N_10839,N_9170,N_8961);
and U10840 (N_10840,N_8241,N_8160);
or U10841 (N_10841,N_9051,N_9593);
or U10842 (N_10842,N_8349,N_8567);
and U10843 (N_10843,N_9586,N_8917);
xor U10844 (N_10844,N_8945,N_9655);
nor U10845 (N_10845,N_8378,N_8289);
and U10846 (N_10846,N_8960,N_9590);
nor U10847 (N_10847,N_9094,N_9521);
nand U10848 (N_10848,N_8876,N_8504);
nand U10849 (N_10849,N_9398,N_8421);
xor U10850 (N_10850,N_8853,N_9113);
nand U10851 (N_10851,N_8776,N_8329);
nand U10852 (N_10852,N_8181,N_9733);
nand U10853 (N_10853,N_9235,N_9580);
xnor U10854 (N_10854,N_8272,N_8320);
nor U10855 (N_10855,N_9765,N_9577);
and U10856 (N_10856,N_9384,N_8984);
or U10857 (N_10857,N_9450,N_8522);
nand U10858 (N_10858,N_8484,N_9967);
and U10859 (N_10859,N_8881,N_9527);
nand U10860 (N_10860,N_9141,N_8006);
nand U10861 (N_10861,N_9473,N_9406);
and U10862 (N_10862,N_9710,N_9685);
nand U10863 (N_10863,N_8455,N_9921);
and U10864 (N_10864,N_9059,N_8119);
or U10865 (N_10865,N_9024,N_8636);
nor U10866 (N_10866,N_8610,N_9945);
and U10867 (N_10867,N_8200,N_9358);
or U10868 (N_10868,N_9791,N_8107);
or U10869 (N_10869,N_8491,N_8238);
or U10870 (N_10870,N_9591,N_9072);
nand U10871 (N_10871,N_9602,N_8483);
and U10872 (N_10872,N_8746,N_8981);
nand U10873 (N_10873,N_8502,N_9429);
nand U10874 (N_10874,N_8409,N_8169);
and U10875 (N_10875,N_9861,N_9093);
and U10876 (N_10876,N_8019,N_9968);
nand U10877 (N_10877,N_9064,N_9470);
or U10878 (N_10878,N_9482,N_9226);
and U10879 (N_10879,N_9547,N_9948);
nor U10880 (N_10880,N_9017,N_9692);
or U10881 (N_10881,N_9778,N_8353);
nor U10882 (N_10882,N_9008,N_8433);
xor U10883 (N_10883,N_9905,N_9478);
nand U10884 (N_10884,N_8162,N_9252);
nor U10885 (N_10885,N_8753,N_9869);
nand U10886 (N_10886,N_9526,N_9011);
and U10887 (N_10887,N_9636,N_9422);
and U10888 (N_10888,N_8265,N_9700);
or U10889 (N_10889,N_8071,N_9410);
nand U10890 (N_10890,N_8326,N_9169);
nor U10891 (N_10891,N_9052,N_8311);
nand U10892 (N_10892,N_9983,N_9485);
nor U10893 (N_10893,N_8015,N_9974);
nand U10894 (N_10894,N_8475,N_9690);
nor U10895 (N_10895,N_9504,N_8888);
and U10896 (N_10896,N_8098,N_9413);
nor U10897 (N_10897,N_8964,N_9424);
and U10898 (N_10898,N_8167,N_9038);
nand U10899 (N_10899,N_9082,N_9399);
xnor U10900 (N_10900,N_8978,N_9205);
or U10901 (N_10901,N_8303,N_8045);
or U10902 (N_10902,N_9639,N_9106);
or U10903 (N_10903,N_8615,N_9777);
or U10904 (N_10904,N_9301,N_8657);
and U10905 (N_10905,N_9287,N_8647);
xor U10906 (N_10906,N_8346,N_9666);
or U10907 (N_10907,N_8760,N_8094);
nand U10908 (N_10908,N_9714,N_8489);
and U10909 (N_10909,N_9435,N_8685);
or U10910 (N_10910,N_9074,N_9532);
nor U10911 (N_10911,N_9566,N_9523);
nand U10912 (N_10912,N_9395,N_8497);
nand U10913 (N_10913,N_9296,N_9895);
or U10914 (N_10914,N_9176,N_9558);
nor U10915 (N_10915,N_8032,N_9989);
or U10916 (N_10916,N_9010,N_8488);
nand U10917 (N_10917,N_8086,N_8829);
or U10918 (N_10918,N_9635,N_8444);
and U10919 (N_10919,N_9797,N_9557);
or U10920 (N_10920,N_8832,N_8955);
nand U10921 (N_10921,N_9615,N_8785);
nor U10922 (N_10922,N_9986,N_9662);
nand U10923 (N_10923,N_8603,N_8141);
and U10924 (N_10924,N_9721,N_8982);
nor U10925 (N_10925,N_8807,N_8543);
or U10926 (N_10926,N_8498,N_9564);
nor U10927 (N_10927,N_8139,N_8131);
and U10928 (N_10928,N_8788,N_8347);
or U10929 (N_10929,N_9671,N_8002);
and U10930 (N_10930,N_8384,N_8205);
or U10931 (N_10931,N_8280,N_8293);
nor U10932 (N_10932,N_9560,N_8764);
nand U10933 (N_10933,N_8432,N_8867);
and U10934 (N_10934,N_9330,N_8835);
nand U10935 (N_10935,N_8797,N_9678);
xor U10936 (N_10936,N_9850,N_8739);
nor U10937 (N_10937,N_9922,N_8531);
nand U10938 (N_10938,N_8364,N_9432);
or U10939 (N_10939,N_8544,N_9266);
and U10940 (N_10940,N_9092,N_8866);
nor U10941 (N_10941,N_9982,N_9400);
xor U10942 (N_10942,N_9935,N_8573);
nor U10943 (N_10943,N_8825,N_8055);
or U10944 (N_10944,N_9456,N_9544);
nand U10945 (N_10945,N_8327,N_8650);
nand U10946 (N_10946,N_8929,N_9321);
xnor U10947 (N_10947,N_9522,N_8910);
xnor U10948 (N_10948,N_9581,N_9686);
nor U10949 (N_10949,N_8276,N_8622);
or U10950 (N_10950,N_8242,N_9288);
and U10951 (N_10951,N_8547,N_8198);
nor U10952 (N_10952,N_9260,N_9938);
xnor U10953 (N_10953,N_8003,N_8712);
nand U10954 (N_10954,N_8670,N_9031);
and U10955 (N_10955,N_8770,N_8282);
nor U10956 (N_10956,N_9161,N_9313);
or U10957 (N_10957,N_9391,N_8939);
and U10958 (N_10958,N_9139,N_9768);
nand U10959 (N_10959,N_8114,N_8514);
nor U10960 (N_10960,N_8855,N_9451);
xor U10961 (N_10961,N_9941,N_8649);
nor U10962 (N_10962,N_9929,N_8072);
nand U10963 (N_10963,N_8463,N_9457);
nand U10964 (N_10964,N_9423,N_9940);
nand U10965 (N_10965,N_8301,N_8022);
xnor U10966 (N_10966,N_9873,N_8872);
or U10967 (N_10967,N_9548,N_9769);
nand U10968 (N_10968,N_9360,N_8791);
xnor U10969 (N_10969,N_8891,N_8117);
and U10970 (N_10970,N_9466,N_8171);
nor U10971 (N_10971,N_9248,N_8363);
and U10972 (N_10972,N_9803,N_9931);
nor U10973 (N_10973,N_9893,N_8744);
and U10974 (N_10974,N_9944,N_8044);
nand U10975 (N_10975,N_9421,N_8075);
nor U10976 (N_10976,N_8560,N_8710);
or U10977 (N_10977,N_9969,N_9356);
or U10978 (N_10978,N_9272,N_9341);
nand U10979 (N_10979,N_9720,N_9019);
and U10980 (N_10980,N_8030,N_8352);
nand U10981 (N_10981,N_8527,N_9062);
and U10982 (N_10982,N_9876,N_8995);
and U10983 (N_10983,N_8815,N_9387);
nand U10984 (N_10984,N_9044,N_8461);
or U10985 (N_10985,N_8604,N_9594);
nor U10986 (N_10986,N_8322,N_8058);
xor U10987 (N_10987,N_8823,N_9109);
and U10988 (N_10988,N_8878,N_9253);
xor U10989 (N_10989,N_9614,N_8512);
or U10990 (N_10990,N_8593,N_9605);
or U10991 (N_10991,N_8494,N_9087);
nand U10992 (N_10992,N_8651,N_9325);
nand U10993 (N_10993,N_9366,N_9277);
or U10994 (N_10994,N_9393,N_9225);
and U10995 (N_10995,N_9070,N_8496);
and U10996 (N_10996,N_9467,N_9689);
or U10997 (N_10997,N_9822,N_9309);
or U10998 (N_10998,N_9270,N_8243);
nand U10999 (N_10999,N_9828,N_9529);
nor U11000 (N_11000,N_8248,N_9159);
nand U11001 (N_11001,N_8462,N_8327);
nor U11002 (N_11002,N_9765,N_9678);
nor U11003 (N_11003,N_9572,N_9631);
and U11004 (N_11004,N_9892,N_9360);
nand U11005 (N_11005,N_8757,N_9709);
nor U11006 (N_11006,N_8158,N_9922);
nand U11007 (N_11007,N_9522,N_8067);
nor U11008 (N_11008,N_8679,N_9869);
xor U11009 (N_11009,N_8324,N_9475);
and U11010 (N_11010,N_9649,N_8132);
nor U11011 (N_11011,N_9897,N_9624);
nand U11012 (N_11012,N_8716,N_9139);
and U11013 (N_11013,N_9251,N_9775);
nor U11014 (N_11014,N_9317,N_9830);
nor U11015 (N_11015,N_9421,N_9910);
nor U11016 (N_11016,N_9671,N_8305);
nor U11017 (N_11017,N_8140,N_9387);
nand U11018 (N_11018,N_8651,N_9708);
and U11019 (N_11019,N_9859,N_8613);
nand U11020 (N_11020,N_8094,N_8548);
nand U11021 (N_11021,N_9325,N_9833);
nand U11022 (N_11022,N_8546,N_8391);
nand U11023 (N_11023,N_8990,N_8528);
nor U11024 (N_11024,N_9234,N_9192);
xnor U11025 (N_11025,N_8980,N_8525);
or U11026 (N_11026,N_9126,N_8451);
nand U11027 (N_11027,N_8877,N_9392);
and U11028 (N_11028,N_9932,N_9388);
or U11029 (N_11029,N_8311,N_9442);
or U11030 (N_11030,N_8206,N_9568);
xnor U11031 (N_11031,N_8290,N_9725);
and U11032 (N_11032,N_8573,N_9798);
nand U11033 (N_11033,N_8478,N_9257);
nand U11034 (N_11034,N_9542,N_9677);
or U11035 (N_11035,N_8460,N_9467);
or U11036 (N_11036,N_8803,N_9908);
and U11037 (N_11037,N_8678,N_9330);
nand U11038 (N_11038,N_8403,N_9554);
nand U11039 (N_11039,N_9707,N_9736);
and U11040 (N_11040,N_9987,N_9556);
and U11041 (N_11041,N_8666,N_8344);
and U11042 (N_11042,N_9531,N_8897);
nor U11043 (N_11043,N_9901,N_9898);
nor U11044 (N_11044,N_8819,N_9006);
and U11045 (N_11045,N_9719,N_9383);
xnor U11046 (N_11046,N_8525,N_9146);
or U11047 (N_11047,N_9869,N_8606);
nand U11048 (N_11048,N_9757,N_9664);
or U11049 (N_11049,N_9513,N_8668);
or U11050 (N_11050,N_9956,N_8349);
or U11051 (N_11051,N_8837,N_9980);
nand U11052 (N_11052,N_8216,N_9668);
or U11053 (N_11053,N_9645,N_9476);
and U11054 (N_11054,N_8974,N_9510);
and U11055 (N_11055,N_8320,N_9612);
nand U11056 (N_11056,N_9694,N_8106);
nor U11057 (N_11057,N_9968,N_9133);
and U11058 (N_11058,N_9728,N_9382);
nand U11059 (N_11059,N_9497,N_8781);
nor U11060 (N_11060,N_8773,N_8648);
xnor U11061 (N_11061,N_8565,N_9205);
xnor U11062 (N_11062,N_8645,N_8334);
and U11063 (N_11063,N_8313,N_9858);
xnor U11064 (N_11064,N_8950,N_9815);
nand U11065 (N_11065,N_8786,N_9798);
or U11066 (N_11066,N_9073,N_8995);
nand U11067 (N_11067,N_9979,N_8133);
and U11068 (N_11068,N_9175,N_9209);
nor U11069 (N_11069,N_9341,N_9150);
nor U11070 (N_11070,N_8784,N_9942);
nand U11071 (N_11071,N_9809,N_8553);
or U11072 (N_11072,N_8362,N_8462);
nor U11073 (N_11073,N_9546,N_8045);
or U11074 (N_11074,N_9723,N_9287);
or U11075 (N_11075,N_9119,N_8441);
xor U11076 (N_11076,N_9614,N_9590);
xnor U11077 (N_11077,N_8678,N_9191);
xor U11078 (N_11078,N_9894,N_9861);
and U11079 (N_11079,N_8436,N_9190);
and U11080 (N_11080,N_8309,N_8013);
nand U11081 (N_11081,N_8639,N_8150);
nand U11082 (N_11082,N_8655,N_9245);
xnor U11083 (N_11083,N_8818,N_8217);
nand U11084 (N_11084,N_9319,N_8728);
nand U11085 (N_11085,N_9156,N_8577);
nand U11086 (N_11086,N_9471,N_8034);
xor U11087 (N_11087,N_8020,N_9180);
xor U11088 (N_11088,N_9266,N_9719);
nand U11089 (N_11089,N_9549,N_9780);
nand U11090 (N_11090,N_8756,N_8091);
xor U11091 (N_11091,N_8847,N_8454);
xor U11092 (N_11092,N_9795,N_9917);
nor U11093 (N_11093,N_9540,N_9786);
nor U11094 (N_11094,N_9038,N_9854);
and U11095 (N_11095,N_9476,N_8695);
xnor U11096 (N_11096,N_9521,N_8544);
or U11097 (N_11097,N_8735,N_9220);
nor U11098 (N_11098,N_8472,N_9177);
nor U11099 (N_11099,N_9643,N_8776);
nand U11100 (N_11100,N_8058,N_8131);
nor U11101 (N_11101,N_8988,N_8285);
nand U11102 (N_11102,N_9123,N_9719);
nor U11103 (N_11103,N_9869,N_8009);
nor U11104 (N_11104,N_9832,N_8835);
nor U11105 (N_11105,N_9555,N_8762);
or U11106 (N_11106,N_8375,N_8781);
nand U11107 (N_11107,N_9283,N_9899);
and U11108 (N_11108,N_8266,N_8390);
and U11109 (N_11109,N_8253,N_9852);
and U11110 (N_11110,N_9543,N_8574);
xnor U11111 (N_11111,N_8505,N_9380);
and U11112 (N_11112,N_8395,N_9325);
or U11113 (N_11113,N_9950,N_8861);
nor U11114 (N_11114,N_9731,N_8400);
nand U11115 (N_11115,N_8470,N_9796);
nand U11116 (N_11116,N_8537,N_8177);
or U11117 (N_11117,N_9198,N_9279);
nand U11118 (N_11118,N_9728,N_9443);
xor U11119 (N_11119,N_8741,N_8419);
and U11120 (N_11120,N_9823,N_9228);
nand U11121 (N_11121,N_9277,N_9453);
nor U11122 (N_11122,N_9881,N_8298);
xor U11123 (N_11123,N_9547,N_8620);
nand U11124 (N_11124,N_9726,N_9282);
or U11125 (N_11125,N_9803,N_8891);
nand U11126 (N_11126,N_9223,N_8865);
or U11127 (N_11127,N_8504,N_9157);
xor U11128 (N_11128,N_9760,N_8901);
xnor U11129 (N_11129,N_8443,N_8881);
and U11130 (N_11130,N_9981,N_9401);
or U11131 (N_11131,N_9629,N_9759);
nor U11132 (N_11132,N_9411,N_9711);
and U11133 (N_11133,N_8809,N_9880);
xnor U11134 (N_11134,N_8251,N_8552);
nor U11135 (N_11135,N_8489,N_9744);
and U11136 (N_11136,N_8253,N_8782);
nand U11137 (N_11137,N_8442,N_8408);
nand U11138 (N_11138,N_8280,N_9217);
and U11139 (N_11139,N_9455,N_8967);
nor U11140 (N_11140,N_8810,N_8106);
or U11141 (N_11141,N_8172,N_8951);
nor U11142 (N_11142,N_8401,N_9391);
nand U11143 (N_11143,N_9081,N_8280);
and U11144 (N_11144,N_8240,N_8994);
and U11145 (N_11145,N_8393,N_9120);
and U11146 (N_11146,N_8801,N_8912);
nor U11147 (N_11147,N_9643,N_9088);
nand U11148 (N_11148,N_9203,N_8022);
and U11149 (N_11149,N_9733,N_9381);
xnor U11150 (N_11150,N_9080,N_9892);
and U11151 (N_11151,N_8336,N_8702);
nor U11152 (N_11152,N_8117,N_8598);
and U11153 (N_11153,N_8084,N_9440);
or U11154 (N_11154,N_9795,N_9889);
nand U11155 (N_11155,N_8342,N_8656);
nand U11156 (N_11156,N_8272,N_9256);
nor U11157 (N_11157,N_9061,N_9725);
or U11158 (N_11158,N_8672,N_9589);
or U11159 (N_11159,N_9060,N_9633);
and U11160 (N_11160,N_8394,N_9645);
and U11161 (N_11161,N_8198,N_9868);
nand U11162 (N_11162,N_8125,N_9212);
xor U11163 (N_11163,N_8329,N_8990);
and U11164 (N_11164,N_8128,N_8154);
nor U11165 (N_11165,N_8559,N_9386);
xor U11166 (N_11166,N_8551,N_9277);
or U11167 (N_11167,N_8342,N_9248);
or U11168 (N_11168,N_9013,N_9273);
or U11169 (N_11169,N_8411,N_9297);
nand U11170 (N_11170,N_8668,N_8168);
nor U11171 (N_11171,N_8028,N_9761);
and U11172 (N_11172,N_8103,N_9568);
nor U11173 (N_11173,N_9894,N_9485);
and U11174 (N_11174,N_9972,N_9692);
nand U11175 (N_11175,N_9957,N_9541);
nor U11176 (N_11176,N_8253,N_9552);
xor U11177 (N_11177,N_9718,N_8433);
or U11178 (N_11178,N_9718,N_9960);
or U11179 (N_11179,N_9849,N_8392);
or U11180 (N_11180,N_8805,N_8957);
nor U11181 (N_11181,N_8728,N_9028);
nor U11182 (N_11182,N_8368,N_8720);
or U11183 (N_11183,N_9813,N_9731);
nand U11184 (N_11184,N_8288,N_8736);
or U11185 (N_11185,N_8414,N_9436);
nand U11186 (N_11186,N_9339,N_9670);
or U11187 (N_11187,N_8864,N_9868);
xnor U11188 (N_11188,N_9491,N_8635);
nand U11189 (N_11189,N_9503,N_8036);
nand U11190 (N_11190,N_8708,N_8750);
and U11191 (N_11191,N_8804,N_9909);
nor U11192 (N_11192,N_9422,N_9198);
or U11193 (N_11193,N_9240,N_8076);
and U11194 (N_11194,N_9076,N_9822);
and U11195 (N_11195,N_9879,N_8881);
nor U11196 (N_11196,N_9282,N_8170);
and U11197 (N_11197,N_8292,N_9857);
nor U11198 (N_11198,N_9974,N_9643);
and U11199 (N_11199,N_9266,N_8598);
or U11200 (N_11200,N_9544,N_8230);
or U11201 (N_11201,N_8824,N_8551);
or U11202 (N_11202,N_9266,N_8370);
or U11203 (N_11203,N_9901,N_9579);
nor U11204 (N_11204,N_8731,N_8409);
or U11205 (N_11205,N_8550,N_8411);
nor U11206 (N_11206,N_9151,N_9314);
nand U11207 (N_11207,N_9758,N_9997);
or U11208 (N_11208,N_8232,N_8669);
or U11209 (N_11209,N_8353,N_8113);
and U11210 (N_11210,N_8612,N_9710);
or U11211 (N_11211,N_8164,N_9712);
and U11212 (N_11212,N_9020,N_9121);
and U11213 (N_11213,N_8290,N_9397);
or U11214 (N_11214,N_8367,N_9554);
nor U11215 (N_11215,N_8324,N_9267);
or U11216 (N_11216,N_9235,N_9642);
and U11217 (N_11217,N_8491,N_8508);
or U11218 (N_11218,N_8932,N_8104);
nand U11219 (N_11219,N_9976,N_8463);
nor U11220 (N_11220,N_8396,N_9219);
nor U11221 (N_11221,N_9706,N_8135);
and U11222 (N_11222,N_8973,N_9967);
xor U11223 (N_11223,N_8575,N_9638);
or U11224 (N_11224,N_8493,N_8661);
nor U11225 (N_11225,N_8335,N_9160);
nand U11226 (N_11226,N_8591,N_9737);
nand U11227 (N_11227,N_8530,N_8841);
nand U11228 (N_11228,N_8536,N_8526);
xnor U11229 (N_11229,N_9160,N_8742);
or U11230 (N_11230,N_9596,N_9984);
nand U11231 (N_11231,N_9641,N_8548);
nor U11232 (N_11232,N_8770,N_8652);
nand U11233 (N_11233,N_8418,N_8440);
or U11234 (N_11234,N_8824,N_9596);
or U11235 (N_11235,N_8855,N_9180);
and U11236 (N_11236,N_8828,N_8096);
nor U11237 (N_11237,N_8774,N_9439);
nor U11238 (N_11238,N_8010,N_9958);
xnor U11239 (N_11239,N_9336,N_8380);
nand U11240 (N_11240,N_8251,N_8119);
and U11241 (N_11241,N_8636,N_9084);
nand U11242 (N_11242,N_9780,N_8237);
xor U11243 (N_11243,N_9991,N_8455);
nand U11244 (N_11244,N_9993,N_9745);
nand U11245 (N_11245,N_8827,N_8857);
and U11246 (N_11246,N_9325,N_9614);
nor U11247 (N_11247,N_9653,N_9901);
or U11248 (N_11248,N_8877,N_8831);
and U11249 (N_11249,N_8850,N_8800);
or U11250 (N_11250,N_8813,N_8070);
nor U11251 (N_11251,N_8625,N_8732);
nand U11252 (N_11252,N_8238,N_8734);
nand U11253 (N_11253,N_9796,N_9981);
xor U11254 (N_11254,N_9949,N_8891);
and U11255 (N_11255,N_9695,N_9421);
nand U11256 (N_11256,N_8781,N_8002);
and U11257 (N_11257,N_9807,N_9283);
or U11258 (N_11258,N_8360,N_8683);
xnor U11259 (N_11259,N_9083,N_9171);
nand U11260 (N_11260,N_9241,N_8970);
or U11261 (N_11261,N_8005,N_9792);
nor U11262 (N_11262,N_9923,N_9021);
nor U11263 (N_11263,N_8682,N_8450);
nand U11264 (N_11264,N_8622,N_8828);
or U11265 (N_11265,N_9398,N_9249);
or U11266 (N_11266,N_8212,N_8583);
nand U11267 (N_11267,N_8610,N_8867);
or U11268 (N_11268,N_8007,N_8311);
or U11269 (N_11269,N_8313,N_8586);
xor U11270 (N_11270,N_9912,N_9547);
nand U11271 (N_11271,N_8474,N_9970);
nand U11272 (N_11272,N_8933,N_9183);
or U11273 (N_11273,N_8609,N_9811);
nor U11274 (N_11274,N_8443,N_9618);
nor U11275 (N_11275,N_8520,N_8397);
nand U11276 (N_11276,N_8181,N_9050);
or U11277 (N_11277,N_9480,N_8955);
xnor U11278 (N_11278,N_8755,N_9905);
nor U11279 (N_11279,N_8892,N_8204);
and U11280 (N_11280,N_8106,N_8210);
nor U11281 (N_11281,N_8879,N_9300);
nand U11282 (N_11282,N_9138,N_9778);
xor U11283 (N_11283,N_8434,N_9817);
or U11284 (N_11284,N_9828,N_8012);
or U11285 (N_11285,N_9421,N_9599);
nor U11286 (N_11286,N_8698,N_8184);
nor U11287 (N_11287,N_9440,N_8057);
nand U11288 (N_11288,N_9356,N_8915);
nor U11289 (N_11289,N_8773,N_9448);
nand U11290 (N_11290,N_9625,N_8814);
nand U11291 (N_11291,N_8982,N_9776);
nand U11292 (N_11292,N_8199,N_8117);
nor U11293 (N_11293,N_9257,N_9170);
xnor U11294 (N_11294,N_9794,N_9529);
nor U11295 (N_11295,N_8856,N_9963);
nor U11296 (N_11296,N_8621,N_8527);
and U11297 (N_11297,N_8811,N_8726);
xor U11298 (N_11298,N_8939,N_8946);
nor U11299 (N_11299,N_9309,N_9810);
nand U11300 (N_11300,N_8871,N_8433);
or U11301 (N_11301,N_8589,N_8030);
nand U11302 (N_11302,N_8565,N_8205);
nor U11303 (N_11303,N_9105,N_9160);
xor U11304 (N_11304,N_8957,N_8627);
and U11305 (N_11305,N_9633,N_9959);
nand U11306 (N_11306,N_9264,N_9553);
xnor U11307 (N_11307,N_8919,N_9027);
and U11308 (N_11308,N_9513,N_8201);
nand U11309 (N_11309,N_9026,N_8096);
or U11310 (N_11310,N_8051,N_9937);
nand U11311 (N_11311,N_9667,N_8524);
or U11312 (N_11312,N_9529,N_9701);
and U11313 (N_11313,N_8514,N_8571);
nand U11314 (N_11314,N_9708,N_9501);
nor U11315 (N_11315,N_8095,N_8120);
nand U11316 (N_11316,N_9270,N_8238);
and U11317 (N_11317,N_8805,N_9929);
xor U11318 (N_11318,N_8001,N_9451);
and U11319 (N_11319,N_8096,N_9641);
nand U11320 (N_11320,N_9763,N_8271);
and U11321 (N_11321,N_9616,N_9405);
nor U11322 (N_11322,N_9930,N_8039);
nand U11323 (N_11323,N_9459,N_8259);
xnor U11324 (N_11324,N_9596,N_9088);
and U11325 (N_11325,N_8187,N_9741);
and U11326 (N_11326,N_8763,N_9440);
or U11327 (N_11327,N_8659,N_8073);
and U11328 (N_11328,N_8327,N_8257);
nand U11329 (N_11329,N_8883,N_9608);
nand U11330 (N_11330,N_9816,N_8671);
and U11331 (N_11331,N_9832,N_8887);
and U11332 (N_11332,N_9072,N_9756);
nor U11333 (N_11333,N_9700,N_8643);
and U11334 (N_11334,N_9590,N_9501);
and U11335 (N_11335,N_8189,N_9746);
nor U11336 (N_11336,N_9245,N_9180);
or U11337 (N_11337,N_9832,N_9989);
nand U11338 (N_11338,N_9927,N_8989);
or U11339 (N_11339,N_9808,N_9860);
nand U11340 (N_11340,N_8329,N_8600);
nor U11341 (N_11341,N_9057,N_8520);
or U11342 (N_11342,N_8156,N_9290);
nor U11343 (N_11343,N_9554,N_9673);
nor U11344 (N_11344,N_9902,N_8982);
nand U11345 (N_11345,N_8635,N_9921);
and U11346 (N_11346,N_9993,N_9487);
nand U11347 (N_11347,N_9882,N_9261);
and U11348 (N_11348,N_8888,N_8153);
nor U11349 (N_11349,N_9704,N_8903);
or U11350 (N_11350,N_8600,N_8882);
or U11351 (N_11351,N_9152,N_8597);
nor U11352 (N_11352,N_9439,N_8507);
and U11353 (N_11353,N_8370,N_8690);
or U11354 (N_11354,N_8188,N_9387);
nor U11355 (N_11355,N_8306,N_8707);
and U11356 (N_11356,N_9182,N_8613);
nand U11357 (N_11357,N_9645,N_9433);
nand U11358 (N_11358,N_8036,N_8644);
nor U11359 (N_11359,N_8164,N_9833);
nand U11360 (N_11360,N_8393,N_9710);
and U11361 (N_11361,N_9276,N_8587);
nor U11362 (N_11362,N_8647,N_9476);
nor U11363 (N_11363,N_9018,N_8268);
nor U11364 (N_11364,N_8693,N_8190);
nor U11365 (N_11365,N_8010,N_8649);
or U11366 (N_11366,N_8980,N_8669);
and U11367 (N_11367,N_9156,N_8469);
or U11368 (N_11368,N_8183,N_8539);
nand U11369 (N_11369,N_9390,N_8491);
nor U11370 (N_11370,N_9695,N_8713);
or U11371 (N_11371,N_9354,N_9316);
and U11372 (N_11372,N_9146,N_9522);
nand U11373 (N_11373,N_9600,N_9329);
nand U11374 (N_11374,N_9100,N_9546);
and U11375 (N_11375,N_9650,N_9870);
nand U11376 (N_11376,N_8908,N_8420);
xnor U11377 (N_11377,N_9085,N_9141);
nand U11378 (N_11378,N_9611,N_9581);
nand U11379 (N_11379,N_9204,N_9841);
nor U11380 (N_11380,N_9602,N_9263);
nand U11381 (N_11381,N_9541,N_9971);
nand U11382 (N_11382,N_8423,N_8970);
nor U11383 (N_11383,N_8669,N_8389);
or U11384 (N_11384,N_9139,N_9509);
xor U11385 (N_11385,N_8844,N_9708);
nand U11386 (N_11386,N_9258,N_8332);
or U11387 (N_11387,N_9170,N_8389);
or U11388 (N_11388,N_9133,N_8151);
or U11389 (N_11389,N_9043,N_8030);
nor U11390 (N_11390,N_8636,N_9725);
and U11391 (N_11391,N_8480,N_9052);
nor U11392 (N_11392,N_9031,N_8241);
and U11393 (N_11393,N_9936,N_9911);
nor U11394 (N_11394,N_8255,N_9793);
xor U11395 (N_11395,N_8280,N_9314);
nand U11396 (N_11396,N_8308,N_9727);
nor U11397 (N_11397,N_8789,N_8632);
nand U11398 (N_11398,N_8229,N_9591);
or U11399 (N_11399,N_8797,N_8454);
nor U11400 (N_11400,N_8635,N_8333);
nor U11401 (N_11401,N_8382,N_8634);
nand U11402 (N_11402,N_9570,N_9263);
and U11403 (N_11403,N_8683,N_8103);
and U11404 (N_11404,N_9067,N_8075);
nand U11405 (N_11405,N_8175,N_9853);
nor U11406 (N_11406,N_9448,N_9562);
nor U11407 (N_11407,N_9826,N_9890);
nand U11408 (N_11408,N_8729,N_8870);
or U11409 (N_11409,N_9957,N_9493);
or U11410 (N_11410,N_9660,N_9879);
nand U11411 (N_11411,N_9294,N_8771);
nor U11412 (N_11412,N_8967,N_9362);
xor U11413 (N_11413,N_9596,N_8779);
nor U11414 (N_11414,N_9069,N_9767);
nand U11415 (N_11415,N_9256,N_8435);
nor U11416 (N_11416,N_8109,N_9259);
and U11417 (N_11417,N_8415,N_8635);
or U11418 (N_11418,N_8833,N_9747);
xor U11419 (N_11419,N_8980,N_9379);
xor U11420 (N_11420,N_9625,N_9217);
nand U11421 (N_11421,N_8464,N_8694);
and U11422 (N_11422,N_9247,N_8197);
xor U11423 (N_11423,N_8544,N_9493);
and U11424 (N_11424,N_8141,N_8959);
or U11425 (N_11425,N_9313,N_8955);
and U11426 (N_11426,N_8071,N_8431);
nand U11427 (N_11427,N_8045,N_9399);
or U11428 (N_11428,N_9387,N_9661);
nor U11429 (N_11429,N_8118,N_8253);
nor U11430 (N_11430,N_8045,N_8627);
or U11431 (N_11431,N_8236,N_8385);
nand U11432 (N_11432,N_9131,N_9985);
nor U11433 (N_11433,N_9164,N_8028);
or U11434 (N_11434,N_9676,N_8533);
nand U11435 (N_11435,N_9839,N_9974);
nand U11436 (N_11436,N_8515,N_8203);
nor U11437 (N_11437,N_9458,N_8708);
nor U11438 (N_11438,N_8747,N_8424);
xor U11439 (N_11439,N_8414,N_9351);
xor U11440 (N_11440,N_9362,N_8989);
nand U11441 (N_11441,N_9798,N_8288);
and U11442 (N_11442,N_8126,N_9629);
and U11443 (N_11443,N_9062,N_8974);
nand U11444 (N_11444,N_9075,N_8444);
and U11445 (N_11445,N_8704,N_8535);
nand U11446 (N_11446,N_9006,N_8228);
or U11447 (N_11447,N_9808,N_9765);
or U11448 (N_11448,N_8693,N_8179);
nand U11449 (N_11449,N_8028,N_9313);
and U11450 (N_11450,N_9024,N_9779);
or U11451 (N_11451,N_8259,N_9183);
nand U11452 (N_11452,N_8545,N_9865);
nor U11453 (N_11453,N_9032,N_8097);
nand U11454 (N_11454,N_8606,N_9781);
or U11455 (N_11455,N_8771,N_8538);
xor U11456 (N_11456,N_9564,N_8104);
nor U11457 (N_11457,N_8841,N_9639);
nor U11458 (N_11458,N_8177,N_8841);
or U11459 (N_11459,N_9428,N_9319);
nor U11460 (N_11460,N_9702,N_9033);
nor U11461 (N_11461,N_8465,N_8666);
and U11462 (N_11462,N_9739,N_8693);
or U11463 (N_11463,N_8209,N_8036);
nor U11464 (N_11464,N_9660,N_9240);
nand U11465 (N_11465,N_8068,N_9131);
nand U11466 (N_11466,N_9935,N_8390);
nor U11467 (N_11467,N_9933,N_8889);
and U11468 (N_11468,N_9334,N_9810);
or U11469 (N_11469,N_9561,N_9054);
and U11470 (N_11470,N_8847,N_9301);
nand U11471 (N_11471,N_8792,N_8702);
nand U11472 (N_11472,N_8765,N_8498);
xnor U11473 (N_11473,N_9512,N_8327);
and U11474 (N_11474,N_8235,N_8640);
nand U11475 (N_11475,N_9170,N_8340);
nor U11476 (N_11476,N_9738,N_8596);
nand U11477 (N_11477,N_9209,N_8784);
nand U11478 (N_11478,N_9447,N_9907);
nor U11479 (N_11479,N_8784,N_9327);
nor U11480 (N_11480,N_8407,N_9880);
nand U11481 (N_11481,N_8475,N_9293);
nand U11482 (N_11482,N_9128,N_8850);
nand U11483 (N_11483,N_9355,N_9334);
nand U11484 (N_11484,N_9173,N_9363);
and U11485 (N_11485,N_8637,N_9588);
xor U11486 (N_11486,N_9703,N_8381);
nor U11487 (N_11487,N_9687,N_8221);
and U11488 (N_11488,N_9779,N_9035);
nor U11489 (N_11489,N_8664,N_8324);
nor U11490 (N_11490,N_8065,N_8636);
xor U11491 (N_11491,N_9848,N_9123);
and U11492 (N_11492,N_9367,N_8281);
nand U11493 (N_11493,N_9005,N_9862);
nor U11494 (N_11494,N_9096,N_9602);
nand U11495 (N_11495,N_8379,N_8414);
or U11496 (N_11496,N_9826,N_8078);
nor U11497 (N_11497,N_8841,N_9961);
nor U11498 (N_11498,N_9055,N_9899);
nand U11499 (N_11499,N_9204,N_8880);
and U11500 (N_11500,N_9220,N_8207);
nand U11501 (N_11501,N_8677,N_8535);
xnor U11502 (N_11502,N_8075,N_9745);
or U11503 (N_11503,N_8488,N_9808);
xor U11504 (N_11504,N_9511,N_9826);
or U11505 (N_11505,N_8818,N_8935);
or U11506 (N_11506,N_9195,N_9557);
and U11507 (N_11507,N_9480,N_8375);
nor U11508 (N_11508,N_9166,N_8433);
and U11509 (N_11509,N_8963,N_8381);
nor U11510 (N_11510,N_9914,N_9867);
nor U11511 (N_11511,N_9285,N_8015);
or U11512 (N_11512,N_8783,N_8218);
nand U11513 (N_11513,N_9147,N_9802);
nor U11514 (N_11514,N_8117,N_8691);
and U11515 (N_11515,N_8408,N_8986);
nand U11516 (N_11516,N_8914,N_8376);
xor U11517 (N_11517,N_9813,N_8105);
nand U11518 (N_11518,N_8075,N_9671);
nand U11519 (N_11519,N_8590,N_9951);
xnor U11520 (N_11520,N_9478,N_9615);
nand U11521 (N_11521,N_8429,N_8802);
or U11522 (N_11522,N_8963,N_8288);
and U11523 (N_11523,N_8784,N_8188);
nand U11524 (N_11524,N_9182,N_9301);
nor U11525 (N_11525,N_9832,N_8579);
nand U11526 (N_11526,N_8607,N_8685);
nand U11527 (N_11527,N_8214,N_8964);
or U11528 (N_11528,N_8558,N_9401);
nor U11529 (N_11529,N_9136,N_8015);
nor U11530 (N_11530,N_9884,N_8773);
or U11531 (N_11531,N_8386,N_8563);
or U11532 (N_11532,N_9879,N_9626);
or U11533 (N_11533,N_9569,N_8545);
nand U11534 (N_11534,N_9631,N_8002);
nand U11535 (N_11535,N_8994,N_8000);
and U11536 (N_11536,N_8969,N_8240);
and U11537 (N_11537,N_8224,N_8152);
nor U11538 (N_11538,N_9492,N_8161);
or U11539 (N_11539,N_9429,N_9229);
and U11540 (N_11540,N_8991,N_8834);
or U11541 (N_11541,N_8417,N_9026);
xor U11542 (N_11542,N_9663,N_9721);
nor U11543 (N_11543,N_9507,N_8092);
nand U11544 (N_11544,N_8008,N_8997);
nor U11545 (N_11545,N_9141,N_9901);
or U11546 (N_11546,N_8342,N_9623);
nor U11547 (N_11547,N_9119,N_9710);
xor U11548 (N_11548,N_8122,N_9687);
nand U11549 (N_11549,N_9410,N_9282);
nand U11550 (N_11550,N_9552,N_9595);
and U11551 (N_11551,N_8697,N_8213);
or U11552 (N_11552,N_8238,N_9504);
nand U11553 (N_11553,N_8350,N_8166);
and U11554 (N_11554,N_8752,N_8763);
nor U11555 (N_11555,N_9629,N_8285);
and U11556 (N_11556,N_9257,N_8859);
or U11557 (N_11557,N_8168,N_8459);
nand U11558 (N_11558,N_8443,N_9633);
or U11559 (N_11559,N_8671,N_9212);
and U11560 (N_11560,N_9656,N_9888);
nand U11561 (N_11561,N_9552,N_9669);
nor U11562 (N_11562,N_9382,N_8350);
nor U11563 (N_11563,N_9927,N_9238);
or U11564 (N_11564,N_8413,N_9092);
and U11565 (N_11565,N_9513,N_9529);
and U11566 (N_11566,N_9438,N_8475);
nor U11567 (N_11567,N_8760,N_8752);
nor U11568 (N_11568,N_8431,N_9424);
xnor U11569 (N_11569,N_8437,N_8188);
or U11570 (N_11570,N_8374,N_9866);
nand U11571 (N_11571,N_8278,N_9649);
or U11572 (N_11572,N_9279,N_9317);
nand U11573 (N_11573,N_9450,N_8680);
nand U11574 (N_11574,N_9485,N_9734);
or U11575 (N_11575,N_8547,N_8045);
nor U11576 (N_11576,N_8770,N_9521);
nand U11577 (N_11577,N_8280,N_8764);
nand U11578 (N_11578,N_9020,N_8571);
and U11579 (N_11579,N_9481,N_9425);
nor U11580 (N_11580,N_8716,N_8247);
and U11581 (N_11581,N_9465,N_9840);
nand U11582 (N_11582,N_9533,N_8359);
nor U11583 (N_11583,N_8978,N_8749);
and U11584 (N_11584,N_9499,N_8959);
and U11585 (N_11585,N_9030,N_8598);
nor U11586 (N_11586,N_8386,N_9871);
and U11587 (N_11587,N_9221,N_8617);
nand U11588 (N_11588,N_8019,N_8077);
and U11589 (N_11589,N_8487,N_8910);
and U11590 (N_11590,N_9991,N_8991);
nor U11591 (N_11591,N_9954,N_9051);
or U11592 (N_11592,N_9579,N_9813);
or U11593 (N_11593,N_9731,N_8567);
or U11594 (N_11594,N_8161,N_9621);
nand U11595 (N_11595,N_8525,N_9724);
and U11596 (N_11596,N_9083,N_9401);
and U11597 (N_11597,N_9857,N_9318);
xnor U11598 (N_11598,N_9683,N_8199);
nor U11599 (N_11599,N_8100,N_8379);
and U11600 (N_11600,N_8660,N_9442);
nor U11601 (N_11601,N_8116,N_9361);
and U11602 (N_11602,N_9796,N_9822);
xnor U11603 (N_11603,N_8294,N_9106);
nor U11604 (N_11604,N_8943,N_8515);
nand U11605 (N_11605,N_9387,N_8209);
xnor U11606 (N_11606,N_8979,N_9938);
or U11607 (N_11607,N_9207,N_9522);
or U11608 (N_11608,N_9685,N_9564);
nor U11609 (N_11609,N_8808,N_8636);
nand U11610 (N_11610,N_8287,N_9298);
or U11611 (N_11611,N_8000,N_9779);
or U11612 (N_11612,N_9456,N_8676);
and U11613 (N_11613,N_9916,N_9382);
or U11614 (N_11614,N_9013,N_8535);
nand U11615 (N_11615,N_9805,N_9022);
nor U11616 (N_11616,N_8749,N_9815);
and U11617 (N_11617,N_9237,N_8815);
or U11618 (N_11618,N_8763,N_8559);
or U11619 (N_11619,N_8357,N_8282);
nor U11620 (N_11620,N_8836,N_8270);
and U11621 (N_11621,N_8300,N_9092);
nor U11622 (N_11622,N_9500,N_8560);
nand U11623 (N_11623,N_8744,N_9815);
nand U11624 (N_11624,N_9121,N_8094);
nor U11625 (N_11625,N_9802,N_8909);
nand U11626 (N_11626,N_9199,N_8168);
or U11627 (N_11627,N_8560,N_8494);
nand U11628 (N_11628,N_8504,N_8489);
nand U11629 (N_11629,N_9599,N_8747);
nand U11630 (N_11630,N_9664,N_8112);
nor U11631 (N_11631,N_9379,N_9551);
nor U11632 (N_11632,N_9345,N_8164);
nor U11633 (N_11633,N_9526,N_8558);
or U11634 (N_11634,N_9575,N_9131);
or U11635 (N_11635,N_8491,N_9560);
or U11636 (N_11636,N_8020,N_9475);
or U11637 (N_11637,N_9994,N_8967);
nand U11638 (N_11638,N_8522,N_9655);
xor U11639 (N_11639,N_9497,N_8071);
and U11640 (N_11640,N_8864,N_8487);
and U11641 (N_11641,N_8494,N_9111);
or U11642 (N_11642,N_9277,N_8771);
xnor U11643 (N_11643,N_9466,N_9153);
xor U11644 (N_11644,N_8121,N_9404);
or U11645 (N_11645,N_8322,N_8349);
and U11646 (N_11646,N_9675,N_8615);
nor U11647 (N_11647,N_8701,N_8358);
xor U11648 (N_11648,N_9353,N_8159);
and U11649 (N_11649,N_9088,N_9809);
nand U11650 (N_11650,N_8475,N_9572);
and U11651 (N_11651,N_9052,N_8459);
nor U11652 (N_11652,N_8790,N_9660);
or U11653 (N_11653,N_9392,N_9482);
nor U11654 (N_11654,N_8997,N_8285);
nand U11655 (N_11655,N_9123,N_9325);
nand U11656 (N_11656,N_9006,N_9359);
nand U11657 (N_11657,N_9165,N_9818);
nand U11658 (N_11658,N_9542,N_8387);
or U11659 (N_11659,N_8148,N_9403);
or U11660 (N_11660,N_9991,N_8008);
nor U11661 (N_11661,N_8299,N_8071);
or U11662 (N_11662,N_9686,N_9713);
nor U11663 (N_11663,N_9963,N_8063);
or U11664 (N_11664,N_9418,N_9871);
or U11665 (N_11665,N_9974,N_9222);
or U11666 (N_11666,N_8254,N_8054);
xnor U11667 (N_11667,N_9839,N_9242);
nand U11668 (N_11668,N_8747,N_8421);
nand U11669 (N_11669,N_8665,N_9072);
nor U11670 (N_11670,N_9808,N_8605);
or U11671 (N_11671,N_8648,N_9125);
xnor U11672 (N_11672,N_8926,N_9646);
nand U11673 (N_11673,N_9925,N_9151);
and U11674 (N_11674,N_9612,N_8675);
or U11675 (N_11675,N_8806,N_9641);
xor U11676 (N_11676,N_8731,N_9678);
and U11677 (N_11677,N_9301,N_8912);
nand U11678 (N_11678,N_8111,N_8108);
nand U11679 (N_11679,N_9384,N_9327);
nor U11680 (N_11680,N_8020,N_9892);
or U11681 (N_11681,N_9753,N_8660);
or U11682 (N_11682,N_8745,N_9336);
and U11683 (N_11683,N_9943,N_8400);
or U11684 (N_11684,N_9658,N_8164);
or U11685 (N_11685,N_9898,N_9469);
nand U11686 (N_11686,N_8010,N_9542);
or U11687 (N_11687,N_8406,N_8127);
or U11688 (N_11688,N_9744,N_8986);
nand U11689 (N_11689,N_9247,N_9628);
and U11690 (N_11690,N_8030,N_9662);
or U11691 (N_11691,N_9902,N_9588);
nor U11692 (N_11692,N_9760,N_8160);
nand U11693 (N_11693,N_9403,N_9582);
and U11694 (N_11694,N_8215,N_8513);
nor U11695 (N_11695,N_9050,N_9594);
and U11696 (N_11696,N_9715,N_8365);
xnor U11697 (N_11697,N_9884,N_9542);
nor U11698 (N_11698,N_8748,N_9008);
nor U11699 (N_11699,N_9041,N_9273);
and U11700 (N_11700,N_8945,N_8610);
and U11701 (N_11701,N_8373,N_9616);
and U11702 (N_11702,N_9940,N_8240);
nand U11703 (N_11703,N_9564,N_9624);
and U11704 (N_11704,N_9644,N_9742);
nand U11705 (N_11705,N_8331,N_8387);
xor U11706 (N_11706,N_9992,N_9879);
and U11707 (N_11707,N_8661,N_9875);
nor U11708 (N_11708,N_9221,N_9709);
nand U11709 (N_11709,N_8086,N_9773);
nand U11710 (N_11710,N_8672,N_8341);
or U11711 (N_11711,N_9222,N_9566);
nor U11712 (N_11712,N_9635,N_8241);
or U11713 (N_11713,N_9452,N_8015);
nor U11714 (N_11714,N_8196,N_8816);
or U11715 (N_11715,N_8461,N_8987);
nor U11716 (N_11716,N_9347,N_9855);
and U11717 (N_11717,N_8397,N_9403);
nand U11718 (N_11718,N_8394,N_9578);
and U11719 (N_11719,N_9617,N_8498);
nor U11720 (N_11720,N_8081,N_8852);
nand U11721 (N_11721,N_9324,N_9694);
nor U11722 (N_11722,N_9729,N_8097);
and U11723 (N_11723,N_8783,N_8870);
nand U11724 (N_11724,N_9372,N_8125);
and U11725 (N_11725,N_9283,N_9661);
and U11726 (N_11726,N_9538,N_9010);
nand U11727 (N_11727,N_8396,N_9574);
nor U11728 (N_11728,N_9821,N_8033);
nor U11729 (N_11729,N_9059,N_8570);
nor U11730 (N_11730,N_9588,N_9114);
nand U11731 (N_11731,N_8280,N_9764);
xor U11732 (N_11732,N_8080,N_8628);
and U11733 (N_11733,N_9733,N_8778);
or U11734 (N_11734,N_9984,N_9987);
nor U11735 (N_11735,N_9392,N_9857);
nor U11736 (N_11736,N_8638,N_8860);
nor U11737 (N_11737,N_9351,N_9847);
xor U11738 (N_11738,N_9218,N_9981);
or U11739 (N_11739,N_9165,N_8226);
nor U11740 (N_11740,N_9397,N_8024);
nor U11741 (N_11741,N_9723,N_8160);
nand U11742 (N_11742,N_9400,N_8179);
nor U11743 (N_11743,N_9372,N_9593);
or U11744 (N_11744,N_9087,N_8960);
and U11745 (N_11745,N_8537,N_8706);
or U11746 (N_11746,N_8302,N_9289);
xor U11747 (N_11747,N_9567,N_9159);
xor U11748 (N_11748,N_8116,N_8185);
nor U11749 (N_11749,N_8812,N_8826);
and U11750 (N_11750,N_9866,N_8611);
nand U11751 (N_11751,N_8393,N_8722);
xnor U11752 (N_11752,N_9261,N_8499);
nor U11753 (N_11753,N_9248,N_9736);
and U11754 (N_11754,N_9825,N_8154);
or U11755 (N_11755,N_9290,N_8932);
nor U11756 (N_11756,N_8217,N_8869);
nand U11757 (N_11757,N_9704,N_8609);
nor U11758 (N_11758,N_8079,N_9774);
nand U11759 (N_11759,N_8414,N_9531);
and U11760 (N_11760,N_8339,N_8507);
or U11761 (N_11761,N_9810,N_9983);
or U11762 (N_11762,N_9517,N_8784);
or U11763 (N_11763,N_8227,N_9182);
and U11764 (N_11764,N_8872,N_9972);
nor U11765 (N_11765,N_9137,N_8969);
or U11766 (N_11766,N_9951,N_8918);
xor U11767 (N_11767,N_9213,N_8820);
or U11768 (N_11768,N_9010,N_9257);
or U11769 (N_11769,N_8332,N_9878);
nand U11770 (N_11770,N_8344,N_9239);
or U11771 (N_11771,N_8569,N_9905);
nand U11772 (N_11772,N_8278,N_9225);
or U11773 (N_11773,N_9116,N_9337);
nor U11774 (N_11774,N_8935,N_8977);
and U11775 (N_11775,N_9902,N_9815);
or U11776 (N_11776,N_9198,N_9300);
nor U11777 (N_11777,N_8854,N_9097);
nand U11778 (N_11778,N_8986,N_9194);
nand U11779 (N_11779,N_8373,N_9060);
or U11780 (N_11780,N_9077,N_9832);
and U11781 (N_11781,N_9970,N_9725);
or U11782 (N_11782,N_8112,N_8981);
xor U11783 (N_11783,N_9169,N_8236);
nor U11784 (N_11784,N_8947,N_8500);
or U11785 (N_11785,N_9581,N_9393);
nor U11786 (N_11786,N_9151,N_8800);
nor U11787 (N_11787,N_9029,N_9525);
or U11788 (N_11788,N_9683,N_9496);
or U11789 (N_11789,N_8534,N_8564);
nor U11790 (N_11790,N_9180,N_9008);
nor U11791 (N_11791,N_9694,N_8148);
or U11792 (N_11792,N_8385,N_9306);
nor U11793 (N_11793,N_8059,N_8828);
or U11794 (N_11794,N_8410,N_8151);
nor U11795 (N_11795,N_9888,N_9496);
nand U11796 (N_11796,N_9829,N_9084);
nand U11797 (N_11797,N_8046,N_9243);
or U11798 (N_11798,N_8928,N_9162);
and U11799 (N_11799,N_9603,N_9532);
nor U11800 (N_11800,N_9007,N_8937);
nand U11801 (N_11801,N_8624,N_9082);
nor U11802 (N_11802,N_9674,N_8589);
and U11803 (N_11803,N_9399,N_8395);
xnor U11804 (N_11804,N_9774,N_8978);
or U11805 (N_11805,N_8297,N_8773);
or U11806 (N_11806,N_8509,N_8914);
or U11807 (N_11807,N_8313,N_9694);
nor U11808 (N_11808,N_9828,N_8955);
nor U11809 (N_11809,N_9253,N_9693);
or U11810 (N_11810,N_9569,N_8265);
and U11811 (N_11811,N_8681,N_9420);
or U11812 (N_11812,N_8912,N_8080);
and U11813 (N_11813,N_8288,N_9439);
or U11814 (N_11814,N_8936,N_9634);
nor U11815 (N_11815,N_8099,N_9736);
or U11816 (N_11816,N_9821,N_8217);
nand U11817 (N_11817,N_9014,N_8105);
or U11818 (N_11818,N_9795,N_9028);
or U11819 (N_11819,N_8933,N_9844);
nor U11820 (N_11820,N_9869,N_9327);
and U11821 (N_11821,N_9729,N_8753);
and U11822 (N_11822,N_8753,N_8609);
or U11823 (N_11823,N_8741,N_9513);
and U11824 (N_11824,N_9124,N_8567);
nand U11825 (N_11825,N_9269,N_9481);
and U11826 (N_11826,N_8005,N_8563);
or U11827 (N_11827,N_9744,N_9536);
nor U11828 (N_11828,N_9047,N_8624);
xnor U11829 (N_11829,N_9533,N_9715);
and U11830 (N_11830,N_9315,N_8746);
nor U11831 (N_11831,N_8963,N_8129);
nand U11832 (N_11832,N_9066,N_9883);
and U11833 (N_11833,N_8632,N_8571);
or U11834 (N_11834,N_9997,N_8160);
or U11835 (N_11835,N_9957,N_8602);
or U11836 (N_11836,N_9840,N_8891);
nand U11837 (N_11837,N_9954,N_9781);
and U11838 (N_11838,N_9848,N_8294);
nand U11839 (N_11839,N_8614,N_9459);
and U11840 (N_11840,N_9980,N_8768);
or U11841 (N_11841,N_8747,N_9326);
and U11842 (N_11842,N_8944,N_8601);
xor U11843 (N_11843,N_8727,N_9073);
or U11844 (N_11844,N_9953,N_9317);
and U11845 (N_11845,N_8582,N_9388);
nor U11846 (N_11846,N_8964,N_9205);
or U11847 (N_11847,N_9213,N_9534);
and U11848 (N_11848,N_8714,N_9597);
and U11849 (N_11849,N_8596,N_8185);
and U11850 (N_11850,N_8175,N_8169);
nand U11851 (N_11851,N_9373,N_8243);
nor U11852 (N_11852,N_8270,N_8233);
xnor U11853 (N_11853,N_9357,N_8648);
nand U11854 (N_11854,N_9050,N_9978);
or U11855 (N_11855,N_9406,N_8451);
and U11856 (N_11856,N_8191,N_8404);
or U11857 (N_11857,N_8997,N_9808);
nand U11858 (N_11858,N_9560,N_8086);
nor U11859 (N_11859,N_9643,N_8664);
nand U11860 (N_11860,N_9372,N_8775);
and U11861 (N_11861,N_9604,N_9517);
and U11862 (N_11862,N_8602,N_8606);
and U11863 (N_11863,N_9843,N_9549);
or U11864 (N_11864,N_9429,N_9650);
nor U11865 (N_11865,N_9934,N_8032);
xnor U11866 (N_11866,N_9958,N_9653);
or U11867 (N_11867,N_8075,N_9744);
and U11868 (N_11868,N_8728,N_8011);
and U11869 (N_11869,N_9213,N_9110);
nand U11870 (N_11870,N_8383,N_8258);
nand U11871 (N_11871,N_9040,N_8635);
nor U11872 (N_11872,N_9093,N_9016);
xor U11873 (N_11873,N_8767,N_8711);
or U11874 (N_11874,N_8994,N_8144);
or U11875 (N_11875,N_9861,N_9255);
nand U11876 (N_11876,N_9958,N_9117);
and U11877 (N_11877,N_8539,N_9075);
nor U11878 (N_11878,N_9737,N_9986);
nor U11879 (N_11879,N_9257,N_9650);
and U11880 (N_11880,N_9127,N_8705);
xor U11881 (N_11881,N_9389,N_8861);
nand U11882 (N_11882,N_8145,N_8314);
nand U11883 (N_11883,N_9600,N_9444);
or U11884 (N_11884,N_9236,N_9055);
nor U11885 (N_11885,N_8776,N_9536);
xnor U11886 (N_11886,N_8863,N_8497);
and U11887 (N_11887,N_9097,N_8623);
and U11888 (N_11888,N_8745,N_9078);
nor U11889 (N_11889,N_9084,N_9431);
or U11890 (N_11890,N_8267,N_8281);
nand U11891 (N_11891,N_8092,N_8155);
and U11892 (N_11892,N_9966,N_8052);
or U11893 (N_11893,N_9956,N_8873);
nand U11894 (N_11894,N_9864,N_8415);
xor U11895 (N_11895,N_9299,N_9052);
nor U11896 (N_11896,N_8658,N_9156);
or U11897 (N_11897,N_9163,N_8071);
or U11898 (N_11898,N_8144,N_9201);
or U11899 (N_11899,N_8354,N_9958);
or U11900 (N_11900,N_9548,N_9128);
nor U11901 (N_11901,N_9066,N_9838);
xnor U11902 (N_11902,N_9387,N_9718);
or U11903 (N_11903,N_8701,N_8263);
and U11904 (N_11904,N_8305,N_9163);
nor U11905 (N_11905,N_9944,N_9110);
nor U11906 (N_11906,N_9198,N_9954);
or U11907 (N_11907,N_8112,N_8404);
and U11908 (N_11908,N_9408,N_8332);
and U11909 (N_11909,N_9147,N_9094);
nor U11910 (N_11910,N_8260,N_8266);
xnor U11911 (N_11911,N_8346,N_9920);
nand U11912 (N_11912,N_9981,N_9991);
and U11913 (N_11913,N_8753,N_9688);
nor U11914 (N_11914,N_8373,N_8770);
nand U11915 (N_11915,N_9129,N_9610);
and U11916 (N_11916,N_9310,N_8459);
or U11917 (N_11917,N_9016,N_9434);
and U11918 (N_11918,N_9739,N_8290);
or U11919 (N_11919,N_9002,N_8599);
or U11920 (N_11920,N_8952,N_8817);
or U11921 (N_11921,N_8269,N_9067);
nor U11922 (N_11922,N_8542,N_8416);
xor U11923 (N_11923,N_8950,N_8149);
or U11924 (N_11924,N_8230,N_8759);
and U11925 (N_11925,N_9508,N_9032);
nand U11926 (N_11926,N_9390,N_9834);
or U11927 (N_11927,N_9424,N_8559);
or U11928 (N_11928,N_8028,N_9615);
or U11929 (N_11929,N_9670,N_8646);
or U11930 (N_11930,N_9794,N_8989);
xor U11931 (N_11931,N_8016,N_9419);
nand U11932 (N_11932,N_9195,N_8199);
nand U11933 (N_11933,N_9634,N_8281);
or U11934 (N_11934,N_8240,N_8054);
or U11935 (N_11935,N_9279,N_9709);
or U11936 (N_11936,N_9985,N_9108);
nor U11937 (N_11937,N_9808,N_8057);
or U11938 (N_11938,N_9461,N_9764);
or U11939 (N_11939,N_8440,N_8108);
nor U11940 (N_11940,N_9054,N_9078);
nand U11941 (N_11941,N_8035,N_8750);
nand U11942 (N_11942,N_9980,N_9770);
nand U11943 (N_11943,N_8195,N_8259);
or U11944 (N_11944,N_9641,N_8986);
and U11945 (N_11945,N_8073,N_9877);
and U11946 (N_11946,N_9611,N_8244);
nand U11947 (N_11947,N_8047,N_9728);
xnor U11948 (N_11948,N_8971,N_9461);
and U11949 (N_11949,N_9148,N_8644);
or U11950 (N_11950,N_8239,N_8912);
nor U11951 (N_11951,N_9054,N_9975);
xnor U11952 (N_11952,N_8755,N_8262);
nor U11953 (N_11953,N_9101,N_9287);
or U11954 (N_11954,N_9478,N_9744);
xnor U11955 (N_11955,N_8856,N_8120);
nor U11956 (N_11956,N_9500,N_9970);
or U11957 (N_11957,N_8669,N_9067);
nand U11958 (N_11958,N_8887,N_9057);
nand U11959 (N_11959,N_9392,N_8113);
nor U11960 (N_11960,N_8574,N_9683);
or U11961 (N_11961,N_8126,N_9184);
xor U11962 (N_11962,N_8737,N_8330);
nor U11963 (N_11963,N_8871,N_9643);
nand U11964 (N_11964,N_9046,N_9963);
nor U11965 (N_11965,N_9072,N_8188);
or U11966 (N_11966,N_9810,N_9091);
nand U11967 (N_11967,N_9570,N_8291);
and U11968 (N_11968,N_9298,N_9268);
and U11969 (N_11969,N_8836,N_8714);
and U11970 (N_11970,N_9789,N_8128);
nand U11971 (N_11971,N_9223,N_9555);
and U11972 (N_11972,N_9319,N_9869);
or U11973 (N_11973,N_8410,N_8208);
and U11974 (N_11974,N_9904,N_8642);
nor U11975 (N_11975,N_9792,N_8035);
nand U11976 (N_11976,N_8093,N_9498);
nand U11977 (N_11977,N_8082,N_9068);
or U11978 (N_11978,N_8547,N_9613);
and U11979 (N_11979,N_9356,N_9959);
or U11980 (N_11980,N_8888,N_8456);
and U11981 (N_11981,N_8811,N_9429);
xor U11982 (N_11982,N_9951,N_9650);
or U11983 (N_11983,N_9518,N_9052);
nor U11984 (N_11984,N_8148,N_9471);
and U11985 (N_11985,N_8723,N_8190);
and U11986 (N_11986,N_9356,N_8148);
and U11987 (N_11987,N_8637,N_8397);
nand U11988 (N_11988,N_9769,N_9509);
and U11989 (N_11989,N_9986,N_9361);
or U11990 (N_11990,N_8881,N_8001);
nand U11991 (N_11991,N_8970,N_8209);
xnor U11992 (N_11992,N_9549,N_9822);
or U11993 (N_11993,N_8231,N_9388);
nor U11994 (N_11994,N_8770,N_8157);
nor U11995 (N_11995,N_9222,N_9383);
xnor U11996 (N_11996,N_8742,N_9559);
nand U11997 (N_11997,N_9990,N_9863);
or U11998 (N_11998,N_8746,N_8900);
or U11999 (N_11999,N_9810,N_8652);
and U12000 (N_12000,N_10679,N_11922);
nand U12001 (N_12001,N_10139,N_10171);
nor U12002 (N_12002,N_10158,N_11287);
nand U12003 (N_12003,N_10697,N_11798);
nor U12004 (N_12004,N_11305,N_10882);
or U12005 (N_12005,N_11279,N_10685);
nand U12006 (N_12006,N_11396,N_10179);
or U12007 (N_12007,N_10982,N_11884);
nand U12008 (N_12008,N_11224,N_10452);
or U12009 (N_12009,N_10116,N_10612);
nand U12010 (N_12010,N_10125,N_11523);
nand U12011 (N_12011,N_11852,N_11945);
xnor U12012 (N_12012,N_11119,N_10188);
nor U12013 (N_12013,N_11792,N_10665);
xnor U12014 (N_12014,N_10102,N_11465);
and U12015 (N_12015,N_11032,N_11811);
nand U12016 (N_12016,N_10716,N_11069);
and U12017 (N_12017,N_11607,N_11347);
nor U12018 (N_12018,N_11251,N_10199);
nand U12019 (N_12019,N_11961,N_10549);
and U12020 (N_12020,N_10531,N_10253);
and U12021 (N_12021,N_10178,N_11797);
nand U12022 (N_12022,N_10321,N_11664);
nand U12023 (N_12023,N_11901,N_10114);
or U12024 (N_12024,N_10422,N_11947);
nor U12025 (N_12025,N_11550,N_11856);
nand U12026 (N_12026,N_11848,N_10820);
and U12027 (N_12027,N_11565,N_11991);
nand U12028 (N_12028,N_11244,N_11053);
nand U12029 (N_12029,N_11990,N_10790);
or U12030 (N_12030,N_10216,N_11660);
nor U12031 (N_12031,N_11923,N_10985);
or U12032 (N_12032,N_11615,N_10659);
or U12033 (N_12033,N_11822,N_10758);
nor U12034 (N_12034,N_11042,N_11795);
or U12035 (N_12035,N_11059,N_11268);
xnor U12036 (N_12036,N_11013,N_11681);
and U12037 (N_12037,N_10973,N_10807);
nor U12038 (N_12038,N_11211,N_10718);
nor U12039 (N_12039,N_11579,N_10595);
nor U12040 (N_12040,N_11734,N_11161);
nand U12041 (N_12041,N_11238,N_11919);
nand U12042 (N_12042,N_10104,N_11432);
nor U12043 (N_12043,N_11930,N_10954);
nor U12044 (N_12044,N_11446,N_10379);
or U12045 (N_12045,N_10023,N_10992);
nor U12046 (N_12046,N_11235,N_10359);
nor U12047 (N_12047,N_10911,N_11997);
xor U12048 (N_12048,N_10100,N_10852);
nand U12049 (N_12049,N_11541,N_11704);
or U12050 (N_12050,N_10515,N_11338);
nand U12051 (N_12051,N_11916,N_11584);
nand U12052 (N_12052,N_10305,N_10520);
nand U12053 (N_12053,N_11241,N_10941);
and U12054 (N_12054,N_10785,N_10907);
nor U12055 (N_12055,N_10480,N_10996);
or U12056 (N_12056,N_10356,N_10908);
and U12057 (N_12057,N_11685,N_10621);
nand U12058 (N_12058,N_10817,N_10878);
and U12059 (N_12059,N_11767,N_10172);
and U12060 (N_12060,N_11741,N_10898);
nor U12061 (N_12061,N_11184,N_11789);
nand U12062 (N_12062,N_10150,N_11989);
and U12063 (N_12063,N_10358,N_11199);
and U12064 (N_12064,N_11146,N_11124);
nand U12065 (N_12065,N_11783,N_10101);
or U12066 (N_12066,N_10486,N_11849);
nand U12067 (N_12067,N_10344,N_10195);
nor U12068 (N_12068,N_11622,N_10768);
and U12069 (N_12069,N_11967,N_11526);
or U12070 (N_12070,N_10862,N_11955);
and U12071 (N_12071,N_10582,N_10575);
or U12072 (N_12072,N_10489,N_11495);
nand U12073 (N_12073,N_10748,N_11595);
or U12074 (N_12074,N_10826,N_11179);
and U12075 (N_12075,N_10162,N_11599);
or U12076 (N_12076,N_11344,N_10956);
nor U12077 (N_12077,N_11556,N_11654);
xnor U12078 (N_12078,N_11571,N_10970);
nor U12079 (N_12079,N_10739,N_11312);
and U12080 (N_12080,N_10066,N_10279);
and U12081 (N_12081,N_11727,N_11775);
and U12082 (N_12082,N_11477,N_10299);
and U12083 (N_12083,N_10043,N_11794);
nor U12084 (N_12084,N_11838,N_10666);
and U12085 (N_12085,N_10326,N_11158);
and U12086 (N_12086,N_11038,N_11826);
and U12087 (N_12087,N_10792,N_11005);
nand U12088 (N_12088,N_10075,N_10008);
nand U12089 (N_12089,N_10459,N_10581);
nor U12090 (N_12090,N_10533,N_11024);
or U12091 (N_12091,N_11330,N_10387);
nor U12092 (N_12092,N_10057,N_11230);
xor U12093 (N_12093,N_10141,N_11958);
and U12094 (N_12094,N_10444,N_11953);
and U12095 (N_12095,N_10889,N_10461);
nor U12096 (N_12096,N_11335,N_11083);
and U12097 (N_12097,N_11204,N_11263);
or U12098 (N_12098,N_11751,N_10738);
or U12099 (N_12099,N_10845,N_10926);
and U12100 (N_12100,N_11918,N_11293);
nor U12101 (N_12101,N_10841,N_10513);
and U12102 (N_12102,N_11248,N_11193);
nor U12103 (N_12103,N_11682,N_10236);
and U12104 (N_12104,N_11907,N_11129);
nand U12105 (N_12105,N_11192,N_11687);
and U12106 (N_12106,N_11484,N_10373);
nand U12107 (N_12107,N_10416,N_11318);
and U12108 (N_12108,N_10923,N_11937);
and U12109 (N_12109,N_11628,N_10784);
and U12110 (N_12110,N_10003,N_10725);
xnor U12111 (N_12111,N_10977,N_11208);
nor U12112 (N_12112,N_11392,N_11698);
nand U12113 (N_12113,N_10537,N_11650);
xnor U12114 (N_12114,N_10498,N_10564);
and U12115 (N_12115,N_10747,N_10890);
nor U12116 (N_12116,N_10028,N_10746);
and U12117 (N_12117,N_11610,N_11168);
nand U12118 (N_12118,N_10056,N_10225);
or U12119 (N_12119,N_11864,N_11639);
or U12120 (N_12120,N_10756,N_11017);
or U12121 (N_12121,N_10558,N_10834);
nor U12122 (N_12122,N_10511,N_11067);
nor U12123 (N_12123,N_11706,N_10660);
nor U12124 (N_12124,N_11957,N_11411);
nor U12125 (N_12125,N_11466,N_10074);
or U12126 (N_12126,N_11755,N_11434);
nand U12127 (N_12127,N_10302,N_11536);
and U12128 (N_12128,N_11941,N_10385);
nor U12129 (N_12129,N_10163,N_10546);
nand U12130 (N_12130,N_10363,N_10080);
nand U12131 (N_12131,N_11212,N_10384);
nand U12132 (N_12132,N_10005,N_10556);
xor U12133 (N_12133,N_11342,N_10068);
and U12134 (N_12134,N_11505,N_11225);
nand U12135 (N_12135,N_10691,N_10092);
nand U12136 (N_12136,N_10935,N_11090);
or U12137 (N_12137,N_10978,N_11878);
nand U12138 (N_12138,N_10257,N_10041);
xor U12139 (N_12139,N_10534,N_10512);
nand U12140 (N_12140,N_11563,N_10181);
nor U12141 (N_12141,N_10953,N_10223);
or U12142 (N_12142,N_11135,N_10979);
nand U12143 (N_12143,N_10864,N_11463);
and U12144 (N_12144,N_10069,N_11290);
xnor U12145 (N_12145,N_11637,N_11606);
nand U12146 (N_12146,N_10110,N_10336);
nand U12147 (N_12147,N_10667,N_11012);
or U12148 (N_12148,N_11104,N_11334);
or U12149 (N_12149,N_11869,N_10166);
or U12150 (N_12150,N_10270,N_11060);
nor U12151 (N_12151,N_10500,N_11868);
or U12152 (N_12152,N_10990,N_10504);
or U12153 (N_12153,N_11862,N_11167);
or U12154 (N_12154,N_10961,N_10588);
xnor U12155 (N_12155,N_11617,N_10428);
nand U12156 (N_12156,N_11044,N_11814);
nand U12157 (N_12157,N_10983,N_10352);
nor U12158 (N_12158,N_10087,N_10340);
or U12159 (N_12159,N_10316,N_10076);
nor U12160 (N_12160,N_11236,N_10773);
and U12161 (N_12161,N_11623,N_11968);
nand U12162 (N_12162,N_11420,N_11883);
xor U12163 (N_12163,N_11793,N_10433);
nor U12164 (N_12164,N_11596,N_11367);
nand U12165 (N_12165,N_10620,N_10629);
and U12166 (N_12166,N_11162,N_10369);
and U12167 (N_12167,N_10154,N_10813);
nand U12168 (N_12168,N_10070,N_11631);
nand U12169 (N_12169,N_10847,N_10176);
xnor U12170 (N_12170,N_10222,N_11562);
or U12171 (N_12171,N_11742,N_11640);
nor U12172 (N_12172,N_10276,N_10951);
xnor U12173 (N_12173,N_10699,N_10338);
nor U12174 (N_12174,N_10728,N_11075);
nand U12175 (N_12175,N_10371,N_11252);
and U12176 (N_12176,N_11188,N_11450);
or U12177 (N_12177,N_11289,N_10891);
xor U12178 (N_12178,N_10020,N_10776);
and U12179 (N_12179,N_11871,N_10925);
or U12180 (N_12180,N_11944,N_11790);
and U12181 (N_12181,N_11616,N_11581);
nand U12182 (N_12182,N_11286,N_10200);
nand U12183 (N_12183,N_11394,N_11813);
and U12184 (N_12184,N_10732,N_11999);
nor U12185 (N_12185,N_11406,N_11771);
or U12186 (N_12186,N_10849,N_10083);
nor U12187 (N_12187,N_11532,N_11476);
nor U12188 (N_12188,N_11904,N_10378);
and U12189 (N_12189,N_11243,N_10330);
and U12190 (N_12190,N_11048,N_10895);
and U12191 (N_12191,N_10710,N_10314);
or U12192 (N_12192,N_10458,N_10372);
nor U12193 (N_12193,N_10475,N_10910);
nor U12194 (N_12194,N_11041,N_10945);
xnor U12195 (N_12195,N_10532,N_10243);
and U12196 (N_12196,N_10542,N_11545);
nor U12197 (N_12197,N_10399,N_10196);
and U12198 (N_12198,N_10551,N_10774);
or U12199 (N_12199,N_11982,N_10840);
nor U12200 (N_12200,N_11386,N_11850);
or U12201 (N_12201,N_11732,N_11121);
nand U12202 (N_12202,N_10654,N_11739);
and U12203 (N_12203,N_10467,N_11511);
nor U12204 (N_12204,N_10980,N_11084);
and U12205 (N_12205,N_10212,N_10850);
and U12206 (N_12206,N_11490,N_11159);
and U12207 (N_12207,N_11352,N_10194);
xor U12208 (N_12208,N_10942,N_10191);
nor U12209 (N_12209,N_10800,N_10674);
and U12210 (N_12210,N_11554,N_11035);
or U12211 (N_12211,N_10788,N_11353);
and U12212 (N_12212,N_10055,N_11102);
nor U12213 (N_12213,N_10355,N_11309);
nand U12214 (N_12214,N_11343,N_10863);
nand U12215 (N_12215,N_11875,N_11444);
and U12216 (N_12216,N_10109,N_10657);
nor U12217 (N_12217,N_10730,N_10811);
and U12218 (N_12218,N_11418,N_11542);
or U12219 (N_12219,N_10259,N_10397);
nor U12220 (N_12220,N_10692,N_10038);
nand U12221 (N_12221,N_10569,N_11061);
or U12222 (N_12222,N_11058,N_10888);
nand U12223 (N_12223,N_11171,N_10086);
nor U12224 (N_12224,N_10409,N_11592);
and U12225 (N_12225,N_10616,N_11026);
nor U12226 (N_12226,N_11578,N_10887);
nor U12227 (N_12227,N_10830,N_11488);
xor U12228 (N_12228,N_10142,N_11777);
nor U12229 (N_12229,N_11151,N_11717);
nand U12230 (N_12230,N_11298,N_11614);
nor U12231 (N_12231,N_10204,N_11594);
nand U12232 (N_12232,N_11763,N_10345);
or U12233 (N_12233,N_10376,N_11210);
nor U12234 (N_12234,N_11003,N_10389);
nor U12235 (N_12235,N_11697,N_10587);
xor U12236 (N_12236,N_11667,N_11952);
or U12237 (N_12237,N_10851,N_10445);
or U12238 (N_12238,N_11454,N_10866);
nand U12239 (N_12239,N_11770,N_10280);
xnor U12240 (N_12240,N_10708,N_10117);
and U12241 (N_12241,N_10735,N_11395);
nand U12242 (N_12242,N_10555,N_10391);
nand U12243 (N_12243,N_11802,N_11576);
xnor U12244 (N_12244,N_11835,N_11521);
nor U12245 (N_12245,N_11683,N_10234);
nor U12246 (N_12246,N_11841,N_10468);
xor U12247 (N_12247,N_10062,N_11984);
nor U12248 (N_12248,N_11675,N_10174);
nand U12249 (N_12249,N_10205,N_11321);
nor U12250 (N_12250,N_11625,N_10880);
and U12251 (N_12251,N_10221,N_10192);
xnor U12252 (N_12252,N_11206,N_10957);
xor U12253 (N_12253,N_10170,N_10897);
and U12254 (N_12254,N_10173,N_10939);
or U12255 (N_12255,N_11470,N_10917);
and U12256 (N_12256,N_10476,N_10896);
and U12257 (N_12257,N_10869,N_11361);
and U12258 (N_12258,N_10411,N_11045);
nor U12259 (N_12259,N_11401,N_10916);
or U12260 (N_12260,N_10715,N_10599);
nor U12261 (N_12261,N_10698,N_11949);
or U12262 (N_12262,N_10517,N_11220);
nand U12263 (N_12263,N_10095,N_10541);
nor U12264 (N_12264,N_10169,N_10250);
xor U12265 (N_12265,N_11823,N_10669);
xnor U12266 (N_12266,N_11668,N_11034);
nand U12267 (N_12267,N_11141,N_11340);
or U12268 (N_12268,N_10443,N_11138);
xor U12269 (N_12269,N_11057,N_10473);
nand U12270 (N_12270,N_11331,N_11014);
and U12271 (N_12271,N_10318,N_11493);
and U12272 (N_12272,N_10606,N_11265);
nand U12273 (N_12273,N_11339,N_10677);
xor U12274 (N_12274,N_11326,N_10272);
nor U12275 (N_12275,N_11388,N_10543);
nand U12276 (N_12276,N_10596,N_10510);
nor U12277 (N_12277,N_11501,N_10161);
nor U12278 (N_12278,N_10012,N_11445);
xnor U12279 (N_12279,N_10947,N_11147);
and U12280 (N_12280,N_11665,N_11890);
nand U12281 (N_12281,N_11183,N_11633);
nand U12282 (N_12282,N_11085,N_10632);
nor U12283 (N_12283,N_11588,N_11707);
and U12284 (N_12284,N_11266,N_10044);
nor U12285 (N_12285,N_11936,N_11711);
nand U12286 (N_12286,N_11538,N_11604);
and U12287 (N_12287,N_11002,N_11986);
xnor U12288 (N_12288,N_11087,N_11929);
or U12289 (N_12289,N_11106,N_11441);
and U12290 (N_12290,N_11605,N_10529);
nand U12291 (N_12291,N_11063,N_11173);
or U12292 (N_12292,N_11859,N_11376);
or U12293 (N_12293,N_10454,N_11701);
nor U12294 (N_12294,N_10334,N_10392);
and U12295 (N_12295,N_11296,N_11357);
nand U12296 (N_12296,N_11653,N_11166);
and U12297 (N_12297,N_10915,N_10576);
or U12298 (N_12298,N_11139,N_11978);
nand U12299 (N_12299,N_10207,N_10165);
nor U12300 (N_12300,N_10837,N_11421);
nor U12301 (N_12301,N_10635,N_10427);
nand U12302 (N_12302,N_11776,N_11245);
or U12303 (N_12303,N_10563,N_11229);
nor U12304 (N_12304,N_10812,N_11174);
nor U12305 (N_12305,N_10557,N_10655);
nand U12306 (N_12306,N_11079,N_10782);
nor U12307 (N_12307,N_10337,N_11165);
xor U12308 (N_12308,N_10821,N_11863);
xnor U12309 (N_12309,N_11692,N_10554);
nor U12310 (N_12310,N_10112,N_10600);
and U12311 (N_12311,N_10810,N_10304);
xor U12312 (N_12312,N_11377,N_10877);
or U12313 (N_12313,N_10932,N_11384);
nand U12314 (N_12314,N_10430,N_10501);
and U12315 (N_12315,N_11496,N_11479);
or U12316 (N_12316,N_11773,N_11825);
nor U12317 (N_12317,N_10091,N_10783);
nor U12318 (N_12318,N_11010,N_11127);
and U12319 (N_12319,N_11663,N_11935);
nor U12320 (N_12320,N_11435,N_10122);
or U12321 (N_12321,N_10856,N_11708);
or U12322 (N_12322,N_11438,N_11757);
nand U12323 (N_12323,N_11729,N_11155);
and U12324 (N_12324,N_11283,N_11720);
nand U12325 (N_12325,N_10309,N_10435);
nand U12326 (N_12326,N_10137,N_11148);
nor U12327 (N_12327,N_10663,N_10843);
xnor U12328 (N_12328,N_11738,N_11927);
nand U12329 (N_12329,N_11055,N_11422);
or U12330 (N_12330,N_11867,N_10108);
or U12331 (N_12331,N_10607,N_10668);
nand U12332 (N_12332,N_11761,N_10146);
xnor U12333 (N_12333,N_10107,N_11200);
nor U12334 (N_12334,N_10022,N_10651);
nand U12335 (N_12335,N_10502,N_10333);
nor U12336 (N_12336,N_10140,N_10871);
and U12337 (N_12337,N_10085,N_11679);
nor U12338 (N_12338,N_10263,N_10124);
and U12339 (N_12339,N_11740,N_10421);
and U12340 (N_12340,N_10567,N_11855);
or U12341 (N_12341,N_11626,N_11943);
nor U12342 (N_12342,N_11191,N_11194);
nor U12343 (N_12343,N_10943,N_11695);
nand U12344 (N_12344,N_10151,N_10902);
nor U12345 (N_12345,N_11497,N_11915);
nand U12346 (N_12346,N_11844,N_10870);
and U12347 (N_12347,N_11702,N_11804);
and U12348 (N_12348,N_10293,N_10670);
or U12349 (N_12349,N_11749,N_10471);
and U12350 (N_12350,N_11602,N_10374);
or U12351 (N_12351,N_11934,N_11355);
and U12352 (N_12352,N_11778,N_11591);
nor U12353 (N_12353,N_11924,N_10335);
and U12354 (N_12354,N_10781,N_11994);
or U12355 (N_12355,N_10465,N_11509);
or U12356 (N_12356,N_10254,N_11673);
or U12357 (N_12357,N_10721,N_10009);
nor U12358 (N_12358,N_10865,N_11100);
nor U12359 (N_12359,N_10548,N_11369);
nand U12360 (N_12360,N_10235,N_10661);
or U12361 (N_12361,N_10455,N_10818);
or U12362 (N_12362,N_10760,N_11115);
or U12363 (N_12363,N_11025,N_10120);
or U12364 (N_12364,N_11328,N_10129);
nand U12365 (N_12365,N_10573,N_11195);
nor U12366 (N_12366,N_10159,N_10297);
nand U12367 (N_12367,N_10252,N_10545);
and U12368 (N_12368,N_10743,N_11471);
xnor U12369 (N_12369,N_10462,N_10904);
nand U12370 (N_12370,N_11282,N_11970);
and U12371 (N_12371,N_10929,N_10988);
nand U12372 (N_12372,N_11082,N_10088);
xor U12373 (N_12373,N_11264,N_10368);
nor U12374 (N_12374,N_10245,N_10641);
or U12375 (N_12375,N_10719,N_11068);
and U12376 (N_12376,N_11537,N_10571);
nor U12377 (N_12377,N_11072,N_10255);
nor U12378 (N_12378,N_11891,N_10625);
or U12379 (N_12379,N_10779,N_11762);
xnor U12380 (N_12380,N_11428,N_10029);
nor U12381 (N_12381,N_11215,N_11834);
nor U12382 (N_12382,N_10019,N_11782);
nor U12383 (N_12383,N_11791,N_11391);
nor U12384 (N_12384,N_10793,N_10404);
or U12385 (N_12385,N_10410,N_10364);
and U12386 (N_12386,N_10496,N_10182);
or U12387 (N_12387,N_11066,N_10271);
or U12388 (N_12388,N_10342,N_11996);
nor U12389 (N_12389,N_11051,N_10282);
xnor U12390 (N_12390,N_10965,N_10395);
nor U12391 (N_12391,N_10562,N_10283);
or U12392 (N_12392,N_11513,N_10247);
nand U12393 (N_12393,N_10138,N_11319);
nor U12394 (N_12394,N_11921,N_11725);
or U12395 (N_12395,N_11015,N_11661);
nand U12396 (N_12396,N_11586,N_11424);
nand U12397 (N_12397,N_10126,N_11004);
nand U12398 (N_12398,N_10906,N_11568);
nor U12399 (N_12399,N_10523,N_11569);
and U12400 (N_12400,N_11656,N_10396);
and U12401 (N_12401,N_10042,N_10197);
nand U12402 (N_12402,N_10806,N_10883);
or U12403 (N_12403,N_11570,N_10975);
and U12404 (N_12404,N_10997,N_11888);
nand U12405 (N_12405,N_10727,N_11735);
and U12406 (N_12406,N_10366,N_11574);
or U12407 (N_12407,N_10959,N_10298);
nor U12408 (N_12408,N_10365,N_11203);
or U12409 (N_12409,N_10361,N_10998);
xor U12410 (N_12410,N_11154,N_10002);
nor U12411 (N_12411,N_10367,N_11081);
and U12412 (N_12412,N_11690,N_11504);
and U12413 (N_12413,N_11239,N_11178);
nand U12414 (N_12414,N_10647,N_10025);
nand U12415 (N_12415,N_11436,N_10754);
nor U12416 (N_12416,N_10689,N_10325);
or U12417 (N_12417,N_10561,N_11327);
nor U12418 (N_12418,N_11381,N_11197);
xnor U12419 (N_12419,N_11976,N_10287);
nor U12420 (N_12420,N_10604,N_10672);
nand U12421 (N_12421,N_10791,N_10375);
or U12422 (N_12422,N_11294,N_10819);
xnor U12423 (N_12423,N_10412,N_11107);
and U12424 (N_12424,N_11828,N_10742);
nor U12425 (N_12425,N_11295,N_11145);
xnor U12426 (N_12426,N_10936,N_10265);
nor U12427 (N_12427,N_11877,N_11096);
nor U12428 (N_12428,N_11582,N_10099);
and U12429 (N_12429,N_11311,N_11905);
nor U12430 (N_12430,N_11817,N_11644);
or U12431 (N_12431,N_11801,N_11473);
or U12432 (N_12432,N_11387,N_11860);
nand U12433 (N_12433,N_10553,N_11910);
nand U12434 (N_12434,N_10798,N_10963);
and U12435 (N_12435,N_11858,N_10522);
and U12436 (N_12436,N_11756,N_10823);
and U12437 (N_12437,N_11443,N_10351);
nor U12438 (N_12438,N_11979,N_10406);
or U12439 (N_12439,N_10853,N_11472);
nor U12440 (N_12440,N_10426,N_11985);
nand U12441 (N_12441,N_11152,N_11299);
nand U12442 (N_12442,N_10772,N_10483);
nor U12443 (N_12443,N_11112,N_10780);
nor U12444 (N_12444,N_10180,N_11360);
xor U12445 (N_12445,N_11525,N_11468);
or U12446 (N_12446,N_10268,N_10921);
nand U12447 (N_12447,N_10627,N_10722);
or U12448 (N_12448,N_10652,N_10815);
and U12449 (N_12449,N_10229,N_10431);
xnor U12450 (N_12450,N_11950,N_10574);
or U12451 (N_12451,N_10231,N_10206);
and U12452 (N_12452,N_11078,N_11689);
or U12453 (N_12453,N_10892,N_10040);
nand U12454 (N_12454,N_11462,N_10269);
nand U12455 (N_12455,N_10566,N_10186);
nand U12456 (N_12456,N_11733,N_11678);
and U12457 (N_12457,N_11815,N_10311);
or U12458 (N_12458,N_10113,N_10673);
nand U12459 (N_12459,N_10147,N_11371);
nor U12460 (N_12460,N_11356,N_10855);
or U12461 (N_12461,N_11136,N_11250);
nand U12462 (N_12462,N_10145,N_10717);
and U12463 (N_12463,N_10063,N_10645);
and U12464 (N_12464,N_11587,N_11109);
nor U12465 (N_12465,N_11170,N_10017);
or U12466 (N_12466,N_11113,N_10696);
nor U12467 (N_12467,N_11033,N_10766);
nand U12468 (N_12468,N_10550,N_11995);
nand U12469 (N_12469,N_11840,N_10278);
nor U12470 (N_12470,N_11185,N_10777);
nor U12471 (N_12471,N_10377,N_11758);
or U12472 (N_12472,N_11634,N_10609);
and U12473 (N_12473,N_10049,N_10755);
and U12474 (N_12474,N_11306,N_10027);
and U12475 (N_12475,N_11753,N_10185);
nor U12476 (N_12476,N_11933,N_11694);
and U12477 (N_12477,N_10051,N_10347);
or U12478 (N_12478,N_11125,N_11364);
and U12479 (N_12479,N_10237,N_11442);
nand U12480 (N_12480,N_10884,N_11736);
and U12481 (N_12481,N_11419,N_11948);
or U12482 (N_12482,N_10676,N_11023);
or U12483 (N_12483,N_10745,N_11799);
and U12484 (N_12484,N_10649,N_10128);
xnor U12485 (N_12485,N_11478,N_10300);
nor U12486 (N_12486,N_11612,N_11743);
and U12487 (N_12487,N_10516,N_11226);
nor U12488 (N_12488,N_10816,N_11071);
or U12489 (N_12489,N_11691,N_10157);
and U12490 (N_12490,N_11885,N_10838);
nand U12491 (N_12491,N_11372,N_11508);
nor U12492 (N_12492,N_11564,N_11531);
or U12493 (N_12493,N_10859,N_11580);
nand U12494 (N_12494,N_11812,N_11276);
nor U12495 (N_12495,N_11142,N_11431);
and U12496 (N_12496,N_11054,N_11433);
nand U12497 (N_12497,N_11651,N_11160);
xnor U12498 (N_12498,N_11009,N_11175);
and U12499 (N_12499,N_10434,N_11029);
nand U12500 (N_12500,N_10796,N_11348);
nor U12501 (N_12501,N_11261,N_11474);
or U12502 (N_12502,N_11676,N_11108);
or U12503 (N_12503,N_11140,N_10230);
or U12504 (N_12504,N_11647,N_10519);
nor U12505 (N_12505,N_11116,N_10857);
or U12506 (N_12506,N_11832,N_11359);
and U12507 (N_12507,N_11404,N_10011);
or U12508 (N_12508,N_11280,N_10624);
or U12509 (N_12509,N_11558,N_10134);
or U12510 (N_12510,N_10492,N_11427);
or U12511 (N_12511,N_11785,N_10995);
or U12512 (N_12512,N_11713,N_11255);
nor U12513 (N_12513,N_10030,N_10922);
nor U12514 (N_12514,N_11091,N_11609);
or U12515 (N_12515,N_11964,N_10281);
or U12516 (N_12516,N_11262,N_11585);
or U12517 (N_12517,N_11959,N_10920);
or U12518 (N_12518,N_10289,N_10808);
or U12519 (N_12519,N_11894,N_11201);
nand U12520 (N_12520,N_10644,N_10803);
and U12521 (N_12521,N_11632,N_11120);
xnor U12522 (N_12522,N_10795,N_11228);
nor U12523 (N_12523,N_10643,N_10653);
and U12524 (N_12524,N_11354,N_10227);
nand U12525 (N_12525,N_11768,N_11627);
nor U12526 (N_12526,N_10438,N_10615);
nor U12527 (N_12527,N_10499,N_11040);
or U12528 (N_12528,N_10261,N_11202);
or U12529 (N_12529,N_10175,N_11567);
and U12530 (N_12530,N_11020,N_11099);
nand U12531 (N_12531,N_10702,N_11350);
or U12532 (N_12532,N_10341,N_11939);
and U12533 (N_12533,N_10054,N_10881);
or U12534 (N_12534,N_11358,N_10418);
or U12535 (N_12535,N_11560,N_11487);
nor U12536 (N_12536,N_10328,N_11819);
nand U12537 (N_12537,N_11643,N_11962);
xnor U12538 (N_12538,N_11455,N_10536);
nand U12539 (N_12539,N_11074,N_11593);
nor U12540 (N_12540,N_11169,N_11629);
nand U12541 (N_12541,N_10767,N_10061);
and U12542 (N_12542,N_11182,N_11070);
nor U12543 (N_12543,N_11399,N_10414);
nor U12544 (N_12544,N_11851,N_10695);
nand U12545 (N_12545,N_11414,N_10598);
nand U12546 (N_12546,N_10106,N_11341);
or U12547 (N_12547,N_11153,N_11385);
nor U12548 (N_12548,N_10900,N_10168);
and U12549 (N_12549,N_11983,N_10955);
xor U12550 (N_12550,N_11366,N_10429);
or U12551 (N_12551,N_10383,N_10111);
nor U12552 (N_12552,N_11400,N_10711);
or U12553 (N_12553,N_10703,N_10686);
nor U12554 (N_12554,N_11854,N_10202);
and U12555 (N_12555,N_10705,N_10241);
nand U12556 (N_12556,N_10403,N_11969);
xor U12557 (N_12557,N_10559,N_10918);
nand U12558 (N_12558,N_10353,N_10474);
or U12559 (N_12559,N_10682,N_10966);
or U12560 (N_12560,N_10634,N_11530);
and U12561 (N_12561,N_11837,N_10485);
or U12562 (N_12562,N_10589,N_11180);
xor U12563 (N_12563,N_10246,N_10687);
and U12564 (N_12564,N_10872,N_10130);
and U12565 (N_12565,N_10681,N_11575);
nor U12566 (N_12566,N_10277,N_10034);
and U12567 (N_12567,N_10420,N_10065);
nand U12568 (N_12568,N_11745,N_11143);
and U12569 (N_12569,N_10984,N_10786);
nor U12570 (N_12570,N_11429,N_10242);
and U12571 (N_12571,N_10481,N_10144);
nand U12572 (N_12572,N_11260,N_10152);
and U12573 (N_12573,N_11249,N_10301);
nor U12574 (N_12574,N_11007,N_10037);
or U12575 (N_12575,N_10805,N_10858);
nand U12576 (N_12576,N_11270,N_11423);
and U12577 (N_12577,N_11426,N_11412);
and U12578 (N_12578,N_11506,N_10233);
and U12579 (N_12579,N_11437,N_10183);
xnor U12580 (N_12580,N_10733,N_10714);
nand U12581 (N_12581,N_10630,N_10944);
nor U12582 (N_12582,N_10622,N_10933);
and U12583 (N_12583,N_10210,N_10209);
or U12584 (N_12584,N_11598,N_11784);
nor U12585 (N_12585,N_10382,N_11365);
nand U12586 (N_12586,N_11351,N_11889);
or U12587 (N_12587,N_11095,N_10464);
and U12588 (N_12588,N_11413,N_11666);
nand U12589 (N_12589,N_11908,N_11464);
nor U12590 (N_12590,N_10081,N_11512);
and U12591 (N_12591,N_11769,N_11754);
nor U12592 (N_12592,N_11449,N_11274);
and U12593 (N_12593,N_10240,N_11719);
nor U12594 (N_12594,N_10605,N_11900);
nand U12595 (N_12595,N_10931,N_11402);
nor U12596 (N_12596,N_11130,N_10286);
nor U12597 (N_12597,N_11920,N_10577);
or U12598 (N_12598,N_10690,N_10741);
nor U12599 (N_12599,N_11648,N_10115);
and U12600 (N_12600,N_10000,N_11577);
and U12601 (N_12601,N_11094,N_11006);
and U12602 (N_12602,N_10494,N_11809);
or U12603 (N_12603,N_11323,N_10879);
xor U12604 (N_12604,N_11325,N_10618);
nor U12605 (N_12605,N_10224,N_10319);
or U12606 (N_12606,N_11942,N_10761);
or U12607 (N_12607,N_10423,N_11552);
and U12608 (N_12608,N_11672,N_11917);
nand U12609 (N_12609,N_10976,N_11103);
and U12610 (N_12610,N_11642,N_11886);
and U12611 (N_12611,N_10704,N_11275);
nand U12612 (N_12612,N_10131,N_11737);
nand U12613 (N_12613,N_11540,N_10313);
and U12614 (N_12614,N_10078,N_11539);
nor U12615 (N_12615,N_11561,N_11172);
and U12616 (N_12616,N_11430,N_10950);
nand U12617 (N_12617,N_11253,N_10839);
nor U12618 (N_12618,N_10320,N_11382);
nand U12619 (N_12619,N_11721,N_10380);
nand U12620 (N_12620,N_10912,N_10193);
or U12621 (N_12621,N_11963,N_11214);
nor U12622 (N_12622,N_11134,N_11903);
nor U12623 (N_12623,N_11726,N_10460);
or U12624 (N_12624,N_10927,N_10032);
or U12625 (N_12625,N_11489,N_11684);
nor U12626 (N_12626,N_11881,N_11345);
nor U12627 (N_12627,N_11895,N_11873);
or U12628 (N_12628,N_11601,N_11774);
nand U12629 (N_12629,N_10968,N_10160);
nand U12630 (N_12630,N_11049,N_11416);
and U12631 (N_12631,N_11073,N_10084);
or U12632 (N_12632,N_10528,N_11329);
or U12633 (N_12633,N_10093,N_10794);
nor U12634 (N_12634,N_11649,N_10357);
xor U12635 (N_12635,N_10439,N_11398);
nor U12636 (N_12636,N_11149,N_10327);
nor U12637 (N_12637,N_11780,N_10628);
nand U12638 (N_12638,N_11619,N_11370);
and U12639 (N_12639,N_11256,N_10981);
nand U12640 (N_12640,N_10343,N_10349);
nand U12641 (N_12641,N_10713,N_11213);
nand U12642 (N_12642,N_11829,N_10348);
and U12643 (N_12643,N_11218,N_11544);
and U12644 (N_12644,N_10258,N_10765);
or U12645 (N_12645,N_10213,N_10388);
nand U12646 (N_12646,N_10867,N_10266);
or U12647 (N_12647,N_11645,N_11808);
nand U12648 (N_12648,N_10184,N_11221);
nor U12649 (N_12649,N_10324,N_10928);
and U12650 (N_12650,N_10608,N_11310);
nand U12651 (N_12651,N_10381,N_10924);
nor U12652 (N_12652,N_11677,N_11408);
nor U12653 (N_12653,N_11548,N_11332);
nor U12654 (N_12654,N_11092,N_11240);
xor U12655 (N_12655,N_11893,N_11630);
xor U12656 (N_12656,N_10763,N_10886);
or U12657 (N_12657,N_10586,N_10132);
nand U12658 (N_12658,N_10021,N_10010);
and U12659 (N_12659,N_11980,N_11047);
and U12660 (N_12660,N_10514,N_10201);
or U12661 (N_12661,N_11658,N_10799);
and U12662 (N_12662,N_11818,N_10539);
nor U12663 (N_12663,N_11638,N_10143);
nor U12664 (N_12664,N_10457,N_11118);
and U12665 (N_12665,N_11491,N_11302);
and U12666 (N_12666,N_10974,N_11646);
and U12667 (N_12667,N_10873,N_10288);
nor U12668 (N_12668,N_10940,N_11362);
and U12669 (N_12669,N_11861,N_11635);
xor U12670 (N_12670,N_10322,N_10899);
and U12671 (N_12671,N_10119,N_11590);
nand U12672 (N_12672,N_10024,N_11998);
nand U12673 (N_12673,N_11000,N_10493);
and U12674 (N_12674,N_11709,N_10033);
nand U12675 (N_12675,N_11258,N_11805);
and U12676 (N_12676,N_11759,N_11911);
nand U12677 (N_12677,N_10291,N_11453);
nand U12678 (N_12678,N_11787,N_10013);
nand U12679 (N_12679,N_10294,N_11712);
or U12680 (N_12680,N_10611,N_11830);
nor U12681 (N_12681,N_10442,N_10836);
or U12682 (N_12682,N_11219,N_11492);
xnor U12683 (N_12683,N_10832,N_11297);
nor U12684 (N_12684,N_11516,N_10495);
nand U12685 (N_12685,N_11037,N_10913);
nor U12686 (N_12686,N_10031,N_10787);
nand U12687 (N_12687,N_10720,N_11992);
nand U12688 (N_12688,N_11016,N_10723);
nand U12689 (N_12689,N_10306,N_11527);
nor U12690 (N_12690,N_11322,N_11699);
or U12691 (N_12691,N_11234,N_10764);
and U12692 (N_12692,N_11227,N_10824);
nand U12693 (N_12693,N_11374,N_10413);
nand U12694 (N_12694,N_10967,N_11077);
xnor U12695 (N_12695,N_11451,N_11613);
or U12696 (N_12696,N_11028,N_11242);
nand U12697 (N_12697,N_10530,N_11304);
or U12698 (N_12698,N_10700,N_10015);
xnor U12699 (N_12699,N_10636,N_11460);
and U12700 (N_12700,N_11529,N_10479);
xnor U12701 (N_12701,N_10217,N_11126);
nor U12702 (N_12702,N_10453,N_11483);
nor U12703 (N_12703,N_11272,N_11368);
nand U12704 (N_12704,N_10740,N_11050);
and U12705 (N_12705,N_10570,N_10354);
and U12706 (N_12706,N_11336,N_11975);
xor U12707 (N_12707,N_11507,N_10506);
and U12708 (N_12708,N_10752,N_11960);
and U12709 (N_12709,N_11246,N_11011);
nand U12710 (N_12710,N_10436,N_10393);
nand U12711 (N_12711,N_10133,N_10903);
nand U12712 (N_12712,N_10712,N_11467);
and U12713 (N_12713,N_10469,N_10290);
nand U12714 (N_12714,N_11181,N_11233);
nand U12715 (N_12715,N_11439,N_11659);
and U12716 (N_12716,N_11528,N_10058);
and U12717 (N_12717,N_11951,N_11600);
nand U12718 (N_12718,N_11284,N_10518);
nand U12719 (N_12719,N_10658,N_10905);
and U12720 (N_12720,N_10310,N_10047);
nand U12721 (N_12721,N_10082,N_11086);
nand U12722 (N_12722,N_10308,N_11405);
nand U12723 (N_12723,N_11641,N_10408);
xor U12724 (N_12724,N_10149,N_11966);
or U12725 (N_12725,N_11553,N_10415);
or U12726 (N_12726,N_10417,N_11820);
or U12727 (N_12727,N_10312,N_10488);
and U12728 (N_12728,N_11485,N_10482);
xor U12729 (N_12729,N_10626,N_11076);
xor U12730 (N_12730,N_11974,N_10706);
nand U12731 (N_12731,N_10449,N_11724);
nand U12732 (N_12732,N_10874,N_11748);
and U12733 (N_12733,N_11292,N_11899);
nor U12734 (N_12734,N_11696,N_11988);
or U12735 (N_12735,N_10637,N_10778);
nand U12736 (N_12736,N_11052,N_10524);
or U12737 (N_12737,N_11186,N_10709);
nand U12738 (N_12738,N_10684,N_11196);
nor U12739 (N_12739,N_10267,N_10731);
nor U12740 (N_12740,N_10045,N_10478);
nor U12741 (N_12741,N_11043,N_11909);
or U12742 (N_12742,N_10284,N_10962);
nand U12743 (N_12743,N_11824,N_10707);
nor U12744 (N_12744,N_10729,N_11620);
and U12745 (N_12745,N_11946,N_10987);
and U12746 (N_12746,N_11494,N_11046);
and U12747 (N_12747,N_10831,N_11836);
nand U12748 (N_12748,N_10487,N_10249);
nand U12749 (N_12749,N_10505,N_10219);
nor U12750 (N_12750,N_11021,N_10232);
nand U12751 (N_12751,N_11499,N_10952);
and U12752 (N_12752,N_10339,N_10829);
or U12753 (N_12753,N_11475,N_11132);
or U12754 (N_12754,N_10801,N_11972);
xor U12755 (N_12755,N_11393,N_11190);
or U12756 (N_12756,N_10260,N_11397);
or U12757 (N_12757,N_11482,N_10190);
nand U12758 (N_12758,N_10680,N_10544);
or U12759 (N_12759,N_11843,N_10835);
nand U12760 (N_12760,N_11301,N_10136);
and U12761 (N_12761,N_10105,N_11914);
nand U12762 (N_12762,N_10650,N_10934);
or U12763 (N_12763,N_10508,N_10538);
or U12764 (N_12764,N_10854,N_11557);
nand U12765 (N_12765,N_10527,N_11036);
and U12766 (N_12766,N_11217,N_10509);
nand U12767 (N_12767,N_11857,N_10701);
or U12768 (N_12768,N_11803,N_10248);
nor U12769 (N_12769,N_10208,N_11440);
xor U12770 (N_12770,N_11971,N_10451);
or U12771 (N_12771,N_10762,N_11655);
or U12772 (N_12772,N_10189,N_10244);
or U12773 (N_12773,N_10472,N_11624);
or U12774 (N_12774,N_10901,N_11137);
xor U12775 (N_12775,N_10156,N_11027);
nand U12776 (N_12776,N_11380,N_11407);
nor U12777 (N_12777,N_10067,N_10583);
nand U12778 (N_12778,N_11765,N_10089);
and U12779 (N_12779,N_10228,N_10614);
nand U12780 (N_12780,N_11931,N_10994);
and U12781 (N_12781,N_10096,N_10949);
and U12782 (N_12782,N_11731,N_11001);
nand U12783 (N_12783,N_11752,N_10597);
or U12784 (N_12784,N_10894,N_11209);
and U12785 (N_12785,N_11271,N_11874);
or U12786 (N_12786,N_11898,N_11546);
nand U12787 (N_12787,N_10633,N_11417);
or U12788 (N_12788,N_11231,N_11308);
nand U12789 (N_12789,N_10050,N_10946);
nand U12790 (N_12790,N_10121,N_11498);
nand U12791 (N_12791,N_11693,N_10285);
and U12792 (N_12792,N_10833,N_10734);
nor U12793 (N_12793,N_11456,N_10503);
nor U12794 (N_12794,N_10360,N_10256);
or U12795 (N_12795,N_11566,N_10437);
or U12796 (N_12796,N_10211,N_10394);
nand U12797 (N_12797,N_11534,N_10448);
nand U12798 (N_12798,N_10639,N_10048);
nor U12799 (N_12799,N_11897,N_10678);
nand U12800 (N_12800,N_11880,N_10405);
or U12801 (N_12801,N_11008,N_10751);
nor U12802 (N_12802,N_10307,N_10971);
or U12803 (N_12803,N_10346,N_10425);
nor U12804 (N_12804,N_11117,N_11728);
nor U12805 (N_12805,N_11324,N_10007);
and U12806 (N_12806,N_10579,N_11333);
and U12807 (N_12807,N_10275,N_11018);
nand U12808 (N_12808,N_11772,N_11415);
and U12809 (N_12809,N_10664,N_11896);
nor U12810 (N_12810,N_11853,N_11486);
nor U12811 (N_12811,N_11636,N_11810);
nor U12812 (N_12812,N_10052,N_11781);
nand U12813 (N_12813,N_10547,N_11403);
nand U12814 (N_12814,N_11176,N_10187);
and U12815 (N_12815,N_11956,N_10619);
nor U12816 (N_12816,N_10590,N_11993);
nor U12817 (N_12817,N_10239,N_10757);
nand U12818 (N_12818,N_10770,N_11913);
and U12819 (N_12819,N_11547,N_11480);
nand U12820 (N_12820,N_11111,N_10675);
nand U12821 (N_12821,N_11705,N_11788);
and U12822 (N_12822,N_10560,N_10938);
nand U12823 (N_12823,N_11870,N_10930);
nand U12824 (N_12824,N_11300,N_10585);
nor U12825 (N_12825,N_11156,N_10398);
and U12826 (N_12826,N_10617,N_11912);
or U12827 (N_12827,N_10402,N_10804);
xor U12828 (N_12828,N_10103,N_10771);
or U12829 (N_12829,N_11796,N_10868);
xor U12830 (N_12830,N_10914,N_10724);
nand U12831 (N_12831,N_11288,N_10424);
or U12832 (N_12832,N_11520,N_10759);
and U12833 (N_12833,N_11458,N_11267);
nor U12834 (N_12834,N_11065,N_11123);
nor U12835 (N_12835,N_10006,N_10090);
nor U12836 (N_12836,N_10631,N_11816);
and U12837 (N_12837,N_10001,N_11062);
and U12838 (N_12838,N_10848,N_10053);
and U12839 (N_12839,N_11237,N_10466);
or U12840 (N_12840,N_11097,N_10749);
nor U12841 (N_12841,N_11669,N_10986);
nand U12842 (N_12842,N_11902,N_11410);
nand U12843 (N_12843,N_11965,N_10578);
nand U12844 (N_12844,N_11954,N_11105);
nor U12845 (N_12845,N_10602,N_11320);
nor U12846 (N_12846,N_10164,N_11621);
and U12847 (N_12847,N_10842,N_11189);
nand U12848 (N_12848,N_10802,N_11981);
xnor U12849 (N_12849,N_11887,N_11730);
and U12850 (N_12850,N_11827,N_11503);
or U12851 (N_12851,N_10432,N_11680);
or U12852 (N_12852,N_11157,N_11457);
nor U12853 (N_12853,N_10552,N_11746);
nor U12854 (N_12854,N_10135,N_10737);
nor U12855 (N_12855,N_10419,N_11674);
and U12856 (N_12856,N_10958,N_11517);
nand U12857 (N_12857,N_10238,N_10441);
nor U12858 (N_12858,N_10036,N_10584);
or U12859 (N_12859,N_11205,N_11314);
or U12860 (N_12860,N_11806,N_10814);
xor U12861 (N_12861,N_11662,N_11089);
and U12862 (N_12862,N_10177,N_10893);
or U12863 (N_12863,N_10123,N_11611);
xor U12864 (N_12864,N_11164,N_11573);
nor U12865 (N_12865,N_10885,N_10753);
nand U12866 (N_12866,N_11459,N_10860);
nand U12867 (N_12867,N_10463,N_10535);
and U12868 (N_12868,N_10750,N_10014);
or U12869 (N_12869,N_11926,N_11187);
nor U12870 (N_12870,N_11088,N_10937);
nand U12871 (N_12871,N_11925,N_11257);
or U12872 (N_12872,N_10642,N_10662);
nor U12873 (N_12873,N_11535,N_11865);
nand U12874 (N_12874,N_11500,N_11022);
xor U12875 (N_12875,N_10215,N_10118);
xnor U12876 (N_12876,N_11779,N_10484);
and U12877 (N_12877,N_10315,N_11163);
and U12878 (N_12878,N_10646,N_10572);
nand U12879 (N_12879,N_10525,N_10991);
nor U12880 (N_12880,N_10688,N_11879);
and U12881 (N_12881,N_11216,N_10565);
nand U12882 (N_12882,N_10825,N_10251);
and U12883 (N_12883,N_11317,N_10909);
or U12884 (N_12884,N_10744,N_10329);
nor U12885 (N_12885,N_10214,N_11269);
or U12886 (N_12886,N_10526,N_11101);
or U12887 (N_12887,N_10203,N_10960);
and U12888 (N_12888,N_10603,N_10317);
nor U12889 (N_12889,N_11510,N_10769);
nor U12890 (N_12890,N_10071,N_10993);
nor U12891 (N_12891,N_11254,N_10060);
nor U12892 (N_12892,N_11222,N_10262);
and U12893 (N_12893,N_11800,N_11128);
nand U12894 (N_12894,N_11278,N_10876);
nor U12895 (N_12895,N_11572,N_11093);
and U12896 (N_12896,N_11502,N_10440);
or U12897 (N_12897,N_11114,N_11316);
or U12898 (N_12898,N_11131,N_11291);
nand U12899 (N_12899,N_11098,N_11122);
nor U12900 (N_12900,N_11390,N_10601);
nand U12901 (N_12901,N_11519,N_10789);
and U12902 (N_12902,N_10736,N_10127);
or U12903 (N_12903,N_11700,N_11031);
nand U12904 (N_12904,N_10580,N_11543);
and U12905 (N_12905,N_10822,N_11766);
and U12906 (N_12906,N_10079,N_10568);
and U12907 (N_12907,N_11703,N_10726);
nand U12908 (N_12908,N_11514,N_11110);
nor U12909 (N_12909,N_11977,N_10400);
or U12910 (N_12910,N_11807,N_11688);
and U12911 (N_12911,N_11524,N_10026);
and U12912 (N_12912,N_10390,N_11551);
xnor U12913 (N_12913,N_11315,N_10401);
xor U12914 (N_12914,N_10035,N_11349);
and U12915 (N_12915,N_11223,N_10332);
and U12916 (N_12916,N_11039,N_11447);
or U12917 (N_12917,N_10591,N_11425);
nand U12918 (N_12918,N_11608,N_11846);
nand U12919 (N_12919,N_10016,N_10875);
and U12920 (N_12920,N_10972,N_10450);
or U12921 (N_12921,N_10274,N_10059);
nand U12922 (N_12922,N_11715,N_11764);
and U12923 (N_12923,N_11281,N_10098);
xnor U12924 (N_12924,N_11555,N_10861);
nand U12925 (N_12925,N_11379,N_10683);
xnor U12926 (N_12926,N_11448,N_11373);
and U12927 (N_12927,N_11718,N_10775);
nand U12928 (N_12928,N_11518,N_10989);
nor U12929 (N_12929,N_11906,N_10521);
nand U12930 (N_12930,N_11938,N_10948);
or U12931 (N_12931,N_10656,N_11760);
and U12932 (N_12932,N_10220,N_10827);
nor U12933 (N_12933,N_11892,N_10064);
or U12934 (N_12934,N_10490,N_11389);
nand U12935 (N_12935,N_11247,N_11303);
xnor U12936 (N_12936,N_11747,N_11273);
nor U12937 (N_12937,N_11750,N_10447);
or U12938 (N_12938,N_10072,N_11932);
nor U12939 (N_12939,N_11469,N_10969);
nand U12940 (N_12940,N_10693,N_11346);
nand U12941 (N_12941,N_10456,N_11842);
and U12942 (N_12942,N_10610,N_11559);
and U12943 (N_12943,N_11821,N_10809);
nand U12944 (N_12944,N_10292,N_11597);
and U12945 (N_12945,N_10999,N_10362);
nand U12946 (N_12946,N_11714,N_10167);
or U12947 (N_12947,N_10846,N_11716);
nand U12948 (N_12948,N_11285,N_11056);
nand U12949 (N_12949,N_10593,N_11313);
or U12950 (N_12950,N_11481,N_11940);
and U12951 (N_12951,N_11845,N_10046);
nand U12952 (N_12952,N_10273,N_10094);
and U12953 (N_12953,N_10797,N_10295);
nor U12954 (N_12954,N_11882,N_11277);
and U12955 (N_12955,N_10331,N_10155);
nand U12956 (N_12956,N_10507,N_11198);
and U12957 (N_12957,N_10919,N_11337);
nand U12958 (N_12958,N_11670,N_10226);
xor U12959 (N_12959,N_10004,N_10828);
and U12960 (N_12960,N_11307,N_10540);
nor U12961 (N_12961,N_11177,N_11064);
or U12962 (N_12962,N_11378,N_11833);
xor U12963 (N_12963,N_11522,N_10303);
or U12964 (N_12964,N_10296,N_11831);
xnor U12965 (N_12965,N_10386,N_11876);
and U12966 (N_12966,N_11652,N_11839);
or U12967 (N_12967,N_11847,N_11549);
or U12968 (N_12968,N_10640,N_11686);
nor U12969 (N_12969,N_11207,N_10198);
or U12970 (N_12970,N_10446,N_10153);
or U12971 (N_12971,N_10844,N_11866);
nand U12972 (N_12972,N_10264,N_10323);
nand U12973 (N_12973,N_11722,N_10370);
nand U12974 (N_12974,N_10039,N_11452);
nand U12975 (N_12975,N_11144,N_11515);
nor U12976 (N_12976,N_10671,N_11019);
or U12977 (N_12977,N_11744,N_11657);
xnor U12978 (N_12978,N_10623,N_10964);
or U12979 (N_12979,N_11533,N_10018);
nor U12980 (N_12980,N_10148,N_10097);
nor U12981 (N_12981,N_10350,N_10592);
or U12982 (N_12982,N_10638,N_11618);
xor U12983 (N_12983,N_11080,N_11786);
nor U12984 (N_12984,N_10497,N_10613);
nor U12985 (N_12985,N_11030,N_11872);
nor U12986 (N_12986,N_11409,N_11363);
nand U12987 (N_12987,N_10470,N_11150);
or U12988 (N_12988,N_11133,N_11671);
xor U12989 (N_12989,N_10477,N_10648);
xor U12990 (N_12990,N_11461,N_11603);
nand U12991 (N_12991,N_10077,N_11583);
nor U12992 (N_12992,N_11928,N_10491);
or U12993 (N_12993,N_11723,N_10694);
and U12994 (N_12994,N_11375,N_10218);
or U12995 (N_12995,N_11259,N_11232);
or U12996 (N_12996,N_10073,N_11383);
nand U12997 (N_12997,N_11987,N_10594);
nand U12998 (N_12998,N_11710,N_10407);
xnor U12999 (N_12999,N_11589,N_11973);
nand U13000 (N_13000,N_11380,N_11906);
and U13001 (N_13001,N_11371,N_10019);
nand U13002 (N_13002,N_10696,N_11033);
nand U13003 (N_13003,N_10265,N_11202);
nand U13004 (N_13004,N_10781,N_11362);
xor U13005 (N_13005,N_11582,N_11713);
nand U13006 (N_13006,N_10021,N_10632);
nor U13007 (N_13007,N_11571,N_11419);
or U13008 (N_13008,N_10382,N_10502);
or U13009 (N_13009,N_11485,N_10060);
or U13010 (N_13010,N_11181,N_11764);
and U13011 (N_13011,N_11776,N_11102);
nor U13012 (N_13012,N_11579,N_10859);
or U13013 (N_13013,N_10192,N_11775);
and U13014 (N_13014,N_11720,N_11673);
nand U13015 (N_13015,N_11593,N_11433);
and U13016 (N_13016,N_11379,N_10621);
and U13017 (N_13017,N_11974,N_10786);
nor U13018 (N_13018,N_11453,N_10153);
or U13019 (N_13019,N_10204,N_11084);
or U13020 (N_13020,N_11608,N_10526);
nand U13021 (N_13021,N_10436,N_10493);
nor U13022 (N_13022,N_10519,N_10225);
or U13023 (N_13023,N_10039,N_11389);
or U13024 (N_13024,N_10031,N_11137);
nand U13025 (N_13025,N_10627,N_10121);
nor U13026 (N_13026,N_10439,N_11324);
nor U13027 (N_13027,N_11124,N_10595);
xor U13028 (N_13028,N_11578,N_10580);
xnor U13029 (N_13029,N_10856,N_10657);
or U13030 (N_13030,N_10229,N_10277);
xnor U13031 (N_13031,N_11974,N_10674);
or U13032 (N_13032,N_11999,N_11274);
nand U13033 (N_13033,N_10921,N_10072);
and U13034 (N_13034,N_10344,N_11487);
and U13035 (N_13035,N_10449,N_11346);
nor U13036 (N_13036,N_11226,N_11887);
and U13037 (N_13037,N_10738,N_10899);
or U13038 (N_13038,N_11427,N_10038);
or U13039 (N_13039,N_10395,N_11593);
nand U13040 (N_13040,N_10228,N_10315);
nand U13041 (N_13041,N_11139,N_11054);
or U13042 (N_13042,N_11652,N_10413);
nor U13043 (N_13043,N_11340,N_11443);
nor U13044 (N_13044,N_10322,N_10912);
and U13045 (N_13045,N_10737,N_11060);
and U13046 (N_13046,N_10501,N_10270);
nand U13047 (N_13047,N_10432,N_11029);
or U13048 (N_13048,N_11111,N_11228);
nand U13049 (N_13049,N_10614,N_10501);
nand U13050 (N_13050,N_11492,N_11125);
xnor U13051 (N_13051,N_10382,N_11820);
nand U13052 (N_13052,N_10216,N_10269);
nand U13053 (N_13053,N_10158,N_11870);
xnor U13054 (N_13054,N_10830,N_11478);
nor U13055 (N_13055,N_10053,N_10065);
nand U13056 (N_13056,N_10938,N_10032);
and U13057 (N_13057,N_10425,N_10582);
nor U13058 (N_13058,N_10328,N_11789);
nand U13059 (N_13059,N_10812,N_10123);
nor U13060 (N_13060,N_11399,N_11076);
nand U13061 (N_13061,N_11360,N_11972);
nor U13062 (N_13062,N_11926,N_10124);
and U13063 (N_13063,N_10948,N_11144);
or U13064 (N_13064,N_10928,N_11502);
nand U13065 (N_13065,N_10317,N_10798);
xnor U13066 (N_13066,N_10525,N_11999);
nand U13067 (N_13067,N_10629,N_11450);
and U13068 (N_13068,N_11668,N_10792);
and U13069 (N_13069,N_10083,N_11991);
nor U13070 (N_13070,N_10701,N_11440);
and U13071 (N_13071,N_11364,N_10916);
and U13072 (N_13072,N_10880,N_11002);
and U13073 (N_13073,N_10655,N_10621);
or U13074 (N_13074,N_10490,N_10398);
nor U13075 (N_13075,N_11488,N_11212);
nor U13076 (N_13076,N_10534,N_11699);
nand U13077 (N_13077,N_11917,N_11894);
and U13078 (N_13078,N_11902,N_10874);
nor U13079 (N_13079,N_10584,N_10364);
nor U13080 (N_13080,N_10831,N_11824);
nand U13081 (N_13081,N_11593,N_10150);
or U13082 (N_13082,N_11141,N_10887);
nor U13083 (N_13083,N_11409,N_10979);
or U13084 (N_13084,N_11875,N_11244);
nand U13085 (N_13085,N_11595,N_11611);
nor U13086 (N_13086,N_10233,N_11075);
xor U13087 (N_13087,N_10649,N_11838);
nand U13088 (N_13088,N_10472,N_11931);
or U13089 (N_13089,N_10242,N_11831);
nor U13090 (N_13090,N_11384,N_10076);
or U13091 (N_13091,N_10006,N_10289);
and U13092 (N_13092,N_11552,N_11850);
or U13093 (N_13093,N_10093,N_11427);
or U13094 (N_13094,N_11103,N_10601);
and U13095 (N_13095,N_10666,N_11004);
nand U13096 (N_13096,N_11658,N_10756);
nand U13097 (N_13097,N_10325,N_11646);
and U13098 (N_13098,N_11935,N_11450);
or U13099 (N_13099,N_11066,N_10656);
nor U13100 (N_13100,N_10029,N_11854);
and U13101 (N_13101,N_11435,N_11287);
or U13102 (N_13102,N_11195,N_11072);
xnor U13103 (N_13103,N_11420,N_11581);
or U13104 (N_13104,N_10632,N_10038);
xnor U13105 (N_13105,N_10689,N_11148);
or U13106 (N_13106,N_10406,N_11003);
and U13107 (N_13107,N_10034,N_10891);
nand U13108 (N_13108,N_10755,N_11163);
nand U13109 (N_13109,N_11284,N_11034);
nand U13110 (N_13110,N_11729,N_11457);
nand U13111 (N_13111,N_11824,N_10996);
or U13112 (N_13112,N_10254,N_11443);
nor U13113 (N_13113,N_10974,N_10544);
nor U13114 (N_13114,N_10171,N_11441);
nand U13115 (N_13115,N_10428,N_11221);
nand U13116 (N_13116,N_10393,N_10286);
nor U13117 (N_13117,N_11810,N_11245);
and U13118 (N_13118,N_10879,N_10799);
nor U13119 (N_13119,N_10487,N_11200);
nand U13120 (N_13120,N_10787,N_10934);
and U13121 (N_13121,N_11065,N_11743);
nand U13122 (N_13122,N_11599,N_11758);
nor U13123 (N_13123,N_10753,N_11082);
or U13124 (N_13124,N_11010,N_10986);
nand U13125 (N_13125,N_10299,N_11854);
xor U13126 (N_13126,N_10009,N_10414);
xnor U13127 (N_13127,N_11852,N_10395);
xnor U13128 (N_13128,N_10622,N_10454);
and U13129 (N_13129,N_10725,N_10651);
or U13130 (N_13130,N_11311,N_11143);
and U13131 (N_13131,N_11182,N_10101);
nand U13132 (N_13132,N_10594,N_11557);
nor U13133 (N_13133,N_10487,N_11935);
xor U13134 (N_13134,N_11189,N_11206);
nor U13135 (N_13135,N_11093,N_10278);
nand U13136 (N_13136,N_10138,N_10342);
nand U13137 (N_13137,N_10717,N_11093);
nand U13138 (N_13138,N_11719,N_10033);
and U13139 (N_13139,N_10697,N_10552);
or U13140 (N_13140,N_10864,N_11905);
nand U13141 (N_13141,N_11723,N_10169);
nand U13142 (N_13142,N_11952,N_11742);
and U13143 (N_13143,N_11954,N_11991);
and U13144 (N_13144,N_11195,N_10649);
or U13145 (N_13145,N_10877,N_11596);
nand U13146 (N_13146,N_10778,N_10998);
nand U13147 (N_13147,N_11212,N_11470);
nand U13148 (N_13148,N_10156,N_11415);
or U13149 (N_13149,N_11484,N_10726);
nor U13150 (N_13150,N_10581,N_10564);
and U13151 (N_13151,N_10164,N_10111);
or U13152 (N_13152,N_10731,N_10311);
and U13153 (N_13153,N_10875,N_10812);
and U13154 (N_13154,N_11210,N_10060);
or U13155 (N_13155,N_11159,N_11408);
and U13156 (N_13156,N_10975,N_11398);
and U13157 (N_13157,N_11145,N_10210);
or U13158 (N_13158,N_11985,N_10697);
nand U13159 (N_13159,N_11150,N_11160);
nor U13160 (N_13160,N_10969,N_10186);
nand U13161 (N_13161,N_11597,N_11493);
xnor U13162 (N_13162,N_10822,N_10777);
xor U13163 (N_13163,N_11205,N_11873);
or U13164 (N_13164,N_11914,N_10631);
nor U13165 (N_13165,N_10037,N_10996);
or U13166 (N_13166,N_10580,N_11390);
nand U13167 (N_13167,N_11120,N_10593);
nand U13168 (N_13168,N_10318,N_11137);
nor U13169 (N_13169,N_11559,N_11636);
nor U13170 (N_13170,N_10200,N_11000);
nand U13171 (N_13171,N_11163,N_11557);
or U13172 (N_13172,N_11562,N_10334);
and U13173 (N_13173,N_11584,N_11482);
nor U13174 (N_13174,N_10999,N_11328);
or U13175 (N_13175,N_10551,N_10395);
or U13176 (N_13176,N_11595,N_11144);
nand U13177 (N_13177,N_10531,N_10639);
or U13178 (N_13178,N_11412,N_10037);
nor U13179 (N_13179,N_11382,N_10223);
nand U13180 (N_13180,N_10121,N_11486);
and U13181 (N_13181,N_11285,N_10831);
nor U13182 (N_13182,N_10130,N_11622);
nand U13183 (N_13183,N_11568,N_11348);
and U13184 (N_13184,N_11779,N_10498);
or U13185 (N_13185,N_10206,N_10564);
or U13186 (N_13186,N_10544,N_11120);
nand U13187 (N_13187,N_10134,N_10347);
nor U13188 (N_13188,N_10024,N_10650);
nor U13189 (N_13189,N_10911,N_11466);
nand U13190 (N_13190,N_10920,N_11379);
or U13191 (N_13191,N_11740,N_10213);
nand U13192 (N_13192,N_11777,N_10942);
nor U13193 (N_13193,N_11051,N_10663);
or U13194 (N_13194,N_11183,N_11464);
nand U13195 (N_13195,N_11383,N_11054);
nor U13196 (N_13196,N_10844,N_11735);
nand U13197 (N_13197,N_10518,N_11416);
and U13198 (N_13198,N_11129,N_11323);
and U13199 (N_13199,N_10419,N_11265);
nor U13200 (N_13200,N_10486,N_11398);
or U13201 (N_13201,N_11854,N_10649);
and U13202 (N_13202,N_11757,N_10087);
and U13203 (N_13203,N_10303,N_10637);
or U13204 (N_13204,N_10474,N_11470);
nand U13205 (N_13205,N_11303,N_10944);
nand U13206 (N_13206,N_10440,N_10470);
or U13207 (N_13207,N_11265,N_11019);
nand U13208 (N_13208,N_11888,N_10627);
or U13209 (N_13209,N_11592,N_11289);
nand U13210 (N_13210,N_11703,N_10760);
nor U13211 (N_13211,N_10048,N_11214);
nor U13212 (N_13212,N_10129,N_10034);
nand U13213 (N_13213,N_11292,N_11035);
nand U13214 (N_13214,N_10213,N_11906);
nor U13215 (N_13215,N_10173,N_11633);
and U13216 (N_13216,N_10712,N_11553);
or U13217 (N_13217,N_11873,N_11414);
xnor U13218 (N_13218,N_11353,N_11975);
nand U13219 (N_13219,N_10935,N_10319);
nor U13220 (N_13220,N_11603,N_10337);
or U13221 (N_13221,N_10732,N_10027);
xnor U13222 (N_13222,N_10003,N_10679);
or U13223 (N_13223,N_10800,N_10716);
and U13224 (N_13224,N_11827,N_10745);
and U13225 (N_13225,N_10425,N_11495);
nor U13226 (N_13226,N_11707,N_11679);
nand U13227 (N_13227,N_10353,N_11353);
xor U13228 (N_13228,N_11112,N_11960);
nor U13229 (N_13229,N_10676,N_10394);
or U13230 (N_13230,N_11802,N_11034);
nor U13231 (N_13231,N_10853,N_11494);
xnor U13232 (N_13232,N_10952,N_10575);
nor U13233 (N_13233,N_10639,N_10448);
nand U13234 (N_13234,N_10607,N_10597);
or U13235 (N_13235,N_10915,N_11754);
nand U13236 (N_13236,N_11066,N_11340);
and U13237 (N_13237,N_10456,N_10978);
and U13238 (N_13238,N_10481,N_10449);
and U13239 (N_13239,N_11117,N_11215);
and U13240 (N_13240,N_11318,N_11894);
nor U13241 (N_13241,N_11049,N_11824);
nor U13242 (N_13242,N_10466,N_11348);
nor U13243 (N_13243,N_10734,N_11658);
or U13244 (N_13244,N_11760,N_11335);
or U13245 (N_13245,N_11063,N_10134);
nor U13246 (N_13246,N_10393,N_11930);
and U13247 (N_13247,N_10937,N_10603);
nor U13248 (N_13248,N_10294,N_11896);
nand U13249 (N_13249,N_11101,N_10797);
or U13250 (N_13250,N_10277,N_11555);
and U13251 (N_13251,N_11833,N_11484);
or U13252 (N_13252,N_11258,N_11375);
nor U13253 (N_13253,N_10772,N_10045);
nand U13254 (N_13254,N_10651,N_10917);
and U13255 (N_13255,N_10688,N_11233);
or U13256 (N_13256,N_11357,N_11726);
nor U13257 (N_13257,N_11494,N_11071);
nor U13258 (N_13258,N_10064,N_11593);
nor U13259 (N_13259,N_11789,N_10821);
or U13260 (N_13260,N_10269,N_11065);
or U13261 (N_13261,N_11697,N_10030);
nand U13262 (N_13262,N_11714,N_10899);
nor U13263 (N_13263,N_10335,N_11057);
xor U13264 (N_13264,N_10050,N_10288);
xnor U13265 (N_13265,N_11488,N_10195);
nor U13266 (N_13266,N_11784,N_10302);
xor U13267 (N_13267,N_11984,N_11928);
and U13268 (N_13268,N_11996,N_10832);
nor U13269 (N_13269,N_10030,N_10055);
nand U13270 (N_13270,N_10567,N_11998);
nand U13271 (N_13271,N_11418,N_10372);
nor U13272 (N_13272,N_10372,N_10716);
nand U13273 (N_13273,N_11696,N_11948);
or U13274 (N_13274,N_11750,N_10161);
or U13275 (N_13275,N_11003,N_10662);
and U13276 (N_13276,N_10195,N_10604);
nor U13277 (N_13277,N_10319,N_10734);
xor U13278 (N_13278,N_10825,N_11520);
and U13279 (N_13279,N_10319,N_11314);
nand U13280 (N_13280,N_10781,N_11182);
nor U13281 (N_13281,N_11252,N_11394);
nand U13282 (N_13282,N_11764,N_10685);
or U13283 (N_13283,N_11634,N_10053);
and U13284 (N_13284,N_10068,N_11781);
nor U13285 (N_13285,N_10550,N_11784);
nor U13286 (N_13286,N_10523,N_11174);
and U13287 (N_13287,N_10181,N_11386);
and U13288 (N_13288,N_11851,N_11249);
or U13289 (N_13289,N_10433,N_10101);
or U13290 (N_13290,N_10226,N_11818);
nand U13291 (N_13291,N_10741,N_11516);
nor U13292 (N_13292,N_10316,N_10924);
nand U13293 (N_13293,N_10363,N_11261);
and U13294 (N_13294,N_11307,N_10717);
nor U13295 (N_13295,N_11184,N_11361);
and U13296 (N_13296,N_11478,N_11740);
nand U13297 (N_13297,N_10828,N_11254);
or U13298 (N_13298,N_11943,N_11278);
nand U13299 (N_13299,N_10503,N_11582);
or U13300 (N_13300,N_10987,N_10991);
and U13301 (N_13301,N_10712,N_11707);
nor U13302 (N_13302,N_10373,N_11356);
or U13303 (N_13303,N_11637,N_10602);
and U13304 (N_13304,N_10637,N_11606);
nand U13305 (N_13305,N_11172,N_11166);
nor U13306 (N_13306,N_11677,N_11691);
nor U13307 (N_13307,N_11330,N_11236);
or U13308 (N_13308,N_10316,N_11814);
and U13309 (N_13309,N_10815,N_10169);
nand U13310 (N_13310,N_10937,N_11949);
nor U13311 (N_13311,N_10540,N_10058);
and U13312 (N_13312,N_10965,N_11705);
nor U13313 (N_13313,N_11803,N_11095);
nor U13314 (N_13314,N_10766,N_10080);
or U13315 (N_13315,N_11232,N_10954);
or U13316 (N_13316,N_10310,N_10834);
and U13317 (N_13317,N_10465,N_11943);
and U13318 (N_13318,N_10539,N_10729);
and U13319 (N_13319,N_11716,N_11732);
nor U13320 (N_13320,N_10130,N_11007);
nand U13321 (N_13321,N_10827,N_10501);
and U13322 (N_13322,N_11910,N_11246);
nand U13323 (N_13323,N_10449,N_11298);
nor U13324 (N_13324,N_11812,N_10479);
or U13325 (N_13325,N_11244,N_10406);
or U13326 (N_13326,N_10093,N_11476);
xor U13327 (N_13327,N_10050,N_10721);
nor U13328 (N_13328,N_10603,N_11903);
xnor U13329 (N_13329,N_11247,N_11651);
or U13330 (N_13330,N_10731,N_11181);
nor U13331 (N_13331,N_10236,N_11176);
and U13332 (N_13332,N_11850,N_10705);
xor U13333 (N_13333,N_11926,N_11027);
xor U13334 (N_13334,N_10502,N_10760);
nand U13335 (N_13335,N_11058,N_10732);
nor U13336 (N_13336,N_11960,N_11943);
nand U13337 (N_13337,N_11285,N_10920);
nor U13338 (N_13338,N_11690,N_11664);
and U13339 (N_13339,N_11698,N_11218);
nor U13340 (N_13340,N_11009,N_11246);
and U13341 (N_13341,N_11919,N_10996);
nand U13342 (N_13342,N_10266,N_10803);
nand U13343 (N_13343,N_11786,N_10636);
and U13344 (N_13344,N_10527,N_11029);
nor U13345 (N_13345,N_11494,N_10633);
nor U13346 (N_13346,N_10332,N_11489);
xor U13347 (N_13347,N_10025,N_11409);
or U13348 (N_13348,N_10307,N_11154);
nor U13349 (N_13349,N_11758,N_11483);
and U13350 (N_13350,N_11932,N_11627);
nor U13351 (N_13351,N_10896,N_11561);
nand U13352 (N_13352,N_11302,N_10343);
nand U13353 (N_13353,N_11811,N_11329);
or U13354 (N_13354,N_10288,N_11057);
nand U13355 (N_13355,N_10480,N_10453);
nor U13356 (N_13356,N_11106,N_11752);
or U13357 (N_13357,N_11847,N_11554);
nand U13358 (N_13358,N_10397,N_11865);
and U13359 (N_13359,N_11850,N_10572);
or U13360 (N_13360,N_10546,N_10597);
and U13361 (N_13361,N_10709,N_10684);
nor U13362 (N_13362,N_10132,N_10826);
nand U13363 (N_13363,N_10619,N_11503);
xor U13364 (N_13364,N_11607,N_10750);
and U13365 (N_13365,N_10817,N_11051);
or U13366 (N_13366,N_10749,N_11684);
nor U13367 (N_13367,N_10828,N_11354);
or U13368 (N_13368,N_10836,N_11738);
nor U13369 (N_13369,N_11961,N_11441);
nor U13370 (N_13370,N_11138,N_11427);
or U13371 (N_13371,N_10647,N_11589);
nand U13372 (N_13372,N_10501,N_10909);
or U13373 (N_13373,N_11510,N_11300);
and U13374 (N_13374,N_11161,N_11079);
nor U13375 (N_13375,N_10351,N_11920);
and U13376 (N_13376,N_10455,N_10794);
xor U13377 (N_13377,N_11132,N_11075);
or U13378 (N_13378,N_10159,N_10509);
nand U13379 (N_13379,N_10085,N_10599);
nor U13380 (N_13380,N_10282,N_10608);
nor U13381 (N_13381,N_10197,N_11258);
or U13382 (N_13382,N_10349,N_10258);
and U13383 (N_13383,N_10105,N_10223);
xnor U13384 (N_13384,N_11934,N_10236);
nand U13385 (N_13385,N_11835,N_10361);
or U13386 (N_13386,N_11948,N_10704);
and U13387 (N_13387,N_11945,N_10879);
or U13388 (N_13388,N_10184,N_10687);
xor U13389 (N_13389,N_11028,N_11757);
or U13390 (N_13390,N_11777,N_10316);
or U13391 (N_13391,N_10477,N_11254);
or U13392 (N_13392,N_11758,N_10552);
and U13393 (N_13393,N_10116,N_11272);
and U13394 (N_13394,N_11431,N_11417);
and U13395 (N_13395,N_11679,N_11829);
nor U13396 (N_13396,N_10360,N_11373);
nand U13397 (N_13397,N_11429,N_11520);
xor U13398 (N_13398,N_11554,N_10446);
or U13399 (N_13399,N_11070,N_11037);
and U13400 (N_13400,N_11850,N_11179);
or U13401 (N_13401,N_11864,N_11027);
nor U13402 (N_13402,N_11685,N_11132);
and U13403 (N_13403,N_10817,N_11083);
and U13404 (N_13404,N_10371,N_10386);
and U13405 (N_13405,N_11801,N_10175);
nor U13406 (N_13406,N_10166,N_10479);
or U13407 (N_13407,N_10550,N_11000);
nand U13408 (N_13408,N_10468,N_10779);
or U13409 (N_13409,N_10479,N_10833);
or U13410 (N_13410,N_11545,N_11709);
or U13411 (N_13411,N_11858,N_10976);
nor U13412 (N_13412,N_11260,N_10083);
and U13413 (N_13413,N_11763,N_10655);
nand U13414 (N_13414,N_10497,N_11183);
and U13415 (N_13415,N_10051,N_11135);
and U13416 (N_13416,N_11328,N_10035);
nand U13417 (N_13417,N_11861,N_10660);
xnor U13418 (N_13418,N_11517,N_10785);
xnor U13419 (N_13419,N_10345,N_10712);
xor U13420 (N_13420,N_11992,N_11821);
or U13421 (N_13421,N_11225,N_10734);
nand U13422 (N_13422,N_10967,N_11848);
nor U13423 (N_13423,N_11857,N_10166);
and U13424 (N_13424,N_10367,N_11982);
nor U13425 (N_13425,N_11681,N_10097);
nor U13426 (N_13426,N_11250,N_10125);
and U13427 (N_13427,N_10717,N_10604);
or U13428 (N_13428,N_11626,N_11592);
nor U13429 (N_13429,N_10725,N_10010);
nand U13430 (N_13430,N_11207,N_11116);
nand U13431 (N_13431,N_10995,N_10668);
xor U13432 (N_13432,N_11027,N_11852);
nor U13433 (N_13433,N_11395,N_11096);
and U13434 (N_13434,N_10519,N_11768);
nor U13435 (N_13435,N_11368,N_10782);
or U13436 (N_13436,N_11579,N_10019);
or U13437 (N_13437,N_10037,N_10294);
or U13438 (N_13438,N_11508,N_10875);
nand U13439 (N_13439,N_11395,N_11563);
and U13440 (N_13440,N_10848,N_11343);
and U13441 (N_13441,N_11805,N_10574);
nor U13442 (N_13442,N_11972,N_10290);
xor U13443 (N_13443,N_11023,N_10848);
and U13444 (N_13444,N_11305,N_11429);
nor U13445 (N_13445,N_10467,N_10277);
and U13446 (N_13446,N_10027,N_10548);
or U13447 (N_13447,N_10469,N_11065);
nand U13448 (N_13448,N_11611,N_11835);
and U13449 (N_13449,N_11271,N_10281);
nand U13450 (N_13450,N_10048,N_11523);
nor U13451 (N_13451,N_10699,N_11275);
and U13452 (N_13452,N_10571,N_11590);
and U13453 (N_13453,N_11303,N_11084);
and U13454 (N_13454,N_10035,N_10875);
and U13455 (N_13455,N_11278,N_10470);
or U13456 (N_13456,N_11121,N_11927);
or U13457 (N_13457,N_11430,N_11263);
and U13458 (N_13458,N_10874,N_10794);
nor U13459 (N_13459,N_10646,N_10900);
nand U13460 (N_13460,N_10797,N_10355);
and U13461 (N_13461,N_11976,N_11196);
and U13462 (N_13462,N_10519,N_11584);
xnor U13463 (N_13463,N_10419,N_11667);
or U13464 (N_13464,N_10661,N_10166);
nor U13465 (N_13465,N_11853,N_10449);
or U13466 (N_13466,N_10489,N_10648);
or U13467 (N_13467,N_11407,N_11223);
and U13468 (N_13468,N_10465,N_11681);
and U13469 (N_13469,N_10220,N_11247);
xor U13470 (N_13470,N_11058,N_10960);
nor U13471 (N_13471,N_10602,N_11073);
and U13472 (N_13472,N_10267,N_11517);
nand U13473 (N_13473,N_10545,N_11750);
or U13474 (N_13474,N_11818,N_11479);
and U13475 (N_13475,N_11776,N_11648);
nand U13476 (N_13476,N_11591,N_10092);
nor U13477 (N_13477,N_11736,N_10433);
or U13478 (N_13478,N_11264,N_11937);
nor U13479 (N_13479,N_11454,N_11206);
xor U13480 (N_13480,N_11083,N_10512);
or U13481 (N_13481,N_11076,N_11780);
or U13482 (N_13482,N_10726,N_11922);
nor U13483 (N_13483,N_10554,N_10836);
or U13484 (N_13484,N_10894,N_10726);
and U13485 (N_13485,N_11517,N_11379);
nand U13486 (N_13486,N_10959,N_10709);
or U13487 (N_13487,N_11613,N_11394);
nor U13488 (N_13488,N_10243,N_11065);
or U13489 (N_13489,N_10538,N_11200);
nor U13490 (N_13490,N_11698,N_10881);
nor U13491 (N_13491,N_11706,N_11177);
and U13492 (N_13492,N_11270,N_10099);
nand U13493 (N_13493,N_10310,N_10167);
and U13494 (N_13494,N_10601,N_10974);
nand U13495 (N_13495,N_10331,N_11053);
nand U13496 (N_13496,N_10204,N_11290);
or U13497 (N_13497,N_11273,N_10734);
and U13498 (N_13498,N_10291,N_10363);
and U13499 (N_13499,N_11183,N_10919);
nand U13500 (N_13500,N_10954,N_11235);
and U13501 (N_13501,N_10545,N_11723);
or U13502 (N_13502,N_11645,N_10937);
or U13503 (N_13503,N_11212,N_10632);
and U13504 (N_13504,N_10194,N_11693);
nor U13505 (N_13505,N_10972,N_11048);
or U13506 (N_13506,N_11767,N_10074);
xor U13507 (N_13507,N_11355,N_11948);
and U13508 (N_13508,N_10310,N_10741);
or U13509 (N_13509,N_11117,N_11111);
nor U13510 (N_13510,N_11693,N_10888);
nor U13511 (N_13511,N_11368,N_11035);
or U13512 (N_13512,N_11760,N_10679);
nand U13513 (N_13513,N_10918,N_10219);
and U13514 (N_13514,N_11201,N_10268);
and U13515 (N_13515,N_11578,N_10834);
or U13516 (N_13516,N_10531,N_11729);
and U13517 (N_13517,N_11816,N_10877);
xnor U13518 (N_13518,N_11043,N_10149);
nand U13519 (N_13519,N_11403,N_10232);
xor U13520 (N_13520,N_10107,N_10132);
and U13521 (N_13521,N_11698,N_11476);
and U13522 (N_13522,N_11173,N_10639);
nand U13523 (N_13523,N_11921,N_10038);
nor U13524 (N_13524,N_10186,N_11920);
nand U13525 (N_13525,N_11160,N_11460);
or U13526 (N_13526,N_10628,N_10474);
or U13527 (N_13527,N_11247,N_10727);
nor U13528 (N_13528,N_10873,N_10906);
nor U13529 (N_13529,N_10294,N_10219);
xor U13530 (N_13530,N_11124,N_11910);
or U13531 (N_13531,N_11808,N_11816);
nor U13532 (N_13532,N_10456,N_10730);
nor U13533 (N_13533,N_11474,N_10270);
nand U13534 (N_13534,N_10831,N_10012);
and U13535 (N_13535,N_11621,N_10421);
and U13536 (N_13536,N_10703,N_10220);
nor U13537 (N_13537,N_10665,N_11682);
nor U13538 (N_13538,N_11032,N_10280);
and U13539 (N_13539,N_11725,N_11343);
nor U13540 (N_13540,N_11782,N_11780);
nor U13541 (N_13541,N_11152,N_10151);
xor U13542 (N_13542,N_11837,N_10889);
nor U13543 (N_13543,N_10018,N_11936);
xor U13544 (N_13544,N_11626,N_10983);
nand U13545 (N_13545,N_10607,N_10184);
xor U13546 (N_13546,N_11213,N_11684);
or U13547 (N_13547,N_10883,N_11371);
nand U13548 (N_13548,N_11887,N_10967);
or U13549 (N_13549,N_11583,N_10914);
or U13550 (N_13550,N_10828,N_10601);
xor U13551 (N_13551,N_11470,N_10205);
xor U13552 (N_13552,N_11314,N_10553);
nand U13553 (N_13553,N_10560,N_10290);
or U13554 (N_13554,N_10280,N_10952);
xor U13555 (N_13555,N_11846,N_11578);
nor U13556 (N_13556,N_11250,N_10709);
and U13557 (N_13557,N_11299,N_11228);
nor U13558 (N_13558,N_10105,N_10828);
nor U13559 (N_13559,N_11933,N_10424);
nor U13560 (N_13560,N_11112,N_10655);
or U13561 (N_13561,N_11696,N_10730);
xor U13562 (N_13562,N_10750,N_11778);
nor U13563 (N_13563,N_10994,N_10096);
nand U13564 (N_13564,N_11743,N_10795);
or U13565 (N_13565,N_10391,N_10560);
nand U13566 (N_13566,N_10911,N_11528);
and U13567 (N_13567,N_11288,N_10341);
and U13568 (N_13568,N_11241,N_11994);
and U13569 (N_13569,N_11224,N_11971);
or U13570 (N_13570,N_10101,N_11963);
or U13571 (N_13571,N_11287,N_11447);
and U13572 (N_13572,N_11532,N_10293);
nor U13573 (N_13573,N_10916,N_10716);
and U13574 (N_13574,N_11104,N_10197);
or U13575 (N_13575,N_11508,N_10567);
nand U13576 (N_13576,N_11941,N_10930);
or U13577 (N_13577,N_10092,N_10542);
nand U13578 (N_13578,N_11603,N_10166);
nor U13579 (N_13579,N_11149,N_11393);
and U13580 (N_13580,N_11662,N_10071);
or U13581 (N_13581,N_10732,N_11165);
nand U13582 (N_13582,N_11570,N_11950);
xor U13583 (N_13583,N_11399,N_10277);
nor U13584 (N_13584,N_10946,N_10358);
nand U13585 (N_13585,N_10408,N_10014);
nor U13586 (N_13586,N_10099,N_10055);
nand U13587 (N_13587,N_11649,N_11444);
nor U13588 (N_13588,N_11273,N_10990);
nor U13589 (N_13589,N_11034,N_11977);
nand U13590 (N_13590,N_10673,N_11297);
or U13591 (N_13591,N_10817,N_11111);
xor U13592 (N_13592,N_11808,N_10872);
or U13593 (N_13593,N_10125,N_11758);
nand U13594 (N_13594,N_10116,N_10803);
nand U13595 (N_13595,N_10345,N_10486);
or U13596 (N_13596,N_11823,N_10852);
nand U13597 (N_13597,N_10388,N_10810);
or U13598 (N_13598,N_11495,N_11940);
nor U13599 (N_13599,N_11972,N_11168);
and U13600 (N_13600,N_10280,N_10855);
and U13601 (N_13601,N_10584,N_11940);
and U13602 (N_13602,N_10487,N_11045);
nor U13603 (N_13603,N_11703,N_11201);
and U13604 (N_13604,N_10202,N_10961);
and U13605 (N_13605,N_10849,N_10175);
or U13606 (N_13606,N_11634,N_11576);
nor U13607 (N_13607,N_11198,N_10804);
and U13608 (N_13608,N_10047,N_11628);
or U13609 (N_13609,N_11712,N_10928);
nand U13610 (N_13610,N_10944,N_11698);
and U13611 (N_13611,N_10093,N_11196);
nor U13612 (N_13612,N_10678,N_11195);
nand U13613 (N_13613,N_11072,N_10370);
nand U13614 (N_13614,N_10183,N_11222);
or U13615 (N_13615,N_10164,N_11406);
xor U13616 (N_13616,N_10961,N_10772);
xor U13617 (N_13617,N_11901,N_11729);
and U13618 (N_13618,N_10420,N_10249);
and U13619 (N_13619,N_10308,N_10588);
nand U13620 (N_13620,N_10041,N_11446);
nor U13621 (N_13621,N_11989,N_10660);
nand U13622 (N_13622,N_11635,N_10603);
nor U13623 (N_13623,N_11243,N_11070);
and U13624 (N_13624,N_10705,N_11083);
nor U13625 (N_13625,N_10635,N_10392);
nor U13626 (N_13626,N_11002,N_11109);
or U13627 (N_13627,N_11202,N_11864);
and U13628 (N_13628,N_11069,N_11159);
nand U13629 (N_13629,N_10741,N_11890);
nor U13630 (N_13630,N_10257,N_11592);
nand U13631 (N_13631,N_10810,N_10597);
nor U13632 (N_13632,N_11125,N_10461);
nand U13633 (N_13633,N_11602,N_10847);
and U13634 (N_13634,N_10264,N_10019);
xnor U13635 (N_13635,N_11971,N_10419);
and U13636 (N_13636,N_11492,N_10316);
nor U13637 (N_13637,N_10897,N_11009);
and U13638 (N_13638,N_10671,N_11010);
nor U13639 (N_13639,N_11464,N_11249);
and U13640 (N_13640,N_10917,N_10918);
nor U13641 (N_13641,N_11023,N_10030);
and U13642 (N_13642,N_10588,N_11640);
nand U13643 (N_13643,N_11266,N_10983);
nor U13644 (N_13644,N_11058,N_10104);
nand U13645 (N_13645,N_11374,N_11139);
nor U13646 (N_13646,N_11461,N_10155);
nand U13647 (N_13647,N_11649,N_11241);
or U13648 (N_13648,N_10682,N_10220);
and U13649 (N_13649,N_10127,N_11968);
and U13650 (N_13650,N_10888,N_11973);
nand U13651 (N_13651,N_11543,N_10180);
or U13652 (N_13652,N_11000,N_11639);
nand U13653 (N_13653,N_10123,N_10226);
and U13654 (N_13654,N_11330,N_10933);
nand U13655 (N_13655,N_11174,N_11724);
and U13656 (N_13656,N_11328,N_11382);
nand U13657 (N_13657,N_11882,N_11808);
nor U13658 (N_13658,N_11912,N_10260);
or U13659 (N_13659,N_11270,N_10332);
nor U13660 (N_13660,N_10334,N_10474);
or U13661 (N_13661,N_10859,N_10127);
xnor U13662 (N_13662,N_11050,N_11900);
or U13663 (N_13663,N_10385,N_10838);
nand U13664 (N_13664,N_10131,N_10758);
or U13665 (N_13665,N_11083,N_10531);
xnor U13666 (N_13666,N_11110,N_10548);
or U13667 (N_13667,N_11136,N_10696);
nand U13668 (N_13668,N_10817,N_11237);
and U13669 (N_13669,N_10069,N_11851);
nand U13670 (N_13670,N_10288,N_11637);
nor U13671 (N_13671,N_11429,N_11899);
xnor U13672 (N_13672,N_10693,N_10171);
and U13673 (N_13673,N_10194,N_10522);
nand U13674 (N_13674,N_10889,N_11691);
nand U13675 (N_13675,N_10893,N_11464);
xnor U13676 (N_13676,N_10637,N_11518);
nand U13677 (N_13677,N_10495,N_11352);
or U13678 (N_13678,N_11374,N_11780);
and U13679 (N_13679,N_10640,N_11286);
nor U13680 (N_13680,N_10791,N_11552);
or U13681 (N_13681,N_10349,N_10218);
nand U13682 (N_13682,N_10813,N_11029);
nand U13683 (N_13683,N_10442,N_11669);
or U13684 (N_13684,N_10316,N_11369);
or U13685 (N_13685,N_11728,N_10831);
nor U13686 (N_13686,N_10192,N_10646);
xor U13687 (N_13687,N_11287,N_11387);
nor U13688 (N_13688,N_11794,N_11930);
xnor U13689 (N_13689,N_11610,N_10562);
or U13690 (N_13690,N_11357,N_10653);
nor U13691 (N_13691,N_10131,N_10568);
nand U13692 (N_13692,N_10716,N_10605);
or U13693 (N_13693,N_11070,N_10107);
nor U13694 (N_13694,N_10945,N_11099);
nor U13695 (N_13695,N_10581,N_11758);
nand U13696 (N_13696,N_11927,N_11408);
nor U13697 (N_13697,N_11928,N_10194);
or U13698 (N_13698,N_10655,N_10282);
nand U13699 (N_13699,N_11129,N_10499);
nor U13700 (N_13700,N_10821,N_10996);
nor U13701 (N_13701,N_10287,N_10471);
and U13702 (N_13702,N_11463,N_10782);
or U13703 (N_13703,N_10004,N_11346);
or U13704 (N_13704,N_10675,N_11924);
and U13705 (N_13705,N_11477,N_11439);
xor U13706 (N_13706,N_10274,N_10652);
and U13707 (N_13707,N_11265,N_10181);
nand U13708 (N_13708,N_10053,N_11473);
and U13709 (N_13709,N_10836,N_10585);
and U13710 (N_13710,N_10503,N_10255);
nor U13711 (N_13711,N_11690,N_10547);
nor U13712 (N_13712,N_11325,N_10007);
nor U13713 (N_13713,N_11042,N_10181);
or U13714 (N_13714,N_10519,N_10638);
nand U13715 (N_13715,N_10501,N_11325);
and U13716 (N_13716,N_10720,N_11926);
or U13717 (N_13717,N_11351,N_10287);
or U13718 (N_13718,N_10246,N_11981);
and U13719 (N_13719,N_11515,N_11542);
and U13720 (N_13720,N_10793,N_11822);
nor U13721 (N_13721,N_11630,N_11327);
nand U13722 (N_13722,N_10835,N_10939);
or U13723 (N_13723,N_10048,N_11288);
nor U13724 (N_13724,N_10685,N_11440);
nor U13725 (N_13725,N_11231,N_11460);
nand U13726 (N_13726,N_11129,N_10363);
nand U13727 (N_13727,N_10076,N_11910);
or U13728 (N_13728,N_10685,N_10275);
xnor U13729 (N_13729,N_10653,N_11481);
nor U13730 (N_13730,N_10715,N_11137);
and U13731 (N_13731,N_10968,N_10304);
nand U13732 (N_13732,N_10602,N_11915);
or U13733 (N_13733,N_10014,N_11900);
nand U13734 (N_13734,N_11318,N_11707);
nor U13735 (N_13735,N_11097,N_11570);
nand U13736 (N_13736,N_11290,N_10633);
or U13737 (N_13737,N_11831,N_11746);
nand U13738 (N_13738,N_10302,N_11568);
nand U13739 (N_13739,N_10480,N_11832);
nor U13740 (N_13740,N_10426,N_11139);
nand U13741 (N_13741,N_10966,N_11125);
xor U13742 (N_13742,N_11789,N_10238);
nor U13743 (N_13743,N_11013,N_10777);
nor U13744 (N_13744,N_11071,N_10677);
nand U13745 (N_13745,N_11163,N_10037);
nor U13746 (N_13746,N_10256,N_11745);
and U13747 (N_13747,N_10400,N_11566);
or U13748 (N_13748,N_10472,N_11197);
or U13749 (N_13749,N_10503,N_11157);
and U13750 (N_13750,N_10239,N_11310);
nand U13751 (N_13751,N_11324,N_10199);
and U13752 (N_13752,N_10821,N_10072);
or U13753 (N_13753,N_11920,N_10438);
and U13754 (N_13754,N_10655,N_10619);
nand U13755 (N_13755,N_11985,N_10926);
and U13756 (N_13756,N_11068,N_11316);
or U13757 (N_13757,N_10087,N_10277);
xnor U13758 (N_13758,N_10073,N_11481);
and U13759 (N_13759,N_10501,N_11368);
and U13760 (N_13760,N_10657,N_10787);
and U13761 (N_13761,N_11306,N_10271);
nor U13762 (N_13762,N_10174,N_11541);
or U13763 (N_13763,N_11918,N_11826);
nor U13764 (N_13764,N_10421,N_11071);
nand U13765 (N_13765,N_11368,N_10719);
nor U13766 (N_13766,N_11652,N_11111);
or U13767 (N_13767,N_11365,N_11143);
and U13768 (N_13768,N_10460,N_10805);
and U13769 (N_13769,N_10837,N_11263);
nand U13770 (N_13770,N_11570,N_10740);
nor U13771 (N_13771,N_11975,N_11269);
nor U13772 (N_13772,N_11229,N_11257);
nand U13773 (N_13773,N_10428,N_10959);
and U13774 (N_13774,N_10332,N_11519);
nand U13775 (N_13775,N_11862,N_10300);
nor U13776 (N_13776,N_11950,N_11532);
xnor U13777 (N_13777,N_11605,N_11587);
and U13778 (N_13778,N_11047,N_10258);
nand U13779 (N_13779,N_10180,N_11549);
nand U13780 (N_13780,N_10677,N_11577);
or U13781 (N_13781,N_10988,N_10857);
xnor U13782 (N_13782,N_11481,N_11394);
xnor U13783 (N_13783,N_10347,N_10091);
and U13784 (N_13784,N_11869,N_11276);
and U13785 (N_13785,N_10769,N_10500);
or U13786 (N_13786,N_10434,N_11493);
nor U13787 (N_13787,N_10447,N_10664);
nor U13788 (N_13788,N_11940,N_10124);
nand U13789 (N_13789,N_10447,N_11015);
or U13790 (N_13790,N_10913,N_10768);
nand U13791 (N_13791,N_10888,N_11689);
nor U13792 (N_13792,N_11755,N_10755);
and U13793 (N_13793,N_11486,N_11805);
xor U13794 (N_13794,N_11769,N_11950);
xnor U13795 (N_13795,N_10466,N_10032);
nand U13796 (N_13796,N_10986,N_10544);
or U13797 (N_13797,N_11359,N_10451);
nor U13798 (N_13798,N_11034,N_10956);
xor U13799 (N_13799,N_10308,N_11616);
or U13800 (N_13800,N_11040,N_10710);
nand U13801 (N_13801,N_11275,N_11282);
or U13802 (N_13802,N_10602,N_10572);
nand U13803 (N_13803,N_11998,N_10950);
xor U13804 (N_13804,N_10655,N_11651);
or U13805 (N_13805,N_11619,N_10983);
nor U13806 (N_13806,N_10515,N_11397);
nor U13807 (N_13807,N_11338,N_10417);
or U13808 (N_13808,N_10153,N_10179);
and U13809 (N_13809,N_11379,N_10639);
and U13810 (N_13810,N_11863,N_11573);
xor U13811 (N_13811,N_11185,N_11278);
nor U13812 (N_13812,N_11952,N_10156);
nor U13813 (N_13813,N_10792,N_10032);
nand U13814 (N_13814,N_11346,N_11747);
nand U13815 (N_13815,N_10738,N_11011);
or U13816 (N_13816,N_11487,N_11879);
nand U13817 (N_13817,N_11582,N_10971);
and U13818 (N_13818,N_11581,N_11915);
nor U13819 (N_13819,N_11437,N_11849);
and U13820 (N_13820,N_10613,N_10729);
or U13821 (N_13821,N_10366,N_11692);
and U13822 (N_13822,N_11277,N_11373);
or U13823 (N_13823,N_10350,N_10670);
and U13824 (N_13824,N_10577,N_11718);
xnor U13825 (N_13825,N_11021,N_11796);
nand U13826 (N_13826,N_10141,N_11883);
or U13827 (N_13827,N_11225,N_11559);
or U13828 (N_13828,N_10121,N_10085);
or U13829 (N_13829,N_11609,N_11758);
or U13830 (N_13830,N_11460,N_10484);
nor U13831 (N_13831,N_10886,N_10026);
nor U13832 (N_13832,N_10029,N_11585);
or U13833 (N_13833,N_10684,N_11772);
nor U13834 (N_13834,N_10502,N_11174);
or U13835 (N_13835,N_11473,N_11899);
nor U13836 (N_13836,N_10641,N_10717);
nor U13837 (N_13837,N_10569,N_10984);
and U13838 (N_13838,N_10389,N_11054);
nor U13839 (N_13839,N_11315,N_10575);
or U13840 (N_13840,N_11913,N_10145);
nor U13841 (N_13841,N_10047,N_11094);
or U13842 (N_13842,N_10863,N_10716);
and U13843 (N_13843,N_10658,N_10655);
or U13844 (N_13844,N_11756,N_11442);
or U13845 (N_13845,N_10843,N_11312);
and U13846 (N_13846,N_11864,N_10953);
nand U13847 (N_13847,N_10004,N_11914);
or U13848 (N_13848,N_11927,N_10881);
xnor U13849 (N_13849,N_10274,N_10715);
or U13850 (N_13850,N_10349,N_11957);
or U13851 (N_13851,N_11523,N_10380);
nor U13852 (N_13852,N_11932,N_10544);
and U13853 (N_13853,N_10116,N_11735);
and U13854 (N_13854,N_10592,N_11096);
nand U13855 (N_13855,N_11677,N_10103);
xnor U13856 (N_13856,N_11888,N_10859);
nand U13857 (N_13857,N_10005,N_10386);
nand U13858 (N_13858,N_11979,N_11544);
or U13859 (N_13859,N_11867,N_11396);
and U13860 (N_13860,N_11780,N_10648);
and U13861 (N_13861,N_10302,N_11884);
nor U13862 (N_13862,N_11217,N_10140);
or U13863 (N_13863,N_11855,N_10266);
or U13864 (N_13864,N_10921,N_10975);
and U13865 (N_13865,N_11274,N_11489);
nand U13866 (N_13866,N_10922,N_11349);
or U13867 (N_13867,N_10844,N_10318);
and U13868 (N_13868,N_11805,N_10933);
xnor U13869 (N_13869,N_10781,N_10575);
nor U13870 (N_13870,N_10306,N_11827);
or U13871 (N_13871,N_10508,N_10179);
or U13872 (N_13872,N_11245,N_11505);
or U13873 (N_13873,N_10945,N_11924);
or U13874 (N_13874,N_11990,N_10735);
and U13875 (N_13875,N_11265,N_11429);
nor U13876 (N_13876,N_10666,N_10917);
or U13877 (N_13877,N_10375,N_11297);
xor U13878 (N_13878,N_11745,N_10602);
and U13879 (N_13879,N_10098,N_10534);
nor U13880 (N_13880,N_11553,N_10476);
nor U13881 (N_13881,N_11943,N_10305);
nor U13882 (N_13882,N_11917,N_11772);
nor U13883 (N_13883,N_10508,N_10615);
nand U13884 (N_13884,N_11058,N_11272);
nor U13885 (N_13885,N_10557,N_11612);
nand U13886 (N_13886,N_11339,N_10265);
nand U13887 (N_13887,N_11761,N_11924);
and U13888 (N_13888,N_11379,N_11343);
nand U13889 (N_13889,N_10110,N_10832);
nor U13890 (N_13890,N_10927,N_10782);
nor U13891 (N_13891,N_11931,N_10580);
nor U13892 (N_13892,N_11092,N_11136);
and U13893 (N_13893,N_11122,N_11171);
xor U13894 (N_13894,N_10199,N_11334);
nand U13895 (N_13895,N_10702,N_11341);
nor U13896 (N_13896,N_10378,N_11547);
or U13897 (N_13897,N_11553,N_11712);
and U13898 (N_13898,N_10634,N_11308);
nand U13899 (N_13899,N_10298,N_11765);
or U13900 (N_13900,N_11065,N_11086);
or U13901 (N_13901,N_10579,N_11930);
or U13902 (N_13902,N_11746,N_11148);
nor U13903 (N_13903,N_10648,N_10819);
nand U13904 (N_13904,N_11390,N_11415);
or U13905 (N_13905,N_11974,N_11217);
nor U13906 (N_13906,N_10857,N_11377);
or U13907 (N_13907,N_10506,N_10404);
and U13908 (N_13908,N_11991,N_11089);
nand U13909 (N_13909,N_11246,N_11938);
or U13910 (N_13910,N_10540,N_11845);
nor U13911 (N_13911,N_10707,N_10051);
or U13912 (N_13912,N_10165,N_10263);
nor U13913 (N_13913,N_10951,N_10379);
nor U13914 (N_13914,N_11854,N_11170);
or U13915 (N_13915,N_11885,N_10866);
nand U13916 (N_13916,N_11180,N_10848);
nor U13917 (N_13917,N_10979,N_11979);
nand U13918 (N_13918,N_10069,N_10828);
nand U13919 (N_13919,N_10755,N_10579);
nor U13920 (N_13920,N_11096,N_10364);
xor U13921 (N_13921,N_10650,N_10866);
and U13922 (N_13922,N_11524,N_11183);
nor U13923 (N_13923,N_10461,N_10350);
nor U13924 (N_13924,N_10743,N_11470);
and U13925 (N_13925,N_10523,N_11111);
nand U13926 (N_13926,N_11661,N_11554);
or U13927 (N_13927,N_10688,N_10750);
and U13928 (N_13928,N_10749,N_10645);
nand U13929 (N_13929,N_11836,N_10054);
nor U13930 (N_13930,N_10538,N_11515);
and U13931 (N_13931,N_11752,N_10017);
nor U13932 (N_13932,N_10113,N_10325);
and U13933 (N_13933,N_11499,N_10424);
or U13934 (N_13934,N_11400,N_10685);
nand U13935 (N_13935,N_10821,N_11390);
xnor U13936 (N_13936,N_11390,N_10914);
nor U13937 (N_13937,N_10436,N_11647);
or U13938 (N_13938,N_10109,N_10802);
or U13939 (N_13939,N_11182,N_11262);
nor U13940 (N_13940,N_10342,N_11916);
nor U13941 (N_13941,N_11700,N_10153);
nor U13942 (N_13942,N_10830,N_10378);
nor U13943 (N_13943,N_10013,N_11760);
nand U13944 (N_13944,N_11632,N_10793);
nand U13945 (N_13945,N_10065,N_11590);
or U13946 (N_13946,N_10300,N_11458);
nand U13947 (N_13947,N_10342,N_11987);
xor U13948 (N_13948,N_11298,N_10919);
nand U13949 (N_13949,N_10902,N_10589);
and U13950 (N_13950,N_10707,N_11122);
nor U13951 (N_13951,N_11772,N_11036);
and U13952 (N_13952,N_11842,N_11548);
nor U13953 (N_13953,N_11989,N_11862);
or U13954 (N_13954,N_11278,N_10415);
or U13955 (N_13955,N_11280,N_10632);
or U13956 (N_13956,N_10632,N_11526);
nor U13957 (N_13957,N_10148,N_11936);
nand U13958 (N_13958,N_11353,N_11275);
or U13959 (N_13959,N_11170,N_10851);
xor U13960 (N_13960,N_10477,N_10499);
nor U13961 (N_13961,N_11897,N_10314);
and U13962 (N_13962,N_11553,N_11831);
nand U13963 (N_13963,N_11526,N_11842);
nor U13964 (N_13964,N_11673,N_11670);
nand U13965 (N_13965,N_11891,N_11775);
or U13966 (N_13966,N_10711,N_11274);
and U13967 (N_13967,N_11485,N_11124);
nand U13968 (N_13968,N_11378,N_11101);
xnor U13969 (N_13969,N_11714,N_11393);
nor U13970 (N_13970,N_10390,N_10787);
nor U13971 (N_13971,N_11974,N_10316);
nor U13972 (N_13972,N_11497,N_11496);
and U13973 (N_13973,N_11425,N_10772);
and U13974 (N_13974,N_11925,N_11133);
xnor U13975 (N_13975,N_11401,N_10867);
xnor U13976 (N_13976,N_10443,N_11861);
or U13977 (N_13977,N_11597,N_10891);
and U13978 (N_13978,N_11046,N_11312);
or U13979 (N_13979,N_10689,N_11269);
nand U13980 (N_13980,N_10746,N_10549);
nor U13981 (N_13981,N_11421,N_11460);
and U13982 (N_13982,N_10936,N_11728);
nand U13983 (N_13983,N_10838,N_11530);
nor U13984 (N_13984,N_10857,N_11574);
nor U13985 (N_13985,N_10021,N_10024);
or U13986 (N_13986,N_11401,N_11598);
xor U13987 (N_13987,N_10548,N_11450);
and U13988 (N_13988,N_10693,N_10579);
nor U13989 (N_13989,N_10824,N_10345);
and U13990 (N_13990,N_10848,N_11673);
nand U13991 (N_13991,N_11413,N_11287);
nor U13992 (N_13992,N_10164,N_10130);
nor U13993 (N_13993,N_10783,N_10406);
and U13994 (N_13994,N_10861,N_11875);
xnor U13995 (N_13995,N_10436,N_11702);
nand U13996 (N_13996,N_11912,N_11647);
xnor U13997 (N_13997,N_11599,N_11794);
or U13998 (N_13998,N_11717,N_10592);
nand U13999 (N_13999,N_10013,N_10553);
nor U14000 (N_14000,N_13363,N_12142);
or U14001 (N_14001,N_12084,N_13548);
or U14002 (N_14002,N_12076,N_13440);
or U14003 (N_14003,N_13874,N_13504);
or U14004 (N_14004,N_12549,N_12005);
nor U14005 (N_14005,N_12199,N_13514);
nor U14006 (N_14006,N_12056,N_13312);
and U14007 (N_14007,N_12995,N_12013);
nor U14008 (N_14008,N_12854,N_12976);
nor U14009 (N_14009,N_12702,N_12593);
xor U14010 (N_14010,N_13478,N_13193);
nor U14011 (N_14011,N_13642,N_12295);
or U14012 (N_14012,N_12647,N_12031);
and U14013 (N_14013,N_13802,N_13528);
or U14014 (N_14014,N_12639,N_13487);
nand U14015 (N_14015,N_12413,N_13347);
and U14016 (N_14016,N_12307,N_13643);
nor U14017 (N_14017,N_12725,N_12676);
and U14018 (N_14018,N_13667,N_13554);
nor U14019 (N_14019,N_13865,N_12172);
nand U14020 (N_14020,N_13190,N_13673);
or U14021 (N_14021,N_13819,N_12883);
nand U14022 (N_14022,N_13062,N_13453);
and U14023 (N_14023,N_12646,N_13796);
nand U14024 (N_14024,N_13463,N_13414);
nand U14025 (N_14025,N_12360,N_13471);
and U14026 (N_14026,N_13403,N_13023);
nand U14027 (N_14027,N_12182,N_12934);
and U14028 (N_14028,N_12001,N_13131);
and U14029 (N_14029,N_13812,N_12843);
and U14030 (N_14030,N_13174,N_12048);
or U14031 (N_14031,N_12327,N_13701);
nor U14032 (N_14032,N_12969,N_13452);
and U14033 (N_14033,N_13218,N_12657);
nor U14034 (N_14034,N_13176,N_13445);
nor U14035 (N_14035,N_12195,N_13637);
xor U14036 (N_14036,N_12675,N_12978);
nand U14037 (N_14037,N_12903,N_12718);
nand U14038 (N_14038,N_13575,N_12203);
and U14039 (N_14039,N_12214,N_13014);
xnor U14040 (N_14040,N_13232,N_13607);
nor U14041 (N_14041,N_12333,N_13003);
nor U14042 (N_14042,N_13310,N_12479);
nor U14043 (N_14043,N_12656,N_12862);
or U14044 (N_14044,N_12276,N_13682);
or U14045 (N_14045,N_13481,N_12755);
nor U14046 (N_14046,N_12108,N_13596);
nor U14047 (N_14047,N_12543,N_13676);
or U14048 (N_14048,N_13692,N_13343);
nor U14049 (N_14049,N_13542,N_12074);
or U14050 (N_14050,N_13266,N_12486);
or U14051 (N_14051,N_13231,N_13904);
nand U14052 (N_14052,N_12762,N_13513);
nand U14053 (N_14053,N_12223,N_12331);
nand U14054 (N_14054,N_13495,N_13731);
or U14055 (N_14055,N_12390,N_12292);
nand U14056 (N_14056,N_13750,N_12796);
and U14057 (N_14057,N_13316,N_13457);
nor U14058 (N_14058,N_12899,N_13708);
xor U14059 (N_14059,N_12985,N_13748);
nand U14060 (N_14060,N_12437,N_13636);
nand U14061 (N_14061,N_13256,N_12080);
xnor U14062 (N_14062,N_12627,N_13612);
xor U14063 (N_14063,N_12316,N_13725);
nand U14064 (N_14064,N_13461,N_12283);
and U14065 (N_14065,N_12527,N_13561);
and U14066 (N_14066,N_12880,N_13129);
xor U14067 (N_14067,N_12558,N_12528);
or U14068 (N_14068,N_12085,N_12610);
xor U14069 (N_14069,N_12401,N_12253);
xnor U14070 (N_14070,N_13292,N_13286);
and U14071 (N_14071,N_12918,N_13976);
or U14072 (N_14072,N_12981,N_13301);
nand U14073 (N_14073,N_12857,N_12187);
or U14074 (N_14074,N_12984,N_12865);
or U14075 (N_14075,N_12665,N_13743);
and U14076 (N_14076,N_12119,N_13931);
nor U14077 (N_14077,N_13936,N_12383);
or U14078 (N_14078,N_13883,N_13611);
nand U14079 (N_14079,N_12177,N_13588);
or U14080 (N_14080,N_13520,N_13794);
and U14081 (N_14081,N_12622,N_13905);
or U14082 (N_14082,N_12106,N_12440);
or U14083 (N_14083,N_13069,N_13184);
or U14084 (N_14084,N_12035,N_12231);
and U14085 (N_14085,N_12278,N_12240);
nand U14086 (N_14086,N_13253,N_12094);
nand U14087 (N_14087,N_13727,N_13724);
and U14088 (N_14088,N_13859,N_12291);
or U14089 (N_14089,N_13267,N_13064);
nand U14090 (N_14090,N_12894,N_12033);
nor U14091 (N_14091,N_13776,N_12197);
nor U14092 (N_14092,N_12595,N_12808);
and U14093 (N_14093,N_12208,N_12280);
nand U14094 (N_14094,N_12888,N_12044);
nor U14095 (N_14095,N_13858,N_12858);
or U14096 (N_14096,N_12666,N_12161);
and U14097 (N_14097,N_12576,N_12889);
nor U14098 (N_14098,N_13506,N_12124);
or U14099 (N_14099,N_12077,N_13764);
and U14100 (N_14100,N_12530,N_12949);
and U14101 (N_14101,N_13132,N_13467);
and U14102 (N_14102,N_13001,N_13926);
and U14103 (N_14103,N_12620,N_12709);
nor U14104 (N_14104,N_13470,N_12767);
or U14105 (N_14105,N_12038,N_13744);
nor U14106 (N_14106,N_13918,N_13718);
nand U14107 (N_14107,N_13421,N_12986);
or U14108 (N_14108,N_13197,N_12046);
and U14109 (N_14109,N_12042,N_13043);
nand U14110 (N_14110,N_13067,N_13328);
and U14111 (N_14111,N_13112,N_13051);
nand U14112 (N_14112,N_12990,N_13071);
or U14113 (N_14113,N_13780,N_12310);
nor U14114 (N_14114,N_13818,N_13582);
and U14115 (N_14115,N_13877,N_12623);
or U14116 (N_14116,N_13547,N_13208);
or U14117 (N_14117,N_13843,N_12293);
nor U14118 (N_14118,N_13978,N_13412);
xor U14119 (N_14119,N_13498,N_12554);
nor U14120 (N_14120,N_12600,N_12839);
nor U14121 (N_14121,N_12217,N_13095);
nand U14122 (N_14122,N_13034,N_13657);
or U14123 (N_14123,N_12111,N_12163);
and U14124 (N_14124,N_12251,N_13924);
or U14125 (N_14125,N_13117,N_12658);
or U14126 (N_14126,N_13140,N_12287);
or U14127 (N_14127,N_13177,N_13317);
nand U14128 (N_14128,N_13852,N_13035);
and U14129 (N_14129,N_13885,N_12218);
and U14130 (N_14130,N_12348,N_12375);
nand U14131 (N_14131,N_12999,N_12419);
nand U14132 (N_14132,N_12186,N_12215);
nand U14133 (N_14133,N_13124,N_12777);
nand U14134 (N_14134,N_12745,N_12881);
nor U14135 (N_14135,N_13960,N_12550);
or U14136 (N_14136,N_12257,N_12015);
nor U14137 (N_14137,N_12460,N_12022);
nor U14138 (N_14138,N_13222,N_12536);
nor U14139 (N_14139,N_13333,N_12566);
or U14140 (N_14140,N_12249,N_12443);
and U14141 (N_14141,N_12176,N_13148);
xor U14142 (N_14142,N_12737,N_13494);
nand U14143 (N_14143,N_12313,N_13969);
and U14144 (N_14144,N_13653,N_13015);
xnor U14145 (N_14145,N_13223,N_13703);
nor U14146 (N_14146,N_13128,N_12628);
nor U14147 (N_14147,N_12933,N_12897);
and U14148 (N_14148,N_13961,N_12556);
xnor U14149 (N_14149,N_13161,N_12258);
nand U14150 (N_14150,N_13726,N_12655);
nor U14151 (N_14151,N_12043,N_12006);
nand U14152 (N_14152,N_13754,N_13785);
or U14153 (N_14153,N_13675,N_12630);
or U14154 (N_14154,N_13138,N_13915);
and U14155 (N_14155,N_12326,N_13787);
or U14156 (N_14156,N_12099,N_12389);
nor U14157 (N_14157,N_13056,N_12606);
and U14158 (N_14158,N_12029,N_13398);
nand U14159 (N_14159,N_13534,N_13570);
and U14160 (N_14160,N_13334,N_13932);
xnor U14161 (N_14161,N_12194,N_12241);
nor U14162 (N_14162,N_12863,N_12663);
nand U14163 (N_14163,N_13766,N_12830);
nand U14164 (N_14164,N_13974,N_13850);
and U14165 (N_14165,N_13216,N_12707);
nor U14166 (N_14166,N_12040,N_13006);
nand U14167 (N_14167,N_12359,N_12632);
nand U14168 (N_14168,N_13214,N_12114);
nor U14169 (N_14169,N_12886,N_13991);
nor U14170 (N_14170,N_12403,N_13171);
nor U14171 (N_14171,N_12004,N_13650);
or U14172 (N_14172,N_12497,N_13428);
xor U14173 (N_14173,N_13597,N_12008);
nand U14174 (N_14174,N_13426,N_13121);
nand U14175 (N_14175,N_12588,N_12929);
nor U14176 (N_14176,N_13104,N_13631);
nand U14177 (N_14177,N_13450,N_13389);
or U14178 (N_14178,N_12580,N_12466);
nand U14179 (N_14179,N_12651,N_12578);
and U14180 (N_14180,N_13097,N_13691);
nor U14181 (N_14181,N_12757,N_12132);
nand U14182 (N_14182,N_12164,N_13359);
xor U14183 (N_14183,N_13045,N_13666);
and U14184 (N_14184,N_13011,N_13665);
or U14185 (N_14185,N_12175,N_13732);
or U14186 (N_14186,N_13878,N_12159);
nor U14187 (N_14187,N_13116,N_13309);
nor U14188 (N_14188,N_12621,N_13620);
nand U14189 (N_14189,N_12242,N_12394);
and U14190 (N_14190,N_12225,N_13917);
nand U14191 (N_14191,N_12179,N_13734);
or U14192 (N_14192,N_12871,N_13801);
xnor U14193 (N_14193,N_12642,N_12321);
xnor U14194 (N_14194,N_13145,N_13322);
nand U14195 (N_14195,N_13984,N_12786);
nor U14196 (N_14196,N_12547,N_13122);
and U14197 (N_14197,N_12488,N_12330);
and U14198 (N_14198,N_13981,N_12815);
or U14199 (N_14199,N_12461,N_12724);
nand U14200 (N_14200,N_13605,N_12983);
xnor U14201 (N_14201,N_12589,N_12407);
nand U14202 (N_14202,N_13916,N_12431);
and U14203 (N_14203,N_12396,N_12067);
xor U14204 (N_14204,N_12607,N_12664);
or U14205 (N_14205,N_13661,N_12212);
and U14206 (N_14206,N_12958,N_12055);
xor U14207 (N_14207,N_12246,N_13871);
xor U14208 (N_14208,N_12797,N_12299);
nor U14209 (N_14209,N_13873,N_13304);
xnor U14210 (N_14210,N_13532,N_12935);
or U14211 (N_14211,N_13672,N_13048);
and U14212 (N_14212,N_12244,N_12446);
xnor U14213 (N_14213,N_13459,N_12727);
and U14214 (N_14214,N_12802,N_12343);
nand U14215 (N_14215,N_12229,N_12157);
xor U14216 (N_14216,N_13963,N_12977);
nor U14217 (N_14217,N_12311,N_13261);
nand U14218 (N_14218,N_12350,N_13540);
xnor U14219 (N_14219,N_13385,N_13390);
or U14220 (N_14220,N_13375,N_13060);
nand U14221 (N_14221,N_12063,N_12890);
xor U14222 (N_14222,N_12648,N_12422);
nand U14223 (N_14223,N_12155,N_13146);
or U14224 (N_14224,N_13427,N_13752);
and U14225 (N_14225,N_13294,N_13560);
nor U14226 (N_14226,N_13861,N_13980);
or U14227 (N_14227,N_12129,N_12586);
nand U14228 (N_14228,N_13770,N_12332);
nor U14229 (N_14229,N_13930,N_12139);
and U14230 (N_14230,N_13629,N_13654);
or U14231 (N_14231,N_13757,N_13272);
and U14232 (N_14232,N_13568,N_13903);
nand U14233 (N_14233,N_12785,N_13751);
nor U14234 (N_14234,N_12388,N_12480);
nor U14235 (N_14235,N_12661,N_13464);
and U14236 (N_14236,N_12104,N_12418);
or U14237 (N_14237,N_12659,N_12420);
nor U14238 (N_14238,N_12302,N_12109);
or U14239 (N_14239,N_13920,N_12495);
or U14240 (N_14240,N_13603,N_13625);
and U14241 (N_14241,N_13585,N_12377);
nor U14242 (N_14242,N_12211,N_13287);
nand U14243 (N_14243,N_12478,N_13712);
or U14244 (N_14244,N_12714,N_13279);
and U14245 (N_14245,N_13408,N_12914);
xor U14246 (N_14246,N_12510,N_13892);
nor U14247 (N_14247,N_13762,N_13291);
nand U14248 (N_14248,N_12694,N_12619);
or U14249 (N_14249,N_12361,N_13820);
or U14250 (N_14250,N_12517,N_13063);
and U14251 (N_14251,N_12684,N_12943);
nand U14252 (N_14252,N_12784,N_12732);
nor U14253 (N_14253,N_13736,N_12692);
nor U14254 (N_14254,N_12054,N_13400);
nand U14255 (N_14255,N_13477,N_12425);
nand U14256 (N_14256,N_12384,N_12221);
nor U14257 (N_14257,N_12456,N_13943);
nand U14258 (N_14258,N_13350,N_12266);
or U14259 (N_14259,N_13810,N_13988);
nor U14260 (N_14260,N_13302,N_13678);
xor U14261 (N_14261,N_13613,N_12907);
and U14262 (N_14262,N_12970,N_13944);
or U14263 (N_14263,N_13690,N_12449);
and U14264 (N_14264,N_12393,N_13900);
and U14265 (N_14265,N_12220,N_13893);
and U14266 (N_14266,N_13289,N_13965);
or U14267 (N_14267,N_13402,N_13424);
nor U14268 (N_14268,N_12546,N_12645);
and U14269 (N_14269,N_13630,N_12275);
and U14270 (N_14270,N_13220,N_13601);
and U14271 (N_14271,N_13243,N_13996);
nor U14272 (N_14272,N_12806,N_12509);
xnor U14273 (N_14273,N_13881,N_12465);
and U14274 (N_14274,N_12412,N_12135);
nand U14275 (N_14275,N_13016,N_13986);
nor U14276 (N_14276,N_12216,N_13880);
and U14277 (N_14277,N_12869,N_12994);
nand U14278 (N_14278,N_12859,N_13913);
and U14279 (N_14279,N_12710,N_12640);
and U14280 (N_14280,N_12234,N_13795);
and U14281 (N_14281,N_13137,N_12691);
or U14282 (N_14282,N_12496,N_13999);
nand U14283 (N_14283,N_13441,N_12152);
xor U14284 (N_14284,N_13444,N_13153);
nor U14285 (N_14285,N_12968,N_13349);
and U14286 (N_14286,N_13092,N_12930);
and U14287 (N_14287,N_13353,N_13182);
and U14288 (N_14288,N_12128,N_12565);
nor U14289 (N_14289,N_13434,N_12491);
xnor U14290 (N_14290,N_12356,N_13686);
xor U14291 (N_14291,N_12344,N_13499);
xor U14292 (N_14292,N_12531,N_13150);
nor U14293 (N_14293,N_12374,N_13431);
or U14294 (N_14294,N_12391,N_13717);
or U14295 (N_14295,N_12538,N_13152);
nand U14296 (N_14296,N_13189,N_12967);
nor U14297 (N_14297,N_13953,N_13646);
and U14298 (N_14298,N_13527,N_13501);
nand U14299 (N_14299,N_12942,N_13055);
nand U14300 (N_14300,N_13524,N_13175);
or U14301 (N_14301,N_12748,N_13536);
nand U14302 (N_14302,N_12272,N_12758);
and U14303 (N_14303,N_13720,N_13922);
or U14304 (N_14304,N_12505,N_12825);
nor U14305 (N_14305,N_13533,N_13139);
nand U14306 (N_14306,N_12909,N_12467);
nand U14307 (N_14307,N_13998,N_12147);
and U14308 (N_14308,N_12312,N_13283);
nor U14309 (N_14309,N_13816,N_12107);
nor U14310 (N_14310,N_13545,N_12637);
nor U14311 (N_14311,N_12036,N_12644);
nand U14312 (N_14312,N_13049,N_13664);
or U14313 (N_14313,N_12790,N_12007);
nand U14314 (N_14314,N_12734,N_13373);
nand U14315 (N_14315,N_12069,N_12463);
nor U14316 (N_14316,N_12701,N_12794);
nor U14317 (N_14317,N_13484,N_12913);
or U14318 (N_14318,N_12392,N_13549);
or U14319 (N_14319,N_12582,N_12030);
and U14320 (N_14320,N_12366,N_13992);
nor U14321 (N_14321,N_13899,N_12851);
and U14322 (N_14322,N_12364,N_12045);
and U14323 (N_14323,N_13050,N_13580);
and U14324 (N_14324,N_12801,N_12116);
or U14325 (N_14325,N_13149,N_12834);
nor U14326 (N_14326,N_12956,N_13107);
nand U14327 (N_14327,N_13094,N_12068);
or U14328 (N_14328,N_12818,N_13351);
nand U14329 (N_14329,N_13352,N_13479);
nand U14330 (N_14330,N_13215,N_13674);
and U14331 (N_14331,N_13233,N_12925);
and U14332 (N_14332,N_13962,N_13017);
or U14333 (N_14333,N_12592,N_12112);
and U14334 (N_14334,N_13516,N_12948);
nor U14335 (N_14335,N_12708,N_12329);
xor U14336 (N_14336,N_13677,N_12338);
nand U14337 (N_14337,N_12000,N_12695);
nor U14338 (N_14338,N_12803,N_12928);
or U14339 (N_14339,N_13746,N_13144);
or U14340 (N_14340,N_13429,N_12380);
and U14341 (N_14341,N_12539,N_12951);
nand U14342 (N_14342,N_12282,N_13659);
nor U14343 (N_14343,N_13250,N_13556);
nand U14344 (N_14344,N_12148,N_13707);
nand U14345 (N_14345,N_13927,N_13244);
and U14346 (N_14346,N_12457,N_12997);
nand U14347 (N_14347,N_13410,N_13699);
nand U14348 (N_14348,N_13123,N_12146);
nand U14349 (N_14349,N_13957,N_12776);
xnor U14350 (N_14350,N_13307,N_12996);
or U14351 (N_14351,N_13245,N_12821);
nand U14352 (N_14352,N_13401,N_12088);
nand U14353 (N_14353,N_13866,N_13010);
nor U14354 (N_14354,N_13374,N_13822);
and U14355 (N_14355,N_13221,N_12832);
nand U14356 (N_14356,N_13258,N_12433);
nor U14357 (N_14357,N_12770,N_12852);
and U14358 (N_14358,N_13476,N_13407);
nand U14359 (N_14359,N_13809,N_12057);
and U14360 (N_14360,N_13046,N_13013);
xnor U14361 (N_14361,N_12097,N_12489);
and U14362 (N_14362,N_13075,N_12095);
xor U14363 (N_14363,N_13337,N_13587);
or U14364 (N_14364,N_12870,N_12091);
xor U14365 (N_14365,N_12286,N_13281);
nor U14366 (N_14366,N_13562,N_13163);
nor U14367 (N_14367,N_13806,N_13681);
nor U14368 (N_14368,N_13005,N_13940);
or U14369 (N_14369,N_12483,N_12256);
and U14370 (N_14370,N_12557,N_13838);
and U14371 (N_14371,N_12542,N_13126);
nor U14372 (N_14372,N_12247,N_13336);
nor U14373 (N_14373,N_12298,N_12733);
nor U14374 (N_14374,N_12974,N_13022);
nor U14375 (N_14375,N_13769,N_13158);
nor U14376 (N_14376,N_13798,N_13381);
or U14377 (N_14377,N_13041,N_13837);
or U14378 (N_14378,N_13827,N_13964);
and U14379 (N_14379,N_12860,N_12945);
or U14380 (N_14380,N_12502,N_12126);
nand U14381 (N_14381,N_13790,N_13781);
nor U14382 (N_14382,N_12923,N_13934);
nor U14383 (N_14383,N_12936,N_12932);
or U14384 (N_14384,N_13951,N_12314);
or U14385 (N_14385,N_13465,N_13552);
xnor U14386 (N_14386,N_12472,N_12868);
or U14387 (N_14387,N_12122,N_13296);
nor U14388 (N_14388,N_12625,N_12156);
nand U14389 (N_14389,N_13950,N_13212);
and U14390 (N_14390,N_12653,N_13308);
or U14391 (N_14391,N_12798,N_13647);
nand U14392 (N_14392,N_12363,N_12255);
or U14393 (N_14393,N_13529,N_13518);
or U14394 (N_14394,N_13098,N_13143);
nand U14395 (N_14395,N_12322,N_12873);
nor U14396 (N_14396,N_12369,N_12494);
nand U14397 (N_14397,N_12944,N_12305);
and U14398 (N_14398,N_12613,N_13517);
or U14399 (N_14399,N_13604,N_12345);
or U14400 (N_14400,N_13007,N_13432);
nand U14401 (N_14401,N_13772,N_12568);
nor U14402 (N_14402,N_13648,N_13417);
nand U14403 (N_14403,N_12540,N_13593);
and U14404 (N_14404,N_13774,N_13728);
nor U14405 (N_14405,N_13422,N_13285);
xnor U14406 (N_14406,N_13468,N_12908);
or U14407 (N_14407,N_13119,N_12477);
and U14408 (N_14408,N_12901,N_13036);
or U14409 (N_14409,N_13165,N_13987);
xor U14410 (N_14410,N_12840,N_13857);
nand U14411 (N_14411,N_13854,N_13592);
nand U14412 (N_14412,N_13070,N_12699);
or U14413 (N_14413,N_13338,N_13270);
nand U14414 (N_14414,N_12533,N_13535);
and U14415 (N_14415,N_13832,N_13366);
or U14416 (N_14416,N_12756,N_13955);
or U14417 (N_14417,N_13945,N_12082);
xor U14418 (N_14418,N_13004,N_12508);
nor U14419 (N_14419,N_12782,N_13037);
or U14420 (N_14420,N_12336,N_13656);
and U14421 (N_14421,N_12975,N_13651);
or U14422 (N_14422,N_13906,N_13155);
and U14423 (N_14423,N_13558,N_13632);
nor U14424 (N_14424,N_13318,N_12768);
nand U14425 (N_14425,N_13571,N_13680);
and U14426 (N_14426,N_12451,N_12026);
nand U14427 (N_14427,N_13668,N_13305);
or U14428 (N_14428,N_12778,N_13644);
and U14429 (N_14429,N_13438,N_13492);
or U14430 (N_14430,N_12749,N_12598);
or U14431 (N_14431,N_13433,N_12306);
xor U14432 (N_14432,N_12219,N_12213);
or U14433 (N_14433,N_12115,N_13888);
and U14434 (N_14434,N_12849,N_13065);
and U14435 (N_14435,N_13559,N_13225);
and U14436 (N_14436,N_13541,N_13685);
xor U14437 (N_14437,N_13509,N_13473);
nor U14438 (N_14438,N_12910,N_13027);
and U14439 (N_14439,N_13073,N_12414);
and U14440 (N_14440,N_12261,N_13357);
or U14441 (N_14441,N_13572,N_12265);
xor U14442 (N_14442,N_12053,N_12340);
nand U14443 (N_14443,N_13392,N_13164);
or U14444 (N_14444,N_12470,N_13263);
or U14445 (N_14445,N_13907,N_12696);
or U14446 (N_14446,N_13324,N_12402);
nand U14447 (N_14447,N_12828,N_13265);
and U14448 (N_14448,N_12826,N_12650);
and U14449 (N_14449,N_13863,N_12300);
and U14450 (N_14450,N_13649,N_12683);
nand U14451 (N_14451,N_13714,N_13199);
nand U14452 (N_14452,N_12188,N_12473);
nand U14453 (N_14453,N_12227,N_13077);
nand U14454 (N_14454,N_12569,N_12847);
or U14455 (N_14455,N_12049,N_13995);
nand U14456 (N_14456,N_13621,N_13971);
nand U14457 (N_14457,N_12183,N_12263);
nand U14458 (N_14458,N_12423,N_12416);
and U14459 (N_14459,N_13130,N_13876);
or U14460 (N_14460,N_12089,N_13723);
and U14461 (N_14461,N_13187,N_12937);
nor U14462 (N_14462,N_12946,N_13985);
nor U14463 (N_14463,N_13230,N_13188);
nor U14464 (N_14464,N_13531,N_13925);
or U14465 (N_14465,N_13135,N_12877);
and U14466 (N_14466,N_12677,N_12285);
xnor U14467 (N_14467,N_13480,N_12406);
nand U14468 (N_14468,N_13949,N_13844);
or U14469 (N_14469,N_12071,N_12075);
and U14470 (N_14470,N_12669,N_12224);
xor U14471 (N_14471,N_12365,N_12952);
or U14472 (N_14472,N_12845,N_12891);
xnor U14473 (N_14473,N_12920,N_12201);
nand U14474 (N_14474,N_12824,N_12501);
xnor U14475 (N_14475,N_13255,N_13923);
nand U14476 (N_14476,N_13713,N_12717);
nand U14477 (N_14477,N_13458,N_12587);
and U14478 (N_14478,N_13160,N_12158);
nand U14479 (N_14479,N_13679,N_12960);
or U14480 (N_14480,N_12602,N_13793);
or U14481 (N_14481,N_12476,N_12562);
nand U14482 (N_14482,N_12335,N_13800);
or U14483 (N_14483,N_12896,N_12130);
or U14484 (N_14484,N_13442,N_13314);
or U14485 (N_14485,N_12079,N_12817);
or U14486 (N_14486,N_12464,N_12713);
or U14487 (N_14487,N_12911,N_12941);
and U14488 (N_14488,N_12515,N_13248);
nand U14489 (N_14489,N_13526,N_13074);
nand U14490 (N_14490,N_13808,N_13078);
nand U14491 (N_14491,N_13898,N_13344);
and U14492 (N_14492,N_13608,N_13271);
or U14493 (N_14493,N_12180,N_12434);
nand U14494 (N_14494,N_12047,N_12017);
nor U14495 (N_14495,N_13490,N_12173);
and U14496 (N_14496,N_13937,N_13044);
nand U14497 (N_14497,N_12585,N_12519);
nor U14498 (N_14498,N_12723,N_12349);
and U14499 (N_14499,N_13869,N_13696);
or U14500 (N_14500,N_12616,N_13275);
xor U14501 (N_14501,N_13186,N_12700);
nand U14502 (N_14502,N_12236,N_13297);
nor U14503 (N_14503,N_12541,N_12685);
or U14504 (N_14504,N_12050,N_13586);
nand U14505 (N_14505,N_13689,N_12222);
and U14506 (N_14506,N_13061,N_12876);
nor U14507 (N_14507,N_12604,N_12424);
nand U14508 (N_14508,N_12511,N_13610);
and U14509 (N_14509,N_12800,N_12237);
nor U14510 (N_14510,N_13142,N_12117);
nor U14511 (N_14511,N_12759,N_13615);
nand U14512 (N_14512,N_13606,N_13404);
or U14513 (N_14513,N_13066,N_13089);
nand U14514 (N_14514,N_12512,N_13977);
or U14515 (N_14515,N_12783,N_13569);
and U14516 (N_14516,N_13823,N_12579);
nand U14517 (N_14517,N_12032,N_13972);
nand U14518 (N_14518,N_12136,N_13093);
or U14519 (N_14519,N_12061,N_13191);
and U14520 (N_14520,N_12636,N_12417);
nor U14521 (N_14521,N_13565,N_12746);
or U14522 (N_14522,N_13979,N_13767);
nand U14523 (N_14523,N_12882,N_12284);
nor U14524 (N_14524,N_13360,N_13747);
nand U14525 (N_14525,N_12105,N_12635);
or U14526 (N_14526,N_13368,N_12697);
nand U14527 (N_14527,N_13765,N_13252);
nor U14528 (N_14528,N_12410,N_12372);
nand U14529 (N_14529,N_13997,N_12917);
and U14530 (N_14530,N_13890,N_12601);
or U14531 (N_14531,N_13466,N_12867);
or U14532 (N_14532,N_13209,N_12319);
and U14533 (N_14533,N_12200,N_12740);
nand U14534 (N_14534,N_12339,N_12864);
and U14535 (N_14535,N_12649,N_12445);
nor U14536 (N_14536,N_12688,N_12181);
and U14537 (N_14537,N_12435,N_12673);
nor U14538 (N_14538,N_12788,N_12207);
and U14539 (N_14539,N_12706,N_12453);
nand U14540 (N_14540,N_12544,N_13180);
and U14541 (N_14541,N_13617,N_13895);
or U14542 (N_14542,N_13614,N_13183);
nand U14543 (N_14543,N_12703,N_13897);
or U14544 (N_14544,N_12705,N_12792);
and U14545 (N_14545,N_13356,N_13326);
and U14546 (N_14546,N_13990,N_13577);
nor U14547 (N_14547,N_13566,N_12320);
or U14548 (N_14548,N_12603,N_12426);
and U14549 (N_14549,N_12002,N_13544);
and U14550 (N_14550,N_12421,N_13099);
or U14551 (N_14551,N_13573,N_12772);
and U14552 (N_14552,N_12334,N_13179);
nor U14553 (N_14553,N_13740,N_13578);
or U14554 (N_14554,N_12317,N_13460);
or U14555 (N_14555,N_12151,N_12775);
or U14556 (N_14556,N_12900,N_12034);
nand U14557 (N_14557,N_13111,N_12513);
nor U14558 (N_14558,N_13340,N_12764);
or U14559 (N_14559,N_13113,N_13273);
and U14560 (N_14560,N_12113,N_13567);
nand U14561 (N_14561,N_13523,N_12092);
or U14562 (N_14562,N_12353,N_12475);
nor U14563 (N_14563,N_12140,N_12638);
and U14564 (N_14564,N_13009,N_12634);
or U14565 (N_14565,N_12552,N_12023);
and U14566 (N_14566,N_12535,N_13393);
nand U14567 (N_14567,N_13362,N_13589);
xnor U14568 (N_14568,N_13154,N_12874);
nor U14569 (N_14569,N_13364,N_13634);
nor U14570 (N_14570,N_13378,N_13238);
nor U14571 (N_14571,N_12822,N_12230);
and U14572 (N_14572,N_13911,N_12982);
and U14573 (N_14573,N_13595,N_13815);
or U14574 (N_14574,N_13213,N_13715);
and U14575 (N_14575,N_12243,N_13475);
nand U14576 (N_14576,N_12009,N_12872);
nor U14577 (N_14577,N_13409,N_13327);
nand U14578 (N_14578,N_12855,N_13346);
xnor U14579 (N_14579,N_12884,N_13002);
nand U14580 (N_14580,N_13008,N_13519);
nand U14581 (N_14581,N_13076,N_12016);
nand U14582 (N_14582,N_13594,N_13599);
nor U14583 (N_14583,N_12432,N_13115);
nand U14584 (N_14584,N_12459,N_13737);
or U14585 (N_14585,N_13628,N_13710);
and U14586 (N_14586,N_12325,N_12529);
nor U14587 (N_14587,N_12059,N_13395);
xnor U14588 (N_14588,N_12728,N_13102);
or U14589 (N_14589,N_12083,N_12609);
nor U14590 (N_14590,N_12730,N_13884);
and U14591 (N_14591,N_12351,N_13345);
and U14592 (N_14592,N_12668,N_13387);
nor U14593 (N_14593,N_12354,N_12245);
and U14594 (N_14594,N_12532,N_13942);
and U14595 (N_14595,N_13939,N_12081);
nand U14596 (N_14596,N_12672,N_13025);
or U14597 (N_14597,N_13454,N_13031);
nor U14598 (N_14598,N_13012,N_13797);
nand U14599 (N_14599,N_13227,N_13862);
and U14600 (N_14600,N_13640,N_12827);
nor U14601 (N_14601,N_12596,N_13170);
nor U14602 (N_14602,N_12373,N_12507);
and U14603 (N_14603,N_12526,N_12101);
nand U14604 (N_14604,N_13510,N_12485);
and U14605 (N_14605,N_13226,N_13032);
and U14606 (N_14606,N_13598,N_13619);
nand U14607 (N_14607,N_12210,N_13086);
and U14608 (N_14608,N_12819,N_13719);
xnor U14609 (N_14609,N_12385,N_13280);
and U14610 (N_14610,N_13777,N_13018);
and U14611 (N_14611,N_13211,N_13768);
or U14612 (N_14612,N_12259,N_13488);
xor U14613 (N_14613,N_12612,N_12992);
or U14614 (N_14614,N_12328,N_13331);
nor U14615 (N_14615,N_13057,N_13841);
nor U14616 (N_14616,N_13655,N_13446);
nor U14617 (N_14617,N_12964,N_12720);
nor U14618 (N_14618,N_13928,N_12352);
and U14619 (N_14619,N_13339,N_12617);
and U14620 (N_14620,N_13383,N_12206);
or U14621 (N_14621,N_13497,N_12957);
xnor U14622 (N_14622,N_12003,N_12963);
xor U14623 (N_14623,N_13396,N_13354);
nand U14624 (N_14624,N_13782,N_13616);
or U14625 (N_14625,N_13207,N_13125);
and U14626 (N_14626,N_12814,N_12769);
or U14627 (N_14627,N_12739,N_12583);
nor U14628 (N_14628,N_12838,N_13399);
nand U14629 (N_14629,N_13276,N_13834);
nand U14630 (N_14630,N_13583,N_12209);
nand U14631 (N_14631,N_13083,N_13042);
nand U14632 (N_14632,N_12309,N_13821);
nand U14633 (N_14633,N_13779,N_13716);
and U14634 (N_14634,N_13684,N_13947);
nor U14635 (N_14635,N_12011,N_12831);
and U14636 (N_14636,N_12927,N_12438);
or U14637 (N_14637,N_12503,N_13753);
nor U14638 (N_14638,N_12520,N_13742);
or U14639 (N_14639,N_13448,N_12471);
or U14640 (N_14640,N_12138,N_13749);
nor U14641 (N_14641,N_12027,N_12747);
nor U14642 (N_14642,N_13096,N_13167);
or U14643 (N_14643,N_12973,N_12308);
and U14644 (N_14644,N_13839,N_12678);
or U14645 (N_14645,N_12121,N_12462);
and U14646 (N_14646,N_12409,N_13830);
nand U14647 (N_14647,N_12682,N_12680);
nor U14648 (N_14648,N_12898,N_12875);
and U14649 (N_14649,N_13257,N_13910);
nor U14650 (N_14650,N_12681,N_13386);
and U14651 (N_14651,N_12090,N_13687);
nor U14652 (N_14652,N_12893,N_13688);
nor U14653 (N_14653,N_12143,N_13958);
nor U14654 (N_14654,N_12912,N_13807);
nor U14655 (N_14655,N_12789,N_13472);
xnor U14656 (N_14656,N_12919,N_13994);
or U14657 (N_14657,N_12921,N_13704);
and U14658 (N_14658,N_13376,N_13306);
nand U14659 (N_14659,N_13040,N_13879);
nor U14660 (N_14660,N_13833,N_13938);
nor U14661 (N_14661,N_13786,N_12277);
or U14662 (N_14662,N_13329,N_12025);
nor U14663 (N_14663,N_12885,N_13335);
or U14664 (N_14664,N_13405,N_12185);
and U14665 (N_14665,N_12378,N_12654);
and U14666 (N_14666,N_12807,N_12367);
and U14667 (N_14667,N_12752,N_12563);
and U14668 (N_14668,N_12841,N_12820);
nand U14669 (N_14669,N_13106,N_13705);
nand U14670 (N_14670,N_13553,N_13236);
and U14671 (N_14671,N_13602,N_13038);
and U14672 (N_14672,N_13415,N_13159);
nor U14673 (N_14673,N_13966,N_12358);
and U14674 (N_14674,N_13799,N_13970);
or U14675 (N_14675,N_13730,N_12805);
and U14676 (N_14676,N_12922,N_12110);
nor U14677 (N_14677,N_13537,N_13663);
nor U14678 (N_14678,N_12850,N_13447);
or U14679 (N_14679,N_12368,N_13320);
nand U14680 (N_14680,N_12448,N_12481);
nor U14681 (N_14681,N_12386,N_12341);
and U14682 (N_14682,N_12271,N_13254);
nand U14683 (N_14683,N_13219,N_12584);
nand U14684 (N_14684,N_13711,N_13455);
nor U14685 (N_14685,N_13058,N_13127);
nand U14686 (N_14686,N_13321,N_13729);
or U14687 (N_14687,N_13872,N_12235);
and U14688 (N_14688,N_12987,N_12267);
and U14689 (N_14689,N_12493,N_12738);
and U14690 (N_14690,N_12518,N_13835);
or U14691 (N_14691,N_12490,N_13842);
and U14692 (N_14692,N_12051,N_12452);
and U14693 (N_14693,N_12765,N_12264);
xnor U14694 (N_14694,N_13982,N_12064);
nor U14695 (N_14695,N_12773,N_13557);
nor U14696 (N_14696,N_13456,N_12039);
or U14697 (N_14697,N_13300,N_13550);
and U14698 (N_14698,N_12743,N_12395);
xnor U14699 (N_14699,N_13848,N_13700);
and U14700 (N_14700,N_13901,N_12915);
and U14701 (N_14701,N_12014,N_12611);
and U14702 (N_14702,N_12905,N_13217);
nand U14703 (N_14703,N_13192,N_13436);
or U14704 (N_14704,N_12581,N_12170);
or U14705 (N_14705,N_13581,N_12131);
nand U14706 (N_14706,N_13469,N_12953);
nor U14707 (N_14707,N_13671,N_13068);
nor U14708 (N_14708,N_13914,N_12268);
nand U14709 (N_14709,N_12980,N_12506);
and U14710 (N_14710,N_12629,N_12561);
nand U14711 (N_14711,N_13909,N_12741);
or U14712 (N_14712,N_13406,N_13278);
nor U14713 (N_14713,N_12498,N_12525);
nand U14714 (N_14714,N_13288,N_12123);
or U14715 (N_14715,N_12904,N_12761);
nor U14716 (N_14716,N_13311,N_13775);
or U14717 (N_14717,N_13627,N_13298);
nor U14718 (N_14718,N_13206,N_12428);
and U14719 (N_14719,N_12545,N_13493);
xor U14720 (N_14720,N_12371,N_12078);
nand U14721 (N_14721,N_12816,N_13855);
or U14722 (N_14722,N_13348,N_12020);
nor U14723 (N_14723,N_13449,N_13954);
or U14724 (N_14724,N_12398,N_12174);
nand U14725 (N_14725,N_12149,N_12193);
and U14726 (N_14726,N_12252,N_13251);
or U14727 (N_14727,N_12835,N_13539);
xor U14728 (N_14728,N_13948,N_13846);
nor U14729 (N_14729,N_12381,N_12763);
or U14730 (N_14730,N_12754,N_12297);
nand U14731 (N_14731,N_13959,N_12861);
nand U14732 (N_14732,N_13262,N_13973);
nand U14733 (N_14733,N_12548,N_13935);
nor U14734 (N_14734,N_13543,N_12399);
nor U14735 (N_14735,N_13662,N_13956);
nor U14736 (N_14736,N_12066,N_13829);
and U14737 (N_14737,N_13169,N_13147);
nand U14738 (N_14738,N_13435,N_12346);
nor U14739 (N_14739,N_12189,N_12662);
or U14740 (N_14740,N_12288,N_13683);
nor U14741 (N_14741,N_12560,N_13882);
or U14742 (N_14742,N_12400,N_12735);
nor U14743 (N_14743,N_12966,N_13443);
or U14744 (N_14744,N_13201,N_13551);
xnor U14745 (N_14745,N_13847,N_13079);
nor U14746 (N_14746,N_12450,N_13763);
or U14747 (N_14747,N_13024,N_12134);
and U14748 (N_14748,N_13864,N_12833);
or U14749 (N_14749,N_13875,N_12906);
nor U14750 (N_14750,N_13355,N_12093);
nor U14751 (N_14751,N_12184,N_12404);
nand U14752 (N_14752,N_12631,N_13411);
or U14753 (N_14753,N_12774,N_12771);
xor U14754 (N_14754,N_13052,N_12166);
and U14755 (N_14755,N_12940,N_12690);
nor U14756 (N_14756,N_12924,N_12301);
nand U14757 (N_14757,N_12150,N_13641);
and U14758 (N_14758,N_12813,N_13284);
and U14759 (N_14759,N_13109,N_12524);
and U14760 (N_14760,N_13849,N_13805);
and U14761 (N_14761,N_12070,N_12098);
xor U14762 (N_14762,N_12687,N_13521);
nor U14763 (N_14763,N_12514,N_12127);
and U14764 (N_14764,N_12988,N_13921);
or U14765 (N_14765,N_13639,N_13856);
nand U14766 (N_14766,N_12742,N_12028);
and U14767 (N_14767,N_12296,N_13778);
and U14768 (N_14768,N_12469,N_12991);
nor U14769 (N_14769,N_12671,N_12073);
and U14770 (N_14770,N_12021,N_13303);
nand U14771 (N_14771,N_12290,N_13546);
and U14772 (N_14772,N_13622,N_13087);
nand U14773 (N_14773,N_13047,N_13803);
and U14774 (N_14774,N_12590,N_13237);
or U14775 (N_14775,N_13983,N_12153);
nand U14776 (N_14776,N_13451,N_12679);
xor U14777 (N_14777,N_12559,N_13946);
and U14778 (N_14778,N_12721,N_13085);
and U14779 (N_14779,N_12019,N_12643);
or U14780 (N_14780,N_13379,N_13228);
nand U14781 (N_14781,N_12608,N_13204);
or U14782 (N_14782,N_12704,N_12171);
nor U14783 (N_14783,N_13323,N_12787);
and U14784 (N_14784,N_12376,N_12641);
xor U14785 (N_14785,N_13788,N_13235);
or U14786 (N_14786,N_12804,N_12137);
xor U14787 (N_14787,N_12484,N_13397);
nor U14788 (N_14788,N_13110,N_12522);
or U14789 (N_14789,N_13290,N_13249);
nor U14790 (N_14790,N_13889,N_12823);
nand U14791 (N_14791,N_12751,N_13836);
nand U14792 (N_14792,N_12753,N_12411);
nor U14793 (N_14793,N_13755,N_12499);
nor U14794 (N_14794,N_13108,N_13391);
nand U14795 (N_14795,N_13919,N_13845);
xnor U14796 (N_14796,N_12979,N_13826);
or U14797 (N_14797,N_12102,N_13332);
or U14798 (N_14798,N_13162,N_13157);
and U14799 (N_14799,N_12415,N_13054);
nor U14800 (N_14800,N_12196,N_12564);
xor U14801 (N_14801,N_13773,N_12304);
and U14802 (N_14802,N_12504,N_12971);
or U14803 (N_14803,N_13029,N_13814);
or U14804 (N_14804,N_13082,N_13416);
xnor U14805 (N_14805,N_13507,N_13658);
or U14806 (N_14806,N_13388,N_13342);
xor U14807 (N_14807,N_13293,N_13771);
xnor U14808 (N_14808,N_13496,N_13172);
nor U14809 (N_14809,N_13824,N_12444);
nor U14810 (N_14810,N_13319,N_12041);
and U14811 (N_14811,N_13886,N_13600);
nand U14812 (N_14812,N_13229,N_13522);
and U14813 (N_14813,N_12715,N_12248);
nand U14814 (N_14814,N_13330,N_12315);
nor U14815 (N_14815,N_13735,N_12719);
nand U14816 (N_14816,N_13502,N_13538);
or U14817 (N_14817,N_12947,N_13828);
nor U14818 (N_14818,N_13259,N_12144);
nor U14819 (N_14819,N_13084,N_12262);
xnor U14820 (N_14820,N_13804,N_12442);
xnor U14821 (N_14821,N_12058,N_13313);
and U14822 (N_14822,N_13891,N_13579);
nor U14823 (N_14823,N_13246,N_12289);
or U14824 (N_14824,N_12439,N_12848);
or U14825 (N_14825,N_12052,N_12712);
and U14826 (N_14826,N_12534,N_13439);
nor U14827 (N_14827,N_13500,N_13840);
and U14828 (N_14828,N_13369,N_12811);
xor U14829 (N_14829,N_13420,N_13028);
nand U14830 (N_14830,N_12178,N_12689);
nor U14831 (N_14831,N_12024,N_12455);
and U14832 (N_14832,N_13020,N_13196);
and U14833 (N_14833,N_13555,N_12793);
or U14834 (N_14834,N_12204,N_13134);
nor U14835 (N_14835,N_12780,N_12998);
xnor U14836 (N_14836,N_13299,N_13260);
xnor U14837 (N_14837,N_12516,N_12430);
and U14838 (N_14838,N_12100,N_12318);
nand U14839 (N_14839,N_12162,N_13738);
or U14840 (N_14840,N_12760,N_12118);
nor U14841 (N_14841,N_13817,N_12429);
or U14842 (N_14842,N_12674,N_13791);
nor U14843 (N_14843,N_12693,N_13091);
nor U14844 (N_14844,N_13745,N_13512);
nor U14845 (N_14845,N_12303,N_12594);
nor U14846 (N_14846,N_13242,N_12145);
nand U14847 (N_14847,N_12744,N_12190);
xnor U14848 (N_14848,N_13792,N_13853);
nand U14849 (N_14849,N_12955,N_12273);
nand U14850 (N_14850,N_13105,N_12686);
xnor U14851 (N_14851,N_12574,N_13194);
nor U14852 (N_14852,N_13133,N_12408);
and U14853 (N_14853,N_13574,N_13341);
nor U14854 (N_14854,N_13968,N_12591);
or U14855 (N_14855,N_13059,N_12614);
nand U14856 (N_14856,N_12938,N_12037);
nand U14857 (N_14857,N_12939,N_13722);
nor U14858 (N_14858,N_13413,N_12362);
nand U14859 (N_14859,N_13693,N_12096);
nor U14860 (N_14860,N_13365,N_13000);
or U14861 (N_14861,N_12087,N_12781);
or U14862 (N_14862,N_12120,N_13491);
nor U14863 (N_14863,N_13367,N_12324);
nand U14864 (N_14864,N_12895,N_13706);
nor U14865 (N_14865,N_12103,N_12167);
and U14866 (N_14866,N_13181,N_13315);
nor U14867 (N_14867,N_13896,N_13274);
or U14868 (N_14868,N_13168,N_12323);
or U14869 (N_14869,N_13623,N_12279);
nand U14870 (N_14870,N_13825,N_13173);
or U14871 (N_14871,N_12698,N_13989);
nand U14872 (N_14872,N_12766,N_12624);
and U14873 (N_14873,N_12573,N_13277);
and U14874 (N_14874,N_13384,N_13645);
or U14875 (N_14875,N_13241,N_12487);
or U14876 (N_14876,N_13090,N_12626);
or U14877 (N_14877,N_13761,N_12337);
nor U14878 (N_14878,N_12141,N_13239);
nor U14879 (N_14879,N_13026,N_13030);
or U14880 (N_14880,N_13198,N_13660);
nand U14881 (N_14881,N_13166,N_13503);
and U14882 (N_14882,N_13633,N_12233);
nor U14883 (N_14883,N_12065,N_12812);
or U14884 (N_14884,N_12887,N_13205);
nand U14885 (N_14885,N_13697,N_12270);
nor U14886 (N_14886,N_12436,N_13887);
nand U14887 (N_14887,N_12916,N_13462);
nor U14888 (N_14888,N_12260,N_13425);
nor U14889 (N_14889,N_13894,N_13624);
nor U14890 (N_14890,N_12567,N_12160);
xnor U14891 (N_14891,N_12447,N_13377);
xnor U14892 (N_14892,N_12599,N_12670);
or U14893 (N_14893,N_13789,N_12125);
nor U14894 (N_14894,N_13505,N_13269);
nand U14895 (N_14895,N_12018,N_12192);
and U14896 (N_14896,N_12468,N_13698);
xnor U14897 (N_14897,N_12667,N_13702);
or U14898 (N_14898,N_13072,N_13993);
xnor U14899 (N_14899,N_12878,N_12228);
nand U14900 (N_14900,N_12853,N_13860);
xnor U14901 (N_14901,N_13372,N_13361);
and U14902 (N_14902,N_13576,N_13967);
or U14903 (N_14903,N_13902,N_13394);
and U14904 (N_14904,N_12474,N_12405);
nand U14905 (N_14905,N_12555,N_13721);
nand U14906 (N_14906,N_13114,N_13423);
and U14907 (N_14907,N_12731,N_12269);
nand U14908 (N_14908,N_13870,N_13136);
or U14909 (N_14909,N_13088,N_12198);
nor U14910 (N_14910,N_13525,N_12856);
nand U14911 (N_14911,N_12799,N_12012);
nand U14912 (N_14912,N_12810,N_12846);
nand U14913 (N_14913,N_12716,N_13564);
xnor U14914 (N_14914,N_12355,N_12482);
or U14915 (N_14915,N_12086,N_13831);
nand U14916 (N_14916,N_13419,N_13638);
nand U14917 (N_14917,N_12226,N_12010);
nand U14918 (N_14918,N_12294,N_13952);
nor U14919 (N_14919,N_13185,N_12342);
and U14920 (N_14920,N_13590,N_13511);
nor U14921 (N_14921,N_12570,N_12729);
nor U14922 (N_14922,N_13234,N_12993);
nor U14923 (N_14923,N_13609,N_13100);
nand U14924 (N_14924,N_13482,N_12072);
nor U14925 (N_14925,N_13584,N_13485);
nand U14926 (N_14926,N_12842,N_12926);
nor U14927 (N_14927,N_13867,N_12633);
and U14928 (N_14928,N_12779,N_12521);
nand U14929 (N_14929,N_12597,N_12837);
and U14930 (N_14930,N_12618,N_12954);
nand U14931 (N_14931,N_13733,N_13695);
and U14932 (N_14932,N_12454,N_13975);
nor U14933 (N_14933,N_12441,N_13515);
xor U14934 (N_14934,N_12711,N_13120);
and U14935 (N_14935,N_13430,N_12060);
nor U14936 (N_14936,N_13295,N_13813);
nand U14937 (N_14937,N_12722,N_13033);
nor U14938 (N_14938,N_13039,N_12357);
or U14939 (N_14939,N_12572,N_13380);
xor U14940 (N_14940,N_12492,N_13210);
nand U14941 (N_14941,N_13268,N_13240);
nor U14942 (N_14942,N_12551,N_12726);
or U14943 (N_14943,N_12154,N_13739);
or U14944 (N_14944,N_12062,N_12205);
or U14945 (N_14945,N_12133,N_13933);
nor U14946 (N_14946,N_13811,N_12605);
xnor U14947 (N_14947,N_13200,N_12829);
or U14948 (N_14948,N_13635,N_12250);
nand U14949 (N_14949,N_13382,N_12169);
nor U14950 (N_14950,N_13741,N_12931);
nand U14951 (N_14951,N_12866,N_12165);
and U14952 (N_14952,N_13195,N_13912);
nand U14953 (N_14953,N_12961,N_13941);
xnor U14954 (N_14954,N_13202,N_13486);
nand U14955 (N_14955,N_12962,N_13929);
or U14956 (N_14956,N_12959,N_12950);
nand U14957 (N_14957,N_12660,N_12382);
nand U14958 (N_14958,N_13080,N_12879);
nand U14959 (N_14959,N_12902,N_12274);
or U14960 (N_14960,N_12571,N_12537);
xnor U14961 (N_14961,N_13652,N_12791);
xnor U14962 (N_14962,N_12836,N_13618);
and U14963 (N_14963,N_12844,N_12281);
or U14964 (N_14964,N_13053,N_12615);
nand U14965 (N_14965,N_12347,N_12795);
and U14966 (N_14966,N_13669,N_13626);
or U14967 (N_14967,N_12972,N_12370);
and U14968 (N_14968,N_13591,N_13264);
nand U14969 (N_14969,N_13325,N_13483);
or U14970 (N_14970,N_13370,N_13437);
nand U14971 (N_14971,N_13759,N_13908);
and U14972 (N_14972,N_13530,N_13563);
and U14973 (N_14973,N_13868,N_13670);
nand U14974 (N_14974,N_13760,N_12652);
xor U14975 (N_14975,N_12168,N_12191);
nand U14976 (N_14976,N_13019,N_13371);
nor U14977 (N_14977,N_12523,N_13474);
xnor U14978 (N_14978,N_12254,N_13758);
nor U14979 (N_14979,N_13151,N_13203);
and U14980 (N_14980,N_12965,N_13101);
or U14981 (N_14981,N_12458,N_13709);
nand U14982 (N_14982,N_12892,N_12427);
or U14983 (N_14983,N_13118,N_13021);
nand U14984 (N_14984,N_13851,N_12736);
nor U14985 (N_14985,N_12575,N_12387);
and U14986 (N_14986,N_13224,N_13081);
nand U14987 (N_14987,N_12989,N_12500);
nand U14988 (N_14988,N_13783,N_12232);
nor U14989 (N_14989,N_12379,N_13489);
nor U14990 (N_14990,N_12750,N_12577);
or U14991 (N_14991,N_13156,N_13141);
nor U14992 (N_14992,N_12553,N_13103);
and U14993 (N_14993,N_13178,N_12397);
nand U14994 (N_14994,N_13282,N_13756);
and U14995 (N_14995,N_12238,N_13358);
or U14996 (N_14996,N_12809,N_12202);
nor U14997 (N_14997,N_13508,N_12239);
and U14998 (N_14998,N_13694,N_13418);
and U14999 (N_14999,N_13247,N_13784);
and U15000 (N_15000,N_12897,N_12872);
nor U15001 (N_15001,N_13714,N_12399);
xor U15002 (N_15002,N_12600,N_13150);
and U15003 (N_15003,N_12326,N_12082);
or U15004 (N_15004,N_13518,N_13129);
nor U15005 (N_15005,N_13520,N_12727);
and U15006 (N_15006,N_12640,N_13312);
and U15007 (N_15007,N_12395,N_12989);
nor U15008 (N_15008,N_12602,N_12549);
nor U15009 (N_15009,N_12711,N_13978);
or U15010 (N_15010,N_13290,N_12094);
or U15011 (N_15011,N_13787,N_12668);
and U15012 (N_15012,N_13005,N_12211);
nand U15013 (N_15013,N_12919,N_12954);
nor U15014 (N_15014,N_12189,N_13152);
or U15015 (N_15015,N_12089,N_13828);
nor U15016 (N_15016,N_13802,N_12077);
nand U15017 (N_15017,N_12232,N_12298);
nand U15018 (N_15018,N_12095,N_12733);
xor U15019 (N_15019,N_13753,N_12421);
or U15020 (N_15020,N_12348,N_13352);
or U15021 (N_15021,N_12541,N_13657);
or U15022 (N_15022,N_12508,N_12100);
nand U15023 (N_15023,N_12569,N_12783);
nor U15024 (N_15024,N_13664,N_12776);
or U15025 (N_15025,N_12903,N_13206);
nand U15026 (N_15026,N_12807,N_12653);
and U15027 (N_15027,N_13428,N_12601);
or U15028 (N_15028,N_12175,N_13789);
nor U15029 (N_15029,N_13484,N_13554);
nor U15030 (N_15030,N_13702,N_12359);
xnor U15031 (N_15031,N_13837,N_12798);
nor U15032 (N_15032,N_12823,N_13833);
or U15033 (N_15033,N_12397,N_12907);
nand U15034 (N_15034,N_13790,N_13884);
nand U15035 (N_15035,N_12938,N_12884);
nor U15036 (N_15036,N_13955,N_12588);
nand U15037 (N_15037,N_12943,N_13199);
nor U15038 (N_15038,N_12519,N_12314);
and U15039 (N_15039,N_13863,N_13242);
or U15040 (N_15040,N_12620,N_12903);
nand U15041 (N_15041,N_12366,N_13535);
or U15042 (N_15042,N_12585,N_13963);
and U15043 (N_15043,N_13250,N_12224);
xor U15044 (N_15044,N_12041,N_13996);
nand U15045 (N_15045,N_12045,N_12970);
xnor U15046 (N_15046,N_12702,N_12787);
or U15047 (N_15047,N_13956,N_12624);
nor U15048 (N_15048,N_13534,N_13548);
nand U15049 (N_15049,N_13316,N_13364);
nand U15050 (N_15050,N_13414,N_12662);
nor U15051 (N_15051,N_13482,N_13718);
xnor U15052 (N_15052,N_13785,N_13489);
and U15053 (N_15053,N_12165,N_13963);
nand U15054 (N_15054,N_12890,N_12970);
nand U15055 (N_15055,N_12429,N_13783);
nand U15056 (N_15056,N_13249,N_13233);
nand U15057 (N_15057,N_12442,N_12925);
and U15058 (N_15058,N_12672,N_12090);
nor U15059 (N_15059,N_12594,N_13258);
or U15060 (N_15060,N_13227,N_13779);
nand U15061 (N_15061,N_12818,N_12810);
and U15062 (N_15062,N_13577,N_13526);
and U15063 (N_15063,N_12053,N_13469);
or U15064 (N_15064,N_13496,N_13637);
nand U15065 (N_15065,N_13936,N_13619);
and U15066 (N_15066,N_13136,N_13875);
nor U15067 (N_15067,N_12361,N_12107);
nand U15068 (N_15068,N_13156,N_13650);
and U15069 (N_15069,N_13481,N_12310);
xnor U15070 (N_15070,N_12643,N_13368);
or U15071 (N_15071,N_13327,N_12229);
or U15072 (N_15072,N_13083,N_13840);
nor U15073 (N_15073,N_12700,N_13543);
and U15074 (N_15074,N_12344,N_12884);
xor U15075 (N_15075,N_12511,N_13788);
nor U15076 (N_15076,N_13701,N_13067);
or U15077 (N_15077,N_13297,N_13400);
nor U15078 (N_15078,N_13293,N_13250);
xnor U15079 (N_15079,N_12378,N_13590);
nor U15080 (N_15080,N_13006,N_12144);
or U15081 (N_15081,N_13737,N_12129);
or U15082 (N_15082,N_13769,N_12968);
and U15083 (N_15083,N_12550,N_13791);
or U15084 (N_15084,N_13050,N_13383);
nor U15085 (N_15085,N_13949,N_12089);
and U15086 (N_15086,N_12271,N_13916);
and U15087 (N_15087,N_12917,N_12259);
nor U15088 (N_15088,N_12306,N_13542);
xor U15089 (N_15089,N_12655,N_13492);
nor U15090 (N_15090,N_13704,N_13891);
nand U15091 (N_15091,N_12820,N_13976);
nor U15092 (N_15092,N_12518,N_13580);
nand U15093 (N_15093,N_12260,N_13697);
nor U15094 (N_15094,N_13346,N_12194);
or U15095 (N_15095,N_12546,N_13785);
nand U15096 (N_15096,N_12443,N_12357);
and U15097 (N_15097,N_13614,N_13700);
and U15098 (N_15098,N_12734,N_13310);
or U15099 (N_15099,N_13488,N_13743);
and U15100 (N_15100,N_12794,N_12375);
nand U15101 (N_15101,N_13255,N_13544);
xnor U15102 (N_15102,N_13386,N_13445);
nor U15103 (N_15103,N_13582,N_13525);
nor U15104 (N_15104,N_13830,N_13819);
or U15105 (N_15105,N_12696,N_13790);
nand U15106 (N_15106,N_13482,N_12463);
or U15107 (N_15107,N_13525,N_12792);
nand U15108 (N_15108,N_12867,N_13310);
and U15109 (N_15109,N_12865,N_13273);
and U15110 (N_15110,N_13580,N_12726);
and U15111 (N_15111,N_13623,N_12616);
or U15112 (N_15112,N_13802,N_12931);
nor U15113 (N_15113,N_13678,N_13006);
and U15114 (N_15114,N_12152,N_12621);
or U15115 (N_15115,N_13672,N_13133);
nand U15116 (N_15116,N_12232,N_12320);
nor U15117 (N_15117,N_12335,N_12742);
nor U15118 (N_15118,N_12089,N_12384);
nor U15119 (N_15119,N_13197,N_13564);
and U15120 (N_15120,N_12931,N_12492);
nand U15121 (N_15121,N_13952,N_13023);
or U15122 (N_15122,N_13881,N_12296);
nor U15123 (N_15123,N_13980,N_13067);
nor U15124 (N_15124,N_13072,N_12765);
and U15125 (N_15125,N_13788,N_13874);
and U15126 (N_15126,N_13912,N_12464);
nor U15127 (N_15127,N_13179,N_12860);
nand U15128 (N_15128,N_13280,N_12143);
nor U15129 (N_15129,N_12428,N_12123);
nor U15130 (N_15130,N_12953,N_13262);
and U15131 (N_15131,N_13427,N_12567);
nor U15132 (N_15132,N_13070,N_13759);
nor U15133 (N_15133,N_13734,N_12803);
nor U15134 (N_15134,N_12620,N_12777);
or U15135 (N_15135,N_13970,N_13158);
nor U15136 (N_15136,N_12300,N_12864);
and U15137 (N_15137,N_12993,N_13159);
xor U15138 (N_15138,N_13261,N_12494);
and U15139 (N_15139,N_13813,N_12389);
or U15140 (N_15140,N_12037,N_12237);
and U15141 (N_15141,N_12305,N_12328);
nand U15142 (N_15142,N_12929,N_13811);
or U15143 (N_15143,N_12191,N_13985);
xor U15144 (N_15144,N_13306,N_12014);
or U15145 (N_15145,N_12764,N_12985);
or U15146 (N_15146,N_13899,N_12678);
nor U15147 (N_15147,N_13669,N_12260);
xnor U15148 (N_15148,N_12348,N_13181);
nor U15149 (N_15149,N_12837,N_12417);
xor U15150 (N_15150,N_13034,N_12514);
or U15151 (N_15151,N_12613,N_13840);
or U15152 (N_15152,N_12779,N_12316);
nand U15153 (N_15153,N_12775,N_13100);
nor U15154 (N_15154,N_12910,N_12599);
or U15155 (N_15155,N_13667,N_13203);
nor U15156 (N_15156,N_13886,N_13252);
or U15157 (N_15157,N_12810,N_12511);
xor U15158 (N_15158,N_13448,N_13706);
nand U15159 (N_15159,N_13162,N_12192);
nor U15160 (N_15160,N_12790,N_13688);
and U15161 (N_15161,N_12468,N_13680);
or U15162 (N_15162,N_12114,N_12827);
and U15163 (N_15163,N_13283,N_13015);
nand U15164 (N_15164,N_13537,N_12020);
and U15165 (N_15165,N_12478,N_12623);
or U15166 (N_15166,N_12002,N_13806);
and U15167 (N_15167,N_13827,N_12715);
and U15168 (N_15168,N_13916,N_13689);
and U15169 (N_15169,N_12126,N_12501);
nor U15170 (N_15170,N_13459,N_12009);
nor U15171 (N_15171,N_12133,N_13091);
nor U15172 (N_15172,N_12563,N_13054);
nand U15173 (N_15173,N_13463,N_13733);
nand U15174 (N_15174,N_13293,N_13816);
and U15175 (N_15175,N_12284,N_12527);
or U15176 (N_15176,N_13001,N_13133);
and U15177 (N_15177,N_13321,N_12666);
nor U15178 (N_15178,N_13165,N_12769);
nand U15179 (N_15179,N_13233,N_12163);
or U15180 (N_15180,N_12672,N_13643);
and U15181 (N_15181,N_12790,N_13882);
and U15182 (N_15182,N_12523,N_12621);
nor U15183 (N_15183,N_12217,N_13197);
nand U15184 (N_15184,N_12037,N_13815);
nand U15185 (N_15185,N_12415,N_13005);
xor U15186 (N_15186,N_12531,N_12524);
nor U15187 (N_15187,N_13030,N_12704);
or U15188 (N_15188,N_13464,N_12089);
or U15189 (N_15189,N_12457,N_13720);
or U15190 (N_15190,N_13437,N_13007);
and U15191 (N_15191,N_13237,N_12762);
or U15192 (N_15192,N_12015,N_13364);
xnor U15193 (N_15193,N_13995,N_12431);
nor U15194 (N_15194,N_13524,N_13941);
nor U15195 (N_15195,N_12856,N_13188);
nor U15196 (N_15196,N_12699,N_12880);
and U15197 (N_15197,N_12286,N_13810);
nand U15198 (N_15198,N_12006,N_13893);
nand U15199 (N_15199,N_12076,N_13583);
nand U15200 (N_15200,N_13324,N_12142);
and U15201 (N_15201,N_12971,N_12784);
nand U15202 (N_15202,N_13893,N_13008);
nor U15203 (N_15203,N_12795,N_12176);
nor U15204 (N_15204,N_12575,N_13787);
nand U15205 (N_15205,N_12958,N_13265);
nor U15206 (N_15206,N_13651,N_13446);
xor U15207 (N_15207,N_13795,N_12244);
nand U15208 (N_15208,N_12202,N_13162);
or U15209 (N_15209,N_12390,N_12442);
and U15210 (N_15210,N_12059,N_13439);
nor U15211 (N_15211,N_13542,N_13547);
nor U15212 (N_15212,N_12419,N_13438);
nor U15213 (N_15213,N_12765,N_13145);
and U15214 (N_15214,N_13652,N_13481);
and U15215 (N_15215,N_12324,N_12515);
xnor U15216 (N_15216,N_12865,N_12348);
or U15217 (N_15217,N_13630,N_13278);
or U15218 (N_15218,N_12883,N_12372);
and U15219 (N_15219,N_13956,N_13199);
nor U15220 (N_15220,N_13475,N_12034);
nand U15221 (N_15221,N_12016,N_12673);
nor U15222 (N_15222,N_12062,N_12004);
nor U15223 (N_15223,N_12075,N_13236);
and U15224 (N_15224,N_13156,N_12864);
or U15225 (N_15225,N_13218,N_12810);
nand U15226 (N_15226,N_13416,N_13759);
and U15227 (N_15227,N_12085,N_13475);
xor U15228 (N_15228,N_12098,N_12264);
xnor U15229 (N_15229,N_13824,N_12782);
nor U15230 (N_15230,N_12766,N_13461);
nor U15231 (N_15231,N_12367,N_13777);
nand U15232 (N_15232,N_13784,N_12195);
and U15233 (N_15233,N_13030,N_12425);
and U15234 (N_15234,N_12098,N_12632);
nand U15235 (N_15235,N_13853,N_13241);
nor U15236 (N_15236,N_13344,N_12289);
or U15237 (N_15237,N_13573,N_13164);
xnor U15238 (N_15238,N_12472,N_12774);
and U15239 (N_15239,N_12216,N_12467);
nor U15240 (N_15240,N_12870,N_12984);
or U15241 (N_15241,N_12416,N_12659);
and U15242 (N_15242,N_12920,N_13167);
nand U15243 (N_15243,N_12683,N_13562);
or U15244 (N_15244,N_12139,N_12801);
or U15245 (N_15245,N_12052,N_12438);
nand U15246 (N_15246,N_12520,N_12936);
nand U15247 (N_15247,N_12119,N_12752);
and U15248 (N_15248,N_12346,N_13097);
nor U15249 (N_15249,N_12247,N_12396);
or U15250 (N_15250,N_13457,N_13209);
and U15251 (N_15251,N_13873,N_13488);
nand U15252 (N_15252,N_12585,N_12651);
nor U15253 (N_15253,N_13763,N_12840);
nand U15254 (N_15254,N_13734,N_12258);
nand U15255 (N_15255,N_12288,N_12050);
nand U15256 (N_15256,N_13150,N_13245);
or U15257 (N_15257,N_13122,N_13296);
and U15258 (N_15258,N_12976,N_13471);
nand U15259 (N_15259,N_12533,N_12681);
and U15260 (N_15260,N_12334,N_13130);
nor U15261 (N_15261,N_12746,N_13805);
xnor U15262 (N_15262,N_12459,N_13011);
or U15263 (N_15263,N_13239,N_12757);
and U15264 (N_15264,N_12851,N_12887);
nand U15265 (N_15265,N_13372,N_12645);
nand U15266 (N_15266,N_12462,N_12619);
xnor U15267 (N_15267,N_12599,N_13472);
and U15268 (N_15268,N_13118,N_12881);
and U15269 (N_15269,N_13298,N_12257);
xor U15270 (N_15270,N_12107,N_12328);
and U15271 (N_15271,N_12692,N_13646);
and U15272 (N_15272,N_12337,N_13013);
and U15273 (N_15273,N_12080,N_13517);
nand U15274 (N_15274,N_12814,N_13987);
or U15275 (N_15275,N_13569,N_13003);
and U15276 (N_15276,N_13123,N_13890);
nor U15277 (N_15277,N_12992,N_13317);
or U15278 (N_15278,N_13101,N_12431);
xnor U15279 (N_15279,N_13026,N_13144);
nor U15280 (N_15280,N_13183,N_13742);
nand U15281 (N_15281,N_13516,N_12286);
and U15282 (N_15282,N_13737,N_13079);
nor U15283 (N_15283,N_12001,N_12954);
and U15284 (N_15284,N_13894,N_12230);
nand U15285 (N_15285,N_12476,N_13100);
nor U15286 (N_15286,N_13879,N_13487);
nor U15287 (N_15287,N_12592,N_12403);
nand U15288 (N_15288,N_13035,N_12022);
or U15289 (N_15289,N_13208,N_13970);
or U15290 (N_15290,N_12175,N_13042);
nor U15291 (N_15291,N_13050,N_12270);
and U15292 (N_15292,N_12339,N_12835);
or U15293 (N_15293,N_12720,N_13065);
and U15294 (N_15294,N_13035,N_12924);
nor U15295 (N_15295,N_12031,N_12610);
nand U15296 (N_15296,N_13228,N_13507);
nor U15297 (N_15297,N_13548,N_12531);
or U15298 (N_15298,N_13688,N_13463);
or U15299 (N_15299,N_12681,N_12355);
xnor U15300 (N_15300,N_12261,N_13978);
and U15301 (N_15301,N_12891,N_12104);
nand U15302 (N_15302,N_13733,N_13713);
nor U15303 (N_15303,N_12574,N_12911);
and U15304 (N_15304,N_13228,N_12069);
or U15305 (N_15305,N_13864,N_13544);
xor U15306 (N_15306,N_13579,N_13313);
nor U15307 (N_15307,N_12644,N_13836);
and U15308 (N_15308,N_13220,N_12327);
and U15309 (N_15309,N_13313,N_13338);
and U15310 (N_15310,N_12548,N_13972);
nand U15311 (N_15311,N_13638,N_13843);
and U15312 (N_15312,N_12865,N_13271);
nand U15313 (N_15313,N_12043,N_12477);
and U15314 (N_15314,N_13121,N_12511);
or U15315 (N_15315,N_13307,N_13484);
and U15316 (N_15316,N_12008,N_13883);
nand U15317 (N_15317,N_12403,N_13682);
and U15318 (N_15318,N_12324,N_13499);
or U15319 (N_15319,N_13453,N_12220);
nor U15320 (N_15320,N_13195,N_13338);
and U15321 (N_15321,N_13398,N_12292);
or U15322 (N_15322,N_13814,N_12237);
nor U15323 (N_15323,N_13587,N_12823);
or U15324 (N_15324,N_12252,N_12645);
xor U15325 (N_15325,N_13112,N_13108);
or U15326 (N_15326,N_13094,N_13247);
nand U15327 (N_15327,N_13705,N_12268);
and U15328 (N_15328,N_13125,N_12183);
nor U15329 (N_15329,N_12853,N_13150);
nand U15330 (N_15330,N_12535,N_13955);
nand U15331 (N_15331,N_12363,N_12814);
nand U15332 (N_15332,N_13648,N_12213);
nand U15333 (N_15333,N_12321,N_13711);
nand U15334 (N_15334,N_13575,N_12309);
nor U15335 (N_15335,N_13162,N_12129);
nor U15336 (N_15336,N_13340,N_13437);
nand U15337 (N_15337,N_13286,N_13059);
nand U15338 (N_15338,N_12644,N_13001);
and U15339 (N_15339,N_12673,N_13544);
nand U15340 (N_15340,N_13907,N_13951);
xnor U15341 (N_15341,N_12094,N_13188);
nand U15342 (N_15342,N_12598,N_12892);
nor U15343 (N_15343,N_13753,N_12169);
and U15344 (N_15344,N_13842,N_13743);
nor U15345 (N_15345,N_12475,N_12058);
nor U15346 (N_15346,N_12522,N_13612);
or U15347 (N_15347,N_12697,N_13720);
nor U15348 (N_15348,N_12746,N_12984);
xor U15349 (N_15349,N_13751,N_13354);
and U15350 (N_15350,N_13041,N_12125);
nor U15351 (N_15351,N_12225,N_12232);
and U15352 (N_15352,N_12898,N_12017);
and U15353 (N_15353,N_13974,N_12135);
nand U15354 (N_15354,N_12887,N_13635);
and U15355 (N_15355,N_13111,N_13711);
and U15356 (N_15356,N_12404,N_13260);
nor U15357 (N_15357,N_12068,N_13623);
or U15358 (N_15358,N_13202,N_12025);
or U15359 (N_15359,N_12352,N_12018);
and U15360 (N_15360,N_12750,N_13906);
nor U15361 (N_15361,N_12653,N_12457);
or U15362 (N_15362,N_13906,N_13697);
and U15363 (N_15363,N_13013,N_12654);
nand U15364 (N_15364,N_13422,N_13287);
and U15365 (N_15365,N_12103,N_13189);
nor U15366 (N_15366,N_12858,N_12389);
nor U15367 (N_15367,N_12040,N_13659);
nor U15368 (N_15368,N_12296,N_13178);
nor U15369 (N_15369,N_13669,N_13569);
or U15370 (N_15370,N_13752,N_13277);
and U15371 (N_15371,N_13935,N_12893);
nor U15372 (N_15372,N_12580,N_13910);
and U15373 (N_15373,N_12658,N_13066);
or U15374 (N_15374,N_13213,N_13314);
or U15375 (N_15375,N_12006,N_13969);
or U15376 (N_15376,N_13206,N_13022);
nor U15377 (N_15377,N_12741,N_12965);
nor U15378 (N_15378,N_13849,N_12102);
nand U15379 (N_15379,N_13142,N_12706);
nor U15380 (N_15380,N_12783,N_13622);
or U15381 (N_15381,N_13706,N_12167);
nand U15382 (N_15382,N_12552,N_13330);
or U15383 (N_15383,N_12229,N_12939);
and U15384 (N_15384,N_13577,N_13640);
and U15385 (N_15385,N_12269,N_13776);
xor U15386 (N_15386,N_13410,N_12334);
or U15387 (N_15387,N_12765,N_12115);
nor U15388 (N_15388,N_12151,N_13972);
and U15389 (N_15389,N_13548,N_13064);
nand U15390 (N_15390,N_12255,N_12019);
nor U15391 (N_15391,N_13913,N_13325);
or U15392 (N_15392,N_12737,N_12191);
and U15393 (N_15393,N_13326,N_13933);
or U15394 (N_15394,N_12304,N_12295);
and U15395 (N_15395,N_13463,N_12370);
and U15396 (N_15396,N_12044,N_13062);
xor U15397 (N_15397,N_12636,N_12411);
nor U15398 (N_15398,N_13331,N_12892);
nor U15399 (N_15399,N_13352,N_13760);
nand U15400 (N_15400,N_12868,N_12722);
nand U15401 (N_15401,N_13995,N_12553);
xnor U15402 (N_15402,N_13380,N_12648);
nand U15403 (N_15403,N_12368,N_12362);
and U15404 (N_15404,N_13213,N_13293);
nand U15405 (N_15405,N_13849,N_13186);
nand U15406 (N_15406,N_13887,N_13351);
nor U15407 (N_15407,N_12661,N_13117);
xor U15408 (N_15408,N_13943,N_13226);
or U15409 (N_15409,N_12227,N_13149);
nor U15410 (N_15410,N_13678,N_13146);
or U15411 (N_15411,N_12573,N_13197);
nand U15412 (N_15412,N_12126,N_12653);
nor U15413 (N_15413,N_12853,N_12353);
or U15414 (N_15414,N_13869,N_12258);
or U15415 (N_15415,N_13679,N_12262);
or U15416 (N_15416,N_13626,N_12026);
or U15417 (N_15417,N_13251,N_13713);
or U15418 (N_15418,N_12958,N_12626);
nand U15419 (N_15419,N_13419,N_12088);
and U15420 (N_15420,N_13063,N_12074);
or U15421 (N_15421,N_12080,N_12556);
and U15422 (N_15422,N_12466,N_12140);
nand U15423 (N_15423,N_13800,N_13899);
nand U15424 (N_15424,N_12551,N_12143);
and U15425 (N_15425,N_12465,N_12511);
nand U15426 (N_15426,N_12714,N_13190);
or U15427 (N_15427,N_12845,N_13878);
nand U15428 (N_15428,N_13466,N_12183);
nand U15429 (N_15429,N_12397,N_13944);
xnor U15430 (N_15430,N_12956,N_13063);
xnor U15431 (N_15431,N_12328,N_13577);
or U15432 (N_15432,N_12202,N_13992);
and U15433 (N_15433,N_12141,N_13443);
nand U15434 (N_15434,N_12198,N_12804);
nand U15435 (N_15435,N_12699,N_13620);
nand U15436 (N_15436,N_12646,N_12750);
and U15437 (N_15437,N_13801,N_12601);
or U15438 (N_15438,N_12375,N_12180);
nand U15439 (N_15439,N_13773,N_13954);
or U15440 (N_15440,N_12296,N_12811);
and U15441 (N_15441,N_12036,N_13040);
or U15442 (N_15442,N_12108,N_13747);
and U15443 (N_15443,N_12713,N_13965);
and U15444 (N_15444,N_12332,N_12867);
xor U15445 (N_15445,N_13971,N_13139);
or U15446 (N_15446,N_13046,N_13275);
nor U15447 (N_15447,N_13395,N_12144);
and U15448 (N_15448,N_13327,N_13898);
and U15449 (N_15449,N_12343,N_12889);
nor U15450 (N_15450,N_13649,N_12587);
and U15451 (N_15451,N_13969,N_13782);
nand U15452 (N_15452,N_13529,N_13116);
nor U15453 (N_15453,N_12371,N_13092);
and U15454 (N_15454,N_13847,N_13676);
or U15455 (N_15455,N_13759,N_13083);
or U15456 (N_15456,N_12381,N_13813);
and U15457 (N_15457,N_13537,N_12599);
or U15458 (N_15458,N_13204,N_12213);
nand U15459 (N_15459,N_12211,N_13548);
and U15460 (N_15460,N_12641,N_12446);
and U15461 (N_15461,N_12660,N_13637);
nor U15462 (N_15462,N_12536,N_13292);
xnor U15463 (N_15463,N_13461,N_13957);
nor U15464 (N_15464,N_13041,N_13235);
or U15465 (N_15465,N_12828,N_13778);
xor U15466 (N_15466,N_12357,N_12568);
or U15467 (N_15467,N_12714,N_12964);
nand U15468 (N_15468,N_12425,N_13886);
and U15469 (N_15469,N_13798,N_13482);
or U15470 (N_15470,N_12127,N_13267);
xnor U15471 (N_15471,N_13516,N_12034);
nor U15472 (N_15472,N_12108,N_13525);
and U15473 (N_15473,N_12935,N_13556);
nand U15474 (N_15474,N_12471,N_12710);
and U15475 (N_15475,N_12806,N_13368);
nand U15476 (N_15476,N_13609,N_13938);
xnor U15477 (N_15477,N_13118,N_12254);
nand U15478 (N_15478,N_12389,N_13126);
nor U15479 (N_15479,N_12441,N_12687);
and U15480 (N_15480,N_13202,N_12641);
and U15481 (N_15481,N_13101,N_13535);
nand U15482 (N_15482,N_12657,N_12903);
nand U15483 (N_15483,N_12480,N_12865);
xor U15484 (N_15484,N_13958,N_13425);
nand U15485 (N_15485,N_12380,N_12702);
xnor U15486 (N_15486,N_13199,N_12211);
or U15487 (N_15487,N_12623,N_13956);
xor U15488 (N_15488,N_13804,N_13149);
or U15489 (N_15489,N_13647,N_13615);
xor U15490 (N_15490,N_12753,N_12717);
nor U15491 (N_15491,N_12524,N_13975);
and U15492 (N_15492,N_13968,N_13954);
nor U15493 (N_15493,N_13821,N_12799);
or U15494 (N_15494,N_13339,N_12108);
and U15495 (N_15495,N_13551,N_13186);
and U15496 (N_15496,N_12788,N_13659);
xnor U15497 (N_15497,N_13900,N_12366);
and U15498 (N_15498,N_12407,N_12943);
or U15499 (N_15499,N_12664,N_12193);
and U15500 (N_15500,N_12286,N_13712);
nand U15501 (N_15501,N_12984,N_13389);
nor U15502 (N_15502,N_13334,N_12658);
or U15503 (N_15503,N_13229,N_12542);
nor U15504 (N_15504,N_13458,N_12823);
xnor U15505 (N_15505,N_13102,N_13874);
nor U15506 (N_15506,N_12198,N_12384);
and U15507 (N_15507,N_12399,N_12741);
and U15508 (N_15508,N_13903,N_12213);
nand U15509 (N_15509,N_12324,N_13542);
nor U15510 (N_15510,N_12326,N_13795);
nor U15511 (N_15511,N_13693,N_13505);
and U15512 (N_15512,N_12206,N_13627);
or U15513 (N_15513,N_13867,N_13301);
and U15514 (N_15514,N_13746,N_13273);
and U15515 (N_15515,N_13225,N_13660);
nor U15516 (N_15516,N_13429,N_12887);
or U15517 (N_15517,N_12596,N_13843);
and U15518 (N_15518,N_12175,N_12742);
xor U15519 (N_15519,N_12640,N_13077);
nor U15520 (N_15520,N_12917,N_12415);
or U15521 (N_15521,N_13009,N_12979);
and U15522 (N_15522,N_13590,N_13213);
nor U15523 (N_15523,N_12607,N_12569);
and U15524 (N_15524,N_12153,N_12080);
nand U15525 (N_15525,N_13883,N_13636);
or U15526 (N_15526,N_12464,N_12523);
or U15527 (N_15527,N_12644,N_13330);
or U15528 (N_15528,N_13997,N_13197);
xnor U15529 (N_15529,N_12738,N_13490);
nand U15530 (N_15530,N_12566,N_13875);
nand U15531 (N_15531,N_13785,N_13881);
xor U15532 (N_15532,N_13018,N_13637);
xor U15533 (N_15533,N_13674,N_13694);
or U15534 (N_15534,N_13497,N_13548);
and U15535 (N_15535,N_13474,N_13646);
and U15536 (N_15536,N_12528,N_12057);
and U15537 (N_15537,N_13759,N_13708);
and U15538 (N_15538,N_12150,N_12609);
or U15539 (N_15539,N_13595,N_13541);
nand U15540 (N_15540,N_13838,N_12204);
nor U15541 (N_15541,N_13217,N_12847);
and U15542 (N_15542,N_12371,N_12097);
xor U15543 (N_15543,N_13106,N_13371);
nand U15544 (N_15544,N_13116,N_13136);
nor U15545 (N_15545,N_12017,N_12597);
and U15546 (N_15546,N_12785,N_12661);
nor U15547 (N_15547,N_13226,N_13095);
and U15548 (N_15548,N_12907,N_12492);
nor U15549 (N_15549,N_12222,N_13759);
nor U15550 (N_15550,N_13164,N_12975);
xnor U15551 (N_15551,N_12435,N_13350);
xor U15552 (N_15552,N_13451,N_12801);
xor U15553 (N_15553,N_12595,N_13839);
nand U15554 (N_15554,N_12653,N_12570);
nor U15555 (N_15555,N_13092,N_12148);
or U15556 (N_15556,N_13280,N_12992);
nor U15557 (N_15557,N_12633,N_12099);
or U15558 (N_15558,N_13872,N_13099);
and U15559 (N_15559,N_13825,N_12648);
and U15560 (N_15560,N_13684,N_12342);
and U15561 (N_15561,N_13275,N_12793);
nand U15562 (N_15562,N_12286,N_12468);
nand U15563 (N_15563,N_13741,N_13294);
and U15564 (N_15564,N_13645,N_12133);
nand U15565 (N_15565,N_12892,N_13297);
nand U15566 (N_15566,N_13107,N_12713);
nor U15567 (N_15567,N_13264,N_12495);
or U15568 (N_15568,N_13891,N_13195);
and U15569 (N_15569,N_13635,N_13368);
nand U15570 (N_15570,N_13170,N_13413);
or U15571 (N_15571,N_13420,N_12623);
nand U15572 (N_15572,N_12564,N_12382);
and U15573 (N_15573,N_13134,N_13155);
nand U15574 (N_15574,N_13200,N_12522);
and U15575 (N_15575,N_12933,N_12342);
nor U15576 (N_15576,N_12940,N_12653);
nor U15577 (N_15577,N_12055,N_13638);
nand U15578 (N_15578,N_13368,N_13406);
xnor U15579 (N_15579,N_13900,N_13555);
nor U15580 (N_15580,N_12462,N_13211);
nor U15581 (N_15581,N_12520,N_12530);
nand U15582 (N_15582,N_13391,N_12149);
or U15583 (N_15583,N_13737,N_13485);
and U15584 (N_15584,N_12588,N_13539);
or U15585 (N_15585,N_12309,N_12336);
nand U15586 (N_15586,N_13752,N_13693);
xor U15587 (N_15587,N_13892,N_13261);
nand U15588 (N_15588,N_12962,N_13684);
and U15589 (N_15589,N_13819,N_12558);
and U15590 (N_15590,N_12770,N_13109);
xor U15591 (N_15591,N_13566,N_12809);
nor U15592 (N_15592,N_12652,N_13748);
nor U15593 (N_15593,N_12590,N_13570);
and U15594 (N_15594,N_12377,N_12067);
and U15595 (N_15595,N_12923,N_12130);
nor U15596 (N_15596,N_12177,N_13152);
or U15597 (N_15597,N_12568,N_13020);
nand U15598 (N_15598,N_13115,N_12320);
nand U15599 (N_15599,N_13346,N_12667);
or U15600 (N_15600,N_13266,N_13115);
nand U15601 (N_15601,N_13569,N_13558);
or U15602 (N_15602,N_12717,N_12462);
nor U15603 (N_15603,N_12774,N_12952);
xor U15604 (N_15604,N_13048,N_13062);
and U15605 (N_15605,N_13361,N_13425);
nor U15606 (N_15606,N_13915,N_13911);
or U15607 (N_15607,N_12271,N_13370);
or U15608 (N_15608,N_12572,N_13857);
xnor U15609 (N_15609,N_12337,N_13858);
nor U15610 (N_15610,N_12438,N_12379);
or U15611 (N_15611,N_13644,N_13403);
or U15612 (N_15612,N_13820,N_13954);
and U15613 (N_15613,N_13422,N_12183);
nor U15614 (N_15614,N_12960,N_12172);
nand U15615 (N_15615,N_12071,N_12920);
and U15616 (N_15616,N_13311,N_13950);
or U15617 (N_15617,N_12496,N_13325);
and U15618 (N_15618,N_12032,N_13653);
or U15619 (N_15619,N_13465,N_12785);
nand U15620 (N_15620,N_12574,N_12676);
nand U15621 (N_15621,N_12842,N_12680);
and U15622 (N_15622,N_12101,N_13305);
or U15623 (N_15623,N_12687,N_12403);
and U15624 (N_15624,N_12906,N_12202);
and U15625 (N_15625,N_13603,N_13572);
and U15626 (N_15626,N_13466,N_13662);
nor U15627 (N_15627,N_13128,N_12808);
nor U15628 (N_15628,N_12318,N_12928);
or U15629 (N_15629,N_12290,N_12862);
nor U15630 (N_15630,N_13607,N_12769);
or U15631 (N_15631,N_13387,N_13138);
xor U15632 (N_15632,N_12401,N_12858);
or U15633 (N_15633,N_12340,N_13800);
nand U15634 (N_15634,N_13672,N_13516);
or U15635 (N_15635,N_12491,N_13913);
or U15636 (N_15636,N_13476,N_13539);
nor U15637 (N_15637,N_13969,N_12632);
xor U15638 (N_15638,N_12621,N_12317);
and U15639 (N_15639,N_12040,N_12431);
or U15640 (N_15640,N_13456,N_12769);
nand U15641 (N_15641,N_12845,N_12260);
nand U15642 (N_15642,N_12370,N_12875);
and U15643 (N_15643,N_12113,N_13114);
nand U15644 (N_15644,N_13023,N_13274);
xor U15645 (N_15645,N_12854,N_13312);
nor U15646 (N_15646,N_12186,N_13590);
nor U15647 (N_15647,N_13969,N_12112);
nor U15648 (N_15648,N_12082,N_12475);
and U15649 (N_15649,N_12556,N_12447);
or U15650 (N_15650,N_13211,N_13866);
or U15651 (N_15651,N_12425,N_12164);
nor U15652 (N_15652,N_13872,N_12736);
and U15653 (N_15653,N_13387,N_13185);
or U15654 (N_15654,N_12481,N_12236);
and U15655 (N_15655,N_12123,N_12595);
nand U15656 (N_15656,N_12953,N_13875);
nand U15657 (N_15657,N_13164,N_12929);
nor U15658 (N_15658,N_12000,N_13684);
and U15659 (N_15659,N_12304,N_13492);
xor U15660 (N_15660,N_13170,N_12186);
and U15661 (N_15661,N_13128,N_12973);
nand U15662 (N_15662,N_12160,N_12584);
or U15663 (N_15663,N_13845,N_13604);
and U15664 (N_15664,N_12724,N_13316);
and U15665 (N_15665,N_12573,N_12984);
nand U15666 (N_15666,N_12016,N_13806);
and U15667 (N_15667,N_12496,N_12744);
nor U15668 (N_15668,N_12099,N_12536);
nand U15669 (N_15669,N_13328,N_12370);
and U15670 (N_15670,N_12426,N_13082);
or U15671 (N_15671,N_12071,N_12309);
or U15672 (N_15672,N_13109,N_13657);
and U15673 (N_15673,N_13534,N_12100);
nand U15674 (N_15674,N_12124,N_13196);
nand U15675 (N_15675,N_12577,N_13388);
or U15676 (N_15676,N_13198,N_13964);
xnor U15677 (N_15677,N_12982,N_12940);
nand U15678 (N_15678,N_13185,N_12439);
nand U15679 (N_15679,N_12658,N_13657);
nor U15680 (N_15680,N_13186,N_12295);
and U15681 (N_15681,N_12326,N_12510);
or U15682 (N_15682,N_12659,N_13015);
nand U15683 (N_15683,N_12163,N_12897);
nor U15684 (N_15684,N_13858,N_12036);
xor U15685 (N_15685,N_12961,N_12172);
nand U15686 (N_15686,N_13053,N_12411);
and U15687 (N_15687,N_12118,N_12778);
or U15688 (N_15688,N_13719,N_13618);
nand U15689 (N_15689,N_13344,N_12351);
or U15690 (N_15690,N_12159,N_12484);
and U15691 (N_15691,N_13810,N_13265);
and U15692 (N_15692,N_12359,N_13087);
and U15693 (N_15693,N_13443,N_12831);
nor U15694 (N_15694,N_12998,N_13016);
nand U15695 (N_15695,N_12442,N_13244);
nor U15696 (N_15696,N_13359,N_13979);
or U15697 (N_15697,N_13753,N_13756);
nand U15698 (N_15698,N_12102,N_12326);
or U15699 (N_15699,N_13272,N_13201);
xnor U15700 (N_15700,N_13337,N_12413);
nor U15701 (N_15701,N_12048,N_13705);
and U15702 (N_15702,N_13116,N_12895);
and U15703 (N_15703,N_12186,N_13285);
nor U15704 (N_15704,N_13041,N_13276);
nand U15705 (N_15705,N_12153,N_12301);
nand U15706 (N_15706,N_13796,N_13825);
nor U15707 (N_15707,N_12873,N_13327);
or U15708 (N_15708,N_13336,N_13000);
and U15709 (N_15709,N_12678,N_12844);
or U15710 (N_15710,N_12034,N_13830);
and U15711 (N_15711,N_13459,N_13849);
xnor U15712 (N_15712,N_13788,N_13082);
xnor U15713 (N_15713,N_13521,N_12259);
and U15714 (N_15714,N_12611,N_13860);
and U15715 (N_15715,N_13821,N_12526);
nand U15716 (N_15716,N_13994,N_13528);
nand U15717 (N_15717,N_13460,N_12069);
or U15718 (N_15718,N_12921,N_12493);
nand U15719 (N_15719,N_12763,N_13670);
and U15720 (N_15720,N_13595,N_12501);
and U15721 (N_15721,N_13774,N_12205);
xor U15722 (N_15722,N_13111,N_13184);
nand U15723 (N_15723,N_13954,N_13740);
xor U15724 (N_15724,N_12016,N_12203);
xor U15725 (N_15725,N_13498,N_13594);
and U15726 (N_15726,N_13341,N_13308);
and U15727 (N_15727,N_13819,N_13809);
nand U15728 (N_15728,N_12087,N_13623);
nor U15729 (N_15729,N_12984,N_12553);
and U15730 (N_15730,N_12146,N_12722);
or U15731 (N_15731,N_13200,N_12642);
or U15732 (N_15732,N_13818,N_12087);
or U15733 (N_15733,N_13726,N_13890);
nand U15734 (N_15734,N_13933,N_12650);
and U15735 (N_15735,N_12247,N_12626);
and U15736 (N_15736,N_13328,N_12093);
or U15737 (N_15737,N_12059,N_13645);
nand U15738 (N_15738,N_12910,N_12590);
or U15739 (N_15739,N_12720,N_12565);
and U15740 (N_15740,N_12838,N_13472);
and U15741 (N_15741,N_12114,N_13969);
and U15742 (N_15742,N_13388,N_12497);
or U15743 (N_15743,N_13173,N_12750);
xor U15744 (N_15744,N_12068,N_13919);
nand U15745 (N_15745,N_12412,N_12984);
nand U15746 (N_15746,N_12480,N_13702);
and U15747 (N_15747,N_12014,N_13799);
or U15748 (N_15748,N_13692,N_13254);
nand U15749 (N_15749,N_12870,N_13335);
nand U15750 (N_15750,N_12328,N_12651);
and U15751 (N_15751,N_12371,N_12720);
xor U15752 (N_15752,N_12255,N_13241);
or U15753 (N_15753,N_12854,N_13110);
nor U15754 (N_15754,N_12732,N_12361);
nor U15755 (N_15755,N_12848,N_12222);
and U15756 (N_15756,N_13266,N_12061);
and U15757 (N_15757,N_13597,N_13347);
or U15758 (N_15758,N_12327,N_13704);
nand U15759 (N_15759,N_12888,N_13636);
or U15760 (N_15760,N_13650,N_13782);
or U15761 (N_15761,N_13645,N_12461);
nor U15762 (N_15762,N_12312,N_12151);
or U15763 (N_15763,N_13775,N_12204);
nand U15764 (N_15764,N_13975,N_12353);
nor U15765 (N_15765,N_13503,N_13665);
or U15766 (N_15766,N_13902,N_12143);
nor U15767 (N_15767,N_13233,N_12311);
nand U15768 (N_15768,N_13360,N_12820);
nand U15769 (N_15769,N_12905,N_13940);
nor U15770 (N_15770,N_13283,N_12877);
and U15771 (N_15771,N_13677,N_12356);
and U15772 (N_15772,N_13515,N_12525);
nand U15773 (N_15773,N_13696,N_12268);
or U15774 (N_15774,N_13819,N_12028);
xor U15775 (N_15775,N_12667,N_13229);
or U15776 (N_15776,N_12283,N_13968);
or U15777 (N_15777,N_13456,N_13286);
and U15778 (N_15778,N_13608,N_12818);
xnor U15779 (N_15779,N_13026,N_12265);
and U15780 (N_15780,N_13933,N_13552);
nand U15781 (N_15781,N_13142,N_12341);
nand U15782 (N_15782,N_13496,N_12927);
or U15783 (N_15783,N_13771,N_13043);
nand U15784 (N_15784,N_12841,N_12485);
and U15785 (N_15785,N_13659,N_12360);
and U15786 (N_15786,N_13541,N_13959);
or U15787 (N_15787,N_12656,N_12047);
nor U15788 (N_15788,N_12194,N_12662);
nor U15789 (N_15789,N_13670,N_13717);
and U15790 (N_15790,N_13735,N_13240);
and U15791 (N_15791,N_12311,N_12659);
or U15792 (N_15792,N_12478,N_12043);
nor U15793 (N_15793,N_12645,N_12927);
and U15794 (N_15794,N_12087,N_13867);
or U15795 (N_15795,N_13597,N_13791);
nand U15796 (N_15796,N_13138,N_12894);
nand U15797 (N_15797,N_12800,N_12792);
or U15798 (N_15798,N_13338,N_13328);
nor U15799 (N_15799,N_13264,N_13374);
and U15800 (N_15800,N_12030,N_12948);
and U15801 (N_15801,N_12827,N_12954);
nand U15802 (N_15802,N_12831,N_13545);
nand U15803 (N_15803,N_13640,N_13035);
or U15804 (N_15804,N_13974,N_12945);
and U15805 (N_15805,N_12908,N_13150);
nand U15806 (N_15806,N_13281,N_12458);
xnor U15807 (N_15807,N_12081,N_13231);
xor U15808 (N_15808,N_12304,N_13651);
nand U15809 (N_15809,N_13662,N_12132);
nand U15810 (N_15810,N_13724,N_13288);
or U15811 (N_15811,N_12707,N_12288);
nand U15812 (N_15812,N_12208,N_13042);
nand U15813 (N_15813,N_13038,N_13163);
xor U15814 (N_15814,N_13021,N_12494);
nor U15815 (N_15815,N_12020,N_13499);
nand U15816 (N_15816,N_13637,N_12966);
xor U15817 (N_15817,N_13255,N_12237);
xor U15818 (N_15818,N_13731,N_12366);
nor U15819 (N_15819,N_13894,N_13764);
and U15820 (N_15820,N_13879,N_12879);
or U15821 (N_15821,N_12039,N_13330);
nor U15822 (N_15822,N_13762,N_12451);
nand U15823 (N_15823,N_12766,N_13093);
or U15824 (N_15824,N_12350,N_13242);
or U15825 (N_15825,N_12312,N_12947);
nor U15826 (N_15826,N_13585,N_13638);
nor U15827 (N_15827,N_12447,N_12175);
xor U15828 (N_15828,N_13716,N_13954);
nand U15829 (N_15829,N_13488,N_12099);
nor U15830 (N_15830,N_12272,N_12198);
nand U15831 (N_15831,N_13289,N_13670);
nor U15832 (N_15832,N_13785,N_12582);
and U15833 (N_15833,N_13603,N_13626);
or U15834 (N_15834,N_13532,N_12075);
or U15835 (N_15835,N_13987,N_13698);
nor U15836 (N_15836,N_12611,N_13259);
or U15837 (N_15837,N_13059,N_12615);
nor U15838 (N_15838,N_12053,N_13228);
and U15839 (N_15839,N_13914,N_12345);
nand U15840 (N_15840,N_12460,N_13285);
nor U15841 (N_15841,N_12535,N_13016);
or U15842 (N_15842,N_12285,N_13909);
nand U15843 (N_15843,N_13184,N_13823);
xor U15844 (N_15844,N_13988,N_12672);
and U15845 (N_15845,N_12231,N_13957);
xor U15846 (N_15846,N_12901,N_13727);
nand U15847 (N_15847,N_12552,N_13187);
nand U15848 (N_15848,N_13724,N_13315);
xor U15849 (N_15849,N_12205,N_12257);
or U15850 (N_15850,N_13764,N_13612);
xnor U15851 (N_15851,N_13644,N_12484);
and U15852 (N_15852,N_13959,N_13690);
or U15853 (N_15853,N_12819,N_13331);
nor U15854 (N_15854,N_13320,N_13582);
or U15855 (N_15855,N_13535,N_12405);
nor U15856 (N_15856,N_12977,N_13351);
xnor U15857 (N_15857,N_13090,N_12453);
or U15858 (N_15858,N_13949,N_12676);
nand U15859 (N_15859,N_13236,N_12346);
nor U15860 (N_15860,N_12388,N_12247);
or U15861 (N_15861,N_13294,N_13166);
or U15862 (N_15862,N_13480,N_13493);
nor U15863 (N_15863,N_13924,N_13103);
and U15864 (N_15864,N_13081,N_13944);
xnor U15865 (N_15865,N_12751,N_13980);
or U15866 (N_15866,N_13296,N_12538);
xnor U15867 (N_15867,N_12958,N_12627);
nor U15868 (N_15868,N_12343,N_13255);
and U15869 (N_15869,N_12950,N_12454);
or U15870 (N_15870,N_12715,N_12205);
nor U15871 (N_15871,N_13149,N_13898);
xor U15872 (N_15872,N_12877,N_13493);
xnor U15873 (N_15873,N_12107,N_13209);
xor U15874 (N_15874,N_12788,N_12300);
or U15875 (N_15875,N_12992,N_12761);
xor U15876 (N_15876,N_12658,N_13518);
or U15877 (N_15877,N_12899,N_13019);
nand U15878 (N_15878,N_13652,N_12209);
xor U15879 (N_15879,N_12118,N_13908);
nor U15880 (N_15880,N_13195,N_13403);
and U15881 (N_15881,N_13118,N_13716);
nand U15882 (N_15882,N_13351,N_13592);
or U15883 (N_15883,N_12259,N_12814);
or U15884 (N_15884,N_13134,N_12169);
and U15885 (N_15885,N_12284,N_12653);
nand U15886 (N_15886,N_12623,N_12527);
nor U15887 (N_15887,N_12260,N_13115);
and U15888 (N_15888,N_13298,N_12271);
and U15889 (N_15889,N_12560,N_13904);
nand U15890 (N_15890,N_12218,N_13523);
xor U15891 (N_15891,N_12866,N_13109);
or U15892 (N_15892,N_13353,N_13293);
nor U15893 (N_15893,N_13332,N_13108);
or U15894 (N_15894,N_13144,N_12351);
xnor U15895 (N_15895,N_13476,N_12209);
nor U15896 (N_15896,N_12571,N_13034);
nor U15897 (N_15897,N_13123,N_13803);
and U15898 (N_15898,N_13639,N_13086);
nand U15899 (N_15899,N_13586,N_12113);
and U15900 (N_15900,N_12699,N_13575);
and U15901 (N_15901,N_13265,N_13352);
nor U15902 (N_15902,N_13153,N_13466);
and U15903 (N_15903,N_12537,N_12818);
nand U15904 (N_15904,N_13127,N_12608);
and U15905 (N_15905,N_12389,N_13521);
or U15906 (N_15906,N_13166,N_13563);
nand U15907 (N_15907,N_13702,N_13894);
nor U15908 (N_15908,N_13783,N_12598);
and U15909 (N_15909,N_12855,N_12753);
and U15910 (N_15910,N_13142,N_13695);
or U15911 (N_15911,N_12548,N_13124);
nand U15912 (N_15912,N_12017,N_12775);
or U15913 (N_15913,N_12565,N_13210);
xnor U15914 (N_15914,N_12424,N_12842);
and U15915 (N_15915,N_12342,N_12955);
nand U15916 (N_15916,N_13045,N_13569);
or U15917 (N_15917,N_12405,N_13549);
xnor U15918 (N_15918,N_12535,N_13279);
nand U15919 (N_15919,N_12681,N_12836);
or U15920 (N_15920,N_13563,N_13320);
or U15921 (N_15921,N_12488,N_12744);
or U15922 (N_15922,N_12149,N_12597);
nand U15923 (N_15923,N_13683,N_12499);
nor U15924 (N_15924,N_13540,N_13867);
or U15925 (N_15925,N_12783,N_12171);
or U15926 (N_15926,N_12689,N_13864);
nand U15927 (N_15927,N_13991,N_12387);
and U15928 (N_15928,N_12539,N_13901);
nand U15929 (N_15929,N_13670,N_13666);
and U15930 (N_15930,N_13791,N_12775);
xnor U15931 (N_15931,N_12260,N_13456);
or U15932 (N_15932,N_13114,N_12324);
nor U15933 (N_15933,N_13019,N_13070);
or U15934 (N_15934,N_13186,N_12060);
or U15935 (N_15935,N_12343,N_12389);
nor U15936 (N_15936,N_13040,N_12102);
nor U15937 (N_15937,N_13552,N_13376);
xnor U15938 (N_15938,N_13084,N_12968);
or U15939 (N_15939,N_12670,N_13225);
or U15940 (N_15940,N_13550,N_13811);
xnor U15941 (N_15941,N_12320,N_12310);
or U15942 (N_15942,N_13505,N_12725);
or U15943 (N_15943,N_12239,N_13041);
or U15944 (N_15944,N_13579,N_12748);
or U15945 (N_15945,N_13785,N_13842);
xnor U15946 (N_15946,N_13453,N_12560);
and U15947 (N_15947,N_13725,N_12022);
or U15948 (N_15948,N_13280,N_12389);
xor U15949 (N_15949,N_13042,N_12174);
or U15950 (N_15950,N_13758,N_12798);
or U15951 (N_15951,N_13572,N_12726);
or U15952 (N_15952,N_12673,N_12973);
nand U15953 (N_15953,N_12608,N_13283);
or U15954 (N_15954,N_12924,N_12357);
and U15955 (N_15955,N_13044,N_13370);
or U15956 (N_15956,N_13159,N_12755);
xor U15957 (N_15957,N_13519,N_12241);
nand U15958 (N_15958,N_12985,N_13992);
nand U15959 (N_15959,N_13640,N_13610);
nand U15960 (N_15960,N_13069,N_12082);
and U15961 (N_15961,N_13359,N_12519);
xnor U15962 (N_15962,N_13490,N_13565);
nand U15963 (N_15963,N_13124,N_13200);
or U15964 (N_15964,N_13392,N_13608);
nor U15965 (N_15965,N_13249,N_12712);
nor U15966 (N_15966,N_13234,N_13274);
or U15967 (N_15967,N_13243,N_12270);
or U15968 (N_15968,N_13573,N_13558);
and U15969 (N_15969,N_13760,N_12940);
and U15970 (N_15970,N_13227,N_12529);
nor U15971 (N_15971,N_12916,N_12080);
nand U15972 (N_15972,N_12622,N_12464);
xnor U15973 (N_15973,N_12385,N_13041);
nand U15974 (N_15974,N_12790,N_12907);
or U15975 (N_15975,N_12978,N_12317);
or U15976 (N_15976,N_12798,N_12206);
or U15977 (N_15977,N_13395,N_12470);
and U15978 (N_15978,N_13666,N_12390);
or U15979 (N_15979,N_13927,N_13609);
nand U15980 (N_15980,N_13519,N_13443);
and U15981 (N_15981,N_13557,N_12371);
nand U15982 (N_15982,N_13167,N_12777);
or U15983 (N_15983,N_12440,N_12882);
or U15984 (N_15984,N_12937,N_12073);
and U15985 (N_15985,N_12314,N_12370);
or U15986 (N_15986,N_13807,N_13496);
nand U15987 (N_15987,N_12025,N_12016);
and U15988 (N_15988,N_12280,N_12219);
and U15989 (N_15989,N_13252,N_12446);
or U15990 (N_15990,N_13344,N_12158);
nand U15991 (N_15991,N_12951,N_13286);
nand U15992 (N_15992,N_13835,N_13907);
and U15993 (N_15993,N_12186,N_13582);
nand U15994 (N_15994,N_13688,N_13022);
and U15995 (N_15995,N_12387,N_12038);
and U15996 (N_15996,N_12898,N_12974);
nand U15997 (N_15997,N_12026,N_13749);
nand U15998 (N_15998,N_13768,N_13742);
nor U15999 (N_15999,N_12120,N_12448);
and U16000 (N_16000,N_14616,N_15754);
nor U16001 (N_16001,N_14354,N_14974);
and U16002 (N_16002,N_14217,N_14803);
nor U16003 (N_16003,N_15716,N_14006);
and U16004 (N_16004,N_14174,N_15484);
nand U16005 (N_16005,N_15791,N_14847);
or U16006 (N_16006,N_14129,N_14558);
or U16007 (N_16007,N_14885,N_14482);
or U16008 (N_16008,N_14066,N_14267);
nand U16009 (N_16009,N_14492,N_15919);
xnor U16010 (N_16010,N_15102,N_14117);
xnor U16011 (N_16011,N_15275,N_15011);
or U16012 (N_16012,N_14528,N_14125);
and U16013 (N_16013,N_14569,N_14346);
and U16014 (N_16014,N_15836,N_15849);
or U16015 (N_16015,N_15835,N_14464);
nor U16016 (N_16016,N_15580,N_15493);
nand U16017 (N_16017,N_14008,N_15370);
and U16018 (N_16018,N_14199,N_15680);
xnor U16019 (N_16019,N_15342,N_14962);
nor U16020 (N_16020,N_15780,N_15413);
nor U16021 (N_16021,N_14868,N_15952);
nor U16022 (N_16022,N_15734,N_14817);
and U16023 (N_16023,N_15550,N_15447);
nand U16024 (N_16024,N_14138,N_15776);
and U16025 (N_16025,N_14251,N_14243);
xor U16026 (N_16026,N_14925,N_15705);
nand U16027 (N_16027,N_14115,N_14619);
and U16028 (N_16028,N_14203,N_15647);
or U16029 (N_16029,N_14358,N_14990);
xnor U16030 (N_16030,N_15984,N_15203);
nor U16031 (N_16031,N_15278,N_14854);
or U16032 (N_16032,N_14047,N_14696);
nor U16033 (N_16033,N_14542,N_14357);
or U16034 (N_16034,N_15380,N_14554);
or U16035 (N_16035,N_14336,N_15172);
and U16036 (N_16036,N_14015,N_15093);
nand U16037 (N_16037,N_15824,N_14525);
xor U16038 (N_16038,N_15440,N_15329);
nor U16039 (N_16039,N_15988,N_15477);
nand U16040 (N_16040,N_15527,N_14802);
or U16041 (N_16041,N_14794,N_15910);
nor U16042 (N_16042,N_14595,N_14845);
and U16043 (N_16043,N_14750,N_14036);
or U16044 (N_16044,N_15639,N_14074);
nand U16045 (N_16045,N_15389,N_14530);
nor U16046 (N_16046,N_14213,N_14252);
and U16047 (N_16047,N_14122,N_15348);
and U16048 (N_16048,N_15872,N_14145);
xnor U16049 (N_16049,N_15686,N_14055);
or U16050 (N_16050,N_15977,N_15608);
and U16051 (N_16051,N_14037,N_15973);
or U16052 (N_16052,N_14475,N_15135);
nand U16053 (N_16053,N_15251,N_15596);
nor U16054 (N_16054,N_15597,N_14276);
nand U16055 (N_16055,N_14620,N_14501);
nor U16056 (N_16056,N_14488,N_14083);
nand U16057 (N_16057,N_14773,N_15526);
or U16058 (N_16058,N_14721,N_14818);
nand U16059 (N_16059,N_15212,N_14812);
nand U16060 (N_16060,N_14449,N_15291);
xnor U16061 (N_16061,N_15163,N_15523);
nand U16062 (N_16062,N_15843,N_15844);
and U16063 (N_16063,N_14720,N_15373);
or U16064 (N_16064,N_14978,N_14755);
and U16065 (N_16065,N_15941,N_15092);
and U16066 (N_16066,N_14127,N_15558);
and U16067 (N_16067,N_14333,N_14472);
or U16068 (N_16068,N_15006,N_14255);
xor U16069 (N_16069,N_15226,N_15012);
or U16070 (N_16070,N_14386,N_15954);
or U16071 (N_16071,N_14997,N_15248);
or U16072 (N_16072,N_14577,N_15846);
nand U16073 (N_16073,N_15213,N_15360);
xor U16074 (N_16074,N_15677,N_14702);
or U16075 (N_16075,N_15332,N_14426);
nand U16076 (N_16076,N_15086,N_15967);
nand U16077 (N_16077,N_15584,N_14284);
or U16078 (N_16078,N_14096,N_14949);
or U16079 (N_16079,N_14784,N_14939);
and U16080 (N_16080,N_14335,N_14261);
or U16081 (N_16081,N_14685,N_14470);
nor U16082 (N_16082,N_14069,N_14305);
or U16083 (N_16083,N_15416,N_14900);
xnor U16084 (N_16084,N_14988,N_14653);
nand U16085 (N_16085,N_14581,N_15082);
xor U16086 (N_16086,N_15581,N_14937);
and U16087 (N_16087,N_14564,N_14474);
nor U16088 (N_16088,N_14423,N_15729);
nand U16089 (N_16089,N_15191,N_14591);
or U16090 (N_16090,N_14486,N_14436);
nand U16091 (N_16091,N_14932,N_14979);
nand U16092 (N_16092,N_15839,N_14376);
nor U16093 (N_16093,N_14409,N_15299);
nor U16094 (N_16094,N_15888,N_14231);
or U16095 (N_16095,N_14296,N_15271);
and U16096 (N_16096,N_14337,N_15217);
nand U16097 (N_16097,N_15439,N_15870);
xor U16098 (N_16098,N_14571,N_15150);
and U16099 (N_16099,N_15946,N_15508);
nor U16100 (N_16100,N_15475,N_14146);
nand U16101 (N_16101,N_15821,N_14807);
and U16102 (N_16102,N_15205,N_15145);
or U16103 (N_16103,N_14038,N_14902);
and U16104 (N_16104,N_14529,N_15438);
nor U16105 (N_16105,N_14016,N_14930);
xnor U16106 (N_16106,N_15805,N_15820);
and U16107 (N_16107,N_14730,N_15784);
nand U16108 (N_16108,N_14250,N_15346);
and U16109 (N_16109,N_14945,N_15173);
or U16110 (N_16110,N_15797,N_15551);
xnor U16111 (N_16111,N_15790,N_15985);
nor U16112 (N_16112,N_14662,N_14809);
nor U16113 (N_16113,N_15991,N_14921);
and U16114 (N_16114,N_15769,N_15909);
xnor U16115 (N_16115,N_14167,N_14188);
xor U16116 (N_16116,N_15316,N_14084);
nand U16117 (N_16117,N_15147,N_14090);
xnor U16118 (N_16118,N_15867,N_15625);
nand U16119 (N_16119,N_15615,N_15325);
xnor U16120 (N_16120,N_14227,N_14447);
or U16121 (N_16121,N_14873,N_14981);
or U16122 (N_16122,N_15617,N_15982);
or U16123 (N_16123,N_15502,N_14442);
or U16124 (N_16124,N_14947,N_15353);
nor U16125 (N_16125,N_15386,N_15607);
and U16126 (N_16126,N_14642,N_15043);
or U16127 (N_16127,N_15133,N_14164);
nor U16128 (N_16128,N_15243,N_15959);
or U16129 (N_16129,N_14003,N_15005);
or U16130 (N_16130,N_14288,N_15732);
nand U16131 (N_16131,N_14406,N_14839);
nand U16132 (N_16132,N_15727,N_15045);
or U16133 (N_16133,N_14832,N_14030);
or U16134 (N_16134,N_15013,N_15265);
nand U16135 (N_16135,N_14814,N_15307);
xor U16136 (N_16136,N_15337,N_15047);
nand U16137 (N_16137,N_15968,N_15363);
or U16138 (N_16138,N_15741,N_14029);
xnor U16139 (N_16139,N_15823,N_15130);
xnor U16140 (N_16140,N_15219,N_14630);
nor U16141 (N_16141,N_14293,N_14269);
or U16142 (N_16142,N_14883,N_15423);
or U16143 (N_16143,N_15588,N_14104);
nor U16144 (N_16144,N_14633,N_15852);
xor U16145 (N_16145,N_15932,N_15736);
xor U16146 (N_16146,N_14739,N_14858);
or U16147 (N_16147,N_15218,N_15454);
nand U16148 (N_16148,N_15533,N_14441);
nand U16149 (N_16149,N_15328,N_15041);
nor U16150 (N_16150,N_14212,N_14260);
and U16151 (N_16151,N_14189,N_14095);
nor U16152 (N_16152,N_14867,N_14957);
and U16153 (N_16153,N_15281,N_14065);
and U16154 (N_16154,N_15379,N_15886);
and U16155 (N_16155,N_14737,N_14229);
nand U16156 (N_16156,N_14326,N_15300);
and U16157 (N_16157,N_14140,N_15992);
nor U16158 (N_16158,N_15890,N_14209);
and U16159 (N_16159,N_15490,N_14905);
and U16160 (N_16160,N_14157,N_15951);
nor U16161 (N_16161,N_14300,N_15312);
nor U16162 (N_16162,N_15055,N_14823);
or U16163 (N_16163,N_14070,N_14332);
nor U16164 (N_16164,N_15787,N_14808);
nor U16165 (N_16165,N_14454,N_15322);
nand U16166 (N_16166,N_14109,N_14225);
nor U16167 (N_16167,N_15514,N_14621);
and U16168 (N_16168,N_15488,N_15960);
xnor U16169 (N_16169,N_15557,N_15189);
nand U16170 (N_16170,N_15916,N_15906);
and U16171 (N_16171,N_15883,N_14600);
nand U16172 (N_16172,N_14214,N_15878);
or U16173 (N_16173,N_14859,N_15063);
or U16174 (N_16174,N_15088,N_15031);
and U16175 (N_16175,N_14113,N_14909);
nor U16176 (N_16176,N_15225,N_15998);
or U16177 (N_16177,N_15297,N_14215);
and U16178 (N_16178,N_15943,N_15552);
xor U16179 (N_16179,N_14513,N_15602);
nor U16180 (N_16180,N_15320,N_14594);
nor U16181 (N_16181,N_14926,N_15507);
nand U16182 (N_16182,N_14718,N_14013);
and U16183 (N_16183,N_14100,N_15080);
nand U16184 (N_16184,N_15192,N_15200);
xnor U16185 (N_16185,N_14646,N_14541);
nand U16186 (N_16186,N_15465,N_15476);
nor U16187 (N_16187,N_15532,N_14636);
xnor U16188 (N_16188,N_15623,N_14353);
nor U16189 (N_16189,N_15813,N_14399);
or U16190 (N_16190,N_15216,N_14674);
or U16191 (N_16191,N_15873,N_15594);
nand U16192 (N_16192,N_14712,N_14461);
and U16193 (N_16193,N_14548,N_15249);
xnor U16194 (N_16194,N_15270,N_15864);
and U16195 (N_16195,N_15343,N_14230);
xor U16196 (N_16196,N_14366,N_15350);
and U16197 (N_16197,N_15518,N_15953);
and U16198 (N_16198,N_15091,N_15897);
nor U16199 (N_16199,N_14890,N_15035);
nor U16200 (N_16200,N_15310,N_14537);
and U16201 (N_16201,N_14891,N_15289);
nor U16202 (N_16202,N_15175,N_14428);
nand U16203 (N_16203,N_14610,N_15381);
and U16204 (N_16204,N_15800,N_15355);
xor U16205 (N_16205,N_14079,N_14405);
and U16206 (N_16206,N_14310,N_15905);
and U16207 (N_16207,N_15482,N_15802);
or U16208 (N_16208,N_15728,N_14012);
nand U16209 (N_16209,N_14745,N_15692);
nor U16210 (N_16210,N_14018,N_14330);
and U16211 (N_16211,N_15298,N_14843);
or U16212 (N_16212,N_14747,N_15649);
nand U16213 (N_16213,N_15364,N_14913);
nand U16214 (N_16214,N_14343,N_14311);
and U16215 (N_16215,N_14879,N_15609);
nor U16216 (N_16216,N_15450,N_15485);
or U16217 (N_16217,N_15395,N_14958);
or U16218 (N_16218,N_14815,N_15923);
or U16219 (N_16219,N_14093,N_14158);
nor U16220 (N_16220,N_14322,N_14959);
xor U16221 (N_16221,N_14089,N_14897);
or U16222 (N_16222,N_14289,N_15230);
or U16223 (N_16223,N_15929,N_15573);
nand U16224 (N_16224,N_14190,N_15947);
and U16225 (N_16225,N_14738,N_15881);
nor U16226 (N_16226,N_15798,N_15255);
or U16227 (N_16227,N_15614,N_14384);
or U16228 (N_16228,N_15981,N_15109);
nand U16229 (N_16229,N_14994,N_14453);
nand U16230 (N_16230,N_14235,N_14272);
nor U16231 (N_16231,N_14292,N_15834);
nor U16232 (N_16232,N_14221,N_15900);
and U16233 (N_16233,N_15713,N_14224);
or U16234 (N_16234,N_14657,N_15566);
nand U16235 (N_16235,N_14800,N_15308);
nor U16236 (N_16236,N_14050,N_14911);
or U16237 (N_16237,N_14906,N_14848);
nor U16238 (N_16238,N_14368,N_15687);
or U16239 (N_16239,N_14506,N_15865);
and U16240 (N_16240,N_14220,N_15100);
nor U16241 (N_16241,N_14306,N_14114);
xnor U16242 (N_16242,N_15453,N_15809);
and U16243 (N_16243,N_15869,N_14950);
nand U16244 (N_16244,N_15948,N_14105);
and U16245 (N_16245,N_14075,N_14560);
nor U16246 (N_16246,N_14363,N_15315);
or U16247 (N_16247,N_15574,N_14816);
xor U16248 (N_16248,N_15585,N_15717);
nand U16249 (N_16249,N_15252,N_14451);
and U16250 (N_16250,N_15361,N_15085);
nand U16251 (N_16251,N_15165,N_14236);
or U16252 (N_16252,N_15633,N_14044);
nand U16253 (N_16253,N_14367,N_14473);
nor U16254 (N_16254,N_15975,N_15345);
nor U16255 (N_16255,N_15026,N_15643);
or U16256 (N_16256,N_14836,N_15096);
xnor U16257 (N_16257,N_15724,N_14103);
nand U16258 (N_16258,N_15666,N_15903);
and U16259 (N_16259,N_15496,N_14732);
nand U16260 (N_16260,N_14054,N_15851);
nor U16261 (N_16261,N_15449,N_14497);
and U16262 (N_16262,N_14121,N_15876);
nor U16263 (N_16263,N_14187,N_15369);
nand U16264 (N_16264,N_15338,N_15668);
nor U16265 (N_16265,N_14341,N_14304);
nor U16266 (N_16266,N_14924,N_15101);
nor U16267 (N_16267,N_15994,N_14724);
and U16268 (N_16268,N_15928,N_14578);
nand U16269 (N_16269,N_15704,N_14345);
or U16270 (N_16270,N_14896,N_14680);
nor U16271 (N_16271,N_14223,N_14785);
and U16272 (N_16272,N_15700,N_14362);
nor U16273 (N_16273,N_14118,N_14494);
and U16274 (N_16274,N_14379,N_14675);
nand U16275 (N_16275,N_15044,N_14862);
or U16276 (N_16276,N_14101,N_15725);
nor U16277 (N_16277,N_15187,N_15256);
and U16278 (N_16278,N_15356,N_14186);
or U16279 (N_16279,N_15286,N_14419);
xor U16280 (N_16280,N_14234,N_14299);
nor U16281 (N_16281,N_14701,N_15319);
nand U16282 (N_16282,N_15738,N_14694);
nand U16283 (N_16283,N_14489,N_14881);
or U16284 (N_16284,N_15164,N_14788);
nand U16285 (N_16285,N_15061,N_14589);
nor U16286 (N_16286,N_15153,N_15521);
and U16287 (N_16287,N_14850,N_14643);
nor U16288 (N_16288,N_14603,N_15742);
nor U16289 (N_16289,N_14071,N_15323);
nand U16290 (N_16290,N_15682,N_15415);
and U16291 (N_16291,N_15140,N_15000);
xor U16292 (N_16292,N_15891,N_15658);
nor U16293 (N_16293,N_14351,N_15431);
and U16294 (N_16294,N_14647,N_15534);
nor U16295 (N_16295,N_15481,N_14328);
or U16296 (N_16296,N_15253,N_14758);
and U16297 (N_16297,N_14584,N_15371);
and U16298 (N_16298,N_14886,N_15194);
nand U16299 (N_16299,N_15313,N_15987);
or U16300 (N_16300,N_15193,N_14045);
nor U16301 (N_16301,N_15448,N_15616);
nand U16302 (N_16302,N_14205,N_15749);
xnor U16303 (N_16303,N_14699,N_15944);
or U16304 (N_16304,N_14964,N_15254);
nor U16305 (N_16305,N_15889,N_15422);
or U16306 (N_16306,N_14705,N_15758);
nor U16307 (N_16307,N_15083,N_14064);
and U16308 (N_16308,N_15801,N_14601);
nand U16309 (N_16309,N_14178,N_14842);
or U16310 (N_16310,N_14431,N_14731);
xnor U16311 (N_16311,N_14557,N_14391);
nor U16312 (N_16312,N_15103,N_15577);
nand U16313 (N_16313,N_15160,N_15884);
nand U16314 (N_16314,N_14144,N_15123);
nand U16315 (N_16315,N_14496,N_15040);
or U16316 (N_16316,N_15284,N_15620);
and U16317 (N_16317,N_14752,N_14700);
and U16318 (N_16318,N_14659,N_15050);
nor U16319 (N_16319,N_15238,N_15917);
and U16320 (N_16320,N_14182,N_14028);
nor U16321 (N_16321,N_15408,N_14727);
and U16322 (N_16322,N_15858,N_14632);
nand U16323 (N_16323,N_14435,N_14155);
and U16324 (N_16324,N_14264,N_15779);
and U16325 (N_16325,N_15376,N_14347);
nand U16326 (N_16326,N_15304,N_15010);
or U16327 (N_16327,N_14938,N_14796);
nand U16328 (N_16328,N_14606,N_14573);
nor U16329 (N_16329,N_14534,N_14500);
and U16330 (N_16330,N_14654,N_15246);
nand U16331 (N_16331,N_14767,N_15007);
and U16332 (N_16332,N_14108,N_14927);
and U16333 (N_16333,N_15171,N_14042);
nand U16334 (N_16334,N_15462,N_15277);
nand U16335 (N_16335,N_15087,N_14546);
nor U16336 (N_16336,N_15303,N_15764);
and U16337 (N_16337,N_14691,N_15621);
xor U16338 (N_16338,N_14931,N_15979);
nor U16339 (N_16339,N_15186,N_14201);
nand U16340 (N_16340,N_15712,N_14314);
xor U16341 (N_16341,N_15236,N_14671);
or U16342 (N_16342,N_15957,N_14059);
nand U16343 (N_16343,N_14919,N_15520);
nor U16344 (N_16344,N_14869,N_14277);
xnor U16345 (N_16345,N_14370,N_15555);
nor U16346 (N_16346,N_14819,N_14283);
nor U16347 (N_16347,N_15403,N_14057);
nor U16348 (N_16348,N_14545,N_14966);
or U16349 (N_16349,N_15469,N_15997);
xnor U16350 (N_16350,N_14527,N_14786);
nor U16351 (N_16351,N_15174,N_14116);
nor U16352 (N_16352,N_14413,N_14725);
or U16353 (N_16353,N_15333,N_14309);
nand U16354 (N_16354,N_14717,N_14339);
and U16355 (N_16355,N_15511,N_14871);
nor U16356 (N_16356,N_15201,N_14266);
nand U16357 (N_16357,N_15512,N_14198);
nand U16358 (N_16358,N_15519,N_14491);
or U16359 (N_16359,N_15144,N_14572);
nand U16360 (N_16360,N_15377,N_15487);
or U16361 (N_16361,N_15626,N_15018);
or U16362 (N_16362,N_14687,N_15646);
or U16363 (N_16363,N_15719,N_15209);
or U16364 (N_16364,N_14855,N_14445);
or U16365 (N_16365,N_14805,N_14552);
or U16366 (N_16366,N_14373,N_15847);
or U16367 (N_16367,N_15405,N_14485);
xnor U16368 (N_16368,N_15108,N_14723);
nand U16369 (N_16369,N_14736,N_14661);
and U16370 (N_16370,N_14387,N_15019);
nand U16371 (N_16371,N_15073,N_15781);
and U16372 (N_16372,N_15875,N_14320);
nor U16373 (N_16373,N_14953,N_14519);
nand U16374 (N_16374,N_14644,N_14318);
and U16375 (N_16375,N_14137,N_15927);
or U16376 (N_16376,N_15782,N_15258);
nand U16377 (N_16377,N_14888,N_15460);
and U16378 (N_16378,N_15024,N_14826);
nand U16379 (N_16379,N_15842,N_15458);
and U16380 (N_16380,N_15950,N_15848);
or U16381 (N_16381,N_15904,N_15359);
and U16382 (N_16382,N_15095,N_14682);
nor U16383 (N_16383,N_14237,N_15115);
or U16384 (N_16384,N_14514,N_14033);
or U16385 (N_16385,N_15179,N_14627);
nor U16386 (N_16386,N_15015,N_14171);
xor U16387 (N_16387,N_15470,N_15400);
and U16388 (N_16388,N_15134,N_14658);
nor U16389 (N_16389,N_15136,N_14798);
and U16390 (N_16390,N_14998,N_15444);
or U16391 (N_16391,N_15401,N_15962);
nand U16392 (N_16392,N_15028,N_14141);
and U16393 (N_16393,N_14995,N_14996);
nor U16394 (N_16394,N_14392,N_15601);
nand U16395 (N_16395,N_15675,N_15168);
or U16396 (N_16396,N_14110,N_15283);
or U16397 (N_16397,N_14751,N_15651);
nor U16398 (N_16398,N_15606,N_15435);
and U16399 (N_16399,N_14588,N_14004);
nor U16400 (N_16400,N_15089,N_15358);
and U16401 (N_16401,N_14835,N_14286);
or U16402 (N_16402,N_15335,N_15034);
xor U16403 (N_16403,N_14863,N_14211);
nor U16404 (N_16404,N_15750,N_15180);
or U16405 (N_16405,N_15622,N_15722);
and U16406 (N_16406,N_15344,N_14099);
nor U16407 (N_16407,N_15806,N_15156);
and U16408 (N_16408,N_14856,N_14463);
nand U16409 (N_16409,N_15016,N_14550);
nand U16410 (N_16410,N_14946,N_15743);
nor U16411 (N_16411,N_14400,N_15279);
and U16412 (N_16412,N_14761,N_15306);
or U16413 (N_16413,N_14077,N_15056);
nor U16414 (N_16414,N_14087,N_14510);
and U16415 (N_16415,N_15397,N_14143);
and U16416 (N_16416,N_15197,N_14348);
and U16417 (N_16417,N_15190,N_15425);
and U16418 (N_16418,N_15427,N_15907);
xor U16419 (N_16419,N_15372,N_14692);
or U16420 (N_16420,N_15042,N_15816);
nor U16421 (N_16421,N_15263,N_15911);
nor U16422 (N_16422,N_14393,N_15861);
or U16423 (N_16423,N_15378,N_15081);
nor U16424 (N_16424,N_14793,N_14973);
and U16425 (N_16425,N_15268,N_15347);
xnor U16426 (N_16426,N_15457,N_15826);
nor U16427 (N_16427,N_14324,N_15114);
xor U16428 (N_16428,N_14574,N_15819);
and U16429 (N_16429,N_15778,N_15763);
or U16430 (N_16430,N_15681,N_15652);
and U16431 (N_16431,N_15783,N_14698);
nor U16432 (N_16432,N_14418,N_15983);
nand U16433 (N_16433,N_14424,N_14583);
and U16434 (N_16434,N_14303,N_14714);
nand U16435 (N_16435,N_14512,N_15463);
nand U16436 (N_16436,N_14350,N_14285);
nor U16437 (N_16437,N_14302,N_15468);
xor U16438 (N_16438,N_14663,N_14416);
nor U16439 (N_16439,N_14648,N_14618);
nand U16440 (N_16440,N_14163,N_15498);
nand U16441 (N_16441,N_14982,N_15543);
nand U16442 (N_16442,N_14360,N_14437);
nor U16443 (N_16443,N_15167,N_14034);
nand U16444 (N_16444,N_14085,N_14968);
nor U16445 (N_16445,N_15336,N_15990);
or U16446 (N_16446,N_14669,N_15935);
nand U16447 (N_16447,N_14408,N_14281);
xor U16448 (N_16448,N_14980,N_15940);
nand U16449 (N_16449,N_14860,N_14617);
and U16450 (N_16450,N_14607,N_15099);
or U16451 (N_16451,N_15365,N_15945);
nand U16452 (N_16452,N_15610,N_14908);
and U16453 (N_16453,N_15961,N_15768);
nand U16454 (N_16454,N_15925,N_15466);
and U16455 (N_16455,N_14895,N_14287);
and U16456 (N_16456,N_14889,N_14342);
nand U16457 (N_16457,N_14520,N_14670);
or U16458 (N_16458,N_15892,N_14238);
xnor U16459 (N_16459,N_15793,N_15837);
nor U16460 (N_16460,N_14443,N_15046);
and U16461 (N_16461,N_15479,N_14719);
xnor U16462 (N_16462,N_14652,N_15424);
xor U16463 (N_16463,N_15036,N_14407);
nor U16464 (N_16464,N_15124,N_15445);
nor U16465 (N_16465,N_14587,N_15544);
nand U16466 (N_16466,N_14076,N_14623);
and U16467 (N_16467,N_14999,N_15301);
or U16468 (N_16468,N_14778,N_14851);
or U16469 (N_16469,N_14273,N_14200);
nand U16470 (N_16470,N_14216,N_15748);
and U16471 (N_16471,N_15321,N_15362);
xnor U16472 (N_16472,N_14726,N_14765);
nand U16473 (N_16473,N_15845,N_14124);
nor U16474 (N_16474,N_14639,N_15565);
nor U16475 (N_16475,N_15659,N_14660);
nor U16476 (N_16476,N_15208,N_15351);
nand U16477 (N_16477,N_14608,N_15942);
and U16478 (N_16478,N_15695,N_14352);
nor U16479 (N_16479,N_15170,N_15474);
nand U16480 (N_16480,N_14315,N_15121);
nand U16481 (N_16481,N_15421,N_14951);
and U16482 (N_16482,N_15214,N_15922);
nor U16483 (N_16483,N_15547,N_14498);
xor U16484 (N_16484,N_15368,N_14060);
or U16485 (N_16485,N_15357,N_15811);
nor U16486 (N_16486,N_15324,N_15472);
or U16487 (N_16487,N_14467,N_15107);
nand U16488 (N_16488,N_14870,N_15676);
nor U16489 (N_16489,N_14063,N_15070);
nor U16490 (N_16490,N_14058,N_14152);
nand U16491 (N_16491,N_14611,N_15505);
nand U16492 (N_16492,N_14983,N_14703);
nand U16493 (N_16493,N_14344,N_14002);
xor U16494 (N_16494,N_14361,N_15582);
nand U16495 (N_16495,N_15603,N_14414);
and U16496 (N_16496,N_15402,N_14954);
nor U16497 (N_16497,N_15866,N_15926);
xor U16498 (N_16498,N_15696,N_14476);
or U16499 (N_16499,N_14041,N_15459);
nand U16500 (N_16500,N_14651,N_15745);
or U16501 (N_16501,N_14177,N_15025);
nand U16502 (N_16502,N_14233,N_15387);
and U16503 (N_16503,N_15760,N_15934);
or U16504 (N_16504,N_14874,N_14676);
nand U16505 (N_16505,N_15915,N_14704);
and U16506 (N_16506,N_15434,N_15517);
xor U16507 (N_16507,N_15292,N_15912);
nor U16508 (N_16508,N_14395,N_14614);
nor U16509 (N_16509,N_15810,N_14555);
nor U16510 (N_16510,N_14148,N_14134);
nor U16511 (N_16511,N_15556,N_14697);
nor U16512 (N_16512,N_15840,N_14774);
and U16513 (N_16513,N_14294,N_15385);
or U16514 (N_16514,N_15827,N_15531);
nor U16515 (N_16515,N_14515,N_14450);
nand U16516 (N_16516,N_14480,N_14120);
or U16517 (N_16517,N_15509,N_14678);
and U16518 (N_16518,N_14410,N_15296);
nand U16519 (N_16519,N_15830,N_14970);
nor U16520 (N_16520,N_15568,N_14323);
and U16521 (N_16521,N_14374,N_15612);
nor U16522 (N_16522,N_15032,N_15720);
or U16523 (N_16523,N_14567,N_14061);
nor U16524 (N_16524,N_14046,N_15037);
or U16525 (N_16525,N_15030,N_14517);
nor U16526 (N_16526,N_15210,N_15288);
and U16527 (N_16527,N_15491,N_15691);
xor U16528 (N_16528,N_14715,N_14649);
and U16529 (N_16529,N_15559,N_15812);
xor U16530 (N_16530,N_15721,N_15525);
nand U16531 (N_16531,N_15318,N_15499);
nor U16532 (N_16532,N_15500,N_14052);
or U16533 (N_16533,N_15349,N_14181);
nand U16534 (N_16534,N_15269,N_14133);
nand U16535 (N_16535,N_15492,N_14729);
nand U16536 (N_16536,N_15125,N_15599);
nor U16537 (N_16537,N_14775,N_14317);
nor U16538 (N_16538,N_15391,N_14955);
nor U16539 (N_16539,N_15241,N_14377);
or U16540 (N_16540,N_14622,N_14420);
xor U16541 (N_16541,N_14629,N_15261);
nor U16542 (N_16542,N_14438,N_15222);
nand U16543 (N_16543,N_14484,N_15414);
or U16544 (N_16544,N_14677,N_15204);
nor U16545 (N_16545,N_14713,N_15267);
nand U16546 (N_16546,N_15117,N_14067);
and U16547 (N_16547,N_14683,N_15250);
nand U16548 (N_16548,N_15151,N_14992);
nand U16549 (N_16549,N_14493,N_15841);
and U16550 (N_16550,N_14032,N_15685);
nand U16551 (N_16551,N_15618,N_14811);
nor U16552 (N_16552,N_14106,N_15570);
nor U16553 (N_16553,N_14505,N_14929);
nor U16554 (N_16554,N_14690,N_15120);
and U16555 (N_16555,N_14433,N_14923);
xnor U16556 (N_16556,N_15966,N_15503);
nor U16557 (N_16557,N_15663,N_14456);
nand U16558 (N_16558,N_14733,N_14638);
xnor U16559 (N_16559,N_14766,N_15767);
or U16560 (N_16560,N_15233,N_15564);
nand U16561 (N_16561,N_15887,N_15964);
or U16562 (N_16562,N_15282,N_14777);
nor U16563 (N_16563,N_15437,N_14961);
nor U16564 (N_16564,N_14204,N_15773);
nand U16565 (N_16565,N_15393,N_15980);
nand U16566 (N_16566,N_15882,N_15650);
xor U16567 (N_16567,N_14760,N_14846);
nand U16568 (N_16568,N_14086,N_14686);
or U16569 (N_16569,N_15228,N_15569);
nand U16570 (N_16570,N_15562,N_15079);
nor U16571 (N_16571,N_14568,N_15902);
xnor U16572 (N_16572,N_14894,N_15317);
and U16573 (N_16573,N_15069,N_14469);
or U16574 (N_16574,N_14605,N_14131);
nand U16575 (N_16575,N_14882,N_15832);
nand U16576 (N_16576,N_15708,N_15772);
xor U16577 (N_16577,N_14176,N_14634);
nor U16578 (N_16578,N_15850,N_14402);
and U16579 (N_16579,N_14389,N_14790);
or U16580 (N_16580,N_14185,N_15074);
and U16581 (N_16581,N_14831,N_14975);
xor U16582 (N_16582,N_14184,N_15879);
or U16583 (N_16583,N_15149,N_15285);
nand U16584 (N_16584,N_15896,N_15075);
nor U16585 (N_16585,N_14985,N_14521);
nand U16586 (N_16586,N_15627,N_15139);
or U16587 (N_16587,N_15038,N_15828);
nand U16588 (N_16588,N_14375,N_15661);
or U16589 (N_16589,N_14080,N_14503);
nor U16590 (N_16590,N_15723,N_14401);
or U16591 (N_16591,N_14355,N_14722);
and U16592 (N_16592,N_15159,N_14772);
and U16593 (N_16593,N_14789,N_14837);
nor U16594 (N_16594,N_15118,N_14340);
or U16595 (N_16595,N_15223,N_14245);
nor U16596 (N_16596,N_15066,N_14740);
nand U16597 (N_16597,N_14532,N_15703);
nand U16598 (N_16598,N_14479,N_15877);
and U16599 (N_16599,N_14385,N_14828);
nand U16600 (N_16600,N_14801,N_14840);
nand U16601 (N_16601,N_15999,N_14708);
or U16602 (N_16602,N_15516,N_15644);
and U16603 (N_16603,N_14904,N_15595);
or U16604 (N_16604,N_14097,N_15058);
and U16605 (N_16605,N_14684,N_15645);
nand U16606 (N_16606,N_15198,N_15451);
nand U16607 (N_16607,N_15662,N_14597);
or U16608 (N_16608,N_14128,N_14928);
nand U16609 (N_16609,N_15656,N_14936);
nand U16610 (N_16610,N_15693,N_14210);
nand U16611 (N_16611,N_14422,N_15112);
or U16612 (N_16612,N_15930,N_15936);
nor U16613 (N_16613,N_15937,N_15394);
nand U16614 (N_16614,N_15489,N_15808);
and U16615 (N_16615,N_15287,N_14716);
nand U16616 (N_16616,N_14609,N_15920);
nor U16617 (N_16617,N_14378,N_14987);
nand U16618 (N_16618,N_15406,N_15195);
nor U16619 (N_16619,N_15965,N_14139);
or U16620 (N_16620,N_14068,N_15589);
and U16621 (N_16621,N_15995,N_15817);
xor U16622 (N_16622,N_15799,N_15077);
or U16623 (N_16623,N_14613,N_15996);
nor U16624 (N_16624,N_14153,N_15057);
nand U16625 (N_16625,N_15127,N_15259);
nand U16626 (N_16626,N_14989,N_14312);
and U16627 (N_16627,N_15726,N_15137);
nor U16628 (N_16628,N_15536,N_14914);
and U16629 (N_16629,N_15684,N_14244);
nor U16630 (N_16630,N_14098,N_15262);
nand U16631 (N_16631,N_15235,N_14556);
nor U16632 (N_16632,N_14147,N_14170);
nand U16633 (N_16633,N_14673,N_15366);
nor U16634 (N_16634,N_15672,N_15632);
nor U16635 (N_16635,N_15611,N_15885);
and U16636 (N_16636,N_15539,N_14960);
nor U16637 (N_16637,N_14681,N_14417);
xor U16638 (N_16638,N_15428,N_14017);
nor U16639 (N_16639,N_15383,N_15382);
nand U16640 (N_16640,N_15648,N_15860);
nand U16641 (N_16641,N_15874,N_14094);
xnor U16642 (N_16642,N_15737,N_14536);
nand U16643 (N_16643,N_15575,N_14693);
or U16644 (N_16644,N_14459,N_15280);
and U16645 (N_16645,N_14265,N_14524);
nor U16646 (N_16646,N_15855,N_14976);
and U16647 (N_16647,N_14645,N_15554);
nand U16648 (N_16648,N_15549,N_14162);
and U16649 (N_16649,N_15631,N_15094);
nor U16650 (N_16650,N_14365,N_14728);
nand U16651 (N_16651,N_15908,N_15613);
or U16652 (N_16652,N_15938,N_15247);
and U16653 (N_16653,N_15796,N_15048);
nand U16654 (N_16654,N_15314,N_14993);
nand U16655 (N_16655,N_14027,N_14969);
nand U16656 (N_16656,N_14637,N_15986);
nand U16657 (N_16657,N_14194,N_15567);
nor U16658 (N_16658,N_15561,N_15829);
and U16659 (N_16659,N_14707,N_15181);
or U16660 (N_16660,N_14844,N_14709);
nor U16661 (N_16661,N_15067,N_14490);
nand U16662 (N_16662,N_14531,N_14258);
or U16663 (N_16663,N_14666,N_14971);
or U16664 (N_16664,N_14448,N_14967);
or U16665 (N_16665,N_15105,N_15237);
xnor U16666 (N_16666,N_15529,N_15642);
nand U16667 (N_16667,N_14746,N_15899);
nand U16668 (N_16668,N_15110,N_14783);
nor U16669 (N_16669,N_14849,N_15143);
nand U16670 (N_16670,N_14540,N_15452);
or U16671 (N_16671,N_14887,N_15515);
nor U16672 (N_16672,N_15326,N_14056);
nand U16673 (N_16673,N_14585,N_15694);
xor U16674 (N_16674,N_15545,N_15412);
nor U16675 (N_16675,N_14757,N_14829);
or U16676 (N_16676,N_14172,N_14313);
nand U16677 (N_16677,N_15478,N_15546);
or U16678 (N_16678,N_14943,N_14465);
nor U16679 (N_16679,N_15240,N_14256);
or U16680 (N_16680,N_15637,N_15029);
nor U16681 (N_16681,N_15524,N_14942);
nand U16682 (N_16682,N_15786,N_14689);
nand U16683 (N_16683,N_14403,N_15868);
xor U16684 (N_16684,N_14197,N_14898);
or U16685 (N_16685,N_14791,N_15062);
nand U16686 (N_16686,N_15775,N_15746);
or U16687 (N_16687,N_15640,N_14561);
and U16688 (N_16688,N_14040,N_14833);
nor U16689 (N_16689,N_14543,N_15939);
and U16690 (N_16690,N_14107,N_14319);
nand U16691 (N_16691,N_14242,N_15211);
nor U16692 (N_16692,N_14159,N_14986);
xnor U16693 (N_16693,N_14329,N_15106);
or U16694 (N_16694,N_14754,N_14460);
nand U16695 (N_16695,N_14667,N_15715);
and U16696 (N_16696,N_15290,N_15017);
xnor U16697 (N_16697,N_15154,N_14102);
nand U16698 (N_16698,N_15753,N_14356);
nor U16699 (N_16699,N_14780,N_15894);
nor U16700 (N_16700,N_14744,N_15098);
nand U16701 (N_16701,N_14741,N_15859);
nand U16702 (N_16702,N_15718,N_14830);
and U16703 (N_16703,N_15302,N_14412);
and U16704 (N_16704,N_14282,N_15711);
and U16705 (N_16705,N_15513,N_14910);
nor U16706 (N_16706,N_14518,N_15804);
nor U16707 (N_16707,N_15417,N_15122);
and U16708 (N_16708,N_15461,N_15956);
and U16709 (N_16709,N_14523,N_15678);
and U16710 (N_16710,N_15506,N_14813);
or U16711 (N_16711,N_15976,N_15730);
nand U16712 (N_16712,N_14544,N_14711);
nor U16713 (N_16713,N_14446,N_15774);
or U16714 (N_16714,N_15548,N_15898);
nor U16715 (N_16715,N_14156,N_15049);
and U16716 (N_16716,N_14135,N_14504);
nand U16717 (N_16717,N_14232,N_15244);
or U16718 (N_16718,N_14776,N_15733);
nand U16719 (N_16719,N_14195,N_15455);
and U16720 (N_16720,N_15004,N_14226);
or U16721 (N_16721,N_14566,N_15969);
nor U16722 (N_16722,N_15785,N_15399);
and U16723 (N_16723,N_15542,N_15535);
or U16724 (N_16724,N_14806,N_14191);
and U16725 (N_16725,N_15600,N_14119);
nand U16726 (N_16726,N_15162,N_15739);
nand U16727 (N_16727,N_15586,N_15051);
nor U16728 (N_16728,N_14820,N_15054);
nand U16729 (N_16729,N_15014,N_14838);
xor U16730 (N_16730,N_15432,N_14380);
and U16731 (N_16731,N_14262,N_14522);
nand U16732 (N_16732,N_15234,N_14877);
or U16733 (N_16733,N_14009,N_15311);
or U16734 (N_16734,N_14246,N_15196);
nor U16735 (N_16735,N_14665,N_15924);
nor U16736 (N_16736,N_14088,N_15053);
nand U16737 (N_16737,N_14248,N_15598);
xor U16738 (N_16738,N_15714,N_15528);
nand U16739 (N_16739,N_15331,N_14136);
and U16740 (N_16740,N_15530,N_14081);
and U16741 (N_16741,N_15392,N_14743);
or U16742 (N_16742,N_15702,N_14656);
xnor U16743 (N_16743,N_14965,N_14834);
nand U16744 (N_16744,N_14321,N_14604);
and U16745 (N_16745,N_15410,N_15119);
xnor U16746 (N_16746,N_14861,N_14948);
or U16747 (N_16747,N_14547,N_14624);
nand U16748 (N_16748,N_14404,N_15949);
or U16749 (N_16749,N_14549,N_15762);
or U16750 (N_16750,N_15111,N_15215);
nor U16751 (N_16751,N_14278,N_15815);
nor U16752 (N_16752,N_14092,N_15657);
or U16753 (N_16753,N_14598,N_15177);
nor U16754 (N_16754,N_14130,N_15022);
nand U16755 (N_16755,N_14468,N_14875);
nand U16756 (N_16756,N_14526,N_14483);
or U16757 (N_16757,N_15002,N_15146);
or U16758 (N_16758,N_14169,N_15456);
nor U16759 (N_16759,N_15653,N_15327);
or U16760 (N_16760,N_14364,N_15305);
and U16761 (N_16761,N_15697,N_15683);
or U16762 (N_16762,N_15390,N_14878);
xor U16763 (N_16763,N_15274,N_15751);
nor U16764 (N_16764,N_14562,N_15264);
or U16765 (N_16765,N_14916,N_14672);
nor U16766 (N_16766,N_15731,N_14415);
nand U16767 (N_16767,N_15814,N_14570);
or U16768 (N_16768,N_14020,N_15128);
nor U16769 (N_16769,N_15673,N_15918);
or U16770 (N_16770,N_15113,N_15199);
or U16771 (N_16771,N_14901,N_15220);
xor U16772 (N_16772,N_14759,N_14021);
nand U16773 (N_16773,N_15132,N_14072);
nor U16774 (N_16774,N_15634,N_15341);
or U16775 (N_16775,N_15538,N_14039);
and U16776 (N_16776,N_15407,N_14275);
nor U16777 (N_16777,N_15522,N_15065);
nor U16778 (N_16778,N_15624,N_14688);
nand U16779 (N_16779,N_14538,N_14779);
and U16780 (N_16780,N_14011,N_15483);
and U16781 (N_16781,N_14565,N_15396);
xnor U16782 (N_16782,N_14756,N_15744);
and U16783 (N_16783,N_15690,N_14586);
or U16784 (N_16784,N_14023,N_14787);
nand U16785 (N_16785,N_14381,N_15667);
xor U16786 (N_16786,N_15334,N_14397);
xnor U16787 (N_16787,N_14533,N_14173);
nand U16788 (N_16788,N_14196,N_14664);
or U16789 (N_16789,N_15021,N_14142);
or U16790 (N_16790,N_14922,N_14308);
and U16791 (N_16791,N_15974,N_14625);
nand U16792 (N_16792,N_14477,N_15404);
or U16793 (N_16793,N_15221,N_15579);
nand U16794 (N_16794,N_15242,N_14179);
nor U16795 (N_16795,N_15831,N_14334);
and U16796 (N_16796,N_14253,N_14612);
and U16797 (N_16797,N_15426,N_15989);
nor U16798 (N_16798,N_15418,N_15818);
nor U16799 (N_16799,N_14035,N_14782);
or U16800 (N_16800,N_15970,N_14301);
and U16801 (N_16801,N_14154,N_15486);
nand U16802 (N_16802,N_14183,N_14762);
or U16803 (N_16803,N_14563,N_15553);
nor U16804 (N_16804,N_14907,N_14241);
nor U16805 (N_16805,N_14753,N_15182);
and U16806 (N_16806,N_15354,N_14165);
and U16807 (N_16807,N_15229,N_14263);
or U16808 (N_16808,N_14825,N_15757);
xor U16809 (N_16809,N_15352,N_15771);
nor U16810 (N_16810,N_14192,N_15803);
nand U16811 (N_16811,N_15188,N_15330);
nand U16812 (N_16812,N_14481,N_14383);
and U16813 (N_16813,N_15504,N_15388);
nand U16814 (N_16814,N_14903,N_14411);
or U16815 (N_16815,N_14439,N_15740);
or U16816 (N_16816,N_15914,N_15429);
nand U16817 (N_16817,N_15068,N_14291);
nor U16818 (N_16818,N_15138,N_14010);
nand U16819 (N_16819,N_14580,N_15071);
nor U16820 (N_16820,N_14427,N_15710);
xor U16821 (N_16821,N_14257,N_15593);
or U16822 (N_16822,N_14274,N_14372);
xor U16823 (N_16823,N_15629,N_14559);
nor U16824 (N_16824,N_15157,N_14429);
and U16825 (N_16825,N_14920,N_14325);
nor U16826 (N_16826,N_15295,N_15591);
xor U16827 (N_16827,N_15895,N_15576);
xor U16828 (N_16828,N_15958,N_15104);
and U16829 (N_16829,N_15155,N_15294);
and U16830 (N_16830,N_14073,N_15224);
or U16831 (N_16831,N_14049,N_15020);
or U16832 (N_16832,N_15563,N_14615);
xor U16833 (N_16833,N_14892,N_15245);
xor U16834 (N_16834,N_14771,N_14022);
nand U16835 (N_16835,N_15166,N_15635);
or U16836 (N_16836,N_15788,N_14599);
and U16837 (N_16837,N_15495,N_14944);
and U16838 (N_16838,N_15059,N_15441);
nand U16839 (N_16839,N_14933,N_14940);
and U16840 (N_16840,N_14749,N_14576);
and U16841 (N_16841,N_14421,N_14748);
nand U16842 (N_16842,N_15755,N_14487);
and U16843 (N_16843,N_15023,N_15972);
nor U16844 (N_16844,N_14952,N_14168);
xnor U16845 (N_16845,N_15792,N_14626);
and U16846 (N_16846,N_14679,N_14602);
or U16847 (N_16847,N_15375,N_15541);
or U16848 (N_16848,N_15232,N_14592);
nand U16849 (N_16849,N_14295,N_15411);
nor U16850 (N_16850,N_14478,N_15862);
nor U16851 (N_16851,N_15178,N_15497);
and U16852 (N_16852,N_14208,N_14280);
or U16853 (N_16853,N_14972,N_14872);
nor U16854 (N_16854,N_15825,N_14180);
nor U16855 (N_16855,N_15467,N_14864);
or U16856 (N_16856,N_15854,N_14371);
nand U16857 (N_16857,N_14382,N_15765);
xor U16858 (N_16858,N_14430,N_15374);
nor U16859 (N_16859,N_14734,N_15913);
or U16860 (N_16860,N_15590,N_14218);
or U16861 (N_16861,N_15674,N_14166);
nor U16862 (N_16862,N_15706,N_15807);
nor U16863 (N_16863,N_14507,N_14051);
and U16864 (N_16864,N_15072,N_14963);
and U16865 (N_16865,N_14768,N_15578);
and U16866 (N_16866,N_14764,N_14466);
nor U16867 (N_16867,N_15756,N_15933);
nand U16868 (N_16868,N_15227,N_14641);
or U16869 (N_16869,N_14628,N_14917);
nand U16870 (N_16870,N_15688,N_15009);
and U16871 (N_16871,N_15893,N_14640);
and U16872 (N_16872,N_15510,N_15398);
nand U16873 (N_16873,N_14509,N_15367);
nand U16874 (N_16874,N_15880,N_14458);
or U16875 (N_16875,N_15231,N_15184);
nand U16876 (N_16876,N_15664,N_14024);
or U16877 (N_16877,N_14338,N_14511);
nor U16878 (N_16878,N_15419,N_14668);
and U16879 (N_16879,N_14781,N_15052);
or U16880 (N_16880,N_15473,N_14579);
and U16881 (N_16881,N_15001,N_15709);
or U16882 (N_16882,N_14123,N_15931);
xnor U16883 (N_16883,N_14452,N_14853);
nor U16884 (N_16884,N_15592,N_14575);
nor U16885 (N_16885,N_15604,N_15097);
or U16886 (N_16886,N_15076,N_15309);
nand U16887 (N_16887,N_15636,N_14582);
or U16888 (N_16888,N_14254,N_14007);
nor U16889 (N_16889,N_14048,N_14001);
and U16890 (N_16890,N_15759,N_14390);
or U16891 (N_16891,N_15587,N_15464);
or U16892 (N_16892,N_15671,N_15039);
nand U16893 (N_16893,N_15206,N_14852);
nor U16894 (N_16894,N_14207,N_15471);
nand U16895 (N_16895,N_14279,N_14956);
or U16896 (N_16896,N_15572,N_14934);
and U16897 (N_16897,N_14991,N_15856);
xor U16898 (N_16898,N_15833,N_14271);
or U16899 (N_16899,N_15148,N_14149);
or U16900 (N_16900,N_14150,N_14297);
and U16901 (N_16901,N_14918,N_15064);
xor U16902 (N_16902,N_14508,N_14865);
and U16903 (N_16903,N_14792,N_14082);
nand U16904 (N_16904,N_15701,N_15084);
and U16905 (N_16905,N_15789,N_15794);
nand U16906 (N_16906,N_15628,N_15630);
nor U16907 (N_16907,N_14298,N_15480);
and U16908 (N_16908,N_14000,N_15239);
nor U16909 (N_16909,N_14349,N_14735);
xnor U16910 (N_16910,N_15443,N_15863);
and U16911 (N_16911,N_14499,N_15183);
nor U16912 (N_16912,N_14935,N_15766);
and U16913 (N_16913,N_14111,N_14495);
and U16914 (N_16914,N_14053,N_14193);
and U16915 (N_16915,N_14327,N_15655);
nor U16916 (N_16916,N_14857,N_14240);
xnor U16917 (N_16917,N_14650,N_14219);
and U16918 (N_16918,N_14804,N_14539);
xnor U16919 (N_16919,N_14596,N_15955);
nand U16920 (N_16920,N_14043,N_15971);
or U16921 (N_16921,N_14175,N_15141);
nor U16922 (N_16922,N_15202,N_14091);
and U16923 (N_16923,N_14899,N_14425);
nor U16924 (N_16924,N_14206,N_15735);
nand U16925 (N_16925,N_14014,N_15857);
nor U16926 (N_16926,N_14866,N_15273);
and U16927 (N_16927,N_14247,N_15339);
or U16928 (N_16928,N_14078,N_14590);
and U16929 (N_16929,N_15078,N_15003);
and U16930 (N_16930,N_15619,N_14290);
and U16931 (N_16931,N_15272,N_14369);
nand U16932 (N_16932,N_15689,N_14884);
nor U16933 (N_16933,N_15660,N_14827);
nand U16934 (N_16934,N_14396,N_15921);
nand U16935 (N_16935,N_15409,N_14388);
or U16936 (N_16936,N_14822,N_15761);
nand U16937 (N_16937,N_15207,N_15654);
nand U16938 (N_16938,N_14593,N_15698);
nor U16939 (N_16939,N_15158,N_14270);
and U16940 (N_16940,N_14706,N_15978);
or U16941 (N_16941,N_14799,N_14797);
nand U16942 (N_16942,N_15670,N_14160);
and U16943 (N_16943,N_14239,N_15560);
xor U16944 (N_16944,N_14880,N_15571);
or U16945 (N_16945,N_15747,N_15822);
nor U16946 (N_16946,N_14062,N_14770);
xor U16947 (N_16947,N_14126,N_15266);
nor U16948 (N_16948,N_15641,N_14394);
and U16949 (N_16949,N_15838,N_14977);
or U16950 (N_16950,N_14893,N_14151);
or U16951 (N_16951,N_14307,N_14795);
and U16952 (N_16952,N_15993,N_15494);
nor U16953 (N_16953,N_14553,N_15770);
nand U16954 (N_16954,N_14005,N_14444);
and U16955 (N_16955,N_14202,N_14941);
and U16956 (N_16956,N_15605,N_14516);
and U16957 (N_16957,N_14268,N_15142);
or U16958 (N_16958,N_14432,N_15257);
nand U16959 (N_16959,N_14398,N_14631);
nand U16960 (N_16960,N_14502,N_15540);
nor U16961 (N_16961,N_15420,N_14535);
nor U16962 (N_16962,N_15795,N_15537);
nor U16963 (N_16963,N_15090,N_14026);
and U16964 (N_16964,N_15777,N_15176);
nor U16965 (N_16965,N_15442,N_14821);
or U16966 (N_16966,N_14455,N_15033);
or U16967 (N_16967,N_14359,N_14161);
or U16968 (N_16968,N_15853,N_14912);
xor U16969 (N_16969,N_14915,N_15901);
or U16970 (N_16970,N_15436,N_15008);
xnor U16971 (N_16971,N_15293,N_15027);
nor U16972 (N_16972,N_14984,N_15384);
or U16973 (N_16973,N_15126,N_15260);
or U16974 (N_16974,N_15707,N_15340);
nor U16975 (N_16975,N_14019,N_14635);
nand U16976 (N_16976,N_14259,N_14331);
and U16977 (N_16977,N_15669,N_14025);
or U16978 (N_16978,N_15129,N_14316);
nor U16979 (N_16979,N_14132,N_15060);
nor U16980 (N_16980,N_14471,N_14434);
and U16981 (N_16981,N_15161,N_15501);
or U16982 (N_16982,N_15583,N_14222);
and U16983 (N_16983,N_15433,N_15963);
or U16984 (N_16984,N_14112,N_14228);
nor U16985 (N_16985,N_15679,N_14440);
nor U16986 (N_16986,N_14031,N_14457);
nand U16987 (N_16987,N_15699,N_14824);
or U16988 (N_16988,N_15276,N_14841);
xor U16989 (N_16989,N_14655,N_15185);
nor U16990 (N_16990,N_14695,N_14769);
or U16991 (N_16991,N_15638,N_15665);
xnor U16992 (N_16992,N_15131,N_14876);
and U16993 (N_16993,N_14249,N_14742);
and U16994 (N_16994,N_15169,N_14551);
or U16995 (N_16995,N_14462,N_15871);
nor U16996 (N_16996,N_14810,N_15752);
and U16997 (N_16997,N_15446,N_15116);
xor U16998 (N_16998,N_14710,N_15430);
nand U16999 (N_16999,N_15152,N_14763);
and U17000 (N_17000,N_14206,N_15657);
or U17001 (N_17001,N_15097,N_14222);
or U17002 (N_17002,N_15981,N_14104);
or U17003 (N_17003,N_14014,N_15771);
and U17004 (N_17004,N_15282,N_15027);
and U17005 (N_17005,N_14542,N_15077);
nand U17006 (N_17006,N_15782,N_15411);
nand U17007 (N_17007,N_14387,N_15900);
or U17008 (N_17008,N_14716,N_15326);
nand U17009 (N_17009,N_14417,N_15034);
or U17010 (N_17010,N_15553,N_14086);
nand U17011 (N_17011,N_14755,N_14954);
xor U17012 (N_17012,N_15241,N_14627);
or U17013 (N_17013,N_14540,N_15934);
and U17014 (N_17014,N_15946,N_15859);
nor U17015 (N_17015,N_14613,N_14934);
or U17016 (N_17016,N_14860,N_14877);
nand U17017 (N_17017,N_14742,N_14478);
and U17018 (N_17018,N_15777,N_15249);
or U17019 (N_17019,N_14971,N_15290);
or U17020 (N_17020,N_14866,N_15494);
xor U17021 (N_17021,N_14316,N_14420);
nor U17022 (N_17022,N_14937,N_14543);
and U17023 (N_17023,N_14418,N_15207);
nand U17024 (N_17024,N_14093,N_14282);
or U17025 (N_17025,N_15560,N_14091);
or U17026 (N_17026,N_15147,N_14091);
nor U17027 (N_17027,N_14499,N_14032);
nand U17028 (N_17028,N_14555,N_14720);
and U17029 (N_17029,N_15143,N_15905);
nor U17030 (N_17030,N_15185,N_15096);
xnor U17031 (N_17031,N_14543,N_15469);
and U17032 (N_17032,N_15420,N_14713);
or U17033 (N_17033,N_15892,N_15124);
or U17034 (N_17034,N_14434,N_15645);
and U17035 (N_17035,N_15380,N_15711);
nor U17036 (N_17036,N_15693,N_14798);
xnor U17037 (N_17037,N_14379,N_15583);
nor U17038 (N_17038,N_14595,N_14603);
and U17039 (N_17039,N_15237,N_14200);
nor U17040 (N_17040,N_14971,N_14386);
or U17041 (N_17041,N_14300,N_14373);
or U17042 (N_17042,N_15287,N_14893);
nor U17043 (N_17043,N_15068,N_15762);
nor U17044 (N_17044,N_14595,N_15328);
and U17045 (N_17045,N_15478,N_14894);
or U17046 (N_17046,N_15913,N_14825);
or U17047 (N_17047,N_14096,N_14600);
or U17048 (N_17048,N_14411,N_14209);
or U17049 (N_17049,N_15997,N_15499);
nand U17050 (N_17050,N_14441,N_14959);
and U17051 (N_17051,N_14682,N_14478);
nor U17052 (N_17052,N_15098,N_14474);
xor U17053 (N_17053,N_14562,N_14950);
nor U17054 (N_17054,N_14368,N_15424);
nor U17055 (N_17055,N_15450,N_15215);
nand U17056 (N_17056,N_14209,N_14824);
and U17057 (N_17057,N_14163,N_15401);
nand U17058 (N_17058,N_15875,N_15017);
or U17059 (N_17059,N_14962,N_14879);
nand U17060 (N_17060,N_15651,N_14890);
and U17061 (N_17061,N_15640,N_14913);
and U17062 (N_17062,N_14384,N_14557);
xnor U17063 (N_17063,N_15354,N_15424);
or U17064 (N_17064,N_15926,N_15067);
and U17065 (N_17065,N_14405,N_14989);
and U17066 (N_17066,N_15235,N_14009);
xnor U17067 (N_17067,N_15945,N_14347);
or U17068 (N_17068,N_15884,N_14590);
and U17069 (N_17069,N_15814,N_15516);
nor U17070 (N_17070,N_15662,N_15714);
nor U17071 (N_17071,N_14315,N_15442);
nor U17072 (N_17072,N_15803,N_14340);
nand U17073 (N_17073,N_15662,N_15548);
nand U17074 (N_17074,N_14757,N_14219);
or U17075 (N_17075,N_15916,N_15386);
xnor U17076 (N_17076,N_15451,N_14147);
nand U17077 (N_17077,N_15216,N_15375);
nand U17078 (N_17078,N_14664,N_14974);
and U17079 (N_17079,N_14698,N_15480);
nor U17080 (N_17080,N_14409,N_14326);
and U17081 (N_17081,N_14165,N_14425);
and U17082 (N_17082,N_14340,N_15019);
and U17083 (N_17083,N_15140,N_15186);
or U17084 (N_17084,N_14900,N_14805);
and U17085 (N_17085,N_15038,N_15490);
nor U17086 (N_17086,N_14893,N_14624);
or U17087 (N_17087,N_15175,N_15886);
nand U17088 (N_17088,N_15728,N_14663);
or U17089 (N_17089,N_15415,N_14783);
nand U17090 (N_17090,N_14567,N_15178);
nand U17091 (N_17091,N_15101,N_14887);
xnor U17092 (N_17092,N_14421,N_15749);
xnor U17093 (N_17093,N_15767,N_14341);
nor U17094 (N_17094,N_14231,N_15681);
and U17095 (N_17095,N_14703,N_15890);
nand U17096 (N_17096,N_15387,N_14182);
or U17097 (N_17097,N_14484,N_14031);
or U17098 (N_17098,N_15485,N_15568);
and U17099 (N_17099,N_15539,N_15296);
nand U17100 (N_17100,N_14977,N_14970);
nor U17101 (N_17101,N_15227,N_15978);
or U17102 (N_17102,N_14634,N_15578);
nand U17103 (N_17103,N_15691,N_14407);
xor U17104 (N_17104,N_15334,N_14363);
or U17105 (N_17105,N_15226,N_14560);
and U17106 (N_17106,N_15365,N_14236);
nor U17107 (N_17107,N_14693,N_14600);
nand U17108 (N_17108,N_15999,N_15136);
nand U17109 (N_17109,N_15606,N_14753);
and U17110 (N_17110,N_14729,N_14851);
and U17111 (N_17111,N_15260,N_15216);
nand U17112 (N_17112,N_15522,N_14848);
or U17113 (N_17113,N_15633,N_14958);
and U17114 (N_17114,N_14148,N_14703);
nor U17115 (N_17115,N_15779,N_14501);
or U17116 (N_17116,N_15604,N_15319);
or U17117 (N_17117,N_14052,N_14108);
and U17118 (N_17118,N_15025,N_14566);
xnor U17119 (N_17119,N_14450,N_15198);
nand U17120 (N_17120,N_15099,N_14394);
nor U17121 (N_17121,N_14055,N_15788);
nor U17122 (N_17122,N_14750,N_14187);
and U17123 (N_17123,N_14405,N_14373);
or U17124 (N_17124,N_15040,N_15475);
and U17125 (N_17125,N_15637,N_15343);
nand U17126 (N_17126,N_14733,N_15655);
nand U17127 (N_17127,N_15765,N_15955);
and U17128 (N_17128,N_15530,N_14042);
and U17129 (N_17129,N_15110,N_15317);
nand U17130 (N_17130,N_15821,N_15939);
nor U17131 (N_17131,N_15640,N_15611);
xor U17132 (N_17132,N_14288,N_15857);
nor U17133 (N_17133,N_14701,N_15311);
nor U17134 (N_17134,N_14197,N_14493);
nand U17135 (N_17135,N_15757,N_14167);
nor U17136 (N_17136,N_14297,N_15774);
nor U17137 (N_17137,N_15662,N_15945);
nand U17138 (N_17138,N_14370,N_14827);
xor U17139 (N_17139,N_14374,N_14372);
and U17140 (N_17140,N_14757,N_15786);
and U17141 (N_17141,N_14508,N_14504);
or U17142 (N_17142,N_14703,N_14270);
and U17143 (N_17143,N_15402,N_14820);
nor U17144 (N_17144,N_14098,N_14024);
or U17145 (N_17145,N_15075,N_15551);
nand U17146 (N_17146,N_15240,N_15201);
nand U17147 (N_17147,N_15381,N_14115);
nor U17148 (N_17148,N_15125,N_15095);
nor U17149 (N_17149,N_15282,N_15658);
xnor U17150 (N_17150,N_14244,N_14950);
nand U17151 (N_17151,N_14379,N_15012);
nand U17152 (N_17152,N_14021,N_15044);
or U17153 (N_17153,N_14880,N_15009);
or U17154 (N_17154,N_15609,N_14643);
xor U17155 (N_17155,N_15327,N_15032);
nor U17156 (N_17156,N_15504,N_15656);
and U17157 (N_17157,N_14141,N_15560);
or U17158 (N_17158,N_14978,N_14048);
or U17159 (N_17159,N_15320,N_14698);
nand U17160 (N_17160,N_15825,N_15383);
and U17161 (N_17161,N_14859,N_15680);
or U17162 (N_17162,N_15395,N_14854);
nand U17163 (N_17163,N_15119,N_15582);
or U17164 (N_17164,N_14580,N_14921);
and U17165 (N_17165,N_14227,N_15011);
nand U17166 (N_17166,N_15226,N_14418);
and U17167 (N_17167,N_15130,N_14736);
xor U17168 (N_17168,N_15407,N_15001);
or U17169 (N_17169,N_14521,N_15602);
or U17170 (N_17170,N_14637,N_14421);
nand U17171 (N_17171,N_15943,N_14381);
or U17172 (N_17172,N_15537,N_14686);
nand U17173 (N_17173,N_14007,N_14391);
nor U17174 (N_17174,N_14851,N_15933);
and U17175 (N_17175,N_14967,N_14705);
xnor U17176 (N_17176,N_14200,N_14796);
nand U17177 (N_17177,N_14696,N_14905);
or U17178 (N_17178,N_15298,N_15572);
nor U17179 (N_17179,N_15739,N_15126);
nand U17180 (N_17180,N_14985,N_15218);
nor U17181 (N_17181,N_15418,N_14640);
nand U17182 (N_17182,N_14747,N_14038);
nor U17183 (N_17183,N_14285,N_14385);
and U17184 (N_17184,N_15716,N_15260);
xor U17185 (N_17185,N_15982,N_14274);
and U17186 (N_17186,N_15755,N_14842);
nand U17187 (N_17187,N_14559,N_15515);
and U17188 (N_17188,N_15950,N_14073);
and U17189 (N_17189,N_15113,N_14247);
nor U17190 (N_17190,N_14252,N_14099);
nor U17191 (N_17191,N_15126,N_15296);
or U17192 (N_17192,N_15558,N_14017);
or U17193 (N_17193,N_14261,N_15803);
nor U17194 (N_17194,N_14627,N_15364);
and U17195 (N_17195,N_14093,N_15484);
nor U17196 (N_17196,N_14104,N_14584);
nor U17197 (N_17197,N_14135,N_15144);
xor U17198 (N_17198,N_14420,N_15138);
xor U17199 (N_17199,N_14844,N_15324);
and U17200 (N_17200,N_15731,N_14337);
or U17201 (N_17201,N_15982,N_15937);
and U17202 (N_17202,N_14530,N_15461);
and U17203 (N_17203,N_15709,N_15274);
nand U17204 (N_17204,N_14462,N_15181);
nor U17205 (N_17205,N_14922,N_15577);
nand U17206 (N_17206,N_15131,N_14145);
nand U17207 (N_17207,N_15010,N_15051);
and U17208 (N_17208,N_15335,N_15205);
xor U17209 (N_17209,N_15441,N_14025);
nor U17210 (N_17210,N_15533,N_14933);
nand U17211 (N_17211,N_14178,N_14512);
nor U17212 (N_17212,N_14649,N_15678);
nand U17213 (N_17213,N_15843,N_14935);
or U17214 (N_17214,N_14677,N_15792);
or U17215 (N_17215,N_15090,N_14259);
and U17216 (N_17216,N_14442,N_14145);
and U17217 (N_17217,N_15747,N_14247);
or U17218 (N_17218,N_14370,N_14377);
or U17219 (N_17219,N_14626,N_14716);
or U17220 (N_17220,N_14289,N_14648);
and U17221 (N_17221,N_15654,N_15492);
nor U17222 (N_17222,N_15762,N_14101);
nand U17223 (N_17223,N_14458,N_14610);
nand U17224 (N_17224,N_14459,N_15252);
xnor U17225 (N_17225,N_14300,N_15876);
or U17226 (N_17226,N_15892,N_15126);
xor U17227 (N_17227,N_14053,N_15317);
or U17228 (N_17228,N_14091,N_14286);
nor U17229 (N_17229,N_15283,N_15228);
and U17230 (N_17230,N_15948,N_14766);
nand U17231 (N_17231,N_15278,N_14031);
and U17232 (N_17232,N_14854,N_14497);
nand U17233 (N_17233,N_14146,N_15131);
nor U17234 (N_17234,N_15991,N_15552);
nor U17235 (N_17235,N_14036,N_15964);
or U17236 (N_17236,N_14832,N_14591);
and U17237 (N_17237,N_15006,N_14682);
and U17238 (N_17238,N_15316,N_15308);
and U17239 (N_17239,N_15914,N_15808);
nand U17240 (N_17240,N_14819,N_14824);
or U17241 (N_17241,N_14930,N_15699);
nor U17242 (N_17242,N_14378,N_15546);
and U17243 (N_17243,N_14737,N_15508);
nor U17244 (N_17244,N_15981,N_14797);
nor U17245 (N_17245,N_15087,N_15754);
xnor U17246 (N_17246,N_15096,N_15383);
or U17247 (N_17247,N_15966,N_15111);
or U17248 (N_17248,N_14607,N_14816);
nand U17249 (N_17249,N_15268,N_15842);
nor U17250 (N_17250,N_14673,N_15598);
xnor U17251 (N_17251,N_15010,N_15982);
or U17252 (N_17252,N_14629,N_14807);
nor U17253 (N_17253,N_14923,N_14009);
nand U17254 (N_17254,N_15173,N_14994);
and U17255 (N_17255,N_15231,N_15698);
and U17256 (N_17256,N_14193,N_15764);
nor U17257 (N_17257,N_14203,N_14145);
nand U17258 (N_17258,N_15454,N_15138);
and U17259 (N_17259,N_15273,N_14686);
nor U17260 (N_17260,N_15530,N_14126);
nand U17261 (N_17261,N_14910,N_15871);
or U17262 (N_17262,N_15252,N_15526);
and U17263 (N_17263,N_14401,N_15037);
or U17264 (N_17264,N_15006,N_14999);
and U17265 (N_17265,N_15778,N_14137);
or U17266 (N_17266,N_14453,N_14455);
nor U17267 (N_17267,N_15969,N_14778);
or U17268 (N_17268,N_15811,N_15267);
nand U17269 (N_17269,N_15482,N_14695);
nand U17270 (N_17270,N_15046,N_15174);
and U17271 (N_17271,N_14899,N_15761);
and U17272 (N_17272,N_14141,N_15607);
and U17273 (N_17273,N_15634,N_15192);
and U17274 (N_17274,N_15276,N_15545);
and U17275 (N_17275,N_15811,N_15100);
nand U17276 (N_17276,N_14248,N_15265);
nor U17277 (N_17277,N_15253,N_14440);
and U17278 (N_17278,N_15080,N_15023);
or U17279 (N_17279,N_14559,N_14906);
nand U17280 (N_17280,N_15071,N_15058);
or U17281 (N_17281,N_15788,N_14524);
nor U17282 (N_17282,N_15576,N_14558);
or U17283 (N_17283,N_15752,N_15901);
nand U17284 (N_17284,N_15041,N_14337);
nand U17285 (N_17285,N_15482,N_15029);
xor U17286 (N_17286,N_14479,N_14903);
nand U17287 (N_17287,N_14793,N_14899);
xor U17288 (N_17288,N_15100,N_14063);
nor U17289 (N_17289,N_15335,N_15141);
and U17290 (N_17290,N_14872,N_15241);
nand U17291 (N_17291,N_15973,N_15278);
nand U17292 (N_17292,N_14785,N_15782);
and U17293 (N_17293,N_14089,N_15361);
and U17294 (N_17294,N_14117,N_14051);
or U17295 (N_17295,N_15211,N_15699);
xnor U17296 (N_17296,N_14254,N_14343);
and U17297 (N_17297,N_15547,N_14614);
xnor U17298 (N_17298,N_15584,N_15353);
and U17299 (N_17299,N_15508,N_14831);
and U17300 (N_17300,N_14491,N_15089);
nor U17301 (N_17301,N_14889,N_15669);
nor U17302 (N_17302,N_15426,N_14758);
or U17303 (N_17303,N_14454,N_14897);
or U17304 (N_17304,N_14311,N_14252);
nor U17305 (N_17305,N_14028,N_15824);
nor U17306 (N_17306,N_14480,N_15861);
nand U17307 (N_17307,N_14060,N_15360);
or U17308 (N_17308,N_14754,N_14331);
or U17309 (N_17309,N_15289,N_15861);
or U17310 (N_17310,N_15161,N_15553);
nand U17311 (N_17311,N_14005,N_14290);
nand U17312 (N_17312,N_14858,N_15580);
nand U17313 (N_17313,N_14697,N_14306);
or U17314 (N_17314,N_14896,N_15295);
and U17315 (N_17315,N_15496,N_15158);
or U17316 (N_17316,N_14871,N_14103);
or U17317 (N_17317,N_14765,N_15509);
or U17318 (N_17318,N_15047,N_14080);
and U17319 (N_17319,N_15417,N_15372);
and U17320 (N_17320,N_14628,N_15894);
and U17321 (N_17321,N_15362,N_14009);
or U17322 (N_17322,N_14054,N_15119);
and U17323 (N_17323,N_14074,N_14100);
and U17324 (N_17324,N_14319,N_15832);
and U17325 (N_17325,N_14154,N_14036);
nand U17326 (N_17326,N_14408,N_14938);
and U17327 (N_17327,N_14847,N_14539);
nor U17328 (N_17328,N_15827,N_15213);
xnor U17329 (N_17329,N_15583,N_14228);
nor U17330 (N_17330,N_15345,N_15548);
xnor U17331 (N_17331,N_15202,N_14736);
or U17332 (N_17332,N_15658,N_14485);
or U17333 (N_17333,N_15729,N_15344);
or U17334 (N_17334,N_14813,N_15885);
or U17335 (N_17335,N_15824,N_15847);
or U17336 (N_17336,N_14967,N_14592);
and U17337 (N_17337,N_15993,N_15552);
or U17338 (N_17338,N_14060,N_14340);
and U17339 (N_17339,N_14712,N_14986);
and U17340 (N_17340,N_15381,N_15201);
nand U17341 (N_17341,N_15204,N_14066);
nor U17342 (N_17342,N_15610,N_15179);
and U17343 (N_17343,N_14767,N_14495);
or U17344 (N_17344,N_14377,N_15404);
xnor U17345 (N_17345,N_14176,N_14103);
nor U17346 (N_17346,N_15066,N_15709);
nor U17347 (N_17347,N_14443,N_15957);
nand U17348 (N_17348,N_15874,N_15876);
nor U17349 (N_17349,N_14966,N_15494);
nand U17350 (N_17350,N_15892,N_14423);
and U17351 (N_17351,N_14587,N_14640);
xor U17352 (N_17352,N_15570,N_15999);
nand U17353 (N_17353,N_14134,N_14125);
nand U17354 (N_17354,N_15952,N_14589);
xor U17355 (N_17355,N_15216,N_15587);
nand U17356 (N_17356,N_15116,N_15934);
or U17357 (N_17357,N_15395,N_15933);
nand U17358 (N_17358,N_14327,N_14512);
nor U17359 (N_17359,N_14300,N_14435);
and U17360 (N_17360,N_14920,N_14591);
nand U17361 (N_17361,N_15414,N_14915);
and U17362 (N_17362,N_14169,N_15081);
and U17363 (N_17363,N_14636,N_14443);
and U17364 (N_17364,N_15069,N_15355);
nor U17365 (N_17365,N_15423,N_14779);
or U17366 (N_17366,N_15924,N_15341);
nand U17367 (N_17367,N_14983,N_14153);
nor U17368 (N_17368,N_15763,N_14081);
nand U17369 (N_17369,N_15128,N_15061);
and U17370 (N_17370,N_15366,N_15870);
and U17371 (N_17371,N_15905,N_14269);
and U17372 (N_17372,N_15115,N_15459);
nor U17373 (N_17373,N_14039,N_14855);
nand U17374 (N_17374,N_15893,N_15565);
nand U17375 (N_17375,N_14893,N_14904);
or U17376 (N_17376,N_14310,N_14627);
or U17377 (N_17377,N_15622,N_14903);
and U17378 (N_17378,N_14102,N_14624);
nor U17379 (N_17379,N_14988,N_14429);
nand U17380 (N_17380,N_14982,N_15424);
xor U17381 (N_17381,N_14276,N_14467);
or U17382 (N_17382,N_14071,N_14432);
nor U17383 (N_17383,N_14752,N_14829);
or U17384 (N_17384,N_15370,N_15255);
nand U17385 (N_17385,N_14150,N_15623);
nor U17386 (N_17386,N_15902,N_14852);
nor U17387 (N_17387,N_15898,N_14955);
or U17388 (N_17388,N_15918,N_15798);
and U17389 (N_17389,N_14648,N_15251);
nand U17390 (N_17390,N_14133,N_15294);
and U17391 (N_17391,N_14511,N_14481);
and U17392 (N_17392,N_14687,N_15129);
xnor U17393 (N_17393,N_15708,N_14719);
and U17394 (N_17394,N_15069,N_15681);
and U17395 (N_17395,N_14774,N_14540);
xor U17396 (N_17396,N_15688,N_14676);
or U17397 (N_17397,N_14764,N_14400);
xor U17398 (N_17398,N_15943,N_14074);
and U17399 (N_17399,N_15601,N_14441);
nor U17400 (N_17400,N_14313,N_14770);
and U17401 (N_17401,N_14836,N_14394);
and U17402 (N_17402,N_15493,N_15063);
nor U17403 (N_17403,N_15240,N_14866);
or U17404 (N_17404,N_14611,N_14283);
and U17405 (N_17405,N_14695,N_14665);
nor U17406 (N_17406,N_15568,N_14829);
and U17407 (N_17407,N_14827,N_14092);
nand U17408 (N_17408,N_15251,N_14400);
xnor U17409 (N_17409,N_15339,N_14043);
or U17410 (N_17410,N_15249,N_14392);
nand U17411 (N_17411,N_15885,N_14693);
nand U17412 (N_17412,N_15706,N_15784);
nand U17413 (N_17413,N_14124,N_14787);
or U17414 (N_17414,N_14625,N_15951);
nor U17415 (N_17415,N_15952,N_14990);
nand U17416 (N_17416,N_14525,N_14452);
nand U17417 (N_17417,N_15777,N_15820);
and U17418 (N_17418,N_15745,N_15795);
nand U17419 (N_17419,N_14497,N_15936);
xnor U17420 (N_17420,N_15640,N_15405);
xnor U17421 (N_17421,N_15157,N_15533);
nor U17422 (N_17422,N_15183,N_14667);
or U17423 (N_17423,N_14022,N_14451);
nor U17424 (N_17424,N_14022,N_14982);
nor U17425 (N_17425,N_14424,N_15268);
nand U17426 (N_17426,N_14406,N_14287);
and U17427 (N_17427,N_14728,N_15395);
and U17428 (N_17428,N_14773,N_14847);
nand U17429 (N_17429,N_15863,N_14535);
or U17430 (N_17430,N_15448,N_14133);
or U17431 (N_17431,N_15674,N_14273);
and U17432 (N_17432,N_15011,N_14101);
or U17433 (N_17433,N_15929,N_14969);
nor U17434 (N_17434,N_14342,N_14574);
and U17435 (N_17435,N_15839,N_15900);
nor U17436 (N_17436,N_14644,N_15308);
xnor U17437 (N_17437,N_15745,N_15271);
nand U17438 (N_17438,N_14353,N_15049);
nor U17439 (N_17439,N_14749,N_15037);
nor U17440 (N_17440,N_14082,N_15819);
or U17441 (N_17441,N_14042,N_15710);
and U17442 (N_17442,N_14793,N_14349);
nand U17443 (N_17443,N_14256,N_14183);
nand U17444 (N_17444,N_14416,N_14150);
or U17445 (N_17445,N_14484,N_15909);
and U17446 (N_17446,N_14534,N_15328);
nor U17447 (N_17447,N_15781,N_15455);
nor U17448 (N_17448,N_14849,N_15084);
nand U17449 (N_17449,N_14856,N_15606);
nor U17450 (N_17450,N_15802,N_15498);
nor U17451 (N_17451,N_15351,N_15547);
nor U17452 (N_17452,N_15481,N_14026);
nand U17453 (N_17453,N_14560,N_14359);
nand U17454 (N_17454,N_15548,N_14630);
and U17455 (N_17455,N_15404,N_14818);
and U17456 (N_17456,N_14790,N_15603);
or U17457 (N_17457,N_15271,N_15251);
or U17458 (N_17458,N_14098,N_14261);
nor U17459 (N_17459,N_15648,N_14988);
or U17460 (N_17460,N_14217,N_14062);
and U17461 (N_17461,N_14387,N_15690);
or U17462 (N_17462,N_14085,N_15778);
or U17463 (N_17463,N_15279,N_14729);
nand U17464 (N_17464,N_15459,N_14793);
nor U17465 (N_17465,N_14066,N_15089);
and U17466 (N_17466,N_15012,N_15308);
and U17467 (N_17467,N_14724,N_15357);
or U17468 (N_17468,N_14925,N_14096);
nor U17469 (N_17469,N_14501,N_14217);
nand U17470 (N_17470,N_15561,N_15768);
xnor U17471 (N_17471,N_14326,N_15775);
nand U17472 (N_17472,N_14378,N_14727);
nand U17473 (N_17473,N_14177,N_15751);
or U17474 (N_17474,N_14873,N_15010);
or U17475 (N_17475,N_15166,N_15037);
nand U17476 (N_17476,N_14222,N_14942);
and U17477 (N_17477,N_14406,N_14940);
nor U17478 (N_17478,N_14300,N_14990);
nand U17479 (N_17479,N_14363,N_15485);
and U17480 (N_17480,N_15722,N_14684);
or U17481 (N_17481,N_15585,N_14642);
nand U17482 (N_17482,N_14540,N_15594);
or U17483 (N_17483,N_15163,N_15856);
and U17484 (N_17484,N_14567,N_15558);
or U17485 (N_17485,N_14533,N_14621);
and U17486 (N_17486,N_14375,N_14868);
and U17487 (N_17487,N_15305,N_15752);
nand U17488 (N_17488,N_15000,N_14525);
nand U17489 (N_17489,N_14714,N_15415);
and U17490 (N_17490,N_14366,N_15498);
nand U17491 (N_17491,N_14031,N_15534);
or U17492 (N_17492,N_14935,N_15361);
nand U17493 (N_17493,N_14357,N_15365);
nor U17494 (N_17494,N_15115,N_14057);
nor U17495 (N_17495,N_14398,N_15149);
and U17496 (N_17496,N_14717,N_15779);
nor U17497 (N_17497,N_15135,N_15603);
xnor U17498 (N_17498,N_14025,N_15085);
or U17499 (N_17499,N_15871,N_14372);
and U17500 (N_17500,N_15719,N_15751);
nand U17501 (N_17501,N_14918,N_14675);
or U17502 (N_17502,N_14351,N_14536);
or U17503 (N_17503,N_14463,N_15886);
nor U17504 (N_17504,N_14083,N_14697);
or U17505 (N_17505,N_15700,N_14064);
or U17506 (N_17506,N_15453,N_15600);
and U17507 (N_17507,N_15956,N_14282);
nand U17508 (N_17508,N_15313,N_15851);
and U17509 (N_17509,N_15004,N_14815);
nor U17510 (N_17510,N_14863,N_15056);
and U17511 (N_17511,N_14010,N_14854);
nor U17512 (N_17512,N_15825,N_14319);
nand U17513 (N_17513,N_15298,N_15316);
or U17514 (N_17514,N_15846,N_14699);
nor U17515 (N_17515,N_14351,N_15873);
or U17516 (N_17516,N_14101,N_15007);
and U17517 (N_17517,N_15783,N_14983);
and U17518 (N_17518,N_15359,N_14101);
nor U17519 (N_17519,N_14770,N_15575);
nand U17520 (N_17520,N_15097,N_15394);
nor U17521 (N_17521,N_14021,N_14554);
or U17522 (N_17522,N_14598,N_14802);
nand U17523 (N_17523,N_14818,N_15399);
or U17524 (N_17524,N_14038,N_15369);
xor U17525 (N_17525,N_15979,N_15512);
and U17526 (N_17526,N_14786,N_14262);
xnor U17527 (N_17527,N_15013,N_14514);
or U17528 (N_17528,N_15396,N_15289);
nor U17529 (N_17529,N_14546,N_14442);
nor U17530 (N_17530,N_14713,N_15347);
nand U17531 (N_17531,N_14198,N_14386);
nand U17532 (N_17532,N_14076,N_15484);
xnor U17533 (N_17533,N_15644,N_15118);
and U17534 (N_17534,N_14160,N_15480);
nor U17535 (N_17535,N_14106,N_14832);
or U17536 (N_17536,N_15082,N_15464);
xor U17537 (N_17537,N_14190,N_15660);
and U17538 (N_17538,N_15179,N_14548);
nand U17539 (N_17539,N_15182,N_14339);
and U17540 (N_17540,N_15652,N_15444);
or U17541 (N_17541,N_14438,N_14080);
xnor U17542 (N_17542,N_15214,N_14291);
or U17543 (N_17543,N_14669,N_15957);
or U17544 (N_17544,N_15206,N_14834);
nor U17545 (N_17545,N_15355,N_15058);
or U17546 (N_17546,N_14671,N_15728);
or U17547 (N_17547,N_14298,N_14700);
and U17548 (N_17548,N_14780,N_14915);
nor U17549 (N_17549,N_14953,N_15290);
nand U17550 (N_17550,N_15850,N_14108);
nand U17551 (N_17551,N_15077,N_15777);
or U17552 (N_17552,N_14806,N_14484);
xor U17553 (N_17553,N_15326,N_14460);
nand U17554 (N_17554,N_15841,N_15671);
xnor U17555 (N_17555,N_15844,N_14734);
or U17556 (N_17556,N_14697,N_14456);
or U17557 (N_17557,N_14116,N_14746);
xnor U17558 (N_17558,N_14848,N_15687);
nand U17559 (N_17559,N_15505,N_15655);
nand U17560 (N_17560,N_15198,N_15077);
nor U17561 (N_17561,N_15405,N_14123);
or U17562 (N_17562,N_15117,N_14014);
and U17563 (N_17563,N_14174,N_15011);
nor U17564 (N_17564,N_15067,N_14356);
nor U17565 (N_17565,N_15058,N_15225);
or U17566 (N_17566,N_15039,N_14271);
and U17567 (N_17567,N_14281,N_14734);
nor U17568 (N_17568,N_15059,N_14460);
and U17569 (N_17569,N_14361,N_14538);
and U17570 (N_17570,N_14401,N_15428);
nor U17571 (N_17571,N_15510,N_15136);
nor U17572 (N_17572,N_14306,N_15805);
xnor U17573 (N_17573,N_15313,N_14995);
nor U17574 (N_17574,N_15317,N_14992);
or U17575 (N_17575,N_15068,N_14511);
and U17576 (N_17576,N_15529,N_15687);
or U17577 (N_17577,N_14473,N_15836);
nand U17578 (N_17578,N_14704,N_14174);
nor U17579 (N_17579,N_14990,N_15136);
xnor U17580 (N_17580,N_14235,N_14660);
nand U17581 (N_17581,N_14746,N_14885);
and U17582 (N_17582,N_15481,N_14623);
nor U17583 (N_17583,N_14043,N_15774);
nand U17584 (N_17584,N_15160,N_14059);
and U17585 (N_17585,N_14535,N_14714);
or U17586 (N_17586,N_15720,N_14992);
and U17587 (N_17587,N_14454,N_15696);
nand U17588 (N_17588,N_15208,N_15625);
and U17589 (N_17589,N_15201,N_15046);
xnor U17590 (N_17590,N_14201,N_15868);
and U17591 (N_17591,N_14415,N_15356);
and U17592 (N_17592,N_15580,N_14461);
or U17593 (N_17593,N_14638,N_14863);
or U17594 (N_17594,N_14802,N_15210);
nand U17595 (N_17595,N_15176,N_14214);
nor U17596 (N_17596,N_15585,N_15416);
nand U17597 (N_17597,N_15939,N_14461);
nor U17598 (N_17598,N_14462,N_15732);
nand U17599 (N_17599,N_15696,N_14220);
or U17600 (N_17600,N_14271,N_14621);
and U17601 (N_17601,N_14139,N_14641);
nand U17602 (N_17602,N_15059,N_14949);
and U17603 (N_17603,N_15211,N_14789);
or U17604 (N_17604,N_15169,N_14439);
or U17605 (N_17605,N_14572,N_14440);
xnor U17606 (N_17606,N_14957,N_15326);
or U17607 (N_17607,N_15202,N_15262);
or U17608 (N_17608,N_14568,N_14946);
or U17609 (N_17609,N_14076,N_14239);
and U17610 (N_17610,N_14184,N_15440);
or U17611 (N_17611,N_15593,N_14005);
and U17612 (N_17612,N_15007,N_15212);
nand U17613 (N_17613,N_14809,N_14095);
xor U17614 (N_17614,N_14499,N_14365);
nor U17615 (N_17615,N_15544,N_15918);
and U17616 (N_17616,N_14171,N_15675);
nor U17617 (N_17617,N_14565,N_14527);
and U17618 (N_17618,N_15573,N_15926);
and U17619 (N_17619,N_15767,N_14143);
and U17620 (N_17620,N_15279,N_14475);
and U17621 (N_17621,N_14679,N_15834);
nor U17622 (N_17622,N_15779,N_15563);
nor U17623 (N_17623,N_14684,N_14190);
nand U17624 (N_17624,N_14682,N_15552);
or U17625 (N_17625,N_14407,N_15126);
nand U17626 (N_17626,N_14938,N_14233);
and U17627 (N_17627,N_14510,N_15665);
and U17628 (N_17628,N_15091,N_15449);
xor U17629 (N_17629,N_15241,N_15230);
and U17630 (N_17630,N_14921,N_14353);
or U17631 (N_17631,N_15260,N_14838);
nand U17632 (N_17632,N_14668,N_14821);
nand U17633 (N_17633,N_15024,N_14709);
nor U17634 (N_17634,N_14204,N_15497);
and U17635 (N_17635,N_14584,N_14905);
nor U17636 (N_17636,N_15062,N_15012);
nand U17637 (N_17637,N_14204,N_14250);
nor U17638 (N_17638,N_14304,N_14122);
or U17639 (N_17639,N_15369,N_15955);
xnor U17640 (N_17640,N_15572,N_15713);
xor U17641 (N_17641,N_15734,N_14932);
and U17642 (N_17642,N_15866,N_14218);
nor U17643 (N_17643,N_14325,N_14578);
nand U17644 (N_17644,N_15136,N_14614);
nand U17645 (N_17645,N_15644,N_14688);
or U17646 (N_17646,N_14753,N_15996);
and U17647 (N_17647,N_15851,N_14516);
or U17648 (N_17648,N_14271,N_15145);
or U17649 (N_17649,N_15516,N_14313);
and U17650 (N_17650,N_15025,N_15616);
nor U17651 (N_17651,N_15861,N_15911);
nand U17652 (N_17652,N_15907,N_15194);
xor U17653 (N_17653,N_15368,N_15537);
nor U17654 (N_17654,N_14843,N_14208);
or U17655 (N_17655,N_14626,N_14832);
or U17656 (N_17656,N_15271,N_15710);
and U17657 (N_17657,N_14457,N_15071);
or U17658 (N_17658,N_15947,N_14375);
nand U17659 (N_17659,N_15648,N_14518);
or U17660 (N_17660,N_15317,N_15348);
nor U17661 (N_17661,N_14866,N_14193);
and U17662 (N_17662,N_14382,N_15880);
xor U17663 (N_17663,N_14768,N_15348);
xor U17664 (N_17664,N_14233,N_14527);
and U17665 (N_17665,N_14270,N_15973);
and U17666 (N_17666,N_14954,N_15888);
xnor U17667 (N_17667,N_14479,N_14748);
nand U17668 (N_17668,N_15424,N_15198);
nor U17669 (N_17669,N_14032,N_14240);
xnor U17670 (N_17670,N_14859,N_14124);
xnor U17671 (N_17671,N_15845,N_15995);
and U17672 (N_17672,N_14904,N_15796);
nor U17673 (N_17673,N_15741,N_14655);
or U17674 (N_17674,N_15889,N_14738);
and U17675 (N_17675,N_14091,N_14989);
xor U17676 (N_17676,N_14199,N_14811);
and U17677 (N_17677,N_15316,N_15135);
or U17678 (N_17678,N_14266,N_15151);
nand U17679 (N_17679,N_15746,N_14610);
or U17680 (N_17680,N_14762,N_15581);
nor U17681 (N_17681,N_14784,N_14641);
and U17682 (N_17682,N_15251,N_14180);
xnor U17683 (N_17683,N_15254,N_14001);
nor U17684 (N_17684,N_15812,N_15856);
xor U17685 (N_17685,N_15291,N_14016);
and U17686 (N_17686,N_14741,N_15595);
nand U17687 (N_17687,N_15903,N_15703);
nor U17688 (N_17688,N_14089,N_15910);
nand U17689 (N_17689,N_15201,N_15181);
and U17690 (N_17690,N_14212,N_14055);
and U17691 (N_17691,N_15397,N_15746);
nand U17692 (N_17692,N_14066,N_14037);
or U17693 (N_17693,N_15289,N_14591);
or U17694 (N_17694,N_14892,N_14549);
or U17695 (N_17695,N_15907,N_15419);
nand U17696 (N_17696,N_14089,N_14169);
nand U17697 (N_17697,N_14008,N_15845);
nor U17698 (N_17698,N_15750,N_15945);
and U17699 (N_17699,N_14711,N_15661);
nand U17700 (N_17700,N_15160,N_15288);
nand U17701 (N_17701,N_14884,N_14674);
xnor U17702 (N_17702,N_15583,N_15485);
nor U17703 (N_17703,N_15199,N_14853);
nor U17704 (N_17704,N_15818,N_15352);
or U17705 (N_17705,N_15030,N_14068);
and U17706 (N_17706,N_15444,N_14803);
nor U17707 (N_17707,N_14491,N_14241);
or U17708 (N_17708,N_15459,N_14862);
or U17709 (N_17709,N_15651,N_14499);
or U17710 (N_17710,N_15623,N_14941);
nor U17711 (N_17711,N_14245,N_15871);
xor U17712 (N_17712,N_15781,N_15673);
nand U17713 (N_17713,N_15107,N_15464);
and U17714 (N_17714,N_15424,N_14953);
or U17715 (N_17715,N_14026,N_14288);
nand U17716 (N_17716,N_15696,N_15973);
nor U17717 (N_17717,N_15632,N_15469);
nand U17718 (N_17718,N_15820,N_15468);
xor U17719 (N_17719,N_14307,N_14439);
or U17720 (N_17720,N_15885,N_14157);
nand U17721 (N_17721,N_15084,N_14523);
or U17722 (N_17722,N_14951,N_14065);
and U17723 (N_17723,N_14669,N_14570);
nor U17724 (N_17724,N_15716,N_14184);
nor U17725 (N_17725,N_15079,N_14267);
nor U17726 (N_17726,N_15098,N_15370);
nor U17727 (N_17727,N_15383,N_15484);
and U17728 (N_17728,N_15670,N_15451);
nand U17729 (N_17729,N_15715,N_15519);
and U17730 (N_17730,N_15724,N_15229);
and U17731 (N_17731,N_15616,N_14567);
nor U17732 (N_17732,N_14055,N_15544);
or U17733 (N_17733,N_15496,N_14269);
nand U17734 (N_17734,N_14427,N_14734);
nand U17735 (N_17735,N_15108,N_15316);
nand U17736 (N_17736,N_15851,N_14617);
or U17737 (N_17737,N_14584,N_14102);
nor U17738 (N_17738,N_14530,N_15365);
xor U17739 (N_17739,N_14562,N_14786);
xnor U17740 (N_17740,N_14030,N_15486);
and U17741 (N_17741,N_14064,N_14554);
and U17742 (N_17742,N_15653,N_14018);
nand U17743 (N_17743,N_15699,N_14822);
or U17744 (N_17744,N_14301,N_14052);
and U17745 (N_17745,N_14879,N_14529);
xor U17746 (N_17746,N_14703,N_15294);
xor U17747 (N_17747,N_14905,N_15359);
and U17748 (N_17748,N_15216,N_15461);
or U17749 (N_17749,N_14073,N_14007);
nor U17750 (N_17750,N_14719,N_14045);
or U17751 (N_17751,N_15523,N_15610);
nor U17752 (N_17752,N_14458,N_15789);
nand U17753 (N_17753,N_14181,N_14946);
nor U17754 (N_17754,N_15025,N_14557);
nor U17755 (N_17755,N_14008,N_15693);
nor U17756 (N_17756,N_15344,N_14777);
and U17757 (N_17757,N_15300,N_15161);
or U17758 (N_17758,N_14085,N_14426);
and U17759 (N_17759,N_14963,N_14490);
or U17760 (N_17760,N_15433,N_15153);
or U17761 (N_17761,N_14072,N_15730);
and U17762 (N_17762,N_14223,N_15142);
xor U17763 (N_17763,N_14399,N_14580);
nor U17764 (N_17764,N_15650,N_15428);
nor U17765 (N_17765,N_15674,N_15456);
nor U17766 (N_17766,N_15409,N_14032);
or U17767 (N_17767,N_14047,N_14623);
nor U17768 (N_17768,N_14936,N_14477);
nand U17769 (N_17769,N_15372,N_15732);
xnor U17770 (N_17770,N_14613,N_15313);
or U17771 (N_17771,N_14417,N_15174);
xor U17772 (N_17772,N_14256,N_15809);
nor U17773 (N_17773,N_15598,N_14958);
nor U17774 (N_17774,N_15288,N_14586);
or U17775 (N_17775,N_14364,N_14262);
and U17776 (N_17776,N_14859,N_15868);
nor U17777 (N_17777,N_15162,N_14490);
nor U17778 (N_17778,N_14840,N_14393);
or U17779 (N_17779,N_14716,N_15484);
or U17780 (N_17780,N_14180,N_15997);
xnor U17781 (N_17781,N_15446,N_14430);
or U17782 (N_17782,N_15294,N_15161);
nand U17783 (N_17783,N_15074,N_14220);
or U17784 (N_17784,N_14480,N_15014);
nand U17785 (N_17785,N_15012,N_14786);
or U17786 (N_17786,N_14494,N_15843);
and U17787 (N_17787,N_15978,N_15756);
xnor U17788 (N_17788,N_15069,N_15075);
xor U17789 (N_17789,N_14350,N_15267);
nor U17790 (N_17790,N_15266,N_15814);
nand U17791 (N_17791,N_15943,N_14952);
nand U17792 (N_17792,N_15783,N_15732);
and U17793 (N_17793,N_15432,N_15566);
nor U17794 (N_17794,N_14200,N_15741);
xor U17795 (N_17795,N_14133,N_15164);
and U17796 (N_17796,N_14980,N_15990);
xor U17797 (N_17797,N_15154,N_15757);
nand U17798 (N_17798,N_14749,N_15750);
nor U17799 (N_17799,N_14179,N_15841);
xnor U17800 (N_17800,N_15006,N_14593);
xnor U17801 (N_17801,N_14701,N_15522);
nand U17802 (N_17802,N_15440,N_15379);
and U17803 (N_17803,N_14309,N_15641);
nand U17804 (N_17804,N_14495,N_15872);
nor U17805 (N_17805,N_15889,N_15406);
or U17806 (N_17806,N_15294,N_15765);
nand U17807 (N_17807,N_15205,N_15915);
or U17808 (N_17808,N_15897,N_14350);
or U17809 (N_17809,N_15115,N_15747);
and U17810 (N_17810,N_14697,N_14142);
nor U17811 (N_17811,N_15616,N_14687);
nor U17812 (N_17812,N_14290,N_15321);
xor U17813 (N_17813,N_15583,N_15797);
and U17814 (N_17814,N_14941,N_15857);
and U17815 (N_17815,N_15941,N_14696);
xnor U17816 (N_17816,N_15561,N_15731);
nor U17817 (N_17817,N_15954,N_15982);
nor U17818 (N_17818,N_15747,N_14680);
and U17819 (N_17819,N_15092,N_15376);
or U17820 (N_17820,N_14688,N_14328);
nor U17821 (N_17821,N_15504,N_14703);
and U17822 (N_17822,N_14076,N_14707);
and U17823 (N_17823,N_14877,N_14053);
and U17824 (N_17824,N_14523,N_14130);
and U17825 (N_17825,N_15178,N_14139);
nand U17826 (N_17826,N_14848,N_15139);
xor U17827 (N_17827,N_15554,N_15578);
and U17828 (N_17828,N_14183,N_15046);
or U17829 (N_17829,N_15112,N_14361);
and U17830 (N_17830,N_15853,N_15172);
nand U17831 (N_17831,N_14180,N_14385);
nand U17832 (N_17832,N_14458,N_14705);
or U17833 (N_17833,N_15132,N_14226);
nor U17834 (N_17834,N_15122,N_14343);
nand U17835 (N_17835,N_14151,N_14519);
or U17836 (N_17836,N_15264,N_14882);
or U17837 (N_17837,N_15431,N_15394);
nor U17838 (N_17838,N_14858,N_14548);
or U17839 (N_17839,N_15769,N_15263);
nand U17840 (N_17840,N_14428,N_14247);
nor U17841 (N_17841,N_15995,N_14656);
or U17842 (N_17842,N_14586,N_14009);
nor U17843 (N_17843,N_15817,N_15527);
or U17844 (N_17844,N_14138,N_14258);
nand U17845 (N_17845,N_14087,N_14529);
and U17846 (N_17846,N_14142,N_14149);
xnor U17847 (N_17847,N_14838,N_15279);
nor U17848 (N_17848,N_14985,N_15831);
and U17849 (N_17849,N_15546,N_15711);
and U17850 (N_17850,N_14009,N_15742);
nand U17851 (N_17851,N_14477,N_14101);
or U17852 (N_17852,N_15703,N_14041);
nor U17853 (N_17853,N_15872,N_14878);
or U17854 (N_17854,N_15856,N_14316);
nand U17855 (N_17855,N_15914,N_15573);
or U17856 (N_17856,N_15466,N_14906);
or U17857 (N_17857,N_14143,N_15499);
and U17858 (N_17858,N_15635,N_14937);
or U17859 (N_17859,N_14392,N_15538);
and U17860 (N_17860,N_14362,N_14094);
and U17861 (N_17861,N_14956,N_14712);
or U17862 (N_17862,N_14401,N_14877);
or U17863 (N_17863,N_14080,N_14911);
and U17864 (N_17864,N_14526,N_15389);
nor U17865 (N_17865,N_14479,N_14447);
nand U17866 (N_17866,N_15504,N_15381);
nor U17867 (N_17867,N_14724,N_15302);
and U17868 (N_17868,N_14688,N_14222);
and U17869 (N_17869,N_15463,N_14018);
nor U17870 (N_17870,N_15321,N_15599);
and U17871 (N_17871,N_15778,N_14581);
nand U17872 (N_17872,N_14375,N_15894);
nand U17873 (N_17873,N_14583,N_14926);
xnor U17874 (N_17874,N_14252,N_15455);
nand U17875 (N_17875,N_14998,N_15181);
nor U17876 (N_17876,N_15688,N_15637);
nor U17877 (N_17877,N_15155,N_15137);
and U17878 (N_17878,N_14267,N_14880);
nor U17879 (N_17879,N_14225,N_14319);
and U17880 (N_17880,N_14274,N_14984);
and U17881 (N_17881,N_14983,N_14882);
or U17882 (N_17882,N_15400,N_14399);
nor U17883 (N_17883,N_14988,N_14801);
and U17884 (N_17884,N_14128,N_15343);
xnor U17885 (N_17885,N_14194,N_15498);
and U17886 (N_17886,N_15698,N_14384);
nor U17887 (N_17887,N_15529,N_14505);
nand U17888 (N_17888,N_14546,N_15959);
xor U17889 (N_17889,N_14398,N_14420);
nor U17890 (N_17890,N_15748,N_15781);
nand U17891 (N_17891,N_15230,N_15770);
and U17892 (N_17892,N_14639,N_15156);
nor U17893 (N_17893,N_15319,N_15641);
or U17894 (N_17894,N_15247,N_14618);
nand U17895 (N_17895,N_15168,N_14500);
and U17896 (N_17896,N_14850,N_14909);
nor U17897 (N_17897,N_14747,N_14497);
and U17898 (N_17898,N_15524,N_15287);
or U17899 (N_17899,N_15169,N_15403);
or U17900 (N_17900,N_15892,N_15275);
and U17901 (N_17901,N_14661,N_14345);
nand U17902 (N_17902,N_14866,N_14079);
nor U17903 (N_17903,N_15181,N_15452);
nand U17904 (N_17904,N_15933,N_15215);
nand U17905 (N_17905,N_14726,N_14688);
and U17906 (N_17906,N_14119,N_15111);
or U17907 (N_17907,N_15968,N_14941);
xor U17908 (N_17908,N_15928,N_14018);
xor U17909 (N_17909,N_14641,N_14686);
or U17910 (N_17910,N_15133,N_15357);
and U17911 (N_17911,N_15923,N_15530);
and U17912 (N_17912,N_15121,N_15652);
xnor U17913 (N_17913,N_14752,N_15597);
nor U17914 (N_17914,N_14283,N_15789);
nor U17915 (N_17915,N_14463,N_14366);
or U17916 (N_17916,N_15850,N_15798);
nand U17917 (N_17917,N_14734,N_15753);
nor U17918 (N_17918,N_14120,N_14594);
nor U17919 (N_17919,N_15097,N_15386);
nor U17920 (N_17920,N_14459,N_14529);
and U17921 (N_17921,N_15398,N_14643);
nand U17922 (N_17922,N_15668,N_15268);
or U17923 (N_17923,N_15137,N_14050);
nand U17924 (N_17924,N_15478,N_14127);
and U17925 (N_17925,N_14136,N_14794);
and U17926 (N_17926,N_14520,N_14489);
nor U17927 (N_17927,N_14608,N_14517);
and U17928 (N_17928,N_15782,N_15615);
and U17929 (N_17929,N_14462,N_15854);
nor U17930 (N_17930,N_14776,N_15174);
nor U17931 (N_17931,N_15118,N_15968);
and U17932 (N_17932,N_15657,N_15442);
xnor U17933 (N_17933,N_15214,N_14829);
nor U17934 (N_17934,N_14580,N_14165);
and U17935 (N_17935,N_14586,N_15123);
xor U17936 (N_17936,N_14288,N_14704);
nand U17937 (N_17937,N_15270,N_15519);
and U17938 (N_17938,N_14870,N_14704);
nand U17939 (N_17939,N_15866,N_15267);
nand U17940 (N_17940,N_15263,N_15906);
or U17941 (N_17941,N_14467,N_15044);
and U17942 (N_17942,N_15180,N_14015);
nand U17943 (N_17943,N_14951,N_15064);
nand U17944 (N_17944,N_15432,N_15685);
and U17945 (N_17945,N_14821,N_14793);
and U17946 (N_17946,N_15707,N_15735);
and U17947 (N_17947,N_14523,N_14775);
nand U17948 (N_17948,N_14960,N_14527);
nor U17949 (N_17949,N_15683,N_14913);
nand U17950 (N_17950,N_14046,N_14209);
and U17951 (N_17951,N_15608,N_15702);
nand U17952 (N_17952,N_15061,N_15902);
xnor U17953 (N_17953,N_14019,N_15564);
xor U17954 (N_17954,N_14464,N_14944);
nor U17955 (N_17955,N_15511,N_14915);
xor U17956 (N_17956,N_15741,N_15341);
nand U17957 (N_17957,N_14189,N_14956);
nor U17958 (N_17958,N_15555,N_15077);
or U17959 (N_17959,N_14151,N_15299);
and U17960 (N_17960,N_15659,N_14819);
nand U17961 (N_17961,N_14633,N_15141);
nor U17962 (N_17962,N_14127,N_14765);
or U17963 (N_17963,N_14077,N_14726);
or U17964 (N_17964,N_14951,N_14702);
or U17965 (N_17965,N_15482,N_15579);
nor U17966 (N_17966,N_15812,N_15043);
nor U17967 (N_17967,N_15433,N_15629);
or U17968 (N_17968,N_15746,N_15161);
xor U17969 (N_17969,N_15270,N_14165);
and U17970 (N_17970,N_15781,N_14084);
nor U17971 (N_17971,N_14204,N_14811);
xor U17972 (N_17972,N_15245,N_14848);
or U17973 (N_17973,N_14592,N_14537);
xor U17974 (N_17974,N_14193,N_14488);
or U17975 (N_17975,N_15090,N_14907);
or U17976 (N_17976,N_15911,N_15889);
nand U17977 (N_17977,N_14085,N_15427);
or U17978 (N_17978,N_15372,N_14846);
nand U17979 (N_17979,N_15760,N_14773);
or U17980 (N_17980,N_15193,N_14072);
or U17981 (N_17981,N_15125,N_14295);
nor U17982 (N_17982,N_15475,N_14175);
or U17983 (N_17983,N_14445,N_15667);
or U17984 (N_17984,N_15931,N_14890);
and U17985 (N_17985,N_14019,N_14507);
nand U17986 (N_17986,N_15326,N_15596);
or U17987 (N_17987,N_14186,N_15164);
nand U17988 (N_17988,N_15411,N_15347);
nand U17989 (N_17989,N_14241,N_15545);
nor U17990 (N_17990,N_14257,N_14651);
or U17991 (N_17991,N_14734,N_14327);
nor U17992 (N_17992,N_15057,N_14335);
and U17993 (N_17993,N_15580,N_14804);
and U17994 (N_17994,N_15783,N_14885);
and U17995 (N_17995,N_14250,N_14883);
or U17996 (N_17996,N_14701,N_15344);
and U17997 (N_17997,N_14261,N_14466);
and U17998 (N_17998,N_14552,N_14860);
nand U17999 (N_17999,N_14735,N_15622);
or U18000 (N_18000,N_16051,N_17372);
xnor U18001 (N_18001,N_17580,N_16583);
and U18002 (N_18002,N_16373,N_16034);
nor U18003 (N_18003,N_16570,N_16790);
or U18004 (N_18004,N_16385,N_16947);
or U18005 (N_18005,N_17857,N_17116);
and U18006 (N_18006,N_17245,N_16736);
nand U18007 (N_18007,N_17640,N_16552);
nor U18008 (N_18008,N_17668,N_17191);
nand U18009 (N_18009,N_17928,N_16620);
and U18010 (N_18010,N_16329,N_16337);
nor U18011 (N_18011,N_17330,N_17209);
nand U18012 (N_18012,N_16954,N_16355);
nand U18013 (N_18013,N_17195,N_17218);
nor U18014 (N_18014,N_17427,N_17146);
and U18015 (N_18015,N_17441,N_16461);
or U18016 (N_18016,N_17738,N_16435);
nand U18017 (N_18017,N_17243,N_17981);
nand U18018 (N_18018,N_17530,N_17314);
and U18019 (N_18019,N_17112,N_17135);
xor U18020 (N_18020,N_16619,N_17302);
xnor U18021 (N_18021,N_17154,N_17782);
nand U18022 (N_18022,N_16036,N_17123);
or U18023 (N_18023,N_16543,N_17333);
xnor U18024 (N_18024,N_17560,N_16952);
or U18025 (N_18025,N_17194,N_17617);
or U18026 (N_18026,N_17970,N_16161);
nor U18027 (N_18027,N_17674,N_17309);
nand U18028 (N_18028,N_16926,N_17865);
and U18029 (N_18029,N_16976,N_17358);
or U18030 (N_18030,N_17371,N_17327);
nor U18031 (N_18031,N_16037,N_17238);
nor U18032 (N_18032,N_17190,N_16382);
nor U18033 (N_18033,N_16213,N_17517);
nand U18034 (N_18034,N_17284,N_16399);
or U18035 (N_18035,N_17702,N_16727);
nand U18036 (N_18036,N_16520,N_16705);
nand U18037 (N_18037,N_16966,N_17055);
or U18038 (N_18038,N_16669,N_16055);
nand U18039 (N_18039,N_17043,N_16794);
nor U18040 (N_18040,N_16428,N_16141);
or U18041 (N_18041,N_16609,N_17313);
or U18042 (N_18042,N_16652,N_16556);
and U18043 (N_18043,N_17585,N_16606);
or U18044 (N_18044,N_16121,N_17077);
nor U18045 (N_18045,N_17616,N_16944);
nor U18046 (N_18046,N_16978,N_17815);
nand U18047 (N_18047,N_16804,N_17796);
xor U18048 (N_18048,N_17794,N_16054);
nand U18049 (N_18049,N_16714,N_17628);
nand U18050 (N_18050,N_17395,N_17021);
nand U18051 (N_18051,N_16144,N_16601);
or U18052 (N_18052,N_16759,N_16352);
nor U18053 (N_18053,N_16394,N_17162);
nand U18054 (N_18054,N_16529,N_17268);
nand U18055 (N_18055,N_16292,N_16080);
nand U18056 (N_18056,N_16668,N_16995);
nor U18057 (N_18057,N_17932,N_16143);
or U18058 (N_18058,N_16236,N_17801);
or U18059 (N_18059,N_17786,N_17565);
or U18060 (N_18060,N_16047,N_16949);
and U18061 (N_18061,N_17233,N_17375);
and U18062 (N_18062,N_16238,N_17224);
and U18063 (N_18063,N_16380,N_17673);
and U18064 (N_18064,N_17849,N_17927);
nand U18065 (N_18065,N_17282,N_17011);
nand U18066 (N_18066,N_16354,N_17956);
and U18067 (N_18067,N_17365,N_17509);
nand U18068 (N_18068,N_17856,N_16634);
or U18069 (N_18069,N_17340,N_17472);
and U18070 (N_18070,N_16659,N_16776);
xnor U18071 (N_18071,N_16280,N_17665);
nor U18072 (N_18072,N_17113,N_16683);
nand U18073 (N_18073,N_17120,N_17009);
nor U18074 (N_18074,N_17583,N_16499);
and U18075 (N_18075,N_16965,N_16909);
nor U18076 (N_18076,N_17418,N_17939);
nor U18077 (N_18077,N_16426,N_17017);
nand U18078 (N_18078,N_16192,N_17273);
and U18079 (N_18079,N_17553,N_17539);
xor U18080 (N_18080,N_16523,N_16469);
nor U18081 (N_18081,N_17103,N_16734);
nand U18082 (N_18082,N_16119,N_17609);
xor U18083 (N_18083,N_17424,N_16123);
nor U18084 (N_18084,N_16827,N_17745);
nand U18085 (N_18085,N_17290,N_17437);
nor U18086 (N_18086,N_17248,N_16240);
and U18087 (N_18087,N_16819,N_16842);
or U18088 (N_18088,N_17513,N_16877);
nor U18089 (N_18089,N_17608,N_16530);
nand U18090 (N_18090,N_16235,N_16832);
nand U18091 (N_18091,N_16189,N_16190);
nand U18092 (N_18092,N_16470,N_17597);
and U18093 (N_18093,N_17543,N_16968);
and U18094 (N_18094,N_16664,N_16277);
nand U18095 (N_18095,N_16741,N_16745);
nor U18096 (N_18096,N_17386,N_16089);
or U18097 (N_18097,N_17459,N_16546);
and U18098 (N_18098,N_17831,N_17707);
nand U18099 (N_18099,N_17873,N_16950);
nand U18100 (N_18100,N_16961,N_16694);
and U18101 (N_18101,N_17752,N_17571);
or U18102 (N_18102,N_17911,N_16281);
or U18103 (N_18103,N_17312,N_17064);
and U18104 (N_18104,N_16211,N_16140);
or U18105 (N_18105,N_16891,N_17540);
nor U18106 (N_18106,N_17983,N_17883);
nand U18107 (N_18107,N_17817,N_17769);
and U18108 (N_18108,N_16622,N_16107);
or U18109 (N_18109,N_16624,N_16414);
or U18110 (N_18110,N_17357,N_16490);
nand U18111 (N_18111,N_16838,N_17534);
nand U18112 (N_18112,N_17071,N_16974);
nand U18113 (N_18113,N_17014,N_16628);
or U18114 (N_18114,N_16287,N_17023);
nor U18115 (N_18115,N_17980,N_16605);
and U18116 (N_18116,N_16333,N_17955);
and U18117 (N_18117,N_16406,N_16769);
and U18118 (N_18118,N_16715,N_16707);
nand U18119 (N_18119,N_16188,N_16320);
nand U18120 (N_18120,N_17004,N_16166);
and U18121 (N_18121,N_17464,N_16805);
nor U18122 (N_18122,N_16489,N_16308);
xor U18123 (N_18123,N_16990,N_17034);
xnor U18124 (N_18124,N_16222,N_17723);
xnor U18125 (N_18125,N_17754,N_17767);
nand U18126 (N_18126,N_17966,N_16996);
or U18127 (N_18127,N_17364,N_17991);
nand U18128 (N_18128,N_17184,N_16039);
nor U18129 (N_18129,N_16148,N_17404);
xor U18130 (N_18130,N_16972,N_16104);
and U18131 (N_18131,N_16049,N_16288);
and U18132 (N_18132,N_16510,N_17703);
and U18133 (N_18133,N_17076,N_16366);
nor U18134 (N_18134,N_16205,N_16969);
nor U18135 (N_18135,N_16883,N_17353);
or U18136 (N_18136,N_16336,N_16252);
nor U18137 (N_18137,N_16194,N_16370);
and U18138 (N_18138,N_17163,N_17827);
nor U18139 (N_18139,N_16822,N_16106);
or U18140 (N_18140,N_17507,N_17699);
nor U18141 (N_18141,N_16914,N_17015);
and U18142 (N_18142,N_17285,N_17943);
nand U18143 (N_18143,N_17663,N_17447);
xor U18144 (N_18144,N_17689,N_17721);
and U18145 (N_18145,N_16591,N_16022);
nor U18146 (N_18146,N_17893,N_17761);
or U18147 (N_18147,N_17806,N_17568);
or U18148 (N_18148,N_17957,N_16063);
or U18149 (N_18149,N_17858,N_16390);
and U18150 (N_18150,N_16882,N_17770);
xor U18151 (N_18151,N_17638,N_16766);
nor U18152 (N_18152,N_16691,N_16689);
and U18153 (N_18153,N_17920,N_17910);
and U18154 (N_18154,N_17522,N_17915);
or U18155 (N_18155,N_17025,N_17953);
nand U18156 (N_18156,N_16450,N_16532);
or U18157 (N_18157,N_17101,N_17755);
nor U18158 (N_18158,N_16654,N_16456);
or U18159 (N_18159,N_17105,N_16483);
or U18160 (N_18160,N_16468,N_17267);
or U18161 (N_18161,N_17486,N_17881);
nor U18162 (N_18162,N_17153,N_16574);
nor U18163 (N_18163,N_16015,N_16756);
or U18164 (N_18164,N_17111,N_17188);
nand U18165 (N_18165,N_17283,N_16580);
and U18166 (N_18166,N_17298,N_17215);
nand U18167 (N_18167,N_17853,N_17474);
and U18168 (N_18168,N_17808,N_17639);
nor U18169 (N_18169,N_17297,N_17637);
nor U18170 (N_18170,N_16071,N_17288);
and U18171 (N_18171,N_16930,N_17338);
nand U18172 (N_18172,N_17524,N_16294);
or U18173 (N_18173,N_16757,N_16774);
nor U18174 (N_18174,N_16072,N_16230);
nor U18175 (N_18175,N_16191,N_17150);
nand U18176 (N_18176,N_16372,N_17501);
nor U18177 (N_18177,N_17660,N_17065);
or U18178 (N_18178,N_17232,N_17158);
nand U18179 (N_18179,N_16183,N_17337);
nor U18180 (N_18180,N_16344,N_17867);
or U18181 (N_18181,N_17537,N_16872);
or U18182 (N_18182,N_16245,N_16186);
or U18183 (N_18183,N_17842,N_17266);
and U18184 (N_18184,N_17716,N_16444);
and U18185 (N_18185,N_17406,N_16541);
nor U18186 (N_18186,N_17973,N_17926);
or U18187 (N_18187,N_17933,N_17480);
and U18188 (N_18188,N_16193,N_17705);
xnor U18189 (N_18189,N_16335,N_17516);
or U18190 (N_18190,N_16993,N_16043);
and U18191 (N_18191,N_16557,N_17694);
nor U18192 (N_18192,N_16296,N_17332);
xnor U18193 (N_18193,N_16395,N_16695);
or U18194 (N_18194,N_16270,N_17145);
or U18195 (N_18195,N_16844,N_17590);
nor U18196 (N_18196,N_17013,N_16740);
and U18197 (N_18197,N_17774,N_17361);
nand U18198 (N_18198,N_17747,N_16475);
nor U18199 (N_18199,N_16587,N_17316);
and U18200 (N_18200,N_16871,N_17342);
and U18201 (N_18201,N_16900,N_16272);
nand U18202 (N_18202,N_16777,N_17343);
or U18203 (N_18203,N_17087,N_17142);
and U18204 (N_18204,N_17156,N_16274);
xnor U18205 (N_18205,N_16565,N_17737);
nor U18206 (N_18206,N_17848,N_16105);
xor U18207 (N_18207,N_17578,N_16368);
nand U18208 (N_18208,N_17899,N_16685);
and U18209 (N_18209,N_17697,N_17659);
or U18210 (N_18210,N_17311,N_16712);
nor U18211 (N_18211,N_17003,N_17781);
and U18212 (N_18212,N_16798,N_17830);
nor U18213 (N_18213,N_17129,N_17802);
and U18214 (N_18214,N_16403,N_16657);
nor U18215 (N_18215,N_17666,N_16566);
or U18216 (N_18216,N_16062,N_16160);
and U18217 (N_18217,N_17086,N_17743);
and U18218 (N_18218,N_16509,N_16137);
nand U18219 (N_18219,N_17036,N_16760);
nor U18220 (N_18220,N_16935,N_16687);
nand U18221 (N_18221,N_16793,N_17347);
or U18222 (N_18222,N_16257,N_17890);
or U18223 (N_18223,N_16568,N_17477);
xnor U18224 (N_18224,N_17591,N_16316);
nand U18225 (N_18225,N_17681,N_17531);
nor U18226 (N_18226,N_16400,N_17099);
nor U18227 (N_18227,N_17108,N_16377);
nand U18228 (N_18228,N_16494,N_16861);
or U18229 (N_18229,N_17061,N_16251);
nor U18230 (N_18230,N_17670,N_16815);
xor U18231 (N_18231,N_17440,N_17898);
nand U18232 (N_18232,N_17614,N_16970);
nand U18233 (N_18233,N_17506,N_16491);
or U18234 (N_18234,N_17633,N_17725);
and U18235 (N_18235,N_17054,N_16964);
nor U18236 (N_18236,N_16214,N_16421);
xor U18237 (N_18237,N_17914,N_16873);
and U18238 (N_18238,N_16441,N_16538);
and U18239 (N_18239,N_16807,N_16847);
xnor U18240 (N_18240,N_17683,N_17244);
and U18241 (N_18241,N_17829,N_16868);
xor U18242 (N_18242,N_17002,N_17435);
nor U18243 (N_18243,N_16402,N_17149);
xnor U18244 (N_18244,N_16291,N_17907);
nand U18245 (N_18245,N_16755,N_16630);
nand U18246 (N_18246,N_16640,N_16026);
or U18247 (N_18247,N_16639,N_16613);
and U18248 (N_18248,N_17428,N_17059);
nor U18249 (N_18249,N_17541,N_16265);
or U18250 (N_18250,N_16535,N_17586);
xor U18251 (N_18251,N_16531,N_17859);
nor U18252 (N_18252,N_17535,N_17515);
nor U18253 (N_18253,N_17741,N_16481);
xnor U18254 (N_18254,N_17878,N_17596);
nand U18255 (N_18255,N_16748,N_17947);
xor U18256 (N_18256,N_16651,N_17151);
or U18257 (N_18257,N_17366,N_17676);
xor U18258 (N_18258,N_16721,N_16463);
nor U18259 (N_18259,N_17429,N_16162);
or U18260 (N_18260,N_16332,N_17478);
xnor U18261 (N_18261,N_16901,N_16473);
nand U18262 (N_18262,N_17056,N_16076);
and U18263 (N_18263,N_17554,N_16381);
nand U18264 (N_18264,N_17648,N_16300);
nor U18265 (N_18265,N_17465,N_17387);
and U18266 (N_18266,N_16744,N_17897);
nand U18267 (N_18267,N_16563,N_17612);
nand U18268 (N_18268,N_17033,N_16889);
nand U18269 (N_18269,N_17466,N_17321);
or U18270 (N_18270,N_16439,N_17895);
nand U18271 (N_18271,N_16152,N_16464);
nor U18272 (N_18272,N_16467,N_16813);
and U18273 (N_18273,N_17582,N_17130);
xor U18274 (N_18274,N_17828,N_17028);
nand U18275 (N_18275,N_17784,N_17679);
and U18276 (N_18276,N_17623,N_17324);
nor U18277 (N_18277,N_17044,N_17511);
nor U18278 (N_18278,N_16876,N_16242);
and U18279 (N_18279,N_17923,N_17669);
nor U18280 (N_18280,N_16146,N_17481);
nand U18281 (N_18281,N_17869,N_17967);
or U18282 (N_18282,N_17775,N_17595);
or U18283 (N_18283,N_16020,N_16008);
nor U18284 (N_18284,N_17326,N_16396);
or U18285 (N_18285,N_17179,N_17714);
or U18286 (N_18286,N_17320,N_16479);
nor U18287 (N_18287,N_17989,N_17498);
nand U18288 (N_18288,N_16553,N_16711);
nand U18289 (N_18289,N_16220,N_17984);
xor U18290 (N_18290,N_16578,N_16156);
xor U18291 (N_18291,N_17846,N_16644);
and U18292 (N_18292,N_17237,N_16921);
nor U18293 (N_18293,N_16413,N_16180);
and U18294 (N_18294,N_16004,N_16837);
and U18295 (N_18295,N_16933,N_16597);
xnor U18296 (N_18296,N_16855,N_16348);
and U18297 (N_18297,N_17969,N_17909);
nand U18298 (N_18298,N_16809,N_17529);
nand U18299 (N_18299,N_17097,N_17308);
xnor U18300 (N_18300,N_16998,N_17247);
nand U18301 (N_18301,N_16702,N_17490);
nor U18302 (N_18302,N_16931,N_16646);
xnor U18303 (N_18303,N_17976,N_16739);
and U18304 (N_18304,N_16111,N_16869);
nand U18305 (N_18305,N_16934,N_16482);
nand U18306 (N_18306,N_16703,N_16069);
nand U18307 (N_18307,N_17363,N_17937);
nor U18308 (N_18308,N_16132,N_16607);
or U18309 (N_18309,N_17000,N_17916);
or U18310 (N_18310,N_17667,N_17075);
or U18311 (N_18311,N_16174,N_17147);
nor U18312 (N_18312,N_17174,N_16330);
and U18313 (N_18313,N_17675,N_16313);
nand U18314 (N_18314,N_16514,N_17814);
or U18315 (N_18315,N_17852,N_16910);
nor U18316 (N_18316,N_17505,N_17572);
or U18317 (N_18317,N_17854,N_16719);
nand U18318 (N_18318,N_16139,N_17467);
nand U18319 (N_18319,N_16264,N_16612);
or U18320 (N_18320,N_16981,N_17323);
xnor U18321 (N_18321,N_17255,N_17208);
and U18322 (N_18322,N_17005,N_16641);
xnor U18323 (N_18323,N_16319,N_17488);
nor U18324 (N_18324,N_16500,N_17252);
or U18325 (N_18325,N_17305,N_17095);
nor U18326 (N_18326,N_16024,N_17791);
nand U18327 (N_18327,N_16547,N_17396);
nor U18328 (N_18328,N_17994,N_16655);
xnor U18329 (N_18329,N_16415,N_17520);
or U18330 (N_18330,N_17074,N_17348);
nand U18331 (N_18331,N_17487,N_17550);
nand U18332 (N_18332,N_16369,N_17685);
nor U18333 (N_18333,N_17952,N_16893);
and U18334 (N_18334,N_16851,N_16902);
nand U18335 (N_18335,N_17664,N_16692);
nor U18336 (N_18336,N_17936,N_16885);
or U18337 (N_18337,N_16818,N_16600);
or U18338 (N_18338,N_17930,N_16027);
or U18339 (N_18339,N_17204,N_16658);
nor U18340 (N_18340,N_16309,N_17442);
and U18341 (N_18341,N_16536,N_17922);
and U18342 (N_18342,N_17325,N_16434);
xor U18343 (N_18343,N_16779,N_17655);
and U18344 (N_18344,N_17415,N_16005);
nor U18345 (N_18345,N_17225,N_17300);
nand U18346 (N_18346,N_17945,N_16207);
nor U18347 (N_18347,N_17606,N_16735);
or U18348 (N_18348,N_17615,N_16411);
nand U18349 (N_18349,N_16710,N_17341);
and U18350 (N_18350,N_17140,N_17496);
nor U18351 (N_18351,N_16347,N_16098);
or U18352 (N_18352,N_16324,N_16073);
nor U18353 (N_18353,N_17189,N_16290);
and U18354 (N_18354,N_16086,N_17278);
xor U18355 (N_18355,N_17497,N_16345);
xor U18356 (N_18356,N_17089,N_16932);
or U18357 (N_18357,N_17289,N_17152);
nand U18358 (N_18358,N_17772,N_17251);
xnor U18359 (N_18359,N_17837,N_17403);
xnor U18360 (N_18360,N_17924,N_17339);
xnor U18361 (N_18361,N_17157,N_16386);
or U18362 (N_18362,N_17523,N_17602);
nand U18363 (N_18363,N_17768,N_16364);
xnor U18364 (N_18364,N_17840,N_16065);
nand U18365 (N_18365,N_16077,N_16716);
or U18366 (N_18366,N_17888,N_17500);
nand U18367 (N_18367,N_16116,N_17407);
nand U18368 (N_18368,N_17131,N_17100);
xor U18369 (N_18369,N_16349,N_17992);
nor U18370 (N_18370,N_17731,N_16584);
nand U18371 (N_18371,N_16895,N_17722);
and U18372 (N_18372,N_16064,N_17192);
or U18373 (N_18373,N_17029,N_17450);
nor U18374 (N_18374,N_17183,N_16233);
nor U18375 (N_18375,N_17730,N_16244);
xor U18376 (N_18376,N_17085,N_16824);
nand U18377 (N_18377,N_16133,N_16157);
nand U18378 (N_18378,N_17078,N_16800);
nor U18379 (N_18379,N_17281,N_16185);
and U18380 (N_18380,N_16425,N_17734);
nor U18381 (N_18381,N_16458,N_16454);
nand U18382 (N_18382,N_16986,N_17999);
nand U18383 (N_18383,N_16810,N_16629);
nand U18384 (N_18384,N_17636,N_17397);
or U18385 (N_18385,N_17102,N_17303);
nand U18386 (N_18386,N_17729,N_16447);
nor U18387 (N_18387,N_16814,N_17793);
and U18388 (N_18388,N_17294,N_17438);
nor U18389 (N_18389,N_16283,N_16356);
nand U18390 (N_18390,N_16266,N_17692);
nor U18391 (N_18391,N_16789,N_16821);
xor U18392 (N_18392,N_17035,N_17336);
or U18393 (N_18393,N_16874,N_16195);
nand U18394 (N_18394,N_16544,N_16788);
and U18395 (N_18395,N_16884,N_17409);
or U18396 (N_18396,N_16564,N_17136);
xnor U18397 (N_18397,N_16223,N_16228);
nand U18398 (N_18398,N_16163,N_17845);
xnor U18399 (N_18399,N_17046,N_17635);
or U18400 (N_18400,N_16853,N_16241);
and U18401 (N_18401,N_16199,N_16379);
and U18402 (N_18402,N_16360,N_16854);
and U18403 (N_18403,N_17448,N_17053);
nor U18404 (N_18404,N_17287,N_17049);
nand U18405 (N_18405,N_16690,N_16341);
nor U18406 (N_18406,N_16560,N_17318);
nor U18407 (N_18407,N_16023,N_16224);
nand U18408 (N_18408,N_16151,N_17941);
or U18409 (N_18409,N_17820,N_17780);
and U18410 (N_18410,N_16585,N_16082);
xor U18411 (N_18411,N_17489,N_16124);
nand U18412 (N_18412,N_16340,N_17121);
nor U18413 (N_18413,N_16250,N_17401);
or U18414 (N_18414,N_17356,N_17626);
nor U18415 (N_18415,N_16674,N_17621);
or U18416 (N_18416,N_16145,N_17205);
nor U18417 (N_18417,N_16526,N_16696);
xor U18418 (N_18418,N_16032,N_16429);
or U18419 (N_18419,N_17677,N_16169);
xor U18420 (N_18420,N_16598,N_17452);
and U18421 (N_18421,N_17826,N_17106);
or U18422 (N_18422,N_16326,N_17700);
or U18423 (N_18423,N_16212,N_16351);
nor U18424 (N_18424,N_16061,N_17744);
and U18425 (N_18425,N_16941,N_17695);
and U18426 (N_18426,N_16058,N_16167);
xnor U18427 (N_18427,N_17217,N_16795);
and U18428 (N_18428,N_17172,N_16924);
nand U18429 (N_18429,N_16991,N_16471);
xnor U18430 (N_18430,N_16019,N_17870);
or U18431 (N_18431,N_16198,N_16787);
nor U18432 (N_18432,N_17264,N_16325);
and U18433 (N_18433,N_17126,N_16904);
nand U18434 (N_18434,N_16030,N_16052);
nor U18435 (N_18435,N_16120,N_17576);
or U18436 (N_18436,N_17902,N_17368);
or U18437 (N_18437,N_16953,N_16911);
nor U18438 (N_18438,N_17649,N_17276);
nand U18439 (N_18439,N_16289,N_16828);
nand U18440 (N_18440,N_16457,N_16496);
nand U18441 (N_18441,N_16256,N_16206);
and U18442 (N_18442,N_16219,N_16187);
nand U18443 (N_18443,N_17824,N_16610);
nor U18444 (N_18444,N_16263,N_16903);
nand U18445 (N_18445,N_16773,N_17797);
and U18446 (N_18446,N_16480,N_17763);
and U18447 (N_18447,N_17168,N_17657);
or U18448 (N_18448,N_16357,N_16864);
xnor U18449 (N_18449,N_17417,N_16525);
and U18450 (N_18450,N_17254,N_16260);
nand U18451 (N_18451,N_16617,N_16713);
and U18452 (N_18452,N_17471,N_17625);
nand U18453 (N_18453,N_16765,N_16142);
or U18454 (N_18454,N_17735,N_17350);
and U18455 (N_18455,N_16596,N_16476);
nor U18456 (N_18456,N_17068,N_16099);
or U18457 (N_18457,N_17581,N_16168);
nor U18458 (N_18458,N_16009,N_17605);
nor U18459 (N_18459,N_16656,N_17027);
and U18460 (N_18460,N_17080,N_17166);
nor U18461 (N_18461,N_16906,N_16684);
xor U18462 (N_18462,N_17349,N_17260);
nand U18463 (N_18463,N_17258,N_17998);
or U18464 (N_18464,N_16196,N_16367);
and U18465 (N_18465,N_16165,N_17528);
and U18466 (N_18466,N_16172,N_17381);
or U18467 (N_18467,N_17222,N_16792);
nand U18468 (N_18468,N_16392,N_17850);
or U18469 (N_18469,N_17485,N_16006);
and U18470 (N_18470,N_16074,N_16865);
nor U18471 (N_18471,N_17887,N_17082);
or U18472 (N_18472,N_17391,N_16937);
or U18473 (N_18473,N_16427,N_16477);
nor U18474 (N_18474,N_17720,N_16555);
nor U18475 (N_18475,N_17178,N_17944);
nor U18476 (N_18476,N_16548,N_16249);
nand U18477 (N_18477,N_16182,N_17634);
or U18478 (N_18478,N_17132,N_16176);
and U18479 (N_18479,N_16550,N_17579);
nand U18480 (N_18480,N_16775,N_17825);
nor U18481 (N_18481,N_17161,N_16661);
and U18482 (N_18482,N_16841,N_16484);
xor U18483 (N_18483,N_16361,N_17037);
nor U18484 (N_18484,N_17518,N_17024);
xnor U18485 (N_18485,N_17834,N_17426);
and U18486 (N_18486,N_17167,N_16016);
xor U18487 (N_18487,N_17019,N_17611);
and U18488 (N_18488,N_17610,N_16181);
xor U18489 (N_18489,N_16963,N_17020);
or U18490 (N_18490,N_17399,N_16449);
and U18491 (N_18491,N_16539,N_17913);
nand U18492 (N_18492,N_16753,N_17929);
xor U18493 (N_18493,N_17390,N_17274);
nand U18494 (N_18494,N_16575,N_17841);
nor U18495 (N_18495,N_16383,N_17042);
and U18496 (N_18496,N_16398,N_16511);
or U18497 (N_18497,N_17862,N_17833);
or U18498 (N_18498,N_16331,N_17645);
nor U18499 (N_18499,N_16778,N_16401);
nor U18500 (N_18500,N_16913,N_16374);
nand U18501 (N_18501,N_17411,N_17795);
xnor U18502 (N_18502,N_17062,N_16067);
and U18503 (N_18503,N_17010,N_16229);
nand U18504 (N_18504,N_16973,N_17016);
xnor U18505 (N_18505,N_16916,N_16923);
nor U18506 (N_18506,N_16768,N_17202);
nor U18507 (N_18507,N_17169,N_16977);
and U18508 (N_18508,N_16431,N_16147);
and U18509 (N_18509,N_16358,N_17642);
nand U18510 (N_18510,N_17709,N_17652);
and U18511 (N_18511,N_16042,N_17094);
nand U18512 (N_18512,N_17272,N_17170);
or U18513 (N_18513,N_16259,N_16772);
or U18514 (N_18514,N_16611,N_17098);
and U18515 (N_18515,N_16307,N_17476);
and U18516 (N_18516,N_17921,N_17249);
or U18517 (N_18517,N_16267,N_16524);
or U18518 (N_18518,N_16155,N_16025);
or U18519 (N_18519,N_16149,N_16638);
or U18520 (N_18520,N_16870,N_16310);
or U18521 (N_18521,N_16549,N_17394);
nand U18522 (N_18522,N_17446,N_16801);
nand U18523 (N_18523,N_16840,N_17732);
nor U18524 (N_18524,N_17879,N_17974);
or U18525 (N_18525,N_17299,N_16938);
nand U18526 (N_18526,N_17026,N_17201);
and U18527 (N_18527,N_17413,N_17119);
or U18528 (N_18528,N_17958,N_17564);
or U18529 (N_18529,N_16594,N_17367);
or U18530 (N_18530,N_17220,N_16846);
or U18531 (N_18531,N_17987,N_16718);
or U18532 (N_18532,N_17414,N_16816);
nor U18533 (N_18533,N_17599,N_17661);
or U18534 (N_18534,N_16096,N_16359);
and U18535 (N_18535,N_17384,N_16699);
and U18536 (N_18536,N_16725,N_17963);
nor U18537 (N_18537,N_17577,N_17985);
and U18538 (N_18538,N_16127,N_16164);
or U18539 (N_18539,N_17370,N_17454);
and U18540 (N_18540,N_16338,N_16436);
or U18541 (N_18541,N_17589,N_17587);
nand U18542 (N_18542,N_17022,N_17491);
or U18543 (N_18543,N_17777,N_17373);
nand U18544 (N_18544,N_16045,N_16586);
or U18545 (N_18545,N_16079,N_16722);
nor U18546 (N_18546,N_17656,N_16134);
or U18547 (N_18547,N_16592,N_16232);
nand U18548 (N_18548,N_17083,N_16635);
nand U18549 (N_18549,N_16175,N_17443);
nor U18550 (N_18550,N_16733,N_17547);
and U18551 (N_18551,N_16208,N_16985);
or U18552 (N_18552,N_17889,N_16097);
nand U18553 (N_18553,N_16781,N_16432);
nor U18554 (N_18554,N_16754,N_17548);
nand U18555 (N_18555,N_16959,N_16090);
nor U18556 (N_18556,N_17090,N_16171);
or U18557 (N_18557,N_16410,N_17792);
and U18558 (N_18558,N_17643,N_16093);
and U18559 (N_18559,N_16297,N_17425);
nand U18560 (N_18560,N_16424,N_16730);
nand U18561 (N_18561,N_17618,N_17960);
nand U18562 (N_18562,N_17964,N_16771);
or U18563 (N_18563,N_17461,N_16936);
xnor U18564 (N_18564,N_16960,N_17684);
nand U18565 (N_18565,N_17253,N_16738);
and U18566 (N_18566,N_16672,N_17280);
nand U18567 (N_18567,N_17510,N_16057);
nor U18568 (N_18568,N_17726,N_16749);
nand U18569 (N_18569,N_16742,N_16273);
or U18570 (N_18570,N_17647,N_16825);
nand U18571 (N_18571,N_16826,N_16955);
or U18572 (N_18572,N_17710,N_17533);
or U18573 (N_18573,N_16677,N_16551);
or U18574 (N_18574,N_16627,N_16762);
xor U18575 (N_18575,N_17434,N_16227);
and U18576 (N_18576,N_17047,N_17884);
or U18577 (N_18577,N_17632,N_17122);
and U18578 (N_18578,N_16302,N_16767);
or U18579 (N_18579,N_16138,N_17069);
and U18580 (N_18580,N_16334,N_17227);
nand U18581 (N_18581,N_16321,N_16092);
and U18582 (N_18582,N_16159,N_17712);
or U18583 (N_18583,N_17301,N_16237);
nand U18584 (N_18584,N_16875,N_17405);
nand U18585 (N_18585,N_17051,N_16000);
and U18586 (N_18586,N_17001,N_17688);
or U18587 (N_18587,N_17213,N_16537);
and U18588 (N_18588,N_17239,N_16033);
nor U18589 (N_18589,N_16676,N_17436);
nor U18590 (N_18590,N_16673,N_16501);
nor U18591 (N_18591,N_16817,N_16059);
or U18592 (N_18592,N_17750,N_17641);
nand U18593 (N_18593,N_16118,N_16204);
and U18594 (N_18594,N_17882,N_16602);
or U18595 (N_18595,N_16850,N_16764);
nor U18596 (N_18596,N_17352,N_16704);
and U18597 (N_18597,N_16279,N_17420);
and U18598 (N_18598,N_17903,N_17110);
or U18599 (N_18599,N_17601,N_17766);
nor U18600 (N_18600,N_16899,N_16750);
xor U18601 (N_18601,N_16528,N_16849);
xnor U18602 (N_18602,N_17598,N_17271);
or U18603 (N_18603,N_16521,N_16243);
nand U18604 (N_18604,N_16013,N_17503);
nor U18605 (N_18605,N_16271,N_17091);
or U18606 (N_18606,N_17378,N_16866);
nor U18607 (N_18607,N_16478,N_17822);
xor U18608 (N_18608,N_17954,N_16782);
or U18609 (N_18609,N_17092,N_16011);
nand U18610 (N_18610,N_16670,N_16724);
or U18611 (N_18611,N_16085,N_17538);
and U18612 (N_18612,N_16423,N_16533);
nand U18613 (N_18613,N_16018,N_17482);
and U18614 (N_18614,N_17749,N_16512);
nand U18615 (N_18615,N_17724,N_17453);
or U18616 (N_18616,N_17479,N_16306);
and U18617 (N_18617,N_17717,N_16616);
nand U18618 (N_18618,N_16679,N_17512);
nor U18619 (N_18619,N_17449,N_17549);
and U18620 (N_18620,N_17751,N_17346);
and U18621 (N_18621,N_16577,N_16633);
nor U18622 (N_18622,N_16021,N_16517);
nor U18623 (N_18623,N_17187,N_17680);
xor U18624 (N_18624,N_17832,N_16091);
nor U18625 (N_18625,N_17234,N_16154);
xnor U18626 (N_18626,N_16590,N_16647);
xor U18627 (N_18627,N_17757,N_17650);
nand U18628 (N_18628,N_16448,N_16522);
xnor U18629 (N_18629,N_16044,N_16675);
nor U18630 (N_18630,N_17573,N_17315);
or U18631 (N_18631,N_17671,N_16409);
xnor U18632 (N_18632,N_17603,N_17779);
xnor U18633 (N_18633,N_17270,N_17925);
xor U18634 (N_18634,N_16897,N_17295);
and U18635 (N_18635,N_17736,N_17277);
nand U18636 (N_18636,N_16806,N_17463);
nor U18637 (N_18637,N_17455,N_17293);
xnor U18638 (N_18638,N_17296,N_17940);
nand U18639 (N_18639,N_17369,N_16908);
or U18640 (N_18640,N_16083,N_17687);
nand U18641 (N_18641,N_17160,N_16365);
and U18642 (N_18642,N_16100,N_17354);
xnor U18643 (N_18643,N_17962,N_16125);
and U18644 (N_18644,N_17462,N_16928);
and U18645 (N_18645,N_17408,N_16487);
nand U18646 (N_18646,N_16417,N_17223);
and U18647 (N_18647,N_16278,N_17388);
and U18648 (N_18648,N_16506,N_16126);
and U18649 (N_18649,N_16796,N_16746);
or U18650 (N_18650,N_16068,N_16299);
nor U18651 (N_18651,N_16508,N_16363);
or U18652 (N_18652,N_17765,N_17176);
nand U18653 (N_18653,N_17935,N_17400);
or U18654 (N_18654,N_16502,N_17758);
and U18655 (N_18655,N_16261,N_16315);
or U18656 (N_18656,N_16982,N_16110);
nor U18657 (N_18657,N_17526,N_17836);
or U18658 (N_18658,N_16226,N_16678);
and U18659 (N_18659,N_17040,N_17872);
nor U18660 (N_18660,N_17275,N_17226);
nand U18661 (N_18661,N_17031,N_16576);
or U18662 (N_18662,N_16393,N_17457);
or U18663 (N_18663,N_16136,N_16102);
or U18664 (N_18664,N_17979,N_16275);
nand U18665 (N_18665,N_17379,N_16465);
or U18666 (N_18666,N_17230,N_17114);
xor U18667 (N_18667,N_16650,N_16388);
xor U18668 (N_18668,N_16247,N_17052);
nand U18669 (N_18669,N_16665,N_16983);
nand U18670 (N_18670,N_17557,N_17460);
nand U18671 (N_18671,N_16412,N_16618);
nor U18672 (N_18672,N_17978,N_17622);
nand U18673 (N_18673,N_17331,N_17785);
nor U18674 (N_18674,N_17996,N_17919);
nor U18675 (N_18675,N_16708,N_17783);
and U18676 (N_18676,N_16726,N_16571);
or U18677 (N_18677,N_16967,N_17335);
and U18678 (N_18678,N_17144,N_17574);
xor U18679 (N_18679,N_16942,N_16327);
nor U18680 (N_18680,N_17050,N_16599);
xor U18681 (N_18681,N_17439,N_16007);
or U18682 (N_18682,N_16014,N_17521);
xor U18683 (N_18683,N_16070,N_16845);
nand U18684 (N_18684,N_17892,N_16892);
or U18685 (N_18685,N_17359,N_16095);
nand U18686 (N_18686,N_16919,N_17193);
and U18687 (N_18687,N_17875,N_16170);
and U18688 (N_18688,N_17555,N_17197);
nand U18689 (N_18689,N_16636,N_17819);
nor U18690 (N_18690,N_16087,N_16857);
or U18691 (N_18691,N_17558,N_16108);
nor U18692 (N_18692,N_16179,N_17682);
nor U18693 (N_18693,N_16318,N_16109);
or U18694 (N_18694,N_16709,N_17708);
or U18695 (N_18695,N_16231,N_16802);
or U18696 (N_18696,N_16623,N_16682);
or U18697 (N_18697,N_16527,N_16763);
nand U18698 (N_18698,N_16579,N_16615);
nand U18699 (N_18699,N_16907,N_17398);
nand U18700 (N_18700,N_17057,N_17701);
nor U18701 (N_18701,N_16197,N_17392);
nand U18702 (N_18702,N_17986,N_16455);
and U18703 (N_18703,N_16920,N_17306);
and U18704 (N_18704,N_17334,N_16437);
and U18705 (N_18705,N_16939,N_17778);
or U18706 (N_18706,N_16561,N_17304);
and U18707 (N_18707,N_16625,N_16582);
and U18708 (N_18708,N_17128,N_17345);
nor U18709 (N_18709,N_17292,N_17117);
and U18710 (N_18710,N_17988,N_16799);
and U18711 (N_18711,N_17084,N_16791);
nor U18712 (N_18712,N_16879,N_17214);
or U18713 (N_18713,N_16305,N_17259);
or U18714 (N_18714,N_17096,N_16416);
nor U18715 (N_18715,N_16642,N_16648);
and U18716 (N_18716,N_16375,N_17246);
and U18717 (N_18717,N_16589,N_17982);
and U18718 (N_18718,N_16202,N_17115);
nor U18719 (N_18719,N_16971,N_17256);
and U18720 (N_18720,N_17653,N_17048);
nand U18721 (N_18721,N_17876,N_16925);
nor U18722 (N_18722,N_16298,N_17698);
or U18723 (N_18723,N_17948,N_16649);
nor U18724 (N_18724,N_16066,N_16515);
nand U18725 (N_18725,N_16003,N_16459);
or U18726 (N_18726,N_17164,N_17803);
or U18727 (N_18727,N_16135,N_16785);
nand U18728 (N_18728,N_17066,N_16859);
nand U18729 (N_18729,N_17600,N_16829);
nor U18730 (N_18730,N_16940,N_16001);
xor U18731 (N_18731,N_17807,N_17328);
xnor U18732 (N_18732,N_17629,N_17072);
nand U18733 (N_18733,N_17393,N_16081);
nor U18734 (N_18734,N_17198,N_16215);
nor U18735 (N_18735,N_17739,N_17776);
nand U18736 (N_18736,N_16002,N_16028);
nand U18737 (N_18737,N_16201,N_17658);
nor U18738 (N_18738,N_16405,N_17199);
and U18739 (N_18739,N_17279,N_17317);
or U18740 (N_18740,N_17383,N_16686);
nor U18741 (N_18741,N_17133,N_17727);
and U18742 (N_18742,N_17322,N_17360);
and U18743 (N_18743,N_17917,N_17265);
xnor U18744 (N_18744,N_16980,N_16833);
or U18745 (N_18745,N_17362,N_16084);
nand U18746 (N_18746,N_16397,N_17107);
nand U18747 (N_18747,N_16698,N_16784);
nand U18748 (N_18748,N_17207,N_16225);
or U18749 (N_18749,N_16445,N_17423);
nor U18750 (N_18750,N_17219,N_17900);
and U18751 (N_18751,N_17262,N_16917);
or U18752 (N_18752,N_16632,N_16662);
nor U18753 (N_18753,N_16808,N_16737);
or U18754 (N_18754,N_17672,N_16284);
and U18755 (N_18755,N_16440,N_17844);
nor U18756 (N_18756,N_16680,N_17030);
nor U18757 (N_18757,N_17760,N_17310);
and U18758 (N_18758,N_17211,N_17561);
nor U18759 (N_18759,N_17137,N_16323);
and U18760 (N_18760,N_16088,N_17196);
or U18761 (N_18761,N_16046,N_17127);
or U18762 (N_18762,N_16328,N_17759);
or U18763 (N_18763,N_17813,N_16505);
or U18764 (N_18764,N_16994,N_17070);
nand U18765 (N_18765,N_16217,N_16486);
nand U18766 (N_18766,N_16706,N_17536);
nor U18767 (N_18767,N_16780,N_16286);
or U18768 (N_18768,N_17307,N_16103);
and U18769 (N_18769,N_17291,N_17686);
nor U18770 (N_18770,N_16581,N_16803);
nand U18771 (N_18771,N_16158,N_17868);
and U18772 (N_18772,N_16117,N_17319);
nor U18773 (N_18773,N_16843,N_17968);
nand U18774 (N_18774,N_17631,N_16422);
and U18775 (N_18775,N_17951,N_17173);
nand U18776 (N_18776,N_17206,N_17861);
nand U18777 (N_18777,N_17382,N_17965);
and U18778 (N_18778,N_17007,N_17008);
nor U18779 (N_18779,N_17620,N_17567);
and U18780 (N_18780,N_17104,N_16221);
nor U18781 (N_18781,N_16322,N_17410);
or U18782 (N_18782,N_17886,N_16075);
nand U18783 (N_18783,N_16017,N_16389);
nand U18784 (N_18784,N_17918,N_17143);
nand U18785 (N_18785,N_16927,N_16783);
or U18786 (N_18786,N_17790,N_17504);
nor U18787 (N_18787,N_17613,N_16943);
nor U18788 (N_18788,N_17950,N_16430);
or U18789 (N_18789,N_16572,N_16860);
or U18790 (N_18790,N_16681,N_17855);
xnor U18791 (N_18791,N_16958,N_17039);
or U18792 (N_18792,N_17433,N_16452);
or U18793 (N_18793,N_16770,N_16637);
nand U18794 (N_18794,N_17456,N_16350);
nand U18795 (N_18795,N_17901,N_17931);
nor U18796 (N_18796,N_17594,N_16451);
xor U18797 (N_18797,N_17551,N_17866);
nand U18798 (N_18798,N_16988,N_16890);
nand U18799 (N_18799,N_16418,N_17118);
nor U18800 (N_18800,N_16101,N_17961);
xnor U18801 (N_18801,N_16446,N_16700);
xor U18802 (N_18802,N_17733,N_16717);
nand U18803 (N_18803,N_17514,N_17809);
nand U18804 (N_18804,N_16761,N_17835);
or U18805 (N_18805,N_16060,N_16848);
or U18806 (N_18806,N_17570,N_17374);
or U18807 (N_18807,N_17257,N_16823);
nand U18808 (N_18808,N_17451,N_16173);
and U18809 (N_18809,N_17838,N_16384);
nor U18810 (N_18810,N_17045,N_16688);
nor U18811 (N_18811,N_17402,N_16752);
nand U18812 (N_18812,N_17971,N_16534);
or U18813 (N_18813,N_16442,N_16836);
and U18814 (N_18814,N_16573,N_17216);
nand U18815 (N_18815,N_16945,N_16276);
nor U18816 (N_18816,N_16376,N_16293);
nand U18817 (N_18817,N_17469,N_17242);
nand U18818 (N_18818,N_17041,N_16407);
nor U18819 (N_18819,N_16956,N_17380);
nand U18820 (N_18820,N_16041,N_17495);
or U18821 (N_18821,N_17493,N_16758);
nand U18822 (N_18822,N_17546,N_16554);
xor U18823 (N_18823,N_17946,N_17552);
nor U18824 (N_18824,N_16951,N_16371);
nor U18825 (N_18825,N_17492,N_17788);
nor U18826 (N_18826,N_16558,N_16604);
nor U18827 (N_18827,N_17527,N_16631);
xnor U18828 (N_18828,N_17139,N_16419);
and U18829 (N_18829,N_16503,N_16239);
nor U18830 (N_18830,N_17894,N_16253);
xnor U18831 (N_18831,N_16888,N_17860);
nand U18832 (N_18832,N_16569,N_17756);
and U18833 (N_18833,N_16894,N_16831);
or U18834 (N_18834,N_17604,N_16603);
nand U18835 (N_18835,N_17221,N_16255);
nand U18836 (N_18836,N_17412,N_17851);
nor U18837 (N_18837,N_17588,N_17748);
or U18838 (N_18838,N_17385,N_17229);
nor U18839 (N_18839,N_17880,N_16729);
nand U18840 (N_18840,N_17344,N_17175);
and U18841 (N_18841,N_17468,N_17762);
nand U18842 (N_18842,N_16835,N_16203);
or U18843 (N_18843,N_17693,N_16957);
nand U18844 (N_18844,N_16177,N_16862);
nor U18845 (N_18845,N_17200,N_16056);
and U18846 (N_18846,N_17871,N_17430);
xnor U18847 (N_18847,N_17995,N_17032);
xnor U18848 (N_18848,N_17422,N_17787);
nand U18849 (N_18849,N_17993,N_16643);
nand U18850 (N_18850,N_16747,N_16728);
nor U18851 (N_18851,N_17812,N_17250);
nor U18852 (N_18852,N_17715,N_16867);
or U18853 (N_18853,N_17789,N_17261);
nor U18854 (N_18854,N_17843,N_17376);
nor U18855 (N_18855,N_16830,N_16346);
nor U18856 (N_18856,N_17678,N_16128);
or U18857 (N_18857,N_17713,N_16811);
xor U18858 (N_18858,N_17155,N_16218);
and U18859 (N_18859,N_16929,N_17990);
and U18860 (N_18860,N_17719,N_16498);
nor U18861 (N_18861,N_16122,N_17180);
xnor U18862 (N_18862,N_16608,N_17231);
nand U18863 (N_18863,N_16472,N_16992);
nand U18864 (N_18864,N_17241,N_17269);
nand U18865 (N_18865,N_17773,N_16723);
nand U18866 (N_18866,N_17148,N_16881);
nand U18867 (N_18867,N_17171,N_17810);
and U18868 (N_18868,N_16150,N_16671);
or U18869 (N_18869,N_17630,N_17742);
nor U18870 (N_18870,N_17972,N_16200);
or U18871 (N_18871,N_16317,N_16050);
xor U18872 (N_18872,N_16131,N_17771);
xor U18873 (N_18873,N_16269,N_17159);
nor U18874 (N_18874,N_17949,N_16667);
and U18875 (N_18875,N_16731,N_16038);
nor U18876 (N_18876,N_17499,N_17228);
xnor U18877 (N_18877,N_16387,N_17811);
nand U18878 (N_18878,N_17483,N_17093);
nor U18879 (N_18879,N_16153,N_17804);
nor U18880 (N_18880,N_17544,N_17977);
nand U18881 (N_18881,N_16653,N_17646);
nor U18882 (N_18882,N_16262,N_17718);
nor U18883 (N_18883,N_16339,N_16497);
nand U18884 (N_18884,N_16880,N_17067);
nand U18885 (N_18885,N_16246,N_16312);
nand U18886 (N_18886,N_16130,N_16975);
or U18887 (N_18887,N_16645,N_17416);
or U18888 (N_18888,N_16495,N_17818);
nor U18889 (N_18889,N_16887,N_16285);
or U18890 (N_18890,N_17210,N_17746);
and U18891 (N_18891,N_17942,N_17079);
nor U18892 (N_18892,N_17654,N_17377);
xor U18893 (N_18893,N_16234,N_17038);
nand U18894 (N_18894,N_17938,N_17286);
nor U18895 (N_18895,N_16012,N_17975);
or U18896 (N_18896,N_16743,N_17556);
nand U18897 (N_18897,N_16408,N_17445);
or U18898 (N_18898,N_16304,N_16595);
nor U18899 (N_18899,N_16031,N_17519);
nor U18900 (N_18900,N_16540,N_16391);
nand U18901 (N_18901,N_17134,N_16029);
nor U18902 (N_18902,N_17458,N_16896);
nand U18903 (N_18903,N_16040,N_16314);
xnor U18904 (N_18904,N_16094,N_17235);
nor U18905 (N_18905,N_17896,N_17839);
nand U18906 (N_18906,N_16433,N_16462);
or U18907 (N_18907,N_17125,N_16614);
nand U18908 (N_18908,N_16559,N_16268);
or U18909 (N_18909,N_16010,N_16922);
nor U18910 (N_18910,N_17182,N_16519);
and U18911 (N_18911,N_16562,N_17644);
xnor U18912 (N_18912,N_16542,N_16210);
or U18913 (N_18913,N_17419,N_17904);
nand U18914 (N_18914,N_17088,N_16666);
xor U18915 (N_18915,N_16812,N_17997);
or U18916 (N_18916,N_17891,N_17141);
nor U18917 (N_18917,N_17593,N_17569);
and U18918 (N_18918,N_16858,N_16258);
nor U18919 (N_18919,N_16918,N_17563);
nor U18920 (N_18920,N_16878,N_17566);
or U18921 (N_18921,N_17018,N_17212);
and U18922 (N_18922,N_17706,N_16999);
nor U18923 (N_18923,N_17081,N_17502);
nand U18924 (N_18924,N_17662,N_17905);
and U18925 (N_18925,N_16295,N_17431);
nand U18926 (N_18926,N_16732,N_16362);
nand U18927 (N_18927,N_16443,N_17885);
nor U18928 (N_18928,N_16989,N_17177);
xor U18929 (N_18929,N_17959,N_17592);
and U18930 (N_18930,N_17764,N_16997);
or U18931 (N_18931,N_16460,N_16621);
and U18932 (N_18932,N_16353,N_16178);
nand U18933 (N_18933,N_17203,N_16660);
nand U18934 (N_18934,N_17823,N_16839);
nor U18935 (N_18935,N_16488,N_17627);
or U18936 (N_18936,N_17063,N_17562);
or U18937 (N_18937,N_17470,N_17109);
nand U18938 (N_18938,N_17821,N_16303);
nand U18939 (N_18939,N_16786,N_16693);
nand U18940 (N_18940,N_16820,N_16343);
nor U18941 (N_18941,N_17351,N_16129);
and U18942 (N_18942,N_16545,N_16987);
and U18943 (N_18943,N_17545,N_17494);
nand U18944 (N_18944,N_16518,N_17575);
nand U18945 (N_18945,N_17421,N_17607);
nand U18946 (N_18946,N_17934,N_17012);
or U18947 (N_18947,N_17389,N_16474);
or U18948 (N_18948,N_17508,N_17651);
nor U18949 (N_18949,N_16466,N_16492);
nand U18950 (N_18950,N_16593,N_16588);
nand U18951 (N_18951,N_16504,N_16863);
nand U18952 (N_18952,N_16946,N_16701);
or U18953 (N_18953,N_17874,N_17691);
and U18954 (N_18954,N_17181,N_17186);
or U18955 (N_18955,N_17236,N_17690);
or U18956 (N_18956,N_16663,N_16626);
or U18957 (N_18957,N_17165,N_17542);
or U18958 (N_18958,N_17525,N_17711);
nor U18959 (N_18959,N_17800,N_17863);
nor U18960 (N_18960,N_16115,N_16311);
nand U18961 (N_18961,N_17799,N_17060);
nor U18962 (N_18962,N_17624,N_16886);
nand U18963 (N_18963,N_16751,N_16962);
nand U18964 (N_18964,N_16048,N_16282);
nor U18965 (N_18965,N_16905,N_16984);
nor U18966 (N_18966,N_17432,N_16420);
and U18967 (N_18967,N_16113,N_16209);
or U18968 (N_18968,N_16184,N_16856);
and U18969 (N_18969,N_16797,N_16453);
or U18970 (N_18970,N_17532,N_16248);
xnor U18971 (N_18971,N_17740,N_17475);
nand U18972 (N_18972,N_17263,N_17138);
nand U18973 (N_18973,N_17058,N_17877);
nand U18974 (N_18974,N_17559,N_16438);
and U18975 (N_18975,N_16035,N_17006);
or U18976 (N_18976,N_16948,N_17185);
or U18977 (N_18977,N_17444,N_17906);
nor U18978 (N_18978,N_16915,N_16720);
nand U18979 (N_18979,N_17728,N_16507);
or U18980 (N_18980,N_17240,N_16053);
and U18981 (N_18981,N_16493,N_17753);
nand U18982 (N_18982,N_17908,N_16516);
or U18983 (N_18983,N_17847,N_17355);
nor U18984 (N_18984,N_17798,N_16254);
nor U18985 (N_18985,N_16852,N_17329);
and U18986 (N_18986,N_16378,N_16216);
or U18987 (N_18987,N_17696,N_17124);
and U18988 (N_18988,N_17816,N_17484);
and U18989 (N_18989,N_16979,N_16485);
and U18990 (N_18990,N_17704,N_17473);
nand U18991 (N_18991,N_16697,N_16567);
nand U18992 (N_18992,N_16078,N_16112);
and U18993 (N_18993,N_16834,N_17073);
or U18994 (N_18994,N_17912,N_17584);
nand U18995 (N_18995,N_16898,N_17864);
xnor U18996 (N_18996,N_16301,N_16342);
nor U18997 (N_18997,N_16513,N_17619);
and U18998 (N_18998,N_16404,N_17805);
or U18999 (N_18999,N_16912,N_16114);
nor U19000 (N_19000,N_17609,N_16981);
xnor U19001 (N_19001,N_17197,N_16992);
or U19002 (N_19002,N_16704,N_17926);
and U19003 (N_19003,N_17269,N_16473);
nand U19004 (N_19004,N_17790,N_16453);
or U19005 (N_19005,N_16406,N_17364);
nand U19006 (N_19006,N_16568,N_17382);
or U19007 (N_19007,N_17436,N_17328);
nand U19008 (N_19008,N_17066,N_16182);
nand U19009 (N_19009,N_17172,N_17018);
and U19010 (N_19010,N_16593,N_17650);
or U19011 (N_19011,N_17896,N_17255);
or U19012 (N_19012,N_17689,N_17405);
nor U19013 (N_19013,N_16365,N_16459);
nor U19014 (N_19014,N_16814,N_17449);
and U19015 (N_19015,N_17892,N_16117);
nand U19016 (N_19016,N_16861,N_17641);
and U19017 (N_19017,N_17717,N_17582);
nand U19018 (N_19018,N_17175,N_17802);
nand U19019 (N_19019,N_17236,N_17377);
nand U19020 (N_19020,N_17595,N_17199);
nand U19021 (N_19021,N_16149,N_16716);
nor U19022 (N_19022,N_16230,N_16788);
and U19023 (N_19023,N_17778,N_16304);
or U19024 (N_19024,N_16502,N_16928);
nand U19025 (N_19025,N_17072,N_17086);
and U19026 (N_19026,N_17554,N_16712);
nor U19027 (N_19027,N_16752,N_17987);
or U19028 (N_19028,N_17835,N_16202);
and U19029 (N_19029,N_17768,N_17278);
xor U19030 (N_19030,N_16125,N_17798);
and U19031 (N_19031,N_16726,N_17417);
or U19032 (N_19032,N_17801,N_16905);
nor U19033 (N_19033,N_16887,N_17344);
and U19034 (N_19034,N_16969,N_17975);
nand U19035 (N_19035,N_16857,N_17337);
nor U19036 (N_19036,N_16025,N_16613);
nor U19037 (N_19037,N_16342,N_17898);
nor U19038 (N_19038,N_16876,N_16885);
nor U19039 (N_19039,N_17329,N_17480);
and U19040 (N_19040,N_17629,N_16729);
nor U19041 (N_19041,N_16763,N_17878);
nand U19042 (N_19042,N_16868,N_17782);
and U19043 (N_19043,N_17306,N_17677);
nand U19044 (N_19044,N_16369,N_17969);
nor U19045 (N_19045,N_17189,N_17463);
and U19046 (N_19046,N_17298,N_17356);
and U19047 (N_19047,N_16303,N_17305);
nand U19048 (N_19048,N_17700,N_17331);
or U19049 (N_19049,N_17205,N_17556);
or U19050 (N_19050,N_16379,N_17046);
nand U19051 (N_19051,N_16458,N_16883);
nor U19052 (N_19052,N_16682,N_16382);
or U19053 (N_19053,N_17273,N_17698);
nand U19054 (N_19054,N_16942,N_17043);
nand U19055 (N_19055,N_16614,N_16923);
or U19056 (N_19056,N_17931,N_16172);
and U19057 (N_19057,N_17033,N_16231);
nand U19058 (N_19058,N_17212,N_17454);
or U19059 (N_19059,N_16875,N_16353);
nor U19060 (N_19060,N_16312,N_17698);
and U19061 (N_19061,N_16717,N_17323);
nor U19062 (N_19062,N_17673,N_17484);
and U19063 (N_19063,N_16166,N_16634);
nand U19064 (N_19064,N_16105,N_16505);
or U19065 (N_19065,N_16002,N_17420);
or U19066 (N_19066,N_16593,N_16711);
and U19067 (N_19067,N_16032,N_16075);
nor U19068 (N_19068,N_17403,N_17469);
and U19069 (N_19069,N_17434,N_16379);
and U19070 (N_19070,N_16491,N_16255);
nand U19071 (N_19071,N_17843,N_16360);
or U19072 (N_19072,N_16124,N_17837);
xnor U19073 (N_19073,N_17833,N_16511);
nand U19074 (N_19074,N_16819,N_16373);
or U19075 (N_19075,N_16799,N_16501);
or U19076 (N_19076,N_17259,N_17412);
or U19077 (N_19077,N_17188,N_16742);
nand U19078 (N_19078,N_16680,N_17810);
xnor U19079 (N_19079,N_17300,N_17937);
and U19080 (N_19080,N_17661,N_17387);
nor U19081 (N_19081,N_16349,N_16584);
nor U19082 (N_19082,N_16860,N_17484);
xor U19083 (N_19083,N_16737,N_17177);
or U19084 (N_19084,N_16286,N_17508);
or U19085 (N_19085,N_17872,N_17935);
and U19086 (N_19086,N_17329,N_16225);
or U19087 (N_19087,N_16412,N_17323);
and U19088 (N_19088,N_16838,N_17172);
nand U19089 (N_19089,N_17618,N_17095);
and U19090 (N_19090,N_17063,N_16610);
and U19091 (N_19091,N_17708,N_16529);
nor U19092 (N_19092,N_16289,N_17072);
and U19093 (N_19093,N_17084,N_16463);
or U19094 (N_19094,N_16862,N_17575);
and U19095 (N_19095,N_17124,N_17755);
nor U19096 (N_19096,N_17725,N_17741);
or U19097 (N_19097,N_17692,N_16647);
and U19098 (N_19098,N_17254,N_17671);
and U19099 (N_19099,N_17240,N_17159);
nand U19100 (N_19100,N_16934,N_16933);
nand U19101 (N_19101,N_17152,N_16945);
and U19102 (N_19102,N_16479,N_16755);
nand U19103 (N_19103,N_17234,N_17137);
nor U19104 (N_19104,N_16193,N_16933);
nand U19105 (N_19105,N_17610,N_16729);
nor U19106 (N_19106,N_17651,N_16013);
nand U19107 (N_19107,N_16509,N_16256);
nor U19108 (N_19108,N_16068,N_17517);
nor U19109 (N_19109,N_17617,N_17487);
xor U19110 (N_19110,N_16319,N_17362);
and U19111 (N_19111,N_17899,N_17869);
nand U19112 (N_19112,N_17122,N_17874);
or U19113 (N_19113,N_17291,N_17886);
nand U19114 (N_19114,N_17845,N_17757);
nor U19115 (N_19115,N_17198,N_16755);
and U19116 (N_19116,N_16978,N_17476);
and U19117 (N_19117,N_17635,N_17157);
xor U19118 (N_19118,N_16216,N_16668);
nor U19119 (N_19119,N_17504,N_17221);
nand U19120 (N_19120,N_16620,N_16361);
xor U19121 (N_19121,N_16584,N_17193);
and U19122 (N_19122,N_16152,N_17683);
and U19123 (N_19123,N_16151,N_17175);
or U19124 (N_19124,N_16889,N_16460);
nor U19125 (N_19125,N_16279,N_16294);
nand U19126 (N_19126,N_17399,N_17138);
and U19127 (N_19127,N_17458,N_16107);
or U19128 (N_19128,N_17327,N_16239);
nor U19129 (N_19129,N_17091,N_17459);
nor U19130 (N_19130,N_16156,N_16828);
nor U19131 (N_19131,N_16492,N_17784);
nor U19132 (N_19132,N_16049,N_17124);
xnor U19133 (N_19133,N_16103,N_16146);
nor U19134 (N_19134,N_16992,N_17801);
nor U19135 (N_19135,N_16363,N_17122);
and U19136 (N_19136,N_16513,N_16732);
and U19137 (N_19137,N_17727,N_17721);
and U19138 (N_19138,N_17715,N_17244);
or U19139 (N_19139,N_17014,N_17587);
xnor U19140 (N_19140,N_17469,N_16019);
and U19141 (N_19141,N_17019,N_16005);
nand U19142 (N_19142,N_16011,N_16973);
nor U19143 (N_19143,N_17986,N_17813);
nor U19144 (N_19144,N_17472,N_16667);
nor U19145 (N_19145,N_17169,N_17274);
or U19146 (N_19146,N_16294,N_16864);
and U19147 (N_19147,N_17609,N_16166);
xnor U19148 (N_19148,N_16149,N_16928);
and U19149 (N_19149,N_17660,N_17375);
nor U19150 (N_19150,N_17533,N_17351);
and U19151 (N_19151,N_17795,N_16980);
or U19152 (N_19152,N_16810,N_17756);
or U19153 (N_19153,N_17725,N_16964);
and U19154 (N_19154,N_17885,N_17438);
nor U19155 (N_19155,N_16839,N_16319);
nand U19156 (N_19156,N_17212,N_16296);
nand U19157 (N_19157,N_16796,N_16733);
nand U19158 (N_19158,N_16228,N_16721);
and U19159 (N_19159,N_16713,N_17101);
and U19160 (N_19160,N_17473,N_16327);
or U19161 (N_19161,N_17845,N_16661);
xor U19162 (N_19162,N_16175,N_17839);
nor U19163 (N_19163,N_17903,N_17185);
or U19164 (N_19164,N_16165,N_17401);
xor U19165 (N_19165,N_16455,N_16058);
nand U19166 (N_19166,N_17593,N_17624);
or U19167 (N_19167,N_17703,N_16438);
nor U19168 (N_19168,N_17712,N_16266);
nor U19169 (N_19169,N_17711,N_17840);
nor U19170 (N_19170,N_17133,N_17216);
nand U19171 (N_19171,N_16947,N_17979);
nand U19172 (N_19172,N_16066,N_17082);
or U19173 (N_19173,N_17697,N_16171);
and U19174 (N_19174,N_16037,N_17924);
and U19175 (N_19175,N_17501,N_16368);
nand U19176 (N_19176,N_17705,N_16145);
xnor U19177 (N_19177,N_16739,N_16417);
nor U19178 (N_19178,N_16431,N_16104);
or U19179 (N_19179,N_17864,N_16859);
nand U19180 (N_19180,N_16018,N_16855);
or U19181 (N_19181,N_16955,N_17952);
and U19182 (N_19182,N_17516,N_16998);
or U19183 (N_19183,N_17782,N_17560);
or U19184 (N_19184,N_17862,N_16547);
nor U19185 (N_19185,N_17482,N_16270);
and U19186 (N_19186,N_16768,N_16732);
nor U19187 (N_19187,N_16753,N_17243);
nor U19188 (N_19188,N_17713,N_16323);
nor U19189 (N_19189,N_17305,N_16606);
and U19190 (N_19190,N_17964,N_17699);
or U19191 (N_19191,N_16816,N_17624);
xnor U19192 (N_19192,N_16272,N_17427);
xnor U19193 (N_19193,N_17542,N_16304);
or U19194 (N_19194,N_17734,N_17908);
or U19195 (N_19195,N_16202,N_17358);
nand U19196 (N_19196,N_17062,N_16604);
and U19197 (N_19197,N_16615,N_17559);
nand U19198 (N_19198,N_16318,N_16522);
or U19199 (N_19199,N_16520,N_16442);
nand U19200 (N_19200,N_17348,N_16248);
nor U19201 (N_19201,N_16484,N_17224);
or U19202 (N_19202,N_16428,N_16508);
nand U19203 (N_19203,N_16434,N_16669);
nand U19204 (N_19204,N_17606,N_16591);
and U19205 (N_19205,N_16378,N_16564);
nor U19206 (N_19206,N_16324,N_16879);
or U19207 (N_19207,N_16787,N_17556);
nor U19208 (N_19208,N_16081,N_16605);
and U19209 (N_19209,N_16266,N_17410);
and U19210 (N_19210,N_16807,N_16658);
or U19211 (N_19211,N_16571,N_16231);
nor U19212 (N_19212,N_16411,N_16618);
xor U19213 (N_19213,N_17816,N_17528);
and U19214 (N_19214,N_17132,N_16443);
nand U19215 (N_19215,N_16523,N_16706);
xor U19216 (N_19216,N_17240,N_17832);
nand U19217 (N_19217,N_17523,N_17450);
xor U19218 (N_19218,N_16870,N_16050);
and U19219 (N_19219,N_17757,N_17056);
or U19220 (N_19220,N_17449,N_17725);
nor U19221 (N_19221,N_16742,N_16381);
nand U19222 (N_19222,N_17269,N_17152);
nor U19223 (N_19223,N_17523,N_17107);
nor U19224 (N_19224,N_17190,N_16468);
and U19225 (N_19225,N_17212,N_17707);
nor U19226 (N_19226,N_16175,N_16396);
xor U19227 (N_19227,N_16344,N_16562);
or U19228 (N_19228,N_16598,N_16384);
nand U19229 (N_19229,N_16819,N_16504);
nor U19230 (N_19230,N_17011,N_17874);
or U19231 (N_19231,N_17915,N_17382);
nand U19232 (N_19232,N_16824,N_16419);
nor U19233 (N_19233,N_16024,N_16882);
xor U19234 (N_19234,N_16366,N_17033);
and U19235 (N_19235,N_17317,N_16474);
nor U19236 (N_19236,N_17606,N_17908);
or U19237 (N_19237,N_16523,N_17474);
nor U19238 (N_19238,N_16685,N_17712);
and U19239 (N_19239,N_16233,N_16522);
or U19240 (N_19240,N_16885,N_17901);
nand U19241 (N_19241,N_17514,N_16502);
nor U19242 (N_19242,N_17348,N_16268);
nor U19243 (N_19243,N_16076,N_17744);
nor U19244 (N_19244,N_16150,N_16182);
nor U19245 (N_19245,N_17888,N_17129);
and U19246 (N_19246,N_16942,N_17659);
nand U19247 (N_19247,N_17332,N_16648);
nand U19248 (N_19248,N_16163,N_16673);
nor U19249 (N_19249,N_17748,N_17918);
and U19250 (N_19250,N_17607,N_16922);
nor U19251 (N_19251,N_16790,N_17593);
or U19252 (N_19252,N_17515,N_17611);
nand U19253 (N_19253,N_16878,N_16954);
nand U19254 (N_19254,N_16383,N_16986);
and U19255 (N_19255,N_16924,N_17871);
and U19256 (N_19256,N_16810,N_17460);
xor U19257 (N_19257,N_17599,N_17195);
nor U19258 (N_19258,N_16804,N_16467);
and U19259 (N_19259,N_16612,N_16973);
nor U19260 (N_19260,N_16984,N_17140);
nand U19261 (N_19261,N_16228,N_17566);
nor U19262 (N_19262,N_17589,N_16915);
xor U19263 (N_19263,N_17946,N_16685);
or U19264 (N_19264,N_16762,N_17874);
and U19265 (N_19265,N_17956,N_16126);
xor U19266 (N_19266,N_17312,N_17549);
nand U19267 (N_19267,N_16333,N_16845);
nand U19268 (N_19268,N_16654,N_17759);
xnor U19269 (N_19269,N_17197,N_17067);
or U19270 (N_19270,N_17537,N_16814);
nor U19271 (N_19271,N_16974,N_16906);
nand U19272 (N_19272,N_16972,N_16279);
or U19273 (N_19273,N_16558,N_16133);
and U19274 (N_19274,N_16128,N_16031);
and U19275 (N_19275,N_17316,N_16069);
or U19276 (N_19276,N_17180,N_16089);
xnor U19277 (N_19277,N_16356,N_16193);
or U19278 (N_19278,N_17608,N_17304);
nor U19279 (N_19279,N_17168,N_16692);
nor U19280 (N_19280,N_16206,N_16761);
and U19281 (N_19281,N_17183,N_17371);
or U19282 (N_19282,N_16802,N_17817);
and U19283 (N_19283,N_16224,N_16871);
and U19284 (N_19284,N_16831,N_16200);
xor U19285 (N_19285,N_16053,N_17043);
or U19286 (N_19286,N_17006,N_16425);
and U19287 (N_19287,N_17504,N_17340);
and U19288 (N_19288,N_17371,N_16891);
xnor U19289 (N_19289,N_16740,N_17951);
and U19290 (N_19290,N_16067,N_17588);
nand U19291 (N_19291,N_16215,N_16424);
and U19292 (N_19292,N_17744,N_17686);
and U19293 (N_19293,N_16780,N_17441);
nor U19294 (N_19294,N_16629,N_16127);
or U19295 (N_19295,N_17137,N_17855);
nor U19296 (N_19296,N_17283,N_17996);
nor U19297 (N_19297,N_17699,N_16045);
nand U19298 (N_19298,N_17685,N_17773);
nor U19299 (N_19299,N_16766,N_16102);
nor U19300 (N_19300,N_16820,N_17858);
xnor U19301 (N_19301,N_17480,N_17351);
xor U19302 (N_19302,N_16718,N_17991);
and U19303 (N_19303,N_17001,N_17173);
nor U19304 (N_19304,N_17310,N_17579);
nand U19305 (N_19305,N_16748,N_16713);
and U19306 (N_19306,N_16578,N_16163);
and U19307 (N_19307,N_16370,N_17513);
nand U19308 (N_19308,N_17082,N_16689);
and U19309 (N_19309,N_17426,N_17145);
and U19310 (N_19310,N_17456,N_17904);
nand U19311 (N_19311,N_16624,N_16069);
or U19312 (N_19312,N_16830,N_17600);
nor U19313 (N_19313,N_16438,N_16561);
nand U19314 (N_19314,N_17239,N_16929);
or U19315 (N_19315,N_17404,N_17291);
or U19316 (N_19316,N_17606,N_17400);
or U19317 (N_19317,N_16857,N_16942);
and U19318 (N_19318,N_17487,N_16943);
or U19319 (N_19319,N_17778,N_17475);
or U19320 (N_19320,N_16778,N_17270);
xnor U19321 (N_19321,N_17435,N_16639);
nor U19322 (N_19322,N_16564,N_16732);
nor U19323 (N_19323,N_17440,N_16709);
nor U19324 (N_19324,N_17747,N_16439);
nand U19325 (N_19325,N_16855,N_17020);
or U19326 (N_19326,N_17610,N_17562);
nand U19327 (N_19327,N_17302,N_17215);
or U19328 (N_19328,N_16922,N_17428);
xnor U19329 (N_19329,N_17363,N_16512);
nand U19330 (N_19330,N_17232,N_16245);
nor U19331 (N_19331,N_16606,N_17754);
or U19332 (N_19332,N_16780,N_17067);
and U19333 (N_19333,N_17936,N_16385);
nor U19334 (N_19334,N_17847,N_17375);
and U19335 (N_19335,N_17004,N_16434);
or U19336 (N_19336,N_17378,N_16523);
or U19337 (N_19337,N_16113,N_16675);
nand U19338 (N_19338,N_17292,N_16099);
nor U19339 (N_19339,N_17529,N_17331);
and U19340 (N_19340,N_16184,N_16949);
or U19341 (N_19341,N_16928,N_17613);
or U19342 (N_19342,N_17360,N_16050);
nand U19343 (N_19343,N_16478,N_17365);
nand U19344 (N_19344,N_17930,N_17710);
or U19345 (N_19345,N_17510,N_17337);
xnor U19346 (N_19346,N_17351,N_17148);
nor U19347 (N_19347,N_17801,N_17321);
or U19348 (N_19348,N_17953,N_16811);
nor U19349 (N_19349,N_17164,N_16667);
nor U19350 (N_19350,N_16681,N_17400);
or U19351 (N_19351,N_16798,N_16983);
and U19352 (N_19352,N_17759,N_17819);
nor U19353 (N_19353,N_17089,N_17581);
or U19354 (N_19354,N_17440,N_17264);
nand U19355 (N_19355,N_17890,N_17612);
and U19356 (N_19356,N_17566,N_16996);
nand U19357 (N_19357,N_17131,N_16131);
and U19358 (N_19358,N_17308,N_16325);
nand U19359 (N_19359,N_17609,N_17848);
and U19360 (N_19360,N_16377,N_16602);
or U19361 (N_19361,N_17397,N_17682);
and U19362 (N_19362,N_16952,N_16144);
and U19363 (N_19363,N_17126,N_16895);
nor U19364 (N_19364,N_17822,N_16851);
nand U19365 (N_19365,N_17280,N_17423);
nand U19366 (N_19366,N_16875,N_17046);
and U19367 (N_19367,N_17540,N_16031);
nand U19368 (N_19368,N_17643,N_17523);
or U19369 (N_19369,N_17637,N_17565);
and U19370 (N_19370,N_16688,N_17980);
nand U19371 (N_19371,N_17913,N_16528);
nor U19372 (N_19372,N_17918,N_17180);
nand U19373 (N_19373,N_17572,N_16096);
nand U19374 (N_19374,N_17362,N_17906);
nor U19375 (N_19375,N_16803,N_17439);
nor U19376 (N_19376,N_17367,N_17581);
and U19377 (N_19377,N_17018,N_17700);
nand U19378 (N_19378,N_16039,N_17614);
nand U19379 (N_19379,N_17973,N_17889);
or U19380 (N_19380,N_17248,N_16591);
nand U19381 (N_19381,N_16433,N_16002);
nor U19382 (N_19382,N_16560,N_17586);
or U19383 (N_19383,N_16013,N_16454);
nor U19384 (N_19384,N_17593,N_16809);
nand U19385 (N_19385,N_16595,N_17435);
nor U19386 (N_19386,N_17523,N_17775);
and U19387 (N_19387,N_17259,N_16240);
or U19388 (N_19388,N_16256,N_17478);
nor U19389 (N_19389,N_16146,N_17299);
xnor U19390 (N_19390,N_17003,N_16780);
nand U19391 (N_19391,N_17431,N_17232);
or U19392 (N_19392,N_17297,N_17687);
nor U19393 (N_19393,N_16376,N_16881);
nand U19394 (N_19394,N_17916,N_17345);
nor U19395 (N_19395,N_17021,N_16030);
nor U19396 (N_19396,N_17331,N_17406);
nor U19397 (N_19397,N_17782,N_16569);
nand U19398 (N_19398,N_16967,N_16627);
nor U19399 (N_19399,N_17490,N_17191);
and U19400 (N_19400,N_16766,N_17051);
xor U19401 (N_19401,N_17906,N_16619);
and U19402 (N_19402,N_17167,N_17577);
or U19403 (N_19403,N_17384,N_17362);
xor U19404 (N_19404,N_17413,N_17494);
and U19405 (N_19405,N_16179,N_17382);
nand U19406 (N_19406,N_17114,N_17017);
and U19407 (N_19407,N_16500,N_16655);
and U19408 (N_19408,N_16905,N_17059);
and U19409 (N_19409,N_17418,N_17081);
nor U19410 (N_19410,N_16845,N_16311);
nand U19411 (N_19411,N_17265,N_17848);
or U19412 (N_19412,N_16683,N_17539);
or U19413 (N_19413,N_17215,N_16798);
nor U19414 (N_19414,N_17995,N_17609);
or U19415 (N_19415,N_17121,N_17520);
or U19416 (N_19416,N_16038,N_17686);
nand U19417 (N_19417,N_17963,N_16495);
xor U19418 (N_19418,N_16078,N_16659);
nand U19419 (N_19419,N_17244,N_17354);
or U19420 (N_19420,N_16366,N_17027);
nand U19421 (N_19421,N_16163,N_17509);
or U19422 (N_19422,N_16806,N_17065);
nor U19423 (N_19423,N_17846,N_16598);
nand U19424 (N_19424,N_16107,N_17482);
xnor U19425 (N_19425,N_16846,N_16863);
or U19426 (N_19426,N_16272,N_17364);
and U19427 (N_19427,N_16611,N_16110);
and U19428 (N_19428,N_16632,N_16450);
xor U19429 (N_19429,N_16423,N_17829);
and U19430 (N_19430,N_16168,N_17248);
or U19431 (N_19431,N_17355,N_16225);
nand U19432 (N_19432,N_16873,N_17742);
nor U19433 (N_19433,N_16065,N_16913);
nand U19434 (N_19434,N_17670,N_16954);
or U19435 (N_19435,N_16250,N_16191);
or U19436 (N_19436,N_16068,N_16439);
nand U19437 (N_19437,N_17239,N_16553);
nor U19438 (N_19438,N_16569,N_16817);
nor U19439 (N_19439,N_17367,N_16786);
nand U19440 (N_19440,N_16451,N_17220);
nor U19441 (N_19441,N_17012,N_16462);
nand U19442 (N_19442,N_16485,N_16539);
or U19443 (N_19443,N_17352,N_16294);
nor U19444 (N_19444,N_16503,N_17143);
nor U19445 (N_19445,N_17854,N_17067);
and U19446 (N_19446,N_17760,N_16457);
nor U19447 (N_19447,N_17050,N_16295);
nor U19448 (N_19448,N_17626,N_16838);
or U19449 (N_19449,N_16333,N_16276);
nor U19450 (N_19450,N_17524,N_17721);
and U19451 (N_19451,N_17507,N_16670);
or U19452 (N_19452,N_17323,N_17390);
or U19453 (N_19453,N_17099,N_16456);
or U19454 (N_19454,N_16450,N_16681);
and U19455 (N_19455,N_16461,N_17158);
nor U19456 (N_19456,N_16028,N_17707);
nand U19457 (N_19457,N_17029,N_17156);
nand U19458 (N_19458,N_17174,N_17036);
or U19459 (N_19459,N_17561,N_16129);
nand U19460 (N_19460,N_17659,N_16335);
or U19461 (N_19461,N_16934,N_17093);
and U19462 (N_19462,N_17571,N_16817);
or U19463 (N_19463,N_16123,N_16013);
nand U19464 (N_19464,N_16474,N_16444);
xor U19465 (N_19465,N_16909,N_17726);
and U19466 (N_19466,N_17312,N_16793);
nor U19467 (N_19467,N_16487,N_16941);
and U19468 (N_19468,N_17008,N_16963);
nand U19469 (N_19469,N_17609,N_16431);
or U19470 (N_19470,N_17679,N_17932);
or U19471 (N_19471,N_17454,N_17028);
and U19472 (N_19472,N_17827,N_17651);
and U19473 (N_19473,N_16410,N_16057);
nor U19474 (N_19474,N_16497,N_16669);
or U19475 (N_19475,N_17051,N_17259);
nand U19476 (N_19476,N_17070,N_16463);
and U19477 (N_19477,N_17985,N_17489);
nand U19478 (N_19478,N_17343,N_17557);
or U19479 (N_19479,N_16707,N_16919);
nand U19480 (N_19480,N_16230,N_17398);
and U19481 (N_19481,N_17308,N_17597);
nand U19482 (N_19482,N_16241,N_17227);
nand U19483 (N_19483,N_17528,N_17922);
nor U19484 (N_19484,N_16588,N_17708);
or U19485 (N_19485,N_16122,N_17681);
nand U19486 (N_19486,N_17980,N_17379);
nand U19487 (N_19487,N_17748,N_16003);
xor U19488 (N_19488,N_17550,N_16909);
or U19489 (N_19489,N_17907,N_17614);
nand U19490 (N_19490,N_16138,N_17151);
and U19491 (N_19491,N_17919,N_17307);
nand U19492 (N_19492,N_17955,N_16998);
or U19493 (N_19493,N_17058,N_16016);
and U19494 (N_19494,N_17766,N_17006);
nor U19495 (N_19495,N_17551,N_17063);
and U19496 (N_19496,N_16419,N_16116);
and U19497 (N_19497,N_17300,N_16413);
nand U19498 (N_19498,N_16370,N_17074);
and U19499 (N_19499,N_17058,N_17376);
nor U19500 (N_19500,N_17905,N_16001);
and U19501 (N_19501,N_17823,N_17573);
or U19502 (N_19502,N_17864,N_17894);
nand U19503 (N_19503,N_16237,N_17914);
and U19504 (N_19504,N_17960,N_17506);
nand U19505 (N_19505,N_17565,N_17139);
nor U19506 (N_19506,N_17182,N_16473);
nor U19507 (N_19507,N_16013,N_16528);
or U19508 (N_19508,N_17244,N_17031);
nand U19509 (N_19509,N_17671,N_17496);
and U19510 (N_19510,N_17011,N_16368);
nor U19511 (N_19511,N_17001,N_16364);
or U19512 (N_19512,N_17592,N_17090);
or U19513 (N_19513,N_17889,N_17108);
xor U19514 (N_19514,N_16669,N_16996);
nand U19515 (N_19515,N_16736,N_16211);
nor U19516 (N_19516,N_17176,N_17655);
nand U19517 (N_19517,N_17318,N_16318);
nand U19518 (N_19518,N_16636,N_17805);
and U19519 (N_19519,N_17362,N_17253);
xnor U19520 (N_19520,N_17399,N_17972);
nor U19521 (N_19521,N_16412,N_17244);
nand U19522 (N_19522,N_17978,N_17504);
nor U19523 (N_19523,N_16740,N_16138);
xnor U19524 (N_19524,N_16442,N_17157);
and U19525 (N_19525,N_17123,N_16779);
and U19526 (N_19526,N_16315,N_17019);
or U19527 (N_19527,N_17992,N_16267);
nor U19528 (N_19528,N_16329,N_16755);
nand U19529 (N_19529,N_16584,N_17877);
nor U19530 (N_19530,N_16236,N_16481);
or U19531 (N_19531,N_17018,N_16854);
nand U19532 (N_19532,N_17445,N_17126);
nor U19533 (N_19533,N_17510,N_16557);
nand U19534 (N_19534,N_17771,N_17626);
xnor U19535 (N_19535,N_16638,N_16357);
and U19536 (N_19536,N_16502,N_16314);
nand U19537 (N_19537,N_16247,N_16565);
nor U19538 (N_19538,N_17527,N_16965);
nand U19539 (N_19539,N_17001,N_17677);
xnor U19540 (N_19540,N_16091,N_16174);
nand U19541 (N_19541,N_16188,N_17160);
nor U19542 (N_19542,N_17178,N_16191);
or U19543 (N_19543,N_16556,N_17319);
nor U19544 (N_19544,N_16464,N_16093);
nor U19545 (N_19545,N_17093,N_17471);
or U19546 (N_19546,N_17731,N_16018);
xor U19547 (N_19547,N_17944,N_16392);
nor U19548 (N_19548,N_17041,N_16109);
nor U19549 (N_19549,N_16762,N_16683);
or U19550 (N_19550,N_16167,N_17660);
or U19551 (N_19551,N_16599,N_16284);
or U19552 (N_19552,N_16027,N_16596);
or U19553 (N_19553,N_17342,N_17124);
or U19554 (N_19554,N_17671,N_16892);
and U19555 (N_19555,N_17774,N_16235);
and U19556 (N_19556,N_16620,N_16768);
or U19557 (N_19557,N_17152,N_16687);
or U19558 (N_19558,N_16114,N_16029);
nor U19559 (N_19559,N_17670,N_16824);
and U19560 (N_19560,N_17728,N_16345);
nand U19561 (N_19561,N_17211,N_17720);
nor U19562 (N_19562,N_17987,N_16800);
xnor U19563 (N_19563,N_16628,N_17674);
or U19564 (N_19564,N_17656,N_16371);
or U19565 (N_19565,N_16474,N_17227);
nand U19566 (N_19566,N_16468,N_17012);
nand U19567 (N_19567,N_17980,N_16642);
xnor U19568 (N_19568,N_17610,N_16368);
or U19569 (N_19569,N_16764,N_16747);
nand U19570 (N_19570,N_16876,N_16129);
nor U19571 (N_19571,N_17081,N_17472);
nand U19572 (N_19572,N_17500,N_17583);
and U19573 (N_19573,N_16494,N_17643);
nor U19574 (N_19574,N_17953,N_17643);
nor U19575 (N_19575,N_17636,N_17328);
and U19576 (N_19576,N_16927,N_16041);
xor U19577 (N_19577,N_17142,N_16192);
nand U19578 (N_19578,N_16090,N_17476);
and U19579 (N_19579,N_17030,N_17092);
nand U19580 (N_19580,N_16677,N_17833);
nand U19581 (N_19581,N_17335,N_17404);
nor U19582 (N_19582,N_17183,N_17093);
nor U19583 (N_19583,N_17528,N_17848);
or U19584 (N_19584,N_16203,N_16487);
nand U19585 (N_19585,N_17790,N_17523);
nor U19586 (N_19586,N_16064,N_17310);
xnor U19587 (N_19587,N_16896,N_17483);
nor U19588 (N_19588,N_17739,N_16158);
or U19589 (N_19589,N_17179,N_17869);
nand U19590 (N_19590,N_17003,N_17052);
nand U19591 (N_19591,N_16087,N_16703);
xnor U19592 (N_19592,N_17878,N_16803);
nand U19593 (N_19593,N_17764,N_16336);
or U19594 (N_19594,N_17657,N_17614);
nor U19595 (N_19595,N_16359,N_17320);
nor U19596 (N_19596,N_16564,N_17754);
nand U19597 (N_19597,N_16914,N_16806);
and U19598 (N_19598,N_17797,N_16293);
and U19599 (N_19599,N_16668,N_17417);
nor U19600 (N_19600,N_16959,N_17603);
xnor U19601 (N_19601,N_17851,N_17986);
nor U19602 (N_19602,N_16390,N_16605);
or U19603 (N_19603,N_16991,N_16462);
and U19604 (N_19604,N_17430,N_17910);
and U19605 (N_19605,N_16304,N_17161);
and U19606 (N_19606,N_17489,N_16920);
nor U19607 (N_19607,N_17035,N_17520);
and U19608 (N_19608,N_16050,N_17642);
nor U19609 (N_19609,N_17317,N_16443);
and U19610 (N_19610,N_17244,N_16154);
and U19611 (N_19611,N_16752,N_17835);
nor U19612 (N_19612,N_17290,N_17214);
and U19613 (N_19613,N_16900,N_17342);
and U19614 (N_19614,N_16346,N_16920);
nor U19615 (N_19615,N_17637,N_16128);
and U19616 (N_19616,N_16132,N_16213);
nand U19617 (N_19617,N_16936,N_17870);
nor U19618 (N_19618,N_16290,N_17868);
nor U19619 (N_19619,N_17428,N_16833);
or U19620 (N_19620,N_17132,N_17349);
nand U19621 (N_19621,N_16086,N_16402);
nand U19622 (N_19622,N_16626,N_16344);
and U19623 (N_19623,N_16094,N_17827);
and U19624 (N_19624,N_17580,N_16324);
or U19625 (N_19625,N_16220,N_17236);
or U19626 (N_19626,N_16170,N_16530);
nor U19627 (N_19627,N_17098,N_17607);
nor U19628 (N_19628,N_17255,N_16614);
and U19629 (N_19629,N_17116,N_16310);
nand U19630 (N_19630,N_17383,N_17230);
nand U19631 (N_19631,N_16972,N_16316);
xnor U19632 (N_19632,N_17246,N_16203);
and U19633 (N_19633,N_16974,N_17443);
nor U19634 (N_19634,N_17540,N_17017);
or U19635 (N_19635,N_17218,N_16768);
or U19636 (N_19636,N_17022,N_16943);
nor U19637 (N_19637,N_17637,N_17201);
or U19638 (N_19638,N_17796,N_16391);
xor U19639 (N_19639,N_16868,N_16622);
nand U19640 (N_19640,N_17623,N_17357);
xnor U19641 (N_19641,N_16881,N_17330);
nand U19642 (N_19642,N_17097,N_16654);
nor U19643 (N_19643,N_17267,N_16915);
or U19644 (N_19644,N_16816,N_16101);
nor U19645 (N_19645,N_16647,N_16902);
nand U19646 (N_19646,N_16459,N_16409);
or U19647 (N_19647,N_16675,N_16693);
and U19648 (N_19648,N_16575,N_17976);
and U19649 (N_19649,N_16290,N_16935);
and U19650 (N_19650,N_17912,N_17531);
nor U19651 (N_19651,N_17816,N_16840);
and U19652 (N_19652,N_16550,N_16659);
nand U19653 (N_19653,N_17877,N_16502);
xor U19654 (N_19654,N_16188,N_16944);
and U19655 (N_19655,N_16680,N_16280);
xor U19656 (N_19656,N_17344,N_17459);
and U19657 (N_19657,N_17605,N_16413);
and U19658 (N_19658,N_16380,N_17593);
and U19659 (N_19659,N_16960,N_16203);
nor U19660 (N_19660,N_17200,N_17158);
and U19661 (N_19661,N_16749,N_17589);
nor U19662 (N_19662,N_16210,N_16194);
or U19663 (N_19663,N_16790,N_17114);
nor U19664 (N_19664,N_16616,N_16790);
and U19665 (N_19665,N_16647,N_16932);
and U19666 (N_19666,N_17316,N_17212);
or U19667 (N_19667,N_16552,N_17549);
and U19668 (N_19668,N_17767,N_16053);
xnor U19669 (N_19669,N_17708,N_17587);
nor U19670 (N_19670,N_17999,N_17605);
and U19671 (N_19671,N_17436,N_17759);
nand U19672 (N_19672,N_17927,N_17992);
xor U19673 (N_19673,N_16154,N_16582);
or U19674 (N_19674,N_17693,N_16791);
nor U19675 (N_19675,N_16177,N_16342);
nor U19676 (N_19676,N_17339,N_17138);
xor U19677 (N_19677,N_17359,N_16444);
nand U19678 (N_19678,N_16911,N_16946);
and U19679 (N_19679,N_16673,N_16933);
or U19680 (N_19680,N_16347,N_17411);
nand U19681 (N_19681,N_17910,N_16714);
nand U19682 (N_19682,N_17083,N_17004);
or U19683 (N_19683,N_17017,N_16443);
nand U19684 (N_19684,N_17234,N_16788);
xnor U19685 (N_19685,N_16315,N_17356);
and U19686 (N_19686,N_16600,N_16678);
and U19687 (N_19687,N_17386,N_16674);
nand U19688 (N_19688,N_16001,N_16581);
nor U19689 (N_19689,N_16189,N_17357);
and U19690 (N_19690,N_16801,N_16720);
nand U19691 (N_19691,N_16119,N_17094);
xor U19692 (N_19692,N_17890,N_16154);
nand U19693 (N_19693,N_16733,N_17117);
and U19694 (N_19694,N_16543,N_16372);
nand U19695 (N_19695,N_17023,N_16154);
nand U19696 (N_19696,N_17139,N_17552);
nand U19697 (N_19697,N_17348,N_17545);
nor U19698 (N_19698,N_17918,N_16120);
nor U19699 (N_19699,N_17429,N_17092);
and U19700 (N_19700,N_17977,N_16023);
xor U19701 (N_19701,N_17097,N_16077);
nand U19702 (N_19702,N_17608,N_16232);
nand U19703 (N_19703,N_17849,N_16909);
nor U19704 (N_19704,N_17069,N_16652);
and U19705 (N_19705,N_17824,N_16115);
xnor U19706 (N_19706,N_16603,N_17061);
or U19707 (N_19707,N_17621,N_16747);
and U19708 (N_19708,N_16425,N_16743);
nand U19709 (N_19709,N_16402,N_17107);
and U19710 (N_19710,N_16212,N_16512);
or U19711 (N_19711,N_16424,N_16555);
xnor U19712 (N_19712,N_16845,N_16332);
and U19713 (N_19713,N_16038,N_16242);
nand U19714 (N_19714,N_16511,N_16170);
or U19715 (N_19715,N_16729,N_17111);
nor U19716 (N_19716,N_16486,N_17994);
or U19717 (N_19717,N_17998,N_16480);
nand U19718 (N_19718,N_17985,N_17866);
or U19719 (N_19719,N_17544,N_17542);
and U19720 (N_19720,N_16135,N_17555);
nand U19721 (N_19721,N_16733,N_17917);
nand U19722 (N_19722,N_16458,N_16242);
nand U19723 (N_19723,N_16738,N_17790);
nor U19724 (N_19724,N_17852,N_17941);
and U19725 (N_19725,N_17886,N_17326);
nor U19726 (N_19726,N_16601,N_17277);
nor U19727 (N_19727,N_16669,N_17003);
nand U19728 (N_19728,N_16716,N_17255);
xnor U19729 (N_19729,N_16727,N_16756);
or U19730 (N_19730,N_16889,N_17495);
or U19731 (N_19731,N_17441,N_17589);
xor U19732 (N_19732,N_17114,N_16887);
nand U19733 (N_19733,N_16561,N_17555);
and U19734 (N_19734,N_17611,N_17280);
nand U19735 (N_19735,N_16779,N_16003);
and U19736 (N_19736,N_16921,N_16139);
xor U19737 (N_19737,N_17572,N_16068);
nand U19738 (N_19738,N_16577,N_16083);
and U19739 (N_19739,N_17269,N_16367);
and U19740 (N_19740,N_17810,N_16242);
xor U19741 (N_19741,N_16960,N_17489);
nor U19742 (N_19742,N_16726,N_16888);
or U19743 (N_19743,N_16604,N_17408);
nand U19744 (N_19744,N_17293,N_16615);
nand U19745 (N_19745,N_17149,N_16618);
and U19746 (N_19746,N_16293,N_16279);
nor U19747 (N_19747,N_16767,N_16705);
xnor U19748 (N_19748,N_17496,N_17588);
and U19749 (N_19749,N_16302,N_17171);
and U19750 (N_19750,N_17291,N_17168);
or U19751 (N_19751,N_16020,N_16164);
and U19752 (N_19752,N_16730,N_17871);
xor U19753 (N_19753,N_16168,N_17575);
nor U19754 (N_19754,N_17875,N_17295);
or U19755 (N_19755,N_16813,N_17789);
nand U19756 (N_19756,N_16629,N_16647);
nor U19757 (N_19757,N_17581,N_17635);
xnor U19758 (N_19758,N_17811,N_16558);
nand U19759 (N_19759,N_16137,N_16481);
and U19760 (N_19760,N_16739,N_17891);
or U19761 (N_19761,N_17961,N_17492);
xnor U19762 (N_19762,N_17248,N_16154);
and U19763 (N_19763,N_16021,N_16356);
and U19764 (N_19764,N_17132,N_16012);
and U19765 (N_19765,N_16451,N_16595);
nor U19766 (N_19766,N_17170,N_16226);
xor U19767 (N_19767,N_17488,N_16629);
nor U19768 (N_19768,N_17700,N_16963);
and U19769 (N_19769,N_16219,N_16063);
nor U19770 (N_19770,N_17896,N_16717);
nand U19771 (N_19771,N_16283,N_17847);
or U19772 (N_19772,N_17538,N_16371);
and U19773 (N_19773,N_17377,N_17431);
nand U19774 (N_19774,N_16505,N_17629);
and U19775 (N_19775,N_17631,N_17698);
or U19776 (N_19776,N_16241,N_16319);
or U19777 (N_19777,N_17099,N_16615);
and U19778 (N_19778,N_17894,N_17396);
nand U19779 (N_19779,N_16632,N_16883);
xnor U19780 (N_19780,N_17106,N_16652);
nand U19781 (N_19781,N_17908,N_16934);
xor U19782 (N_19782,N_16179,N_17182);
nor U19783 (N_19783,N_16276,N_16659);
nor U19784 (N_19784,N_17988,N_17315);
xor U19785 (N_19785,N_16080,N_16923);
nand U19786 (N_19786,N_16162,N_17254);
nor U19787 (N_19787,N_16780,N_16589);
nand U19788 (N_19788,N_16527,N_17143);
nand U19789 (N_19789,N_16394,N_16453);
nor U19790 (N_19790,N_16985,N_16572);
and U19791 (N_19791,N_16527,N_16944);
or U19792 (N_19792,N_16978,N_16629);
or U19793 (N_19793,N_17237,N_17653);
nor U19794 (N_19794,N_16276,N_16772);
or U19795 (N_19795,N_16173,N_17027);
xor U19796 (N_19796,N_16979,N_17086);
xor U19797 (N_19797,N_17560,N_17931);
or U19798 (N_19798,N_17178,N_16302);
nand U19799 (N_19799,N_16037,N_17637);
nor U19800 (N_19800,N_17000,N_16921);
nand U19801 (N_19801,N_17444,N_16617);
or U19802 (N_19802,N_16428,N_16317);
or U19803 (N_19803,N_17298,N_17992);
nand U19804 (N_19804,N_17825,N_17520);
nor U19805 (N_19805,N_16009,N_16135);
or U19806 (N_19806,N_16285,N_17987);
nand U19807 (N_19807,N_16133,N_16755);
xor U19808 (N_19808,N_16897,N_17868);
or U19809 (N_19809,N_16368,N_17590);
nor U19810 (N_19810,N_16994,N_17434);
or U19811 (N_19811,N_16402,N_17486);
or U19812 (N_19812,N_16956,N_16975);
nor U19813 (N_19813,N_17413,N_16897);
and U19814 (N_19814,N_16499,N_16648);
or U19815 (N_19815,N_16364,N_17840);
nand U19816 (N_19816,N_16486,N_16992);
nor U19817 (N_19817,N_16096,N_16904);
nand U19818 (N_19818,N_17087,N_17152);
nor U19819 (N_19819,N_16328,N_16264);
or U19820 (N_19820,N_16445,N_17207);
and U19821 (N_19821,N_17179,N_17420);
nand U19822 (N_19822,N_17067,N_17530);
and U19823 (N_19823,N_16052,N_17416);
nor U19824 (N_19824,N_16474,N_17695);
nor U19825 (N_19825,N_17894,N_16748);
nand U19826 (N_19826,N_17796,N_17690);
or U19827 (N_19827,N_17600,N_17477);
or U19828 (N_19828,N_17436,N_17497);
or U19829 (N_19829,N_16441,N_16950);
nand U19830 (N_19830,N_16112,N_16114);
and U19831 (N_19831,N_16249,N_16055);
nand U19832 (N_19832,N_17902,N_17855);
nor U19833 (N_19833,N_16145,N_16130);
nor U19834 (N_19834,N_16910,N_17938);
nand U19835 (N_19835,N_16796,N_17748);
and U19836 (N_19836,N_17079,N_17070);
or U19837 (N_19837,N_17890,N_17026);
or U19838 (N_19838,N_17661,N_16767);
or U19839 (N_19839,N_17788,N_16693);
or U19840 (N_19840,N_16080,N_16576);
and U19841 (N_19841,N_17880,N_17716);
or U19842 (N_19842,N_16971,N_17579);
nand U19843 (N_19843,N_17502,N_16389);
nand U19844 (N_19844,N_17225,N_17465);
or U19845 (N_19845,N_16419,N_17962);
nor U19846 (N_19846,N_17417,N_17905);
and U19847 (N_19847,N_16316,N_16641);
or U19848 (N_19848,N_17461,N_17030);
xnor U19849 (N_19849,N_16753,N_17255);
nor U19850 (N_19850,N_17483,N_17652);
and U19851 (N_19851,N_17426,N_16981);
nand U19852 (N_19852,N_16547,N_16315);
nor U19853 (N_19853,N_16258,N_17545);
nand U19854 (N_19854,N_16547,N_16787);
nand U19855 (N_19855,N_16417,N_17420);
and U19856 (N_19856,N_17419,N_16186);
or U19857 (N_19857,N_17442,N_17710);
and U19858 (N_19858,N_17985,N_16663);
nor U19859 (N_19859,N_16582,N_16142);
and U19860 (N_19860,N_16572,N_17567);
nand U19861 (N_19861,N_16109,N_17163);
nor U19862 (N_19862,N_16339,N_16388);
nand U19863 (N_19863,N_17686,N_16066);
or U19864 (N_19864,N_17900,N_17747);
xnor U19865 (N_19865,N_17628,N_17858);
and U19866 (N_19866,N_16854,N_17235);
and U19867 (N_19867,N_17404,N_16703);
xor U19868 (N_19868,N_16871,N_17967);
xnor U19869 (N_19869,N_17083,N_17375);
or U19870 (N_19870,N_16155,N_17782);
or U19871 (N_19871,N_17011,N_16661);
nand U19872 (N_19872,N_16420,N_16113);
nor U19873 (N_19873,N_17749,N_17592);
or U19874 (N_19874,N_17023,N_17422);
or U19875 (N_19875,N_17420,N_16137);
nand U19876 (N_19876,N_17047,N_16518);
nand U19877 (N_19877,N_16735,N_16793);
nand U19878 (N_19878,N_17144,N_16995);
or U19879 (N_19879,N_16491,N_17965);
nor U19880 (N_19880,N_17927,N_17721);
or U19881 (N_19881,N_17467,N_17190);
nand U19882 (N_19882,N_16842,N_16061);
or U19883 (N_19883,N_17535,N_16536);
nor U19884 (N_19884,N_17125,N_17879);
nand U19885 (N_19885,N_17218,N_16944);
nor U19886 (N_19886,N_16167,N_16156);
nand U19887 (N_19887,N_17524,N_16359);
and U19888 (N_19888,N_16731,N_16294);
and U19889 (N_19889,N_17708,N_16246);
and U19890 (N_19890,N_17800,N_17301);
and U19891 (N_19891,N_16386,N_17155);
and U19892 (N_19892,N_16541,N_17381);
xnor U19893 (N_19893,N_16916,N_17641);
or U19894 (N_19894,N_17664,N_16640);
xor U19895 (N_19895,N_16223,N_16078);
nor U19896 (N_19896,N_16177,N_16653);
or U19897 (N_19897,N_16728,N_16782);
or U19898 (N_19898,N_16554,N_17378);
nor U19899 (N_19899,N_16607,N_16127);
or U19900 (N_19900,N_16056,N_17857);
or U19901 (N_19901,N_16407,N_17490);
or U19902 (N_19902,N_16446,N_16058);
xnor U19903 (N_19903,N_16551,N_16987);
or U19904 (N_19904,N_17934,N_17980);
nand U19905 (N_19905,N_17251,N_16384);
nor U19906 (N_19906,N_16549,N_17429);
or U19907 (N_19907,N_17681,N_17634);
xnor U19908 (N_19908,N_17238,N_16778);
and U19909 (N_19909,N_16984,N_16065);
nand U19910 (N_19910,N_17583,N_17765);
xor U19911 (N_19911,N_16348,N_16583);
nand U19912 (N_19912,N_17076,N_16546);
or U19913 (N_19913,N_17895,N_17522);
nand U19914 (N_19914,N_17017,N_17482);
nor U19915 (N_19915,N_17461,N_16788);
nand U19916 (N_19916,N_17847,N_17251);
and U19917 (N_19917,N_17737,N_16086);
and U19918 (N_19918,N_17071,N_17076);
or U19919 (N_19919,N_16336,N_16471);
nor U19920 (N_19920,N_17417,N_16599);
and U19921 (N_19921,N_16508,N_17479);
nand U19922 (N_19922,N_17534,N_17112);
nand U19923 (N_19923,N_16062,N_16521);
nor U19924 (N_19924,N_17883,N_17804);
nor U19925 (N_19925,N_17662,N_17208);
or U19926 (N_19926,N_17895,N_16931);
nand U19927 (N_19927,N_16958,N_16309);
nor U19928 (N_19928,N_16942,N_16284);
nor U19929 (N_19929,N_17450,N_16093);
and U19930 (N_19930,N_16340,N_16084);
nand U19931 (N_19931,N_16231,N_16698);
nand U19932 (N_19932,N_16825,N_17747);
nor U19933 (N_19933,N_17801,N_16460);
nand U19934 (N_19934,N_16742,N_16879);
nor U19935 (N_19935,N_17556,N_16624);
and U19936 (N_19936,N_17053,N_16405);
or U19937 (N_19937,N_16539,N_17167);
and U19938 (N_19938,N_16875,N_17326);
or U19939 (N_19939,N_17287,N_16779);
or U19940 (N_19940,N_17231,N_16523);
nor U19941 (N_19941,N_16059,N_17913);
and U19942 (N_19942,N_16571,N_17344);
or U19943 (N_19943,N_16113,N_16623);
nand U19944 (N_19944,N_16641,N_17740);
nor U19945 (N_19945,N_16682,N_17582);
nor U19946 (N_19946,N_17827,N_16560);
nor U19947 (N_19947,N_16023,N_16056);
nor U19948 (N_19948,N_17209,N_16522);
xor U19949 (N_19949,N_16967,N_17142);
and U19950 (N_19950,N_17253,N_16027);
or U19951 (N_19951,N_17102,N_17493);
nand U19952 (N_19952,N_17465,N_17704);
or U19953 (N_19953,N_16827,N_17454);
and U19954 (N_19954,N_16513,N_16687);
nor U19955 (N_19955,N_17508,N_16054);
or U19956 (N_19956,N_17799,N_17356);
and U19957 (N_19957,N_17865,N_17338);
or U19958 (N_19958,N_16953,N_17483);
nand U19959 (N_19959,N_17245,N_17101);
nor U19960 (N_19960,N_16759,N_17752);
xor U19961 (N_19961,N_17828,N_17808);
or U19962 (N_19962,N_17761,N_16624);
xnor U19963 (N_19963,N_17741,N_17019);
nand U19964 (N_19964,N_16792,N_17592);
xor U19965 (N_19965,N_17883,N_17662);
nand U19966 (N_19966,N_17726,N_17061);
and U19967 (N_19967,N_17604,N_17140);
nand U19968 (N_19968,N_16773,N_17269);
nand U19969 (N_19969,N_16748,N_16610);
and U19970 (N_19970,N_16596,N_17240);
and U19971 (N_19971,N_17522,N_16796);
nor U19972 (N_19972,N_17291,N_17267);
and U19973 (N_19973,N_17402,N_17239);
or U19974 (N_19974,N_17982,N_16838);
nand U19975 (N_19975,N_17531,N_16768);
and U19976 (N_19976,N_17919,N_17961);
and U19977 (N_19977,N_17500,N_17297);
or U19978 (N_19978,N_17881,N_17541);
nor U19979 (N_19979,N_17274,N_16049);
and U19980 (N_19980,N_16606,N_17833);
and U19981 (N_19981,N_17690,N_16895);
nor U19982 (N_19982,N_17830,N_16448);
or U19983 (N_19983,N_17575,N_17819);
nand U19984 (N_19984,N_17209,N_17097);
nor U19985 (N_19985,N_16883,N_16405);
and U19986 (N_19986,N_16980,N_16251);
or U19987 (N_19987,N_17772,N_16138);
nor U19988 (N_19988,N_16875,N_17636);
nor U19989 (N_19989,N_17991,N_16369);
xor U19990 (N_19990,N_17197,N_17380);
nor U19991 (N_19991,N_17085,N_16362);
xnor U19992 (N_19992,N_16241,N_16921);
or U19993 (N_19993,N_16067,N_17860);
nor U19994 (N_19994,N_16133,N_16018);
nand U19995 (N_19995,N_17577,N_17955);
nor U19996 (N_19996,N_16513,N_17494);
and U19997 (N_19997,N_17032,N_17645);
or U19998 (N_19998,N_17693,N_17985);
nand U19999 (N_19999,N_17296,N_17018);
xnor UO_0 (O_0,N_19319,N_18117);
and UO_1 (O_1,N_18885,N_18796);
nand UO_2 (O_2,N_19916,N_18116);
or UO_3 (O_3,N_19668,N_19753);
nand UO_4 (O_4,N_18903,N_18257);
nand UO_5 (O_5,N_18002,N_18670);
nor UO_6 (O_6,N_18775,N_19694);
nor UO_7 (O_7,N_18914,N_19229);
nand UO_8 (O_8,N_18440,N_19301);
nand UO_9 (O_9,N_18530,N_19348);
or UO_10 (O_10,N_19852,N_18853);
nor UO_11 (O_11,N_18490,N_18522);
nor UO_12 (O_12,N_19208,N_19130);
nand UO_13 (O_13,N_18733,N_18863);
or UO_14 (O_14,N_18755,N_18327);
and UO_15 (O_15,N_18409,N_19782);
xor UO_16 (O_16,N_18916,N_19031);
and UO_17 (O_17,N_19575,N_19046);
xor UO_18 (O_18,N_18266,N_18553);
xnor UO_19 (O_19,N_19108,N_19883);
nor UO_20 (O_20,N_18587,N_19003);
xor UO_21 (O_21,N_18435,N_18314);
nor UO_22 (O_22,N_19468,N_18546);
and UO_23 (O_23,N_18279,N_18776);
and UO_24 (O_24,N_18230,N_19273);
nor UO_25 (O_25,N_18021,N_19553);
or UO_26 (O_26,N_19503,N_18904);
and UO_27 (O_27,N_19186,N_18337);
nor UO_28 (O_28,N_18235,N_19905);
and UO_29 (O_29,N_18066,N_19739);
and UO_30 (O_30,N_18586,N_19100);
and UO_31 (O_31,N_18098,N_19906);
nor UO_32 (O_32,N_19631,N_19177);
nand UO_33 (O_33,N_18559,N_19429);
xnor UO_34 (O_34,N_19321,N_19630);
nand UO_35 (O_35,N_19640,N_18386);
xnor UO_36 (O_36,N_19029,N_18069);
nor UO_37 (O_37,N_19927,N_18592);
nand UO_38 (O_38,N_19941,N_19014);
or UO_39 (O_39,N_18186,N_19078);
and UO_40 (O_40,N_19970,N_19152);
or UO_41 (O_41,N_19664,N_18560);
nor UO_42 (O_42,N_18537,N_18525);
nand UO_43 (O_43,N_19472,N_19781);
or UO_44 (O_44,N_18182,N_19483);
or UO_45 (O_45,N_19510,N_19785);
nand UO_46 (O_46,N_19792,N_18390);
nor UO_47 (O_47,N_19121,N_19371);
nor UO_48 (O_48,N_18748,N_19691);
and UO_49 (O_49,N_19324,N_18698);
nand UO_50 (O_50,N_19975,N_19891);
and UO_51 (O_51,N_19262,N_19098);
or UO_52 (O_52,N_19387,N_19166);
nor UO_53 (O_53,N_19446,N_19258);
or UO_54 (O_54,N_19300,N_19990);
or UO_55 (O_55,N_19012,N_18271);
nand UO_56 (O_56,N_19635,N_18138);
nor UO_57 (O_57,N_19135,N_18785);
nor UO_58 (O_58,N_19118,N_18237);
nor UO_59 (O_59,N_19577,N_19068);
nand UO_60 (O_60,N_19735,N_18411);
or UO_61 (O_61,N_19616,N_19952);
or UO_62 (O_62,N_18822,N_19185);
and UO_63 (O_63,N_18662,N_18212);
xor UO_64 (O_64,N_18823,N_19707);
or UO_65 (O_65,N_18373,N_19953);
nor UO_66 (O_66,N_18782,N_19778);
nor UO_67 (O_67,N_19661,N_18623);
or UO_68 (O_68,N_19062,N_19642);
or UO_69 (O_69,N_18418,N_18712);
nand UO_70 (O_70,N_18991,N_18943);
nand UO_71 (O_71,N_18244,N_19058);
and UO_72 (O_72,N_18556,N_19085);
or UO_73 (O_73,N_18091,N_19613);
nand UO_74 (O_74,N_18618,N_19687);
xnor UO_75 (O_75,N_19174,N_18264);
and UO_76 (O_76,N_18947,N_19009);
and UO_77 (O_77,N_19458,N_19230);
or UO_78 (O_78,N_18949,N_19362);
xnor UO_79 (O_79,N_19801,N_19469);
xor UO_80 (O_80,N_19690,N_18577);
nor UO_81 (O_81,N_19679,N_18446);
nor UO_82 (O_82,N_19155,N_18584);
nand UO_83 (O_83,N_18864,N_18371);
and UO_84 (O_84,N_19128,N_18836);
nand UO_85 (O_85,N_18974,N_18602);
nor UO_86 (O_86,N_18136,N_19089);
and UO_87 (O_87,N_18201,N_18896);
or UO_88 (O_88,N_19788,N_19482);
and UO_89 (O_89,N_18064,N_18330);
nor UO_90 (O_90,N_19861,N_19084);
nor UO_91 (O_91,N_19154,N_19655);
nor UO_92 (O_92,N_18451,N_18114);
nor UO_93 (O_93,N_18920,N_18517);
nand UO_94 (O_94,N_19450,N_18861);
and UO_95 (O_95,N_18438,N_19996);
nand UO_96 (O_96,N_18535,N_19625);
and UO_97 (O_97,N_19988,N_19485);
and UO_98 (O_98,N_18869,N_18489);
nand UO_99 (O_99,N_18077,N_19382);
nor UO_100 (O_100,N_18470,N_18402);
nor UO_101 (O_101,N_19545,N_19709);
nor UO_102 (O_102,N_19867,N_19604);
xnor UO_103 (O_103,N_19914,N_18888);
nor UO_104 (O_104,N_18448,N_18539);
xnor UO_105 (O_105,N_18263,N_19373);
nor UO_106 (O_106,N_19111,N_18326);
nand UO_107 (O_107,N_18385,N_18282);
nand UO_108 (O_108,N_18648,N_19183);
nand UO_109 (O_109,N_19091,N_19999);
and UO_110 (O_110,N_19017,N_19415);
nor UO_111 (O_111,N_19143,N_18840);
and UO_112 (O_112,N_18778,N_18014);
nor UO_113 (O_113,N_19726,N_18379);
and UO_114 (O_114,N_18959,N_18100);
nor UO_115 (O_115,N_19278,N_18696);
xnor UO_116 (O_116,N_18972,N_18941);
nor UO_117 (O_117,N_18955,N_18012);
nand UO_118 (O_118,N_18514,N_19515);
nor UO_119 (O_119,N_19368,N_18845);
and UO_120 (O_120,N_19203,N_19930);
nor UO_121 (O_121,N_19167,N_19488);
nor UO_122 (O_122,N_19981,N_19391);
and UO_123 (O_123,N_18984,N_19473);
and UO_124 (O_124,N_18819,N_18210);
or UO_125 (O_125,N_18688,N_18042);
nor UO_126 (O_126,N_18258,N_18180);
nand UO_127 (O_127,N_18987,N_19598);
and UO_128 (O_128,N_18601,N_18807);
nand UO_129 (O_129,N_18509,N_18950);
or UO_130 (O_130,N_18147,N_19414);
and UO_131 (O_131,N_18693,N_19431);
nor UO_132 (O_132,N_19833,N_18044);
xor UO_133 (O_133,N_19310,N_18394);
and UO_134 (O_134,N_18301,N_18893);
and UO_135 (O_135,N_19037,N_18028);
xor UO_136 (O_136,N_19856,N_18208);
nor UO_137 (O_137,N_19741,N_19148);
and UO_138 (O_138,N_18083,N_19184);
or UO_139 (O_139,N_18849,N_18550);
nor UO_140 (O_140,N_18225,N_19559);
nor UO_141 (O_141,N_19532,N_18746);
xnor UO_142 (O_142,N_19026,N_18249);
or UO_143 (O_143,N_19369,N_19637);
nand UO_144 (O_144,N_19725,N_18891);
or UO_145 (O_145,N_18882,N_18923);
and UO_146 (O_146,N_19866,N_18469);
and UO_147 (O_147,N_19857,N_18043);
nor UO_148 (O_148,N_19949,N_19983);
nand UO_149 (O_149,N_18039,N_19101);
or UO_150 (O_150,N_18628,N_18273);
xor UO_151 (O_151,N_19090,N_19438);
and UO_152 (O_152,N_19768,N_18484);
nor UO_153 (O_153,N_19823,N_19669);
nand UO_154 (O_154,N_18752,N_18790);
nor UO_155 (O_155,N_18013,N_19169);
or UO_156 (O_156,N_19571,N_18188);
nand UO_157 (O_157,N_19809,N_19752);
or UO_158 (O_158,N_19484,N_18195);
xnor UO_159 (O_159,N_19671,N_18582);
nand UO_160 (O_160,N_18784,N_19918);
nand UO_161 (O_161,N_18524,N_19103);
and UO_162 (O_162,N_19623,N_18604);
and UO_163 (O_163,N_19486,N_19408);
and UO_164 (O_164,N_18770,N_18267);
xnor UO_165 (O_165,N_19743,N_18431);
and UO_166 (O_166,N_19274,N_18133);
nand UO_167 (O_167,N_19194,N_19561);
nand UO_168 (O_168,N_18004,N_19531);
nand UO_169 (O_169,N_18977,N_18088);
nor UO_170 (O_170,N_18757,N_18474);
nor UO_171 (O_171,N_18497,N_19039);
or UO_172 (O_172,N_19182,N_19517);
and UO_173 (O_173,N_19674,N_19693);
and UO_174 (O_174,N_19110,N_18352);
nor UO_175 (O_175,N_19720,N_18001);
or UO_176 (O_176,N_18358,N_19870);
and UO_177 (O_177,N_19609,N_18595);
nor UO_178 (O_178,N_19920,N_19924);
xor UO_179 (O_179,N_18183,N_19765);
and UO_180 (O_180,N_19292,N_18299);
xor UO_181 (O_181,N_19803,N_18175);
nand UO_182 (O_182,N_19233,N_18363);
nand UO_183 (O_183,N_18190,N_19066);
nand UO_184 (O_184,N_18262,N_19897);
nand UO_185 (O_185,N_18009,N_18740);
nor UO_186 (O_186,N_19077,N_18336);
or UO_187 (O_187,N_18049,N_19819);
xor UO_188 (O_188,N_19134,N_19926);
nor UO_189 (O_189,N_19383,N_18905);
nand UO_190 (O_190,N_18983,N_18221);
nand UO_191 (O_191,N_18948,N_18487);
and UO_192 (O_192,N_18513,N_18214);
nand UO_193 (O_193,N_19297,N_18008);
nor UO_194 (O_194,N_19452,N_19699);
nor UO_195 (O_195,N_19296,N_19116);
or UO_196 (O_196,N_18339,N_18593);
nand UO_197 (O_197,N_18838,N_18375);
or UO_198 (O_198,N_18804,N_19762);
nor UO_199 (O_199,N_19276,N_19977);
nand UO_200 (O_200,N_19277,N_19599);
or UO_201 (O_201,N_18806,N_19393);
and UO_202 (O_202,N_18242,N_19961);
nor UO_203 (O_203,N_19147,N_18452);
nand UO_204 (O_204,N_18318,N_19242);
xnor UO_205 (O_205,N_19401,N_18547);
nor UO_206 (O_206,N_18278,N_19427);
or UO_207 (O_207,N_18010,N_18641);
nand UO_208 (O_208,N_19955,N_19298);
or UO_209 (O_209,N_19360,N_19123);
and UO_210 (O_210,N_18055,N_18792);
nor UO_211 (O_211,N_18859,N_18449);
nor UO_212 (O_212,N_19732,N_19567);
or UO_213 (O_213,N_18416,N_18382);
nor UO_214 (O_214,N_19505,N_18189);
or UO_215 (O_215,N_18018,N_19650);
or UO_216 (O_216,N_19295,N_19347);
or UO_217 (O_217,N_18889,N_18989);
and UO_218 (O_218,N_19757,N_19172);
and UO_219 (O_219,N_19322,N_18198);
or UO_220 (O_220,N_19264,N_19652);
nand UO_221 (O_221,N_19774,N_18000);
and UO_222 (O_222,N_18715,N_18518);
xor UO_223 (O_223,N_19855,N_19044);
nor UO_224 (O_224,N_19994,N_18809);
and UO_225 (O_225,N_19754,N_18872);
nand UO_226 (O_226,N_18625,N_19476);
and UO_227 (O_227,N_18824,N_19524);
nand UO_228 (O_228,N_18685,N_19727);
nor UO_229 (O_229,N_19877,N_18516);
nand UO_230 (O_230,N_19795,N_19159);
and UO_231 (O_231,N_18492,N_19263);
or UO_232 (O_232,N_19187,N_19818);
nand UO_233 (O_233,N_19922,N_19943);
or UO_234 (O_234,N_18082,N_19170);
xor UO_235 (O_235,N_19936,N_19326);
nand UO_236 (O_236,N_18324,N_19954);
and UO_237 (O_237,N_18728,N_18291);
or UO_238 (O_238,N_19290,N_19518);
nand UO_239 (O_239,N_19069,N_18458);
nand UO_240 (O_240,N_19848,N_19072);
or UO_241 (O_241,N_18193,N_18684);
nor UO_242 (O_242,N_18050,N_18222);
nand UO_243 (O_243,N_19279,N_19222);
or UO_244 (O_244,N_18570,N_19216);
nand UO_245 (O_245,N_19814,N_18393);
or UO_246 (O_246,N_19911,N_19423);
nor UO_247 (O_247,N_19660,N_19887);
and UO_248 (O_248,N_18202,N_19467);
nor UO_249 (O_249,N_18245,N_19269);
nor UO_250 (O_250,N_18205,N_18852);
and UO_251 (O_251,N_18969,N_19437);
xnor UO_252 (O_252,N_19933,N_19333);
or UO_253 (O_253,N_19620,N_18184);
or UO_254 (O_254,N_18629,N_18229);
or UO_255 (O_255,N_19320,N_19639);
or UO_256 (O_256,N_18437,N_19344);
nor UO_257 (O_257,N_18563,N_19378);
or UO_258 (O_258,N_18313,N_18781);
nor UO_259 (O_259,N_18213,N_18408);
nor UO_260 (O_260,N_19235,N_18999);
nor UO_261 (O_261,N_19251,N_19931);
nor UO_262 (O_262,N_18661,N_19453);
nor UO_263 (O_263,N_18747,N_18059);
and UO_264 (O_264,N_19982,N_19576);
nand UO_265 (O_265,N_19232,N_19049);
and UO_266 (O_266,N_19385,N_18471);
and UO_267 (O_267,N_19428,N_19838);
nor UO_268 (O_268,N_18831,N_19939);
nor UO_269 (O_269,N_19767,N_19481);
nor UO_270 (O_270,N_18721,N_18632);
nor UO_271 (O_271,N_19672,N_18159);
or UO_272 (O_272,N_18125,N_18970);
or UO_273 (O_273,N_19670,N_18366);
nor UO_274 (O_274,N_19534,N_18666);
or UO_275 (O_275,N_18472,N_19711);
or UO_276 (O_276,N_19136,N_18115);
nor UO_277 (O_277,N_18150,N_18857);
nor UO_278 (O_278,N_19247,N_18051);
or UO_279 (O_279,N_19636,N_18504);
nor UO_280 (O_280,N_19379,N_18599);
nor UO_281 (O_281,N_19909,N_19138);
nor UO_282 (O_282,N_18322,N_18585);
nor UO_283 (O_283,N_19761,N_19557);
nor UO_284 (O_284,N_19705,N_18401);
xor UO_285 (O_285,N_19665,N_18142);
nand UO_286 (O_286,N_18260,N_18600);
nand UO_287 (O_287,N_19667,N_19281);
nor UO_288 (O_288,N_18677,N_19738);
xnor UO_289 (O_289,N_18855,N_18040);
and UO_290 (O_290,N_18023,N_18395);
and UO_291 (O_291,N_18668,N_18485);
nor UO_292 (O_292,N_18995,N_19330);
nor UO_293 (O_293,N_18978,N_18298);
or UO_294 (O_294,N_19227,N_18477);
nand UO_295 (O_295,N_18681,N_18376);
nand UO_296 (O_296,N_18777,N_18467);
nand UO_297 (O_297,N_18967,N_19211);
xnor UO_298 (O_298,N_19537,N_18131);
and UO_299 (O_299,N_19219,N_19477);
nand UO_300 (O_300,N_18211,N_18636);
and UO_301 (O_301,N_18749,N_18589);
and UO_302 (O_302,N_19133,N_18152);
nand UO_303 (O_303,N_18323,N_18506);
or UO_304 (O_304,N_19175,N_18925);
xnor UO_305 (O_305,N_18268,N_19878);
nor UO_306 (O_306,N_18483,N_19411);
and UO_307 (O_307,N_18179,N_19032);
nor UO_308 (O_308,N_18694,N_19967);
xnor UO_309 (O_309,N_18439,N_19688);
or UO_310 (O_310,N_18110,N_19126);
xor UO_311 (O_311,N_18562,N_18396);
nor UO_312 (O_312,N_19787,N_18901);
or UO_313 (O_313,N_19614,N_19677);
nand UO_314 (O_314,N_19556,N_19894);
and UO_315 (O_315,N_19099,N_18334);
nor UO_316 (O_316,N_19840,N_18501);
nor UO_317 (O_317,N_19124,N_19606);
nor UO_318 (O_318,N_19755,N_18074);
and UO_319 (O_319,N_18378,N_18276);
or UO_320 (O_320,N_18520,N_19651);
or UO_321 (O_321,N_18015,N_19551);
and UO_322 (O_322,N_18710,N_18555);
nor UO_323 (O_323,N_18342,N_18926);
nor UO_324 (O_324,N_18315,N_19560);
nand UO_325 (O_325,N_18032,N_18206);
and UO_326 (O_326,N_18716,N_18798);
xor UO_327 (O_327,N_18374,N_18960);
nor UO_328 (O_328,N_19195,N_18799);
nor UO_329 (O_329,N_18788,N_18351);
or UO_330 (O_330,N_19797,N_18118);
nor UO_331 (O_331,N_18603,N_19065);
nor UO_332 (O_332,N_18187,N_19053);
and UO_333 (O_333,N_18713,N_19721);
nor UO_334 (O_334,N_19287,N_18417);
or UO_335 (O_335,N_18737,N_18270);
and UO_336 (O_336,N_19835,N_19356);
nor UO_337 (O_337,N_18370,N_18369);
xnor UO_338 (O_338,N_19514,N_19591);
nand UO_339 (O_339,N_18669,N_19956);
and UO_340 (O_340,N_19492,N_19791);
nand UO_341 (O_341,N_18033,N_19658);
or UO_342 (O_342,N_18802,N_18638);
or UO_343 (O_343,N_18054,N_19418);
nor UO_344 (O_344,N_19964,N_18765);
or UO_345 (O_345,N_18392,N_18080);
nand UO_346 (O_346,N_19902,N_18106);
or UO_347 (O_347,N_18557,N_19086);
nand UO_348 (O_348,N_18453,N_19615);
nand UO_349 (O_349,N_18306,N_19831);
or UO_350 (O_350,N_19980,N_18756);
and UO_351 (O_351,N_18252,N_19261);
and UO_352 (O_352,N_19228,N_18588);
nand UO_353 (O_353,N_19789,N_18812);
nand UO_354 (O_354,N_19444,N_18841);
and UO_355 (O_355,N_18934,N_18281);
nor UO_356 (O_356,N_18579,N_18982);
nor UO_357 (O_357,N_19303,N_18456);
nor UO_358 (O_358,N_19603,N_18664);
nor UO_359 (O_359,N_19719,N_18403);
nor UO_360 (O_360,N_18407,N_18507);
and UO_361 (O_361,N_19901,N_19349);
nor UO_362 (O_362,N_19538,N_19236);
or UO_363 (O_363,N_18992,N_19013);
or UO_364 (O_364,N_19162,N_18350);
nor UO_365 (O_365,N_18340,N_19257);
or UO_366 (O_366,N_18736,N_19489);
or UO_367 (O_367,N_19697,N_19662);
nor UO_368 (O_368,N_18283,N_18714);
and UO_369 (O_369,N_19192,N_19610);
xor UO_370 (O_370,N_19449,N_19204);
or UO_371 (O_371,N_18095,N_18380);
or UO_372 (O_372,N_19309,N_19067);
nor UO_373 (O_373,N_18332,N_19565);
nor UO_374 (O_374,N_18762,N_18436);
or UO_375 (O_375,N_19120,N_18063);
and UO_376 (O_376,N_18041,N_18143);
or UO_377 (O_377,N_19663,N_19445);
or UO_378 (O_378,N_18325,N_18622);
and UO_379 (O_379,N_19617,N_18961);
and UO_380 (O_380,N_19254,N_18656);
nand UO_381 (O_381,N_19407,N_18917);
or UO_382 (O_382,N_19470,N_18383);
and UO_383 (O_383,N_19302,N_18174);
xnor UO_384 (O_384,N_18645,N_19199);
or UO_385 (O_385,N_18758,N_18123);
and UO_386 (O_386,N_19267,N_19722);
or UO_387 (O_387,N_18354,N_18912);
nand UO_388 (O_388,N_18647,N_19611);
nor UO_389 (O_389,N_18567,N_19006);
nand UO_390 (O_390,N_18135,N_19354);
nand UO_391 (O_391,N_19872,N_19579);
or UO_392 (O_392,N_19286,N_18674);
nor UO_393 (O_393,N_19076,N_19569);
nor UO_394 (O_394,N_18090,N_18568);
nand UO_395 (O_395,N_18415,N_18827);
and UO_396 (O_396,N_19555,N_18613);
nor UO_397 (O_397,N_19628,N_18521);
or UO_398 (O_398,N_19244,N_18167);
or UO_399 (O_399,N_19384,N_19095);
and UO_400 (O_400,N_19412,N_19406);
nor UO_401 (O_401,N_19751,N_18353);
nor UO_402 (O_402,N_19713,N_18606);
and UO_403 (O_403,N_18265,N_19357);
nor UO_404 (O_404,N_19491,N_18536);
or UO_405 (O_405,N_18346,N_18381);
nor UO_406 (O_406,N_19307,N_18495);
and UO_407 (O_407,N_18695,N_18708);
nor UO_408 (O_408,N_19447,N_19365);
nor UO_409 (O_409,N_19826,N_19837);
nand UO_410 (O_410,N_18387,N_18897);
xor UO_411 (O_411,N_19097,N_19283);
nand UO_412 (O_412,N_18132,N_18973);
or UO_413 (O_413,N_18410,N_19675);
nor UO_414 (O_414,N_19948,N_19769);
nor UO_415 (O_415,N_19986,N_18388);
or UO_416 (O_416,N_18880,N_18047);
or UO_417 (O_417,N_19289,N_19995);
nand UO_418 (O_418,N_18929,N_19581);
nor UO_419 (O_419,N_18005,N_19315);
or UO_420 (O_420,N_19779,N_19638);
nor UO_421 (O_421,N_19018,N_18347);
and UO_422 (O_422,N_18858,N_18833);
nor UO_423 (O_423,N_19564,N_19632);
nand UO_424 (O_424,N_18254,N_19364);
and UO_425 (O_425,N_18031,N_19027);
and UO_426 (O_426,N_19311,N_19156);
nor UO_427 (O_427,N_19417,N_19590);
and UO_428 (O_428,N_19993,N_18486);
or UO_429 (O_429,N_19201,N_19747);
or UO_430 (O_430,N_18990,N_18791);
xor UO_431 (O_431,N_19466,N_19375);
nand UO_432 (O_432,N_18994,N_19821);
or UO_433 (O_433,N_18345,N_18811);
nor UO_434 (O_434,N_19104,N_18199);
or UO_435 (O_435,N_19464,N_18615);
nor UO_436 (O_436,N_19800,N_18312);
nand UO_437 (O_437,N_18572,N_19873);
and UO_438 (O_438,N_19034,N_18581);
nand UO_439 (O_439,N_18073,N_18475);
nand UO_440 (O_440,N_19692,N_18362);
and UO_441 (O_441,N_18726,N_18655);
nand UO_442 (O_442,N_19858,N_19806);
nor UO_443 (O_443,N_19370,N_18902);
nor UO_444 (O_444,N_18731,N_18459);
xnor UO_445 (O_445,N_19701,N_19422);
or UO_446 (O_446,N_18646,N_18921);
or UO_447 (O_447,N_19149,N_19979);
nand UO_448 (O_448,N_18580,N_19758);
nand UO_449 (O_449,N_19844,N_19968);
and UO_450 (O_450,N_18508,N_19893);
nor UO_451 (O_451,N_18985,N_19708);
nor UO_452 (O_452,N_19107,N_18515);
or UO_453 (O_453,N_19448,N_19987);
nor UO_454 (O_454,N_18169,N_19978);
nor UO_455 (O_455,N_19025,N_18156);
and UO_456 (O_456,N_19054,N_18433);
or UO_457 (O_457,N_18119,N_19377);
nor UO_458 (O_458,N_19206,N_18022);
nor UO_459 (O_459,N_18690,N_19359);
nor UO_460 (O_460,N_19361,N_18988);
xnor UO_461 (O_461,N_19327,N_18542);
nand UO_462 (O_462,N_19416,N_18815);
nand UO_463 (O_463,N_18844,N_18886);
nand UO_464 (O_464,N_18006,N_19443);
or UO_465 (O_465,N_19519,N_19329);
nor UO_466 (O_466,N_18687,N_18166);
and UO_467 (O_467,N_19055,N_19678);
nor UO_468 (O_468,N_18605,N_19889);
or UO_469 (O_469,N_19885,N_19112);
xnor UO_470 (O_470,N_19189,N_18450);
nor UO_471 (O_471,N_18928,N_18843);
nand UO_472 (O_472,N_18430,N_18767);
and UO_473 (O_473,N_18966,N_19820);
or UO_474 (O_474,N_19096,N_18224);
nor UO_475 (O_475,N_18389,N_18935);
xor UO_476 (O_476,N_18248,N_19207);
nand UO_477 (O_477,N_18630,N_19060);
nor UO_478 (O_478,N_19325,N_18357);
xnor UO_479 (O_479,N_19511,N_18510);
xor UO_480 (O_480,N_18612,N_19716);
nor UO_481 (O_481,N_18764,N_18384);
nor UO_482 (O_482,N_18335,N_18275);
xnor UO_483 (O_483,N_18061,N_18742);
or UO_484 (O_484,N_18404,N_19572);
xor UO_485 (O_485,N_19225,N_18149);
or UO_486 (O_486,N_18729,N_19352);
or UO_487 (O_487,N_19533,N_18523);
and UO_488 (O_488,N_19210,N_18892);
or UO_489 (O_489,N_18107,N_18161);
xnor UO_490 (O_490,N_18722,N_18652);
xnor UO_491 (O_491,N_19163,N_18130);
nor UO_492 (O_492,N_19546,N_18284);
xor UO_493 (O_493,N_19317,N_19038);
nor UO_494 (O_494,N_18635,N_19850);
nand UO_495 (O_495,N_19442,N_18209);
xnor UO_496 (O_496,N_18078,N_19865);
and UO_497 (O_497,N_19250,N_18675);
nor UO_498 (O_498,N_18364,N_19860);
nor UO_499 (O_499,N_19520,N_18682);
nor UO_500 (O_500,N_18856,N_19910);
nor UO_501 (O_501,N_18128,N_19146);
nand UO_502 (O_502,N_18422,N_19619);
xor UO_503 (O_503,N_19381,N_18246);
or UO_504 (O_504,N_18287,N_18356);
nand UO_505 (O_505,N_18654,N_19395);
or UO_506 (O_506,N_19355,N_18832);
nand UO_507 (O_507,N_18365,N_19724);
or UO_508 (O_508,N_19080,N_19040);
nand UO_509 (O_509,N_19780,N_18825);
or UO_510 (O_510,N_18025,N_19173);
and UO_511 (O_511,N_19213,N_19337);
xnor UO_512 (O_512,N_19413,N_19772);
nand UO_513 (O_513,N_19794,N_18529);
nor UO_514 (O_514,N_18223,N_19051);
or UO_515 (O_515,N_18368,N_19033);
nor UO_516 (O_516,N_18968,N_19552);
and UO_517 (O_517,N_19763,N_19246);
nand UO_518 (O_518,N_19937,N_18979);
nor UO_519 (O_519,N_18134,N_18216);
and UO_520 (O_520,N_19587,N_18660);
xnor UO_521 (O_521,N_19353,N_18423);
xor UO_522 (O_522,N_19386,N_18238);
or UO_523 (O_523,N_19756,N_18558);
xnor UO_524 (O_524,N_19465,N_19525);
or UO_525 (O_525,N_19291,N_18445);
and UO_526 (O_526,N_19063,N_18026);
nand UO_527 (O_527,N_18400,N_19734);
nor UO_528 (O_528,N_18455,N_19374);
nor UO_529 (O_529,N_19178,N_19042);
nor UO_530 (O_530,N_19340,N_18293);
nand UO_531 (O_531,N_19070,N_18952);
nand UO_532 (O_532,N_18294,N_18097);
and UO_533 (O_533,N_18251,N_18112);
and UO_534 (O_534,N_19335,N_18329);
and UO_535 (O_535,N_18482,N_19853);
nand UO_536 (O_536,N_19144,N_18680);
nand UO_537 (O_537,N_19539,N_19548);
or UO_538 (O_538,N_18874,N_19272);
and UO_539 (O_539,N_18763,N_18734);
or UO_540 (O_540,N_18333,N_18532);
nor UO_541 (O_541,N_19313,N_19454);
xnor UO_542 (O_542,N_18019,N_19471);
nor UO_543 (O_543,N_19913,N_18173);
nand UO_544 (O_544,N_19043,N_18259);
or UO_545 (O_545,N_19478,N_18096);
and UO_546 (O_546,N_19938,N_19903);
or UO_547 (O_547,N_18881,N_19334);
nand UO_548 (O_548,N_18709,N_19832);
or UO_549 (O_549,N_19868,N_18348);
or UO_550 (O_550,N_18919,N_18321);
nand UO_551 (O_551,N_19601,N_19500);
nand UO_552 (O_552,N_18727,N_18779);
and UO_553 (O_553,N_19223,N_19849);
and UO_554 (O_554,N_18964,N_19925);
nor UO_555 (O_555,N_19807,N_18093);
and UO_556 (O_556,N_19580,N_19839);
nor UO_557 (O_557,N_19836,N_19602);
nor UO_558 (O_558,N_19859,N_18360);
or UO_559 (O_559,N_19884,N_19245);
or UO_560 (O_560,N_19585,N_19205);
or UO_561 (O_561,N_19389,N_18683);
xor UO_562 (O_562,N_19071,N_19252);
nand UO_563 (O_563,N_19028,N_19589);
and UO_564 (O_564,N_19214,N_18255);
nor UO_565 (O_565,N_18048,N_19946);
or UO_566 (O_566,N_18304,N_18805);
or UO_567 (O_567,N_18465,N_18145);
or UO_568 (O_568,N_18481,N_19958);
or UO_569 (O_569,N_19341,N_18505);
or UO_570 (O_570,N_19728,N_18020);
nor UO_571 (O_571,N_18931,N_18519);
and UO_572 (O_572,N_18511,N_19050);
or UO_573 (O_573,N_19451,N_19597);
and UO_574 (O_574,N_18113,N_19079);
and UO_575 (O_575,N_18850,N_18848);
nand UO_576 (O_576,N_19328,N_19323);
nor UO_577 (O_577,N_19094,N_18653);
nor UO_578 (O_578,N_19529,N_18750);
and UO_579 (O_579,N_18425,N_18847);
or UO_580 (O_580,N_18939,N_19908);
nor UO_581 (O_581,N_19540,N_18540);
and UO_582 (O_582,N_18933,N_19249);
nor UO_583 (O_583,N_18951,N_18793);
xor UO_584 (O_584,N_18141,N_18037);
or UO_585 (O_585,N_18220,N_18704);
nor UO_586 (O_586,N_18168,N_19376);
xnor UO_587 (O_587,N_19197,N_19499);
nor UO_588 (O_588,N_19212,N_19991);
or UO_589 (O_589,N_19816,N_19681);
xor UO_590 (O_590,N_18598,N_19653);
and UO_591 (O_591,N_18735,N_19234);
nor UO_592 (O_592,N_19504,N_18160);
nand UO_593 (O_593,N_19502,N_18975);
nor UO_594 (O_594,N_18871,N_18035);
nand UO_595 (O_595,N_19731,N_19712);
nor UO_596 (O_596,N_18821,N_18620);
or UO_597 (O_597,N_19342,N_19582);
nor UO_598 (O_598,N_18663,N_19951);
xnor UO_599 (O_599,N_19501,N_19649);
nor UO_600 (O_600,N_19388,N_18405);
nor UO_601 (O_601,N_18894,N_18302);
and UO_602 (O_602,N_19896,N_18261);
xnor UO_603 (O_603,N_19509,N_19777);
or UO_604 (O_604,N_19275,N_19191);
xor UO_605 (O_605,N_19456,N_19932);
nor UO_606 (O_606,N_19904,N_19023);
nand UO_607 (O_607,N_18241,N_18122);
xnor UO_608 (O_608,N_19842,N_19237);
and UO_609 (O_609,N_18247,N_18719);
nor UO_610 (O_610,N_18913,N_19770);
and UO_611 (O_611,N_19864,N_19805);
nor UO_612 (O_612,N_18285,N_18480);
or UO_613 (O_613,N_18958,N_19966);
nand UO_614 (O_614,N_19940,N_18773);
and UO_615 (O_615,N_18817,N_19432);
or UO_616 (O_616,N_19284,N_19523);
and UO_617 (O_617,N_19271,N_19209);
nor UO_618 (O_618,N_18232,N_19963);
nor UO_619 (O_619,N_18803,N_18164);
nor UO_620 (O_620,N_19494,N_19396);
nand UO_621 (O_621,N_18918,N_18576);
or UO_622 (O_622,N_18621,N_19224);
nor UO_623 (O_623,N_18940,N_18627);
nand UO_624 (O_624,N_19945,N_19151);
nor UO_625 (O_625,N_19440,N_18191);
nor UO_626 (O_626,N_19621,N_19702);
nor UO_627 (O_627,N_19593,N_18153);
nor UO_628 (O_628,N_19950,N_19266);
nand UO_629 (O_629,N_18030,N_19000);
nor UO_630 (O_630,N_18414,N_19825);
and UO_631 (O_631,N_18591,N_19102);
nand UO_632 (O_632,N_19218,N_18659);
or UO_633 (O_633,N_19190,N_19521);
and UO_634 (O_634,N_18771,N_18176);
or UO_635 (O_635,N_19036,N_19441);
nand UO_636 (O_636,N_18768,N_18068);
and UO_637 (O_637,N_18866,N_18137);
nand UO_638 (O_638,N_19742,N_18538);
xnor UO_639 (O_639,N_18331,N_19600);
nand UO_640 (O_640,N_18200,N_19160);
nor UO_641 (O_641,N_19626,N_18686);
and UO_642 (O_642,N_18637,N_18739);
or UO_643 (O_643,N_18226,N_19784);
and UO_644 (O_644,N_19459,N_18034);
nand UO_645 (O_645,N_19270,N_18759);
or UO_646 (O_646,N_18127,N_19550);
nand UO_647 (O_647,N_19350,N_18441);
nand UO_648 (O_648,N_18087,N_19586);
or UO_649 (O_649,N_18909,N_19083);
and UO_650 (O_650,N_18165,N_19895);
nor UO_651 (O_651,N_18215,N_18789);
nor UO_652 (O_652,N_19139,N_18070);
nand UO_653 (O_653,N_19410,N_18745);
nand UO_654 (O_654,N_18311,N_18181);
or UO_655 (O_655,N_19358,N_18772);
and UO_656 (O_656,N_19117,N_18024);
nand UO_657 (O_657,N_19005,N_18953);
nand UO_658 (O_658,N_19462,N_18962);
or UO_659 (O_659,N_18460,N_18124);
and UO_660 (O_660,N_18932,N_19934);
nand UO_661 (O_661,N_19573,N_19487);
or UO_662 (O_662,N_19882,N_19845);
nor UO_663 (O_663,N_18801,N_19268);
xnor UO_664 (O_664,N_19001,N_18361);
nor UO_665 (O_665,N_18678,N_19748);
nor UO_666 (O_666,N_18094,N_19992);
and UO_667 (O_667,N_19919,N_18060);
or UO_668 (O_668,N_18862,N_18590);
and UO_669 (O_669,N_18657,N_18146);
or UO_670 (O_670,N_19595,N_18464);
nor UO_671 (O_671,N_19962,N_18930);
xor UO_672 (O_672,N_18065,N_18544);
nand UO_673 (O_673,N_18830,N_18597);
nor UO_674 (O_674,N_19841,N_18671);
xor UO_675 (O_675,N_19390,N_18296);
nor UO_676 (O_676,N_19686,N_19704);
nand UO_677 (O_677,N_18924,N_18986);
xor UO_678 (O_678,N_19775,N_19131);
xnor UO_679 (O_679,N_19657,N_18910);
and UO_680 (O_680,N_19513,N_19137);
or UO_681 (O_681,N_19346,N_18527);
xor UO_682 (O_682,N_19339,N_19957);
and UO_683 (O_683,N_19822,N_18017);
nor UO_684 (O_684,N_18101,N_19984);
nand UO_685 (O_685,N_19196,N_19886);
and UO_686 (O_686,N_18056,N_19847);
and UO_687 (O_687,N_18496,N_19744);
xnor UO_688 (O_688,N_18942,N_18443);
xnor UO_689 (O_689,N_18795,N_18526);
nor UO_690 (O_690,N_18946,N_18876);
nand UO_691 (O_691,N_19508,N_19047);
or UO_692 (O_692,N_19288,N_19140);
nand UO_693 (O_693,N_19645,N_19125);
xnor UO_694 (O_694,N_19647,N_19109);
and UO_695 (O_695,N_18608,N_18092);
or UO_696 (O_696,N_19971,N_18320);
and UO_697 (O_697,N_19563,N_19052);
nand UO_698 (O_698,N_19436,N_19659);
nor UO_699 (O_699,N_19256,N_19463);
and UO_700 (O_700,N_19082,N_18541);
nor UO_701 (O_701,N_18148,N_19425);
and UO_702 (O_702,N_18718,N_19776);
nor UO_703 (O_703,N_19202,N_18355);
xnor UO_704 (O_704,N_19802,N_18444);
or UO_705 (O_705,N_18502,N_18289);
nand UO_706 (O_706,N_18705,N_18038);
nor UO_707 (O_707,N_18996,N_18936);
xnor UO_708 (O_708,N_19568,N_18619);
xor UO_709 (O_709,N_18111,N_18829);
nand UO_710 (O_710,N_18665,N_18240);
nor UO_711 (O_711,N_18826,N_18846);
and UO_712 (O_712,N_18870,N_19718);
and UO_713 (O_713,N_19171,N_18503);
or UO_714 (O_714,N_18741,N_18691);
and UO_715 (O_715,N_18290,N_19811);
and UO_716 (O_716,N_18873,N_19929);
nor UO_717 (O_717,N_18089,N_18564);
nand UO_718 (O_718,N_18937,N_18954);
or UO_719 (O_719,N_18614,N_18412);
and UO_720 (O_720,N_19424,N_18155);
xor UO_721 (O_721,N_19729,N_19004);
nor UO_722 (O_722,N_18108,N_18194);
and UO_723 (O_723,N_18867,N_19372);
xor UO_724 (O_724,N_19921,N_19092);
or UO_725 (O_725,N_19153,N_19399);
nor UO_726 (O_726,N_18426,N_18253);
nor UO_727 (O_727,N_19248,N_19627);
nor UO_728 (O_728,N_19308,N_18154);
nand UO_729 (O_729,N_19804,N_19899);
nor UO_730 (O_730,N_19703,N_18828);
nor UO_731 (O_731,N_19016,N_19164);
and UO_732 (O_732,N_19176,N_18543);
and UO_733 (O_733,N_19498,N_18554);
xor UO_734 (O_734,N_18227,N_19188);
nand UO_735 (O_735,N_19455,N_19198);
or UO_736 (O_736,N_18084,N_18679);
nor UO_737 (O_737,N_18029,N_18751);
or UO_738 (O_738,N_19812,N_18887);
and UO_739 (O_739,N_18295,N_19907);
nand UO_740 (O_740,N_19115,N_18574);
and UO_741 (O_741,N_18711,N_19596);
xor UO_742 (O_742,N_18545,N_18911);
nor UO_743 (O_743,N_18288,N_18105);
nand UO_744 (O_744,N_18016,N_18217);
or UO_745 (O_745,N_19624,N_18406);
nor UO_746 (O_746,N_19259,N_18498);
or UO_747 (O_747,N_19592,N_19280);
nor UO_748 (O_748,N_18689,N_19351);
xor UO_749 (O_749,N_19493,N_19656);
nor UO_750 (O_750,N_19002,N_19879);
or UO_751 (O_751,N_18120,N_18754);
or UO_752 (O_752,N_19643,N_19578);
nand UO_753 (O_753,N_18488,N_18644);
and UO_754 (O_754,N_18890,N_18085);
xnor UO_755 (O_755,N_18976,N_19947);
nor UO_756 (O_756,N_18908,N_19542);
nand UO_757 (O_757,N_19409,N_18239);
or UO_758 (O_758,N_18067,N_18720);
nand UO_759 (O_759,N_18800,N_19888);
nand UO_760 (O_760,N_19544,N_18104);
nand UO_761 (O_761,N_19846,N_19654);
nand UO_762 (O_762,N_18309,N_18250);
and UO_763 (O_763,N_19238,N_18571);
or UO_764 (O_764,N_19119,N_19646);
xnor UO_765 (O_765,N_19405,N_18204);
or UO_766 (O_766,N_19730,N_18699);
xnor UO_767 (O_767,N_18697,N_19558);
or UO_768 (O_768,N_19419,N_18071);
or UO_769 (O_769,N_19574,N_19700);
nand UO_770 (O_770,N_19158,N_18162);
nor UO_771 (O_771,N_19871,N_18140);
xor UO_772 (O_772,N_19706,N_18766);
or UO_773 (O_773,N_19843,N_18981);
nand UO_774 (O_774,N_19547,N_19854);
and UO_775 (O_775,N_19129,N_18277);
nand UO_776 (O_776,N_18297,N_18834);
nand UO_777 (O_777,N_18879,N_19019);
and UO_778 (O_778,N_18228,N_19305);
xor UO_779 (O_779,N_19180,N_18725);
nor UO_780 (O_780,N_19398,N_19965);
xnor UO_781 (O_781,N_19526,N_19942);
nand UO_782 (O_782,N_18316,N_18820);
nor UO_783 (O_783,N_18786,N_18878);
nand UO_784 (O_784,N_18317,N_18185);
nor UO_785 (O_785,N_18424,N_18234);
nand UO_786 (O_786,N_19022,N_18397);
or UO_787 (O_787,N_19512,N_19715);
nor UO_788 (O_788,N_18651,N_19255);
nor UO_789 (O_789,N_18706,N_18965);
or UO_790 (O_790,N_19161,N_19426);
and UO_791 (O_791,N_19783,N_18738);
or UO_792 (O_792,N_19928,N_19997);
nor UO_793 (O_793,N_19306,N_18658);
nor UO_794 (O_794,N_19815,N_18927);
nand UO_795 (O_795,N_19285,N_19294);
and UO_796 (O_796,N_18144,N_19698);
and UO_797 (O_797,N_18633,N_19790);
nor UO_798 (O_798,N_18057,N_18157);
and UO_799 (O_799,N_18466,N_19193);
and UO_800 (O_800,N_19397,N_19944);
nor UO_801 (O_801,N_19239,N_19960);
and UO_802 (O_802,N_18769,N_18787);
or UO_803 (O_803,N_19900,N_18676);
nand UO_804 (O_804,N_19874,N_18774);
or UO_805 (O_805,N_19122,N_19240);
or UO_806 (O_806,N_19834,N_19010);
and UO_807 (O_807,N_18569,N_19917);
xor UO_808 (O_808,N_19061,N_18280);
or UO_809 (O_809,N_18573,N_18700);
nand UO_810 (O_810,N_19141,N_18310);
nand UO_811 (O_811,N_19618,N_19045);
xnor UO_812 (O_812,N_19015,N_18207);
xnor UO_813 (O_813,N_18851,N_18170);
nand UO_814 (O_814,N_19392,N_19260);
and UO_815 (O_815,N_18673,N_19915);
nor UO_816 (O_816,N_18286,N_19998);
xor UO_817 (O_817,N_19536,N_19622);
or UO_818 (O_818,N_19400,N_18075);
nand UO_819 (O_819,N_18434,N_18724);
or UO_820 (O_820,N_19976,N_18243);
xnor UO_821 (O_821,N_18461,N_18454);
xnor UO_822 (O_822,N_18163,N_19475);
or UO_823 (O_823,N_18103,N_19562);
and UO_824 (O_824,N_18743,N_18233);
nand UO_825 (O_825,N_19608,N_18895);
nor UO_826 (O_826,N_18703,N_19605);
xnor UO_827 (O_827,N_19093,N_18344);
or UO_828 (O_828,N_18639,N_19402);
or UO_829 (O_829,N_18359,N_19318);
nor UO_830 (O_830,N_19231,N_18898);
xnor UO_831 (O_831,N_19435,N_19810);
xnor UO_832 (O_832,N_19132,N_19226);
nand UO_833 (O_833,N_18447,N_18349);
and UO_834 (O_834,N_18797,N_18842);
xnor UO_835 (O_835,N_18197,N_19105);
and UO_836 (O_836,N_19007,N_19648);
xor UO_837 (O_837,N_19074,N_18341);
or UO_838 (O_838,N_19265,N_19075);
or UO_839 (O_839,N_19527,N_19142);
nand UO_840 (O_840,N_19008,N_19760);
or UO_841 (O_841,N_18196,N_19695);
nand UO_842 (O_842,N_18617,N_19766);
nand UO_843 (O_843,N_18794,N_19641);
or UO_844 (O_844,N_19114,N_18126);
nor UO_845 (O_845,N_18534,N_19666);
nand UO_846 (O_846,N_19217,N_19530);
or UO_847 (O_847,N_19157,N_19253);
or UO_848 (O_848,N_18578,N_19380);
nand UO_849 (O_849,N_19088,N_18058);
and UO_850 (O_850,N_19215,N_19200);
or UO_851 (O_851,N_19607,N_18129);
and UO_852 (O_852,N_18303,N_19460);
nor UO_853 (O_853,N_19179,N_18413);
nor UO_854 (O_854,N_19030,N_18099);
xor UO_855 (O_855,N_18552,N_18300);
nor UO_856 (O_856,N_18860,N_18528);
nor UO_857 (O_857,N_18372,N_19059);
and UO_858 (O_858,N_18491,N_19710);
and UO_859 (O_859,N_18062,N_19304);
or UO_860 (O_860,N_18045,N_18476);
nand UO_861 (O_861,N_19430,N_19064);
nor UO_862 (O_862,N_18753,N_19496);
or UO_863 (O_863,N_19851,N_19829);
and UO_864 (O_864,N_18957,N_18177);
nor UO_865 (O_865,N_19737,N_18650);
nand UO_866 (O_866,N_18478,N_19570);
nor UO_867 (O_867,N_18533,N_18036);
nand UO_868 (O_868,N_19746,N_18915);
xor UO_869 (O_869,N_19020,N_18701);
nor UO_870 (O_870,N_19892,N_18319);
and UO_871 (O_871,N_19336,N_18274);
nor UO_872 (O_872,N_18305,N_18672);
nand UO_873 (O_873,N_19168,N_18236);
nand UO_874 (O_874,N_18640,N_18046);
or UO_875 (O_875,N_19316,N_19676);
or UO_876 (O_876,N_19796,N_19685);
nand UO_877 (O_877,N_19808,N_18500);
and UO_878 (O_878,N_18780,N_18391);
nor UO_879 (O_879,N_19243,N_19516);
or UO_880 (O_880,N_19011,N_19343);
nor UO_881 (O_881,N_18813,N_18377);
nand UO_882 (O_882,N_19745,N_19145);
or UO_883 (O_883,N_18421,N_18007);
xnor UO_884 (O_884,N_18808,N_19314);
and UO_885 (O_885,N_18102,N_18883);
nand UO_886 (O_886,N_18810,N_19181);
and UO_887 (O_887,N_18565,N_19773);
or UO_888 (O_888,N_18575,N_18292);
nor UO_889 (O_889,N_19733,N_19876);
and UO_890 (O_890,N_19057,N_19717);
or UO_891 (O_891,N_18944,N_19331);
and UO_892 (O_892,N_19566,N_18631);
nor UO_893 (O_893,N_18884,N_18203);
xnor UO_894 (O_894,N_18192,N_18499);
or UO_895 (O_895,N_18938,N_18717);
or UO_896 (O_896,N_19629,N_19081);
nor UO_897 (O_897,N_18566,N_19506);
nand UO_898 (O_898,N_19798,N_18634);
nand UO_899 (O_899,N_19474,N_18003);
nand UO_900 (O_900,N_18561,N_19973);
or UO_901 (O_901,N_18730,N_18468);
nand UO_902 (O_902,N_19056,N_18428);
nand UO_903 (O_903,N_18583,N_19535);
nor UO_904 (O_904,N_19594,N_18611);
nand UO_905 (O_905,N_18079,N_19972);
or UO_906 (O_906,N_19479,N_18178);
or UO_907 (O_907,N_19959,N_19495);
xnor UO_908 (O_908,N_19830,N_19367);
nor UO_909 (O_909,N_18906,N_18993);
xor UO_910 (O_910,N_19736,N_19923);
nor UO_911 (O_911,N_19828,N_19749);
or UO_912 (O_912,N_19862,N_19421);
nand UO_913 (O_913,N_19048,N_18783);
xor UO_914 (O_914,N_19881,N_18338);
nand UO_915 (O_915,N_19817,N_19680);
nor UO_916 (O_916,N_18839,N_19898);
nor UO_917 (O_917,N_18907,N_19974);
and UO_918 (O_918,N_19345,N_19024);
and UO_919 (O_919,N_18998,N_19087);
nor UO_920 (O_920,N_19507,N_19869);
nor UO_921 (O_921,N_18723,N_19497);
and UO_922 (O_922,N_18899,N_18109);
or UO_923 (O_923,N_19633,N_18473);
nand UO_924 (O_924,N_19420,N_18956);
or UO_925 (O_925,N_19490,N_19434);
nand UO_926 (O_926,N_19799,N_18643);
nor UO_927 (O_927,N_19985,N_18121);
xor UO_928 (O_928,N_19723,N_18814);
or UO_929 (O_929,N_19073,N_18971);
xnor UO_930 (O_930,N_19750,N_19332);
or UO_931 (O_931,N_18702,N_19543);
nand UO_932 (O_932,N_18171,N_19363);
nand UO_933 (O_933,N_19989,N_18081);
nand UO_934 (O_934,N_18218,N_18158);
nand UO_935 (O_935,N_18053,N_18072);
nand UO_936 (O_936,N_19588,N_18307);
nand UO_937 (O_937,N_19890,N_18432);
nand UO_938 (O_938,N_18076,N_19683);
xnor UO_939 (O_939,N_19759,N_19338);
nor UO_940 (O_940,N_18429,N_18900);
nand UO_941 (O_941,N_18626,N_18624);
and UO_942 (O_942,N_18875,N_18548);
nor UO_943 (O_943,N_19439,N_19554);
nor UO_944 (O_944,N_18649,N_19221);
nor UO_945 (O_945,N_18980,N_18219);
nor UO_946 (O_946,N_19457,N_18420);
nor UO_947 (O_947,N_18308,N_19824);
and UO_948 (O_948,N_18692,N_18744);
and UO_949 (O_949,N_18151,N_18642);
xor UO_950 (O_950,N_19461,N_19583);
nor UO_951 (O_951,N_19241,N_18011);
nand UO_952 (O_952,N_19299,N_19549);
xor UO_953 (O_953,N_18172,N_18854);
or UO_954 (O_954,N_18594,N_18609);
and UO_955 (O_955,N_19021,N_19612);
and UO_956 (O_956,N_19786,N_19584);
and UO_957 (O_957,N_18231,N_19875);
or UO_958 (O_958,N_19793,N_19480);
nand UO_959 (O_959,N_19813,N_18818);
nand UO_960 (O_960,N_18493,N_18607);
nand UO_961 (O_961,N_19106,N_18760);
or UO_962 (O_962,N_19041,N_18816);
and UO_963 (O_963,N_18922,N_19880);
nand UO_964 (O_964,N_19912,N_19969);
nand UO_965 (O_965,N_18963,N_19403);
nand UO_966 (O_966,N_19150,N_18868);
or UO_967 (O_967,N_18549,N_19404);
nand UO_968 (O_968,N_19127,N_18457);
nand UO_969 (O_969,N_18139,N_19541);
xnor UO_970 (O_970,N_19528,N_19165);
xor UO_971 (O_971,N_18479,N_19220);
nor UO_972 (O_972,N_18761,N_19113);
or UO_973 (O_973,N_18945,N_18837);
nand UO_974 (O_974,N_18667,N_19433);
and UO_975 (O_975,N_18463,N_18610);
or UO_976 (O_976,N_18052,N_18616);
nand UO_977 (O_977,N_18494,N_18835);
nor UO_978 (O_978,N_18328,N_18343);
nor UO_979 (O_979,N_19827,N_19935);
xnor UO_980 (O_980,N_18419,N_19682);
nand UO_981 (O_981,N_18512,N_18997);
nand UO_982 (O_982,N_18877,N_18865);
or UO_983 (O_983,N_18596,N_18442);
nand UO_984 (O_984,N_19764,N_19684);
and UO_985 (O_985,N_18707,N_18462);
nor UO_986 (O_986,N_19740,N_19771);
nor UO_987 (O_987,N_18427,N_18269);
nor UO_988 (O_988,N_19522,N_18732);
or UO_989 (O_989,N_19293,N_19673);
and UO_990 (O_990,N_19366,N_19035);
nand UO_991 (O_991,N_18398,N_18551);
nand UO_992 (O_992,N_18399,N_18256);
nand UO_993 (O_993,N_19644,N_18531);
xor UO_994 (O_994,N_19634,N_19689);
and UO_995 (O_995,N_19312,N_19394);
and UO_996 (O_996,N_18272,N_19696);
nor UO_997 (O_997,N_18027,N_18367);
and UO_998 (O_998,N_18086,N_19714);
nor UO_999 (O_999,N_19863,N_19282);
xor UO_1000 (O_1000,N_19356,N_19407);
nor UO_1001 (O_1001,N_18360,N_19663);
nand UO_1002 (O_1002,N_19012,N_18421);
nand UO_1003 (O_1003,N_19040,N_19449);
and UO_1004 (O_1004,N_18616,N_18300);
and UO_1005 (O_1005,N_19947,N_19379);
or UO_1006 (O_1006,N_19270,N_19183);
or UO_1007 (O_1007,N_19011,N_18833);
nand UO_1008 (O_1008,N_19032,N_18156);
nor UO_1009 (O_1009,N_18355,N_19822);
and UO_1010 (O_1010,N_19452,N_18171);
xor UO_1011 (O_1011,N_18806,N_19422);
xor UO_1012 (O_1012,N_19514,N_18036);
nor UO_1013 (O_1013,N_18285,N_19506);
and UO_1014 (O_1014,N_18086,N_19022);
nor UO_1015 (O_1015,N_19525,N_19031);
nor UO_1016 (O_1016,N_19930,N_18172);
nor UO_1017 (O_1017,N_19324,N_18384);
xnor UO_1018 (O_1018,N_18161,N_18451);
nand UO_1019 (O_1019,N_18093,N_19685);
or UO_1020 (O_1020,N_18481,N_18600);
or UO_1021 (O_1021,N_19521,N_18555);
nor UO_1022 (O_1022,N_19478,N_19718);
nor UO_1023 (O_1023,N_18578,N_19193);
and UO_1024 (O_1024,N_19550,N_19628);
nand UO_1025 (O_1025,N_19064,N_18397);
or UO_1026 (O_1026,N_19386,N_19426);
or UO_1027 (O_1027,N_19488,N_19231);
nand UO_1028 (O_1028,N_18223,N_19773);
xnor UO_1029 (O_1029,N_18433,N_19671);
xor UO_1030 (O_1030,N_19215,N_19286);
nor UO_1031 (O_1031,N_19702,N_18831);
and UO_1032 (O_1032,N_19396,N_18139);
nor UO_1033 (O_1033,N_18315,N_19013);
or UO_1034 (O_1034,N_18828,N_18851);
nor UO_1035 (O_1035,N_18876,N_19097);
or UO_1036 (O_1036,N_19345,N_18823);
xnor UO_1037 (O_1037,N_18373,N_19113);
and UO_1038 (O_1038,N_19935,N_18336);
xor UO_1039 (O_1039,N_18772,N_18593);
nor UO_1040 (O_1040,N_19542,N_19068);
nor UO_1041 (O_1041,N_18280,N_19225);
and UO_1042 (O_1042,N_18816,N_18661);
nand UO_1043 (O_1043,N_19640,N_18576);
or UO_1044 (O_1044,N_18234,N_18546);
nor UO_1045 (O_1045,N_19523,N_19876);
xor UO_1046 (O_1046,N_19539,N_18048);
nand UO_1047 (O_1047,N_18728,N_18910);
xor UO_1048 (O_1048,N_18490,N_19145);
or UO_1049 (O_1049,N_18474,N_18345);
and UO_1050 (O_1050,N_18638,N_18383);
nand UO_1051 (O_1051,N_18436,N_18467);
xnor UO_1052 (O_1052,N_18470,N_19765);
nand UO_1053 (O_1053,N_18202,N_18023);
nor UO_1054 (O_1054,N_18837,N_18666);
or UO_1055 (O_1055,N_19287,N_19215);
and UO_1056 (O_1056,N_18434,N_19542);
and UO_1057 (O_1057,N_19442,N_18178);
nor UO_1058 (O_1058,N_18406,N_19051);
and UO_1059 (O_1059,N_19553,N_18792);
nand UO_1060 (O_1060,N_18384,N_19509);
xor UO_1061 (O_1061,N_19163,N_19661);
nand UO_1062 (O_1062,N_19334,N_19949);
nand UO_1063 (O_1063,N_18397,N_18234);
nor UO_1064 (O_1064,N_19179,N_18792);
and UO_1065 (O_1065,N_18332,N_18558);
nand UO_1066 (O_1066,N_19750,N_18109);
nor UO_1067 (O_1067,N_18006,N_18711);
xor UO_1068 (O_1068,N_18407,N_18403);
and UO_1069 (O_1069,N_19545,N_18175);
and UO_1070 (O_1070,N_19224,N_18981);
nand UO_1071 (O_1071,N_19137,N_19657);
nor UO_1072 (O_1072,N_19896,N_18563);
nor UO_1073 (O_1073,N_18182,N_19906);
nand UO_1074 (O_1074,N_18919,N_18617);
nor UO_1075 (O_1075,N_19966,N_19742);
and UO_1076 (O_1076,N_19076,N_19278);
and UO_1077 (O_1077,N_18417,N_19029);
nand UO_1078 (O_1078,N_19324,N_19743);
nor UO_1079 (O_1079,N_18387,N_19132);
nor UO_1080 (O_1080,N_19160,N_18455);
xnor UO_1081 (O_1081,N_19961,N_18840);
nor UO_1082 (O_1082,N_19324,N_19096);
and UO_1083 (O_1083,N_19673,N_18563);
or UO_1084 (O_1084,N_19502,N_19240);
or UO_1085 (O_1085,N_19232,N_18688);
or UO_1086 (O_1086,N_18328,N_18519);
and UO_1087 (O_1087,N_19141,N_18421);
nand UO_1088 (O_1088,N_19343,N_19986);
nor UO_1089 (O_1089,N_19252,N_19293);
and UO_1090 (O_1090,N_18616,N_19407);
and UO_1091 (O_1091,N_19292,N_19632);
nor UO_1092 (O_1092,N_18362,N_18729);
and UO_1093 (O_1093,N_18863,N_19447);
and UO_1094 (O_1094,N_18744,N_18007);
nand UO_1095 (O_1095,N_19385,N_19466);
and UO_1096 (O_1096,N_19686,N_18395);
and UO_1097 (O_1097,N_19688,N_19373);
and UO_1098 (O_1098,N_19808,N_18762);
and UO_1099 (O_1099,N_19650,N_18202);
and UO_1100 (O_1100,N_18263,N_18359);
nand UO_1101 (O_1101,N_18931,N_19170);
nor UO_1102 (O_1102,N_19606,N_19087);
and UO_1103 (O_1103,N_18533,N_19673);
nand UO_1104 (O_1104,N_19475,N_18545);
nor UO_1105 (O_1105,N_19541,N_19166);
or UO_1106 (O_1106,N_19525,N_18899);
or UO_1107 (O_1107,N_19585,N_19684);
or UO_1108 (O_1108,N_19209,N_19087);
nor UO_1109 (O_1109,N_19964,N_18734);
or UO_1110 (O_1110,N_19241,N_19831);
nand UO_1111 (O_1111,N_19813,N_18199);
or UO_1112 (O_1112,N_19147,N_19339);
nor UO_1113 (O_1113,N_19136,N_19584);
and UO_1114 (O_1114,N_18997,N_18014);
xor UO_1115 (O_1115,N_18210,N_19188);
nor UO_1116 (O_1116,N_18051,N_19641);
nor UO_1117 (O_1117,N_19640,N_19175);
nand UO_1118 (O_1118,N_19601,N_19497);
nand UO_1119 (O_1119,N_18142,N_18975);
nor UO_1120 (O_1120,N_19564,N_19952);
nand UO_1121 (O_1121,N_19663,N_19953);
and UO_1122 (O_1122,N_19168,N_18556);
and UO_1123 (O_1123,N_18893,N_18466);
and UO_1124 (O_1124,N_19529,N_19400);
or UO_1125 (O_1125,N_18481,N_19568);
or UO_1126 (O_1126,N_18803,N_18881);
xor UO_1127 (O_1127,N_18174,N_18501);
or UO_1128 (O_1128,N_18404,N_18291);
xor UO_1129 (O_1129,N_19084,N_19266);
nand UO_1130 (O_1130,N_19041,N_19252);
nand UO_1131 (O_1131,N_19483,N_19810);
or UO_1132 (O_1132,N_18495,N_19792);
xnor UO_1133 (O_1133,N_18073,N_18941);
and UO_1134 (O_1134,N_18177,N_19568);
or UO_1135 (O_1135,N_18675,N_18154);
and UO_1136 (O_1136,N_19754,N_18227);
and UO_1137 (O_1137,N_18578,N_19833);
or UO_1138 (O_1138,N_19285,N_18497);
xor UO_1139 (O_1139,N_19963,N_19406);
nand UO_1140 (O_1140,N_19685,N_18605);
nand UO_1141 (O_1141,N_19490,N_19599);
nor UO_1142 (O_1142,N_18980,N_19950);
nor UO_1143 (O_1143,N_18709,N_18130);
nand UO_1144 (O_1144,N_19437,N_18377);
or UO_1145 (O_1145,N_18779,N_18623);
and UO_1146 (O_1146,N_18729,N_19713);
nor UO_1147 (O_1147,N_19596,N_18433);
or UO_1148 (O_1148,N_19375,N_18764);
or UO_1149 (O_1149,N_19616,N_19816);
or UO_1150 (O_1150,N_18194,N_18689);
nand UO_1151 (O_1151,N_19946,N_18594);
and UO_1152 (O_1152,N_18570,N_18868);
and UO_1153 (O_1153,N_19511,N_19131);
or UO_1154 (O_1154,N_19350,N_19877);
nand UO_1155 (O_1155,N_19019,N_19420);
and UO_1156 (O_1156,N_18980,N_18904);
or UO_1157 (O_1157,N_19167,N_18131);
nand UO_1158 (O_1158,N_18478,N_19752);
or UO_1159 (O_1159,N_19350,N_18543);
nand UO_1160 (O_1160,N_18053,N_19286);
and UO_1161 (O_1161,N_18268,N_18640);
nand UO_1162 (O_1162,N_19168,N_19875);
nor UO_1163 (O_1163,N_18512,N_19619);
nand UO_1164 (O_1164,N_19996,N_18895);
nand UO_1165 (O_1165,N_19922,N_19338);
or UO_1166 (O_1166,N_19426,N_18863);
and UO_1167 (O_1167,N_19120,N_19210);
nand UO_1168 (O_1168,N_19592,N_18153);
and UO_1169 (O_1169,N_18417,N_19142);
or UO_1170 (O_1170,N_18236,N_19989);
nor UO_1171 (O_1171,N_18194,N_18248);
or UO_1172 (O_1172,N_19478,N_18376);
or UO_1173 (O_1173,N_18113,N_18250);
nand UO_1174 (O_1174,N_18295,N_19342);
nor UO_1175 (O_1175,N_19238,N_18830);
nand UO_1176 (O_1176,N_18537,N_18932);
nor UO_1177 (O_1177,N_18166,N_19179);
nand UO_1178 (O_1178,N_18654,N_19307);
xor UO_1179 (O_1179,N_19287,N_19545);
and UO_1180 (O_1180,N_18457,N_18523);
or UO_1181 (O_1181,N_18101,N_18087);
nor UO_1182 (O_1182,N_19499,N_18520);
nor UO_1183 (O_1183,N_18468,N_19260);
nand UO_1184 (O_1184,N_19800,N_19856);
nand UO_1185 (O_1185,N_19000,N_18476);
nand UO_1186 (O_1186,N_18606,N_19997);
and UO_1187 (O_1187,N_18471,N_19930);
and UO_1188 (O_1188,N_19380,N_19762);
or UO_1189 (O_1189,N_19772,N_19240);
nor UO_1190 (O_1190,N_19996,N_19257);
xnor UO_1191 (O_1191,N_19279,N_18374);
nand UO_1192 (O_1192,N_18575,N_18324);
nand UO_1193 (O_1193,N_19121,N_19546);
nor UO_1194 (O_1194,N_19137,N_18248);
nor UO_1195 (O_1195,N_18484,N_18306);
or UO_1196 (O_1196,N_18813,N_18106);
and UO_1197 (O_1197,N_19833,N_18566);
nor UO_1198 (O_1198,N_18393,N_18273);
and UO_1199 (O_1199,N_19554,N_19521);
and UO_1200 (O_1200,N_18921,N_18092);
and UO_1201 (O_1201,N_19902,N_18412);
and UO_1202 (O_1202,N_18579,N_18268);
nand UO_1203 (O_1203,N_18701,N_19475);
and UO_1204 (O_1204,N_19351,N_19250);
nor UO_1205 (O_1205,N_18947,N_19581);
nand UO_1206 (O_1206,N_19938,N_18167);
nor UO_1207 (O_1207,N_18350,N_19034);
nand UO_1208 (O_1208,N_19683,N_19350);
nand UO_1209 (O_1209,N_18310,N_19288);
nor UO_1210 (O_1210,N_19974,N_18700);
and UO_1211 (O_1211,N_19375,N_19882);
nor UO_1212 (O_1212,N_19812,N_19486);
nor UO_1213 (O_1213,N_19688,N_18975);
xnor UO_1214 (O_1214,N_18515,N_18182);
nor UO_1215 (O_1215,N_19446,N_19644);
and UO_1216 (O_1216,N_19382,N_19846);
and UO_1217 (O_1217,N_18597,N_18107);
and UO_1218 (O_1218,N_19619,N_18462);
nand UO_1219 (O_1219,N_19379,N_18569);
or UO_1220 (O_1220,N_19233,N_19769);
or UO_1221 (O_1221,N_19349,N_19329);
nand UO_1222 (O_1222,N_19669,N_19107);
nand UO_1223 (O_1223,N_19758,N_18583);
or UO_1224 (O_1224,N_18539,N_18530);
and UO_1225 (O_1225,N_18719,N_19261);
nor UO_1226 (O_1226,N_19620,N_18940);
nor UO_1227 (O_1227,N_18468,N_18594);
or UO_1228 (O_1228,N_19435,N_19769);
xnor UO_1229 (O_1229,N_18784,N_19180);
or UO_1230 (O_1230,N_18567,N_18222);
nand UO_1231 (O_1231,N_18535,N_18300);
nand UO_1232 (O_1232,N_18546,N_18911);
or UO_1233 (O_1233,N_19430,N_19629);
nor UO_1234 (O_1234,N_19332,N_19543);
nor UO_1235 (O_1235,N_19109,N_18034);
and UO_1236 (O_1236,N_18760,N_19217);
or UO_1237 (O_1237,N_18409,N_18293);
nor UO_1238 (O_1238,N_19347,N_18775);
or UO_1239 (O_1239,N_18137,N_19422);
nand UO_1240 (O_1240,N_19329,N_19054);
nor UO_1241 (O_1241,N_18966,N_18008);
and UO_1242 (O_1242,N_18042,N_19599);
nand UO_1243 (O_1243,N_19688,N_18455);
xnor UO_1244 (O_1244,N_19412,N_18018);
xnor UO_1245 (O_1245,N_18168,N_18634);
or UO_1246 (O_1246,N_18103,N_18615);
and UO_1247 (O_1247,N_19349,N_19515);
or UO_1248 (O_1248,N_18073,N_18635);
or UO_1249 (O_1249,N_19424,N_19788);
or UO_1250 (O_1250,N_19243,N_18589);
nor UO_1251 (O_1251,N_18107,N_19036);
and UO_1252 (O_1252,N_19992,N_18474);
and UO_1253 (O_1253,N_18196,N_18402);
or UO_1254 (O_1254,N_18576,N_19082);
nor UO_1255 (O_1255,N_18990,N_18160);
and UO_1256 (O_1256,N_18995,N_18028);
nor UO_1257 (O_1257,N_18717,N_19499);
or UO_1258 (O_1258,N_19665,N_18411);
or UO_1259 (O_1259,N_19511,N_18734);
or UO_1260 (O_1260,N_19865,N_18692);
and UO_1261 (O_1261,N_18106,N_18718);
nor UO_1262 (O_1262,N_18635,N_19454);
and UO_1263 (O_1263,N_19432,N_19101);
or UO_1264 (O_1264,N_19921,N_19320);
and UO_1265 (O_1265,N_18994,N_18776);
and UO_1266 (O_1266,N_18154,N_19932);
xnor UO_1267 (O_1267,N_19848,N_18075);
nor UO_1268 (O_1268,N_19767,N_19359);
and UO_1269 (O_1269,N_19097,N_18040);
nand UO_1270 (O_1270,N_18142,N_18854);
nand UO_1271 (O_1271,N_19823,N_18631);
and UO_1272 (O_1272,N_18979,N_19639);
nand UO_1273 (O_1273,N_18048,N_19830);
or UO_1274 (O_1274,N_18923,N_18449);
nor UO_1275 (O_1275,N_19700,N_18011);
or UO_1276 (O_1276,N_19792,N_18538);
or UO_1277 (O_1277,N_18827,N_19150);
or UO_1278 (O_1278,N_19981,N_18151);
or UO_1279 (O_1279,N_19513,N_18423);
nor UO_1280 (O_1280,N_19232,N_18053);
or UO_1281 (O_1281,N_19410,N_19671);
nand UO_1282 (O_1282,N_19249,N_19944);
or UO_1283 (O_1283,N_19335,N_19068);
and UO_1284 (O_1284,N_18203,N_18586);
xnor UO_1285 (O_1285,N_19521,N_18319);
nand UO_1286 (O_1286,N_18714,N_19994);
nand UO_1287 (O_1287,N_18362,N_19907);
nor UO_1288 (O_1288,N_18149,N_18296);
or UO_1289 (O_1289,N_18090,N_18413);
nor UO_1290 (O_1290,N_19295,N_18779);
xnor UO_1291 (O_1291,N_19485,N_18080);
or UO_1292 (O_1292,N_19219,N_18773);
nor UO_1293 (O_1293,N_19379,N_19284);
and UO_1294 (O_1294,N_18658,N_19417);
nand UO_1295 (O_1295,N_19257,N_19639);
or UO_1296 (O_1296,N_19789,N_18768);
or UO_1297 (O_1297,N_18087,N_19868);
or UO_1298 (O_1298,N_18230,N_18028);
and UO_1299 (O_1299,N_18157,N_19733);
xor UO_1300 (O_1300,N_18857,N_18548);
or UO_1301 (O_1301,N_18210,N_18373);
nand UO_1302 (O_1302,N_18029,N_18105);
nand UO_1303 (O_1303,N_19062,N_18865);
nor UO_1304 (O_1304,N_18035,N_18904);
or UO_1305 (O_1305,N_18679,N_19188);
and UO_1306 (O_1306,N_19692,N_19060);
and UO_1307 (O_1307,N_18138,N_18990);
nand UO_1308 (O_1308,N_19324,N_19959);
and UO_1309 (O_1309,N_18795,N_18125);
nor UO_1310 (O_1310,N_19347,N_18024);
and UO_1311 (O_1311,N_19131,N_18932);
xor UO_1312 (O_1312,N_18868,N_19452);
nor UO_1313 (O_1313,N_18744,N_19334);
xnor UO_1314 (O_1314,N_18163,N_18451);
and UO_1315 (O_1315,N_19929,N_19619);
nand UO_1316 (O_1316,N_18816,N_18364);
nor UO_1317 (O_1317,N_19993,N_18740);
nor UO_1318 (O_1318,N_19001,N_19319);
or UO_1319 (O_1319,N_18465,N_18893);
or UO_1320 (O_1320,N_19645,N_18334);
nand UO_1321 (O_1321,N_19820,N_19320);
nand UO_1322 (O_1322,N_19744,N_19323);
nand UO_1323 (O_1323,N_18074,N_19111);
nor UO_1324 (O_1324,N_19131,N_19387);
xnor UO_1325 (O_1325,N_19827,N_19304);
nor UO_1326 (O_1326,N_18784,N_18698);
nor UO_1327 (O_1327,N_19086,N_18441);
nand UO_1328 (O_1328,N_18965,N_18278);
nand UO_1329 (O_1329,N_18188,N_19200);
xnor UO_1330 (O_1330,N_18079,N_19500);
or UO_1331 (O_1331,N_19288,N_18323);
xnor UO_1332 (O_1332,N_18325,N_18588);
or UO_1333 (O_1333,N_18360,N_18557);
xnor UO_1334 (O_1334,N_18276,N_18967);
and UO_1335 (O_1335,N_19772,N_18050);
and UO_1336 (O_1336,N_18895,N_18072);
nand UO_1337 (O_1337,N_18481,N_18150);
nor UO_1338 (O_1338,N_19181,N_19917);
nand UO_1339 (O_1339,N_18924,N_19568);
or UO_1340 (O_1340,N_19385,N_18986);
or UO_1341 (O_1341,N_18338,N_19924);
or UO_1342 (O_1342,N_19530,N_19873);
nor UO_1343 (O_1343,N_18428,N_18889);
nand UO_1344 (O_1344,N_19846,N_19099);
or UO_1345 (O_1345,N_18357,N_19057);
and UO_1346 (O_1346,N_18412,N_18351);
nor UO_1347 (O_1347,N_18434,N_18305);
nand UO_1348 (O_1348,N_18849,N_19797);
nand UO_1349 (O_1349,N_19044,N_18374);
xnor UO_1350 (O_1350,N_18391,N_18321);
nand UO_1351 (O_1351,N_18308,N_19204);
or UO_1352 (O_1352,N_19850,N_18716);
or UO_1353 (O_1353,N_18799,N_19521);
and UO_1354 (O_1354,N_19905,N_18192);
nand UO_1355 (O_1355,N_18776,N_18839);
xnor UO_1356 (O_1356,N_19154,N_19061);
or UO_1357 (O_1357,N_18309,N_19048);
and UO_1358 (O_1358,N_18448,N_19586);
or UO_1359 (O_1359,N_19394,N_18591);
xnor UO_1360 (O_1360,N_18700,N_18876);
or UO_1361 (O_1361,N_18810,N_18997);
or UO_1362 (O_1362,N_18826,N_18654);
nand UO_1363 (O_1363,N_18042,N_19080);
xor UO_1364 (O_1364,N_19466,N_19182);
nand UO_1365 (O_1365,N_19337,N_18044);
or UO_1366 (O_1366,N_18037,N_18777);
nand UO_1367 (O_1367,N_19542,N_19302);
nor UO_1368 (O_1368,N_18686,N_19131);
nand UO_1369 (O_1369,N_18603,N_19904);
or UO_1370 (O_1370,N_18595,N_19205);
xnor UO_1371 (O_1371,N_19190,N_18681);
xnor UO_1372 (O_1372,N_18235,N_18358);
xor UO_1373 (O_1373,N_19273,N_19077);
and UO_1374 (O_1374,N_18926,N_18162);
nor UO_1375 (O_1375,N_19866,N_18857);
nand UO_1376 (O_1376,N_19563,N_19455);
or UO_1377 (O_1377,N_18014,N_18663);
nand UO_1378 (O_1378,N_19767,N_18607);
and UO_1379 (O_1379,N_19128,N_19015);
and UO_1380 (O_1380,N_19242,N_19590);
or UO_1381 (O_1381,N_18402,N_19143);
or UO_1382 (O_1382,N_18378,N_18911);
nor UO_1383 (O_1383,N_19381,N_18032);
nor UO_1384 (O_1384,N_19577,N_18747);
xor UO_1385 (O_1385,N_19203,N_19003);
and UO_1386 (O_1386,N_18478,N_19371);
nor UO_1387 (O_1387,N_18603,N_18019);
nor UO_1388 (O_1388,N_19022,N_19717);
nand UO_1389 (O_1389,N_18993,N_19542);
and UO_1390 (O_1390,N_19964,N_19911);
and UO_1391 (O_1391,N_19120,N_19746);
or UO_1392 (O_1392,N_19897,N_18865);
or UO_1393 (O_1393,N_18300,N_18836);
or UO_1394 (O_1394,N_18581,N_18288);
nand UO_1395 (O_1395,N_19312,N_19811);
and UO_1396 (O_1396,N_19750,N_19888);
nand UO_1397 (O_1397,N_18900,N_18316);
or UO_1398 (O_1398,N_18874,N_19730);
xor UO_1399 (O_1399,N_18711,N_18131);
or UO_1400 (O_1400,N_19065,N_18483);
and UO_1401 (O_1401,N_19599,N_19003);
nand UO_1402 (O_1402,N_19279,N_19514);
nor UO_1403 (O_1403,N_19653,N_18282);
xor UO_1404 (O_1404,N_18218,N_18502);
nor UO_1405 (O_1405,N_19590,N_18864);
nand UO_1406 (O_1406,N_19999,N_18845);
nor UO_1407 (O_1407,N_18615,N_18782);
nand UO_1408 (O_1408,N_19622,N_19760);
or UO_1409 (O_1409,N_19488,N_19889);
or UO_1410 (O_1410,N_18832,N_18881);
nor UO_1411 (O_1411,N_18255,N_18649);
nand UO_1412 (O_1412,N_19856,N_18945);
nor UO_1413 (O_1413,N_18600,N_18297);
nand UO_1414 (O_1414,N_18490,N_18765);
or UO_1415 (O_1415,N_18001,N_18392);
or UO_1416 (O_1416,N_19691,N_18366);
and UO_1417 (O_1417,N_19024,N_18158);
nor UO_1418 (O_1418,N_18859,N_19931);
xnor UO_1419 (O_1419,N_19886,N_18690);
nand UO_1420 (O_1420,N_18528,N_18080);
and UO_1421 (O_1421,N_19179,N_19669);
nand UO_1422 (O_1422,N_19843,N_18514);
nand UO_1423 (O_1423,N_18566,N_18845);
nand UO_1424 (O_1424,N_19455,N_18890);
and UO_1425 (O_1425,N_19305,N_19396);
nand UO_1426 (O_1426,N_18342,N_19660);
nor UO_1427 (O_1427,N_19118,N_18792);
or UO_1428 (O_1428,N_19379,N_19489);
or UO_1429 (O_1429,N_18177,N_19515);
or UO_1430 (O_1430,N_18087,N_19971);
and UO_1431 (O_1431,N_19167,N_19375);
nor UO_1432 (O_1432,N_18589,N_19193);
nor UO_1433 (O_1433,N_18939,N_18978);
nand UO_1434 (O_1434,N_19228,N_19580);
or UO_1435 (O_1435,N_18105,N_18611);
nor UO_1436 (O_1436,N_18457,N_18567);
nor UO_1437 (O_1437,N_19052,N_18062);
nor UO_1438 (O_1438,N_19436,N_19587);
nand UO_1439 (O_1439,N_18023,N_18059);
or UO_1440 (O_1440,N_19071,N_19193);
and UO_1441 (O_1441,N_18929,N_19034);
and UO_1442 (O_1442,N_19441,N_18200);
and UO_1443 (O_1443,N_19835,N_19734);
and UO_1444 (O_1444,N_19554,N_18258);
and UO_1445 (O_1445,N_18286,N_19195);
nor UO_1446 (O_1446,N_18802,N_18258);
or UO_1447 (O_1447,N_18249,N_18337);
and UO_1448 (O_1448,N_19490,N_18037);
and UO_1449 (O_1449,N_19320,N_19083);
nor UO_1450 (O_1450,N_18972,N_19242);
or UO_1451 (O_1451,N_18464,N_18812);
and UO_1452 (O_1452,N_19828,N_18153);
nand UO_1453 (O_1453,N_19385,N_18139);
or UO_1454 (O_1454,N_19508,N_19490);
and UO_1455 (O_1455,N_19797,N_18357);
and UO_1456 (O_1456,N_18917,N_18164);
nand UO_1457 (O_1457,N_19350,N_19645);
xnor UO_1458 (O_1458,N_19396,N_18796);
nand UO_1459 (O_1459,N_19056,N_18048);
nor UO_1460 (O_1460,N_18936,N_18615);
or UO_1461 (O_1461,N_19299,N_18514);
and UO_1462 (O_1462,N_19569,N_19529);
nand UO_1463 (O_1463,N_19764,N_18111);
nand UO_1464 (O_1464,N_18810,N_19861);
and UO_1465 (O_1465,N_19901,N_19158);
xor UO_1466 (O_1466,N_19046,N_18792);
nor UO_1467 (O_1467,N_18716,N_18207);
nor UO_1468 (O_1468,N_18919,N_19342);
and UO_1469 (O_1469,N_18901,N_18198);
and UO_1470 (O_1470,N_19346,N_18397);
nand UO_1471 (O_1471,N_18103,N_19400);
nand UO_1472 (O_1472,N_19434,N_18787);
and UO_1473 (O_1473,N_19883,N_19084);
nand UO_1474 (O_1474,N_19930,N_19393);
or UO_1475 (O_1475,N_19251,N_19405);
nand UO_1476 (O_1476,N_19261,N_18947);
nand UO_1477 (O_1477,N_19537,N_18062);
and UO_1478 (O_1478,N_18006,N_18662);
and UO_1479 (O_1479,N_19084,N_18565);
and UO_1480 (O_1480,N_18065,N_18305);
xnor UO_1481 (O_1481,N_19429,N_18681);
nor UO_1482 (O_1482,N_19706,N_19962);
nand UO_1483 (O_1483,N_18547,N_18140);
nand UO_1484 (O_1484,N_18078,N_19069);
and UO_1485 (O_1485,N_18563,N_19209);
nor UO_1486 (O_1486,N_19110,N_19544);
nor UO_1487 (O_1487,N_18211,N_19970);
xor UO_1488 (O_1488,N_19989,N_19530);
and UO_1489 (O_1489,N_19814,N_18575);
or UO_1490 (O_1490,N_18547,N_19337);
nor UO_1491 (O_1491,N_18483,N_19400);
nor UO_1492 (O_1492,N_18716,N_19639);
nand UO_1493 (O_1493,N_19335,N_18151);
or UO_1494 (O_1494,N_18938,N_19696);
nor UO_1495 (O_1495,N_18484,N_18611);
nand UO_1496 (O_1496,N_19208,N_18107);
and UO_1497 (O_1497,N_19344,N_19893);
xnor UO_1498 (O_1498,N_18749,N_19633);
and UO_1499 (O_1499,N_18079,N_19093);
and UO_1500 (O_1500,N_18760,N_18361);
and UO_1501 (O_1501,N_18362,N_19674);
or UO_1502 (O_1502,N_18286,N_19690);
or UO_1503 (O_1503,N_18418,N_18742);
nand UO_1504 (O_1504,N_19104,N_19312);
xor UO_1505 (O_1505,N_19408,N_19270);
or UO_1506 (O_1506,N_18991,N_18078);
nor UO_1507 (O_1507,N_19754,N_19044);
and UO_1508 (O_1508,N_19129,N_18282);
nand UO_1509 (O_1509,N_19420,N_19043);
nand UO_1510 (O_1510,N_18736,N_18696);
nor UO_1511 (O_1511,N_18690,N_19073);
and UO_1512 (O_1512,N_19783,N_19241);
nor UO_1513 (O_1513,N_19173,N_19567);
and UO_1514 (O_1514,N_18760,N_19272);
or UO_1515 (O_1515,N_19718,N_18357);
nand UO_1516 (O_1516,N_18625,N_19682);
xnor UO_1517 (O_1517,N_19025,N_19227);
and UO_1518 (O_1518,N_19178,N_18695);
or UO_1519 (O_1519,N_19937,N_18059);
or UO_1520 (O_1520,N_18019,N_18378);
or UO_1521 (O_1521,N_18094,N_19954);
or UO_1522 (O_1522,N_19871,N_18060);
nand UO_1523 (O_1523,N_18070,N_18768);
nand UO_1524 (O_1524,N_19858,N_19813);
and UO_1525 (O_1525,N_18477,N_18189);
nor UO_1526 (O_1526,N_19773,N_19890);
and UO_1527 (O_1527,N_18660,N_19905);
nor UO_1528 (O_1528,N_18728,N_19712);
nand UO_1529 (O_1529,N_19065,N_18817);
and UO_1530 (O_1530,N_19467,N_18051);
nand UO_1531 (O_1531,N_18075,N_18538);
nor UO_1532 (O_1532,N_18655,N_19044);
and UO_1533 (O_1533,N_18670,N_19583);
or UO_1534 (O_1534,N_19584,N_18925);
xnor UO_1535 (O_1535,N_19776,N_19852);
nor UO_1536 (O_1536,N_18897,N_18238);
or UO_1537 (O_1537,N_18549,N_19531);
and UO_1538 (O_1538,N_18244,N_18564);
nand UO_1539 (O_1539,N_18919,N_19346);
nand UO_1540 (O_1540,N_18655,N_19383);
and UO_1541 (O_1541,N_18772,N_19415);
nor UO_1542 (O_1542,N_18077,N_18352);
nor UO_1543 (O_1543,N_19233,N_18006);
or UO_1544 (O_1544,N_18347,N_18767);
xor UO_1545 (O_1545,N_18430,N_19818);
or UO_1546 (O_1546,N_18514,N_18144);
or UO_1547 (O_1547,N_19619,N_19969);
nand UO_1548 (O_1548,N_19582,N_19080);
and UO_1549 (O_1549,N_19073,N_19761);
nand UO_1550 (O_1550,N_19655,N_18749);
nor UO_1551 (O_1551,N_18495,N_18398);
and UO_1552 (O_1552,N_19910,N_19451);
or UO_1553 (O_1553,N_19319,N_18498);
nor UO_1554 (O_1554,N_19261,N_19723);
nor UO_1555 (O_1555,N_18660,N_19537);
and UO_1556 (O_1556,N_19418,N_19669);
nor UO_1557 (O_1557,N_19782,N_19116);
or UO_1558 (O_1558,N_19867,N_19246);
and UO_1559 (O_1559,N_19074,N_19304);
and UO_1560 (O_1560,N_18412,N_19072);
and UO_1561 (O_1561,N_19851,N_18185);
and UO_1562 (O_1562,N_18241,N_18744);
nor UO_1563 (O_1563,N_19006,N_18951);
and UO_1564 (O_1564,N_18871,N_18171);
and UO_1565 (O_1565,N_18078,N_18821);
nor UO_1566 (O_1566,N_18855,N_18524);
xor UO_1567 (O_1567,N_18861,N_19420);
nand UO_1568 (O_1568,N_18689,N_18313);
and UO_1569 (O_1569,N_19413,N_19196);
and UO_1570 (O_1570,N_19455,N_18779);
and UO_1571 (O_1571,N_18164,N_19511);
nor UO_1572 (O_1572,N_19021,N_19602);
or UO_1573 (O_1573,N_19311,N_19914);
or UO_1574 (O_1574,N_18994,N_19012);
or UO_1575 (O_1575,N_19165,N_18505);
or UO_1576 (O_1576,N_19467,N_19072);
or UO_1577 (O_1577,N_19323,N_18303);
and UO_1578 (O_1578,N_19959,N_19595);
nand UO_1579 (O_1579,N_18369,N_18098);
nor UO_1580 (O_1580,N_19817,N_19583);
and UO_1581 (O_1581,N_19926,N_18757);
xnor UO_1582 (O_1582,N_18678,N_19533);
nand UO_1583 (O_1583,N_19655,N_19890);
xor UO_1584 (O_1584,N_19515,N_18282);
nand UO_1585 (O_1585,N_19212,N_19793);
and UO_1586 (O_1586,N_19577,N_18052);
or UO_1587 (O_1587,N_18391,N_18809);
or UO_1588 (O_1588,N_18919,N_18748);
nand UO_1589 (O_1589,N_18799,N_18118);
nor UO_1590 (O_1590,N_19180,N_19574);
and UO_1591 (O_1591,N_19069,N_18434);
nor UO_1592 (O_1592,N_18600,N_18830);
and UO_1593 (O_1593,N_18092,N_18677);
nor UO_1594 (O_1594,N_18740,N_19891);
xor UO_1595 (O_1595,N_19117,N_19291);
nand UO_1596 (O_1596,N_18814,N_18408);
nand UO_1597 (O_1597,N_19501,N_18543);
or UO_1598 (O_1598,N_18082,N_18184);
or UO_1599 (O_1599,N_19464,N_18013);
nand UO_1600 (O_1600,N_19945,N_18182);
and UO_1601 (O_1601,N_19448,N_19058);
nand UO_1602 (O_1602,N_18278,N_19578);
nand UO_1603 (O_1603,N_18078,N_18209);
nor UO_1604 (O_1604,N_19047,N_18855);
or UO_1605 (O_1605,N_18206,N_18714);
nor UO_1606 (O_1606,N_19426,N_19904);
and UO_1607 (O_1607,N_19873,N_18331);
and UO_1608 (O_1608,N_18014,N_18167);
or UO_1609 (O_1609,N_18416,N_18614);
nor UO_1610 (O_1610,N_18839,N_19937);
and UO_1611 (O_1611,N_19130,N_19756);
xor UO_1612 (O_1612,N_18889,N_18527);
and UO_1613 (O_1613,N_19000,N_18946);
xnor UO_1614 (O_1614,N_18590,N_19379);
xnor UO_1615 (O_1615,N_18933,N_19759);
or UO_1616 (O_1616,N_19989,N_19504);
nand UO_1617 (O_1617,N_19871,N_19417);
nor UO_1618 (O_1618,N_19710,N_18094);
and UO_1619 (O_1619,N_18730,N_19596);
or UO_1620 (O_1620,N_18762,N_18185);
xor UO_1621 (O_1621,N_19666,N_18673);
nor UO_1622 (O_1622,N_19108,N_18998);
or UO_1623 (O_1623,N_19701,N_18731);
nand UO_1624 (O_1624,N_19204,N_18566);
or UO_1625 (O_1625,N_19311,N_18158);
nand UO_1626 (O_1626,N_19041,N_18494);
nor UO_1627 (O_1627,N_19875,N_19599);
or UO_1628 (O_1628,N_19304,N_19284);
nand UO_1629 (O_1629,N_19144,N_18349);
nand UO_1630 (O_1630,N_18997,N_18192);
nand UO_1631 (O_1631,N_19505,N_19061);
nand UO_1632 (O_1632,N_19239,N_18484);
and UO_1633 (O_1633,N_19350,N_19322);
or UO_1634 (O_1634,N_19062,N_19173);
or UO_1635 (O_1635,N_19883,N_19128);
nand UO_1636 (O_1636,N_18767,N_18065);
and UO_1637 (O_1637,N_18382,N_18055);
and UO_1638 (O_1638,N_18518,N_18393);
nand UO_1639 (O_1639,N_19830,N_18527);
or UO_1640 (O_1640,N_18590,N_19983);
nor UO_1641 (O_1641,N_18521,N_19204);
nor UO_1642 (O_1642,N_18655,N_18706);
or UO_1643 (O_1643,N_19568,N_19956);
nor UO_1644 (O_1644,N_18846,N_18582);
or UO_1645 (O_1645,N_18912,N_18610);
nor UO_1646 (O_1646,N_18872,N_18023);
or UO_1647 (O_1647,N_19760,N_19324);
or UO_1648 (O_1648,N_18906,N_18130);
nand UO_1649 (O_1649,N_19344,N_18118);
and UO_1650 (O_1650,N_18018,N_18241);
and UO_1651 (O_1651,N_18867,N_18522);
nor UO_1652 (O_1652,N_18982,N_18131);
and UO_1653 (O_1653,N_19198,N_19694);
and UO_1654 (O_1654,N_19620,N_18724);
nand UO_1655 (O_1655,N_19247,N_18234);
nor UO_1656 (O_1656,N_18863,N_19564);
nor UO_1657 (O_1657,N_18100,N_19623);
or UO_1658 (O_1658,N_19595,N_18767);
nor UO_1659 (O_1659,N_19102,N_18751);
or UO_1660 (O_1660,N_18783,N_19247);
and UO_1661 (O_1661,N_19297,N_18362);
nor UO_1662 (O_1662,N_19956,N_19139);
nor UO_1663 (O_1663,N_19785,N_19360);
nand UO_1664 (O_1664,N_18208,N_19487);
nor UO_1665 (O_1665,N_19212,N_19794);
nor UO_1666 (O_1666,N_19476,N_18251);
xnor UO_1667 (O_1667,N_18426,N_18610);
xor UO_1668 (O_1668,N_18639,N_19322);
nand UO_1669 (O_1669,N_18993,N_19406);
or UO_1670 (O_1670,N_18181,N_18045);
and UO_1671 (O_1671,N_18453,N_18316);
nand UO_1672 (O_1672,N_19415,N_19866);
nor UO_1673 (O_1673,N_18535,N_18594);
nand UO_1674 (O_1674,N_18490,N_19839);
nor UO_1675 (O_1675,N_18998,N_18521);
and UO_1676 (O_1676,N_19587,N_19889);
nand UO_1677 (O_1677,N_19278,N_18308);
xnor UO_1678 (O_1678,N_18389,N_19281);
nor UO_1679 (O_1679,N_19361,N_19487);
or UO_1680 (O_1680,N_18757,N_19366);
and UO_1681 (O_1681,N_18295,N_18261);
or UO_1682 (O_1682,N_18218,N_19054);
xor UO_1683 (O_1683,N_19384,N_19670);
and UO_1684 (O_1684,N_18402,N_18337);
or UO_1685 (O_1685,N_19269,N_19777);
and UO_1686 (O_1686,N_18791,N_18820);
and UO_1687 (O_1687,N_18202,N_19504);
nand UO_1688 (O_1688,N_18241,N_19862);
nand UO_1689 (O_1689,N_19305,N_19999);
nor UO_1690 (O_1690,N_19671,N_18163);
and UO_1691 (O_1691,N_18328,N_18940);
nand UO_1692 (O_1692,N_19969,N_18062);
and UO_1693 (O_1693,N_19088,N_19884);
nor UO_1694 (O_1694,N_18851,N_18275);
xor UO_1695 (O_1695,N_19575,N_18677);
nand UO_1696 (O_1696,N_19599,N_19225);
nand UO_1697 (O_1697,N_19195,N_19327);
and UO_1698 (O_1698,N_19689,N_19932);
and UO_1699 (O_1699,N_19807,N_19733);
nand UO_1700 (O_1700,N_18092,N_18213);
or UO_1701 (O_1701,N_19991,N_18740);
nor UO_1702 (O_1702,N_19199,N_18697);
and UO_1703 (O_1703,N_18169,N_19456);
nor UO_1704 (O_1704,N_19962,N_19854);
and UO_1705 (O_1705,N_19878,N_19627);
and UO_1706 (O_1706,N_19205,N_18363);
and UO_1707 (O_1707,N_18245,N_19634);
or UO_1708 (O_1708,N_19427,N_19797);
or UO_1709 (O_1709,N_18074,N_19306);
nor UO_1710 (O_1710,N_18892,N_18336);
nor UO_1711 (O_1711,N_19800,N_18303);
nor UO_1712 (O_1712,N_18333,N_18330);
nand UO_1713 (O_1713,N_19288,N_19276);
nor UO_1714 (O_1714,N_18518,N_18733);
nor UO_1715 (O_1715,N_19930,N_18435);
nor UO_1716 (O_1716,N_18042,N_19298);
nor UO_1717 (O_1717,N_19546,N_18979);
nand UO_1718 (O_1718,N_19211,N_19212);
and UO_1719 (O_1719,N_18669,N_19290);
or UO_1720 (O_1720,N_18578,N_18966);
nand UO_1721 (O_1721,N_19819,N_18365);
nor UO_1722 (O_1722,N_18057,N_18383);
or UO_1723 (O_1723,N_19833,N_19449);
nor UO_1724 (O_1724,N_18084,N_18809);
nand UO_1725 (O_1725,N_19214,N_19180);
or UO_1726 (O_1726,N_18474,N_18432);
or UO_1727 (O_1727,N_19370,N_19345);
nand UO_1728 (O_1728,N_18160,N_18328);
and UO_1729 (O_1729,N_18319,N_18860);
nor UO_1730 (O_1730,N_18917,N_19956);
nand UO_1731 (O_1731,N_19583,N_19675);
nor UO_1732 (O_1732,N_19711,N_19064);
nor UO_1733 (O_1733,N_18079,N_18220);
or UO_1734 (O_1734,N_18080,N_18217);
and UO_1735 (O_1735,N_18429,N_19632);
and UO_1736 (O_1736,N_18672,N_18893);
or UO_1737 (O_1737,N_19172,N_19760);
or UO_1738 (O_1738,N_19813,N_19034);
nand UO_1739 (O_1739,N_18095,N_18657);
or UO_1740 (O_1740,N_19048,N_19125);
and UO_1741 (O_1741,N_19649,N_19299);
xnor UO_1742 (O_1742,N_19156,N_18796);
and UO_1743 (O_1743,N_18624,N_18912);
nand UO_1744 (O_1744,N_18818,N_19717);
nand UO_1745 (O_1745,N_19607,N_19200);
or UO_1746 (O_1746,N_19451,N_19767);
xor UO_1747 (O_1747,N_19136,N_18199);
or UO_1748 (O_1748,N_19656,N_19831);
nor UO_1749 (O_1749,N_19844,N_19946);
or UO_1750 (O_1750,N_19582,N_19464);
xor UO_1751 (O_1751,N_18444,N_18640);
and UO_1752 (O_1752,N_18236,N_19386);
nor UO_1753 (O_1753,N_19279,N_19786);
and UO_1754 (O_1754,N_18790,N_18025);
xor UO_1755 (O_1755,N_19626,N_19637);
or UO_1756 (O_1756,N_19178,N_18078);
nand UO_1757 (O_1757,N_19755,N_18628);
nor UO_1758 (O_1758,N_18635,N_19054);
or UO_1759 (O_1759,N_18416,N_18045);
and UO_1760 (O_1760,N_19806,N_18339);
or UO_1761 (O_1761,N_18635,N_18755);
or UO_1762 (O_1762,N_18097,N_19624);
xnor UO_1763 (O_1763,N_18897,N_18315);
nand UO_1764 (O_1764,N_18094,N_18389);
or UO_1765 (O_1765,N_18767,N_18440);
nand UO_1766 (O_1766,N_19126,N_18262);
nor UO_1767 (O_1767,N_18894,N_19111);
and UO_1768 (O_1768,N_19610,N_18747);
or UO_1769 (O_1769,N_19902,N_19422);
or UO_1770 (O_1770,N_19833,N_18834);
xor UO_1771 (O_1771,N_19355,N_19734);
or UO_1772 (O_1772,N_19920,N_18211);
and UO_1773 (O_1773,N_19936,N_18938);
and UO_1774 (O_1774,N_19925,N_19433);
or UO_1775 (O_1775,N_18963,N_19776);
xor UO_1776 (O_1776,N_18848,N_19449);
nor UO_1777 (O_1777,N_18571,N_19054);
and UO_1778 (O_1778,N_19716,N_19990);
nand UO_1779 (O_1779,N_19943,N_19254);
xnor UO_1780 (O_1780,N_19046,N_19079);
or UO_1781 (O_1781,N_19525,N_18201);
nand UO_1782 (O_1782,N_19813,N_18574);
xnor UO_1783 (O_1783,N_19825,N_19248);
nand UO_1784 (O_1784,N_18499,N_19232);
nand UO_1785 (O_1785,N_19813,N_19426);
nand UO_1786 (O_1786,N_18593,N_18316);
and UO_1787 (O_1787,N_18819,N_19290);
or UO_1788 (O_1788,N_19930,N_19450);
and UO_1789 (O_1789,N_19043,N_19630);
nand UO_1790 (O_1790,N_18822,N_19216);
nand UO_1791 (O_1791,N_18034,N_18731);
nand UO_1792 (O_1792,N_19919,N_18425);
or UO_1793 (O_1793,N_19419,N_18772);
and UO_1794 (O_1794,N_19442,N_18464);
nor UO_1795 (O_1795,N_19302,N_19507);
or UO_1796 (O_1796,N_18617,N_19568);
nor UO_1797 (O_1797,N_18904,N_18136);
or UO_1798 (O_1798,N_19395,N_19073);
xor UO_1799 (O_1799,N_19441,N_19380);
nand UO_1800 (O_1800,N_19055,N_18385);
and UO_1801 (O_1801,N_18044,N_18602);
and UO_1802 (O_1802,N_18378,N_19011);
nor UO_1803 (O_1803,N_18685,N_18100);
xnor UO_1804 (O_1804,N_18485,N_19444);
nand UO_1805 (O_1805,N_18360,N_18738);
or UO_1806 (O_1806,N_18405,N_18851);
nor UO_1807 (O_1807,N_18608,N_19645);
or UO_1808 (O_1808,N_18651,N_19458);
nand UO_1809 (O_1809,N_18231,N_19320);
and UO_1810 (O_1810,N_18457,N_18637);
or UO_1811 (O_1811,N_18191,N_18950);
nor UO_1812 (O_1812,N_19831,N_18942);
nor UO_1813 (O_1813,N_19338,N_18012);
nor UO_1814 (O_1814,N_18083,N_19512);
nor UO_1815 (O_1815,N_19901,N_19511);
nand UO_1816 (O_1816,N_19723,N_19206);
and UO_1817 (O_1817,N_18873,N_19988);
and UO_1818 (O_1818,N_18015,N_18488);
or UO_1819 (O_1819,N_18234,N_19486);
or UO_1820 (O_1820,N_18429,N_18372);
or UO_1821 (O_1821,N_19365,N_18192);
or UO_1822 (O_1822,N_19460,N_19334);
nand UO_1823 (O_1823,N_18406,N_18543);
nor UO_1824 (O_1824,N_18181,N_18273);
nand UO_1825 (O_1825,N_19585,N_18318);
nand UO_1826 (O_1826,N_18027,N_19824);
and UO_1827 (O_1827,N_18225,N_19788);
nand UO_1828 (O_1828,N_19013,N_19793);
nor UO_1829 (O_1829,N_18293,N_18322);
or UO_1830 (O_1830,N_19147,N_19201);
nand UO_1831 (O_1831,N_19757,N_19994);
nand UO_1832 (O_1832,N_18980,N_19804);
or UO_1833 (O_1833,N_19218,N_19463);
and UO_1834 (O_1834,N_18368,N_19107);
and UO_1835 (O_1835,N_19375,N_18561);
nand UO_1836 (O_1836,N_18569,N_19823);
or UO_1837 (O_1837,N_18760,N_19594);
and UO_1838 (O_1838,N_18852,N_18050);
and UO_1839 (O_1839,N_18451,N_18589);
and UO_1840 (O_1840,N_19237,N_18279);
and UO_1841 (O_1841,N_19712,N_19419);
nor UO_1842 (O_1842,N_18967,N_19350);
nor UO_1843 (O_1843,N_19122,N_18632);
or UO_1844 (O_1844,N_19676,N_19992);
or UO_1845 (O_1845,N_19554,N_18001);
and UO_1846 (O_1846,N_19881,N_18164);
nor UO_1847 (O_1847,N_19958,N_18592);
nor UO_1848 (O_1848,N_18427,N_19360);
xor UO_1849 (O_1849,N_19017,N_19347);
nor UO_1850 (O_1850,N_18042,N_18949);
or UO_1851 (O_1851,N_19079,N_19778);
or UO_1852 (O_1852,N_18385,N_19642);
nand UO_1853 (O_1853,N_19343,N_19865);
or UO_1854 (O_1854,N_18665,N_18675);
and UO_1855 (O_1855,N_19563,N_18259);
nand UO_1856 (O_1856,N_19880,N_18944);
or UO_1857 (O_1857,N_19666,N_18897);
and UO_1858 (O_1858,N_18629,N_18757);
or UO_1859 (O_1859,N_18755,N_18357);
xor UO_1860 (O_1860,N_18226,N_19919);
xor UO_1861 (O_1861,N_18224,N_19326);
or UO_1862 (O_1862,N_18087,N_18553);
nand UO_1863 (O_1863,N_19969,N_18097);
nor UO_1864 (O_1864,N_18093,N_19828);
nor UO_1865 (O_1865,N_19722,N_19839);
nor UO_1866 (O_1866,N_19769,N_19462);
nand UO_1867 (O_1867,N_18536,N_19135);
or UO_1868 (O_1868,N_19747,N_18119);
nand UO_1869 (O_1869,N_19687,N_19218);
or UO_1870 (O_1870,N_19962,N_18174);
nor UO_1871 (O_1871,N_19169,N_19303);
and UO_1872 (O_1872,N_19789,N_19503);
nor UO_1873 (O_1873,N_19655,N_19130);
nor UO_1874 (O_1874,N_18609,N_18598);
or UO_1875 (O_1875,N_18124,N_19769);
nand UO_1876 (O_1876,N_18522,N_19179);
xor UO_1877 (O_1877,N_18319,N_18649);
and UO_1878 (O_1878,N_19290,N_19340);
and UO_1879 (O_1879,N_19785,N_18750);
xnor UO_1880 (O_1880,N_18785,N_19853);
nor UO_1881 (O_1881,N_18621,N_19324);
and UO_1882 (O_1882,N_19837,N_18674);
nand UO_1883 (O_1883,N_18555,N_19401);
and UO_1884 (O_1884,N_18518,N_19292);
or UO_1885 (O_1885,N_19428,N_19899);
and UO_1886 (O_1886,N_19388,N_19259);
or UO_1887 (O_1887,N_19742,N_19170);
nor UO_1888 (O_1888,N_18516,N_19120);
nor UO_1889 (O_1889,N_19056,N_18547);
nand UO_1890 (O_1890,N_18322,N_19255);
nand UO_1891 (O_1891,N_19942,N_18882);
or UO_1892 (O_1892,N_18673,N_19817);
nand UO_1893 (O_1893,N_19861,N_18233);
nand UO_1894 (O_1894,N_18081,N_19738);
and UO_1895 (O_1895,N_19456,N_18174);
nor UO_1896 (O_1896,N_19324,N_19671);
nand UO_1897 (O_1897,N_19619,N_19565);
and UO_1898 (O_1898,N_18805,N_19581);
and UO_1899 (O_1899,N_19682,N_18186);
nand UO_1900 (O_1900,N_19958,N_18338);
and UO_1901 (O_1901,N_18760,N_18092);
nand UO_1902 (O_1902,N_18252,N_18163);
nand UO_1903 (O_1903,N_18891,N_18501);
and UO_1904 (O_1904,N_19586,N_19479);
and UO_1905 (O_1905,N_19048,N_18339);
or UO_1906 (O_1906,N_18203,N_19214);
xnor UO_1907 (O_1907,N_18779,N_18142);
nor UO_1908 (O_1908,N_19647,N_18061);
and UO_1909 (O_1909,N_19107,N_18997);
xor UO_1910 (O_1910,N_18764,N_18136);
nand UO_1911 (O_1911,N_18970,N_18160);
nor UO_1912 (O_1912,N_19454,N_19558);
or UO_1913 (O_1913,N_18164,N_19324);
nand UO_1914 (O_1914,N_18357,N_18985);
nand UO_1915 (O_1915,N_19445,N_18577);
nor UO_1916 (O_1916,N_18400,N_18190);
nand UO_1917 (O_1917,N_19942,N_19630);
or UO_1918 (O_1918,N_18662,N_19171);
nand UO_1919 (O_1919,N_19553,N_18899);
nand UO_1920 (O_1920,N_18019,N_18204);
nand UO_1921 (O_1921,N_19174,N_19085);
xnor UO_1922 (O_1922,N_18503,N_19008);
or UO_1923 (O_1923,N_18089,N_18913);
nand UO_1924 (O_1924,N_18737,N_19531);
and UO_1925 (O_1925,N_18110,N_18384);
nand UO_1926 (O_1926,N_18462,N_18977);
or UO_1927 (O_1927,N_19678,N_19816);
or UO_1928 (O_1928,N_18129,N_19346);
nand UO_1929 (O_1929,N_18346,N_19528);
xor UO_1930 (O_1930,N_18700,N_18500);
nand UO_1931 (O_1931,N_18868,N_19627);
nand UO_1932 (O_1932,N_19652,N_18045);
or UO_1933 (O_1933,N_19856,N_19311);
nor UO_1934 (O_1934,N_19898,N_18925);
xor UO_1935 (O_1935,N_19743,N_19539);
and UO_1936 (O_1936,N_19074,N_18474);
xnor UO_1937 (O_1937,N_19361,N_18359);
or UO_1938 (O_1938,N_19104,N_18222);
nand UO_1939 (O_1939,N_19617,N_18402);
or UO_1940 (O_1940,N_19982,N_18166);
nor UO_1941 (O_1941,N_19167,N_18070);
xnor UO_1942 (O_1942,N_19889,N_19009);
or UO_1943 (O_1943,N_18199,N_18084);
and UO_1944 (O_1944,N_19096,N_18215);
nand UO_1945 (O_1945,N_18429,N_19153);
and UO_1946 (O_1946,N_18471,N_18790);
xor UO_1947 (O_1947,N_18383,N_18775);
nand UO_1948 (O_1948,N_19940,N_18697);
and UO_1949 (O_1949,N_19184,N_19094);
nand UO_1950 (O_1950,N_18536,N_19118);
nor UO_1951 (O_1951,N_18989,N_18494);
and UO_1952 (O_1952,N_18161,N_18945);
nor UO_1953 (O_1953,N_19683,N_18908);
nor UO_1954 (O_1954,N_18931,N_18921);
nand UO_1955 (O_1955,N_18357,N_18084);
nor UO_1956 (O_1956,N_18017,N_19303);
nor UO_1957 (O_1957,N_19669,N_19211);
or UO_1958 (O_1958,N_18019,N_18566);
or UO_1959 (O_1959,N_19639,N_19269);
nand UO_1960 (O_1960,N_19661,N_19736);
and UO_1961 (O_1961,N_19108,N_18254);
nor UO_1962 (O_1962,N_19142,N_18059);
or UO_1963 (O_1963,N_19630,N_18679);
or UO_1964 (O_1964,N_19020,N_19604);
nor UO_1965 (O_1965,N_18919,N_18199);
and UO_1966 (O_1966,N_18676,N_18278);
nor UO_1967 (O_1967,N_19665,N_18699);
xnor UO_1968 (O_1968,N_19968,N_18902);
nand UO_1969 (O_1969,N_19457,N_19409);
or UO_1970 (O_1970,N_18106,N_18539);
nor UO_1971 (O_1971,N_18145,N_19056);
nor UO_1972 (O_1972,N_19364,N_19959);
nand UO_1973 (O_1973,N_19673,N_18405);
nor UO_1974 (O_1974,N_19614,N_18577);
nor UO_1975 (O_1975,N_19387,N_18735);
nor UO_1976 (O_1976,N_19065,N_19895);
or UO_1977 (O_1977,N_18903,N_19769);
and UO_1978 (O_1978,N_18754,N_18580);
nand UO_1979 (O_1979,N_19758,N_18260);
nor UO_1980 (O_1980,N_18169,N_18739);
nand UO_1981 (O_1981,N_19853,N_18436);
or UO_1982 (O_1982,N_19603,N_19311);
nand UO_1983 (O_1983,N_18072,N_18798);
or UO_1984 (O_1984,N_18491,N_18294);
or UO_1985 (O_1985,N_19356,N_19015);
nor UO_1986 (O_1986,N_19114,N_19010);
nand UO_1987 (O_1987,N_18512,N_19723);
and UO_1988 (O_1988,N_18151,N_19066);
nor UO_1989 (O_1989,N_19280,N_19293);
nand UO_1990 (O_1990,N_18629,N_18733);
or UO_1991 (O_1991,N_19007,N_18517);
and UO_1992 (O_1992,N_19809,N_18997);
or UO_1993 (O_1993,N_19562,N_18180);
nor UO_1994 (O_1994,N_19329,N_19465);
or UO_1995 (O_1995,N_19891,N_19520);
nor UO_1996 (O_1996,N_19521,N_18900);
and UO_1997 (O_1997,N_19021,N_18859);
or UO_1998 (O_1998,N_19998,N_18757);
nand UO_1999 (O_1999,N_18283,N_19133);
nor UO_2000 (O_2000,N_19333,N_19196);
nand UO_2001 (O_2001,N_19739,N_19618);
or UO_2002 (O_2002,N_18000,N_19364);
nand UO_2003 (O_2003,N_19749,N_19955);
nand UO_2004 (O_2004,N_19096,N_18877);
nor UO_2005 (O_2005,N_18083,N_18977);
or UO_2006 (O_2006,N_18053,N_19261);
nor UO_2007 (O_2007,N_18845,N_19910);
xor UO_2008 (O_2008,N_19238,N_18017);
or UO_2009 (O_2009,N_18176,N_19496);
xnor UO_2010 (O_2010,N_19787,N_19405);
or UO_2011 (O_2011,N_18097,N_19409);
or UO_2012 (O_2012,N_18400,N_19266);
and UO_2013 (O_2013,N_18412,N_18870);
and UO_2014 (O_2014,N_19418,N_18923);
xnor UO_2015 (O_2015,N_18519,N_18197);
and UO_2016 (O_2016,N_18670,N_18379);
nand UO_2017 (O_2017,N_19884,N_19749);
nor UO_2018 (O_2018,N_18656,N_19949);
nor UO_2019 (O_2019,N_19959,N_19511);
nand UO_2020 (O_2020,N_18981,N_18851);
nand UO_2021 (O_2021,N_19190,N_18340);
nand UO_2022 (O_2022,N_19501,N_19003);
xor UO_2023 (O_2023,N_19264,N_19266);
or UO_2024 (O_2024,N_19107,N_18339);
or UO_2025 (O_2025,N_18057,N_19644);
nor UO_2026 (O_2026,N_18499,N_18681);
nand UO_2027 (O_2027,N_19355,N_18742);
xnor UO_2028 (O_2028,N_19672,N_19784);
and UO_2029 (O_2029,N_19093,N_18692);
or UO_2030 (O_2030,N_18934,N_19616);
and UO_2031 (O_2031,N_18208,N_18672);
nor UO_2032 (O_2032,N_18266,N_19068);
and UO_2033 (O_2033,N_18435,N_19070);
nor UO_2034 (O_2034,N_19841,N_19034);
nor UO_2035 (O_2035,N_19928,N_18346);
and UO_2036 (O_2036,N_18438,N_19528);
and UO_2037 (O_2037,N_19930,N_19768);
nor UO_2038 (O_2038,N_19503,N_18334);
and UO_2039 (O_2039,N_19665,N_19087);
nor UO_2040 (O_2040,N_19367,N_18493);
and UO_2041 (O_2041,N_19375,N_18677);
or UO_2042 (O_2042,N_18498,N_19916);
nand UO_2043 (O_2043,N_19826,N_19918);
or UO_2044 (O_2044,N_19077,N_18010);
and UO_2045 (O_2045,N_19861,N_18641);
and UO_2046 (O_2046,N_18097,N_18881);
and UO_2047 (O_2047,N_18246,N_19814);
and UO_2048 (O_2048,N_18610,N_18419);
or UO_2049 (O_2049,N_18193,N_18204);
or UO_2050 (O_2050,N_18874,N_18315);
and UO_2051 (O_2051,N_18580,N_19285);
and UO_2052 (O_2052,N_18434,N_18368);
nand UO_2053 (O_2053,N_18219,N_19330);
or UO_2054 (O_2054,N_19813,N_19094);
xor UO_2055 (O_2055,N_18281,N_18181);
nand UO_2056 (O_2056,N_19574,N_18076);
xnor UO_2057 (O_2057,N_18789,N_18780);
nor UO_2058 (O_2058,N_19364,N_18508);
and UO_2059 (O_2059,N_18003,N_19806);
and UO_2060 (O_2060,N_18377,N_19969);
nor UO_2061 (O_2061,N_19651,N_18058);
or UO_2062 (O_2062,N_19791,N_19772);
or UO_2063 (O_2063,N_18950,N_19981);
nor UO_2064 (O_2064,N_18942,N_18787);
and UO_2065 (O_2065,N_18568,N_19541);
and UO_2066 (O_2066,N_18257,N_18404);
nand UO_2067 (O_2067,N_19783,N_19491);
and UO_2068 (O_2068,N_18018,N_18512);
and UO_2069 (O_2069,N_19056,N_19902);
or UO_2070 (O_2070,N_18529,N_19039);
and UO_2071 (O_2071,N_19063,N_19886);
nor UO_2072 (O_2072,N_18360,N_19079);
nand UO_2073 (O_2073,N_18000,N_18554);
nor UO_2074 (O_2074,N_19041,N_18652);
nand UO_2075 (O_2075,N_19029,N_18493);
or UO_2076 (O_2076,N_18911,N_18450);
nor UO_2077 (O_2077,N_19543,N_18419);
nor UO_2078 (O_2078,N_18804,N_19820);
or UO_2079 (O_2079,N_19911,N_18468);
nand UO_2080 (O_2080,N_19040,N_19337);
nand UO_2081 (O_2081,N_18602,N_18200);
nand UO_2082 (O_2082,N_18508,N_18457);
nand UO_2083 (O_2083,N_18278,N_18128);
or UO_2084 (O_2084,N_19648,N_18318);
xor UO_2085 (O_2085,N_18022,N_19353);
nor UO_2086 (O_2086,N_18458,N_18596);
nor UO_2087 (O_2087,N_19654,N_19407);
or UO_2088 (O_2088,N_18924,N_18039);
and UO_2089 (O_2089,N_18481,N_18711);
and UO_2090 (O_2090,N_18329,N_19838);
xnor UO_2091 (O_2091,N_18839,N_18709);
and UO_2092 (O_2092,N_18011,N_19725);
and UO_2093 (O_2093,N_18315,N_19367);
and UO_2094 (O_2094,N_18953,N_18437);
nor UO_2095 (O_2095,N_18556,N_18039);
or UO_2096 (O_2096,N_18049,N_19948);
and UO_2097 (O_2097,N_18209,N_18772);
nor UO_2098 (O_2098,N_19169,N_19517);
xor UO_2099 (O_2099,N_19638,N_19610);
nand UO_2100 (O_2100,N_19598,N_19614);
nor UO_2101 (O_2101,N_19865,N_18019);
or UO_2102 (O_2102,N_18388,N_19162);
and UO_2103 (O_2103,N_18477,N_18781);
or UO_2104 (O_2104,N_18070,N_18608);
and UO_2105 (O_2105,N_19796,N_18674);
nor UO_2106 (O_2106,N_19346,N_18577);
nand UO_2107 (O_2107,N_19378,N_18577);
and UO_2108 (O_2108,N_19994,N_19637);
nor UO_2109 (O_2109,N_18547,N_19867);
and UO_2110 (O_2110,N_18480,N_18023);
and UO_2111 (O_2111,N_19881,N_19361);
or UO_2112 (O_2112,N_19529,N_19329);
nor UO_2113 (O_2113,N_18489,N_18722);
and UO_2114 (O_2114,N_19965,N_19339);
nor UO_2115 (O_2115,N_18199,N_18128);
or UO_2116 (O_2116,N_19281,N_18332);
nand UO_2117 (O_2117,N_18744,N_19171);
nand UO_2118 (O_2118,N_18745,N_19249);
nor UO_2119 (O_2119,N_19881,N_18839);
nand UO_2120 (O_2120,N_19032,N_19292);
or UO_2121 (O_2121,N_19674,N_19317);
nor UO_2122 (O_2122,N_18671,N_19018);
nor UO_2123 (O_2123,N_18166,N_19784);
or UO_2124 (O_2124,N_18520,N_19255);
nand UO_2125 (O_2125,N_19734,N_19457);
nand UO_2126 (O_2126,N_18380,N_18838);
or UO_2127 (O_2127,N_19656,N_18635);
nand UO_2128 (O_2128,N_19990,N_18011);
nand UO_2129 (O_2129,N_18637,N_18079);
nand UO_2130 (O_2130,N_18044,N_19477);
xnor UO_2131 (O_2131,N_19258,N_19252);
and UO_2132 (O_2132,N_18615,N_19332);
nor UO_2133 (O_2133,N_19956,N_18450);
nand UO_2134 (O_2134,N_19760,N_19110);
nand UO_2135 (O_2135,N_19526,N_18564);
nor UO_2136 (O_2136,N_18568,N_18602);
or UO_2137 (O_2137,N_18376,N_18887);
nor UO_2138 (O_2138,N_18730,N_19793);
nor UO_2139 (O_2139,N_18439,N_19255);
nor UO_2140 (O_2140,N_19417,N_19315);
nand UO_2141 (O_2141,N_19128,N_19343);
and UO_2142 (O_2142,N_18277,N_19140);
and UO_2143 (O_2143,N_18827,N_18282);
nand UO_2144 (O_2144,N_18067,N_18294);
and UO_2145 (O_2145,N_18979,N_18970);
nand UO_2146 (O_2146,N_19245,N_18618);
nor UO_2147 (O_2147,N_18362,N_18415);
or UO_2148 (O_2148,N_19665,N_18328);
nand UO_2149 (O_2149,N_18911,N_19327);
and UO_2150 (O_2150,N_18070,N_18540);
nor UO_2151 (O_2151,N_19054,N_19192);
or UO_2152 (O_2152,N_19048,N_19538);
and UO_2153 (O_2153,N_19175,N_18384);
or UO_2154 (O_2154,N_19043,N_18038);
nor UO_2155 (O_2155,N_19025,N_19452);
and UO_2156 (O_2156,N_19618,N_19602);
nor UO_2157 (O_2157,N_18792,N_19523);
nand UO_2158 (O_2158,N_18450,N_18894);
and UO_2159 (O_2159,N_18586,N_19122);
or UO_2160 (O_2160,N_18210,N_19953);
nor UO_2161 (O_2161,N_19035,N_18476);
or UO_2162 (O_2162,N_19686,N_18905);
nor UO_2163 (O_2163,N_18913,N_18471);
nand UO_2164 (O_2164,N_18066,N_19801);
or UO_2165 (O_2165,N_18318,N_18907);
and UO_2166 (O_2166,N_19870,N_18994);
xor UO_2167 (O_2167,N_18399,N_18919);
and UO_2168 (O_2168,N_19595,N_18511);
nand UO_2169 (O_2169,N_18560,N_18792);
nand UO_2170 (O_2170,N_18155,N_18971);
nor UO_2171 (O_2171,N_18480,N_19752);
nand UO_2172 (O_2172,N_19131,N_18147);
nor UO_2173 (O_2173,N_19115,N_19551);
or UO_2174 (O_2174,N_18351,N_18589);
or UO_2175 (O_2175,N_18616,N_19768);
or UO_2176 (O_2176,N_18441,N_18565);
xor UO_2177 (O_2177,N_19855,N_18176);
or UO_2178 (O_2178,N_18660,N_18874);
nand UO_2179 (O_2179,N_18642,N_19607);
or UO_2180 (O_2180,N_18357,N_18942);
or UO_2181 (O_2181,N_19071,N_19466);
xnor UO_2182 (O_2182,N_18888,N_18345);
xor UO_2183 (O_2183,N_18742,N_18432);
nor UO_2184 (O_2184,N_18247,N_18818);
nor UO_2185 (O_2185,N_19263,N_19671);
or UO_2186 (O_2186,N_18449,N_19982);
and UO_2187 (O_2187,N_19612,N_19847);
and UO_2188 (O_2188,N_19896,N_18866);
nand UO_2189 (O_2189,N_19579,N_18986);
or UO_2190 (O_2190,N_18635,N_18691);
or UO_2191 (O_2191,N_19915,N_18859);
or UO_2192 (O_2192,N_18376,N_19085);
nor UO_2193 (O_2193,N_19775,N_19771);
or UO_2194 (O_2194,N_19172,N_19042);
or UO_2195 (O_2195,N_19693,N_18915);
or UO_2196 (O_2196,N_19039,N_19902);
or UO_2197 (O_2197,N_18216,N_18256);
nor UO_2198 (O_2198,N_18223,N_18586);
nor UO_2199 (O_2199,N_19205,N_19280);
xor UO_2200 (O_2200,N_18141,N_19269);
or UO_2201 (O_2201,N_19642,N_18551);
and UO_2202 (O_2202,N_19077,N_19056);
nor UO_2203 (O_2203,N_18962,N_19243);
nor UO_2204 (O_2204,N_19156,N_19047);
nand UO_2205 (O_2205,N_19775,N_19721);
xnor UO_2206 (O_2206,N_18828,N_18839);
and UO_2207 (O_2207,N_18428,N_18100);
nand UO_2208 (O_2208,N_18061,N_19893);
and UO_2209 (O_2209,N_18024,N_18966);
nand UO_2210 (O_2210,N_18429,N_19063);
xnor UO_2211 (O_2211,N_19844,N_18928);
nor UO_2212 (O_2212,N_18661,N_18304);
and UO_2213 (O_2213,N_19651,N_19097);
nor UO_2214 (O_2214,N_19923,N_18303);
nor UO_2215 (O_2215,N_19831,N_19132);
and UO_2216 (O_2216,N_19408,N_18986);
nand UO_2217 (O_2217,N_19025,N_19654);
nand UO_2218 (O_2218,N_19578,N_19098);
nand UO_2219 (O_2219,N_18962,N_18177);
xor UO_2220 (O_2220,N_18494,N_18697);
nor UO_2221 (O_2221,N_18218,N_19034);
or UO_2222 (O_2222,N_19577,N_18650);
nor UO_2223 (O_2223,N_18308,N_18662);
xor UO_2224 (O_2224,N_19928,N_18218);
nor UO_2225 (O_2225,N_18458,N_19144);
nand UO_2226 (O_2226,N_18516,N_18828);
nor UO_2227 (O_2227,N_18491,N_18120);
and UO_2228 (O_2228,N_19092,N_19176);
nor UO_2229 (O_2229,N_18062,N_19593);
nand UO_2230 (O_2230,N_18326,N_18298);
xnor UO_2231 (O_2231,N_18594,N_19410);
and UO_2232 (O_2232,N_19008,N_19670);
or UO_2233 (O_2233,N_19288,N_19314);
nand UO_2234 (O_2234,N_19695,N_18844);
nor UO_2235 (O_2235,N_18716,N_19147);
nor UO_2236 (O_2236,N_18224,N_18438);
nor UO_2237 (O_2237,N_19477,N_19403);
and UO_2238 (O_2238,N_18263,N_19681);
and UO_2239 (O_2239,N_19678,N_18842);
nand UO_2240 (O_2240,N_18963,N_18462);
or UO_2241 (O_2241,N_18621,N_18807);
and UO_2242 (O_2242,N_19772,N_19177);
nand UO_2243 (O_2243,N_18038,N_18725);
and UO_2244 (O_2244,N_18456,N_18209);
and UO_2245 (O_2245,N_19879,N_19974);
nand UO_2246 (O_2246,N_18655,N_19854);
xnor UO_2247 (O_2247,N_19143,N_18877);
nand UO_2248 (O_2248,N_18414,N_19788);
or UO_2249 (O_2249,N_19039,N_18426);
xnor UO_2250 (O_2250,N_18261,N_19865);
and UO_2251 (O_2251,N_18074,N_19124);
and UO_2252 (O_2252,N_19323,N_18288);
nand UO_2253 (O_2253,N_18656,N_18430);
nor UO_2254 (O_2254,N_18814,N_19687);
or UO_2255 (O_2255,N_19030,N_19079);
nor UO_2256 (O_2256,N_19030,N_18898);
xor UO_2257 (O_2257,N_19761,N_18157);
nand UO_2258 (O_2258,N_19149,N_19937);
nand UO_2259 (O_2259,N_19396,N_19743);
nor UO_2260 (O_2260,N_19553,N_18187);
and UO_2261 (O_2261,N_18201,N_19792);
nor UO_2262 (O_2262,N_18116,N_19351);
and UO_2263 (O_2263,N_18429,N_18840);
xnor UO_2264 (O_2264,N_18416,N_19335);
or UO_2265 (O_2265,N_18061,N_18688);
nand UO_2266 (O_2266,N_19214,N_18798);
nor UO_2267 (O_2267,N_18028,N_18706);
nand UO_2268 (O_2268,N_18186,N_19333);
nor UO_2269 (O_2269,N_18345,N_18609);
xor UO_2270 (O_2270,N_19223,N_19427);
or UO_2271 (O_2271,N_19815,N_19275);
nand UO_2272 (O_2272,N_18438,N_18149);
nor UO_2273 (O_2273,N_18719,N_19212);
nor UO_2274 (O_2274,N_19295,N_19167);
nand UO_2275 (O_2275,N_19812,N_19228);
nor UO_2276 (O_2276,N_19300,N_19077);
and UO_2277 (O_2277,N_18843,N_19689);
and UO_2278 (O_2278,N_18248,N_19201);
and UO_2279 (O_2279,N_18346,N_18004);
and UO_2280 (O_2280,N_18687,N_19972);
nor UO_2281 (O_2281,N_19967,N_19249);
and UO_2282 (O_2282,N_19667,N_19722);
nor UO_2283 (O_2283,N_18694,N_18298);
or UO_2284 (O_2284,N_19225,N_19277);
nor UO_2285 (O_2285,N_19670,N_19724);
and UO_2286 (O_2286,N_19947,N_19583);
nand UO_2287 (O_2287,N_19975,N_18184);
nand UO_2288 (O_2288,N_19638,N_18171);
and UO_2289 (O_2289,N_18204,N_18053);
nand UO_2290 (O_2290,N_19732,N_19144);
nor UO_2291 (O_2291,N_19240,N_18082);
nor UO_2292 (O_2292,N_19293,N_18645);
and UO_2293 (O_2293,N_18717,N_19895);
or UO_2294 (O_2294,N_18347,N_19023);
nand UO_2295 (O_2295,N_18343,N_19975);
nand UO_2296 (O_2296,N_18543,N_18025);
xnor UO_2297 (O_2297,N_18712,N_19059);
nand UO_2298 (O_2298,N_18800,N_19423);
and UO_2299 (O_2299,N_19260,N_18987);
nand UO_2300 (O_2300,N_19399,N_18510);
nor UO_2301 (O_2301,N_19882,N_18693);
nor UO_2302 (O_2302,N_19696,N_19809);
xor UO_2303 (O_2303,N_19884,N_19572);
xnor UO_2304 (O_2304,N_19372,N_18821);
nand UO_2305 (O_2305,N_18881,N_18082);
nor UO_2306 (O_2306,N_19578,N_18795);
or UO_2307 (O_2307,N_19073,N_18719);
nand UO_2308 (O_2308,N_18188,N_19344);
or UO_2309 (O_2309,N_19530,N_19583);
or UO_2310 (O_2310,N_19259,N_18524);
or UO_2311 (O_2311,N_18109,N_18938);
or UO_2312 (O_2312,N_18795,N_18602);
nor UO_2313 (O_2313,N_18025,N_19708);
xor UO_2314 (O_2314,N_19651,N_18936);
or UO_2315 (O_2315,N_19120,N_19875);
xnor UO_2316 (O_2316,N_18797,N_18919);
or UO_2317 (O_2317,N_18069,N_19185);
nor UO_2318 (O_2318,N_19270,N_18712);
or UO_2319 (O_2319,N_19587,N_19210);
or UO_2320 (O_2320,N_19430,N_19662);
nand UO_2321 (O_2321,N_18741,N_19906);
or UO_2322 (O_2322,N_18644,N_19539);
nor UO_2323 (O_2323,N_18945,N_18905);
nor UO_2324 (O_2324,N_19231,N_18852);
nor UO_2325 (O_2325,N_19236,N_19159);
or UO_2326 (O_2326,N_18463,N_18916);
nand UO_2327 (O_2327,N_19466,N_18401);
nand UO_2328 (O_2328,N_18914,N_19056);
nor UO_2329 (O_2329,N_19752,N_18531);
nor UO_2330 (O_2330,N_19396,N_18391);
or UO_2331 (O_2331,N_18236,N_18339);
or UO_2332 (O_2332,N_18145,N_18315);
nor UO_2333 (O_2333,N_18734,N_18348);
and UO_2334 (O_2334,N_18744,N_19037);
or UO_2335 (O_2335,N_18804,N_18366);
nor UO_2336 (O_2336,N_18123,N_19354);
nor UO_2337 (O_2337,N_18431,N_19382);
nor UO_2338 (O_2338,N_18033,N_19588);
or UO_2339 (O_2339,N_18027,N_18164);
and UO_2340 (O_2340,N_18552,N_18792);
nor UO_2341 (O_2341,N_19491,N_19722);
or UO_2342 (O_2342,N_18961,N_18251);
or UO_2343 (O_2343,N_18903,N_18826);
and UO_2344 (O_2344,N_19413,N_18469);
or UO_2345 (O_2345,N_18958,N_18820);
and UO_2346 (O_2346,N_18833,N_18279);
xor UO_2347 (O_2347,N_19280,N_18058);
nor UO_2348 (O_2348,N_19249,N_19852);
nand UO_2349 (O_2349,N_18541,N_19968);
nor UO_2350 (O_2350,N_19041,N_19967);
and UO_2351 (O_2351,N_19583,N_19376);
nor UO_2352 (O_2352,N_18643,N_18062);
and UO_2353 (O_2353,N_18437,N_18718);
or UO_2354 (O_2354,N_19419,N_19551);
nor UO_2355 (O_2355,N_19366,N_19370);
xor UO_2356 (O_2356,N_18723,N_18623);
nor UO_2357 (O_2357,N_19167,N_18794);
and UO_2358 (O_2358,N_19973,N_18045);
and UO_2359 (O_2359,N_19627,N_18249);
nor UO_2360 (O_2360,N_19106,N_18570);
nor UO_2361 (O_2361,N_18970,N_18811);
nand UO_2362 (O_2362,N_19086,N_18515);
or UO_2363 (O_2363,N_18769,N_19338);
and UO_2364 (O_2364,N_19651,N_18199);
nand UO_2365 (O_2365,N_19181,N_18374);
nor UO_2366 (O_2366,N_19914,N_18176);
nor UO_2367 (O_2367,N_18729,N_19098);
xor UO_2368 (O_2368,N_19002,N_18750);
nand UO_2369 (O_2369,N_19999,N_19964);
nor UO_2370 (O_2370,N_18040,N_19520);
or UO_2371 (O_2371,N_18654,N_18920);
nor UO_2372 (O_2372,N_18711,N_19039);
nor UO_2373 (O_2373,N_18893,N_19006);
nand UO_2374 (O_2374,N_18956,N_19412);
xnor UO_2375 (O_2375,N_18330,N_19892);
nor UO_2376 (O_2376,N_18217,N_19788);
nor UO_2377 (O_2377,N_18585,N_18288);
or UO_2378 (O_2378,N_19434,N_18118);
nand UO_2379 (O_2379,N_18370,N_19409);
and UO_2380 (O_2380,N_18051,N_18927);
nand UO_2381 (O_2381,N_19087,N_19104);
nand UO_2382 (O_2382,N_18073,N_19684);
and UO_2383 (O_2383,N_19805,N_19266);
nand UO_2384 (O_2384,N_19436,N_18491);
or UO_2385 (O_2385,N_19325,N_19865);
and UO_2386 (O_2386,N_19179,N_19819);
nand UO_2387 (O_2387,N_18793,N_19601);
nand UO_2388 (O_2388,N_19085,N_19913);
nand UO_2389 (O_2389,N_19144,N_19418);
or UO_2390 (O_2390,N_18947,N_18665);
and UO_2391 (O_2391,N_18673,N_18885);
xor UO_2392 (O_2392,N_19178,N_18479);
or UO_2393 (O_2393,N_19839,N_19503);
nand UO_2394 (O_2394,N_19028,N_19949);
and UO_2395 (O_2395,N_19061,N_18172);
or UO_2396 (O_2396,N_18931,N_18531);
nand UO_2397 (O_2397,N_19607,N_19022);
nor UO_2398 (O_2398,N_19308,N_18674);
nor UO_2399 (O_2399,N_19497,N_18193);
nor UO_2400 (O_2400,N_19582,N_18259);
or UO_2401 (O_2401,N_19125,N_18250);
nor UO_2402 (O_2402,N_18755,N_18212);
and UO_2403 (O_2403,N_18039,N_19817);
or UO_2404 (O_2404,N_19473,N_19639);
or UO_2405 (O_2405,N_19972,N_18638);
or UO_2406 (O_2406,N_18938,N_19281);
and UO_2407 (O_2407,N_18860,N_18578);
xor UO_2408 (O_2408,N_19956,N_18257);
nand UO_2409 (O_2409,N_18084,N_18977);
nor UO_2410 (O_2410,N_19671,N_19453);
nand UO_2411 (O_2411,N_18660,N_19648);
nand UO_2412 (O_2412,N_19884,N_19500);
and UO_2413 (O_2413,N_19812,N_18665);
and UO_2414 (O_2414,N_19813,N_19564);
nor UO_2415 (O_2415,N_18477,N_18117);
nor UO_2416 (O_2416,N_19821,N_18694);
nor UO_2417 (O_2417,N_19696,N_19792);
nand UO_2418 (O_2418,N_18380,N_18736);
nor UO_2419 (O_2419,N_19752,N_18769);
nor UO_2420 (O_2420,N_19168,N_18570);
nor UO_2421 (O_2421,N_19154,N_18078);
nor UO_2422 (O_2422,N_18087,N_18950);
and UO_2423 (O_2423,N_18841,N_19624);
and UO_2424 (O_2424,N_19966,N_18983);
and UO_2425 (O_2425,N_18650,N_19517);
or UO_2426 (O_2426,N_19828,N_18849);
and UO_2427 (O_2427,N_18038,N_19186);
or UO_2428 (O_2428,N_18095,N_18021);
xor UO_2429 (O_2429,N_19995,N_18010);
and UO_2430 (O_2430,N_19374,N_19562);
and UO_2431 (O_2431,N_19265,N_18040);
nand UO_2432 (O_2432,N_18050,N_18810);
and UO_2433 (O_2433,N_18550,N_19257);
nand UO_2434 (O_2434,N_18474,N_19624);
and UO_2435 (O_2435,N_19445,N_18472);
nor UO_2436 (O_2436,N_18550,N_18854);
nor UO_2437 (O_2437,N_19980,N_19302);
nor UO_2438 (O_2438,N_19401,N_19429);
nand UO_2439 (O_2439,N_19150,N_19144);
nand UO_2440 (O_2440,N_19365,N_19324);
and UO_2441 (O_2441,N_19812,N_18152);
nor UO_2442 (O_2442,N_18396,N_18399);
nor UO_2443 (O_2443,N_18692,N_19050);
nand UO_2444 (O_2444,N_18389,N_19627);
or UO_2445 (O_2445,N_18707,N_19047);
xnor UO_2446 (O_2446,N_18833,N_19187);
and UO_2447 (O_2447,N_19442,N_18184);
nand UO_2448 (O_2448,N_19948,N_19897);
or UO_2449 (O_2449,N_18109,N_19076);
xor UO_2450 (O_2450,N_18917,N_19667);
or UO_2451 (O_2451,N_18743,N_18288);
or UO_2452 (O_2452,N_18719,N_18327);
nand UO_2453 (O_2453,N_19876,N_19775);
nor UO_2454 (O_2454,N_19071,N_18805);
and UO_2455 (O_2455,N_18071,N_19646);
nand UO_2456 (O_2456,N_19862,N_18251);
and UO_2457 (O_2457,N_19698,N_19120);
nor UO_2458 (O_2458,N_18889,N_18004);
nor UO_2459 (O_2459,N_18613,N_19582);
nor UO_2460 (O_2460,N_18281,N_18646);
and UO_2461 (O_2461,N_18754,N_19228);
nor UO_2462 (O_2462,N_19574,N_18858);
and UO_2463 (O_2463,N_19814,N_18210);
or UO_2464 (O_2464,N_18160,N_18880);
and UO_2465 (O_2465,N_18114,N_18285);
or UO_2466 (O_2466,N_19610,N_18559);
nand UO_2467 (O_2467,N_19548,N_19252);
or UO_2468 (O_2468,N_19795,N_19316);
nor UO_2469 (O_2469,N_18907,N_18188);
and UO_2470 (O_2470,N_18579,N_19808);
nor UO_2471 (O_2471,N_19941,N_18860);
or UO_2472 (O_2472,N_19534,N_19491);
nor UO_2473 (O_2473,N_19821,N_19425);
nor UO_2474 (O_2474,N_19643,N_18797);
xor UO_2475 (O_2475,N_19563,N_19415);
nand UO_2476 (O_2476,N_18173,N_18138);
nand UO_2477 (O_2477,N_18563,N_18754);
nor UO_2478 (O_2478,N_18391,N_19137);
or UO_2479 (O_2479,N_19651,N_18100);
and UO_2480 (O_2480,N_18832,N_19026);
or UO_2481 (O_2481,N_19706,N_19412);
xor UO_2482 (O_2482,N_18632,N_18093);
nand UO_2483 (O_2483,N_19812,N_18933);
nand UO_2484 (O_2484,N_19224,N_19110);
or UO_2485 (O_2485,N_19025,N_18585);
or UO_2486 (O_2486,N_18571,N_18250);
nand UO_2487 (O_2487,N_19834,N_18644);
nor UO_2488 (O_2488,N_18599,N_18028);
or UO_2489 (O_2489,N_18641,N_18197);
nand UO_2490 (O_2490,N_18983,N_19176);
nand UO_2491 (O_2491,N_19509,N_18798);
nand UO_2492 (O_2492,N_18800,N_18665);
or UO_2493 (O_2493,N_19317,N_19816);
or UO_2494 (O_2494,N_19143,N_19422);
nor UO_2495 (O_2495,N_19733,N_18498);
nor UO_2496 (O_2496,N_18063,N_19715);
nor UO_2497 (O_2497,N_18101,N_19301);
nand UO_2498 (O_2498,N_18083,N_18342);
and UO_2499 (O_2499,N_18411,N_18442);
endmodule