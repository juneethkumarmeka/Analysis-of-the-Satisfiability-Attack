module basic_2000_20000_2500_10_levels_10xor_2(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999;
nor U0 (N_0,In_445,In_1073);
and U1 (N_1,In_1639,In_179);
or U2 (N_2,In_1994,In_879);
or U3 (N_3,In_57,In_1518);
xnor U4 (N_4,In_841,In_21);
xor U5 (N_5,In_85,In_183);
nand U6 (N_6,In_986,In_1059);
nor U7 (N_7,In_1308,In_1752);
nand U8 (N_8,In_1386,In_426);
nor U9 (N_9,In_391,In_814);
and U10 (N_10,In_610,In_1103);
nand U11 (N_11,In_1033,In_586);
nand U12 (N_12,In_608,In_1420);
nor U13 (N_13,In_977,In_1254);
or U14 (N_14,In_538,In_1324);
nor U15 (N_15,In_200,In_431);
or U16 (N_16,In_1086,In_1751);
xor U17 (N_17,In_1924,In_1910);
xnor U18 (N_18,In_1002,In_1432);
and U19 (N_19,In_1301,In_397);
nand U20 (N_20,In_272,In_1045);
xnor U21 (N_21,In_74,In_1605);
nand U22 (N_22,In_1495,In_1366);
and U23 (N_23,In_1126,In_1606);
nor U24 (N_24,In_1703,In_146);
and U25 (N_25,In_1768,In_1271);
nor U26 (N_26,In_1967,In_1593);
and U27 (N_27,In_296,In_1841);
or U28 (N_28,In_725,In_650);
xnor U29 (N_29,In_411,In_1584);
and U30 (N_30,In_845,In_1995);
nor U31 (N_31,In_681,In_522);
nand U32 (N_32,In_498,In_56);
nand U33 (N_33,In_1672,In_679);
and U34 (N_34,In_828,In_1552);
or U35 (N_35,In_1394,In_1705);
and U36 (N_36,In_1160,In_988);
xor U37 (N_37,In_688,In_478);
or U38 (N_38,In_469,In_16);
xor U39 (N_39,In_1834,In_261);
xor U40 (N_40,In_602,In_1999);
and U41 (N_41,In_62,In_1919);
nor U42 (N_42,In_1288,In_1558);
xnor U43 (N_43,In_1978,In_936);
or U44 (N_44,In_784,In_511);
nand U45 (N_45,In_435,In_1296);
nor U46 (N_46,In_1687,In_449);
or U47 (N_47,In_1966,In_744);
nand U48 (N_48,In_121,In_1776);
and U49 (N_49,In_181,In_402);
nor U50 (N_50,In_967,In_849);
and U51 (N_51,In_491,In_790);
and U52 (N_52,In_182,In_1643);
nor U53 (N_53,In_160,In_858);
xnor U54 (N_54,In_1917,In_1772);
and U55 (N_55,In_1057,In_1704);
and U56 (N_56,In_571,In_1803);
nor U57 (N_57,In_769,In_1331);
and U58 (N_58,In_1036,In_554);
or U59 (N_59,In_100,In_924);
and U60 (N_60,In_1303,In_351);
or U61 (N_61,In_606,In_505);
or U62 (N_62,In_526,In_882);
and U63 (N_63,In_980,In_1276);
xnor U64 (N_64,In_477,In_1922);
xor U65 (N_65,In_937,In_990);
nand U66 (N_66,In_1938,In_163);
nand U67 (N_67,In_330,In_532);
nand U68 (N_68,In_1808,In_68);
or U69 (N_69,In_1594,In_177);
and U70 (N_70,In_1476,In_780);
nand U71 (N_71,In_695,In_61);
nor U72 (N_72,In_1670,In_1529);
xor U73 (N_73,In_953,In_1852);
or U74 (N_74,In_5,In_1790);
xor U75 (N_75,In_1202,In_983);
and U76 (N_76,In_765,In_208);
and U77 (N_77,In_22,In_752);
and U78 (N_78,In_1491,In_1141);
and U79 (N_79,In_1031,In_1872);
xnor U80 (N_80,In_1333,In_35);
xnor U81 (N_81,In_1058,In_254);
nand U82 (N_82,In_1167,In_603);
nor U83 (N_83,In_783,In_369);
xnor U84 (N_84,In_859,In_791);
nand U85 (N_85,In_1765,In_1415);
xnor U86 (N_86,In_1983,In_1497);
and U87 (N_87,In_1216,In_1610);
nand U88 (N_88,In_732,In_1480);
nand U89 (N_89,In_572,In_1946);
and U90 (N_90,In_1267,In_394);
and U91 (N_91,In_552,In_617);
or U92 (N_92,In_867,In_689);
and U93 (N_93,In_358,In_1973);
xnor U94 (N_94,In_53,In_1256);
nor U95 (N_95,In_1678,In_1253);
nor U96 (N_96,In_551,In_246);
or U97 (N_97,In_1589,In_865);
nand U98 (N_98,In_1258,In_1169);
nand U99 (N_99,In_1306,In_1121);
nand U100 (N_100,In_837,In_999);
nand U101 (N_101,In_782,In_1475);
nand U102 (N_102,In_388,In_1343);
or U103 (N_103,In_1070,In_1025);
nor U104 (N_104,In_1322,In_143);
nor U105 (N_105,In_1454,In_1578);
nand U106 (N_106,In_805,In_622);
nand U107 (N_107,In_803,In_1088);
and U108 (N_108,In_747,In_103);
nor U109 (N_109,In_1282,In_620);
nor U110 (N_110,In_1375,In_1285);
nand U111 (N_111,In_1876,In_169);
nand U112 (N_112,In_1647,In_777);
nor U113 (N_113,In_1051,In_420);
or U114 (N_114,In_640,In_925);
xor U115 (N_115,In_1812,In_1470);
nor U116 (N_116,In_618,In_1775);
nand U117 (N_117,In_851,In_1094);
and U118 (N_118,In_1758,In_1206);
nor U119 (N_119,In_885,In_901);
or U120 (N_120,In_728,In_675);
xor U121 (N_121,In_140,In_429);
nand U122 (N_122,In_1614,In_318);
or U123 (N_123,In_735,In_408);
and U124 (N_124,In_1311,In_1952);
or U125 (N_125,In_1891,In_648);
or U126 (N_126,In_1223,In_1598);
nor U127 (N_127,In_1419,In_243);
and U128 (N_128,In_40,In_663);
and U129 (N_129,In_1535,In_1753);
or U130 (N_130,In_1185,In_1607);
xor U131 (N_131,In_1747,In_731);
or U132 (N_132,In_952,In_1261);
and U133 (N_133,In_1627,In_1543);
xnor U134 (N_134,In_1871,In_30);
and U135 (N_135,In_709,In_806);
or U136 (N_136,In_1097,In_138);
nand U137 (N_137,In_549,In_1920);
and U138 (N_138,In_1733,In_543);
nand U139 (N_139,In_150,In_1448);
nand U140 (N_140,In_786,In_155);
xnor U141 (N_141,In_1942,In_438);
or U142 (N_142,In_105,In_1136);
xnor U143 (N_143,In_975,In_1909);
or U144 (N_144,In_89,In_935);
and U145 (N_145,In_1717,In_199);
and U146 (N_146,In_1797,In_1958);
nand U147 (N_147,In_1948,In_678);
xor U148 (N_148,In_1934,In_518);
or U149 (N_149,In_1950,In_877);
or U150 (N_150,In_1810,In_1707);
or U151 (N_151,In_993,In_779);
nor U152 (N_152,In_1989,In_934);
xor U153 (N_153,In_587,In_943);
xor U154 (N_154,In_940,In_1645);
nor U155 (N_155,In_792,In_1653);
nor U156 (N_156,In_361,In_1686);
xor U157 (N_157,In_1907,In_298);
and U158 (N_158,In_166,In_497);
nor U159 (N_159,In_24,In_122);
nand U160 (N_160,In_323,In_291);
nand U161 (N_161,In_1894,In_1706);
and U162 (N_162,In_1550,In_1673);
nor U163 (N_163,In_15,In_701);
nor U164 (N_164,In_1874,In_824);
or U165 (N_165,In_1024,In_510);
or U166 (N_166,In_1591,In_613);
nor U167 (N_167,In_718,In_1344);
nor U168 (N_168,In_1561,In_1131);
nand U169 (N_169,In_1338,In_50);
nor U170 (N_170,In_615,In_1755);
nand U171 (N_171,In_37,In_702);
or U172 (N_172,In_674,In_1806);
nand U173 (N_173,In_564,In_185);
nand U174 (N_174,In_338,In_174);
xnor U175 (N_175,In_1538,In_1574);
nand U176 (N_176,In_1179,In_1323);
and U177 (N_177,In_123,In_1139);
nand U178 (N_178,In_1878,In_167);
and U179 (N_179,In_736,In_1349);
nor U180 (N_180,In_1109,In_316);
xnor U181 (N_181,In_1243,In_164);
nor U182 (N_182,In_873,In_631);
xnor U183 (N_183,In_897,In_39);
nor U184 (N_184,In_1161,In_342);
nor U185 (N_185,In_191,In_1230);
nor U186 (N_186,In_868,In_739);
or U187 (N_187,In_34,In_1229);
and U188 (N_188,In_706,In_1882);
and U189 (N_189,In_1617,In_793);
nor U190 (N_190,In_1905,In_1113);
xor U191 (N_191,In_1397,In_1832);
xor U192 (N_192,In_1793,In_946);
nor U193 (N_193,In_1728,In_846);
nor U194 (N_194,In_738,In_748);
and U195 (N_195,In_1547,In_726);
nor U196 (N_196,In_1955,In_515);
nor U197 (N_197,In_1684,In_1210);
nand U198 (N_198,In_1588,In_344);
nor U199 (N_199,In_1052,In_1988);
nand U200 (N_200,In_978,In_1326);
nand U201 (N_201,In_939,In_1744);
xor U202 (N_202,In_447,In_238);
and U203 (N_203,In_651,In_839);
xor U204 (N_204,In_754,In_1177);
and U205 (N_205,In_1587,In_1043);
or U206 (N_206,In_1341,In_1232);
and U207 (N_207,In_161,In_644);
nor U208 (N_208,In_1295,In_1355);
xor U209 (N_209,In_1135,In_1368);
nor U210 (N_210,In_1644,In_813);
xor U211 (N_211,In_1601,In_557);
or U212 (N_212,In_1227,In_1119);
or U213 (N_213,In_1723,In_1899);
and U214 (N_214,In_11,In_1443);
or U215 (N_215,In_1123,In_153);
xor U216 (N_216,In_1219,In_1337);
nor U217 (N_217,In_364,In_821);
and U218 (N_218,In_1925,In_743);
and U219 (N_219,In_1949,In_611);
xnor U220 (N_220,In_470,In_1947);
or U221 (N_221,In_1888,In_114);
nand U222 (N_222,In_1944,In_1661);
nand U223 (N_223,In_365,In_268);
and U224 (N_224,In_1034,In_109);
xor U225 (N_225,In_1399,In_951);
and U226 (N_226,In_1778,In_797);
or U227 (N_227,In_482,In_984);
nor U228 (N_228,In_304,In_1379);
xor U229 (N_229,In_1467,In_1280);
xnor U230 (N_230,In_290,In_267);
nor U231 (N_231,In_1218,In_544);
and U232 (N_232,In_286,In_1464);
nor U233 (N_233,In_1650,In_1545);
or U234 (N_234,In_1204,In_1055);
and U235 (N_235,In_1164,In_959);
and U236 (N_236,In_1275,In_1054);
nor U237 (N_237,In_950,In_833);
and U238 (N_238,In_488,In_830);
nor U239 (N_239,In_1691,In_1151);
nand U240 (N_240,In_1798,In_919);
nand U241 (N_241,In_1396,In_1353);
or U242 (N_242,In_1273,In_152);
or U243 (N_243,In_637,In_698);
nand U244 (N_244,In_1975,In_1367);
or U245 (N_245,In_1245,In_1864);
and U246 (N_246,In_457,In_1390);
nor U247 (N_247,In_1238,In_1101);
nor U248 (N_248,In_46,In_836);
and U249 (N_249,In_1392,In_1609);
and U250 (N_250,In_931,In_1828);
and U251 (N_251,In_319,In_1567);
xnor U252 (N_252,In_1003,In_900);
xor U253 (N_253,In_560,In_1783);
xnor U254 (N_254,In_1608,In_501);
and U255 (N_255,In_1130,In_630);
nor U256 (N_256,In_635,In_374);
nor U257 (N_257,In_619,In_25);
xor U258 (N_258,In_1168,In_1028);
nand U259 (N_259,In_656,In_1377);
or U260 (N_260,In_740,In_759);
xor U261 (N_261,In_1671,In_452);
and U262 (N_262,In_1365,In_1436);
or U263 (N_263,In_1359,In_981);
and U264 (N_264,In_1731,In_1056);
or U265 (N_265,In_1940,In_1496);
nor U266 (N_266,In_1615,In_545);
or U267 (N_267,In_412,In_144);
and U268 (N_268,In_3,In_834);
xnor U269 (N_269,In_43,In_652);
and U270 (N_270,In_72,In_370);
xnor U271 (N_271,In_773,In_712);
and U272 (N_272,In_992,In_948);
nor U273 (N_273,In_400,In_279);
or U274 (N_274,In_1416,In_1340);
or U275 (N_275,In_909,In_1465);
or U276 (N_276,In_1203,In_1603);
nand U277 (N_277,In_1823,In_93);
nor U278 (N_278,In_1431,In_881);
nand U279 (N_279,In_1079,In_1345);
xor U280 (N_280,In_1582,In_550);
nor U281 (N_281,In_755,In_48);
or U282 (N_282,In_87,In_230);
xnor U283 (N_283,In_96,In_1821);
or U284 (N_284,In_434,In_717);
or U285 (N_285,In_801,In_1649);
and U286 (N_286,In_807,In_1725);
and U287 (N_287,In_1679,In_1462);
or U288 (N_288,In_276,In_216);
xnor U289 (N_289,In_1279,In_1968);
nand U290 (N_290,In_1696,In_1176);
nand U291 (N_291,In_1805,In_1885);
or U292 (N_292,In_1861,In_581);
nor U293 (N_293,In_1815,In_1100);
xor U294 (N_294,In_212,In_154);
nand U295 (N_295,In_719,In_1564);
and U296 (N_296,In_1393,In_264);
nor U297 (N_297,In_287,In_1134);
or U298 (N_298,In_585,In_250);
nand U299 (N_299,In_366,In_1847);
or U300 (N_300,In_812,In_927);
and U301 (N_301,In_1076,In_489);
or U302 (N_302,In_471,In_1865);
nand U303 (N_303,In_184,In_1486);
and U304 (N_304,In_680,In_653);
nor U305 (N_305,In_775,In_415);
and U306 (N_306,In_1387,In_20);
xor U307 (N_307,In_1182,In_1674);
xnor U308 (N_308,In_1658,In_235);
and U309 (N_309,In_1921,In_750);
nor U310 (N_310,In_1270,In_513);
nor U311 (N_311,In_1047,In_1314);
nand U312 (N_312,In_1181,In_343);
xor U313 (N_313,In_772,In_1931);
nor U314 (N_314,In_1522,In_789);
xnor U315 (N_315,In_1466,In_159);
and U316 (N_316,In_893,In_26);
and U317 (N_317,In_1050,In_1665);
and U318 (N_318,In_843,In_1620);
xnor U319 (N_319,In_1362,In_938);
or U320 (N_320,In_1493,In_1425);
nor U321 (N_321,In_1423,In_215);
xnor U322 (N_322,In_1657,In_1499);
nand U323 (N_323,In_187,In_69);
or U324 (N_324,In_942,In_1746);
xor U325 (N_325,In_49,In_472);
or U326 (N_326,In_357,In_1640);
nand U327 (N_327,In_1622,In_998);
nand U328 (N_328,In_1896,In_1456);
nand U329 (N_329,In_1022,In_1540);
nor U330 (N_330,In_217,In_7);
xnor U331 (N_331,In_1681,In_1251);
xnor U332 (N_332,In_1265,In_1427);
and U333 (N_333,In_1463,In_1996);
nor U334 (N_334,In_1818,In_1621);
nand U335 (N_335,In_110,In_51);
nor U336 (N_336,In_874,In_1374);
or U337 (N_337,In_1114,In_1690);
xor U338 (N_338,In_328,In_1260);
and U339 (N_339,In_204,In_381);
and U340 (N_340,In_263,In_913);
xnor U341 (N_341,In_730,In_891);
nand U342 (N_342,In_741,In_1831);
xnor U343 (N_343,In_0,In_629);
or U344 (N_344,In_240,In_1906);
nor U345 (N_345,In_1774,In_1128);
nor U346 (N_346,In_90,In_245);
nand U347 (N_347,In_1546,In_1817);
and U348 (N_348,In_219,In_384);
and U349 (N_349,In_141,In_172);
nand U350 (N_350,In_233,In_1277);
nor U351 (N_351,In_1009,In_1811);
xor U352 (N_352,In_1618,In_912);
nand U353 (N_353,In_107,In_292);
nor U354 (N_354,In_816,In_1802);
or U355 (N_355,In_1078,In_521);
xor U356 (N_356,In_173,In_1520);
or U357 (N_357,In_1032,In_1524);
and U358 (N_358,In_205,In_1963);
xnor U359 (N_359,In_294,In_1830);
nor U360 (N_360,In_373,In_300);
or U361 (N_361,In_54,In_607);
nand U362 (N_362,In_1848,In_527);
or U363 (N_363,In_1510,In_353);
nand U364 (N_364,In_1042,In_623);
nor U365 (N_365,In_593,In_1992);
and U366 (N_366,In_1211,In_55);
nand U367 (N_367,In_523,In_525);
nor U368 (N_368,In_295,In_1631);
nand U369 (N_369,In_818,In_98);
xor U370 (N_370,In_742,In_1595);
nand U371 (N_371,In_616,In_1110);
nand U372 (N_372,In_387,In_1590);
or U373 (N_373,In_1422,In_579);
or U374 (N_374,In_1208,In_1249);
xor U375 (N_375,In_1675,In_1976);
nand U376 (N_376,In_809,In_722);
xnor U377 (N_377,In_1129,In_857);
or U378 (N_378,In_178,In_604);
nor U379 (N_379,In_410,In_856);
or U380 (N_380,In_339,In_1702);
nor U381 (N_381,In_414,In_1735);
nand U382 (N_382,In_462,In_380);
nor U383 (N_383,In_1521,In_1859);
nor U384 (N_384,In_371,In_293);
xnor U385 (N_385,In_536,In_850);
nand U386 (N_386,In_1987,In_1274);
or U387 (N_387,In_1483,In_1077);
nand U388 (N_388,In_1556,In_331);
xor U389 (N_389,In_1039,In_991);
xor U390 (N_390,In_262,In_1255);
nor U391 (N_391,In_1759,In_770);
xor U392 (N_392,In_1886,In_1557);
nand U393 (N_393,In_1325,In_1846);
or U394 (N_394,In_788,In_1741);
xor U395 (N_395,In_271,In_1877);
nand U396 (N_396,In_664,In_1660);
nand U397 (N_397,In_1791,In_996);
nor U398 (N_398,In_1668,In_835);
and U399 (N_399,In_766,In_479);
or U400 (N_400,In_1318,In_1626);
and U401 (N_401,In_1289,In_1195);
nand U402 (N_402,In_1585,In_252);
nand U403 (N_403,In_768,In_229);
xor U404 (N_404,In_1482,In_1898);
nor U405 (N_405,In_142,In_320);
or U406 (N_406,In_1069,In_1143);
xnor U407 (N_407,In_1347,In_1514);
and U408 (N_408,In_1586,In_1172);
or U409 (N_409,In_979,In_201);
and U410 (N_410,In_480,In_1575);
nand U411 (N_411,In_944,In_1236);
and U412 (N_412,In_1105,In_1310);
nor U413 (N_413,In_1426,In_91);
xnor U414 (N_414,In_1175,In_186);
and U415 (N_415,In_1373,In_1224);
nor U416 (N_416,In_1091,In_1201);
and U417 (N_417,In_440,In_454);
nand U418 (N_418,In_1980,In_1228);
nor U419 (N_419,In_605,In_335);
nor U420 (N_420,In_227,In_1667);
and U421 (N_421,In_724,In_377);
nor U422 (N_422,In_221,In_125);
or U423 (N_423,In_463,In_1272);
or U424 (N_424,In_1035,In_441);
nor U425 (N_425,In_1320,In_941);
nand U426 (N_426,In_1112,In_1299);
nand U427 (N_427,In_1071,In_1619);
and U428 (N_428,In_28,In_658);
or U429 (N_429,In_1655,In_455);
xnor U430 (N_430,In_251,In_714);
xnor U431 (N_431,In_1484,In_202);
or U432 (N_432,In_1038,In_911);
xor U433 (N_433,In_247,In_493);
xor U434 (N_434,In_802,In_17);
nand U435 (N_435,In_1478,In_665);
xor U436 (N_436,In_546,In_1508);
nand U437 (N_437,In_1321,In_692);
xnor U438 (N_438,In_222,In_982);
and U439 (N_439,In_1727,In_363);
nor U440 (N_440,In_1178,In_907);
nand U441 (N_441,In_1441,In_583);
nand U442 (N_442,In_1889,In_570);
or U443 (N_443,In_425,In_1796);
nand U444 (N_444,In_367,In_1469);
nor U445 (N_445,In_829,In_278);
and U446 (N_446,In_461,In_76);
nand U447 (N_447,In_1074,In_1205);
nand U448 (N_448,In_727,In_1361);
nor U449 (N_449,In_1880,In_1548);
nand U450 (N_450,In_1984,In_6);
nand U451 (N_451,In_337,In_1406);
and U452 (N_452,In_947,In_1554);
nor U453 (N_453,In_1242,In_1838);
nor U454 (N_454,In_347,In_1468);
and U455 (N_455,In_1870,In_285);
or U456 (N_456,In_487,In_890);
and U457 (N_457,In_1066,In_1146);
and U458 (N_458,In_1893,In_1695);
and U459 (N_459,In_534,In_1278);
or U460 (N_460,In_853,In_149);
and U461 (N_461,In_1525,In_474);
nor U462 (N_462,In_1153,In_506);
nand U463 (N_463,In_111,In_1669);
and U464 (N_464,In_10,In_1300);
nand U465 (N_465,In_156,In_1986);
xor U466 (N_466,In_1434,In_737);
nor U467 (N_467,In_1804,In_1352);
nor U468 (N_468,In_1459,In_1000);
and U469 (N_469,In_1246,In_1440);
nand U470 (N_470,In_1264,In_417);
or U471 (N_471,In_641,In_244);
and U472 (N_472,In_1104,In_1965);
and U473 (N_473,In_1157,In_1851);
or U474 (N_474,In_1309,In_962);
and U475 (N_475,In_1715,In_284);
nand U476 (N_476,In_643,In_108);
nor U477 (N_477,In_1807,In_465);
or U478 (N_478,In_1879,In_1395);
xnor U479 (N_479,In_439,In_1633);
and U480 (N_480,In_628,In_450);
nor U481 (N_481,In_1162,In_1090);
and U482 (N_482,In_1531,In_1881);
nand U483 (N_483,In_1287,In_1794);
or U484 (N_484,In_955,In_77);
nor U485 (N_485,In_705,In_1235);
or U486 (N_486,In_1516,In_1080);
nand U487 (N_487,In_423,In_1855);
nor U488 (N_488,In_649,In_1981);
nor U489 (N_489,In_1442,In_270);
xor U490 (N_490,In_1819,In_119);
and U491 (N_491,In_862,In_485);
xnor U492 (N_492,In_466,In_672);
nand U493 (N_493,In_1064,In_1269);
and U494 (N_494,In_1579,In_277);
xor U495 (N_495,In_964,In_1356);
nor U496 (N_496,In_811,In_350);
and U497 (N_497,In_171,In_317);
nand U498 (N_498,In_1754,In_1858);
nand U499 (N_499,In_375,In_228);
nand U500 (N_500,In_1960,In_1029);
nor U501 (N_501,In_869,In_1305);
nor U502 (N_502,In_1936,In_671);
nand U503 (N_503,In_1093,In_12);
nor U504 (N_504,In_1824,In_1890);
or U505 (N_505,In_1785,In_578);
or U506 (N_506,In_1213,In_1358);
nand U507 (N_507,In_1724,In_1664);
or U508 (N_508,In_1676,In_1700);
or U509 (N_509,In_1194,In_27);
nor U510 (N_510,In_1822,In_255);
or U511 (N_511,In_707,In_1472);
nor U512 (N_512,In_1604,In_758);
nand U513 (N_513,In_1625,In_147);
nor U514 (N_514,In_1451,In_914);
or U515 (N_515,In_1542,In_676);
and U516 (N_516,In_257,In_334);
nor U517 (N_517,In_976,In_561);
nand U518 (N_518,In_1062,In_659);
or U519 (N_519,In_883,In_753);
nor U520 (N_520,In_669,In_484);
nor U521 (N_521,In_1656,In_1628);
nor U522 (N_522,In_433,In_1027);
or U523 (N_523,In_269,In_632);
and U524 (N_524,In_396,In_580);
or U525 (N_525,In_517,In_139);
nand U526 (N_526,In_81,In_589);
xor U527 (N_527,In_430,In_733);
or U528 (N_528,In_1685,In_1197);
or U529 (N_529,In_1266,In_1217);
and U530 (N_530,In_905,In_1503);
nand U531 (N_531,In_99,In_647);
xor U532 (N_532,In_646,In_355);
or U533 (N_533,In_442,In_1106);
nand U534 (N_534,In_823,In_315);
xnor U535 (N_535,In_1332,In_1757);
xor U536 (N_536,In_568,In_398);
or U537 (N_537,In_1638,In_127);
nor U538 (N_538,In_1708,In_1600);
nand U539 (N_539,In_1826,In_1901);
nand U540 (N_540,In_1929,In_1458);
xor U541 (N_541,In_958,In_1125);
nor U542 (N_542,In_781,In_1293);
nand U543 (N_543,In_590,In_1430);
and U544 (N_544,In_1869,In_573);
or U545 (N_545,In_1839,In_1061);
and U546 (N_546,In_281,In_1363);
xor U547 (N_547,In_336,In_120);
or U548 (N_548,In_1257,In_1714);
nor U549 (N_549,In_842,In_1187);
nand U550 (N_550,In_776,In_1449);
and U551 (N_551,In_903,In_102);
or U552 (N_552,In_1165,In_866);
nor U553 (N_553,In_1883,In_1350);
nor U554 (N_554,In_1549,In_1099);
or U555 (N_555,In_654,In_1502);
nand U556 (N_556,In_340,In_274);
and U557 (N_557,In_422,In_1750);
nand U558 (N_558,In_508,In_542);
xnor U559 (N_559,In_574,In_468);
xnor U560 (N_560,In_1351,In_1118);
nand U561 (N_561,In_582,In_926);
xnor U562 (N_562,In_1513,In_1207);
nand U563 (N_563,In_729,In_206);
and U564 (N_564,In_1935,In_1401);
and U565 (N_565,In_1215,In_282);
or U566 (N_566,In_313,In_1192);
xnor U567 (N_567,In_1312,In_1654);
nor U568 (N_568,In_224,In_1993);
or U569 (N_569,In_1346,In_1581);
xnor U570 (N_570,In_588,In_595);
xor U571 (N_571,In_1457,In_1756);
nor U572 (N_572,In_1505,In_1364);
nand U573 (N_573,In_1382,In_356);
xor U574 (N_574,In_467,In_763);
or U575 (N_575,In_75,In_1761);
or U576 (N_576,In_1021,In_148);
or U577 (N_577,In_749,In_662);
xnor U578 (N_578,In_1102,In_1792);
nand U579 (N_579,In_453,In_1405);
nand U580 (N_580,In_1711,In_1836);
nor U581 (N_581,In_112,In_870);
nor U582 (N_582,In_157,In_700);
or U583 (N_583,In_1297,In_686);
and U584 (N_584,In_957,In_1536);
nand U585 (N_585,In_1504,In_918);
xnor U586 (N_586,In_537,In_495);
or U587 (N_587,In_910,In_31);
nand U588 (N_588,In_1262,In_660);
xnor U589 (N_589,In_710,In_516);
nand U590 (N_590,In_1250,In_1541);
nor U591 (N_591,In_1414,In_794);
nor U592 (N_592,In_137,In_4);
xor U593 (N_593,In_1418,In_1148);
and U594 (N_594,In_889,In_473);
or U595 (N_595,In_1961,In_1868);
or U596 (N_596,In_464,In_299);
and U597 (N_597,In_97,In_673);
and U598 (N_598,In_1539,In_1718);
xor U599 (N_599,In_825,In_180);
and U600 (N_600,In_1553,In_902);
xnor U601 (N_601,In_66,In_1450);
xor U602 (N_602,In_852,In_1698);
and U603 (N_603,In_972,In_1829);
nor U604 (N_604,In_1012,In_1471);
or U605 (N_605,In_569,In_1391);
nor U606 (N_606,In_418,In_368);
or U607 (N_607,In_389,In_530);
nor U608 (N_608,In_458,In_1500);
and U609 (N_609,In_945,In_1928);
and U610 (N_610,In_1184,In_83);
and U611 (N_611,In_1231,In_18);
or U612 (N_612,In_1460,In_1760);
xor U613 (N_613,In_1298,In_424);
xor U614 (N_614,In_1154,In_1044);
and U615 (N_615,In_1597,In_1138);
or U616 (N_616,In_1651,In_1384);
or U617 (N_617,In_1334,In_540);
xnor U618 (N_618,In_1895,In_1611);
nor U619 (N_619,In_1412,In_1998);
nor U620 (N_620,In_1937,In_1302);
nor U621 (N_621,In_136,In_625);
nand U622 (N_622,In_1122,In_1875);
or U623 (N_623,In_1013,In_884);
xnor U624 (N_624,In_104,In_437);
and U625 (N_625,In_406,In_645);
nor U626 (N_626,In_1190,In_915);
or U627 (N_627,In_819,In_1354);
xor U628 (N_628,In_432,In_887);
nor U629 (N_629,In_1378,In_1939);
xnor U630 (N_630,In_494,In_1962);
nand U631 (N_631,In_1788,In_778);
xor U632 (N_632,In_745,In_1683);
xnor U633 (N_633,In_1511,In_923);
xnor U634 (N_634,In_1927,In_880);
nand U635 (N_635,In_1291,In_405);
xnor U636 (N_636,In_1970,In_1630);
nand U637 (N_637,In_1576,In_1835);
or U638 (N_638,In_242,In_757);
and U639 (N_639,In_1739,In_1912);
nor U640 (N_640,In_1694,In_548);
nor U641 (N_641,In_810,In_1720);
nand U642 (N_642,In_312,In_875);
or U643 (N_643,In_362,In_704);
or U644 (N_644,In_1635,In_597);
nand U645 (N_645,In_1237,In_1085);
nor U646 (N_646,In_333,In_448);
nor U647 (N_647,In_118,In_1918);
nand U648 (N_648,In_994,In_655);
xor U649 (N_649,In_1004,In_44);
nor U650 (N_650,In_198,In_1943);
nor U651 (N_651,In_1209,In_963);
nand U652 (N_652,In_1799,In_1914);
nand U653 (N_653,In_1455,In_209);
xnor U654 (N_654,In_73,In_499);
or U655 (N_655,In_1400,In_427);
or U656 (N_656,In_1072,In_908);
xnor U657 (N_657,In_231,In_1897);
xnor U658 (N_658,In_385,In_1007);
xor U659 (N_659,In_1065,In_1512);
nand U660 (N_660,In_639,In_1501);
nand U661 (N_661,In_409,In_65);
nand U662 (N_662,In_1560,In_1842);
xor U663 (N_663,In_1490,In_311);
nand U664 (N_664,In_168,In_197);
and U665 (N_665,In_1573,In_1116);
or U666 (N_666,In_1599,In_1964);
nor U667 (N_667,In_1402,In_987);
or U668 (N_668,In_624,In_657);
xnor U669 (N_669,In_1166,In_151);
nand U670 (N_670,In_1159,In_1316);
nor U671 (N_671,In_1081,In_932);
and U672 (N_672,In_916,In_642);
and U673 (N_673,In_584,In_133);
or U674 (N_674,In_1284,In_524);
nor U675 (N_675,In_1629,In_541);
or U676 (N_676,In_1833,In_771);
xor U677 (N_677,In_60,In_1329);
nand U678 (N_678,In_971,In_258);
or U679 (N_679,In_1816,In_128);
and U680 (N_680,In_1697,In_1853);
or U681 (N_681,In_19,In_113);
xor U682 (N_682,In_1712,In_596);
or U683 (N_683,In_395,In_1592);
nor U684 (N_684,In_1551,In_2);
xor U685 (N_685,In_1196,In_32);
nor U686 (N_686,In_237,In_1281);
and U687 (N_687,In_1769,In_1777);
nand U688 (N_688,In_360,In_661);
xor U689 (N_689,In_1915,In_1781);
nand U690 (N_690,In_1641,In_1155);
and U691 (N_691,In_594,In_969);
nor U692 (N_692,In_47,In_399);
or U693 (N_693,In_1307,In_382);
nor U694 (N_694,In_1189,In_71);
nor U695 (N_695,In_1404,In_1780);
nor U696 (N_696,In_997,In_259);
or U697 (N_697,In_1506,In_954);
nor U698 (N_698,In_1445,In_459);
xor U699 (N_699,In_131,In_1259);
nor U700 (N_700,In_1360,In_1719);
xor U701 (N_701,In_514,In_124);
nand U702 (N_702,In_88,In_1120);
xor U703 (N_703,In_917,In_822);
or U704 (N_704,In_1095,In_1133);
xnor U705 (N_705,In_1637,In_609);
or U706 (N_706,In_393,In_225);
or U707 (N_707,In_1075,In_1380);
or U708 (N_708,In_1860,In_70);
nand U709 (N_709,In_683,In_1124);
nor U710 (N_710,In_481,In_796);
xnor U711 (N_711,In_1814,In_721);
nand U712 (N_712,In_419,In_1623);
xor U713 (N_713,In_1082,In_116);
and U714 (N_714,In_1163,In_956);
xnor U715 (N_715,In_1447,In_1737);
nor U716 (N_716,In_1659,In_266);
nor U717 (N_717,In_1212,In_787);
and U718 (N_718,In_1489,In_1517);
and U719 (N_719,In_871,In_41);
nor U720 (N_720,In_832,In_241);
nor U721 (N_721,In_1537,In_196);
and U722 (N_722,In_1158,In_1226);
and U723 (N_723,In_504,In_507);
and U724 (N_724,In_1636,In_226);
xnor U725 (N_725,In_1096,In_1477);
nor U726 (N_726,In_175,In_1523);
nor U727 (N_727,In_94,In_170);
and U728 (N_728,In_1068,In_1117);
and U729 (N_729,In_451,In_129);
and U730 (N_730,In_1969,In_685);
xor U731 (N_731,In_519,In_249);
nor U732 (N_732,In_1932,In_421);
xor U733 (N_733,In_1666,In_1049);
nor U734 (N_734,In_1923,In_256);
nor U735 (N_735,In_804,In_1572);
or U736 (N_736,In_1439,In_861);
or U737 (N_737,In_1926,In_288);
and U738 (N_738,In_165,In_132);
or U739 (N_739,In_1429,In_145);
and U740 (N_740,In_1991,In_711);
xor U741 (N_741,In_1559,In_558);
nand U742 (N_742,In_1515,In_130);
nor U743 (N_743,In_354,In_1767);
and U744 (N_744,In_888,In_106);
nor U745 (N_745,In_697,In_345);
xnor U746 (N_746,In_86,In_214);
and U747 (N_747,In_699,In_14);
or U748 (N_748,In_1173,In_496);
nor U749 (N_749,In_1,In_1770);
and U750 (N_750,In_310,In_1234);
or U751 (N_751,In_349,In_1850);
and U752 (N_752,In_876,In_1763);
and U753 (N_753,In_1982,In_193);
nor U754 (N_754,In_1527,In_460);
nor U755 (N_755,In_708,In_1191);
xor U756 (N_756,In_383,In_598);
nand U757 (N_757,In_1037,In_1421);
nand U758 (N_758,In_67,In_1677);
xnor U759 (N_759,In_600,In_547);
nand U760 (N_760,In_677,In_248);
or U761 (N_761,In_929,In_1046);
nand U762 (N_762,In_403,In_79);
or U763 (N_763,In_1010,In_1438);
nor U764 (N_764,In_1145,In_303);
or U765 (N_765,In_1137,In_1108);
nand U766 (N_766,In_64,In_1873);
or U767 (N_767,In_456,In_872);
xor U768 (N_768,In_970,In_1596);
and U769 (N_769,In_1193,In_715);
nand U770 (N_770,In_1916,In_1199);
nand U771 (N_771,In_1140,In_1563);
nand U772 (N_772,In_1292,In_188);
or U773 (N_773,In_966,In_1221);
or U774 (N_774,In_1453,In_1534);
and U775 (N_775,In_346,In_634);
nor U776 (N_776,In_1111,In_668);
nand U777 (N_777,In_1532,In_1825);
nand U778 (N_778,In_1328,In_1845);
or U779 (N_779,In_1016,In_1716);
nand U780 (N_780,In_341,In_1857);
nand U781 (N_781,In_1317,In_1283);
nor U782 (N_782,In_1294,In_314);
or U783 (N_783,In_1682,In_1904);
nor U784 (N_784,In_1263,In_1648);
nor U785 (N_785,In_1766,In_696);
or U786 (N_786,In_808,In_1580);
nand U787 (N_787,In_928,In_1526);
xnor U788 (N_788,In_533,In_985);
and U789 (N_789,In_1498,In_1183);
or U790 (N_790,In_490,In_1959);
xnor U791 (N_791,In_95,In_1411);
and U792 (N_792,In_1555,In_1951);
or U793 (N_793,In_1784,In_575);
nor U794 (N_794,In_1787,In_1507);
and U795 (N_795,In_1789,In_190);
nand U796 (N_796,In_1827,In_848);
nor U797 (N_797,In_682,In_392);
or U798 (N_798,In_189,In_1854);
and U799 (N_799,In_1067,In_1186);
nor U800 (N_800,In_1974,In_1887);
nor U801 (N_801,In_58,In_213);
and U802 (N_802,In_562,In_78);
or U803 (N_803,In_1748,In_309);
nor U804 (N_804,In_1327,In_280);
xnor U805 (N_805,In_767,In_265);
or U806 (N_806,In_563,In_1616);
nand U807 (N_807,In_973,In_1371);
xnor U808 (N_808,In_239,In_1319);
nand U809 (N_809,In_1315,In_1063);
xnor U810 (N_810,In_1844,In_1150);
nor U811 (N_811,In_302,In_1239);
or U812 (N_812,In_633,In_1409);
or U813 (N_813,In_1565,In_1840);
nand U814 (N_814,In_1408,In_232);
nand U815 (N_815,In_860,In_1652);
or U816 (N_816,In_1011,In_855);
and U817 (N_817,In_308,In_638);
or U818 (N_818,In_1180,In_1372);
xnor U819 (N_819,In_1132,In_1562);
xor U820 (N_820,In_922,In_404);
nor U821 (N_821,In_1407,In_1544);
xnor U822 (N_822,In_1107,In_1330);
and U823 (N_823,In_840,In_1268);
and U824 (N_824,In_612,In_785);
xnor U825 (N_825,In_1570,In_1006);
nand U826 (N_826,In_670,In_577);
nor U827 (N_827,In_1689,In_1241);
nor U828 (N_828,In_904,In_1699);
or U829 (N_829,In_390,In_1098);
or U830 (N_830,In_1446,In_1225);
xor U831 (N_831,In_621,In_1800);
nor U832 (N_832,In_1030,In_378);
nand U833 (N_833,In_1481,In_1856);
or U834 (N_834,In_989,In_1680);
xor U835 (N_835,In_1709,In_1997);
nor U836 (N_836,In_1884,In_684);
xnor U837 (N_837,In_1990,In_260);
nand U838 (N_838,In_1485,In_1509);
nand U839 (N_839,In_23,In_1240);
xor U840 (N_840,In_1583,In_1642);
or U841 (N_841,In_1624,In_1149);
nand U842 (N_842,In_694,In_556);
nand U843 (N_843,In_1903,In_1820);
nor U844 (N_844,In_666,In_446);
or U845 (N_845,In_930,In_847);
nand U846 (N_846,In_1381,In_898);
nand U847 (N_847,In_253,In_760);
nor U848 (N_848,In_1688,In_1933);
and U849 (N_849,In_1188,In_553);
and U850 (N_850,In_716,In_1147);
xor U851 (N_851,In_1602,In_1900);
nor U852 (N_852,In_444,In_899);
nand U853 (N_853,In_1220,In_1200);
nor U854 (N_854,In_1142,In_9);
and U855 (N_855,In_1773,In_1252);
nor U856 (N_856,In_1908,In_800);
xor U857 (N_857,In_1304,In_1568);
nand U858 (N_858,In_1632,In_592);
nand U859 (N_859,In_1866,In_827);
and U860 (N_860,In_690,In_1801);
nor U861 (N_861,In_961,In_1740);
nand U862 (N_862,In_372,In_703);
or U863 (N_863,In_1248,In_1084);
and U864 (N_864,In_1479,In_162);
nor U865 (N_865,In_1722,In_1734);
or U866 (N_866,In_329,In_1452);
and U867 (N_867,In_352,In_475);
and U868 (N_868,In_1771,In_1198);
nor U869 (N_869,In_1026,In_1348);
and U870 (N_870,In_1398,In_960);
xor U871 (N_871,In_192,In_1813);
or U872 (N_872,In_407,In_483);
or U873 (N_873,In_1779,In_1745);
or U874 (N_874,In_1433,In_844);
xnor U875 (N_875,In_774,In_1053);
nand U876 (N_876,In_1089,In_1867);
and U877 (N_877,In_626,In_933);
xnor U878 (N_878,In_1786,In_158);
xnor U879 (N_879,In_1018,In_115);
nand U880 (N_880,In_321,In_322);
xnor U881 (N_881,In_1336,In_194);
nor U882 (N_882,In_1487,In_1048);
and U883 (N_883,In_29,In_974);
or U884 (N_884,In_80,In_1530);
nand U885 (N_885,In_503,In_325);
nor U886 (N_886,In_210,In_1435);
and U887 (N_887,In_234,In_1488);
or U888 (N_888,In_1339,In_1403);
nor U889 (N_889,In_117,In_1342);
nand U890 (N_890,In_614,In_1417);
or U891 (N_891,In_486,In_1945);
nand U892 (N_892,In_1892,In_176);
nand U893 (N_893,In_1428,In_1710);
or U894 (N_894,In_566,In_1849);
nor U895 (N_895,In_1410,In_854);
and U896 (N_896,In_762,In_565);
xor U897 (N_897,In_1170,In_667);
nor U898 (N_898,In_1569,In_236);
xor U899 (N_899,In_1214,In_203);
xor U900 (N_900,In_691,In_1577);
nand U901 (N_901,In_1713,In_195);
and U902 (N_902,In_8,In_359);
nand U903 (N_903,In_1171,In_1782);
xnor U904 (N_904,In_1041,In_306);
and U905 (N_905,In_1809,In_134);
or U906 (N_906,In_376,In_1837);
nand U907 (N_907,In_348,In_1290);
or U908 (N_908,In_1954,In_636);
nor U909 (N_909,In_1492,In_838);
xnor U910 (N_910,In_1613,In_82);
nand U911 (N_911,In_1721,In_92);
or U912 (N_912,In_894,In_13);
or U913 (N_913,In_1738,In_1742);
or U914 (N_914,In_36,In_283);
or U915 (N_915,In_305,In_949);
and U916 (N_916,In_273,In_1736);
and U917 (N_917,In_413,In_1749);
nor U918 (N_918,In_601,In_528);
nor U919 (N_919,In_476,In_627);
and U920 (N_920,In_559,In_1370);
nor U921 (N_921,In_1424,In_1020);
xnor U922 (N_922,In_693,In_1244);
and U923 (N_923,In_965,In_1174);
xor U924 (N_924,In_59,In_1863);
nand U925 (N_925,In_1023,In_1730);
or U926 (N_926,In_386,In_1017);
or U927 (N_927,In_599,In_1977);
nand U928 (N_928,In_401,In_436);
nand U929 (N_929,In_1971,In_38);
or U930 (N_930,In_1953,In_761);
and U931 (N_931,In_995,In_1437);
and U932 (N_932,In_1911,In_746);
nand U933 (N_933,In_1972,In_720);
nand U934 (N_934,In_1473,In_1115);
or U935 (N_935,In_512,In_1005);
xnor U936 (N_936,In_509,In_864);
nor U937 (N_937,In_63,In_687);
and U938 (N_938,In_1913,In_307);
or U939 (N_939,In_863,In_1692);
xnor U940 (N_940,In_886,In_326);
nor U941 (N_941,In_906,In_135);
or U942 (N_942,In_576,In_529);
or U943 (N_943,In_1385,In_84);
xnor U944 (N_944,In_126,In_591);
nor U945 (N_945,In_1612,In_1729);
nor U946 (N_946,In_817,In_920);
and U947 (N_947,In_1528,In_799);
nand U948 (N_948,In_968,In_223);
or U949 (N_949,In_831,In_327);
nor U950 (N_950,In_52,In_764);
nor U951 (N_951,In_1389,In_1369);
and U952 (N_952,In_756,In_1413);
xnor U953 (N_953,In_416,In_1663);
and U954 (N_954,In_1533,In_1474);
nand U955 (N_955,In_1494,In_1634);
nand U956 (N_956,In_1985,In_1444);
and U957 (N_957,In_1762,In_892);
or U958 (N_958,In_1127,In_1247);
nand U959 (N_959,In_815,In_207);
nor U960 (N_960,In_535,In_1646);
or U961 (N_961,In_1743,In_713);
or U962 (N_962,In_1795,In_1843);
and U963 (N_963,In_301,In_878);
or U964 (N_964,In_1357,In_1571);
nor U965 (N_965,In_734,In_1957);
nor U966 (N_966,In_1144,In_1092);
nor U967 (N_967,In_795,In_101);
nor U968 (N_968,In_820,In_332);
or U969 (N_969,In_1087,In_520);
nor U970 (N_970,In_1152,In_1014);
xnor U971 (N_971,In_1693,In_921);
and U972 (N_972,In_1313,In_531);
nand U973 (N_973,In_500,In_42);
nor U974 (N_974,In_211,In_1060);
and U975 (N_975,In_297,In_1701);
or U976 (N_976,In_1222,In_1376);
nand U977 (N_977,In_1979,In_1519);
and U978 (N_978,In_1930,In_1566);
or U979 (N_979,In_1862,In_1941);
nor U980 (N_980,In_220,In_1662);
nand U981 (N_981,In_1335,In_1019);
nand U982 (N_982,In_1286,In_428);
and U983 (N_983,In_324,In_1461);
xnor U984 (N_984,In_1156,In_492);
xnor U985 (N_985,In_218,In_379);
xnor U986 (N_986,In_555,In_1732);
xnor U987 (N_987,In_1764,In_895);
and U988 (N_988,In_1015,In_1383);
or U989 (N_989,In_1001,In_1956);
nand U990 (N_990,In_539,In_798);
xor U991 (N_991,In_723,In_1040);
nor U992 (N_992,In_751,In_896);
nand U993 (N_993,In_1902,In_826);
and U994 (N_994,In_275,In_1083);
nand U995 (N_995,In_1233,In_443);
xor U996 (N_996,In_502,In_1388);
and U997 (N_997,In_289,In_45);
nand U998 (N_998,In_33,In_1008);
nand U999 (N_999,In_567,In_1726);
or U1000 (N_1000,In_1410,In_697);
and U1001 (N_1001,In_17,In_1718);
nand U1002 (N_1002,In_982,In_1296);
and U1003 (N_1003,In_1013,In_1288);
nand U1004 (N_1004,In_1537,In_921);
xnor U1005 (N_1005,In_1905,In_1436);
xnor U1006 (N_1006,In_60,In_1556);
xnor U1007 (N_1007,In_30,In_1298);
nor U1008 (N_1008,In_1934,In_906);
and U1009 (N_1009,In_386,In_1617);
or U1010 (N_1010,In_583,In_1044);
or U1011 (N_1011,In_1030,In_197);
nand U1012 (N_1012,In_455,In_636);
nor U1013 (N_1013,In_357,In_1684);
nor U1014 (N_1014,In_183,In_1980);
or U1015 (N_1015,In_510,In_1093);
xor U1016 (N_1016,In_740,In_98);
or U1017 (N_1017,In_387,In_376);
nand U1018 (N_1018,In_1038,In_1492);
xnor U1019 (N_1019,In_154,In_1556);
xor U1020 (N_1020,In_413,In_323);
nand U1021 (N_1021,In_1870,In_1093);
nand U1022 (N_1022,In_1343,In_49);
xor U1023 (N_1023,In_1257,In_617);
nor U1024 (N_1024,In_988,In_267);
xnor U1025 (N_1025,In_661,In_311);
or U1026 (N_1026,In_180,In_231);
nand U1027 (N_1027,In_1648,In_1111);
xnor U1028 (N_1028,In_737,In_609);
xnor U1029 (N_1029,In_1691,In_1878);
nand U1030 (N_1030,In_202,In_18);
nand U1031 (N_1031,In_397,In_1808);
nor U1032 (N_1032,In_1791,In_1826);
nand U1033 (N_1033,In_1667,In_374);
or U1034 (N_1034,In_392,In_242);
nand U1035 (N_1035,In_1413,In_367);
or U1036 (N_1036,In_1117,In_14);
nor U1037 (N_1037,In_1869,In_483);
and U1038 (N_1038,In_724,In_1367);
and U1039 (N_1039,In_103,In_1026);
xor U1040 (N_1040,In_1877,In_1360);
or U1041 (N_1041,In_326,In_848);
and U1042 (N_1042,In_1659,In_480);
nand U1043 (N_1043,In_10,In_461);
xnor U1044 (N_1044,In_1910,In_1149);
xnor U1045 (N_1045,In_1579,In_1961);
nand U1046 (N_1046,In_226,In_1477);
or U1047 (N_1047,In_579,In_1463);
and U1048 (N_1048,In_1876,In_305);
and U1049 (N_1049,In_627,In_400);
and U1050 (N_1050,In_819,In_166);
xnor U1051 (N_1051,In_1750,In_84);
or U1052 (N_1052,In_1548,In_1285);
nor U1053 (N_1053,In_1596,In_1278);
or U1054 (N_1054,In_1443,In_1467);
nand U1055 (N_1055,In_439,In_973);
nor U1056 (N_1056,In_1899,In_1932);
and U1057 (N_1057,In_1485,In_240);
or U1058 (N_1058,In_889,In_1756);
or U1059 (N_1059,In_1407,In_791);
or U1060 (N_1060,In_1856,In_1660);
or U1061 (N_1061,In_1569,In_453);
or U1062 (N_1062,In_459,In_872);
nand U1063 (N_1063,In_1957,In_1139);
nand U1064 (N_1064,In_994,In_1946);
and U1065 (N_1065,In_1702,In_1209);
and U1066 (N_1066,In_48,In_1512);
or U1067 (N_1067,In_325,In_379);
nand U1068 (N_1068,In_755,In_1717);
nand U1069 (N_1069,In_763,In_1184);
and U1070 (N_1070,In_64,In_1568);
xor U1071 (N_1071,In_895,In_1621);
nand U1072 (N_1072,In_1886,In_1589);
or U1073 (N_1073,In_52,In_1968);
xor U1074 (N_1074,In_365,In_713);
xor U1075 (N_1075,In_35,In_1055);
nand U1076 (N_1076,In_694,In_1545);
and U1077 (N_1077,In_994,In_1821);
nor U1078 (N_1078,In_999,In_1003);
and U1079 (N_1079,In_608,In_398);
and U1080 (N_1080,In_173,In_1915);
xor U1081 (N_1081,In_809,In_595);
nand U1082 (N_1082,In_63,In_617);
nor U1083 (N_1083,In_645,In_637);
and U1084 (N_1084,In_1115,In_1841);
or U1085 (N_1085,In_1688,In_1171);
and U1086 (N_1086,In_763,In_1723);
and U1087 (N_1087,In_811,In_325);
and U1088 (N_1088,In_971,In_1689);
and U1089 (N_1089,In_132,In_851);
and U1090 (N_1090,In_59,In_1013);
and U1091 (N_1091,In_596,In_1110);
nor U1092 (N_1092,In_1550,In_2);
nand U1093 (N_1093,In_326,In_1080);
nand U1094 (N_1094,In_807,In_875);
xor U1095 (N_1095,In_241,In_1507);
nor U1096 (N_1096,In_1919,In_1381);
or U1097 (N_1097,In_1158,In_1396);
and U1098 (N_1098,In_1733,In_849);
or U1099 (N_1099,In_120,In_1663);
or U1100 (N_1100,In_1875,In_1649);
and U1101 (N_1101,In_347,In_310);
xnor U1102 (N_1102,In_1448,In_1435);
nand U1103 (N_1103,In_1875,In_1611);
nor U1104 (N_1104,In_166,In_369);
xnor U1105 (N_1105,In_1189,In_63);
nor U1106 (N_1106,In_923,In_1320);
or U1107 (N_1107,In_629,In_52);
xnor U1108 (N_1108,In_857,In_1541);
and U1109 (N_1109,In_355,In_199);
and U1110 (N_1110,In_1408,In_1362);
nand U1111 (N_1111,In_159,In_1105);
and U1112 (N_1112,In_246,In_1820);
and U1113 (N_1113,In_261,In_1197);
nor U1114 (N_1114,In_1696,In_184);
or U1115 (N_1115,In_1375,In_120);
nand U1116 (N_1116,In_804,In_136);
nor U1117 (N_1117,In_724,In_1650);
nand U1118 (N_1118,In_1383,In_1755);
nand U1119 (N_1119,In_363,In_1132);
and U1120 (N_1120,In_791,In_1312);
xor U1121 (N_1121,In_926,In_1230);
xnor U1122 (N_1122,In_1636,In_1258);
nor U1123 (N_1123,In_1988,In_604);
nor U1124 (N_1124,In_176,In_1477);
nor U1125 (N_1125,In_55,In_722);
or U1126 (N_1126,In_1929,In_230);
or U1127 (N_1127,In_36,In_1068);
or U1128 (N_1128,In_1917,In_93);
and U1129 (N_1129,In_772,In_1685);
or U1130 (N_1130,In_655,In_630);
or U1131 (N_1131,In_787,In_1509);
and U1132 (N_1132,In_967,In_1213);
or U1133 (N_1133,In_1275,In_580);
xnor U1134 (N_1134,In_669,In_278);
xnor U1135 (N_1135,In_988,In_294);
nand U1136 (N_1136,In_165,In_1653);
or U1137 (N_1137,In_1780,In_1588);
or U1138 (N_1138,In_1773,In_690);
and U1139 (N_1139,In_1025,In_1718);
nand U1140 (N_1140,In_1623,In_1804);
nor U1141 (N_1141,In_1407,In_1768);
nand U1142 (N_1142,In_555,In_467);
nand U1143 (N_1143,In_392,In_1473);
or U1144 (N_1144,In_1422,In_834);
nand U1145 (N_1145,In_566,In_1430);
nor U1146 (N_1146,In_315,In_1633);
nand U1147 (N_1147,In_434,In_37);
nand U1148 (N_1148,In_1219,In_932);
xnor U1149 (N_1149,In_1731,In_159);
or U1150 (N_1150,In_784,In_1135);
xor U1151 (N_1151,In_1602,In_1370);
xor U1152 (N_1152,In_1947,In_117);
or U1153 (N_1153,In_385,In_84);
xor U1154 (N_1154,In_253,In_1098);
and U1155 (N_1155,In_1647,In_460);
nand U1156 (N_1156,In_725,In_701);
nor U1157 (N_1157,In_1077,In_189);
nor U1158 (N_1158,In_303,In_709);
nand U1159 (N_1159,In_72,In_932);
xor U1160 (N_1160,In_1642,In_259);
nand U1161 (N_1161,In_1929,In_314);
nor U1162 (N_1162,In_1242,In_1996);
or U1163 (N_1163,In_333,In_508);
or U1164 (N_1164,In_956,In_661);
or U1165 (N_1165,In_712,In_686);
nand U1166 (N_1166,In_1428,In_571);
or U1167 (N_1167,In_1141,In_742);
or U1168 (N_1168,In_1538,In_1284);
and U1169 (N_1169,In_1041,In_1967);
xnor U1170 (N_1170,In_1677,In_783);
xor U1171 (N_1171,In_969,In_1295);
and U1172 (N_1172,In_1744,In_104);
or U1173 (N_1173,In_967,In_963);
nand U1174 (N_1174,In_818,In_1713);
xor U1175 (N_1175,In_1611,In_230);
xnor U1176 (N_1176,In_1634,In_814);
and U1177 (N_1177,In_684,In_302);
and U1178 (N_1178,In_1520,In_736);
or U1179 (N_1179,In_1764,In_1664);
xor U1180 (N_1180,In_572,In_1652);
nor U1181 (N_1181,In_466,In_1574);
xor U1182 (N_1182,In_300,In_1648);
nor U1183 (N_1183,In_1518,In_869);
nor U1184 (N_1184,In_1061,In_2);
and U1185 (N_1185,In_936,In_17);
and U1186 (N_1186,In_1067,In_1507);
xnor U1187 (N_1187,In_1577,In_592);
xor U1188 (N_1188,In_824,In_1025);
and U1189 (N_1189,In_940,In_1828);
xnor U1190 (N_1190,In_1506,In_1666);
nor U1191 (N_1191,In_879,In_552);
or U1192 (N_1192,In_963,In_1633);
nor U1193 (N_1193,In_1277,In_472);
nand U1194 (N_1194,In_540,In_841);
or U1195 (N_1195,In_1886,In_272);
xnor U1196 (N_1196,In_1097,In_823);
and U1197 (N_1197,In_1805,In_332);
and U1198 (N_1198,In_1278,In_293);
nand U1199 (N_1199,In_1409,In_1162);
nand U1200 (N_1200,In_882,In_279);
or U1201 (N_1201,In_1267,In_1768);
xnor U1202 (N_1202,In_888,In_894);
nand U1203 (N_1203,In_548,In_1685);
nor U1204 (N_1204,In_49,In_467);
xor U1205 (N_1205,In_1671,In_713);
nor U1206 (N_1206,In_572,In_1835);
nand U1207 (N_1207,In_1445,In_121);
or U1208 (N_1208,In_1578,In_1782);
or U1209 (N_1209,In_606,In_342);
and U1210 (N_1210,In_1387,In_1573);
or U1211 (N_1211,In_1950,In_1260);
nand U1212 (N_1212,In_757,In_458);
nand U1213 (N_1213,In_1197,In_1661);
nand U1214 (N_1214,In_588,In_573);
and U1215 (N_1215,In_795,In_369);
and U1216 (N_1216,In_161,In_1431);
and U1217 (N_1217,In_1070,In_1397);
and U1218 (N_1218,In_1224,In_867);
and U1219 (N_1219,In_1990,In_207);
xnor U1220 (N_1220,In_573,In_1045);
or U1221 (N_1221,In_1714,In_1901);
or U1222 (N_1222,In_418,In_165);
nand U1223 (N_1223,In_1476,In_1014);
and U1224 (N_1224,In_205,In_1527);
and U1225 (N_1225,In_558,In_167);
nand U1226 (N_1226,In_1052,In_1259);
and U1227 (N_1227,In_16,In_553);
nand U1228 (N_1228,In_1409,In_1608);
xnor U1229 (N_1229,In_181,In_1633);
xor U1230 (N_1230,In_674,In_887);
nor U1231 (N_1231,In_1432,In_914);
nand U1232 (N_1232,In_673,In_680);
nor U1233 (N_1233,In_1891,In_872);
or U1234 (N_1234,In_1791,In_792);
xnor U1235 (N_1235,In_925,In_1888);
nand U1236 (N_1236,In_1805,In_1916);
or U1237 (N_1237,In_1402,In_1950);
nor U1238 (N_1238,In_594,In_503);
or U1239 (N_1239,In_1786,In_1589);
and U1240 (N_1240,In_1317,In_966);
nand U1241 (N_1241,In_1310,In_757);
xor U1242 (N_1242,In_1875,In_1551);
and U1243 (N_1243,In_1240,In_720);
and U1244 (N_1244,In_711,In_643);
nand U1245 (N_1245,In_765,In_743);
and U1246 (N_1246,In_614,In_698);
xor U1247 (N_1247,In_78,In_1023);
or U1248 (N_1248,In_445,In_423);
nor U1249 (N_1249,In_1657,In_585);
or U1250 (N_1250,In_707,In_389);
and U1251 (N_1251,In_1936,In_351);
xor U1252 (N_1252,In_804,In_1354);
nor U1253 (N_1253,In_706,In_993);
nor U1254 (N_1254,In_34,In_1251);
nand U1255 (N_1255,In_111,In_1114);
and U1256 (N_1256,In_908,In_730);
nor U1257 (N_1257,In_1110,In_932);
and U1258 (N_1258,In_530,In_176);
and U1259 (N_1259,In_1707,In_161);
and U1260 (N_1260,In_729,In_1095);
nand U1261 (N_1261,In_653,In_1379);
nor U1262 (N_1262,In_1773,In_1750);
nand U1263 (N_1263,In_753,In_1501);
and U1264 (N_1264,In_200,In_842);
nor U1265 (N_1265,In_1677,In_202);
nor U1266 (N_1266,In_1504,In_1737);
and U1267 (N_1267,In_1117,In_1730);
nor U1268 (N_1268,In_230,In_1968);
xor U1269 (N_1269,In_874,In_601);
nand U1270 (N_1270,In_1263,In_1784);
or U1271 (N_1271,In_1598,In_1210);
xor U1272 (N_1272,In_40,In_1210);
nor U1273 (N_1273,In_857,In_1741);
nand U1274 (N_1274,In_437,In_1339);
nand U1275 (N_1275,In_297,In_912);
or U1276 (N_1276,In_1069,In_1723);
nand U1277 (N_1277,In_894,In_326);
nor U1278 (N_1278,In_1382,In_1824);
nor U1279 (N_1279,In_781,In_360);
or U1280 (N_1280,In_74,In_651);
nor U1281 (N_1281,In_1279,In_317);
and U1282 (N_1282,In_1366,In_574);
and U1283 (N_1283,In_887,In_972);
and U1284 (N_1284,In_1797,In_757);
nand U1285 (N_1285,In_339,In_1983);
nor U1286 (N_1286,In_1122,In_938);
xnor U1287 (N_1287,In_596,In_78);
nor U1288 (N_1288,In_524,In_304);
or U1289 (N_1289,In_358,In_813);
and U1290 (N_1290,In_1962,In_1924);
nor U1291 (N_1291,In_1231,In_518);
nand U1292 (N_1292,In_313,In_273);
and U1293 (N_1293,In_1990,In_1786);
nand U1294 (N_1294,In_922,In_516);
xor U1295 (N_1295,In_703,In_1042);
and U1296 (N_1296,In_1855,In_928);
or U1297 (N_1297,In_1739,In_991);
nand U1298 (N_1298,In_679,In_528);
nand U1299 (N_1299,In_1905,In_1947);
or U1300 (N_1300,In_1797,In_767);
nand U1301 (N_1301,In_1959,In_1865);
or U1302 (N_1302,In_1860,In_498);
nor U1303 (N_1303,In_584,In_504);
or U1304 (N_1304,In_1554,In_1391);
or U1305 (N_1305,In_759,In_1794);
and U1306 (N_1306,In_1212,In_105);
nand U1307 (N_1307,In_426,In_861);
or U1308 (N_1308,In_1808,In_491);
nand U1309 (N_1309,In_1498,In_570);
or U1310 (N_1310,In_938,In_6);
nand U1311 (N_1311,In_1404,In_484);
or U1312 (N_1312,In_263,In_751);
nor U1313 (N_1313,In_601,In_357);
nand U1314 (N_1314,In_1437,In_1770);
nand U1315 (N_1315,In_1471,In_53);
nor U1316 (N_1316,In_1923,In_25);
nor U1317 (N_1317,In_1828,In_360);
xor U1318 (N_1318,In_501,In_1616);
xnor U1319 (N_1319,In_915,In_1900);
xor U1320 (N_1320,In_1490,In_1115);
or U1321 (N_1321,In_307,In_910);
or U1322 (N_1322,In_1525,In_710);
xor U1323 (N_1323,In_596,In_1778);
and U1324 (N_1324,In_1257,In_205);
xor U1325 (N_1325,In_584,In_995);
xnor U1326 (N_1326,In_281,In_1140);
or U1327 (N_1327,In_102,In_956);
nand U1328 (N_1328,In_1716,In_537);
and U1329 (N_1329,In_629,In_998);
nor U1330 (N_1330,In_1672,In_437);
xor U1331 (N_1331,In_1790,In_11);
and U1332 (N_1332,In_1187,In_1818);
xnor U1333 (N_1333,In_243,In_1941);
or U1334 (N_1334,In_1668,In_183);
nor U1335 (N_1335,In_1767,In_679);
nor U1336 (N_1336,In_1602,In_451);
and U1337 (N_1337,In_1249,In_933);
nand U1338 (N_1338,In_1832,In_1007);
nor U1339 (N_1339,In_1969,In_690);
nand U1340 (N_1340,In_436,In_1258);
nand U1341 (N_1341,In_1539,In_566);
nor U1342 (N_1342,In_1075,In_1711);
or U1343 (N_1343,In_109,In_1821);
xnor U1344 (N_1344,In_1113,In_1198);
nand U1345 (N_1345,In_473,In_521);
nor U1346 (N_1346,In_603,In_360);
or U1347 (N_1347,In_1961,In_1972);
xor U1348 (N_1348,In_173,In_1958);
nand U1349 (N_1349,In_619,In_1289);
or U1350 (N_1350,In_1114,In_1642);
and U1351 (N_1351,In_1598,In_1771);
or U1352 (N_1352,In_1863,In_1125);
and U1353 (N_1353,In_1970,In_1679);
nor U1354 (N_1354,In_1558,In_1662);
nand U1355 (N_1355,In_594,In_1328);
or U1356 (N_1356,In_113,In_323);
xor U1357 (N_1357,In_1566,In_631);
nor U1358 (N_1358,In_1906,In_1439);
and U1359 (N_1359,In_1870,In_1446);
or U1360 (N_1360,In_97,In_1760);
xor U1361 (N_1361,In_617,In_1593);
nor U1362 (N_1362,In_1201,In_444);
nand U1363 (N_1363,In_464,In_382);
and U1364 (N_1364,In_1,In_391);
or U1365 (N_1365,In_1458,In_571);
or U1366 (N_1366,In_608,In_0);
or U1367 (N_1367,In_827,In_1466);
or U1368 (N_1368,In_1616,In_1166);
nor U1369 (N_1369,In_1649,In_1930);
xor U1370 (N_1370,In_21,In_1611);
and U1371 (N_1371,In_122,In_356);
nand U1372 (N_1372,In_900,In_410);
xor U1373 (N_1373,In_781,In_870);
nor U1374 (N_1374,In_1798,In_1906);
nand U1375 (N_1375,In_1896,In_456);
xor U1376 (N_1376,In_603,In_942);
nor U1377 (N_1377,In_1178,In_1667);
nand U1378 (N_1378,In_799,In_322);
or U1379 (N_1379,In_549,In_1145);
nor U1380 (N_1380,In_1083,In_1293);
or U1381 (N_1381,In_1042,In_1690);
nor U1382 (N_1382,In_1748,In_813);
xor U1383 (N_1383,In_169,In_1936);
and U1384 (N_1384,In_1903,In_178);
xnor U1385 (N_1385,In_419,In_864);
xnor U1386 (N_1386,In_555,In_1212);
xor U1387 (N_1387,In_1650,In_1725);
nand U1388 (N_1388,In_1750,In_1633);
nor U1389 (N_1389,In_960,In_1496);
xor U1390 (N_1390,In_1821,In_1901);
xnor U1391 (N_1391,In_1540,In_621);
and U1392 (N_1392,In_1949,In_605);
nor U1393 (N_1393,In_437,In_1444);
and U1394 (N_1394,In_563,In_900);
and U1395 (N_1395,In_1924,In_1667);
or U1396 (N_1396,In_228,In_1768);
nand U1397 (N_1397,In_1723,In_1010);
xor U1398 (N_1398,In_76,In_1783);
nand U1399 (N_1399,In_1175,In_1481);
xor U1400 (N_1400,In_1963,In_996);
nand U1401 (N_1401,In_859,In_1222);
nor U1402 (N_1402,In_509,In_1042);
xor U1403 (N_1403,In_171,In_1742);
or U1404 (N_1404,In_303,In_848);
xor U1405 (N_1405,In_1828,In_627);
nand U1406 (N_1406,In_1813,In_918);
nand U1407 (N_1407,In_1905,In_779);
xor U1408 (N_1408,In_154,In_874);
xnor U1409 (N_1409,In_389,In_1583);
or U1410 (N_1410,In_1793,In_1393);
nor U1411 (N_1411,In_1260,In_1337);
nand U1412 (N_1412,In_362,In_457);
nand U1413 (N_1413,In_1594,In_714);
or U1414 (N_1414,In_613,In_233);
nand U1415 (N_1415,In_787,In_1794);
nor U1416 (N_1416,In_581,In_1434);
nor U1417 (N_1417,In_1623,In_296);
or U1418 (N_1418,In_942,In_1893);
or U1419 (N_1419,In_812,In_1667);
xor U1420 (N_1420,In_927,In_622);
or U1421 (N_1421,In_500,In_1647);
nand U1422 (N_1422,In_1412,In_691);
nand U1423 (N_1423,In_1007,In_919);
and U1424 (N_1424,In_1970,In_1545);
nor U1425 (N_1425,In_1568,In_1100);
or U1426 (N_1426,In_1517,In_1305);
nor U1427 (N_1427,In_855,In_404);
nor U1428 (N_1428,In_323,In_1837);
nand U1429 (N_1429,In_90,In_423);
nand U1430 (N_1430,In_1898,In_946);
xor U1431 (N_1431,In_1507,In_502);
xor U1432 (N_1432,In_1504,In_78);
and U1433 (N_1433,In_1439,In_1385);
and U1434 (N_1434,In_1943,In_954);
nand U1435 (N_1435,In_25,In_297);
xnor U1436 (N_1436,In_1857,In_326);
or U1437 (N_1437,In_323,In_1823);
xor U1438 (N_1438,In_317,In_1743);
and U1439 (N_1439,In_713,In_1351);
nand U1440 (N_1440,In_1186,In_1214);
nor U1441 (N_1441,In_1538,In_1856);
and U1442 (N_1442,In_1596,In_906);
or U1443 (N_1443,In_94,In_76);
nand U1444 (N_1444,In_998,In_1347);
or U1445 (N_1445,In_984,In_75);
and U1446 (N_1446,In_134,In_1752);
or U1447 (N_1447,In_1500,In_620);
or U1448 (N_1448,In_490,In_88);
nor U1449 (N_1449,In_1319,In_1961);
or U1450 (N_1450,In_1513,In_101);
xor U1451 (N_1451,In_1865,In_1453);
xor U1452 (N_1452,In_1812,In_1860);
xor U1453 (N_1453,In_965,In_1761);
and U1454 (N_1454,In_736,In_940);
or U1455 (N_1455,In_1832,In_1006);
xor U1456 (N_1456,In_865,In_212);
nand U1457 (N_1457,In_413,In_272);
xnor U1458 (N_1458,In_1700,In_1145);
or U1459 (N_1459,In_150,In_876);
or U1460 (N_1460,In_819,In_1876);
nor U1461 (N_1461,In_1764,In_1365);
nor U1462 (N_1462,In_14,In_1613);
and U1463 (N_1463,In_148,In_13);
nor U1464 (N_1464,In_303,In_409);
or U1465 (N_1465,In_1543,In_301);
nand U1466 (N_1466,In_874,In_1704);
nor U1467 (N_1467,In_275,In_91);
and U1468 (N_1468,In_707,In_416);
nand U1469 (N_1469,In_1269,In_1939);
xor U1470 (N_1470,In_551,In_1794);
or U1471 (N_1471,In_984,In_1921);
xor U1472 (N_1472,In_902,In_1226);
xor U1473 (N_1473,In_860,In_741);
nand U1474 (N_1474,In_68,In_1617);
xor U1475 (N_1475,In_1732,In_1108);
or U1476 (N_1476,In_1884,In_1752);
or U1477 (N_1477,In_1964,In_796);
nor U1478 (N_1478,In_1540,In_87);
nand U1479 (N_1479,In_1947,In_540);
and U1480 (N_1480,In_90,In_1639);
xor U1481 (N_1481,In_1834,In_1195);
and U1482 (N_1482,In_1783,In_1085);
or U1483 (N_1483,In_245,In_870);
nor U1484 (N_1484,In_65,In_1031);
nor U1485 (N_1485,In_1400,In_1119);
or U1486 (N_1486,In_199,In_1097);
and U1487 (N_1487,In_1059,In_1029);
or U1488 (N_1488,In_738,In_469);
nand U1489 (N_1489,In_1722,In_1078);
nand U1490 (N_1490,In_624,In_184);
or U1491 (N_1491,In_1492,In_1004);
xnor U1492 (N_1492,In_1047,In_1843);
nand U1493 (N_1493,In_717,In_683);
or U1494 (N_1494,In_316,In_1517);
xnor U1495 (N_1495,In_781,In_564);
or U1496 (N_1496,In_1389,In_958);
nand U1497 (N_1497,In_94,In_1387);
nor U1498 (N_1498,In_1382,In_754);
or U1499 (N_1499,In_412,In_812);
and U1500 (N_1500,In_1294,In_527);
nor U1501 (N_1501,In_1054,In_520);
and U1502 (N_1502,In_271,In_1500);
and U1503 (N_1503,In_40,In_1442);
nor U1504 (N_1504,In_1160,In_1981);
xor U1505 (N_1505,In_32,In_622);
xnor U1506 (N_1506,In_1295,In_1629);
or U1507 (N_1507,In_320,In_404);
nand U1508 (N_1508,In_1084,In_1390);
or U1509 (N_1509,In_1697,In_1407);
nand U1510 (N_1510,In_1929,In_946);
nand U1511 (N_1511,In_1185,In_1896);
nor U1512 (N_1512,In_480,In_297);
nand U1513 (N_1513,In_287,In_1107);
nand U1514 (N_1514,In_455,In_1054);
and U1515 (N_1515,In_325,In_666);
xor U1516 (N_1516,In_28,In_37);
nand U1517 (N_1517,In_380,In_1810);
nor U1518 (N_1518,In_418,In_1221);
nand U1519 (N_1519,In_1901,In_211);
and U1520 (N_1520,In_1431,In_290);
or U1521 (N_1521,In_300,In_844);
nor U1522 (N_1522,In_1590,In_1670);
and U1523 (N_1523,In_1056,In_1064);
xnor U1524 (N_1524,In_141,In_7);
and U1525 (N_1525,In_1302,In_1036);
xnor U1526 (N_1526,In_736,In_1733);
xor U1527 (N_1527,In_1124,In_823);
or U1528 (N_1528,In_711,In_199);
and U1529 (N_1529,In_1796,In_1276);
nor U1530 (N_1530,In_580,In_332);
or U1531 (N_1531,In_1388,In_985);
xor U1532 (N_1532,In_278,In_1395);
xnor U1533 (N_1533,In_1014,In_399);
or U1534 (N_1534,In_1453,In_1753);
or U1535 (N_1535,In_539,In_1181);
xnor U1536 (N_1536,In_1108,In_163);
nand U1537 (N_1537,In_1030,In_108);
or U1538 (N_1538,In_846,In_1872);
nand U1539 (N_1539,In_1913,In_1207);
nand U1540 (N_1540,In_1194,In_1643);
and U1541 (N_1541,In_618,In_289);
nor U1542 (N_1542,In_1411,In_1654);
nor U1543 (N_1543,In_1491,In_122);
and U1544 (N_1544,In_84,In_38);
or U1545 (N_1545,In_1603,In_79);
and U1546 (N_1546,In_229,In_674);
nand U1547 (N_1547,In_1823,In_187);
or U1548 (N_1548,In_791,In_1708);
nand U1549 (N_1549,In_1160,In_382);
or U1550 (N_1550,In_1313,In_1384);
and U1551 (N_1551,In_1505,In_1661);
xor U1552 (N_1552,In_237,In_1539);
or U1553 (N_1553,In_87,In_1565);
or U1554 (N_1554,In_714,In_729);
nand U1555 (N_1555,In_596,In_961);
nand U1556 (N_1556,In_1228,In_272);
and U1557 (N_1557,In_1650,In_1936);
xor U1558 (N_1558,In_185,In_59);
nor U1559 (N_1559,In_1730,In_1620);
nor U1560 (N_1560,In_130,In_377);
nand U1561 (N_1561,In_1602,In_1099);
nand U1562 (N_1562,In_1750,In_1267);
or U1563 (N_1563,In_1331,In_970);
or U1564 (N_1564,In_1276,In_77);
and U1565 (N_1565,In_487,In_376);
or U1566 (N_1566,In_916,In_1425);
nor U1567 (N_1567,In_1097,In_1334);
nor U1568 (N_1568,In_518,In_1429);
nor U1569 (N_1569,In_1309,In_947);
and U1570 (N_1570,In_1149,In_1095);
and U1571 (N_1571,In_1137,In_577);
nand U1572 (N_1572,In_1476,In_846);
xnor U1573 (N_1573,In_934,In_1345);
and U1574 (N_1574,In_1853,In_1060);
or U1575 (N_1575,In_1178,In_498);
or U1576 (N_1576,In_807,In_1504);
xor U1577 (N_1577,In_798,In_212);
and U1578 (N_1578,In_344,In_467);
or U1579 (N_1579,In_441,In_265);
and U1580 (N_1580,In_340,In_1127);
or U1581 (N_1581,In_927,In_368);
or U1582 (N_1582,In_1278,In_1806);
or U1583 (N_1583,In_352,In_1462);
or U1584 (N_1584,In_230,In_206);
nand U1585 (N_1585,In_192,In_98);
xnor U1586 (N_1586,In_805,In_1923);
nand U1587 (N_1587,In_434,In_826);
nor U1588 (N_1588,In_708,In_203);
or U1589 (N_1589,In_1097,In_1399);
nor U1590 (N_1590,In_302,In_976);
and U1591 (N_1591,In_845,In_1391);
or U1592 (N_1592,In_422,In_755);
xnor U1593 (N_1593,In_1323,In_548);
nor U1594 (N_1594,In_1037,In_1012);
or U1595 (N_1595,In_934,In_1809);
xnor U1596 (N_1596,In_563,In_1687);
and U1597 (N_1597,In_1871,In_872);
xnor U1598 (N_1598,In_120,In_1289);
nor U1599 (N_1599,In_628,In_146);
or U1600 (N_1600,In_155,In_1471);
xor U1601 (N_1601,In_718,In_355);
xor U1602 (N_1602,In_1633,In_1700);
nand U1603 (N_1603,In_634,In_1087);
xor U1604 (N_1604,In_1611,In_1921);
or U1605 (N_1605,In_237,In_405);
and U1606 (N_1606,In_430,In_1836);
nor U1607 (N_1607,In_1931,In_1343);
xor U1608 (N_1608,In_490,In_342);
xnor U1609 (N_1609,In_627,In_1313);
xor U1610 (N_1610,In_480,In_797);
nand U1611 (N_1611,In_1814,In_1909);
nand U1612 (N_1612,In_1147,In_1059);
nand U1613 (N_1613,In_971,In_1686);
xor U1614 (N_1614,In_1800,In_814);
or U1615 (N_1615,In_1420,In_1294);
nand U1616 (N_1616,In_1479,In_672);
or U1617 (N_1617,In_922,In_1219);
xnor U1618 (N_1618,In_1977,In_1291);
and U1619 (N_1619,In_1441,In_1594);
xnor U1620 (N_1620,In_1592,In_503);
or U1621 (N_1621,In_1753,In_1245);
nor U1622 (N_1622,In_979,In_1780);
and U1623 (N_1623,In_1639,In_569);
and U1624 (N_1624,In_581,In_1593);
or U1625 (N_1625,In_1937,In_1952);
xnor U1626 (N_1626,In_1356,In_916);
or U1627 (N_1627,In_1766,In_1345);
nor U1628 (N_1628,In_1939,In_975);
xor U1629 (N_1629,In_1134,In_996);
or U1630 (N_1630,In_587,In_1712);
nor U1631 (N_1631,In_1228,In_1198);
nor U1632 (N_1632,In_846,In_995);
or U1633 (N_1633,In_714,In_1895);
nand U1634 (N_1634,In_803,In_1938);
nand U1635 (N_1635,In_1754,In_1955);
and U1636 (N_1636,In_243,In_333);
or U1637 (N_1637,In_1882,In_1455);
and U1638 (N_1638,In_151,In_255);
xnor U1639 (N_1639,In_1557,In_93);
xor U1640 (N_1640,In_608,In_613);
and U1641 (N_1641,In_1399,In_1985);
nand U1642 (N_1642,In_1852,In_11);
xnor U1643 (N_1643,In_110,In_256);
or U1644 (N_1644,In_1083,In_1179);
or U1645 (N_1645,In_725,In_1923);
and U1646 (N_1646,In_423,In_1097);
nand U1647 (N_1647,In_1395,In_604);
nor U1648 (N_1648,In_1685,In_1005);
or U1649 (N_1649,In_180,In_1339);
nand U1650 (N_1650,In_186,In_1557);
and U1651 (N_1651,In_1571,In_259);
and U1652 (N_1652,In_1919,In_408);
and U1653 (N_1653,In_727,In_898);
or U1654 (N_1654,In_1417,In_825);
xnor U1655 (N_1655,In_33,In_857);
xnor U1656 (N_1656,In_1813,In_290);
xor U1657 (N_1657,In_1907,In_1319);
nor U1658 (N_1658,In_1535,In_937);
nor U1659 (N_1659,In_1746,In_1084);
nand U1660 (N_1660,In_1841,In_1730);
or U1661 (N_1661,In_797,In_438);
nand U1662 (N_1662,In_1250,In_1134);
xor U1663 (N_1663,In_1339,In_293);
xnor U1664 (N_1664,In_572,In_902);
xnor U1665 (N_1665,In_130,In_1419);
nand U1666 (N_1666,In_1774,In_1601);
xor U1667 (N_1667,In_1782,In_142);
nor U1668 (N_1668,In_1051,In_561);
nand U1669 (N_1669,In_1466,In_1159);
nand U1670 (N_1670,In_1145,In_1771);
and U1671 (N_1671,In_1157,In_863);
xnor U1672 (N_1672,In_386,In_373);
nor U1673 (N_1673,In_1296,In_1532);
nor U1674 (N_1674,In_1218,In_911);
nand U1675 (N_1675,In_364,In_1527);
xor U1676 (N_1676,In_1193,In_151);
and U1677 (N_1677,In_1752,In_1519);
nor U1678 (N_1678,In_1331,In_1203);
nor U1679 (N_1679,In_1378,In_1849);
xnor U1680 (N_1680,In_1364,In_1414);
nand U1681 (N_1681,In_484,In_958);
nand U1682 (N_1682,In_761,In_478);
and U1683 (N_1683,In_678,In_1912);
xnor U1684 (N_1684,In_641,In_1045);
and U1685 (N_1685,In_344,In_1055);
xnor U1686 (N_1686,In_1506,In_535);
nand U1687 (N_1687,In_1616,In_287);
nor U1688 (N_1688,In_228,In_319);
and U1689 (N_1689,In_1243,In_774);
nand U1690 (N_1690,In_1264,In_1150);
nor U1691 (N_1691,In_1567,In_596);
or U1692 (N_1692,In_1836,In_792);
and U1693 (N_1693,In_665,In_747);
nand U1694 (N_1694,In_800,In_1220);
and U1695 (N_1695,In_1763,In_616);
nor U1696 (N_1696,In_1777,In_1072);
and U1697 (N_1697,In_711,In_497);
or U1698 (N_1698,In_137,In_1459);
and U1699 (N_1699,In_540,In_1271);
nor U1700 (N_1700,In_896,In_1283);
nor U1701 (N_1701,In_709,In_889);
and U1702 (N_1702,In_961,In_1999);
xnor U1703 (N_1703,In_743,In_288);
or U1704 (N_1704,In_1235,In_886);
nor U1705 (N_1705,In_227,In_789);
and U1706 (N_1706,In_1515,In_303);
and U1707 (N_1707,In_729,In_1822);
xor U1708 (N_1708,In_834,In_804);
xor U1709 (N_1709,In_1519,In_311);
or U1710 (N_1710,In_679,In_6);
xnor U1711 (N_1711,In_436,In_398);
nand U1712 (N_1712,In_1348,In_530);
nand U1713 (N_1713,In_707,In_709);
nand U1714 (N_1714,In_1313,In_774);
nor U1715 (N_1715,In_1087,In_843);
and U1716 (N_1716,In_914,In_1002);
xnor U1717 (N_1717,In_733,In_926);
nand U1718 (N_1718,In_47,In_900);
xnor U1719 (N_1719,In_1125,In_432);
xor U1720 (N_1720,In_252,In_1378);
xor U1721 (N_1721,In_1390,In_1448);
or U1722 (N_1722,In_728,In_371);
nor U1723 (N_1723,In_612,In_1847);
nand U1724 (N_1724,In_1037,In_1228);
xnor U1725 (N_1725,In_215,In_1357);
nand U1726 (N_1726,In_134,In_611);
and U1727 (N_1727,In_377,In_1668);
nand U1728 (N_1728,In_593,In_255);
xnor U1729 (N_1729,In_1007,In_1015);
and U1730 (N_1730,In_1027,In_1953);
or U1731 (N_1731,In_1032,In_1416);
or U1732 (N_1732,In_939,In_1897);
nor U1733 (N_1733,In_1781,In_231);
xnor U1734 (N_1734,In_339,In_1086);
nor U1735 (N_1735,In_274,In_392);
nor U1736 (N_1736,In_577,In_151);
xnor U1737 (N_1737,In_1407,In_809);
xnor U1738 (N_1738,In_1643,In_1797);
and U1739 (N_1739,In_782,In_1260);
or U1740 (N_1740,In_1195,In_360);
or U1741 (N_1741,In_1832,In_690);
nor U1742 (N_1742,In_1991,In_1810);
nand U1743 (N_1743,In_166,In_1698);
xor U1744 (N_1744,In_1057,In_1913);
and U1745 (N_1745,In_1557,In_667);
nand U1746 (N_1746,In_1660,In_1294);
nand U1747 (N_1747,In_803,In_237);
nand U1748 (N_1748,In_1028,In_1814);
nor U1749 (N_1749,In_663,In_22);
nand U1750 (N_1750,In_1375,In_1263);
and U1751 (N_1751,In_373,In_450);
and U1752 (N_1752,In_161,In_1560);
xnor U1753 (N_1753,In_1914,In_1470);
and U1754 (N_1754,In_1679,In_1930);
nor U1755 (N_1755,In_1901,In_1166);
and U1756 (N_1756,In_876,In_1162);
xor U1757 (N_1757,In_907,In_346);
nor U1758 (N_1758,In_808,In_1514);
nor U1759 (N_1759,In_1718,In_697);
xor U1760 (N_1760,In_1709,In_1535);
nand U1761 (N_1761,In_640,In_1690);
xnor U1762 (N_1762,In_1209,In_1916);
xor U1763 (N_1763,In_1508,In_842);
nor U1764 (N_1764,In_1849,In_1677);
and U1765 (N_1765,In_949,In_1076);
nor U1766 (N_1766,In_1508,In_302);
and U1767 (N_1767,In_369,In_529);
nand U1768 (N_1768,In_1992,In_49);
nand U1769 (N_1769,In_208,In_513);
xnor U1770 (N_1770,In_1533,In_477);
xor U1771 (N_1771,In_516,In_1791);
xnor U1772 (N_1772,In_1388,In_127);
xnor U1773 (N_1773,In_281,In_960);
nor U1774 (N_1774,In_1509,In_33);
and U1775 (N_1775,In_1253,In_1706);
xor U1776 (N_1776,In_1827,In_1750);
or U1777 (N_1777,In_1912,In_755);
or U1778 (N_1778,In_341,In_394);
nor U1779 (N_1779,In_127,In_768);
or U1780 (N_1780,In_1414,In_1313);
nor U1781 (N_1781,In_1185,In_278);
or U1782 (N_1782,In_850,In_14);
xor U1783 (N_1783,In_1888,In_502);
nor U1784 (N_1784,In_1182,In_792);
or U1785 (N_1785,In_194,In_1084);
xor U1786 (N_1786,In_1127,In_1885);
nand U1787 (N_1787,In_227,In_1905);
nor U1788 (N_1788,In_738,In_746);
xor U1789 (N_1789,In_1731,In_1313);
or U1790 (N_1790,In_1237,In_150);
nor U1791 (N_1791,In_504,In_1598);
nand U1792 (N_1792,In_1111,In_564);
and U1793 (N_1793,In_209,In_971);
nand U1794 (N_1794,In_949,In_1011);
or U1795 (N_1795,In_1326,In_279);
xor U1796 (N_1796,In_878,In_1762);
nor U1797 (N_1797,In_1391,In_1575);
and U1798 (N_1798,In_901,In_838);
nand U1799 (N_1799,In_1640,In_50);
nor U1800 (N_1800,In_779,In_1618);
nand U1801 (N_1801,In_414,In_600);
or U1802 (N_1802,In_610,In_587);
nand U1803 (N_1803,In_360,In_64);
nor U1804 (N_1804,In_936,In_907);
nand U1805 (N_1805,In_1737,In_1084);
nand U1806 (N_1806,In_951,In_1264);
or U1807 (N_1807,In_14,In_825);
and U1808 (N_1808,In_224,In_1030);
nor U1809 (N_1809,In_1389,In_685);
xnor U1810 (N_1810,In_1134,In_1348);
xor U1811 (N_1811,In_1105,In_1983);
or U1812 (N_1812,In_1660,In_1546);
and U1813 (N_1813,In_191,In_1143);
nor U1814 (N_1814,In_1619,In_178);
xnor U1815 (N_1815,In_1345,In_1735);
nand U1816 (N_1816,In_1903,In_1044);
and U1817 (N_1817,In_274,In_1741);
and U1818 (N_1818,In_663,In_1272);
and U1819 (N_1819,In_110,In_920);
nor U1820 (N_1820,In_725,In_732);
and U1821 (N_1821,In_1309,In_695);
xor U1822 (N_1822,In_753,In_1533);
and U1823 (N_1823,In_884,In_1726);
xnor U1824 (N_1824,In_1510,In_1774);
or U1825 (N_1825,In_1040,In_588);
or U1826 (N_1826,In_77,In_966);
xor U1827 (N_1827,In_852,In_603);
xnor U1828 (N_1828,In_937,In_218);
nand U1829 (N_1829,In_1339,In_50);
nor U1830 (N_1830,In_400,In_490);
and U1831 (N_1831,In_1803,In_744);
and U1832 (N_1832,In_1133,In_853);
nand U1833 (N_1833,In_1620,In_75);
nand U1834 (N_1834,In_871,In_1605);
or U1835 (N_1835,In_1968,In_579);
nand U1836 (N_1836,In_1919,In_1663);
nor U1837 (N_1837,In_1950,In_1263);
or U1838 (N_1838,In_1437,In_911);
and U1839 (N_1839,In_1204,In_91);
or U1840 (N_1840,In_95,In_7);
or U1841 (N_1841,In_1304,In_620);
xnor U1842 (N_1842,In_1314,In_477);
xor U1843 (N_1843,In_148,In_1206);
or U1844 (N_1844,In_1585,In_223);
and U1845 (N_1845,In_1996,In_1487);
nor U1846 (N_1846,In_501,In_1769);
or U1847 (N_1847,In_295,In_1588);
nor U1848 (N_1848,In_986,In_1467);
and U1849 (N_1849,In_1573,In_1212);
or U1850 (N_1850,In_1465,In_1090);
nor U1851 (N_1851,In_1031,In_1767);
or U1852 (N_1852,In_1517,In_1910);
and U1853 (N_1853,In_1106,In_657);
nand U1854 (N_1854,In_1815,In_93);
and U1855 (N_1855,In_962,In_1576);
nand U1856 (N_1856,In_1606,In_1957);
and U1857 (N_1857,In_1049,In_134);
nor U1858 (N_1858,In_484,In_828);
xnor U1859 (N_1859,In_903,In_1912);
nor U1860 (N_1860,In_267,In_531);
nor U1861 (N_1861,In_1438,In_386);
and U1862 (N_1862,In_731,In_1234);
and U1863 (N_1863,In_1676,In_678);
xor U1864 (N_1864,In_1195,In_1337);
xnor U1865 (N_1865,In_1171,In_81);
nor U1866 (N_1866,In_430,In_1283);
nor U1867 (N_1867,In_209,In_272);
xnor U1868 (N_1868,In_1477,In_1803);
or U1869 (N_1869,In_778,In_1704);
nor U1870 (N_1870,In_1473,In_724);
or U1871 (N_1871,In_1684,In_966);
nand U1872 (N_1872,In_1365,In_1161);
xnor U1873 (N_1873,In_497,In_1239);
xor U1874 (N_1874,In_859,In_1630);
xnor U1875 (N_1875,In_1909,In_1346);
xor U1876 (N_1876,In_1097,In_436);
or U1877 (N_1877,In_1112,In_1491);
nand U1878 (N_1878,In_153,In_957);
nor U1879 (N_1879,In_1052,In_386);
or U1880 (N_1880,In_370,In_1461);
nand U1881 (N_1881,In_914,In_1706);
and U1882 (N_1882,In_1501,In_468);
xor U1883 (N_1883,In_186,In_1086);
xnor U1884 (N_1884,In_560,In_1147);
or U1885 (N_1885,In_1144,In_188);
and U1886 (N_1886,In_347,In_1797);
xnor U1887 (N_1887,In_875,In_1452);
nand U1888 (N_1888,In_1409,In_227);
nand U1889 (N_1889,In_27,In_1735);
xor U1890 (N_1890,In_1910,In_384);
xnor U1891 (N_1891,In_1271,In_840);
nor U1892 (N_1892,In_585,In_912);
xnor U1893 (N_1893,In_116,In_935);
and U1894 (N_1894,In_473,In_1077);
nor U1895 (N_1895,In_1619,In_1866);
or U1896 (N_1896,In_930,In_1146);
and U1897 (N_1897,In_1026,In_1714);
xor U1898 (N_1898,In_819,In_1486);
xnor U1899 (N_1899,In_1490,In_1689);
nor U1900 (N_1900,In_1412,In_1049);
nor U1901 (N_1901,In_502,In_499);
and U1902 (N_1902,In_1983,In_233);
and U1903 (N_1903,In_672,In_727);
or U1904 (N_1904,In_1373,In_1782);
or U1905 (N_1905,In_1001,In_1341);
or U1906 (N_1906,In_1987,In_1444);
xor U1907 (N_1907,In_1383,In_1864);
nor U1908 (N_1908,In_1703,In_237);
or U1909 (N_1909,In_1742,In_86);
or U1910 (N_1910,In_1103,In_845);
and U1911 (N_1911,In_1210,In_233);
xnor U1912 (N_1912,In_1068,In_1600);
nor U1913 (N_1913,In_762,In_1837);
nor U1914 (N_1914,In_258,In_1851);
or U1915 (N_1915,In_1119,In_67);
or U1916 (N_1916,In_1900,In_1920);
nand U1917 (N_1917,In_459,In_1008);
nand U1918 (N_1918,In_54,In_1330);
xnor U1919 (N_1919,In_1762,In_723);
xnor U1920 (N_1920,In_179,In_975);
or U1921 (N_1921,In_1859,In_1636);
or U1922 (N_1922,In_1574,In_1150);
nor U1923 (N_1923,In_1589,In_1535);
nor U1924 (N_1924,In_541,In_1401);
and U1925 (N_1925,In_904,In_1737);
nand U1926 (N_1926,In_53,In_1809);
and U1927 (N_1927,In_912,In_934);
xnor U1928 (N_1928,In_1423,In_1914);
and U1929 (N_1929,In_486,In_977);
nor U1930 (N_1930,In_1127,In_700);
and U1931 (N_1931,In_286,In_866);
xnor U1932 (N_1932,In_1296,In_799);
nand U1933 (N_1933,In_1086,In_1459);
nor U1934 (N_1934,In_956,In_212);
and U1935 (N_1935,In_190,In_45);
nor U1936 (N_1936,In_1791,In_845);
nor U1937 (N_1937,In_219,In_189);
nor U1938 (N_1938,In_1253,In_1442);
nand U1939 (N_1939,In_1014,In_110);
or U1940 (N_1940,In_129,In_602);
and U1941 (N_1941,In_736,In_1288);
or U1942 (N_1942,In_1484,In_1025);
xnor U1943 (N_1943,In_1141,In_566);
and U1944 (N_1944,In_621,In_1075);
nand U1945 (N_1945,In_748,In_897);
or U1946 (N_1946,In_1733,In_1164);
and U1947 (N_1947,In_1241,In_416);
or U1948 (N_1948,In_635,In_1440);
xnor U1949 (N_1949,In_111,In_849);
nor U1950 (N_1950,In_1771,In_143);
or U1951 (N_1951,In_1499,In_242);
xnor U1952 (N_1952,In_1819,In_1007);
nand U1953 (N_1953,In_375,In_1128);
xnor U1954 (N_1954,In_1048,In_1439);
or U1955 (N_1955,In_820,In_945);
nor U1956 (N_1956,In_1726,In_125);
and U1957 (N_1957,In_1693,In_945);
nor U1958 (N_1958,In_1040,In_1181);
or U1959 (N_1959,In_602,In_291);
and U1960 (N_1960,In_1391,In_1857);
nand U1961 (N_1961,In_1124,In_397);
nand U1962 (N_1962,In_467,In_1802);
and U1963 (N_1963,In_837,In_503);
and U1964 (N_1964,In_156,In_1466);
nand U1965 (N_1965,In_1831,In_1267);
nor U1966 (N_1966,In_1635,In_472);
nand U1967 (N_1967,In_1694,In_705);
nand U1968 (N_1968,In_1896,In_1160);
nand U1969 (N_1969,In_1376,In_1187);
nand U1970 (N_1970,In_304,In_765);
nand U1971 (N_1971,In_1230,In_1446);
xor U1972 (N_1972,In_1899,In_1577);
xnor U1973 (N_1973,In_1670,In_834);
nand U1974 (N_1974,In_1598,In_797);
and U1975 (N_1975,In_903,In_929);
or U1976 (N_1976,In_1043,In_1069);
or U1977 (N_1977,In_1425,In_480);
xor U1978 (N_1978,In_1057,In_1824);
nor U1979 (N_1979,In_1477,In_967);
or U1980 (N_1980,In_1409,In_469);
or U1981 (N_1981,In_811,In_796);
nand U1982 (N_1982,In_616,In_1489);
xnor U1983 (N_1983,In_974,In_1785);
xor U1984 (N_1984,In_441,In_29);
xnor U1985 (N_1985,In_668,In_1479);
or U1986 (N_1986,In_1426,In_1601);
nand U1987 (N_1987,In_1208,In_1968);
nor U1988 (N_1988,In_402,In_1701);
xnor U1989 (N_1989,In_286,In_575);
nor U1990 (N_1990,In_700,In_459);
xor U1991 (N_1991,In_584,In_1946);
nor U1992 (N_1992,In_1344,In_543);
nand U1993 (N_1993,In_1033,In_1880);
or U1994 (N_1994,In_333,In_1596);
xor U1995 (N_1995,In_777,In_105);
and U1996 (N_1996,In_1864,In_1543);
or U1997 (N_1997,In_1432,In_15);
or U1998 (N_1998,In_1836,In_379);
nand U1999 (N_1999,In_254,In_1470);
xor U2000 (N_2000,N_161,N_673);
nor U2001 (N_2001,N_822,N_1654);
xor U2002 (N_2002,N_215,N_1690);
and U2003 (N_2003,N_1463,N_921);
nor U2004 (N_2004,N_230,N_396);
and U2005 (N_2005,N_1960,N_1063);
xor U2006 (N_2006,N_712,N_1619);
or U2007 (N_2007,N_203,N_1649);
and U2008 (N_2008,N_34,N_1651);
or U2009 (N_2009,N_156,N_70);
and U2010 (N_2010,N_66,N_750);
nand U2011 (N_2011,N_113,N_647);
nand U2012 (N_2012,N_666,N_1020);
nor U2013 (N_2013,N_448,N_1609);
nand U2014 (N_2014,N_1676,N_931);
or U2015 (N_2015,N_843,N_1540);
xor U2016 (N_2016,N_1418,N_789);
or U2017 (N_2017,N_13,N_1867);
xor U2018 (N_2018,N_1689,N_516);
or U2019 (N_2019,N_1851,N_801);
xnor U2020 (N_2020,N_0,N_1744);
and U2021 (N_2021,N_414,N_407);
or U2022 (N_2022,N_766,N_233);
or U2023 (N_2023,N_102,N_1179);
xor U2024 (N_2024,N_106,N_1606);
and U2025 (N_2025,N_1094,N_255);
and U2026 (N_2026,N_470,N_1142);
or U2027 (N_2027,N_1764,N_1240);
nor U2028 (N_2028,N_1590,N_1201);
or U2029 (N_2029,N_389,N_1787);
nor U2030 (N_2030,N_648,N_1580);
or U2031 (N_2031,N_88,N_8);
xor U2032 (N_2032,N_1019,N_500);
and U2033 (N_2033,N_1781,N_1388);
nor U2034 (N_2034,N_1014,N_1930);
and U2035 (N_2035,N_744,N_593);
nor U2036 (N_2036,N_1322,N_68);
and U2037 (N_2037,N_1161,N_933);
and U2038 (N_2038,N_914,N_1384);
nor U2039 (N_2039,N_1193,N_1440);
nor U2040 (N_2040,N_915,N_355);
nand U2041 (N_2041,N_780,N_92);
xor U2042 (N_2042,N_1655,N_883);
or U2043 (N_2043,N_968,N_637);
xnor U2044 (N_2044,N_1489,N_1086);
nor U2045 (N_2045,N_1659,N_1458);
xnor U2046 (N_2046,N_511,N_1182);
or U2047 (N_2047,N_179,N_412);
nand U2048 (N_2048,N_1076,N_1919);
nand U2049 (N_2049,N_410,N_891);
xor U2050 (N_2050,N_84,N_1703);
nand U2051 (N_2051,N_54,N_1716);
nor U2052 (N_2052,N_1451,N_1591);
nor U2053 (N_2053,N_674,N_1173);
nand U2054 (N_2054,N_1373,N_1470);
or U2055 (N_2055,N_3,N_258);
nand U2056 (N_2056,N_164,N_1531);
nor U2057 (N_2057,N_746,N_1598);
nand U2058 (N_2058,N_524,N_1243);
nor U2059 (N_2059,N_786,N_1499);
nand U2060 (N_2060,N_1480,N_264);
nand U2061 (N_2061,N_18,N_1761);
nand U2062 (N_2062,N_755,N_52);
nand U2063 (N_2063,N_395,N_1359);
nor U2064 (N_2064,N_21,N_1868);
nand U2065 (N_2065,N_1383,N_1506);
and U2066 (N_2066,N_1091,N_241);
or U2067 (N_2067,N_216,N_1902);
nand U2068 (N_2068,N_28,N_144);
nor U2069 (N_2069,N_1328,N_297);
or U2070 (N_2070,N_979,N_1588);
and U2071 (N_2071,N_1239,N_783);
nor U2072 (N_2072,N_317,N_1369);
nor U2073 (N_2073,N_1999,N_808);
and U2074 (N_2074,N_739,N_279);
nor U2075 (N_2075,N_567,N_145);
and U2076 (N_2076,N_1184,N_1141);
nand U2077 (N_2077,N_1396,N_1560);
and U2078 (N_2078,N_1473,N_114);
nand U2079 (N_2079,N_25,N_486);
nor U2080 (N_2080,N_1840,N_1997);
nand U2081 (N_2081,N_603,N_1062);
and U2082 (N_2082,N_876,N_1414);
nand U2083 (N_2083,N_229,N_1773);
nand U2084 (N_2084,N_575,N_577);
and U2085 (N_2085,N_529,N_303);
or U2086 (N_2086,N_276,N_94);
or U2087 (N_2087,N_1083,N_1484);
nand U2088 (N_2088,N_26,N_1347);
nand U2089 (N_2089,N_227,N_1913);
xor U2090 (N_2090,N_492,N_23);
xor U2091 (N_2091,N_1077,N_731);
or U2092 (N_2092,N_613,N_1252);
and U2093 (N_2093,N_413,N_165);
nand U2094 (N_2094,N_199,N_1089);
and U2095 (N_2095,N_1578,N_526);
nand U2096 (N_2096,N_1981,N_313);
and U2097 (N_2097,N_627,N_865);
nor U2098 (N_2098,N_1650,N_1163);
nor U2099 (N_2099,N_589,N_1582);
xnor U2100 (N_2100,N_1188,N_827);
nand U2101 (N_2101,N_714,N_1080);
xor U2102 (N_2102,N_1425,N_523);
and U2103 (N_2103,N_964,N_1011);
nor U2104 (N_2104,N_1380,N_1284);
nand U2105 (N_2105,N_1259,N_247);
or U2106 (N_2106,N_1174,N_6);
and U2107 (N_2107,N_1250,N_960);
or U2108 (N_2108,N_1952,N_1266);
xor U2109 (N_2109,N_1305,N_1827);
xnor U2110 (N_2110,N_1576,N_820);
and U2111 (N_2111,N_1054,N_61);
nor U2112 (N_2112,N_1330,N_1510);
xor U2113 (N_2113,N_1992,N_1189);
xor U2114 (N_2114,N_1633,N_1724);
nand U2115 (N_2115,N_552,N_792);
or U2116 (N_2116,N_926,N_1736);
xnor U2117 (N_2117,N_244,N_969);
nand U2118 (N_2118,N_392,N_1427);
nor U2119 (N_2119,N_512,N_548);
xnor U2120 (N_2120,N_771,N_275);
or U2121 (N_2121,N_9,N_1759);
nand U2122 (N_2122,N_322,N_1137);
xor U2123 (N_2123,N_1381,N_4);
nand U2124 (N_2124,N_1241,N_1286);
xor U2125 (N_2125,N_759,N_1317);
or U2126 (N_2126,N_1820,N_1100);
and U2127 (N_2127,N_689,N_1394);
nand U2128 (N_2128,N_695,N_184);
xor U2129 (N_2129,N_80,N_812);
xor U2130 (N_2130,N_1740,N_310);
or U2131 (N_2131,N_400,N_1095);
or U2132 (N_2132,N_1911,N_1464);
and U2133 (N_2133,N_1107,N_1623);
or U2134 (N_2134,N_991,N_57);
or U2135 (N_2135,N_1798,N_1908);
and U2136 (N_2136,N_1399,N_483);
xor U2137 (N_2137,N_1012,N_1766);
xnor U2138 (N_2138,N_649,N_1669);
xor U2139 (N_2139,N_967,N_828);
or U2140 (N_2140,N_1513,N_453);
xnor U2141 (N_2141,N_842,N_433);
nor U2142 (N_2142,N_624,N_1356);
and U2143 (N_2143,N_565,N_851);
and U2144 (N_2144,N_955,N_710);
xor U2145 (N_2145,N_111,N_1434);
and U2146 (N_2146,N_560,N_368);
or U2147 (N_2147,N_195,N_1171);
xor U2148 (N_2148,N_840,N_1639);
or U2149 (N_2149,N_631,N_1708);
nand U2150 (N_2150,N_1392,N_1881);
nand U2151 (N_2151,N_667,N_1620);
nand U2152 (N_2152,N_862,N_1946);
nand U2153 (N_2153,N_1051,N_1162);
nand U2154 (N_2154,N_1036,N_1296);
xnor U2155 (N_2155,N_507,N_596);
and U2156 (N_2156,N_1310,N_315);
and U2157 (N_2157,N_265,N_119);
or U2158 (N_2158,N_653,N_974);
nand U2159 (N_2159,N_1,N_956);
and U2160 (N_2160,N_1558,N_605);
or U2161 (N_2161,N_1664,N_1420);
nor U2162 (N_2162,N_540,N_1785);
and U2163 (N_2163,N_234,N_1546);
xor U2164 (N_2164,N_1706,N_1979);
nor U2165 (N_2165,N_569,N_1196);
xnor U2166 (N_2166,N_334,N_1718);
or U2167 (N_2167,N_811,N_1497);
nor U2168 (N_2168,N_570,N_1772);
and U2169 (N_2169,N_617,N_450);
nand U2170 (N_2170,N_494,N_1121);
nand U2171 (N_2171,N_734,N_881);
nand U2172 (N_2172,N_616,N_1857);
and U2173 (N_2173,N_937,N_198);
and U2174 (N_2174,N_1353,N_1180);
nand U2175 (N_2175,N_1789,N_1301);
nor U2176 (N_2176,N_1613,N_882);
nor U2177 (N_2177,N_1711,N_939);
nor U2178 (N_2178,N_1068,N_1871);
xor U2179 (N_2179,N_925,N_1859);
nor U2180 (N_2180,N_623,N_296);
or U2181 (N_2181,N_1666,N_1684);
xor U2182 (N_2182,N_846,N_1360);
xnor U2183 (N_2183,N_573,N_259);
nand U2184 (N_2184,N_290,N_74);
xnor U2185 (N_2185,N_509,N_51);
nor U2186 (N_2186,N_1671,N_1276);
xnor U2187 (N_2187,N_1125,N_920);
nand U2188 (N_2188,N_411,N_541);
and U2189 (N_2189,N_1072,N_455);
nand U2190 (N_2190,N_168,N_778);
and U2191 (N_2191,N_1835,N_1526);
xnor U2192 (N_2192,N_350,N_1505);
and U2193 (N_2193,N_207,N_1528);
xor U2194 (N_2194,N_126,N_1983);
and U2195 (N_2195,N_940,N_711);
nand U2196 (N_2196,N_339,N_1437);
nor U2197 (N_2197,N_277,N_975);
xor U2198 (N_2198,N_534,N_323);
xnor U2199 (N_2199,N_1402,N_1251);
and U2200 (N_2200,N_1765,N_76);
nor U2201 (N_2201,N_127,N_1856);
xor U2202 (N_2202,N_238,N_736);
or U2203 (N_2203,N_42,N_1109);
or U2204 (N_2204,N_452,N_1774);
and U2205 (N_2205,N_1292,N_1041);
and U2206 (N_2206,N_1233,N_1204);
nor U2207 (N_2207,N_428,N_841);
xor U2208 (N_2208,N_1577,N_885);
xor U2209 (N_2209,N_1574,N_1514);
and U2210 (N_2210,N_604,N_489);
xnor U2211 (N_2211,N_340,N_1572);
nor U2212 (N_2212,N_679,N_629);
nand U2213 (N_2213,N_1273,N_397);
nand U2214 (N_2214,N_844,N_966);
and U2215 (N_2215,N_327,N_201);
and U2216 (N_2216,N_359,N_550);
nor U2217 (N_2217,N_1261,N_520);
nor U2218 (N_2218,N_154,N_1185);
nor U2219 (N_2219,N_1167,N_517);
and U2220 (N_2220,N_601,N_497);
nor U2221 (N_2221,N_740,N_1800);
and U2222 (N_2222,N_767,N_1426);
xnor U2223 (N_2223,N_1993,N_1541);
nand U2224 (N_2224,N_283,N_78);
nor U2225 (N_2225,N_430,N_1112);
nor U2226 (N_2226,N_136,N_1755);
nand U2227 (N_2227,N_902,N_1336);
xor U2228 (N_2228,N_930,N_1730);
xnor U2229 (N_2229,N_1575,N_1984);
nor U2230 (N_2230,N_923,N_1404);
xnor U2231 (N_2231,N_1763,N_1652);
xor U2232 (N_2232,N_1753,N_525);
xor U2233 (N_2233,N_157,N_1768);
nor U2234 (N_2234,N_929,N_1551);
nor U2235 (N_2235,N_1750,N_638);
xor U2236 (N_2236,N_549,N_1131);
xnor U2237 (N_2237,N_1677,N_562);
nand U2238 (N_2238,N_1726,N_476);
or U2239 (N_2239,N_950,N_46);
nand U2240 (N_2240,N_1046,N_1621);
nor U2241 (N_2241,N_1879,N_787);
or U2242 (N_2242,N_837,N_1562);
nor U2243 (N_2243,N_898,N_887);
nand U2244 (N_2244,N_943,N_1783);
nor U2245 (N_2245,N_141,N_139);
xor U2246 (N_2246,N_1692,N_1519);
nor U2247 (N_2247,N_532,N_335);
and U2248 (N_2248,N_219,N_1552);
xor U2249 (N_2249,N_1958,N_174);
or U2250 (N_2250,N_1874,N_1729);
or U2251 (N_2251,N_344,N_153);
xor U2252 (N_2252,N_886,N_1738);
nand U2253 (N_2253,N_218,N_374);
and U2254 (N_2254,N_652,N_703);
and U2255 (N_2255,N_1071,N_835);
or U2256 (N_2256,N_522,N_1969);
nand U2257 (N_2257,N_261,N_819);
and U2258 (N_2258,N_938,N_1568);
or U2259 (N_2259,N_1517,N_872);
nand U2260 (N_2260,N_1333,N_1891);
xor U2261 (N_2261,N_1005,N_1038);
and U2262 (N_2262,N_1342,N_375);
xnor U2263 (N_2263,N_1589,N_82);
or U2264 (N_2264,N_346,N_1625);
xor U2265 (N_2265,N_547,N_701);
xnor U2266 (N_2266,N_1731,N_1078);
and U2267 (N_2267,N_326,N_1878);
or U2268 (N_2268,N_704,N_228);
and U2269 (N_2269,N_1147,N_231);
xor U2270 (N_2270,N_650,N_361);
or U2271 (N_2271,N_1592,N_1127);
and U2272 (N_2272,N_607,N_436);
nand U2273 (N_2273,N_542,N_67);
nor U2274 (N_2274,N_100,N_1352);
xnor U2275 (N_2275,N_1246,N_980);
xnor U2276 (N_2276,N_1009,N_1377);
and U2277 (N_2277,N_1767,N_243);
xnor U2278 (N_2278,N_1483,N_1222);
xnor U2279 (N_2279,N_1114,N_875);
and U2280 (N_2280,N_1496,N_702);
nor U2281 (N_2281,N_528,N_566);
nor U2282 (N_2282,N_1618,N_1221);
nor U2283 (N_2283,N_867,N_1269);
or U2284 (N_2284,N_134,N_1897);
nand U2285 (N_2285,N_999,N_316);
and U2286 (N_2286,N_1447,N_1449);
nand U2287 (N_2287,N_636,N_1776);
nor U2288 (N_2288,N_1294,N_1421);
or U2289 (N_2289,N_1285,N_401);
and U2290 (N_2290,N_1031,N_1627);
or U2291 (N_2291,N_1644,N_705);
or U2292 (N_2292,N_1166,N_1103);
nand U2293 (N_2293,N_996,N_1900);
or U2294 (N_2294,N_274,N_663);
nand U2295 (N_2295,N_367,N_1130);
or U2296 (N_2296,N_1436,N_62);
nand U2297 (N_2297,N_1490,N_546);
or U2298 (N_2298,N_661,N_1796);
or U2299 (N_2299,N_1093,N_1733);
or U2300 (N_2300,N_1367,N_1925);
or U2301 (N_2301,N_1863,N_435);
nand U2302 (N_2302,N_1017,N_321);
nand U2303 (N_2303,N_1374,N_65);
xor U2304 (N_2304,N_376,N_1225);
xor U2305 (N_2305,N_572,N_850);
nand U2306 (N_2306,N_1281,N_681);
nand U2307 (N_2307,N_632,N_194);
nor U2308 (N_2308,N_1146,N_557);
and U2309 (N_2309,N_320,N_1673);
or U2310 (N_2310,N_32,N_1197);
or U2311 (N_2311,N_829,N_166);
or U2312 (N_2312,N_1110,N_1824);
nand U2313 (N_2313,N_437,N_1903);
nand U2314 (N_2314,N_912,N_963);
xor U2315 (N_2315,N_1614,N_479);
nand U2316 (N_2316,N_805,N_625);
nand U2317 (N_2317,N_879,N_558);
and U2318 (N_2318,N_694,N_1779);
or U2319 (N_2319,N_1465,N_587);
and U2320 (N_2320,N_237,N_1253);
nand U2321 (N_2321,N_1807,N_1350);
and U2322 (N_2322,N_1536,N_1140);
xor U2323 (N_2323,N_1550,N_15);
or U2324 (N_2324,N_1075,N_1971);
xor U2325 (N_2325,N_877,N_1721);
xor U2326 (N_2326,N_1423,N_1351);
and U2327 (N_2327,N_1149,N_1935);
and U2328 (N_2328,N_1719,N_976);
nand U2329 (N_2329,N_1088,N_609);
or U2330 (N_2330,N_1487,N_1052);
or U2331 (N_2331,N_1821,N_1670);
nand U2332 (N_2332,N_332,N_1608);
nor U2333 (N_2333,N_890,N_1509);
and U2334 (N_2334,N_588,N_793);
xor U2335 (N_2335,N_336,N_285);
or U2336 (N_2336,N_633,N_1694);
and U2337 (N_2337,N_1469,N_1454);
nand U2338 (N_2338,N_254,N_590);
xor U2339 (N_2339,N_490,N_471);
nor U2340 (N_2340,N_742,N_640);
nand U2341 (N_2341,N_845,N_798);
nor U2342 (N_2342,N_718,N_1699);
xnor U2343 (N_2343,N_722,N_348);
nand U2344 (N_2344,N_29,N_1525);
and U2345 (N_2345,N_852,N_1337);
or U2346 (N_2346,N_1954,N_1634);
or U2347 (N_2347,N_386,N_83);
nand U2348 (N_2348,N_725,N_903);
nor U2349 (N_2349,N_466,N_1211);
and U2350 (N_2350,N_1308,N_1688);
and U2351 (N_2351,N_16,N_459);
or U2352 (N_2352,N_698,N_1491);
nand U2353 (N_2353,N_1538,N_1371);
and U2354 (N_2354,N_193,N_1583);
or U2355 (N_2355,N_1771,N_382);
nand U2356 (N_2356,N_1283,N_1869);
or U2357 (N_2357,N_122,N_189);
or U2358 (N_2358,N_1455,N_574);
or U2359 (N_2359,N_1512,N_473);
and U2360 (N_2360,N_676,N_1823);
and U2361 (N_2361,N_257,N_1355);
nand U2362 (N_2362,N_1160,N_833);
or U2363 (N_2363,N_1151,N_138);
xnor U2364 (N_2364,N_752,N_1416);
and U2365 (N_2365,N_871,N_615);
nand U2366 (N_2366,N_1941,N_1864);
nor U2367 (N_2367,N_1963,N_1323);
or U2368 (N_2368,N_112,N_1450);
nor U2369 (N_2369,N_1500,N_343);
and U2370 (N_2370,N_142,N_416);
nor U2371 (N_2371,N_1135,N_543);
or U2372 (N_2372,N_1695,N_176);
and U2373 (N_2373,N_1516,N_85);
or U2374 (N_2374,N_170,N_670);
xnor U2375 (N_2375,N_472,N_1825);
xor U2376 (N_2376,N_1749,N_1111);
and U2377 (N_2377,N_1686,N_592);
nand U2378 (N_2378,N_753,N_642);
nand U2379 (N_2379,N_733,N_684);
or U2380 (N_2380,N_669,N_427);
or U2381 (N_2381,N_456,N_59);
nand U2382 (N_2382,N_1446,N_1048);
or U2383 (N_2383,N_1544,N_236);
and U2384 (N_2384,N_839,N_434);
and U2385 (N_2385,N_1290,N_803);
xnor U2386 (N_2386,N_1553,N_608);
nor U2387 (N_2387,N_656,N_1599);
or U2388 (N_2388,N_319,N_306);
or U2389 (N_2389,N_446,N_175);
nor U2390 (N_2390,N_1375,N_889);
xnor U2391 (N_2391,N_1013,N_458);
xor U2392 (N_2392,N_1808,N_1235);
nor U2393 (N_2393,N_1720,N_724);
or U2394 (N_2394,N_785,N_757);
nor U2395 (N_2395,N_985,N_571);
nor U2396 (N_2396,N_738,N_180);
or U2397 (N_2397,N_796,N_209);
and U2398 (N_2398,N_1084,N_618);
and U2399 (N_2399,N_1065,N_716);
nor U2400 (N_2400,N_1139,N_928);
or U2401 (N_2401,N_1680,N_1725);
nand U2402 (N_2402,N_847,N_1944);
xor U2403 (N_2403,N_1810,N_372);
nand U2404 (N_2404,N_1407,N_1674);
xnor U2405 (N_2405,N_700,N_1501);
and U2406 (N_2406,N_1442,N_1847);
and U2407 (N_2407,N_1543,N_1660);
nand U2408 (N_2408,N_1428,N_1372);
or U2409 (N_2409,N_1980,N_1136);
and U2410 (N_2410,N_1325,N_1461);
xor U2411 (N_2411,N_56,N_794);
nor U2412 (N_2412,N_393,N_1277);
nor U2413 (N_2413,N_905,N_1362);
nand U2414 (N_2414,N_385,N_556);
nor U2415 (N_2415,N_217,N_1630);
xnor U2416 (N_2416,N_1906,N_73);
nor U2417 (N_2417,N_1391,N_38);
and U2418 (N_2418,N_510,N_800);
nor U2419 (N_2419,N_1120,N_423);
nand U2420 (N_2420,N_720,N_868);
and U2421 (N_2421,N_432,N_748);
nor U2422 (N_2422,N_1557,N_672);
and U2423 (N_2423,N_1833,N_1203);
xor U2424 (N_2424,N_1929,N_1368);
and U2425 (N_2425,N_1029,N_1838);
xor U2426 (N_2426,N_1124,N_1662);
xnor U2427 (N_2427,N_1758,N_10);
xor U2428 (N_2428,N_1556,N_1010);
nand U2429 (N_2429,N_1482,N_260);
xnor U2430 (N_2430,N_539,N_72);
and U2431 (N_2431,N_1248,N_299);
xnor U2432 (N_2432,N_272,N_1811);
xnor U2433 (N_2433,N_1683,N_978);
or U2434 (N_2434,N_178,N_1486);
xnor U2435 (N_2435,N_662,N_1306);
nand U2436 (N_2436,N_474,N_1387);
nand U2437 (N_2437,N_1262,N_22);
and U2438 (N_2438,N_696,N_1218);
xnor U2439 (N_2439,N_438,N_946);
nor U2440 (N_2440,N_821,N_1382);
or U2441 (N_2441,N_1492,N_1965);
xnor U2442 (N_2442,N_418,N_1605);
nor U2443 (N_2443,N_977,N_559);
nor U2444 (N_2444,N_1132,N_1886);
xnor U2445 (N_2445,N_1631,N_1697);
xor U2446 (N_2446,N_1852,N_1249);
xnor U2447 (N_2447,N_150,N_641);
and U2448 (N_2448,N_1542,N_1311);
xnor U2449 (N_2449,N_1629,N_1494);
or U2450 (N_2450,N_1928,N_1788);
and U2451 (N_2451,N_916,N_1200);
nand U2452 (N_2452,N_1379,N_768);
nor U2453 (N_2453,N_50,N_1622);
nand U2454 (N_2454,N_1194,N_186);
nand U2455 (N_2455,N_719,N_1309);
or U2456 (N_2456,N_1028,N_1812);
and U2457 (N_2457,N_813,N_461);
and U2458 (N_2458,N_1702,N_1943);
or U2459 (N_2459,N_439,N_788);
nor U2460 (N_2460,N_1803,N_484);
and U2461 (N_2461,N_1433,N_1882);
xnor U2462 (N_2462,N_256,N_419);
xor U2463 (N_2463,N_44,N_1866);
nor U2464 (N_2464,N_1105,N_1667);
and U2465 (N_2465,N_1564,N_1939);
and U2466 (N_2466,N_858,N_1743);
nor U2467 (N_2467,N_1539,N_1157);
xor U2468 (N_2468,N_1467,N_622);
or U2469 (N_2469,N_1303,N_2);
or U2470 (N_2470,N_1060,N_1747);
or U2471 (N_2471,N_103,N_390);
nand U2472 (N_2472,N_727,N_505);
xnor U2473 (N_2473,N_657,N_330);
and U2474 (N_2474,N_1880,N_487);
and U2475 (N_2475,N_1593,N_1507);
xor U2476 (N_2476,N_1116,N_853);
or U2477 (N_2477,N_723,N_1393);
and U2478 (N_2478,N_519,N_1951);
nor U2479 (N_2479,N_140,N_1279);
xnor U2480 (N_2480,N_1242,N_990);
and U2481 (N_2481,N_398,N_1914);
xnor U2482 (N_2482,N_874,N_1527);
nor U2483 (N_2483,N_1186,N_1861);
nand U2484 (N_2484,N_1485,N_1476);
and U2485 (N_2485,N_1175,N_823);
and U2486 (N_2486,N_495,N_799);
nand U2487 (N_2487,N_1701,N_1280);
xnor U2488 (N_2488,N_1901,N_1366);
or U2489 (N_2489,N_1632,N_324);
xor U2490 (N_2490,N_1549,N_709);
nor U2491 (N_2491,N_36,N_1968);
or U2492 (N_2492,N_1797,N_1320);
nand U2493 (N_2493,N_1430,N_1475);
and U2494 (N_2494,N_445,N_287);
or U2495 (N_2495,N_40,N_708);
nand U2496 (N_2496,N_314,N_635);
xor U2497 (N_2497,N_774,N_1961);
or U2498 (N_2498,N_849,N_1950);
nand U2499 (N_2499,N_1271,N_212);
or U2500 (N_2500,N_163,N_266);
xor U2501 (N_2501,N_465,N_123);
nand U2502 (N_2502,N_688,N_1403);
or U2503 (N_2503,N_1601,N_579);
nor U2504 (N_2504,N_1524,N_441);
and U2505 (N_2505,N_1793,N_1904);
nor U2506 (N_2506,N_1734,N_364);
nand U2507 (N_2507,N_816,N_329);
and U2508 (N_2508,N_331,N_779);
or U2509 (N_2509,N_1287,N_1819);
nor U2510 (N_2510,N_564,N_544);
nor U2511 (N_2511,N_791,N_172);
and U2512 (N_2512,N_288,N_1799);
or U2513 (N_2513,N_1830,N_1926);
nor U2514 (N_2514,N_1164,N_451);
and U2515 (N_2515,N_1214,N_535);
or U2516 (N_2516,N_292,N_1899);
or U2517 (N_2517,N_869,N_148);
or U2518 (N_2518,N_1339,N_409);
nand U2519 (N_2519,N_686,N_1079);
nand U2520 (N_2520,N_832,N_294);
nand U2521 (N_2521,N_1818,N_1117);
and U2522 (N_2522,N_878,N_270);
nand U2523 (N_2523,N_1176,N_1663);
nand U2524 (N_2524,N_477,N_1389);
xnor U2525 (N_2525,N_406,N_131);
xor U2526 (N_2526,N_518,N_761);
nand U2527 (N_2527,N_1429,N_1612);
nor U2528 (N_2528,N_268,N_1700);
xor U2529 (N_2529,N_1212,N_1340);
nand U2530 (N_2530,N_1976,N_1782);
xnor U2531 (N_2531,N_1073,N_1587);
or U2532 (N_2532,N_1912,N_404);
nor U2533 (N_2533,N_463,N_919);
nor U2534 (N_2534,N_1033,N_1565);
nor U2535 (N_2535,N_130,N_1872);
nand U2536 (N_2536,N_1829,N_1099);
nor U2537 (N_2537,N_273,N_1682);
or U2538 (N_2538,N_89,N_659);
or U2539 (N_2539,N_1298,N_394);
nor U2540 (N_2540,N_1762,N_1534);
nand U2541 (N_2541,N_1635,N_1931);
or U2542 (N_2542,N_857,N_1408);
xnor U2543 (N_2543,N_870,N_942);
nor U2544 (N_2544,N_252,N_11);
or U2545 (N_2545,N_349,N_1217);
xnor U2546 (N_2546,N_894,N_553);
nand U2547 (N_2547,N_1836,N_69);
nand U2548 (N_2548,N_17,N_1144);
and U2549 (N_2549,N_224,N_1354);
nand U2550 (N_2550,N_1970,N_1945);
xor U2551 (N_2551,N_1626,N_462);
nand U2552 (N_2552,N_90,N_1230);
or U2553 (N_2553,N_1714,N_422);
or U2554 (N_2554,N_1386,N_1917);
nand U2555 (N_2555,N_619,N_415);
and U2556 (N_2556,N_863,N_478);
nand U2557 (N_2557,N_177,N_533);
and U2558 (N_2558,N_305,N_354);
and U2559 (N_2559,N_1806,N_530);
nand U2560 (N_2560,N_424,N_831);
and U2561 (N_2561,N_1304,N_1097);
and U2562 (N_2562,N_1705,N_1169);
and U2563 (N_2563,N_1410,N_1502);
xor U2564 (N_2564,N_1326,N_1295);
xnor U2565 (N_2565,N_1170,N_1918);
and U2566 (N_2566,N_949,N_1302);
nand U2567 (N_2567,N_171,N_884);
and U2568 (N_2568,N_55,N_1696);
xor U2569 (N_2569,N_795,N_1995);
nand U2570 (N_2570,N_347,N_536);
nand U2571 (N_2571,N_146,N_1846);
nand U2572 (N_2572,N_1045,N_1138);
nand U2573 (N_2573,N_1055,N_932);
or U2574 (N_2574,N_1792,N_769);
and U2575 (N_2575,N_1571,N_726);
xnor U2576 (N_2576,N_39,N_356);
and U2577 (N_2577,N_63,N_1845);
xor U2578 (N_2578,N_1967,N_1318);
or U2579 (N_2579,N_110,N_658);
or U2580 (N_2580,N_1101,N_1027);
nor U2581 (N_2581,N_992,N_1511);
or U2582 (N_2582,N_621,N_861);
nor U2583 (N_2583,N_781,N_208);
nor U2584 (N_2584,N_654,N_1113);
xnor U2585 (N_2585,N_31,N_1327);
xor U2586 (N_2586,N_1989,N_280);
xor U2587 (N_2587,N_600,N_1849);
and U2588 (N_2588,N_1554,N_1615);
xnor U2589 (N_2589,N_531,N_1358);
nor U2590 (N_2590,N_595,N_1916);
and U2591 (N_2591,N_1237,N_309);
or U2592 (N_2592,N_1828,N_682);
nor U2593 (N_2593,N_1229,N_1195);
or U2594 (N_2594,N_232,N_606);
or U2595 (N_2595,N_784,N_1831);
and U2596 (N_2596,N_1953,N_1521);
and U2597 (N_2597,N_12,N_1668);
nand U2598 (N_2598,N_1313,N_1289);
xor U2599 (N_2599,N_1348,N_697);
nand U2600 (N_2600,N_1611,N_1723);
nor U2601 (N_2601,N_1441,N_1123);
nor U2602 (N_2602,N_1642,N_1415);
nor U2603 (N_2603,N_1760,N_1223);
or U2604 (N_2604,N_1376,N_271);
nor U2605 (N_2605,N_71,N_1471);
xnor U2606 (N_2606,N_1198,N_1687);
xnor U2607 (N_2607,N_384,N_1457);
or U2608 (N_2608,N_953,N_924);
nand U2609 (N_2609,N_1254,N_910);
xnor U2610 (N_2610,N_1775,N_664);
or U2611 (N_2611,N_341,N_1982);
and U2612 (N_2612,N_1794,N_1887);
nand U2613 (N_2613,N_1804,N_1119);
and U2614 (N_2614,N_895,N_19);
nand U2615 (N_2615,N_169,N_1096);
nand U2616 (N_2616,N_187,N_1444);
xnor U2617 (N_2617,N_1523,N_496);
and U2618 (N_2618,N_1460,N_1949);
or U2619 (N_2619,N_1074,N_360);
or U2620 (N_2620,N_907,N_1535);
nand U2621 (N_2621,N_782,N_934);
or U2622 (N_2622,N_1843,N_1876);
and U2623 (N_2623,N_1624,N_854);
or U2624 (N_2624,N_1937,N_1927);
nor U2625 (N_2625,N_909,N_1640);
and U2626 (N_2626,N_660,N_1332);
nand U2627 (N_2627,N_1877,N_408);
nand U2628 (N_2628,N_1022,N_381);
or U2629 (N_2629,N_1335,N_1602);
xor U2630 (N_2630,N_1938,N_190);
nand U2631 (N_2631,N_634,N_1058);
nand U2632 (N_2632,N_947,N_683);
or U2633 (N_2633,N_124,N_1067);
and U2634 (N_2634,N_901,N_502);
or U2635 (N_2635,N_120,N_289);
and U2636 (N_2636,N_578,N_1658);
nand U2637 (N_2637,N_1047,N_644);
nand U2638 (N_2638,N_1924,N_250);
and U2639 (N_2639,N_152,N_1059);
nand U2640 (N_2640,N_584,N_48);
xor U2641 (N_2641,N_927,N_1448);
nor U2642 (N_2642,N_1893,N_253);
and U2643 (N_2643,N_1648,N_371);
nor U2644 (N_2644,N_1637,N_773);
nor U2645 (N_2645,N_873,N_1190);
xor U2646 (N_2646,N_1737,N_1584);
xor U2647 (N_2647,N_325,N_643);
nand U2648 (N_2648,N_690,N_747);
nor U2649 (N_2649,N_365,N_391);
or U2650 (N_2650,N_1518,N_1988);
nor U2651 (N_2651,N_1940,N_137);
and U2652 (N_2652,N_1754,N_1977);
or U2653 (N_2653,N_680,N_630);
or U2654 (N_2654,N_1152,N_1567);
or U2655 (N_2655,N_1712,N_896);
xnor U2656 (N_2656,N_221,N_35);
xor U2657 (N_2657,N_1357,N_855);
or U2658 (N_2658,N_192,N_1003);
nor U2659 (N_2659,N_1474,N_1090);
and U2660 (N_2660,N_1300,N_1258);
xnor U2661 (N_2661,N_917,N_1270);
nand U2662 (N_2662,N_1936,N_1921);
xor U2663 (N_2663,N_838,N_1638);
or U2664 (N_2664,N_1986,N_506);
nor U2665 (N_2665,N_1363,N_758);
xnor U2666 (N_2666,N_214,N_1907);
nand U2667 (N_2667,N_143,N_1234);
nor U2668 (N_2668,N_225,N_797);
or U2669 (N_2669,N_467,N_514);
xor U2670 (N_2670,N_1975,N_1777);
and U2671 (N_2671,N_307,N_1870);
xnor U2672 (N_2672,N_442,N_1905);
and U2673 (N_2673,N_580,N_1349);
and U2674 (N_2674,N_1616,N_1238);
or U2675 (N_2675,N_101,N_1641);
xor U2676 (N_2676,N_1452,N_599);
or U2677 (N_2677,N_188,N_1035);
nand U2678 (N_2678,N_586,N_685);
nor U2679 (N_2679,N_989,N_1839);
and U2680 (N_2680,N_191,N_155);
xor U2681 (N_2681,N_267,N_1841);
nand U2682 (N_2682,N_460,N_1555);
nor U2683 (N_2683,N_729,N_728);
or U2684 (N_2684,N_1272,N_713);
or U2685 (N_2685,N_1922,N_918);
nor U2686 (N_2686,N_269,N_1257);
or U2687 (N_2687,N_1600,N_687);
xnor U2688 (N_2688,N_815,N_53);
or U2689 (N_2689,N_1443,N_1991);
xor U2690 (N_2690,N_1098,N_1962);
nor U2691 (N_2691,N_183,N_1331);
or U2692 (N_2692,N_1888,N_262);
xor U2693 (N_2693,N_922,N_1156);
xor U2694 (N_2694,N_772,N_1070);
xor U2695 (N_2695,N_1532,N_1573);
nor U2696 (N_2696,N_856,N_1192);
xnor U2697 (N_2697,N_504,N_1653);
or U2698 (N_2698,N_1268,N_1603);
xor U2699 (N_2699,N_1741,N_1685);
xnor U2700 (N_2700,N_1586,N_417);
and U2701 (N_2701,N_1972,N_133);
or U2702 (N_2702,N_481,N_402);
nand U2703 (N_2703,N_1974,N_7);
nor U2704 (N_2704,N_485,N_913);
or U2705 (N_2705,N_1329,N_1092);
xor U2706 (N_2706,N_420,N_1128);
or U2707 (N_2707,N_561,N_735);
and U2708 (N_2708,N_1232,N_1748);
or U2709 (N_2709,N_555,N_302);
and U2710 (N_2710,N_1693,N_1263);
xnor U2711 (N_2711,N_298,N_1008);
nand U2712 (N_2712,N_447,N_1216);
nand U2713 (N_2713,N_1909,N_1481);
and U2714 (N_2714,N_1424,N_99);
nor U2715 (N_2715,N_1202,N_545);
nor U2716 (N_2716,N_1681,N_1814);
and U2717 (N_2717,N_538,N_1081);
or U2718 (N_2718,N_1274,N_749);
xnor U2719 (N_2719,N_936,N_185);
nand U2720 (N_2720,N_1129,N_91);
or U2721 (N_2721,N_1049,N_239);
nand U2722 (N_2722,N_1032,N_981);
or U2723 (N_2723,N_1915,N_1264);
and U2724 (N_2724,N_508,N_197);
or U2725 (N_2725,N_1154,N_1964);
or U2726 (N_2726,N_223,N_1226);
xor U2727 (N_2727,N_1529,N_1037);
nor U2728 (N_2728,N_1236,N_1145);
and U2729 (N_2729,N_378,N_970);
and U2730 (N_2730,N_665,N_97);
xor U2731 (N_2731,N_1873,N_205);
nand U2732 (N_2732,N_1115,N_117);
and U2733 (N_2733,N_1409,N_1401);
or U2734 (N_2734,N_1411,N_959);
nor U2735 (N_2735,N_1044,N_776);
or U2736 (N_2736,N_1207,N_1875);
or U2737 (N_2737,N_1021,N_213);
nand U2738 (N_2738,N_45,N_1594);
or U2739 (N_2739,N_1122,N_1646);
nand U2740 (N_2740,N_1150,N_1778);
or U2741 (N_2741,N_1459,N_1817);
nor U2742 (N_2742,N_318,N_454);
or U2743 (N_2743,N_1439,N_1570);
or U2744 (N_2744,N_1215,N_125);
and U2745 (N_2745,N_972,N_1678);
nor U2746 (N_2746,N_1344,N_668);
xor U2747 (N_2747,N_948,N_1533);
nor U2748 (N_2748,N_1069,N_1334);
and U2749 (N_2749,N_328,N_1739);
nand U2750 (N_2750,N_312,N_1865);
nor U2751 (N_2751,N_814,N_1213);
nor U2752 (N_2752,N_173,N_1260);
nand U2753 (N_2753,N_282,N_1061);
and U2754 (N_2754,N_551,N_1957);
and U2755 (N_2755,N_107,N_1645);
nand U2756 (N_2756,N_1400,N_1102);
xor U2757 (N_2757,N_818,N_443);
nand U2758 (N_2758,N_240,N_762);
nand U2759 (N_2759,N_1848,N_1040);
xnor U2760 (N_2760,N_1343,N_1610);
or U2761 (N_2761,N_431,N_475);
and U2762 (N_2762,N_1030,N_181);
and U2763 (N_2763,N_848,N_362);
xnor U2764 (N_2764,N_1438,N_1985);
nor U2765 (N_2765,N_1002,N_1199);
xnor U2766 (N_2766,N_311,N_30);
or U2767 (N_2767,N_892,N_333);
nor U2768 (N_2768,N_1826,N_1732);
and U2769 (N_2769,N_1822,N_482);
and U2770 (N_2770,N_1884,N_692);
nand U2771 (N_2771,N_286,N_1628);
nand U2772 (N_2772,N_242,N_860);
xnor U2773 (N_2773,N_345,N_1883);
or U2774 (N_2774,N_1698,N_162);
nand U2775 (N_2775,N_741,N_211);
or U2776 (N_2776,N_488,N_1607);
and U2777 (N_2777,N_200,N_988);
xor U2778 (N_2778,N_1106,N_1324);
or U2779 (N_2779,N_958,N_58);
nor U2780 (N_2780,N_79,N_1082);
or U2781 (N_2781,N_1126,N_1026);
and U2782 (N_2782,N_1370,N_1206);
or U2783 (N_2783,N_691,N_941);
and U2784 (N_2784,N_1177,N_830);
xor U2785 (N_2785,N_1210,N_491);
or U2786 (N_2786,N_1933,N_1710);
nor U2787 (N_2787,N_204,N_1431);
or U2788 (N_2788,N_1338,N_1488);
and U2789 (N_2789,N_1291,N_1006);
nor U2790 (N_2790,N_1345,N_775);
or U2791 (N_2791,N_965,N_47);
and U2792 (N_2792,N_1104,N_995);
xor U2793 (N_2793,N_1453,N_388);
and U2794 (N_2794,N_1756,N_291);
or U2795 (N_2795,N_1220,N_1432);
nand U2796 (N_2796,N_1990,N_984);
or U2797 (N_2797,N_352,N_1656);
or U2798 (N_2798,N_897,N_944);
nor U2799 (N_2799,N_993,N_576);
nand U2800 (N_2800,N_675,N_1000);
or U2801 (N_2801,N_1148,N_1837);
and U2802 (N_2802,N_1717,N_1178);
nand U2803 (N_2803,N_1043,N_1001);
and U2804 (N_2804,N_1503,N_1314);
or U2805 (N_2805,N_1548,N_128);
and U2806 (N_2806,N_278,N_1636);
and U2807 (N_2807,N_1537,N_1053);
and U2808 (N_2808,N_935,N_521);
xnor U2809 (N_2809,N_1361,N_1208);
nor U2810 (N_2810,N_1709,N_904);
xnor U2811 (N_2811,N_1784,N_1854);
and U2812 (N_2812,N_1050,N_1495);
and U2813 (N_2813,N_301,N_1722);
or U2814 (N_2814,N_468,N_1024);
and U2815 (N_2815,N_358,N_866);
nor U2816 (N_2816,N_263,N_908);
nand U2817 (N_2817,N_1158,N_1412);
and U2818 (N_2818,N_1769,N_646);
and U2819 (N_2819,N_1691,N_585);
and U2820 (N_2820,N_1155,N_300);
or U2821 (N_2821,N_817,N_383);
xnor U2822 (N_2822,N_763,N_1462);
and U2823 (N_2823,N_1751,N_1405);
or U2824 (N_2824,N_825,N_1889);
nor U2825 (N_2825,N_1498,N_864);
and U2826 (N_2826,N_1947,N_597);
nor U2827 (N_2827,N_1617,N_982);
and U2828 (N_2828,N_602,N_1809);
nand U2829 (N_2829,N_1064,N_1923);
and U2830 (N_2830,N_809,N_824);
nand U2831 (N_2831,N_1023,N_1996);
xnor U2832 (N_2832,N_693,N_1813);
xnor U2833 (N_2833,N_1267,N_1597);
nand U2834 (N_2834,N_806,N_43);
or U2835 (N_2835,N_1942,N_1244);
xor U2836 (N_2836,N_1585,N_27);
or U2837 (N_2837,N_1219,N_581);
nor U2838 (N_2838,N_671,N_1134);
and U2839 (N_2839,N_880,N_1920);
xor U2840 (N_2840,N_370,N_1715);
xnor U2841 (N_2841,N_1315,N_834);
nor U2842 (N_2842,N_1862,N_81);
nand U2843 (N_2843,N_1850,N_1834);
xor U2844 (N_2844,N_293,N_1227);
xor U2845 (N_2845,N_899,N_730);
nand U2846 (N_2846,N_598,N_754);
and U2847 (N_2847,N_611,N_994);
nand U2848 (N_2848,N_353,N_464);
or U2849 (N_2849,N_1665,N_1647);
and U2850 (N_2850,N_1209,N_1932);
nand U2851 (N_2851,N_1057,N_1275);
nor U2852 (N_2852,N_5,N_129);
nor U2853 (N_2853,N_1735,N_1752);
or U2854 (N_2854,N_1245,N_1816);
nor U2855 (N_2855,N_75,N_699);
nor U2856 (N_2856,N_1770,N_1395);
nor U2857 (N_2857,N_49,N_501);
xnor U2858 (N_2858,N_337,N_86);
or U2859 (N_2859,N_1885,N_1445);
nor U2860 (N_2860,N_1479,N_449);
or U2861 (N_2861,N_1547,N_610);
or U2862 (N_2862,N_1346,N_1435);
xnor U2863 (N_2863,N_1472,N_206);
nor U2864 (N_2864,N_1456,N_998);
or U2865 (N_2865,N_1018,N_121);
nor U2866 (N_2866,N_226,N_1312);
and U2867 (N_2867,N_338,N_612);
nor U2868 (N_2868,N_1417,N_1378);
xnor U2869 (N_2869,N_1398,N_1973);
xor U2870 (N_2870,N_678,N_888);
and U2871 (N_2871,N_1802,N_60);
or U2872 (N_2872,N_1278,N_513);
xnor U2873 (N_2873,N_246,N_1530);
or U2874 (N_2874,N_1745,N_1955);
or U2875 (N_2875,N_802,N_1934);
nand U2876 (N_2876,N_1746,N_764);
xor U2877 (N_2877,N_1742,N_639);
nor U2878 (N_2878,N_804,N_1228);
xor U2879 (N_2879,N_41,N_281);
nand U2880 (N_2880,N_1780,N_132);
or U2881 (N_2881,N_1832,N_469);
nor U2882 (N_2882,N_732,N_1508);
nand U2883 (N_2883,N_1133,N_655);
xnor U2884 (N_2884,N_1515,N_1522);
and U2885 (N_2885,N_202,N_1108);
nand U2886 (N_2886,N_1795,N_743);
xor U2887 (N_2887,N_1466,N_425);
xor U2888 (N_2888,N_760,N_1085);
nand U2889 (N_2889,N_20,N_1890);
nor U2890 (N_2890,N_906,N_591);
nand U2891 (N_2891,N_96,N_64);
xnor U2892 (N_2892,N_1419,N_33);
or U2893 (N_2893,N_1790,N_568);
or U2894 (N_2894,N_1118,N_440);
nor U2895 (N_2895,N_756,N_1657);
nor U2896 (N_2896,N_1520,N_554);
nand U2897 (N_2897,N_426,N_810);
nand U2898 (N_2898,N_377,N_1039);
nor U2899 (N_2899,N_135,N_1007);
nand U2900 (N_2900,N_1896,N_620);
and U2901 (N_2901,N_1894,N_1791);
or U2902 (N_2902,N_1056,N_1704);
and U2903 (N_2903,N_1168,N_1801);
and U2904 (N_2904,N_1319,N_444);
nand U2905 (N_2905,N_745,N_1288);
or U2906 (N_2906,N_342,N_628);
nor U2907 (N_2907,N_1728,N_770);
nand U2908 (N_2908,N_24,N_357);
nor U2909 (N_2909,N_158,N_403);
or U2910 (N_2910,N_1643,N_457);
nor U2911 (N_2911,N_304,N_429);
nor U2912 (N_2912,N_108,N_945);
xor U2913 (N_2913,N_582,N_1581);
or U2914 (N_2914,N_1406,N_366);
or U2915 (N_2915,N_1966,N_1231);
nor U2916 (N_2916,N_807,N_98);
or U2917 (N_2917,N_1390,N_147);
xnor U2918 (N_2918,N_1016,N_1321);
nand U2919 (N_2919,N_1165,N_1596);
and U2920 (N_2920,N_1265,N_363);
xnor U2921 (N_2921,N_997,N_1895);
or U2922 (N_2922,N_1559,N_1898);
nor U2923 (N_2923,N_1842,N_1307);
xnor U2924 (N_2924,N_1563,N_715);
nand U2925 (N_2925,N_1579,N_1143);
and U2926 (N_2926,N_379,N_1892);
and U2927 (N_2927,N_706,N_151);
xnor U2928 (N_2928,N_1595,N_1365);
nor U2929 (N_2929,N_182,N_765);
and U2930 (N_2930,N_498,N_1858);
xnor U2931 (N_2931,N_677,N_104);
nor U2932 (N_2932,N_1034,N_1959);
nor U2933 (N_2933,N_405,N_737);
nand U2934 (N_2934,N_961,N_1661);
xor U2935 (N_2935,N_1707,N_1205);
and U2936 (N_2936,N_645,N_421);
and U2937 (N_2937,N_503,N_87);
and U2938 (N_2938,N_220,N_1994);
or U2939 (N_2939,N_1282,N_1757);
xor U2940 (N_2940,N_351,N_387);
nand U2941 (N_2941,N_1910,N_721);
and U2942 (N_2942,N_1948,N_1478);
and U2943 (N_2943,N_614,N_95);
or U2944 (N_2944,N_1860,N_1815);
and U2945 (N_2945,N_118,N_159);
or U2946 (N_2946,N_196,N_836);
or U2947 (N_2947,N_251,N_1978);
and U2948 (N_2948,N_954,N_957);
and U2949 (N_2949,N_1672,N_1015);
nand U2950 (N_2950,N_1675,N_1855);
xor U2951 (N_2951,N_1561,N_1566);
nand U2952 (N_2952,N_1422,N_399);
or U2953 (N_2953,N_651,N_717);
and U2954 (N_2954,N_1805,N_499);
xor U2955 (N_2955,N_563,N_1853);
nor U2956 (N_2956,N_284,N_1224);
or U2957 (N_2957,N_826,N_1679);
nor U2958 (N_2958,N_167,N_1191);
and U2959 (N_2959,N_1604,N_480);
or U2960 (N_2960,N_248,N_583);
xor U2961 (N_2961,N_1956,N_537);
nor U2962 (N_2962,N_369,N_1172);
xor U2963 (N_2963,N_983,N_1493);
nor U2964 (N_2964,N_116,N_893);
or U2965 (N_2965,N_37,N_707);
and U2966 (N_2966,N_527,N_962);
nor U2967 (N_2967,N_987,N_1341);
nand U2968 (N_2968,N_1299,N_900);
xnor U2969 (N_2969,N_1247,N_626);
xnor U2970 (N_2970,N_295,N_1468);
nor U2971 (N_2971,N_115,N_515);
and U2972 (N_2972,N_1181,N_1297);
nand U2973 (N_2973,N_1004,N_1256);
xor U2974 (N_2974,N_777,N_245);
and U2975 (N_2975,N_93,N_308);
and U2976 (N_2976,N_951,N_751);
and U2977 (N_2977,N_380,N_973);
and U2978 (N_2978,N_210,N_971);
xnor U2979 (N_2979,N_1087,N_1727);
nand U2980 (N_2980,N_1545,N_1042);
and U2981 (N_2981,N_911,N_109);
and U2982 (N_2982,N_986,N_249);
xor U2983 (N_2983,N_1786,N_790);
or U2984 (N_2984,N_594,N_493);
nor U2985 (N_2985,N_1569,N_1187);
and U2986 (N_2986,N_1477,N_160);
nand U2987 (N_2987,N_1504,N_952);
or U2988 (N_2988,N_235,N_1397);
xnor U2989 (N_2989,N_1293,N_105);
xnor U2990 (N_2990,N_1998,N_1385);
or U2991 (N_2991,N_149,N_1987);
or U2992 (N_2992,N_859,N_77);
nand U2993 (N_2993,N_1255,N_1025);
nor U2994 (N_2994,N_1413,N_1153);
and U2995 (N_2995,N_373,N_1066);
xnor U2996 (N_2996,N_1713,N_1159);
nand U2997 (N_2997,N_1316,N_1844);
and U2998 (N_2998,N_14,N_222);
nand U2999 (N_2999,N_1364,N_1183);
and U3000 (N_3000,N_655,N_1839);
nor U3001 (N_3001,N_1849,N_1624);
nor U3002 (N_3002,N_1877,N_1045);
nor U3003 (N_3003,N_1216,N_1305);
or U3004 (N_3004,N_714,N_1379);
nor U3005 (N_3005,N_1544,N_982);
xnor U3006 (N_3006,N_160,N_1446);
xnor U3007 (N_3007,N_1425,N_340);
xor U3008 (N_3008,N_76,N_1321);
nor U3009 (N_3009,N_561,N_904);
nand U3010 (N_3010,N_1903,N_533);
nand U3011 (N_3011,N_1526,N_886);
or U3012 (N_3012,N_1589,N_59);
xor U3013 (N_3013,N_397,N_1546);
or U3014 (N_3014,N_1277,N_1458);
or U3015 (N_3015,N_1884,N_161);
and U3016 (N_3016,N_1377,N_1488);
nand U3017 (N_3017,N_291,N_889);
xor U3018 (N_3018,N_1698,N_1234);
nor U3019 (N_3019,N_1576,N_1584);
and U3020 (N_3020,N_1886,N_836);
nand U3021 (N_3021,N_705,N_649);
or U3022 (N_3022,N_1470,N_607);
or U3023 (N_3023,N_1990,N_1662);
xor U3024 (N_3024,N_1568,N_594);
nor U3025 (N_3025,N_1578,N_1427);
and U3026 (N_3026,N_1601,N_586);
nand U3027 (N_3027,N_1984,N_201);
or U3028 (N_3028,N_1075,N_1158);
nor U3029 (N_3029,N_1146,N_76);
nand U3030 (N_3030,N_46,N_133);
nor U3031 (N_3031,N_175,N_1361);
xnor U3032 (N_3032,N_1806,N_1065);
nor U3033 (N_3033,N_791,N_1937);
nand U3034 (N_3034,N_1775,N_1344);
nand U3035 (N_3035,N_561,N_401);
xnor U3036 (N_3036,N_1304,N_1011);
xnor U3037 (N_3037,N_1173,N_1611);
and U3038 (N_3038,N_1767,N_1074);
nor U3039 (N_3039,N_326,N_113);
and U3040 (N_3040,N_1532,N_1743);
nor U3041 (N_3041,N_133,N_1486);
and U3042 (N_3042,N_817,N_1772);
xnor U3043 (N_3043,N_690,N_1137);
or U3044 (N_3044,N_1591,N_851);
xor U3045 (N_3045,N_1708,N_1976);
or U3046 (N_3046,N_814,N_1980);
nand U3047 (N_3047,N_1152,N_657);
or U3048 (N_3048,N_1121,N_567);
or U3049 (N_3049,N_1177,N_968);
nand U3050 (N_3050,N_465,N_1658);
xnor U3051 (N_3051,N_552,N_124);
and U3052 (N_3052,N_21,N_556);
or U3053 (N_3053,N_291,N_1366);
nor U3054 (N_3054,N_616,N_943);
and U3055 (N_3055,N_1081,N_1111);
and U3056 (N_3056,N_543,N_792);
nand U3057 (N_3057,N_846,N_165);
or U3058 (N_3058,N_1714,N_1955);
nor U3059 (N_3059,N_1632,N_1755);
nand U3060 (N_3060,N_1079,N_1382);
nand U3061 (N_3061,N_986,N_707);
nand U3062 (N_3062,N_998,N_1590);
nand U3063 (N_3063,N_1511,N_106);
nand U3064 (N_3064,N_1089,N_827);
nand U3065 (N_3065,N_451,N_153);
and U3066 (N_3066,N_757,N_100);
xor U3067 (N_3067,N_1459,N_33);
xor U3068 (N_3068,N_880,N_1782);
or U3069 (N_3069,N_201,N_576);
or U3070 (N_3070,N_782,N_1488);
xnor U3071 (N_3071,N_1312,N_1755);
nand U3072 (N_3072,N_1354,N_1945);
and U3073 (N_3073,N_1622,N_345);
nor U3074 (N_3074,N_1631,N_582);
or U3075 (N_3075,N_193,N_274);
nand U3076 (N_3076,N_1318,N_1904);
nand U3077 (N_3077,N_429,N_1388);
nor U3078 (N_3078,N_1407,N_718);
xnor U3079 (N_3079,N_1770,N_242);
nand U3080 (N_3080,N_1228,N_1337);
xor U3081 (N_3081,N_0,N_1086);
nand U3082 (N_3082,N_882,N_430);
or U3083 (N_3083,N_1662,N_1351);
or U3084 (N_3084,N_1862,N_297);
xnor U3085 (N_3085,N_1092,N_635);
or U3086 (N_3086,N_617,N_747);
xor U3087 (N_3087,N_371,N_1504);
nand U3088 (N_3088,N_1262,N_1215);
xnor U3089 (N_3089,N_1723,N_677);
and U3090 (N_3090,N_1389,N_200);
and U3091 (N_3091,N_1070,N_1973);
xor U3092 (N_3092,N_1642,N_1197);
or U3093 (N_3093,N_1183,N_1693);
or U3094 (N_3094,N_1099,N_1383);
xnor U3095 (N_3095,N_1141,N_511);
nor U3096 (N_3096,N_1174,N_1741);
or U3097 (N_3097,N_1526,N_1090);
xnor U3098 (N_3098,N_752,N_448);
nor U3099 (N_3099,N_434,N_582);
and U3100 (N_3100,N_1112,N_190);
nor U3101 (N_3101,N_629,N_214);
nand U3102 (N_3102,N_434,N_838);
xor U3103 (N_3103,N_757,N_1737);
nand U3104 (N_3104,N_1424,N_1165);
xor U3105 (N_3105,N_945,N_1515);
nand U3106 (N_3106,N_1741,N_60);
or U3107 (N_3107,N_399,N_704);
nand U3108 (N_3108,N_975,N_289);
nand U3109 (N_3109,N_1436,N_968);
nand U3110 (N_3110,N_648,N_1935);
xnor U3111 (N_3111,N_329,N_1574);
and U3112 (N_3112,N_1044,N_907);
xnor U3113 (N_3113,N_1065,N_786);
xor U3114 (N_3114,N_663,N_829);
nor U3115 (N_3115,N_1921,N_416);
xnor U3116 (N_3116,N_1099,N_1263);
or U3117 (N_3117,N_210,N_1154);
and U3118 (N_3118,N_1003,N_169);
or U3119 (N_3119,N_1812,N_608);
nand U3120 (N_3120,N_1803,N_591);
xor U3121 (N_3121,N_1033,N_913);
xnor U3122 (N_3122,N_1923,N_243);
nor U3123 (N_3123,N_531,N_510);
nor U3124 (N_3124,N_1603,N_1604);
xnor U3125 (N_3125,N_833,N_390);
nor U3126 (N_3126,N_803,N_519);
nand U3127 (N_3127,N_62,N_1655);
or U3128 (N_3128,N_350,N_1498);
or U3129 (N_3129,N_1820,N_456);
nor U3130 (N_3130,N_755,N_681);
nor U3131 (N_3131,N_1846,N_1189);
and U3132 (N_3132,N_1062,N_905);
nand U3133 (N_3133,N_1829,N_1904);
and U3134 (N_3134,N_161,N_1881);
nor U3135 (N_3135,N_535,N_1616);
nand U3136 (N_3136,N_1113,N_530);
and U3137 (N_3137,N_1297,N_199);
nand U3138 (N_3138,N_1389,N_1494);
nor U3139 (N_3139,N_356,N_525);
nand U3140 (N_3140,N_1900,N_1049);
or U3141 (N_3141,N_817,N_1295);
xor U3142 (N_3142,N_730,N_451);
nand U3143 (N_3143,N_1818,N_1973);
nand U3144 (N_3144,N_363,N_796);
or U3145 (N_3145,N_1363,N_1720);
xor U3146 (N_3146,N_1296,N_1403);
nor U3147 (N_3147,N_122,N_539);
and U3148 (N_3148,N_1484,N_227);
and U3149 (N_3149,N_1061,N_873);
and U3150 (N_3150,N_1295,N_1922);
nand U3151 (N_3151,N_1255,N_420);
nor U3152 (N_3152,N_1427,N_960);
nor U3153 (N_3153,N_1846,N_766);
xnor U3154 (N_3154,N_1432,N_863);
and U3155 (N_3155,N_541,N_1820);
or U3156 (N_3156,N_1360,N_1387);
nand U3157 (N_3157,N_1343,N_1540);
or U3158 (N_3158,N_756,N_724);
or U3159 (N_3159,N_259,N_972);
nand U3160 (N_3160,N_1585,N_1186);
xnor U3161 (N_3161,N_538,N_1096);
xnor U3162 (N_3162,N_863,N_286);
or U3163 (N_3163,N_139,N_1956);
nand U3164 (N_3164,N_282,N_345);
nand U3165 (N_3165,N_618,N_186);
xor U3166 (N_3166,N_1408,N_1660);
nor U3167 (N_3167,N_379,N_671);
nor U3168 (N_3168,N_1730,N_588);
nand U3169 (N_3169,N_1286,N_855);
and U3170 (N_3170,N_62,N_309);
xor U3171 (N_3171,N_1020,N_115);
xor U3172 (N_3172,N_1227,N_1919);
or U3173 (N_3173,N_1976,N_1039);
nand U3174 (N_3174,N_432,N_986);
xor U3175 (N_3175,N_206,N_453);
nor U3176 (N_3176,N_1604,N_1681);
or U3177 (N_3177,N_1306,N_476);
and U3178 (N_3178,N_767,N_1197);
nand U3179 (N_3179,N_1364,N_1584);
or U3180 (N_3180,N_1684,N_1300);
nand U3181 (N_3181,N_106,N_1688);
and U3182 (N_3182,N_1034,N_1982);
nand U3183 (N_3183,N_207,N_1958);
nor U3184 (N_3184,N_22,N_1454);
xor U3185 (N_3185,N_348,N_1564);
nand U3186 (N_3186,N_299,N_122);
nor U3187 (N_3187,N_909,N_464);
or U3188 (N_3188,N_73,N_1611);
nor U3189 (N_3189,N_422,N_1117);
and U3190 (N_3190,N_639,N_1413);
or U3191 (N_3191,N_99,N_1981);
nor U3192 (N_3192,N_597,N_116);
nand U3193 (N_3193,N_1345,N_244);
and U3194 (N_3194,N_1162,N_926);
xnor U3195 (N_3195,N_1558,N_607);
xor U3196 (N_3196,N_995,N_1758);
xnor U3197 (N_3197,N_1106,N_1380);
or U3198 (N_3198,N_832,N_1430);
or U3199 (N_3199,N_1311,N_1935);
and U3200 (N_3200,N_678,N_1844);
xnor U3201 (N_3201,N_1342,N_1658);
nand U3202 (N_3202,N_1039,N_890);
or U3203 (N_3203,N_1754,N_85);
and U3204 (N_3204,N_1925,N_822);
or U3205 (N_3205,N_1781,N_1159);
or U3206 (N_3206,N_936,N_460);
or U3207 (N_3207,N_1130,N_1855);
or U3208 (N_3208,N_1173,N_1620);
or U3209 (N_3209,N_201,N_1525);
or U3210 (N_3210,N_1752,N_650);
or U3211 (N_3211,N_1102,N_1233);
nand U3212 (N_3212,N_1364,N_1474);
nor U3213 (N_3213,N_1251,N_1572);
and U3214 (N_3214,N_1809,N_1929);
nand U3215 (N_3215,N_802,N_1272);
and U3216 (N_3216,N_1294,N_1817);
or U3217 (N_3217,N_49,N_899);
nor U3218 (N_3218,N_1990,N_1475);
xor U3219 (N_3219,N_675,N_301);
or U3220 (N_3220,N_813,N_499);
nand U3221 (N_3221,N_1432,N_146);
nand U3222 (N_3222,N_1443,N_891);
xnor U3223 (N_3223,N_1680,N_718);
and U3224 (N_3224,N_696,N_1622);
xnor U3225 (N_3225,N_1099,N_862);
and U3226 (N_3226,N_1073,N_912);
and U3227 (N_3227,N_73,N_1433);
and U3228 (N_3228,N_661,N_352);
nand U3229 (N_3229,N_938,N_456);
nor U3230 (N_3230,N_500,N_931);
or U3231 (N_3231,N_1295,N_468);
xnor U3232 (N_3232,N_125,N_151);
nor U3233 (N_3233,N_1052,N_1106);
or U3234 (N_3234,N_561,N_1042);
nand U3235 (N_3235,N_1155,N_784);
nand U3236 (N_3236,N_1810,N_1880);
and U3237 (N_3237,N_545,N_99);
or U3238 (N_3238,N_1516,N_256);
nand U3239 (N_3239,N_1830,N_364);
or U3240 (N_3240,N_1054,N_1617);
and U3241 (N_3241,N_1143,N_1380);
nand U3242 (N_3242,N_420,N_1965);
nand U3243 (N_3243,N_1124,N_1531);
nor U3244 (N_3244,N_251,N_704);
nor U3245 (N_3245,N_562,N_1903);
xnor U3246 (N_3246,N_577,N_1548);
nand U3247 (N_3247,N_1508,N_1454);
xor U3248 (N_3248,N_1568,N_421);
xor U3249 (N_3249,N_1623,N_1833);
nor U3250 (N_3250,N_1639,N_1101);
xor U3251 (N_3251,N_96,N_872);
or U3252 (N_3252,N_1681,N_1987);
and U3253 (N_3253,N_1944,N_202);
or U3254 (N_3254,N_474,N_1563);
and U3255 (N_3255,N_871,N_251);
or U3256 (N_3256,N_889,N_1779);
or U3257 (N_3257,N_1237,N_270);
nor U3258 (N_3258,N_1383,N_371);
xnor U3259 (N_3259,N_1072,N_418);
and U3260 (N_3260,N_610,N_805);
nand U3261 (N_3261,N_13,N_789);
nand U3262 (N_3262,N_610,N_1799);
xnor U3263 (N_3263,N_1678,N_1543);
or U3264 (N_3264,N_335,N_1368);
and U3265 (N_3265,N_727,N_976);
nor U3266 (N_3266,N_489,N_1074);
or U3267 (N_3267,N_204,N_774);
nor U3268 (N_3268,N_353,N_401);
xor U3269 (N_3269,N_1314,N_298);
and U3270 (N_3270,N_843,N_1905);
nand U3271 (N_3271,N_1663,N_1549);
xnor U3272 (N_3272,N_954,N_1517);
nand U3273 (N_3273,N_855,N_98);
nand U3274 (N_3274,N_1068,N_709);
nor U3275 (N_3275,N_585,N_223);
or U3276 (N_3276,N_1592,N_1192);
nand U3277 (N_3277,N_708,N_1915);
nor U3278 (N_3278,N_1988,N_985);
and U3279 (N_3279,N_387,N_1286);
nor U3280 (N_3280,N_1616,N_306);
nand U3281 (N_3281,N_1443,N_1497);
or U3282 (N_3282,N_474,N_982);
nor U3283 (N_3283,N_108,N_156);
or U3284 (N_3284,N_1489,N_1536);
or U3285 (N_3285,N_858,N_59);
or U3286 (N_3286,N_1361,N_1760);
nand U3287 (N_3287,N_810,N_763);
and U3288 (N_3288,N_1664,N_1533);
nand U3289 (N_3289,N_1409,N_455);
or U3290 (N_3290,N_1242,N_1670);
or U3291 (N_3291,N_1670,N_247);
xnor U3292 (N_3292,N_1172,N_366);
nand U3293 (N_3293,N_1307,N_357);
xor U3294 (N_3294,N_1749,N_1990);
and U3295 (N_3295,N_754,N_1457);
nor U3296 (N_3296,N_1812,N_857);
or U3297 (N_3297,N_290,N_919);
xor U3298 (N_3298,N_476,N_227);
or U3299 (N_3299,N_1847,N_1040);
or U3300 (N_3300,N_895,N_1142);
nand U3301 (N_3301,N_1879,N_206);
or U3302 (N_3302,N_1932,N_1672);
nand U3303 (N_3303,N_1608,N_857);
nor U3304 (N_3304,N_1043,N_1611);
nor U3305 (N_3305,N_1989,N_741);
and U3306 (N_3306,N_1576,N_1082);
nor U3307 (N_3307,N_1843,N_1205);
xor U3308 (N_3308,N_215,N_1865);
nand U3309 (N_3309,N_1121,N_935);
nor U3310 (N_3310,N_1075,N_495);
nand U3311 (N_3311,N_878,N_807);
nand U3312 (N_3312,N_1148,N_1782);
nand U3313 (N_3313,N_1610,N_1435);
or U3314 (N_3314,N_518,N_373);
or U3315 (N_3315,N_398,N_830);
or U3316 (N_3316,N_1753,N_1081);
xnor U3317 (N_3317,N_1020,N_1669);
nor U3318 (N_3318,N_85,N_1701);
nand U3319 (N_3319,N_1495,N_1119);
and U3320 (N_3320,N_399,N_857);
nand U3321 (N_3321,N_859,N_575);
and U3322 (N_3322,N_1750,N_816);
nand U3323 (N_3323,N_465,N_1755);
nor U3324 (N_3324,N_13,N_1018);
nor U3325 (N_3325,N_287,N_1885);
nand U3326 (N_3326,N_1776,N_428);
nor U3327 (N_3327,N_761,N_184);
or U3328 (N_3328,N_1085,N_1791);
and U3329 (N_3329,N_457,N_1251);
nor U3330 (N_3330,N_936,N_1585);
and U3331 (N_3331,N_1240,N_752);
or U3332 (N_3332,N_1550,N_1761);
nor U3333 (N_3333,N_434,N_48);
and U3334 (N_3334,N_159,N_1);
xor U3335 (N_3335,N_605,N_636);
or U3336 (N_3336,N_1592,N_1543);
nand U3337 (N_3337,N_226,N_1328);
xor U3338 (N_3338,N_837,N_804);
nor U3339 (N_3339,N_991,N_1478);
xnor U3340 (N_3340,N_1396,N_1956);
or U3341 (N_3341,N_501,N_274);
and U3342 (N_3342,N_1886,N_1356);
nor U3343 (N_3343,N_323,N_1441);
or U3344 (N_3344,N_1140,N_274);
or U3345 (N_3345,N_1361,N_909);
or U3346 (N_3346,N_1896,N_1197);
xnor U3347 (N_3347,N_16,N_586);
nand U3348 (N_3348,N_1386,N_473);
nor U3349 (N_3349,N_1797,N_974);
xor U3350 (N_3350,N_1165,N_1110);
nor U3351 (N_3351,N_1876,N_1001);
nand U3352 (N_3352,N_1399,N_714);
nor U3353 (N_3353,N_615,N_1008);
xnor U3354 (N_3354,N_226,N_94);
and U3355 (N_3355,N_964,N_1625);
nor U3356 (N_3356,N_1773,N_1142);
nor U3357 (N_3357,N_602,N_937);
nor U3358 (N_3358,N_1589,N_892);
nor U3359 (N_3359,N_1974,N_568);
nand U3360 (N_3360,N_1638,N_770);
nand U3361 (N_3361,N_579,N_1567);
xor U3362 (N_3362,N_839,N_125);
nand U3363 (N_3363,N_1767,N_922);
xor U3364 (N_3364,N_815,N_1587);
and U3365 (N_3365,N_1989,N_1597);
xnor U3366 (N_3366,N_1178,N_345);
and U3367 (N_3367,N_123,N_456);
xor U3368 (N_3368,N_1839,N_1959);
and U3369 (N_3369,N_1815,N_1792);
and U3370 (N_3370,N_1991,N_1978);
xnor U3371 (N_3371,N_642,N_698);
nand U3372 (N_3372,N_1474,N_1121);
and U3373 (N_3373,N_1044,N_717);
nor U3374 (N_3374,N_387,N_1833);
or U3375 (N_3375,N_1938,N_160);
or U3376 (N_3376,N_1245,N_1293);
xnor U3377 (N_3377,N_847,N_2);
or U3378 (N_3378,N_1947,N_452);
nand U3379 (N_3379,N_1263,N_880);
nor U3380 (N_3380,N_843,N_1932);
and U3381 (N_3381,N_525,N_1130);
nand U3382 (N_3382,N_1129,N_1097);
and U3383 (N_3383,N_1637,N_1525);
nor U3384 (N_3384,N_1616,N_416);
or U3385 (N_3385,N_1060,N_1430);
xor U3386 (N_3386,N_623,N_662);
nor U3387 (N_3387,N_72,N_1378);
nor U3388 (N_3388,N_961,N_128);
or U3389 (N_3389,N_835,N_28);
xnor U3390 (N_3390,N_1857,N_781);
xor U3391 (N_3391,N_1106,N_1745);
and U3392 (N_3392,N_35,N_1698);
or U3393 (N_3393,N_1968,N_812);
or U3394 (N_3394,N_1752,N_1704);
nor U3395 (N_3395,N_1999,N_1065);
nor U3396 (N_3396,N_1354,N_1213);
or U3397 (N_3397,N_1976,N_1893);
and U3398 (N_3398,N_657,N_633);
or U3399 (N_3399,N_581,N_391);
or U3400 (N_3400,N_48,N_639);
and U3401 (N_3401,N_1264,N_1912);
xnor U3402 (N_3402,N_400,N_1484);
nor U3403 (N_3403,N_1558,N_1345);
nor U3404 (N_3404,N_1940,N_1279);
nor U3405 (N_3405,N_679,N_191);
and U3406 (N_3406,N_1211,N_563);
or U3407 (N_3407,N_1845,N_1884);
or U3408 (N_3408,N_308,N_875);
xnor U3409 (N_3409,N_1919,N_59);
and U3410 (N_3410,N_1246,N_1076);
nand U3411 (N_3411,N_1599,N_1196);
or U3412 (N_3412,N_403,N_1825);
or U3413 (N_3413,N_1747,N_1013);
nor U3414 (N_3414,N_1060,N_1317);
or U3415 (N_3415,N_43,N_347);
nand U3416 (N_3416,N_1550,N_49);
xor U3417 (N_3417,N_1497,N_221);
and U3418 (N_3418,N_1007,N_1798);
and U3419 (N_3419,N_966,N_1280);
xnor U3420 (N_3420,N_89,N_171);
and U3421 (N_3421,N_1840,N_881);
nor U3422 (N_3422,N_1791,N_79);
or U3423 (N_3423,N_677,N_667);
nor U3424 (N_3424,N_13,N_1697);
or U3425 (N_3425,N_1304,N_804);
and U3426 (N_3426,N_718,N_316);
nand U3427 (N_3427,N_537,N_1851);
or U3428 (N_3428,N_294,N_1498);
and U3429 (N_3429,N_1673,N_1822);
nor U3430 (N_3430,N_701,N_196);
nor U3431 (N_3431,N_526,N_290);
nand U3432 (N_3432,N_436,N_1944);
xnor U3433 (N_3433,N_192,N_491);
nand U3434 (N_3434,N_1815,N_1176);
xnor U3435 (N_3435,N_170,N_1492);
xor U3436 (N_3436,N_1049,N_1279);
nor U3437 (N_3437,N_118,N_1270);
nand U3438 (N_3438,N_1263,N_1235);
and U3439 (N_3439,N_95,N_409);
or U3440 (N_3440,N_618,N_779);
or U3441 (N_3441,N_1439,N_187);
and U3442 (N_3442,N_1067,N_754);
and U3443 (N_3443,N_659,N_1903);
xor U3444 (N_3444,N_64,N_86);
nand U3445 (N_3445,N_1495,N_1117);
nor U3446 (N_3446,N_1617,N_1473);
nor U3447 (N_3447,N_1796,N_106);
nor U3448 (N_3448,N_1160,N_1328);
nor U3449 (N_3449,N_1795,N_1778);
xor U3450 (N_3450,N_62,N_1644);
xor U3451 (N_3451,N_1345,N_1378);
xor U3452 (N_3452,N_886,N_1670);
nand U3453 (N_3453,N_807,N_1886);
and U3454 (N_3454,N_176,N_663);
nor U3455 (N_3455,N_576,N_1075);
nor U3456 (N_3456,N_344,N_616);
nor U3457 (N_3457,N_820,N_998);
and U3458 (N_3458,N_1645,N_1746);
nand U3459 (N_3459,N_837,N_1133);
xnor U3460 (N_3460,N_1265,N_783);
or U3461 (N_3461,N_1270,N_122);
xnor U3462 (N_3462,N_1770,N_1480);
nand U3463 (N_3463,N_1184,N_447);
nand U3464 (N_3464,N_318,N_855);
xor U3465 (N_3465,N_1315,N_1683);
nor U3466 (N_3466,N_1044,N_1169);
nand U3467 (N_3467,N_940,N_196);
nand U3468 (N_3468,N_113,N_186);
and U3469 (N_3469,N_1542,N_1231);
and U3470 (N_3470,N_792,N_1218);
nor U3471 (N_3471,N_943,N_1116);
xor U3472 (N_3472,N_1723,N_1580);
or U3473 (N_3473,N_350,N_1004);
and U3474 (N_3474,N_457,N_260);
or U3475 (N_3475,N_1523,N_945);
xnor U3476 (N_3476,N_786,N_785);
and U3477 (N_3477,N_69,N_242);
xnor U3478 (N_3478,N_1878,N_434);
xor U3479 (N_3479,N_559,N_147);
and U3480 (N_3480,N_1475,N_615);
xnor U3481 (N_3481,N_385,N_1701);
and U3482 (N_3482,N_586,N_80);
nand U3483 (N_3483,N_1428,N_1765);
xor U3484 (N_3484,N_160,N_1421);
or U3485 (N_3485,N_1684,N_1486);
or U3486 (N_3486,N_1317,N_1255);
nand U3487 (N_3487,N_1082,N_556);
nor U3488 (N_3488,N_1074,N_817);
xor U3489 (N_3489,N_73,N_1675);
and U3490 (N_3490,N_1168,N_1866);
or U3491 (N_3491,N_61,N_911);
and U3492 (N_3492,N_1852,N_1391);
and U3493 (N_3493,N_1778,N_1359);
xor U3494 (N_3494,N_915,N_1585);
and U3495 (N_3495,N_1543,N_521);
nand U3496 (N_3496,N_1078,N_364);
xnor U3497 (N_3497,N_620,N_616);
nor U3498 (N_3498,N_33,N_985);
nand U3499 (N_3499,N_1243,N_1304);
nor U3500 (N_3500,N_959,N_1292);
xnor U3501 (N_3501,N_1556,N_1662);
nor U3502 (N_3502,N_1113,N_724);
nand U3503 (N_3503,N_972,N_574);
nand U3504 (N_3504,N_741,N_833);
or U3505 (N_3505,N_1724,N_1400);
and U3506 (N_3506,N_1739,N_163);
nor U3507 (N_3507,N_338,N_133);
or U3508 (N_3508,N_314,N_1008);
and U3509 (N_3509,N_749,N_1161);
or U3510 (N_3510,N_1816,N_1103);
nor U3511 (N_3511,N_477,N_1204);
and U3512 (N_3512,N_1713,N_132);
nand U3513 (N_3513,N_621,N_12);
and U3514 (N_3514,N_1570,N_784);
or U3515 (N_3515,N_1384,N_1725);
or U3516 (N_3516,N_1396,N_1517);
and U3517 (N_3517,N_1501,N_795);
or U3518 (N_3518,N_1792,N_83);
nor U3519 (N_3519,N_1578,N_373);
nor U3520 (N_3520,N_1508,N_823);
or U3521 (N_3521,N_1412,N_1723);
nor U3522 (N_3522,N_708,N_1093);
nor U3523 (N_3523,N_417,N_1472);
or U3524 (N_3524,N_1488,N_1172);
nor U3525 (N_3525,N_528,N_1936);
nor U3526 (N_3526,N_1931,N_1312);
and U3527 (N_3527,N_1898,N_1702);
xnor U3528 (N_3528,N_1518,N_1810);
xnor U3529 (N_3529,N_1837,N_715);
or U3530 (N_3530,N_1113,N_660);
xor U3531 (N_3531,N_1618,N_24);
or U3532 (N_3532,N_1815,N_1967);
and U3533 (N_3533,N_1352,N_1369);
or U3534 (N_3534,N_125,N_1723);
xor U3535 (N_3535,N_123,N_321);
or U3536 (N_3536,N_1353,N_1599);
and U3537 (N_3537,N_959,N_1734);
xnor U3538 (N_3538,N_31,N_596);
nand U3539 (N_3539,N_1455,N_1751);
nand U3540 (N_3540,N_1398,N_545);
nand U3541 (N_3541,N_668,N_972);
or U3542 (N_3542,N_178,N_174);
and U3543 (N_3543,N_1800,N_1357);
nand U3544 (N_3544,N_684,N_833);
nor U3545 (N_3545,N_1534,N_1227);
and U3546 (N_3546,N_1321,N_735);
nand U3547 (N_3547,N_752,N_542);
or U3548 (N_3548,N_453,N_284);
nor U3549 (N_3549,N_1535,N_1037);
nor U3550 (N_3550,N_964,N_1839);
or U3551 (N_3551,N_1359,N_1843);
nand U3552 (N_3552,N_1143,N_894);
and U3553 (N_3553,N_1785,N_421);
and U3554 (N_3554,N_1393,N_1873);
xnor U3555 (N_3555,N_808,N_93);
xor U3556 (N_3556,N_1948,N_1254);
nand U3557 (N_3557,N_705,N_1110);
or U3558 (N_3558,N_1855,N_52);
nand U3559 (N_3559,N_1136,N_253);
nor U3560 (N_3560,N_1138,N_1813);
xor U3561 (N_3561,N_1454,N_718);
xnor U3562 (N_3562,N_1643,N_613);
nand U3563 (N_3563,N_316,N_293);
or U3564 (N_3564,N_296,N_88);
or U3565 (N_3565,N_1748,N_1706);
and U3566 (N_3566,N_558,N_364);
or U3567 (N_3567,N_1239,N_646);
and U3568 (N_3568,N_862,N_1141);
and U3569 (N_3569,N_816,N_803);
xnor U3570 (N_3570,N_1779,N_329);
or U3571 (N_3571,N_917,N_18);
xor U3572 (N_3572,N_66,N_1254);
nor U3573 (N_3573,N_1251,N_1321);
xnor U3574 (N_3574,N_1197,N_1158);
and U3575 (N_3575,N_1662,N_1410);
nor U3576 (N_3576,N_1443,N_134);
nor U3577 (N_3577,N_1671,N_1978);
xor U3578 (N_3578,N_626,N_1153);
xnor U3579 (N_3579,N_902,N_1405);
xor U3580 (N_3580,N_1748,N_928);
nand U3581 (N_3581,N_729,N_1636);
or U3582 (N_3582,N_1278,N_992);
nand U3583 (N_3583,N_594,N_1226);
nand U3584 (N_3584,N_3,N_1807);
xnor U3585 (N_3585,N_841,N_357);
nand U3586 (N_3586,N_1229,N_1517);
nor U3587 (N_3587,N_1030,N_1413);
or U3588 (N_3588,N_987,N_315);
or U3589 (N_3589,N_693,N_955);
xnor U3590 (N_3590,N_684,N_458);
and U3591 (N_3591,N_595,N_270);
and U3592 (N_3592,N_650,N_548);
or U3593 (N_3593,N_1466,N_53);
or U3594 (N_3594,N_867,N_1375);
xor U3595 (N_3595,N_1073,N_1396);
nand U3596 (N_3596,N_896,N_1053);
nand U3597 (N_3597,N_1033,N_724);
or U3598 (N_3598,N_629,N_1422);
and U3599 (N_3599,N_965,N_1234);
or U3600 (N_3600,N_1585,N_1260);
nor U3601 (N_3601,N_1882,N_910);
nor U3602 (N_3602,N_325,N_1811);
nand U3603 (N_3603,N_1944,N_1004);
nand U3604 (N_3604,N_632,N_1015);
nor U3605 (N_3605,N_719,N_794);
nor U3606 (N_3606,N_23,N_1369);
xnor U3607 (N_3607,N_497,N_1935);
xnor U3608 (N_3608,N_369,N_1339);
and U3609 (N_3609,N_794,N_1477);
nor U3610 (N_3610,N_1426,N_642);
xor U3611 (N_3611,N_1074,N_125);
and U3612 (N_3612,N_1579,N_1407);
or U3613 (N_3613,N_1368,N_1956);
xnor U3614 (N_3614,N_918,N_1261);
nor U3615 (N_3615,N_926,N_1145);
xor U3616 (N_3616,N_129,N_390);
or U3617 (N_3617,N_1757,N_1951);
nand U3618 (N_3618,N_1247,N_1121);
nor U3619 (N_3619,N_1320,N_190);
xnor U3620 (N_3620,N_1225,N_551);
or U3621 (N_3621,N_542,N_265);
or U3622 (N_3622,N_1605,N_131);
nand U3623 (N_3623,N_1567,N_212);
nand U3624 (N_3624,N_126,N_778);
nor U3625 (N_3625,N_4,N_635);
and U3626 (N_3626,N_1789,N_382);
nor U3627 (N_3627,N_242,N_1879);
xor U3628 (N_3628,N_1117,N_502);
or U3629 (N_3629,N_282,N_1987);
or U3630 (N_3630,N_1221,N_1848);
and U3631 (N_3631,N_232,N_1572);
xnor U3632 (N_3632,N_1264,N_914);
and U3633 (N_3633,N_607,N_1654);
xor U3634 (N_3634,N_1684,N_265);
xor U3635 (N_3635,N_1986,N_651);
xnor U3636 (N_3636,N_1425,N_266);
nand U3637 (N_3637,N_1703,N_532);
nor U3638 (N_3638,N_1153,N_268);
nor U3639 (N_3639,N_1660,N_1118);
nor U3640 (N_3640,N_1840,N_1603);
and U3641 (N_3641,N_134,N_1063);
nor U3642 (N_3642,N_1293,N_459);
nor U3643 (N_3643,N_1174,N_1959);
nand U3644 (N_3644,N_179,N_270);
or U3645 (N_3645,N_72,N_1394);
and U3646 (N_3646,N_1436,N_722);
xnor U3647 (N_3647,N_1451,N_19);
xor U3648 (N_3648,N_400,N_1975);
nor U3649 (N_3649,N_1982,N_502);
nor U3650 (N_3650,N_156,N_1826);
nand U3651 (N_3651,N_431,N_1214);
xor U3652 (N_3652,N_1754,N_186);
nand U3653 (N_3653,N_275,N_1799);
nand U3654 (N_3654,N_265,N_966);
nor U3655 (N_3655,N_1051,N_67);
nor U3656 (N_3656,N_778,N_1159);
or U3657 (N_3657,N_766,N_88);
xnor U3658 (N_3658,N_1019,N_1440);
nand U3659 (N_3659,N_1936,N_1247);
nand U3660 (N_3660,N_1134,N_1669);
nor U3661 (N_3661,N_616,N_966);
nand U3662 (N_3662,N_441,N_1386);
or U3663 (N_3663,N_336,N_550);
nor U3664 (N_3664,N_1010,N_597);
nand U3665 (N_3665,N_128,N_150);
nand U3666 (N_3666,N_1700,N_1696);
nand U3667 (N_3667,N_1147,N_967);
xnor U3668 (N_3668,N_414,N_1789);
nand U3669 (N_3669,N_1134,N_563);
nor U3670 (N_3670,N_1366,N_1898);
nor U3671 (N_3671,N_893,N_1496);
xnor U3672 (N_3672,N_1515,N_1667);
and U3673 (N_3673,N_958,N_887);
and U3674 (N_3674,N_1049,N_168);
xor U3675 (N_3675,N_587,N_1212);
xor U3676 (N_3676,N_1574,N_1509);
nor U3677 (N_3677,N_1616,N_1641);
xor U3678 (N_3678,N_524,N_119);
nand U3679 (N_3679,N_229,N_1132);
or U3680 (N_3680,N_1336,N_577);
xor U3681 (N_3681,N_1488,N_552);
and U3682 (N_3682,N_103,N_874);
nor U3683 (N_3683,N_1819,N_1809);
nand U3684 (N_3684,N_1579,N_1841);
xnor U3685 (N_3685,N_1791,N_1609);
xnor U3686 (N_3686,N_1741,N_1300);
nor U3687 (N_3687,N_797,N_897);
nor U3688 (N_3688,N_855,N_1194);
xor U3689 (N_3689,N_1844,N_818);
xnor U3690 (N_3690,N_682,N_724);
and U3691 (N_3691,N_309,N_850);
nor U3692 (N_3692,N_579,N_356);
nand U3693 (N_3693,N_1483,N_549);
nor U3694 (N_3694,N_719,N_1306);
xor U3695 (N_3695,N_1737,N_78);
or U3696 (N_3696,N_570,N_1676);
and U3697 (N_3697,N_385,N_1137);
nor U3698 (N_3698,N_1453,N_911);
or U3699 (N_3699,N_775,N_1920);
and U3700 (N_3700,N_116,N_384);
nand U3701 (N_3701,N_623,N_844);
nor U3702 (N_3702,N_839,N_1928);
xor U3703 (N_3703,N_278,N_765);
and U3704 (N_3704,N_977,N_1063);
xor U3705 (N_3705,N_1266,N_510);
xnor U3706 (N_3706,N_35,N_1);
or U3707 (N_3707,N_1014,N_156);
nor U3708 (N_3708,N_925,N_1257);
or U3709 (N_3709,N_385,N_469);
and U3710 (N_3710,N_1177,N_201);
or U3711 (N_3711,N_1741,N_52);
and U3712 (N_3712,N_76,N_1764);
nand U3713 (N_3713,N_476,N_427);
or U3714 (N_3714,N_924,N_977);
or U3715 (N_3715,N_1096,N_1968);
nand U3716 (N_3716,N_1709,N_964);
nor U3717 (N_3717,N_599,N_1873);
nand U3718 (N_3718,N_447,N_1727);
nand U3719 (N_3719,N_852,N_1247);
and U3720 (N_3720,N_1548,N_1104);
nor U3721 (N_3721,N_217,N_560);
or U3722 (N_3722,N_1329,N_1000);
nor U3723 (N_3723,N_927,N_508);
and U3724 (N_3724,N_1804,N_838);
xor U3725 (N_3725,N_962,N_728);
xor U3726 (N_3726,N_1658,N_1316);
and U3727 (N_3727,N_689,N_909);
and U3728 (N_3728,N_652,N_905);
or U3729 (N_3729,N_94,N_428);
nand U3730 (N_3730,N_272,N_939);
or U3731 (N_3731,N_274,N_460);
xnor U3732 (N_3732,N_1499,N_1566);
nand U3733 (N_3733,N_1568,N_996);
or U3734 (N_3734,N_432,N_746);
or U3735 (N_3735,N_1925,N_208);
or U3736 (N_3736,N_1451,N_1744);
xnor U3737 (N_3737,N_311,N_183);
and U3738 (N_3738,N_88,N_1603);
xnor U3739 (N_3739,N_879,N_1069);
or U3740 (N_3740,N_581,N_1977);
xor U3741 (N_3741,N_1026,N_525);
nor U3742 (N_3742,N_813,N_1474);
nand U3743 (N_3743,N_461,N_1426);
nor U3744 (N_3744,N_275,N_1333);
xnor U3745 (N_3745,N_239,N_243);
or U3746 (N_3746,N_1436,N_1557);
xnor U3747 (N_3747,N_1610,N_257);
xor U3748 (N_3748,N_1422,N_1417);
xnor U3749 (N_3749,N_152,N_318);
and U3750 (N_3750,N_1475,N_1879);
nand U3751 (N_3751,N_53,N_350);
or U3752 (N_3752,N_1551,N_221);
and U3753 (N_3753,N_947,N_976);
xor U3754 (N_3754,N_1971,N_1841);
nand U3755 (N_3755,N_128,N_1820);
and U3756 (N_3756,N_188,N_348);
xor U3757 (N_3757,N_1050,N_530);
xor U3758 (N_3758,N_592,N_566);
nor U3759 (N_3759,N_480,N_390);
nor U3760 (N_3760,N_1986,N_1756);
or U3761 (N_3761,N_1255,N_1543);
or U3762 (N_3762,N_1809,N_780);
xor U3763 (N_3763,N_210,N_1527);
or U3764 (N_3764,N_33,N_1766);
and U3765 (N_3765,N_1346,N_1628);
nand U3766 (N_3766,N_1076,N_321);
nor U3767 (N_3767,N_1026,N_403);
nand U3768 (N_3768,N_1500,N_310);
xor U3769 (N_3769,N_1064,N_294);
and U3770 (N_3770,N_1350,N_1577);
or U3771 (N_3771,N_433,N_248);
and U3772 (N_3772,N_66,N_474);
xor U3773 (N_3773,N_631,N_1963);
nor U3774 (N_3774,N_305,N_79);
or U3775 (N_3775,N_261,N_658);
or U3776 (N_3776,N_811,N_234);
and U3777 (N_3777,N_1547,N_1599);
and U3778 (N_3778,N_1737,N_756);
nand U3779 (N_3779,N_1393,N_838);
nand U3780 (N_3780,N_1299,N_1690);
or U3781 (N_3781,N_1772,N_144);
nand U3782 (N_3782,N_513,N_40);
nor U3783 (N_3783,N_234,N_1765);
and U3784 (N_3784,N_78,N_575);
nand U3785 (N_3785,N_1029,N_1654);
nand U3786 (N_3786,N_1047,N_770);
nand U3787 (N_3787,N_884,N_1307);
and U3788 (N_3788,N_1677,N_204);
and U3789 (N_3789,N_1881,N_1469);
nor U3790 (N_3790,N_260,N_965);
nor U3791 (N_3791,N_92,N_1823);
and U3792 (N_3792,N_1622,N_1142);
xor U3793 (N_3793,N_512,N_1067);
nor U3794 (N_3794,N_690,N_162);
nand U3795 (N_3795,N_1058,N_1660);
nand U3796 (N_3796,N_661,N_1529);
nor U3797 (N_3797,N_1773,N_533);
nor U3798 (N_3798,N_471,N_896);
nand U3799 (N_3799,N_1579,N_724);
nor U3800 (N_3800,N_1001,N_445);
or U3801 (N_3801,N_550,N_1931);
or U3802 (N_3802,N_1973,N_746);
nor U3803 (N_3803,N_712,N_102);
or U3804 (N_3804,N_1095,N_1982);
and U3805 (N_3805,N_662,N_1084);
xor U3806 (N_3806,N_0,N_1200);
and U3807 (N_3807,N_104,N_1533);
xnor U3808 (N_3808,N_76,N_1762);
nor U3809 (N_3809,N_1400,N_1437);
xor U3810 (N_3810,N_1443,N_359);
nor U3811 (N_3811,N_1604,N_933);
or U3812 (N_3812,N_94,N_1264);
nand U3813 (N_3813,N_64,N_1211);
or U3814 (N_3814,N_1425,N_1174);
and U3815 (N_3815,N_175,N_342);
xnor U3816 (N_3816,N_90,N_1843);
and U3817 (N_3817,N_329,N_1404);
and U3818 (N_3818,N_533,N_417);
nor U3819 (N_3819,N_484,N_987);
and U3820 (N_3820,N_1208,N_1545);
nor U3821 (N_3821,N_5,N_901);
or U3822 (N_3822,N_623,N_1288);
or U3823 (N_3823,N_1095,N_369);
and U3824 (N_3824,N_1621,N_985);
and U3825 (N_3825,N_1668,N_1956);
xnor U3826 (N_3826,N_715,N_144);
nor U3827 (N_3827,N_1855,N_917);
or U3828 (N_3828,N_696,N_1116);
or U3829 (N_3829,N_1600,N_1988);
nor U3830 (N_3830,N_1478,N_543);
nor U3831 (N_3831,N_704,N_1986);
nor U3832 (N_3832,N_37,N_447);
or U3833 (N_3833,N_112,N_775);
nand U3834 (N_3834,N_35,N_1415);
xnor U3835 (N_3835,N_413,N_1818);
or U3836 (N_3836,N_1234,N_226);
xnor U3837 (N_3837,N_1413,N_1910);
xor U3838 (N_3838,N_221,N_1548);
nand U3839 (N_3839,N_175,N_1611);
xor U3840 (N_3840,N_1559,N_1013);
and U3841 (N_3841,N_909,N_1851);
xor U3842 (N_3842,N_886,N_1728);
and U3843 (N_3843,N_286,N_927);
xnor U3844 (N_3844,N_1528,N_211);
or U3845 (N_3845,N_839,N_1510);
or U3846 (N_3846,N_159,N_684);
xor U3847 (N_3847,N_1165,N_1529);
and U3848 (N_3848,N_1619,N_1602);
or U3849 (N_3849,N_1138,N_287);
and U3850 (N_3850,N_1869,N_1526);
xnor U3851 (N_3851,N_609,N_1409);
and U3852 (N_3852,N_1422,N_453);
or U3853 (N_3853,N_506,N_27);
xnor U3854 (N_3854,N_1189,N_85);
nand U3855 (N_3855,N_1460,N_622);
nand U3856 (N_3856,N_1692,N_509);
nor U3857 (N_3857,N_966,N_585);
xor U3858 (N_3858,N_774,N_1608);
xor U3859 (N_3859,N_600,N_592);
xor U3860 (N_3860,N_595,N_626);
nand U3861 (N_3861,N_1482,N_1483);
nor U3862 (N_3862,N_570,N_613);
nor U3863 (N_3863,N_914,N_1938);
nor U3864 (N_3864,N_1004,N_125);
and U3865 (N_3865,N_659,N_623);
xnor U3866 (N_3866,N_607,N_1591);
nor U3867 (N_3867,N_852,N_243);
nor U3868 (N_3868,N_1923,N_1013);
or U3869 (N_3869,N_1264,N_98);
and U3870 (N_3870,N_1783,N_1901);
or U3871 (N_3871,N_1689,N_189);
nor U3872 (N_3872,N_310,N_1399);
or U3873 (N_3873,N_1002,N_833);
and U3874 (N_3874,N_1962,N_1411);
xnor U3875 (N_3875,N_1124,N_1386);
and U3876 (N_3876,N_1947,N_643);
or U3877 (N_3877,N_1600,N_1553);
xor U3878 (N_3878,N_1687,N_1180);
xnor U3879 (N_3879,N_1707,N_424);
nand U3880 (N_3880,N_1872,N_916);
xnor U3881 (N_3881,N_38,N_559);
and U3882 (N_3882,N_1327,N_1018);
or U3883 (N_3883,N_1977,N_190);
nand U3884 (N_3884,N_533,N_398);
or U3885 (N_3885,N_411,N_388);
and U3886 (N_3886,N_1270,N_1574);
and U3887 (N_3887,N_599,N_939);
or U3888 (N_3888,N_1377,N_598);
nand U3889 (N_3889,N_1869,N_1859);
or U3890 (N_3890,N_1742,N_1765);
and U3891 (N_3891,N_1032,N_338);
or U3892 (N_3892,N_1223,N_20);
xnor U3893 (N_3893,N_1359,N_1413);
nor U3894 (N_3894,N_1467,N_133);
or U3895 (N_3895,N_1463,N_849);
nor U3896 (N_3896,N_204,N_930);
xnor U3897 (N_3897,N_660,N_458);
nand U3898 (N_3898,N_1757,N_829);
nor U3899 (N_3899,N_1915,N_1450);
nand U3900 (N_3900,N_876,N_510);
and U3901 (N_3901,N_1306,N_1214);
nand U3902 (N_3902,N_1483,N_1340);
and U3903 (N_3903,N_429,N_1607);
xnor U3904 (N_3904,N_841,N_527);
and U3905 (N_3905,N_1765,N_1912);
and U3906 (N_3906,N_1935,N_1927);
or U3907 (N_3907,N_1453,N_518);
nand U3908 (N_3908,N_1180,N_230);
nand U3909 (N_3909,N_1112,N_1302);
or U3910 (N_3910,N_293,N_1994);
xor U3911 (N_3911,N_1936,N_884);
xnor U3912 (N_3912,N_226,N_119);
nor U3913 (N_3913,N_1637,N_1279);
and U3914 (N_3914,N_1097,N_354);
xnor U3915 (N_3915,N_672,N_1287);
xnor U3916 (N_3916,N_355,N_1219);
xor U3917 (N_3917,N_524,N_508);
nor U3918 (N_3918,N_1614,N_1244);
and U3919 (N_3919,N_304,N_1614);
or U3920 (N_3920,N_1116,N_1404);
and U3921 (N_3921,N_1695,N_1134);
and U3922 (N_3922,N_47,N_256);
nand U3923 (N_3923,N_1604,N_1916);
xnor U3924 (N_3924,N_316,N_291);
or U3925 (N_3925,N_1117,N_1564);
or U3926 (N_3926,N_153,N_97);
and U3927 (N_3927,N_1673,N_540);
and U3928 (N_3928,N_712,N_414);
xor U3929 (N_3929,N_902,N_1186);
and U3930 (N_3930,N_1885,N_370);
nor U3931 (N_3931,N_504,N_1343);
and U3932 (N_3932,N_377,N_1340);
xnor U3933 (N_3933,N_1490,N_229);
and U3934 (N_3934,N_736,N_305);
nor U3935 (N_3935,N_665,N_1271);
or U3936 (N_3936,N_1149,N_831);
nand U3937 (N_3937,N_1871,N_923);
nor U3938 (N_3938,N_41,N_1444);
xor U3939 (N_3939,N_840,N_1757);
xor U3940 (N_3940,N_1821,N_1752);
or U3941 (N_3941,N_1025,N_1568);
nor U3942 (N_3942,N_815,N_1358);
nor U3943 (N_3943,N_848,N_1470);
and U3944 (N_3944,N_325,N_1962);
or U3945 (N_3945,N_217,N_1378);
and U3946 (N_3946,N_1929,N_1214);
or U3947 (N_3947,N_1469,N_1583);
nor U3948 (N_3948,N_1914,N_1478);
xor U3949 (N_3949,N_1316,N_1054);
nor U3950 (N_3950,N_1673,N_1449);
or U3951 (N_3951,N_47,N_1296);
and U3952 (N_3952,N_856,N_591);
nand U3953 (N_3953,N_917,N_1231);
or U3954 (N_3954,N_437,N_1165);
nand U3955 (N_3955,N_491,N_1775);
or U3956 (N_3956,N_1959,N_802);
or U3957 (N_3957,N_1542,N_1841);
xor U3958 (N_3958,N_396,N_955);
or U3959 (N_3959,N_1045,N_842);
xnor U3960 (N_3960,N_1712,N_702);
nor U3961 (N_3961,N_1764,N_176);
nand U3962 (N_3962,N_242,N_792);
nand U3963 (N_3963,N_339,N_1527);
or U3964 (N_3964,N_718,N_362);
and U3965 (N_3965,N_1701,N_871);
nor U3966 (N_3966,N_722,N_177);
and U3967 (N_3967,N_523,N_861);
xnor U3968 (N_3968,N_782,N_280);
or U3969 (N_3969,N_1522,N_1659);
or U3970 (N_3970,N_1750,N_473);
nand U3971 (N_3971,N_252,N_852);
nor U3972 (N_3972,N_139,N_497);
xnor U3973 (N_3973,N_55,N_1574);
and U3974 (N_3974,N_931,N_987);
or U3975 (N_3975,N_788,N_31);
and U3976 (N_3976,N_365,N_282);
and U3977 (N_3977,N_1910,N_1384);
and U3978 (N_3978,N_1510,N_1149);
and U3979 (N_3979,N_1083,N_303);
nor U3980 (N_3980,N_375,N_319);
xor U3981 (N_3981,N_1254,N_1938);
or U3982 (N_3982,N_1886,N_1273);
xor U3983 (N_3983,N_1444,N_1435);
or U3984 (N_3984,N_472,N_1435);
or U3985 (N_3985,N_969,N_1382);
or U3986 (N_3986,N_90,N_704);
and U3987 (N_3987,N_787,N_1935);
nor U3988 (N_3988,N_1932,N_846);
or U3989 (N_3989,N_366,N_81);
nand U3990 (N_3990,N_1805,N_939);
nand U3991 (N_3991,N_482,N_896);
and U3992 (N_3992,N_1681,N_1410);
nor U3993 (N_3993,N_1263,N_1619);
nor U3994 (N_3994,N_1587,N_741);
and U3995 (N_3995,N_1260,N_535);
nor U3996 (N_3996,N_1462,N_141);
and U3997 (N_3997,N_258,N_1761);
and U3998 (N_3998,N_184,N_1421);
xnor U3999 (N_3999,N_1802,N_716);
and U4000 (N_4000,N_3505,N_3456);
nor U4001 (N_4001,N_3884,N_2132);
nand U4002 (N_4002,N_2416,N_3261);
xor U4003 (N_4003,N_3975,N_2507);
xnor U4004 (N_4004,N_3722,N_2925);
and U4005 (N_4005,N_3155,N_3385);
and U4006 (N_4006,N_3867,N_3855);
nor U4007 (N_4007,N_2640,N_2524);
or U4008 (N_4008,N_2949,N_2633);
and U4009 (N_4009,N_2411,N_2577);
or U4010 (N_4010,N_2141,N_3102);
nor U4011 (N_4011,N_3428,N_3131);
nor U4012 (N_4012,N_2704,N_2923);
nor U4013 (N_4013,N_2555,N_2405);
and U4014 (N_4014,N_2724,N_3213);
xnor U4015 (N_4015,N_3694,N_3984);
or U4016 (N_4016,N_2015,N_2442);
and U4017 (N_4017,N_3240,N_3266);
nand U4018 (N_4018,N_3289,N_2283);
nand U4019 (N_4019,N_3055,N_3317);
nand U4020 (N_4020,N_3424,N_2478);
and U4021 (N_4021,N_3976,N_2368);
xnor U4022 (N_4022,N_3189,N_3046);
nor U4023 (N_4023,N_2615,N_2655);
nor U4024 (N_4024,N_2729,N_2146);
nor U4025 (N_4025,N_2152,N_2398);
nor U4026 (N_4026,N_3246,N_3286);
and U4027 (N_4027,N_3329,N_2552);
or U4028 (N_4028,N_2099,N_3034);
and U4029 (N_4029,N_2224,N_2927);
nor U4030 (N_4030,N_2173,N_2901);
xnor U4031 (N_4031,N_2785,N_3672);
and U4032 (N_4032,N_2847,N_2871);
nor U4033 (N_4033,N_2906,N_3302);
and U4034 (N_4034,N_2907,N_3402);
nor U4035 (N_4035,N_2941,N_3258);
or U4036 (N_4036,N_3490,N_2199);
and U4037 (N_4037,N_2686,N_3190);
nand U4038 (N_4038,N_3099,N_3857);
and U4039 (N_4039,N_2170,N_2497);
nor U4040 (N_4040,N_3212,N_3679);
nand U4041 (N_4041,N_3997,N_2825);
and U4042 (N_4042,N_3335,N_3815);
and U4043 (N_4043,N_3122,N_3520);
xnor U4044 (N_4044,N_3780,N_2761);
or U4045 (N_4045,N_3935,N_3886);
nor U4046 (N_4046,N_3928,N_2214);
xnor U4047 (N_4047,N_2494,N_2360);
xnor U4048 (N_4048,N_3595,N_2365);
or U4049 (N_4049,N_2786,N_3795);
xnor U4050 (N_4050,N_2010,N_2516);
nor U4051 (N_4051,N_2450,N_3382);
nor U4052 (N_4052,N_3929,N_3743);
nor U4053 (N_4053,N_3982,N_2429);
or U4054 (N_4054,N_2008,N_2328);
nor U4055 (N_4055,N_3872,N_3902);
or U4056 (N_4056,N_2462,N_3836);
nor U4057 (N_4057,N_2459,N_3469);
nor U4058 (N_4058,N_3084,N_2805);
nor U4059 (N_4059,N_2568,N_2231);
and U4060 (N_4060,N_2994,N_3360);
or U4061 (N_4061,N_2496,N_3121);
nand U4062 (N_4062,N_2080,N_3254);
or U4063 (N_4063,N_3577,N_3790);
and U4064 (N_4064,N_2620,N_2216);
nand U4065 (N_4065,N_2523,N_2361);
or U4066 (N_4066,N_2610,N_2647);
nand U4067 (N_4067,N_3091,N_2728);
or U4068 (N_4068,N_2066,N_2566);
xnor U4069 (N_4069,N_2409,N_2990);
and U4070 (N_4070,N_3852,N_2591);
and U4071 (N_4071,N_3847,N_2401);
xor U4072 (N_4072,N_2465,N_2318);
nand U4073 (N_4073,N_2322,N_3410);
xor U4074 (N_4074,N_3858,N_2469);
nand U4075 (N_4075,N_2707,N_2626);
or U4076 (N_4076,N_3012,N_3047);
nor U4077 (N_4077,N_2210,N_2977);
nand U4078 (N_4078,N_3863,N_2787);
xnor U4079 (N_4079,N_2940,N_2364);
nand U4080 (N_4080,N_3404,N_3217);
nor U4081 (N_4081,N_3796,N_3590);
nand U4082 (N_4082,N_2747,N_2102);
nor U4083 (N_4083,N_3879,N_2354);
xor U4084 (N_4084,N_3005,N_3609);
and U4085 (N_4085,N_3521,N_2850);
and U4086 (N_4086,N_2054,N_3262);
nand U4087 (N_4087,N_2910,N_3116);
or U4088 (N_4088,N_2315,N_2520);
nand U4089 (N_4089,N_3371,N_2646);
and U4090 (N_4090,N_2154,N_3831);
nand U4091 (N_4091,N_3363,N_3378);
nor U4092 (N_4092,N_2197,N_3088);
and U4093 (N_4093,N_2912,N_3561);
or U4094 (N_4094,N_2206,N_3958);
nand U4095 (N_4095,N_2914,N_2299);
xor U4096 (N_4096,N_2612,N_3175);
nand U4097 (N_4097,N_3808,N_2083);
xor U4098 (N_4098,N_3137,N_2930);
nand U4099 (N_4099,N_3144,N_2426);
xnor U4100 (N_4100,N_3687,N_2684);
and U4101 (N_4101,N_3299,N_2466);
nor U4102 (N_4102,N_2413,N_2456);
or U4103 (N_4103,N_3713,N_3946);
or U4104 (N_4104,N_2943,N_3582);
nand U4105 (N_4105,N_3472,N_2394);
nor U4106 (N_4106,N_2300,N_3560);
nand U4107 (N_4107,N_3032,N_3451);
and U4108 (N_4108,N_2585,N_3650);
xnor U4109 (N_4109,N_2533,N_2603);
and U4110 (N_4110,N_3011,N_2571);
nor U4111 (N_4111,N_3699,N_2040);
nand U4112 (N_4112,N_3653,N_3541);
nor U4113 (N_4113,N_3533,N_2230);
and U4114 (N_4114,N_2195,N_3072);
and U4115 (N_4115,N_2713,N_3550);
nor U4116 (N_4116,N_3422,N_2500);
xor U4117 (N_4117,N_2295,N_2415);
nor U4118 (N_4118,N_2860,N_2498);
and U4119 (N_4119,N_2864,N_2277);
nor U4120 (N_4120,N_2726,N_2350);
nor U4121 (N_4121,N_2447,N_3986);
nand U4122 (N_4122,N_2512,N_2699);
xnor U4123 (N_4123,N_2262,N_3501);
and U4124 (N_4124,N_3898,N_2079);
or U4125 (N_4125,N_2420,N_3369);
and U4126 (N_4126,N_3330,N_2117);
nor U4127 (N_4127,N_3380,N_3983);
and U4128 (N_4128,N_2878,N_2280);
nand U4129 (N_4129,N_2275,N_2103);
nand U4130 (N_4130,N_3700,N_2693);
xor U4131 (N_4131,N_2900,N_3532);
and U4132 (N_4132,N_2888,N_3479);
nor U4133 (N_4133,N_3018,N_2711);
xor U4134 (N_4134,N_3548,N_3803);
nand U4135 (N_4135,N_2880,N_3639);
xor U4136 (N_4136,N_2624,N_2391);
and U4137 (N_4137,N_3773,N_3914);
nand U4138 (N_4138,N_3905,N_2619);
and U4139 (N_4139,N_2959,N_2736);
nand U4140 (N_4140,N_2869,N_3370);
or U4141 (N_4141,N_2379,N_2636);
or U4142 (N_4142,N_3497,N_3324);
or U4143 (N_4143,N_2444,N_3429);
or U4144 (N_4144,N_2521,N_2928);
or U4145 (N_4145,N_2695,N_2944);
and U4146 (N_4146,N_2898,N_3411);
nor U4147 (N_4147,N_3792,N_2667);
nand U4148 (N_4148,N_3513,N_2605);
nor U4149 (N_4149,N_3383,N_2282);
or U4150 (N_4150,N_3333,N_2443);
xnor U4151 (N_4151,N_2313,N_3204);
xor U4152 (N_4152,N_3964,N_2338);
nor U4153 (N_4153,N_2806,N_3089);
nand U4154 (N_4154,N_3060,N_2092);
xnor U4155 (N_4155,N_2219,N_2669);
and U4156 (N_4156,N_2593,N_3887);
nand U4157 (N_4157,N_2168,N_3606);
nand U4158 (N_4158,N_2134,N_3419);
nand U4159 (N_4159,N_3090,N_3970);
nand U4160 (N_4160,N_2376,N_3686);
and U4161 (N_4161,N_3485,N_3148);
nand U4162 (N_4162,N_2233,N_3705);
and U4163 (N_4163,N_2798,N_2588);
nor U4164 (N_4164,N_2094,N_3556);
or U4165 (N_4165,N_2823,N_2853);
or U4166 (N_4166,N_3054,N_2009);
or U4167 (N_4167,N_2471,N_2001);
nand U4168 (N_4168,N_2635,N_2399);
xor U4169 (N_4169,N_2461,N_2085);
nor U4170 (N_4170,N_3519,N_2375);
xor U4171 (N_4171,N_3373,N_2263);
xor U4172 (N_4172,N_3647,N_3197);
xnor U4173 (N_4173,N_3080,N_3656);
or U4174 (N_4174,N_3292,N_2205);
and U4175 (N_4175,N_2664,N_2563);
and U4176 (N_4176,N_2683,N_3587);
nand U4177 (N_4177,N_2039,N_2653);
nand U4178 (N_4178,N_2939,N_2915);
nand U4179 (N_4179,N_2885,N_2631);
xor U4180 (N_4180,N_2169,N_2202);
nand U4181 (N_4181,N_3086,N_2722);
and U4182 (N_4182,N_2858,N_3649);
or U4183 (N_4183,N_2757,N_3515);
xnor U4184 (N_4184,N_3381,N_3284);
and U4185 (N_4185,N_3637,N_2529);
nor U4186 (N_4186,N_2709,N_2830);
or U4187 (N_4187,N_3001,N_3162);
xnor U4188 (N_4188,N_3053,N_2650);
nand U4189 (N_4189,N_2998,N_2922);
nand U4190 (N_4190,N_3807,N_3387);
xnor U4191 (N_4191,N_2799,N_3010);
nor U4192 (N_4192,N_2258,N_3719);
and U4193 (N_4193,N_2019,N_2539);
or U4194 (N_4194,N_2307,N_3889);
and U4195 (N_4195,N_2362,N_2266);
nand U4196 (N_4196,N_2890,N_3526);
nand U4197 (N_4197,N_3483,N_2984);
xor U4198 (N_4198,N_2622,N_3608);
nor U4199 (N_4199,N_3247,N_3978);
or U4200 (N_4200,N_3814,N_3510);
nor U4201 (N_4201,N_2408,N_3017);
xnor U4202 (N_4202,N_2694,N_3095);
and U4203 (N_4203,N_3002,N_2114);
xor U4204 (N_4204,N_3837,N_2034);
or U4205 (N_4205,N_3665,N_3123);
nand U4206 (N_4206,N_2112,N_3899);
nand U4207 (N_4207,N_3165,N_3822);
or U4208 (N_4208,N_2316,N_3124);
and U4209 (N_4209,N_3308,N_3833);
or U4210 (N_4210,N_3025,N_2511);
nand U4211 (N_4211,N_2078,N_3633);
or U4212 (N_4212,N_2983,N_2979);
and U4213 (N_4213,N_2573,N_3912);
or U4214 (N_4214,N_2164,N_2041);
and U4215 (N_4215,N_2732,N_2291);
or U4216 (N_4216,N_3974,N_2887);
and U4217 (N_4217,N_3117,N_3104);
and U4218 (N_4218,N_3127,N_3540);
and U4219 (N_4219,N_3442,N_2175);
or U4220 (N_4220,N_3991,N_3888);
xor U4221 (N_4221,N_3600,N_3136);
or U4222 (N_4222,N_3075,N_2333);
nor U4223 (N_4223,N_3923,N_3006);
or U4224 (N_4224,N_3563,N_3279);
nand U4225 (N_4225,N_2611,N_3253);
nor U4226 (N_4226,N_3830,N_3188);
xnor U4227 (N_4227,N_3498,N_3695);
nand U4228 (N_4228,N_2086,N_3750);
nand U4229 (N_4229,N_2933,N_2926);
nand U4230 (N_4230,N_2562,N_2808);
or U4231 (N_4231,N_3527,N_3846);
nand U4232 (N_4232,N_2011,N_3149);
or U4233 (N_4233,N_3697,N_2658);
or U4234 (N_4234,N_2832,N_3715);
and U4235 (N_4235,N_2119,N_2675);
nand U4236 (N_4236,N_2839,N_2292);
or U4237 (N_4237,N_3584,N_3937);
and U4238 (N_4238,N_2951,N_3871);
and U4239 (N_4239,N_2232,N_2186);
and U4240 (N_4240,N_3542,N_2139);
nor U4241 (N_4241,N_2642,N_3783);
xor U4242 (N_4242,N_3921,N_2337);
xnor U4243 (N_4243,N_2595,N_2198);
or U4244 (N_4244,N_2881,N_3763);
and U4245 (N_4245,N_3023,N_3327);
or U4246 (N_4246,N_3824,N_3314);
xor U4247 (N_4247,N_3666,N_2522);
xor U4248 (N_4248,N_2892,N_2059);
nor U4249 (N_4249,N_3843,N_2953);
nand U4250 (N_4250,N_3000,N_2784);
nor U4251 (N_4251,N_3907,N_3657);
xor U4252 (N_4252,N_3244,N_2921);
xnor U4253 (N_4253,N_3630,N_3667);
nand U4254 (N_4254,N_3446,N_3282);
nor U4255 (N_4255,N_2879,N_2381);
or U4256 (N_4256,N_3441,N_2614);
or U4257 (N_4257,N_2740,N_3225);
nor U4258 (N_4258,N_3932,N_3361);
xnor U4259 (N_4259,N_2848,N_3919);
xor U4260 (N_4260,N_3045,N_3249);
nor U4261 (N_4261,N_2913,N_3374);
xor U4262 (N_4262,N_2489,N_3746);
or U4263 (N_4263,N_2004,N_2816);
and U4264 (N_4264,N_2358,N_3107);
or U4265 (N_4265,N_2666,N_3161);
xor U4266 (N_4266,N_3892,N_2673);
or U4267 (N_4267,N_3063,N_2543);
or U4268 (N_4268,N_2672,N_2731);
and U4269 (N_4269,N_2145,N_3678);
and U4270 (N_4270,N_3029,N_2430);
or U4271 (N_4271,N_2662,N_3627);
and U4272 (N_4272,N_3463,N_3480);
nand U4273 (N_4273,N_2796,N_2135);
xnor U4274 (N_4274,N_2918,N_3328);
or U4275 (N_4275,N_2441,N_3789);
nand U4276 (N_4276,N_2685,N_2730);
xnor U4277 (N_4277,N_2965,N_3942);
or U4278 (N_4278,N_3818,N_3506);
nand U4279 (N_4279,N_3464,N_3893);
nor U4280 (N_4280,N_2661,N_3163);
nor U4281 (N_4281,N_3870,N_3358);
nor U4282 (N_4282,N_3890,N_3239);
and U4283 (N_4283,N_3848,N_2395);
and U4284 (N_4284,N_2764,N_3603);
or U4285 (N_4285,N_3977,N_3557);
xor U4286 (N_4286,N_2826,N_2668);
nor U4287 (N_4287,N_2705,N_3399);
and U4288 (N_4288,N_3634,N_3351);
nor U4289 (N_4289,N_3268,N_2625);
and U4290 (N_4290,N_2517,N_2222);
nor U4291 (N_4291,N_3660,N_2296);
nand U4292 (N_4292,N_2717,N_3431);
nor U4293 (N_4293,N_2963,N_2301);
and U4294 (N_4294,N_3409,N_2437);
or U4295 (N_4295,N_2800,N_2957);
nor U4296 (N_4296,N_2075,N_2213);
nor U4297 (N_4297,N_3841,N_2254);
nand U4298 (N_4298,N_3181,N_2166);
and U4299 (N_4299,N_3891,N_2810);
nand U4300 (N_4300,N_2710,N_2235);
nand U4301 (N_4301,N_2064,N_2968);
nor U4302 (N_4302,N_2209,N_2976);
xnor U4303 (N_4303,N_2087,N_2992);
nor U4304 (N_4304,N_3448,N_2643);
or U4305 (N_4305,N_2884,N_3384);
and U4306 (N_4306,N_3873,N_2062);
or U4307 (N_4307,N_2988,N_2093);
xor U4308 (N_4308,N_3543,N_2618);
xor U4309 (N_4309,N_3176,N_2654);
or U4310 (N_4310,N_3622,N_3341);
or U4311 (N_4311,N_3432,N_3264);
and U4312 (N_4312,N_2767,N_2743);
and U4313 (N_4313,N_3015,N_3294);
or U4314 (N_4314,N_3153,N_2870);
or U4315 (N_4315,N_3169,N_2557);
xnor U4316 (N_4316,N_2273,N_3154);
or U4317 (N_4317,N_2801,N_3486);
nor U4318 (N_4318,N_3069,N_3680);
and U4319 (N_4319,N_3575,N_3337);
nor U4320 (N_4320,N_2423,N_3503);
nor U4321 (N_4321,N_2821,N_2116);
nor U4322 (N_4322,N_3493,N_3979);
xor U4323 (N_4323,N_3273,N_3586);
xor U4324 (N_4324,N_3347,N_3927);
nor U4325 (N_4325,N_3798,N_2644);
or U4326 (N_4326,N_3717,N_3737);
xnor U4327 (N_4327,N_2439,N_3875);
and U4328 (N_4328,N_2783,N_2894);
or U4329 (N_4329,N_2495,N_3911);
xor U4330 (N_4330,N_2025,N_3224);
or U4331 (N_4331,N_3462,N_3305);
xnor U4332 (N_4332,N_2428,N_3613);
and U4333 (N_4333,N_3477,N_3531);
nor U4334 (N_4334,N_2765,N_3635);
nor U4335 (N_4335,N_3570,N_3825);
and U4336 (N_4336,N_3673,N_2440);
nor U4337 (N_4337,N_3955,N_3801);
xnor U4338 (N_4338,N_2842,N_3832);
and U4339 (N_4339,N_2306,N_3147);
nor U4340 (N_4340,N_2274,N_2127);
nor U4341 (N_4341,N_3194,N_2594);
and U4342 (N_4342,N_2128,N_3707);
and U4343 (N_4343,N_2476,N_3767);
nor U4344 (N_4344,N_3934,N_2422);
and U4345 (N_4345,N_3152,N_2929);
nor U4346 (N_4346,N_3571,N_3438);
nor U4347 (N_4347,N_3800,N_2745);
nor U4348 (N_4348,N_2071,N_3476);
or U4349 (N_4349,N_3222,N_2804);
nor U4350 (N_4350,N_2972,N_3396);
nor U4351 (N_4351,N_2560,N_2966);
nor U4352 (N_4352,N_2866,N_3903);
and U4353 (N_4353,N_3035,N_3158);
or U4354 (N_4354,N_3945,N_3272);
and U4355 (N_4355,N_2601,N_3619);
xnor U4356 (N_4356,N_2113,N_2244);
xnor U4357 (N_4357,N_3952,N_3338);
nand U4358 (N_4358,N_3320,N_3732);
xor U4359 (N_4359,N_2122,N_3309);
xor U4360 (N_4360,N_2515,N_2771);
xor U4361 (N_4361,N_2903,N_2063);
nand U4362 (N_4362,N_3598,N_2149);
and U4363 (N_4363,N_3779,N_2329);
xnor U4364 (N_4364,N_3218,N_2479);
and U4365 (N_4365,N_3504,N_2253);
and U4366 (N_4366,N_2242,N_2341);
xor U4367 (N_4367,N_2264,N_2534);
xor U4368 (N_4368,N_2163,N_3953);
nor U4369 (N_4369,N_2617,N_3621);
and U4370 (N_4370,N_2304,N_2788);
or U4371 (N_4371,N_3344,N_2780);
or U4372 (N_4372,N_2490,N_3312);
or U4373 (N_4373,N_2574,N_3760);
and U4374 (N_4374,N_2753,N_3252);
nand U4375 (N_4375,N_3110,N_3459);
nor U4376 (N_4376,N_2446,N_2970);
xor U4377 (N_4377,N_3652,N_2347);
and U4378 (N_4378,N_3706,N_3401);
nor U4379 (N_4379,N_3223,N_3534);
xnor U4380 (N_4380,N_3368,N_3265);
and U4381 (N_4381,N_2969,N_3232);
xnor U4382 (N_4382,N_2817,N_2831);
nand U4383 (N_4383,N_3196,N_3973);
and U4384 (N_4384,N_3031,N_2133);
nor U4385 (N_4385,N_3332,N_2451);
and U4386 (N_4386,N_2532,N_2223);
nor U4387 (N_4387,N_2193,N_2160);
nand U4388 (N_4388,N_2703,N_3944);
xor U4389 (N_4389,N_3812,N_3221);
and U4390 (N_4390,N_2793,N_3766);
xnor U4391 (N_4391,N_2404,N_3051);
or U4392 (N_4392,N_2849,N_3915);
or U4393 (N_4393,N_3962,N_3488);
and U4394 (N_4394,N_2670,N_3597);
nand U4395 (N_4395,N_2370,N_2727);
nand U4396 (N_4396,N_3078,N_3450);
nor U4397 (N_4397,N_3097,N_2572);
and U4398 (N_4398,N_3420,N_3900);
nand U4399 (N_4399,N_2482,N_2311);
nand U4400 (N_4400,N_2060,N_2499);
nor U4401 (N_4401,N_3465,N_3311);
nor U4402 (N_4402,N_3228,N_2602);
nor U4403 (N_4403,N_3164,N_2956);
nand U4404 (N_4404,N_3629,N_2147);
nor U4405 (N_4405,N_3909,N_3828);
nor U4406 (N_4406,N_2592,N_3565);
xnor U4407 (N_4407,N_2934,N_3059);
nor U4408 (N_4408,N_3058,N_3718);
xor U4409 (N_4409,N_2386,N_3740);
nand U4410 (N_4410,N_3400,N_3495);
nor U4411 (N_4411,N_2735,N_2525);
nand U4412 (N_4412,N_2493,N_3177);
nor U4413 (N_4413,N_2445,N_2387);
and U4414 (N_4414,N_3340,N_3115);
or U4415 (N_4415,N_2030,N_3184);
and U4416 (N_4416,N_2245,N_2151);
nor U4417 (N_4417,N_2098,N_2449);
nand U4418 (N_4418,N_3617,N_2854);
nor U4419 (N_4419,N_3781,N_3735);
nor U4420 (N_4420,N_2840,N_2176);
nand U4421 (N_4421,N_3198,N_2582);
and U4422 (N_4422,N_2700,N_2167);
nand U4423 (N_4423,N_2924,N_2586);
nand U4424 (N_4424,N_2140,N_2677);
nand U4425 (N_4425,N_3345,N_2138);
xor U4426 (N_4426,N_2575,N_3236);
or U4427 (N_4427,N_3092,N_2873);
xor U4428 (N_4428,N_3318,N_2841);
nor U4429 (N_4429,N_2088,N_3452);
nor U4430 (N_4430,N_2606,N_2294);
nand U4431 (N_4431,N_3468,N_2150);
xnor U4432 (N_4432,N_2252,N_3851);
and U4433 (N_4433,N_2754,N_2014);
xor U4434 (N_4434,N_2680,N_2121);
nor U4435 (N_4435,N_2580,N_3793);
nor U4436 (N_4436,N_2272,N_2565);
or U4437 (N_4437,N_3453,N_2053);
nor U4438 (N_4438,N_3074,N_2200);
or U4439 (N_4439,N_3685,N_2107);
nor U4440 (N_4440,N_2342,N_2385);
xor U4441 (N_4441,N_2403,N_2803);
nand U4442 (N_4442,N_3961,N_2590);
and U4443 (N_4443,N_2380,N_2425);
nand U4444 (N_4444,N_3394,N_3277);
or U4445 (N_4445,N_2845,N_2974);
or U4446 (N_4446,N_2284,N_2607);
or U4447 (N_4447,N_3992,N_2372);
or U4448 (N_4448,N_3319,N_2208);
or U4449 (N_4449,N_3267,N_3731);
and U4450 (N_4450,N_2920,N_2355);
or U4451 (N_4451,N_3291,N_2396);
xor U4452 (N_4452,N_3734,N_3056);
xor U4453 (N_4453,N_3551,N_3077);
nand U4454 (N_4454,N_2480,N_3199);
and U4455 (N_4455,N_3200,N_3126);
or U4456 (N_4456,N_3414,N_3585);
xor U4457 (N_4457,N_2407,N_3040);
xnor U4458 (N_4458,N_2072,N_2367);
xor U4459 (N_4459,N_2212,N_3210);
nand U4460 (N_4460,N_2074,N_3840);
nand U4461 (N_4461,N_3326,N_2975);
and U4462 (N_4462,N_2211,N_3367);
nor U4463 (N_4463,N_2701,N_2373);
xor U4464 (N_4464,N_3076,N_2589);
or U4465 (N_4465,N_3087,N_3375);
nor U4466 (N_4466,N_3811,N_3616);
xnor U4467 (N_4467,N_3632,N_3057);
and U4468 (N_4468,N_2775,N_3125);
nor U4469 (N_4469,N_3671,N_3461);
or U4470 (N_4470,N_2042,N_2344);
and U4471 (N_4471,N_2967,N_2962);
xor U4472 (N_4472,N_3739,N_3073);
nand U4473 (N_4473,N_2201,N_2882);
nand U4474 (N_4474,N_2221,N_3774);
or U4475 (N_4475,N_2043,N_3693);
nor U4476 (N_4476,N_3810,N_2115);
nor U4477 (N_4477,N_3965,N_3528);
xnor U4478 (N_4478,N_3391,N_3243);
xnor U4479 (N_4479,N_2288,N_2762);
or U4480 (N_4480,N_3105,N_2427);
nor U4481 (N_4481,N_3209,N_2600);
and U4482 (N_4482,N_2542,N_3219);
nand U4483 (N_4483,N_2578,N_3007);
or U4484 (N_4484,N_2985,N_3389);
and U4485 (N_4485,N_3026,N_3416);
and U4486 (N_4486,N_3957,N_3522);
xnor U4487 (N_4487,N_3878,N_2973);
xnor U4488 (N_4488,N_2287,N_2937);
or U4489 (N_4489,N_3297,N_3897);
xor U4490 (N_4490,N_2527,N_3624);
and U4491 (N_4491,N_3193,N_2191);
and U4492 (N_4492,N_2501,N_3646);
nand U4493 (N_4493,N_3500,N_3969);
and U4494 (N_4494,N_2862,N_2790);
and U4495 (N_4495,N_2950,N_2022);
or U4496 (N_4496,N_3742,N_3336);
nor U4497 (N_4497,N_3720,N_3321);
nor U4498 (N_4498,N_3281,N_3093);
or U4499 (N_4499,N_3569,N_2987);
xor U4500 (N_4500,N_2932,N_3854);
nand U4501 (N_4501,N_2297,N_3386);
nor U4502 (N_4502,N_2961,N_2000);
nand U4503 (N_4503,N_2334,N_3064);
and U4504 (N_4504,N_2234,N_2876);
nand U4505 (N_4505,N_3021,N_2795);
nand U4506 (N_4506,N_3775,N_2748);
and U4507 (N_4507,N_3467,N_3436);
nand U4508 (N_4508,N_2768,N_3434);
and U4509 (N_4509,N_2587,N_3166);
nor U4510 (N_4510,N_2936,N_3230);
and U4511 (N_4511,N_3727,N_2773);
and U4512 (N_4512,N_2353,N_2838);
nand U4513 (N_4513,N_3168,N_3733);
nand U4514 (N_4514,N_2818,N_3559);
and U4515 (N_4515,N_2172,N_3203);
or U4516 (N_4516,N_2558,N_3778);
nand U4517 (N_4517,N_2752,N_2559);
xor U4518 (N_4518,N_3736,N_2770);
nor U4519 (N_4519,N_3113,N_2174);
xnor U4520 (N_4520,N_2608,N_3278);
or U4521 (N_4521,N_2598,N_2276);
or U4522 (N_4522,N_2938,N_3112);
and U4523 (N_4523,N_2875,N_3489);
nor U4524 (N_4524,N_2410,N_3202);
nand U4525 (N_4525,N_3956,N_3939);
nor U4526 (N_4526,N_2016,N_2414);
and U4527 (N_4527,N_3537,N_3896);
nor U4528 (N_4528,N_3037,N_2857);
or U4529 (N_4529,N_3625,N_2006);
nor U4530 (N_4530,N_3413,N_2584);
nor U4531 (N_4531,N_3138,N_2049);
nor U4532 (N_4532,N_3922,N_3628);
or U4533 (N_4533,N_2433,N_2217);
nand U4534 (N_4534,N_2551,N_3250);
and U4535 (N_4535,N_2687,N_2303);
nor U4536 (N_4536,N_2491,N_3435);
xor U4537 (N_4537,N_3967,N_3395);
and U4538 (N_4538,N_2844,N_2484);
nand U4539 (N_4539,N_3770,N_3379);
nor U4540 (N_4540,N_2463,N_3407);
nand U4541 (N_4541,N_2369,N_3631);
xnor U4542 (N_4542,N_3701,N_3926);
nor U4543 (N_4543,N_2750,N_2397);
or U4544 (N_4544,N_2548,N_3139);
or U4545 (N_4545,N_2343,N_2402);
xor U4546 (N_4546,N_3313,N_2346);
xnor U4547 (N_4547,N_3640,N_2530);
xor U4548 (N_4548,N_3248,N_2886);
or U4549 (N_4549,N_3885,N_2317);
or U4550 (N_4550,N_3325,N_2013);
nand U4551 (N_4551,N_3388,N_2110);
nand U4552 (N_4552,N_3949,N_2298);
and U4553 (N_4553,N_3256,N_2434);
xnor U4554 (N_4554,N_3723,N_3170);
and U4555 (N_4555,N_3874,N_2581);
xor U4556 (N_4556,N_2681,N_2310);
nand U4557 (N_4557,N_3610,N_3014);
nand U4558 (N_4558,N_3704,N_2819);
nand U4559 (N_4559,N_3579,N_3877);
and U4560 (N_4560,N_3269,N_3356);
nand U4561 (N_4561,N_3868,N_3359);
nand U4562 (N_4562,N_3024,N_2037);
or U4563 (N_4563,N_2243,N_2852);
and U4564 (N_4564,N_3859,N_3842);
and U4565 (N_4565,N_3159,N_3427);
xor U4566 (N_4566,N_2627,N_2108);
nor U4567 (N_4567,N_3804,N_3755);
nand U4568 (N_4568,N_3791,N_3662);
nand U4569 (N_4569,N_2207,N_2851);
nand U4570 (N_4570,N_3690,N_3539);
nor U4571 (N_4571,N_3494,N_2996);
nor U4572 (N_4572,N_3132,N_3067);
xor U4573 (N_4573,N_3782,N_3861);
nand U4574 (N_4574,N_2609,N_2702);
nor U4575 (N_4575,N_2159,N_3516);
and U4576 (N_4576,N_3100,N_3759);
and U4577 (N_4577,N_3160,N_3083);
xnor U4578 (N_4578,N_2432,N_2749);
and U4579 (N_4579,N_2802,N_2374);
nor U4580 (N_4580,N_2286,N_2256);
or U4581 (N_4581,N_2697,N_3643);
and U4582 (N_4582,N_3028,N_2268);
nand U4583 (N_4583,N_2505,N_3454);
or U4584 (N_4584,N_3043,N_3938);
and U4585 (N_4585,N_3729,N_2629);
xor U4586 (N_4586,N_3849,N_2073);
nand U4587 (N_4587,N_2077,N_2545);
and U4588 (N_4588,N_2181,N_3930);
nand U4589 (N_4589,N_3208,N_2746);
xor U4590 (N_4590,N_3604,N_3300);
nor U4591 (N_4591,N_2143,N_3809);
or U4592 (N_4592,N_2241,N_3862);
xor U4593 (N_4593,N_3036,N_2436);
nor U4594 (N_4594,N_3020,N_2359);
xnor U4595 (N_4595,N_3481,N_3114);
xor U4596 (N_4596,N_3853,N_3611);
xnor U4597 (N_4597,N_3761,N_3525);
and U4598 (N_4598,N_2518,N_3157);
or U4599 (N_4599,N_2822,N_2325);
nand U4600 (N_4600,N_3238,N_3508);
or U4601 (N_4601,N_2118,N_3355);
nor U4602 (N_4602,N_2126,N_2487);
and U4603 (N_4603,N_2184,N_3829);
nand U4604 (N_4604,N_3806,N_3140);
or U4605 (N_4605,N_3558,N_3052);
nor U4606 (N_4606,N_3103,N_2579);
nor U4607 (N_4607,N_3931,N_2971);
nand U4608 (N_4608,N_2679,N_2027);
nand U4609 (N_4609,N_2196,N_2836);
nand U4610 (N_4610,N_3178,N_2236);
and U4611 (N_4611,N_3233,N_3787);
xor U4612 (N_4612,N_2047,N_3445);
nor U4613 (N_4613,N_2756,N_2483);
nand U4614 (N_4614,N_3712,N_3354);
and U4615 (N_4615,N_3275,N_3290);
or U4616 (N_4616,N_2911,N_3492);
or U4617 (N_4617,N_2827,N_3216);
xnor U4618 (N_4618,N_2759,N_3572);
xor U4619 (N_4619,N_3623,N_3641);
nor U4620 (N_4620,N_2708,N_2005);
nor U4621 (N_4621,N_2597,N_2513);
nand U4622 (N_4622,N_2349,N_2051);
nor U4623 (N_4623,N_2455,N_3310);
nand U4624 (N_4624,N_3654,N_3499);
nand U4625 (N_4625,N_2247,N_2715);
nor U4626 (N_4626,N_2046,N_2056);
nand U4627 (N_4627,N_3645,N_3393);
or U4628 (N_4628,N_2553,N_3180);
nand U4629 (N_4629,N_3669,N_2400);
and U4630 (N_4630,N_2766,N_2123);
nand U4631 (N_4631,N_2250,N_2531);
and U4632 (N_4632,N_2339,N_2716);
nor U4633 (N_4633,N_3315,N_2238);
and U4634 (N_4634,N_2412,N_2357);
nand U4635 (N_4635,N_3323,N_2909);
and U4636 (N_4636,N_2467,N_3392);
xnor U4637 (N_4637,N_3748,N_2129);
and U4638 (N_4638,N_2096,N_2954);
xor U4639 (N_4639,N_3215,N_2659);
xnor U4640 (N_4640,N_2289,N_2719);
xnor U4641 (N_4641,N_2378,N_3426);
nor U4642 (N_4642,N_3270,N_3372);
nand U4643 (N_4643,N_2421,N_2637);
nor U4644 (N_4644,N_2829,N_2540);
or U4645 (N_4645,N_2377,N_2744);
nor U4646 (N_4646,N_3364,N_3482);
xnor U4647 (N_4647,N_3866,N_3993);
nor U4648 (N_4648,N_3602,N_3995);
nor U4649 (N_4649,N_2792,N_2218);
or U4650 (N_4650,N_2454,N_3710);
nand U4651 (N_4651,N_2097,N_2599);
xnor U4652 (N_4652,N_2665,N_3226);
nand U4653 (N_4653,N_2182,N_3703);
nand U4654 (N_4654,N_2782,N_2741);
xnor U4655 (N_4655,N_2384,N_3530);
nand U4656 (N_4656,N_3764,N_3689);
and U4657 (N_4657,N_2492,N_2738);
or U4658 (N_4658,N_3788,N_2651);
xnor U4659 (N_4659,N_3593,N_2278);
nor U4660 (N_4660,N_2448,N_3183);
or U4661 (N_4661,N_2772,N_2919);
nor U4662 (N_4662,N_3022,N_2714);
and U4663 (N_4663,N_3963,N_3813);
xnor U4664 (N_4664,N_2855,N_3924);
or U4665 (N_4665,N_2038,N_2960);
nand U4666 (N_4666,N_3041,N_3133);
xor U4667 (N_4667,N_2424,N_3688);
or U4668 (N_4668,N_2999,N_2834);
nor U4669 (N_4669,N_3999,N_3589);
nor U4670 (N_4670,N_3220,N_3618);
and U4671 (N_4671,N_3936,N_2569);
or U4672 (N_4672,N_3856,N_3990);
nand U4673 (N_4673,N_2251,N_2124);
nand U4674 (N_4674,N_2136,N_2058);
nor U4675 (N_4675,N_2406,N_2833);
or U4676 (N_4676,N_2007,N_3071);
or U4677 (N_4677,N_3274,N_3994);
xor U4678 (N_4678,N_2229,N_2177);
and U4679 (N_4679,N_3769,N_3950);
and U4680 (N_4680,N_3191,N_3514);
or U4681 (N_4681,N_3296,N_3682);
xor U4682 (N_4682,N_3474,N_2319);
nand U4683 (N_4683,N_2336,N_2105);
and U4684 (N_4684,N_2021,N_2997);
or U4685 (N_4685,N_2874,N_2897);
nor U4686 (N_4686,N_2509,N_3423);
or U4687 (N_4687,N_2226,N_2550);
and U4688 (N_4688,N_3753,N_2789);
nand U4689 (N_4689,N_3642,N_3430);
nor U4690 (N_4690,N_2255,N_3398);
or U4691 (N_4691,N_2309,N_2777);
and U4692 (N_4692,N_2225,N_2541);
xnor U4693 (N_4693,N_3425,N_3553);
nand U4694 (N_4694,N_2781,N_2488);
nand U4695 (N_4695,N_2155,N_3343);
nand U4696 (N_4696,N_3082,N_2980);
nor U4697 (N_4697,N_2050,N_3966);
and U4698 (N_4698,N_2417,N_3663);
and U4699 (N_4699,N_2812,N_2120);
xnor U4700 (N_4700,N_2958,N_3061);
xor U4701 (N_4701,N_2682,N_3651);
xor U4702 (N_4702,N_3821,N_2755);
nand U4703 (N_4703,N_2547,N_3987);
or U4704 (N_4704,N_3214,N_2158);
or U4705 (N_4705,N_3172,N_3555);
nor U4706 (N_4706,N_2623,N_3721);
nor U4707 (N_4707,N_2190,N_3229);
xnor U4708 (N_4708,N_2106,N_3916);
and U4709 (N_4709,N_3918,N_3185);
or U4710 (N_4710,N_2718,N_3397);
or U4711 (N_4711,N_3457,N_3008);
or U4712 (N_4712,N_3206,N_2220);
nor U4713 (N_4713,N_2861,N_3545);
and U4714 (N_4714,N_2893,N_2457);
nand U4715 (N_4715,N_3141,N_3797);
nand U4716 (N_4716,N_3342,N_2326);
xor U4717 (N_4717,N_2185,N_3241);
nand U4718 (N_4718,N_3304,N_2688);
xnor U4719 (N_4719,N_3066,N_3405);
or U4720 (N_4720,N_3758,N_3638);
nand U4721 (N_4721,N_2081,N_2720);
xnor U4722 (N_4722,N_3322,N_3512);
nand U4723 (N_4723,N_2751,N_2458);
xor U4724 (N_4724,N_3471,N_2028);
or U4725 (N_4725,N_2824,N_2712);
nor U4726 (N_4726,N_3048,N_3850);
and U4727 (N_4727,N_3947,N_3179);
xor U4728 (N_4728,N_2026,N_2868);
xor U4729 (N_4729,N_3708,N_3044);
nand U4730 (N_4730,N_3786,N_2203);
nor U4731 (N_4731,N_2634,N_2828);
nand U4732 (N_4732,N_3068,N_2514);
and U4733 (N_4733,N_3507,N_3933);
xor U4734 (N_4734,N_3085,N_2791);
nand U4735 (N_4735,N_2065,N_3306);
nand U4736 (N_4736,N_3151,N_2239);
nor U4737 (N_4737,N_3406,N_2621);
and U4738 (N_4738,N_3255,N_2948);
nand U4739 (N_4739,N_2237,N_3819);
nand U4740 (N_4740,N_3365,N_3511);
nand U4741 (N_4741,N_3757,N_3765);
or U4742 (N_4742,N_3574,N_2576);
and U4743 (N_4743,N_2706,N_2604);
or U4744 (N_4744,N_2157,N_3768);
xor U4745 (N_4745,N_2348,N_3283);
nor U4746 (N_4746,N_2486,N_3607);
xor U4747 (N_4747,N_3466,N_3211);
xor U4748 (N_4748,N_2867,N_3901);
nor U4749 (N_4749,N_3741,N_2660);
nand U4750 (N_4750,N_3301,N_3119);
nand U4751 (N_4751,N_2877,N_2371);
and U4752 (N_4752,N_3747,N_2351);
nor U4753 (N_4753,N_3816,N_2995);
and U4754 (N_4754,N_2815,N_2567);
nand U4755 (N_4755,N_2204,N_2045);
nor U4756 (N_4756,N_2327,N_2002);
or U4757 (N_4757,N_3895,N_3668);
and U4758 (N_4758,N_3186,N_2820);
or U4759 (N_4759,N_3111,N_2689);
xnor U4760 (N_4760,N_3042,N_3016);
or U4761 (N_4761,N_3518,N_2536);
xnor U4762 (N_4762,N_2859,N_3134);
and U4763 (N_4763,N_3744,N_3227);
xnor U4764 (N_4764,N_2240,N_3237);
xor U4765 (N_4765,N_3263,N_2908);
nor U4766 (N_4766,N_3412,N_3205);
nor U4767 (N_4767,N_3985,N_2003);
or U4768 (N_4768,N_3135,N_3817);
xnor U4769 (N_4769,N_2048,N_3745);
and U4770 (N_4770,N_2031,N_3377);
nor U4771 (N_4771,N_2690,N_2510);
xor U4772 (N_4772,N_2392,N_2388);
nor U4773 (N_4773,N_2055,N_2267);
or U4774 (N_4774,N_2320,N_3620);
nand U4775 (N_4775,N_3287,N_2331);
nand U4776 (N_4776,N_2091,N_3567);
nand U4777 (N_4777,N_2069,N_2259);
xnor U4778 (N_4778,N_2335,N_3470);
nand U4779 (N_4779,N_2737,N_3971);
xor U4780 (N_4780,N_3143,N_3908);
xor U4781 (N_4781,N_3940,N_3502);
or U4782 (N_4782,N_3677,N_3544);
nor U4783 (N_4783,N_3805,N_2872);
nor U4784 (N_4784,N_3242,N_2142);
nor U4785 (N_4785,N_3664,N_2678);
or U4786 (N_4786,N_2769,N_2645);
nand U4787 (N_4787,N_2981,N_3594);
nand U4788 (N_4788,N_3065,N_3601);
xnor U4789 (N_4789,N_2012,N_3027);
or U4790 (N_4790,N_3098,N_3728);
nand U4791 (N_4791,N_3331,N_3698);
nand U4792 (N_4792,N_3725,N_3547);
or U4793 (N_4793,N_2438,N_2144);
nor U4794 (N_4794,N_3101,N_2544);
xor U4795 (N_4795,N_2931,N_2366);
and U4796 (N_4796,N_2068,N_3003);
xnor U4797 (N_4797,N_2835,N_2656);
nor U4798 (N_4798,N_2549,N_2228);
nand U4799 (N_4799,N_2023,N_3894);
nand U4800 (N_4800,N_2613,N_2774);
or U4801 (N_4801,N_2192,N_2641);
xnor U4802 (N_4802,N_3280,N_3951);
and U4803 (N_4803,N_3906,N_3173);
xnor U4804 (N_4804,N_2935,N_3981);
xor U4805 (N_4805,N_3376,N_3752);
nand U4806 (N_4806,N_2691,N_2156);
nand U4807 (N_4807,N_3167,N_2017);
nand U4808 (N_4808,N_3009,N_2502);
xnor U4809 (N_4809,N_3998,N_2261);
nor U4810 (N_4810,N_3864,N_3724);
xor U4811 (N_4811,N_3285,N_3583);
or U4812 (N_4812,N_2503,N_2308);
xnor U4813 (N_4813,N_3288,N_2776);
or U4814 (N_4814,N_2100,N_3316);
xor U4815 (N_4815,N_2464,N_2794);
and U4816 (N_4816,N_2082,N_3709);
or U4817 (N_4817,N_3437,N_2917);
nor U4818 (N_4818,N_3195,N_3869);
nor U4819 (N_4819,N_3187,N_2148);
and U4820 (N_4820,N_3612,N_3455);
nand U4821 (N_4821,N_2431,N_2519);
nand U4822 (N_4822,N_3972,N_2758);
xnor U4823 (N_4823,N_3552,N_3681);
and U4824 (N_4824,N_2321,N_3959);
nor U4825 (N_4825,N_2556,N_2964);
nor U4826 (N_4826,N_3838,N_2460);
and U4827 (N_4827,N_2942,N_3417);
xor U4828 (N_4828,N_3118,N_2896);
xor U4829 (N_4829,N_3334,N_2989);
nor U4830 (N_4830,N_2473,N_2044);
xor U4831 (N_4831,N_3079,N_2393);
nor U4832 (N_4832,N_3659,N_3674);
nand U4833 (N_4833,N_2178,N_3295);
nor U4834 (N_4834,N_3776,N_3844);
nand U4835 (N_4835,N_2312,N_2508);
xnor U4836 (N_4836,N_3546,N_3108);
and U4837 (N_4837,N_3478,N_3174);
nand U4838 (N_4838,N_2652,N_2632);
nor U4839 (N_4839,N_2895,N_2778);
nand U4840 (N_4840,N_3716,N_2279);
nor U4841 (N_4841,N_2383,N_3827);
nand U4842 (N_4842,N_3580,N_2475);
nor U4843 (N_4843,N_2269,N_3954);
and U4844 (N_4844,N_3655,N_2215);
and U4845 (N_4845,N_3771,N_3307);
or U4846 (N_4846,N_3033,N_3443);
nor U4847 (N_4847,N_3447,N_2616);
or U4848 (N_4848,N_3799,N_2035);
xor U4849 (N_4849,N_3615,N_3475);
xor U4850 (N_4850,N_3192,N_3038);
nor U4851 (N_4851,N_3257,N_3549);
and U4852 (N_4852,N_2564,N_3865);
xnor U4853 (N_4853,N_3245,N_2352);
nand U4854 (N_4854,N_2153,N_2846);
nor U4855 (N_4855,N_3348,N_2843);
and U4856 (N_4856,N_3968,N_3523);
nand U4857 (N_4857,N_2194,N_2639);
nor U4858 (N_4858,N_3751,N_2453);
and U4859 (N_4859,N_2293,N_3702);
or U4860 (N_4860,N_3989,N_3408);
nor U4861 (N_4861,N_2257,N_2865);
nor U4862 (N_4862,N_2189,N_2648);
nor U4863 (N_4863,N_3605,N_3980);
nor U4864 (N_4864,N_2638,N_3231);
and U4865 (N_4865,N_2537,N_2955);
nor U4866 (N_4866,N_3106,N_2991);
or U4867 (N_4867,N_2982,N_2330);
or U4868 (N_4868,N_2905,N_3536);
or U4869 (N_4869,N_3276,N_3235);
xnor U4870 (N_4870,N_2676,N_3484);
nand U4871 (N_4871,N_2356,N_3150);
nand U4872 (N_4872,N_3403,N_2452);
or U4873 (N_4873,N_3460,N_3573);
xnor U4874 (N_4874,N_3449,N_3835);
xor U4875 (N_4875,N_2435,N_3777);
nor U4876 (N_4876,N_3019,N_2628);
nor U4877 (N_4877,N_3303,N_3293);
or U4878 (N_4878,N_2418,N_3772);
and U4879 (N_4879,N_3925,N_3820);
nor U4880 (N_4880,N_3362,N_2663);
xnor U4881 (N_4881,N_3081,N_3353);
xnor U4882 (N_4882,N_2863,N_2270);
xor U4883 (N_4883,N_3201,N_3754);
and U4884 (N_4884,N_2779,N_2314);
nand U4885 (N_4885,N_2061,N_2076);
nor U4886 (N_4886,N_3496,N_2477);
xor U4887 (N_4887,N_2733,N_3415);
and U4888 (N_4888,N_2070,N_3941);
nor U4889 (N_4889,N_2188,N_2554);
xor U4890 (N_4890,N_3259,N_3696);
xor U4891 (N_4891,N_3182,N_2485);
xor U4892 (N_4892,N_3070,N_3730);
and U4893 (N_4893,N_2389,N_2029);
nor U4894 (N_4894,N_2162,N_2067);
or U4895 (N_4895,N_2382,N_2290);
nand U4896 (N_4896,N_2883,N_3142);
or U4897 (N_4897,N_2899,N_3802);
xor U4898 (N_4898,N_3684,N_3948);
xor U4899 (N_4899,N_3661,N_3860);
nand U4900 (N_4900,N_2171,N_3473);
and U4901 (N_4901,N_2057,N_3711);
and U4902 (N_4902,N_2721,N_3418);
nor U4903 (N_4903,N_3576,N_2671);
nor U4904 (N_4904,N_3785,N_3350);
nor U4905 (N_4905,N_2945,N_3714);
nor U4906 (N_4906,N_2470,N_3726);
nand U4907 (N_4907,N_2763,N_2227);
xor U4908 (N_4908,N_3129,N_3349);
or U4909 (N_4909,N_3578,N_2419);
nor U4910 (N_4910,N_2090,N_3145);
nand U4911 (N_4911,N_3845,N_3120);
or U4912 (N_4912,N_2020,N_2137);
nor U4913 (N_4913,N_3509,N_3904);
xor U4914 (N_4914,N_2285,N_3794);
or U4915 (N_4915,N_2340,N_3913);
nand U4916 (N_4916,N_2734,N_2084);
xor U4917 (N_4917,N_3960,N_3834);
nor U4918 (N_4918,N_2596,N_2246);
xor U4919 (N_4919,N_2904,N_2797);
and U4920 (N_4920,N_2811,N_3566);
and U4921 (N_4921,N_2535,N_2739);
nand U4922 (N_4922,N_2302,N_2363);
xnor U4923 (N_4923,N_2807,N_3756);
nor U4924 (N_4924,N_3030,N_2546);
nor U4925 (N_4925,N_3823,N_3049);
nor U4926 (N_4926,N_3039,N_2993);
or U4927 (N_4927,N_3648,N_2032);
xor U4928 (N_4928,N_3004,N_2324);
nor U4929 (N_4929,N_2165,N_3156);
or U4930 (N_4930,N_3692,N_3538);
and U4931 (N_4931,N_2649,N_3366);
nand U4932 (N_4932,N_3683,N_3050);
xor U4933 (N_4933,N_2504,N_2916);
nand U4934 (N_4934,N_2692,N_3251);
or U4935 (N_4935,N_3554,N_2474);
or U4936 (N_4936,N_2538,N_3491);
and U4937 (N_4937,N_2271,N_3128);
nor U4938 (N_4938,N_3880,N_3592);
and U4939 (N_4939,N_2323,N_2856);
xor U4940 (N_4940,N_2570,N_3614);
nor U4941 (N_4941,N_2814,N_3636);
nor U4942 (N_4942,N_2947,N_2101);
or U4943 (N_4943,N_2130,N_3920);
nor U4944 (N_4944,N_2052,N_2742);
xnor U4945 (N_4945,N_2561,N_3352);
nand U4946 (N_4946,N_3626,N_2674);
or U4947 (N_4947,N_3346,N_2249);
nor U4948 (N_4948,N_2506,N_3439);
nor U4949 (N_4949,N_2305,N_3568);
nor U4950 (N_4950,N_3487,N_2978);
nor U4951 (N_4951,N_3564,N_2332);
nand U4952 (N_4952,N_3591,N_2018);
nor U4953 (N_4953,N_3094,N_3562);
or U4954 (N_4954,N_2248,N_3171);
or U4955 (N_4955,N_3421,N_3339);
xor U4956 (N_4956,N_3762,N_3458);
or U4957 (N_4957,N_3109,N_2583);
xnor U4958 (N_4958,N_3207,N_3433);
nand U4959 (N_4959,N_2698,N_2265);
nor U4960 (N_4960,N_2024,N_3271);
nor U4961 (N_4961,N_2760,N_3784);
nand U4962 (N_4962,N_3146,N_3529);
nor U4963 (N_4963,N_2472,N_3234);
nand U4964 (N_4964,N_3676,N_2111);
and U4965 (N_4965,N_2179,N_3535);
nor U4966 (N_4966,N_2089,N_2526);
nand U4967 (N_4967,N_2725,N_2946);
or U4968 (N_4968,N_2630,N_2696);
or U4969 (N_4969,N_3581,N_3596);
nand U4970 (N_4970,N_2095,N_2161);
xnor U4971 (N_4971,N_3390,N_2390);
nand U4972 (N_4972,N_3876,N_2481);
xor U4973 (N_4973,N_3670,N_3883);
xor U4974 (N_4974,N_2104,N_2109);
xor U4975 (N_4975,N_3599,N_2986);
nand U4976 (N_4976,N_3013,N_3749);
nand U4977 (N_4977,N_3675,N_3917);
or U4978 (N_4978,N_2281,N_2837);
and U4979 (N_4979,N_3691,N_3644);
or U4980 (N_4980,N_3996,N_2468);
xor U4981 (N_4981,N_2952,N_3588);
nor U4982 (N_4982,N_3882,N_3839);
xor U4983 (N_4983,N_3130,N_3440);
or U4984 (N_4984,N_3444,N_2723);
and U4985 (N_4985,N_2813,N_3260);
nor U4986 (N_4986,N_2528,N_2131);
xor U4987 (N_4987,N_2033,N_2187);
xor U4988 (N_4988,N_2183,N_3298);
xnor U4989 (N_4989,N_2891,N_3826);
nor U4990 (N_4990,N_3910,N_3062);
nand U4991 (N_4991,N_2260,N_2902);
nand U4992 (N_4992,N_3943,N_2125);
nor U4993 (N_4993,N_3738,N_2657);
nor U4994 (N_4994,N_2180,N_3357);
or U4995 (N_4995,N_2036,N_2809);
xnor U4996 (N_4996,N_2345,N_2889);
nor U4997 (N_4997,N_3658,N_3517);
nor U4998 (N_4998,N_3524,N_3881);
xor U4999 (N_4999,N_3096,N_3988);
and U5000 (N_5000,N_2630,N_2916);
nand U5001 (N_5001,N_3558,N_3231);
nor U5002 (N_5002,N_3928,N_3701);
or U5003 (N_5003,N_3656,N_2097);
xor U5004 (N_5004,N_2863,N_2897);
xor U5005 (N_5005,N_2723,N_3026);
nand U5006 (N_5006,N_2550,N_3764);
xnor U5007 (N_5007,N_2092,N_2811);
and U5008 (N_5008,N_2731,N_2078);
or U5009 (N_5009,N_2889,N_2957);
nor U5010 (N_5010,N_3091,N_3180);
or U5011 (N_5011,N_3254,N_2501);
xnor U5012 (N_5012,N_3122,N_2772);
nor U5013 (N_5013,N_3051,N_2137);
nand U5014 (N_5014,N_2088,N_2030);
or U5015 (N_5015,N_2121,N_2871);
nand U5016 (N_5016,N_3789,N_3330);
or U5017 (N_5017,N_3369,N_3608);
xnor U5018 (N_5018,N_3599,N_2179);
or U5019 (N_5019,N_2990,N_3811);
and U5020 (N_5020,N_2083,N_2442);
and U5021 (N_5021,N_2629,N_2772);
xnor U5022 (N_5022,N_3399,N_3809);
or U5023 (N_5023,N_3616,N_3286);
nor U5024 (N_5024,N_2504,N_3569);
nand U5025 (N_5025,N_2460,N_3925);
nand U5026 (N_5026,N_3873,N_2717);
and U5027 (N_5027,N_2903,N_2960);
nand U5028 (N_5028,N_2494,N_3612);
and U5029 (N_5029,N_2201,N_3391);
nor U5030 (N_5030,N_3335,N_3853);
nor U5031 (N_5031,N_3338,N_3734);
and U5032 (N_5032,N_3164,N_2997);
nand U5033 (N_5033,N_3835,N_2214);
nor U5034 (N_5034,N_2980,N_3635);
and U5035 (N_5035,N_2738,N_2957);
nor U5036 (N_5036,N_3603,N_2790);
nand U5037 (N_5037,N_3941,N_3038);
xor U5038 (N_5038,N_3726,N_3514);
and U5039 (N_5039,N_3123,N_2670);
nor U5040 (N_5040,N_2634,N_3089);
xor U5041 (N_5041,N_3919,N_3465);
nor U5042 (N_5042,N_3412,N_3035);
and U5043 (N_5043,N_3764,N_3117);
xor U5044 (N_5044,N_3035,N_2859);
xnor U5045 (N_5045,N_2587,N_3084);
xor U5046 (N_5046,N_3580,N_3263);
and U5047 (N_5047,N_3734,N_2550);
and U5048 (N_5048,N_2273,N_2492);
xor U5049 (N_5049,N_2957,N_2008);
nor U5050 (N_5050,N_3452,N_2739);
or U5051 (N_5051,N_2504,N_2935);
or U5052 (N_5052,N_2822,N_2873);
or U5053 (N_5053,N_2248,N_3340);
nor U5054 (N_5054,N_2791,N_2417);
or U5055 (N_5055,N_2047,N_3014);
or U5056 (N_5056,N_2075,N_3784);
and U5057 (N_5057,N_3405,N_2196);
and U5058 (N_5058,N_2809,N_3968);
or U5059 (N_5059,N_2498,N_2134);
and U5060 (N_5060,N_2097,N_3600);
nor U5061 (N_5061,N_3578,N_2493);
nand U5062 (N_5062,N_2844,N_2375);
xnor U5063 (N_5063,N_2038,N_3791);
nand U5064 (N_5064,N_2539,N_2871);
xor U5065 (N_5065,N_2650,N_3538);
nand U5066 (N_5066,N_3973,N_2827);
xor U5067 (N_5067,N_3503,N_2053);
or U5068 (N_5068,N_2410,N_2142);
nor U5069 (N_5069,N_3214,N_3478);
xnor U5070 (N_5070,N_2360,N_2749);
nor U5071 (N_5071,N_3050,N_3915);
and U5072 (N_5072,N_2512,N_2901);
xor U5073 (N_5073,N_3696,N_3354);
xnor U5074 (N_5074,N_2310,N_3436);
or U5075 (N_5075,N_3541,N_2140);
or U5076 (N_5076,N_2612,N_3294);
and U5077 (N_5077,N_2705,N_2421);
and U5078 (N_5078,N_3716,N_2646);
or U5079 (N_5079,N_2409,N_3200);
xor U5080 (N_5080,N_3479,N_3119);
xnor U5081 (N_5081,N_2182,N_3112);
xnor U5082 (N_5082,N_3226,N_2219);
and U5083 (N_5083,N_3865,N_2157);
or U5084 (N_5084,N_2853,N_2597);
and U5085 (N_5085,N_2814,N_2572);
nor U5086 (N_5086,N_3974,N_3998);
xnor U5087 (N_5087,N_2201,N_2504);
or U5088 (N_5088,N_2764,N_2188);
nor U5089 (N_5089,N_3496,N_2287);
nor U5090 (N_5090,N_3102,N_2965);
xnor U5091 (N_5091,N_2899,N_2992);
nor U5092 (N_5092,N_2676,N_2034);
or U5093 (N_5093,N_2003,N_2748);
and U5094 (N_5094,N_3404,N_2051);
nor U5095 (N_5095,N_3179,N_3386);
and U5096 (N_5096,N_3322,N_2401);
nor U5097 (N_5097,N_2995,N_2137);
nor U5098 (N_5098,N_3518,N_2366);
nor U5099 (N_5099,N_3633,N_2100);
nand U5100 (N_5100,N_2562,N_2406);
nor U5101 (N_5101,N_3122,N_2092);
or U5102 (N_5102,N_2548,N_2415);
or U5103 (N_5103,N_2902,N_3318);
nor U5104 (N_5104,N_3217,N_2820);
and U5105 (N_5105,N_2825,N_3162);
and U5106 (N_5106,N_2748,N_3807);
or U5107 (N_5107,N_3616,N_3524);
xnor U5108 (N_5108,N_2162,N_2791);
or U5109 (N_5109,N_2231,N_2318);
nor U5110 (N_5110,N_3651,N_2933);
nand U5111 (N_5111,N_3550,N_3562);
and U5112 (N_5112,N_2881,N_2626);
and U5113 (N_5113,N_3619,N_2300);
xnor U5114 (N_5114,N_3867,N_2026);
nor U5115 (N_5115,N_3347,N_2715);
xnor U5116 (N_5116,N_3029,N_2845);
and U5117 (N_5117,N_2124,N_3364);
xnor U5118 (N_5118,N_2023,N_2848);
xor U5119 (N_5119,N_2008,N_2105);
and U5120 (N_5120,N_3515,N_2911);
and U5121 (N_5121,N_3077,N_2193);
nor U5122 (N_5122,N_2869,N_3332);
nor U5123 (N_5123,N_2906,N_2200);
nand U5124 (N_5124,N_3245,N_3521);
nor U5125 (N_5125,N_2065,N_3288);
xnor U5126 (N_5126,N_2911,N_3129);
nor U5127 (N_5127,N_2192,N_2984);
nand U5128 (N_5128,N_2892,N_3423);
nand U5129 (N_5129,N_2821,N_3667);
nor U5130 (N_5130,N_3630,N_2329);
nor U5131 (N_5131,N_3721,N_2330);
nand U5132 (N_5132,N_2156,N_3743);
xor U5133 (N_5133,N_2670,N_2476);
and U5134 (N_5134,N_3735,N_2551);
xnor U5135 (N_5135,N_3854,N_2050);
nor U5136 (N_5136,N_3764,N_2098);
and U5137 (N_5137,N_3751,N_2978);
xor U5138 (N_5138,N_2803,N_2223);
xnor U5139 (N_5139,N_2356,N_3999);
xor U5140 (N_5140,N_3672,N_3540);
xnor U5141 (N_5141,N_2266,N_3949);
and U5142 (N_5142,N_2167,N_3468);
xor U5143 (N_5143,N_3763,N_3666);
nand U5144 (N_5144,N_2510,N_2568);
nand U5145 (N_5145,N_2315,N_3018);
nand U5146 (N_5146,N_3125,N_2643);
nor U5147 (N_5147,N_3282,N_3881);
nand U5148 (N_5148,N_2651,N_3846);
nand U5149 (N_5149,N_2702,N_3677);
xnor U5150 (N_5150,N_3041,N_2567);
xnor U5151 (N_5151,N_2406,N_3822);
and U5152 (N_5152,N_2978,N_2242);
nor U5153 (N_5153,N_2540,N_2883);
and U5154 (N_5154,N_3048,N_3690);
xor U5155 (N_5155,N_3227,N_2569);
nand U5156 (N_5156,N_2847,N_2067);
xor U5157 (N_5157,N_3545,N_2516);
and U5158 (N_5158,N_3756,N_2588);
xnor U5159 (N_5159,N_3768,N_3004);
or U5160 (N_5160,N_2863,N_3463);
nand U5161 (N_5161,N_3475,N_3049);
or U5162 (N_5162,N_3830,N_2135);
xnor U5163 (N_5163,N_2971,N_2995);
xor U5164 (N_5164,N_3440,N_3166);
nand U5165 (N_5165,N_2998,N_3264);
xnor U5166 (N_5166,N_3783,N_3999);
and U5167 (N_5167,N_3585,N_3876);
nor U5168 (N_5168,N_2821,N_2861);
nand U5169 (N_5169,N_2439,N_3122);
nand U5170 (N_5170,N_2617,N_2094);
nand U5171 (N_5171,N_3381,N_2525);
nor U5172 (N_5172,N_2285,N_2453);
nor U5173 (N_5173,N_2939,N_3590);
and U5174 (N_5174,N_3451,N_2326);
xnor U5175 (N_5175,N_2670,N_3313);
or U5176 (N_5176,N_2701,N_2349);
or U5177 (N_5177,N_2916,N_2996);
nor U5178 (N_5178,N_3666,N_3996);
or U5179 (N_5179,N_2483,N_2936);
or U5180 (N_5180,N_3447,N_2781);
or U5181 (N_5181,N_2863,N_2998);
nand U5182 (N_5182,N_3483,N_3470);
and U5183 (N_5183,N_3522,N_3496);
xor U5184 (N_5184,N_2285,N_3657);
and U5185 (N_5185,N_2243,N_3027);
and U5186 (N_5186,N_3270,N_2670);
xor U5187 (N_5187,N_3293,N_3199);
nand U5188 (N_5188,N_2726,N_2299);
nor U5189 (N_5189,N_2628,N_3922);
xnor U5190 (N_5190,N_3336,N_2970);
nor U5191 (N_5191,N_2787,N_3008);
or U5192 (N_5192,N_2466,N_2323);
and U5193 (N_5193,N_2488,N_2927);
and U5194 (N_5194,N_3618,N_3219);
xor U5195 (N_5195,N_2045,N_3050);
or U5196 (N_5196,N_2437,N_3398);
xor U5197 (N_5197,N_3893,N_2693);
and U5198 (N_5198,N_2776,N_3313);
xor U5199 (N_5199,N_3259,N_3834);
nand U5200 (N_5200,N_2934,N_2869);
or U5201 (N_5201,N_3105,N_2587);
nand U5202 (N_5202,N_2334,N_2378);
nor U5203 (N_5203,N_2940,N_3536);
nand U5204 (N_5204,N_3602,N_2051);
nand U5205 (N_5205,N_2827,N_3623);
xor U5206 (N_5206,N_3621,N_2540);
or U5207 (N_5207,N_3803,N_3810);
xor U5208 (N_5208,N_3169,N_2209);
nor U5209 (N_5209,N_2736,N_2025);
nand U5210 (N_5210,N_2934,N_3471);
and U5211 (N_5211,N_3150,N_2447);
xnor U5212 (N_5212,N_2801,N_2964);
nor U5213 (N_5213,N_3116,N_2289);
xor U5214 (N_5214,N_3212,N_3616);
or U5215 (N_5215,N_2883,N_3010);
nand U5216 (N_5216,N_3672,N_2476);
xor U5217 (N_5217,N_2362,N_2172);
or U5218 (N_5218,N_3919,N_3485);
xor U5219 (N_5219,N_3655,N_3008);
or U5220 (N_5220,N_2694,N_2420);
and U5221 (N_5221,N_3553,N_3969);
xor U5222 (N_5222,N_2257,N_2399);
nand U5223 (N_5223,N_2694,N_2818);
nand U5224 (N_5224,N_2010,N_2703);
nand U5225 (N_5225,N_2132,N_2488);
or U5226 (N_5226,N_3466,N_2776);
nand U5227 (N_5227,N_3709,N_2451);
nor U5228 (N_5228,N_3555,N_2747);
nand U5229 (N_5229,N_2035,N_2728);
nand U5230 (N_5230,N_2394,N_3547);
xnor U5231 (N_5231,N_2981,N_3075);
nor U5232 (N_5232,N_3309,N_3198);
and U5233 (N_5233,N_3602,N_3588);
xor U5234 (N_5234,N_2441,N_2800);
nor U5235 (N_5235,N_2263,N_3606);
nor U5236 (N_5236,N_3684,N_3996);
or U5237 (N_5237,N_2667,N_3426);
and U5238 (N_5238,N_3042,N_2750);
or U5239 (N_5239,N_3741,N_2259);
and U5240 (N_5240,N_2011,N_2117);
nor U5241 (N_5241,N_2368,N_3011);
and U5242 (N_5242,N_3174,N_3446);
or U5243 (N_5243,N_3234,N_2437);
xor U5244 (N_5244,N_2060,N_2016);
nor U5245 (N_5245,N_3668,N_2887);
nand U5246 (N_5246,N_2880,N_3239);
nand U5247 (N_5247,N_3771,N_2361);
or U5248 (N_5248,N_3183,N_2380);
or U5249 (N_5249,N_3357,N_3987);
nor U5250 (N_5250,N_3175,N_2357);
nand U5251 (N_5251,N_3325,N_3492);
xor U5252 (N_5252,N_2216,N_3424);
nand U5253 (N_5253,N_2802,N_3239);
nor U5254 (N_5254,N_2273,N_3930);
xor U5255 (N_5255,N_3399,N_2178);
xnor U5256 (N_5256,N_3749,N_3996);
and U5257 (N_5257,N_2169,N_3358);
nor U5258 (N_5258,N_2954,N_3009);
nor U5259 (N_5259,N_2934,N_3080);
nand U5260 (N_5260,N_3261,N_2518);
and U5261 (N_5261,N_3657,N_2436);
or U5262 (N_5262,N_3181,N_2812);
xnor U5263 (N_5263,N_2713,N_3738);
or U5264 (N_5264,N_3258,N_2676);
nand U5265 (N_5265,N_3207,N_3176);
nor U5266 (N_5266,N_3665,N_2968);
and U5267 (N_5267,N_2828,N_2153);
or U5268 (N_5268,N_3269,N_3380);
nand U5269 (N_5269,N_2878,N_2418);
or U5270 (N_5270,N_3373,N_3587);
or U5271 (N_5271,N_3683,N_2305);
xnor U5272 (N_5272,N_3569,N_2559);
nor U5273 (N_5273,N_2406,N_2516);
and U5274 (N_5274,N_2695,N_2509);
nand U5275 (N_5275,N_3801,N_2159);
or U5276 (N_5276,N_2054,N_2399);
xor U5277 (N_5277,N_3522,N_3242);
nor U5278 (N_5278,N_3363,N_2368);
and U5279 (N_5279,N_3412,N_3647);
nand U5280 (N_5280,N_2439,N_3350);
xor U5281 (N_5281,N_3242,N_3714);
and U5282 (N_5282,N_3062,N_3844);
or U5283 (N_5283,N_3499,N_3381);
nor U5284 (N_5284,N_3598,N_3019);
nand U5285 (N_5285,N_3221,N_2158);
or U5286 (N_5286,N_3249,N_2212);
nand U5287 (N_5287,N_3649,N_3710);
or U5288 (N_5288,N_2819,N_3841);
nor U5289 (N_5289,N_3067,N_2141);
xnor U5290 (N_5290,N_3455,N_3573);
xor U5291 (N_5291,N_3430,N_3742);
nor U5292 (N_5292,N_3252,N_3198);
nand U5293 (N_5293,N_2948,N_3120);
nor U5294 (N_5294,N_2508,N_2423);
or U5295 (N_5295,N_2351,N_3385);
nand U5296 (N_5296,N_2229,N_2162);
nor U5297 (N_5297,N_2927,N_3114);
or U5298 (N_5298,N_3539,N_3165);
nand U5299 (N_5299,N_3333,N_3444);
xnor U5300 (N_5300,N_2812,N_2083);
or U5301 (N_5301,N_3593,N_2318);
and U5302 (N_5302,N_2520,N_3145);
or U5303 (N_5303,N_3745,N_2464);
nand U5304 (N_5304,N_3562,N_3758);
nor U5305 (N_5305,N_3115,N_3654);
xor U5306 (N_5306,N_2683,N_2340);
or U5307 (N_5307,N_2884,N_2281);
xor U5308 (N_5308,N_3781,N_3217);
nand U5309 (N_5309,N_3325,N_3673);
nor U5310 (N_5310,N_3473,N_3649);
nand U5311 (N_5311,N_2495,N_3846);
xnor U5312 (N_5312,N_2166,N_3439);
nor U5313 (N_5313,N_2115,N_3704);
xor U5314 (N_5314,N_3065,N_3028);
or U5315 (N_5315,N_2979,N_3494);
nand U5316 (N_5316,N_2202,N_2097);
or U5317 (N_5317,N_3597,N_3779);
nand U5318 (N_5318,N_3402,N_3335);
or U5319 (N_5319,N_3277,N_3840);
xor U5320 (N_5320,N_2227,N_2326);
or U5321 (N_5321,N_3378,N_2148);
or U5322 (N_5322,N_3288,N_3000);
and U5323 (N_5323,N_3823,N_2753);
or U5324 (N_5324,N_3244,N_2568);
or U5325 (N_5325,N_2471,N_3375);
nor U5326 (N_5326,N_2503,N_3635);
or U5327 (N_5327,N_3592,N_3800);
nand U5328 (N_5328,N_2791,N_3781);
and U5329 (N_5329,N_2773,N_2942);
nor U5330 (N_5330,N_2815,N_3773);
and U5331 (N_5331,N_3231,N_2946);
nand U5332 (N_5332,N_2202,N_2086);
nor U5333 (N_5333,N_2499,N_3581);
or U5334 (N_5334,N_3145,N_3193);
nand U5335 (N_5335,N_2478,N_2308);
or U5336 (N_5336,N_3013,N_2577);
xnor U5337 (N_5337,N_2333,N_3350);
xnor U5338 (N_5338,N_2685,N_2925);
xnor U5339 (N_5339,N_3935,N_3466);
or U5340 (N_5340,N_2394,N_2224);
or U5341 (N_5341,N_2290,N_2909);
nand U5342 (N_5342,N_3225,N_2876);
nor U5343 (N_5343,N_2696,N_2889);
nor U5344 (N_5344,N_3597,N_2068);
xnor U5345 (N_5345,N_3779,N_3994);
nor U5346 (N_5346,N_2603,N_2735);
and U5347 (N_5347,N_3715,N_3148);
or U5348 (N_5348,N_3749,N_3561);
and U5349 (N_5349,N_3180,N_2352);
xnor U5350 (N_5350,N_3647,N_2555);
and U5351 (N_5351,N_2565,N_3101);
and U5352 (N_5352,N_2326,N_3821);
nor U5353 (N_5353,N_3049,N_3245);
nor U5354 (N_5354,N_3851,N_2822);
nor U5355 (N_5355,N_2483,N_2959);
xor U5356 (N_5356,N_2336,N_2719);
nor U5357 (N_5357,N_3123,N_2896);
or U5358 (N_5358,N_3209,N_2166);
or U5359 (N_5359,N_3986,N_3450);
nand U5360 (N_5360,N_3121,N_3611);
and U5361 (N_5361,N_3704,N_2756);
or U5362 (N_5362,N_2200,N_3875);
or U5363 (N_5363,N_2558,N_2934);
nor U5364 (N_5364,N_3949,N_2655);
nor U5365 (N_5365,N_2988,N_3162);
xnor U5366 (N_5366,N_2856,N_3201);
and U5367 (N_5367,N_2373,N_3927);
nand U5368 (N_5368,N_3562,N_2435);
and U5369 (N_5369,N_3876,N_3285);
nand U5370 (N_5370,N_2642,N_2004);
xor U5371 (N_5371,N_3232,N_3517);
nor U5372 (N_5372,N_3243,N_3880);
nand U5373 (N_5373,N_3429,N_2760);
and U5374 (N_5374,N_2749,N_3159);
and U5375 (N_5375,N_3033,N_2057);
and U5376 (N_5376,N_2519,N_3645);
xor U5377 (N_5377,N_3371,N_3984);
and U5378 (N_5378,N_2264,N_3044);
nor U5379 (N_5379,N_2667,N_2922);
xor U5380 (N_5380,N_3510,N_3013);
xor U5381 (N_5381,N_2673,N_3911);
nor U5382 (N_5382,N_2975,N_3371);
or U5383 (N_5383,N_2238,N_2990);
xor U5384 (N_5384,N_3340,N_2724);
nand U5385 (N_5385,N_3301,N_3672);
nor U5386 (N_5386,N_2409,N_3079);
nand U5387 (N_5387,N_2463,N_2331);
nand U5388 (N_5388,N_3972,N_3459);
nand U5389 (N_5389,N_2493,N_2187);
or U5390 (N_5390,N_2720,N_3999);
nor U5391 (N_5391,N_3430,N_2884);
xnor U5392 (N_5392,N_3607,N_2506);
nor U5393 (N_5393,N_2772,N_3146);
and U5394 (N_5394,N_2809,N_2735);
xor U5395 (N_5395,N_3071,N_3991);
nand U5396 (N_5396,N_3526,N_3784);
nand U5397 (N_5397,N_3046,N_3917);
and U5398 (N_5398,N_3207,N_2413);
xnor U5399 (N_5399,N_3241,N_3897);
nor U5400 (N_5400,N_3838,N_2436);
xnor U5401 (N_5401,N_2593,N_2891);
or U5402 (N_5402,N_3608,N_2630);
xor U5403 (N_5403,N_2974,N_2864);
nand U5404 (N_5404,N_3534,N_2827);
nor U5405 (N_5405,N_3607,N_2092);
xnor U5406 (N_5406,N_2388,N_2110);
nand U5407 (N_5407,N_2056,N_3593);
xnor U5408 (N_5408,N_3914,N_2054);
xnor U5409 (N_5409,N_3578,N_3755);
xor U5410 (N_5410,N_3918,N_2284);
xnor U5411 (N_5411,N_3124,N_2380);
nor U5412 (N_5412,N_2966,N_3289);
xnor U5413 (N_5413,N_2643,N_2080);
or U5414 (N_5414,N_2628,N_2177);
and U5415 (N_5415,N_2975,N_3503);
xor U5416 (N_5416,N_2817,N_2049);
xnor U5417 (N_5417,N_3835,N_3373);
or U5418 (N_5418,N_2055,N_2888);
and U5419 (N_5419,N_2810,N_3352);
and U5420 (N_5420,N_2730,N_2125);
and U5421 (N_5421,N_2949,N_2340);
or U5422 (N_5422,N_3285,N_2992);
and U5423 (N_5423,N_3006,N_3183);
nor U5424 (N_5424,N_3995,N_2276);
xor U5425 (N_5425,N_2463,N_3198);
and U5426 (N_5426,N_3797,N_2385);
nand U5427 (N_5427,N_2767,N_3761);
xor U5428 (N_5428,N_3771,N_3956);
xnor U5429 (N_5429,N_2758,N_3736);
xor U5430 (N_5430,N_2448,N_3228);
nor U5431 (N_5431,N_3052,N_2113);
and U5432 (N_5432,N_3258,N_2169);
nand U5433 (N_5433,N_2136,N_2440);
nand U5434 (N_5434,N_3976,N_3138);
nand U5435 (N_5435,N_3893,N_3111);
or U5436 (N_5436,N_2703,N_2099);
and U5437 (N_5437,N_3028,N_2289);
or U5438 (N_5438,N_3110,N_3471);
nor U5439 (N_5439,N_3398,N_3783);
nor U5440 (N_5440,N_2086,N_2781);
nand U5441 (N_5441,N_2257,N_2491);
xor U5442 (N_5442,N_3843,N_3523);
and U5443 (N_5443,N_3939,N_3006);
or U5444 (N_5444,N_3260,N_2739);
and U5445 (N_5445,N_2969,N_3906);
and U5446 (N_5446,N_3713,N_3905);
nor U5447 (N_5447,N_2598,N_3754);
nor U5448 (N_5448,N_2137,N_2980);
and U5449 (N_5449,N_2892,N_2260);
or U5450 (N_5450,N_3386,N_3364);
nor U5451 (N_5451,N_2345,N_3821);
or U5452 (N_5452,N_2546,N_3640);
or U5453 (N_5453,N_2605,N_2620);
xnor U5454 (N_5454,N_3264,N_2853);
nand U5455 (N_5455,N_2692,N_3706);
xor U5456 (N_5456,N_3054,N_3485);
nand U5457 (N_5457,N_3405,N_3152);
nor U5458 (N_5458,N_2402,N_2148);
and U5459 (N_5459,N_3167,N_3301);
or U5460 (N_5460,N_3074,N_3213);
xnor U5461 (N_5461,N_2542,N_3973);
and U5462 (N_5462,N_3830,N_3031);
xnor U5463 (N_5463,N_2320,N_3892);
or U5464 (N_5464,N_2157,N_3287);
nand U5465 (N_5465,N_3975,N_2375);
or U5466 (N_5466,N_3317,N_2599);
nand U5467 (N_5467,N_3763,N_3487);
or U5468 (N_5468,N_2888,N_3089);
or U5469 (N_5469,N_3500,N_2408);
nor U5470 (N_5470,N_3243,N_3725);
or U5471 (N_5471,N_3554,N_3621);
or U5472 (N_5472,N_3996,N_2845);
or U5473 (N_5473,N_3025,N_3624);
and U5474 (N_5474,N_3813,N_3205);
nand U5475 (N_5475,N_3512,N_2793);
xor U5476 (N_5476,N_3834,N_3993);
nand U5477 (N_5477,N_3077,N_2799);
nor U5478 (N_5478,N_3451,N_3083);
and U5479 (N_5479,N_3354,N_2045);
xnor U5480 (N_5480,N_3761,N_2277);
and U5481 (N_5481,N_3849,N_3355);
nand U5482 (N_5482,N_3639,N_2763);
or U5483 (N_5483,N_2601,N_2164);
nor U5484 (N_5484,N_2906,N_2688);
nor U5485 (N_5485,N_3914,N_3749);
and U5486 (N_5486,N_3722,N_2826);
or U5487 (N_5487,N_2388,N_2282);
nand U5488 (N_5488,N_2127,N_2039);
and U5489 (N_5489,N_3518,N_3255);
or U5490 (N_5490,N_3875,N_2172);
nor U5491 (N_5491,N_3792,N_2668);
nor U5492 (N_5492,N_2534,N_2383);
nor U5493 (N_5493,N_2811,N_2944);
nor U5494 (N_5494,N_3552,N_2472);
xor U5495 (N_5495,N_3983,N_3865);
or U5496 (N_5496,N_3174,N_3108);
nand U5497 (N_5497,N_2164,N_2525);
xor U5498 (N_5498,N_2993,N_3071);
and U5499 (N_5499,N_3885,N_2618);
and U5500 (N_5500,N_3086,N_3912);
or U5501 (N_5501,N_2484,N_3887);
or U5502 (N_5502,N_3871,N_2000);
or U5503 (N_5503,N_3879,N_3676);
nand U5504 (N_5504,N_2564,N_2016);
or U5505 (N_5505,N_2212,N_3170);
xnor U5506 (N_5506,N_2320,N_2416);
nor U5507 (N_5507,N_2204,N_3908);
and U5508 (N_5508,N_3771,N_3943);
xor U5509 (N_5509,N_3247,N_3109);
nand U5510 (N_5510,N_2183,N_2219);
nor U5511 (N_5511,N_2919,N_2673);
nand U5512 (N_5512,N_3946,N_3416);
or U5513 (N_5513,N_2146,N_2805);
xnor U5514 (N_5514,N_3875,N_2769);
nand U5515 (N_5515,N_2496,N_2598);
nand U5516 (N_5516,N_2876,N_3357);
or U5517 (N_5517,N_3299,N_3861);
nand U5518 (N_5518,N_3638,N_3983);
nand U5519 (N_5519,N_2591,N_2708);
or U5520 (N_5520,N_2041,N_2725);
xnor U5521 (N_5521,N_2821,N_3766);
or U5522 (N_5522,N_3765,N_3506);
xnor U5523 (N_5523,N_3068,N_2985);
and U5524 (N_5524,N_3367,N_2118);
nor U5525 (N_5525,N_2731,N_2830);
nand U5526 (N_5526,N_2008,N_3152);
nor U5527 (N_5527,N_2894,N_3995);
nand U5528 (N_5528,N_3656,N_2089);
nor U5529 (N_5529,N_3592,N_2766);
or U5530 (N_5530,N_2413,N_2290);
or U5531 (N_5531,N_3028,N_2476);
nor U5532 (N_5532,N_3598,N_2116);
nand U5533 (N_5533,N_3242,N_2398);
and U5534 (N_5534,N_3359,N_2637);
xor U5535 (N_5535,N_3693,N_3688);
nand U5536 (N_5536,N_3392,N_3749);
or U5537 (N_5537,N_2774,N_2501);
xor U5538 (N_5538,N_2033,N_2220);
xor U5539 (N_5539,N_3004,N_3554);
nand U5540 (N_5540,N_2635,N_2514);
nand U5541 (N_5541,N_3279,N_2404);
nor U5542 (N_5542,N_2697,N_2132);
and U5543 (N_5543,N_3693,N_2310);
nor U5544 (N_5544,N_3098,N_2229);
or U5545 (N_5545,N_3569,N_2952);
xnor U5546 (N_5546,N_2198,N_2999);
and U5547 (N_5547,N_3818,N_3786);
or U5548 (N_5548,N_3290,N_3332);
nand U5549 (N_5549,N_2150,N_3828);
xor U5550 (N_5550,N_3522,N_3029);
nor U5551 (N_5551,N_2120,N_2792);
or U5552 (N_5552,N_2640,N_3282);
or U5553 (N_5553,N_3185,N_2950);
nor U5554 (N_5554,N_2990,N_2852);
or U5555 (N_5555,N_2129,N_2867);
nor U5556 (N_5556,N_2746,N_3968);
nor U5557 (N_5557,N_2672,N_3562);
nand U5558 (N_5558,N_2561,N_3303);
and U5559 (N_5559,N_2761,N_2021);
nand U5560 (N_5560,N_3248,N_2030);
and U5561 (N_5561,N_3656,N_3345);
xnor U5562 (N_5562,N_2956,N_3003);
nor U5563 (N_5563,N_3950,N_2591);
and U5564 (N_5564,N_3160,N_3837);
and U5565 (N_5565,N_2697,N_3770);
or U5566 (N_5566,N_2234,N_3070);
and U5567 (N_5567,N_3265,N_2261);
nand U5568 (N_5568,N_2046,N_2859);
nor U5569 (N_5569,N_2820,N_2476);
nor U5570 (N_5570,N_2555,N_3380);
nor U5571 (N_5571,N_3768,N_3762);
nor U5572 (N_5572,N_2395,N_3911);
nor U5573 (N_5573,N_3251,N_2971);
nor U5574 (N_5574,N_2100,N_3407);
nand U5575 (N_5575,N_2222,N_3597);
and U5576 (N_5576,N_2019,N_2248);
nor U5577 (N_5577,N_2995,N_2630);
or U5578 (N_5578,N_3840,N_3966);
or U5579 (N_5579,N_2289,N_2535);
xnor U5580 (N_5580,N_3172,N_3407);
and U5581 (N_5581,N_3104,N_2564);
or U5582 (N_5582,N_2140,N_3041);
nor U5583 (N_5583,N_3502,N_2393);
or U5584 (N_5584,N_2717,N_3478);
and U5585 (N_5585,N_3644,N_3104);
xnor U5586 (N_5586,N_3342,N_3759);
nor U5587 (N_5587,N_3591,N_2380);
or U5588 (N_5588,N_2645,N_2469);
nand U5589 (N_5589,N_3172,N_3670);
xnor U5590 (N_5590,N_3622,N_3429);
nor U5591 (N_5591,N_3509,N_2559);
nor U5592 (N_5592,N_2874,N_2228);
nor U5593 (N_5593,N_3681,N_2901);
nand U5594 (N_5594,N_3847,N_2915);
and U5595 (N_5595,N_2507,N_3927);
nor U5596 (N_5596,N_3261,N_2467);
nand U5597 (N_5597,N_3210,N_3460);
nand U5598 (N_5598,N_2188,N_3749);
xnor U5599 (N_5599,N_3754,N_3032);
nand U5600 (N_5600,N_3991,N_2358);
and U5601 (N_5601,N_2519,N_2243);
and U5602 (N_5602,N_3757,N_3269);
and U5603 (N_5603,N_3335,N_3550);
nor U5604 (N_5604,N_2246,N_3052);
or U5605 (N_5605,N_2808,N_2402);
and U5606 (N_5606,N_2434,N_3971);
xor U5607 (N_5607,N_3995,N_3208);
xnor U5608 (N_5608,N_3143,N_3159);
and U5609 (N_5609,N_2904,N_2630);
nand U5610 (N_5610,N_3167,N_3944);
or U5611 (N_5611,N_2097,N_2075);
nor U5612 (N_5612,N_3834,N_2217);
nand U5613 (N_5613,N_2058,N_3529);
nand U5614 (N_5614,N_2175,N_2862);
xnor U5615 (N_5615,N_2534,N_3293);
or U5616 (N_5616,N_2681,N_3934);
nand U5617 (N_5617,N_3877,N_3788);
xor U5618 (N_5618,N_2434,N_3302);
nor U5619 (N_5619,N_3234,N_3506);
or U5620 (N_5620,N_3698,N_3580);
or U5621 (N_5621,N_2981,N_2537);
nor U5622 (N_5622,N_2460,N_3172);
xor U5623 (N_5623,N_2479,N_2161);
or U5624 (N_5624,N_3846,N_3862);
or U5625 (N_5625,N_3589,N_2577);
nand U5626 (N_5626,N_3136,N_3468);
or U5627 (N_5627,N_2855,N_2302);
and U5628 (N_5628,N_2469,N_3849);
nor U5629 (N_5629,N_2572,N_2620);
nor U5630 (N_5630,N_2889,N_2909);
nor U5631 (N_5631,N_2470,N_3208);
nand U5632 (N_5632,N_2015,N_2456);
nor U5633 (N_5633,N_2318,N_3531);
and U5634 (N_5634,N_2798,N_3477);
xor U5635 (N_5635,N_2137,N_2881);
or U5636 (N_5636,N_3013,N_2034);
nor U5637 (N_5637,N_2835,N_2287);
xor U5638 (N_5638,N_3190,N_2538);
nand U5639 (N_5639,N_2168,N_3544);
xnor U5640 (N_5640,N_3806,N_3394);
or U5641 (N_5641,N_3579,N_3640);
or U5642 (N_5642,N_2361,N_2707);
nand U5643 (N_5643,N_3347,N_3145);
nand U5644 (N_5644,N_3687,N_2040);
and U5645 (N_5645,N_2855,N_3035);
nand U5646 (N_5646,N_2316,N_2058);
and U5647 (N_5647,N_2546,N_3082);
nand U5648 (N_5648,N_3494,N_3647);
nand U5649 (N_5649,N_3377,N_3471);
nand U5650 (N_5650,N_3350,N_2327);
nor U5651 (N_5651,N_3313,N_2092);
nor U5652 (N_5652,N_3441,N_3870);
nand U5653 (N_5653,N_3321,N_2726);
nand U5654 (N_5654,N_3589,N_2562);
or U5655 (N_5655,N_2962,N_2482);
nand U5656 (N_5656,N_2033,N_2078);
nand U5657 (N_5657,N_3133,N_2754);
nor U5658 (N_5658,N_2531,N_2577);
or U5659 (N_5659,N_3597,N_2582);
xnor U5660 (N_5660,N_3442,N_2734);
xnor U5661 (N_5661,N_2191,N_2956);
nand U5662 (N_5662,N_2316,N_2368);
and U5663 (N_5663,N_3548,N_3883);
nor U5664 (N_5664,N_2423,N_3472);
or U5665 (N_5665,N_3611,N_2108);
nor U5666 (N_5666,N_2120,N_2569);
nand U5667 (N_5667,N_3528,N_3868);
nand U5668 (N_5668,N_2292,N_2933);
and U5669 (N_5669,N_3377,N_2472);
nor U5670 (N_5670,N_2472,N_2715);
and U5671 (N_5671,N_3689,N_2440);
or U5672 (N_5672,N_2930,N_2561);
xor U5673 (N_5673,N_3060,N_2123);
or U5674 (N_5674,N_3955,N_3729);
and U5675 (N_5675,N_3790,N_2825);
and U5676 (N_5676,N_3244,N_2261);
nor U5677 (N_5677,N_2883,N_3416);
or U5678 (N_5678,N_3447,N_3860);
nor U5679 (N_5679,N_3497,N_3048);
nand U5680 (N_5680,N_3811,N_2870);
nor U5681 (N_5681,N_3246,N_3823);
nand U5682 (N_5682,N_3792,N_3705);
nand U5683 (N_5683,N_2142,N_2832);
and U5684 (N_5684,N_2025,N_3668);
and U5685 (N_5685,N_2681,N_3040);
or U5686 (N_5686,N_3831,N_2683);
or U5687 (N_5687,N_2170,N_2273);
and U5688 (N_5688,N_3635,N_3932);
nor U5689 (N_5689,N_3293,N_2551);
xnor U5690 (N_5690,N_3199,N_2930);
xor U5691 (N_5691,N_3296,N_2087);
and U5692 (N_5692,N_2069,N_3716);
nand U5693 (N_5693,N_3877,N_2817);
and U5694 (N_5694,N_3853,N_2119);
and U5695 (N_5695,N_3848,N_3320);
nand U5696 (N_5696,N_2211,N_3845);
and U5697 (N_5697,N_3829,N_2798);
and U5698 (N_5698,N_2227,N_3476);
nand U5699 (N_5699,N_3434,N_2129);
xor U5700 (N_5700,N_3669,N_3246);
or U5701 (N_5701,N_3011,N_3335);
xnor U5702 (N_5702,N_3082,N_3123);
or U5703 (N_5703,N_2388,N_2762);
or U5704 (N_5704,N_2652,N_3873);
nor U5705 (N_5705,N_3636,N_3245);
nand U5706 (N_5706,N_3522,N_2054);
and U5707 (N_5707,N_2969,N_3828);
and U5708 (N_5708,N_3597,N_2634);
nor U5709 (N_5709,N_2551,N_3640);
nor U5710 (N_5710,N_3291,N_3258);
or U5711 (N_5711,N_2538,N_3789);
and U5712 (N_5712,N_2964,N_3920);
or U5713 (N_5713,N_3200,N_2211);
xnor U5714 (N_5714,N_3069,N_3952);
nand U5715 (N_5715,N_3379,N_3064);
or U5716 (N_5716,N_2525,N_3611);
nor U5717 (N_5717,N_3680,N_3854);
or U5718 (N_5718,N_2970,N_2925);
nor U5719 (N_5719,N_3404,N_2027);
nand U5720 (N_5720,N_2945,N_3058);
or U5721 (N_5721,N_3180,N_2869);
and U5722 (N_5722,N_2043,N_2489);
or U5723 (N_5723,N_3678,N_2763);
xor U5724 (N_5724,N_3090,N_2793);
and U5725 (N_5725,N_2090,N_2509);
xor U5726 (N_5726,N_2342,N_2045);
and U5727 (N_5727,N_3522,N_3446);
nand U5728 (N_5728,N_3356,N_2947);
xnor U5729 (N_5729,N_2335,N_3269);
or U5730 (N_5730,N_3717,N_2627);
nor U5731 (N_5731,N_2343,N_2644);
nor U5732 (N_5732,N_2351,N_2131);
xnor U5733 (N_5733,N_3814,N_2015);
nand U5734 (N_5734,N_2540,N_2534);
nor U5735 (N_5735,N_3140,N_2008);
nand U5736 (N_5736,N_3204,N_2521);
xor U5737 (N_5737,N_2716,N_2969);
nor U5738 (N_5738,N_3089,N_3227);
xnor U5739 (N_5739,N_2586,N_3715);
or U5740 (N_5740,N_3115,N_3069);
nand U5741 (N_5741,N_3155,N_2515);
or U5742 (N_5742,N_3959,N_2252);
xor U5743 (N_5743,N_3386,N_3953);
xor U5744 (N_5744,N_2033,N_2777);
or U5745 (N_5745,N_2568,N_2847);
and U5746 (N_5746,N_3387,N_3776);
or U5747 (N_5747,N_3550,N_2263);
xnor U5748 (N_5748,N_3239,N_3307);
or U5749 (N_5749,N_2749,N_3824);
nand U5750 (N_5750,N_2238,N_3284);
and U5751 (N_5751,N_2805,N_2375);
and U5752 (N_5752,N_3206,N_2304);
nor U5753 (N_5753,N_3027,N_3710);
xor U5754 (N_5754,N_2628,N_3744);
and U5755 (N_5755,N_2698,N_2019);
xnor U5756 (N_5756,N_2709,N_3230);
or U5757 (N_5757,N_3000,N_3845);
xor U5758 (N_5758,N_2253,N_3091);
and U5759 (N_5759,N_2861,N_3230);
xnor U5760 (N_5760,N_2147,N_2239);
nor U5761 (N_5761,N_3883,N_2965);
and U5762 (N_5762,N_3456,N_3226);
and U5763 (N_5763,N_2505,N_3067);
nor U5764 (N_5764,N_3243,N_3323);
nand U5765 (N_5765,N_3181,N_2135);
or U5766 (N_5766,N_3039,N_3829);
or U5767 (N_5767,N_2531,N_2280);
and U5768 (N_5768,N_2048,N_3059);
or U5769 (N_5769,N_3643,N_2285);
nor U5770 (N_5770,N_3677,N_3321);
xnor U5771 (N_5771,N_2378,N_3243);
and U5772 (N_5772,N_3381,N_2527);
xor U5773 (N_5773,N_2995,N_3508);
xnor U5774 (N_5774,N_2520,N_3004);
or U5775 (N_5775,N_2445,N_3284);
nor U5776 (N_5776,N_2440,N_3239);
and U5777 (N_5777,N_2396,N_3191);
nor U5778 (N_5778,N_3461,N_3542);
xnor U5779 (N_5779,N_2841,N_3908);
or U5780 (N_5780,N_3089,N_3077);
nand U5781 (N_5781,N_3885,N_3082);
and U5782 (N_5782,N_3879,N_2767);
or U5783 (N_5783,N_3928,N_3423);
nor U5784 (N_5784,N_2672,N_2330);
and U5785 (N_5785,N_3685,N_2777);
or U5786 (N_5786,N_2102,N_3906);
xor U5787 (N_5787,N_3195,N_3230);
nor U5788 (N_5788,N_2139,N_3816);
nor U5789 (N_5789,N_3754,N_3962);
or U5790 (N_5790,N_3331,N_3142);
xnor U5791 (N_5791,N_3661,N_2700);
nand U5792 (N_5792,N_3150,N_2100);
nor U5793 (N_5793,N_2705,N_2334);
nand U5794 (N_5794,N_3438,N_3174);
nor U5795 (N_5795,N_3879,N_2969);
nand U5796 (N_5796,N_2450,N_2222);
xor U5797 (N_5797,N_3772,N_3691);
xnor U5798 (N_5798,N_2072,N_2922);
or U5799 (N_5799,N_2042,N_3119);
nand U5800 (N_5800,N_2902,N_3946);
xnor U5801 (N_5801,N_3174,N_3437);
nor U5802 (N_5802,N_3792,N_2519);
and U5803 (N_5803,N_3818,N_2250);
or U5804 (N_5804,N_2940,N_3812);
and U5805 (N_5805,N_3329,N_2618);
nor U5806 (N_5806,N_2607,N_2724);
xor U5807 (N_5807,N_2499,N_2774);
nand U5808 (N_5808,N_2627,N_2581);
nand U5809 (N_5809,N_2600,N_3696);
and U5810 (N_5810,N_2927,N_3788);
nand U5811 (N_5811,N_2238,N_3942);
nand U5812 (N_5812,N_3222,N_3635);
nor U5813 (N_5813,N_3394,N_3056);
and U5814 (N_5814,N_3659,N_3921);
xor U5815 (N_5815,N_2151,N_2674);
xor U5816 (N_5816,N_2504,N_3991);
and U5817 (N_5817,N_2208,N_3787);
nand U5818 (N_5818,N_3097,N_3077);
nor U5819 (N_5819,N_2858,N_3331);
xnor U5820 (N_5820,N_2167,N_3255);
nand U5821 (N_5821,N_3678,N_3832);
or U5822 (N_5822,N_3988,N_2795);
nor U5823 (N_5823,N_2674,N_2393);
and U5824 (N_5824,N_2969,N_3426);
and U5825 (N_5825,N_3297,N_3913);
and U5826 (N_5826,N_3343,N_2483);
nor U5827 (N_5827,N_2796,N_2722);
and U5828 (N_5828,N_3596,N_2865);
nand U5829 (N_5829,N_2668,N_2816);
xnor U5830 (N_5830,N_2630,N_2300);
nand U5831 (N_5831,N_2783,N_2558);
nor U5832 (N_5832,N_3653,N_2299);
nand U5833 (N_5833,N_3788,N_3480);
and U5834 (N_5834,N_3853,N_2049);
xnor U5835 (N_5835,N_2505,N_3206);
nor U5836 (N_5836,N_3222,N_3599);
nand U5837 (N_5837,N_3265,N_3547);
xor U5838 (N_5838,N_3388,N_2403);
nand U5839 (N_5839,N_3026,N_3027);
nor U5840 (N_5840,N_2589,N_3141);
nor U5841 (N_5841,N_2347,N_3653);
nor U5842 (N_5842,N_3430,N_3531);
or U5843 (N_5843,N_2537,N_3950);
xnor U5844 (N_5844,N_3047,N_2367);
nand U5845 (N_5845,N_3474,N_2323);
xnor U5846 (N_5846,N_3196,N_2138);
nor U5847 (N_5847,N_2392,N_2134);
or U5848 (N_5848,N_3444,N_2050);
xor U5849 (N_5849,N_3834,N_2836);
xor U5850 (N_5850,N_3209,N_3931);
nand U5851 (N_5851,N_2461,N_2353);
nand U5852 (N_5852,N_3414,N_3070);
nor U5853 (N_5853,N_3655,N_3486);
nor U5854 (N_5854,N_2963,N_3542);
nor U5855 (N_5855,N_3244,N_3486);
and U5856 (N_5856,N_3515,N_2866);
xor U5857 (N_5857,N_2481,N_2512);
xnor U5858 (N_5858,N_3961,N_2400);
xnor U5859 (N_5859,N_2230,N_2027);
xnor U5860 (N_5860,N_3100,N_2849);
or U5861 (N_5861,N_3568,N_2367);
and U5862 (N_5862,N_3375,N_3062);
nor U5863 (N_5863,N_3912,N_3955);
or U5864 (N_5864,N_2260,N_3383);
and U5865 (N_5865,N_2837,N_3884);
nand U5866 (N_5866,N_2043,N_2821);
and U5867 (N_5867,N_2119,N_2207);
nand U5868 (N_5868,N_3160,N_2974);
and U5869 (N_5869,N_3722,N_2851);
or U5870 (N_5870,N_2342,N_2189);
and U5871 (N_5871,N_2243,N_2322);
xnor U5872 (N_5872,N_2737,N_3816);
nor U5873 (N_5873,N_3051,N_2887);
and U5874 (N_5874,N_2781,N_3203);
and U5875 (N_5875,N_2041,N_2347);
nor U5876 (N_5876,N_3342,N_3758);
and U5877 (N_5877,N_2992,N_2481);
or U5878 (N_5878,N_2858,N_2207);
xor U5879 (N_5879,N_3498,N_3617);
and U5880 (N_5880,N_2984,N_3328);
and U5881 (N_5881,N_3162,N_2263);
and U5882 (N_5882,N_3814,N_3094);
and U5883 (N_5883,N_2937,N_2721);
xnor U5884 (N_5884,N_3226,N_2479);
or U5885 (N_5885,N_3154,N_2525);
nor U5886 (N_5886,N_3066,N_3440);
and U5887 (N_5887,N_3086,N_2428);
xnor U5888 (N_5888,N_2244,N_3775);
or U5889 (N_5889,N_3552,N_3565);
nand U5890 (N_5890,N_3724,N_2924);
nand U5891 (N_5891,N_3805,N_3495);
nand U5892 (N_5892,N_3242,N_2730);
nand U5893 (N_5893,N_3981,N_3829);
nand U5894 (N_5894,N_2794,N_3629);
nand U5895 (N_5895,N_2194,N_2327);
nand U5896 (N_5896,N_3373,N_2907);
xnor U5897 (N_5897,N_2549,N_2016);
or U5898 (N_5898,N_2767,N_3619);
and U5899 (N_5899,N_3195,N_3244);
nor U5900 (N_5900,N_3990,N_3285);
xor U5901 (N_5901,N_2515,N_2056);
and U5902 (N_5902,N_3469,N_3033);
nand U5903 (N_5903,N_3723,N_3929);
nor U5904 (N_5904,N_2686,N_3971);
xor U5905 (N_5905,N_2726,N_3163);
and U5906 (N_5906,N_3226,N_3927);
nor U5907 (N_5907,N_3892,N_2586);
or U5908 (N_5908,N_3302,N_2935);
and U5909 (N_5909,N_2955,N_3472);
xor U5910 (N_5910,N_3934,N_3183);
xnor U5911 (N_5911,N_2451,N_3883);
or U5912 (N_5912,N_2053,N_2841);
nor U5913 (N_5913,N_3425,N_3110);
xnor U5914 (N_5914,N_3261,N_2779);
or U5915 (N_5915,N_2994,N_3487);
or U5916 (N_5916,N_3470,N_2108);
and U5917 (N_5917,N_3219,N_2850);
xor U5918 (N_5918,N_2230,N_2330);
or U5919 (N_5919,N_2690,N_2896);
or U5920 (N_5920,N_3986,N_2354);
xnor U5921 (N_5921,N_3619,N_2968);
or U5922 (N_5922,N_3624,N_2415);
and U5923 (N_5923,N_2458,N_2107);
nor U5924 (N_5924,N_2013,N_2290);
and U5925 (N_5925,N_3171,N_3728);
and U5926 (N_5926,N_2226,N_2863);
xnor U5927 (N_5927,N_2574,N_3740);
and U5928 (N_5928,N_3936,N_2612);
nor U5929 (N_5929,N_3686,N_3243);
and U5930 (N_5930,N_2810,N_2271);
or U5931 (N_5931,N_3297,N_3962);
and U5932 (N_5932,N_3045,N_3223);
nand U5933 (N_5933,N_3809,N_3087);
and U5934 (N_5934,N_2476,N_2750);
or U5935 (N_5935,N_3476,N_2525);
nor U5936 (N_5936,N_3456,N_2490);
nand U5937 (N_5937,N_2720,N_3152);
nor U5938 (N_5938,N_3141,N_2631);
xnor U5939 (N_5939,N_2467,N_3243);
and U5940 (N_5940,N_3362,N_3764);
xnor U5941 (N_5941,N_3324,N_2580);
nand U5942 (N_5942,N_3482,N_2740);
nand U5943 (N_5943,N_3327,N_2728);
xnor U5944 (N_5944,N_3762,N_3772);
nand U5945 (N_5945,N_3918,N_3066);
nand U5946 (N_5946,N_3818,N_2517);
or U5947 (N_5947,N_3280,N_3865);
nor U5948 (N_5948,N_2566,N_3769);
or U5949 (N_5949,N_3478,N_3815);
nand U5950 (N_5950,N_2329,N_3979);
xor U5951 (N_5951,N_3208,N_2589);
or U5952 (N_5952,N_3266,N_2012);
nand U5953 (N_5953,N_2701,N_3098);
and U5954 (N_5954,N_2617,N_2107);
xnor U5955 (N_5955,N_2380,N_3108);
nand U5956 (N_5956,N_2984,N_3794);
and U5957 (N_5957,N_3232,N_3090);
nor U5958 (N_5958,N_3190,N_3858);
or U5959 (N_5959,N_3339,N_2034);
and U5960 (N_5960,N_2279,N_2927);
and U5961 (N_5961,N_2068,N_3252);
nand U5962 (N_5962,N_2454,N_2407);
nor U5963 (N_5963,N_2488,N_2472);
nor U5964 (N_5964,N_3906,N_2895);
or U5965 (N_5965,N_3528,N_2796);
nand U5966 (N_5966,N_3826,N_3577);
nor U5967 (N_5967,N_3592,N_2324);
xnor U5968 (N_5968,N_3002,N_2333);
and U5969 (N_5969,N_2842,N_2428);
nor U5970 (N_5970,N_3753,N_3768);
or U5971 (N_5971,N_3368,N_2729);
xor U5972 (N_5972,N_2851,N_3219);
nor U5973 (N_5973,N_2833,N_3910);
and U5974 (N_5974,N_3742,N_3184);
nand U5975 (N_5975,N_2641,N_3864);
nor U5976 (N_5976,N_2444,N_3485);
or U5977 (N_5977,N_3034,N_3159);
nor U5978 (N_5978,N_3269,N_2430);
and U5979 (N_5979,N_2733,N_2090);
and U5980 (N_5980,N_3331,N_2478);
xor U5981 (N_5981,N_2108,N_3315);
nor U5982 (N_5982,N_2517,N_3056);
nand U5983 (N_5983,N_3568,N_2411);
nand U5984 (N_5984,N_2629,N_2693);
nor U5985 (N_5985,N_2346,N_2059);
xor U5986 (N_5986,N_2004,N_3635);
and U5987 (N_5987,N_2500,N_3747);
xnor U5988 (N_5988,N_3366,N_2498);
and U5989 (N_5989,N_3368,N_2809);
xor U5990 (N_5990,N_3004,N_2685);
xor U5991 (N_5991,N_2713,N_3180);
nor U5992 (N_5992,N_2364,N_2587);
nor U5993 (N_5993,N_2238,N_2135);
and U5994 (N_5994,N_2587,N_3857);
xor U5995 (N_5995,N_3571,N_2003);
and U5996 (N_5996,N_2072,N_3288);
nor U5997 (N_5997,N_2640,N_2864);
nor U5998 (N_5998,N_2375,N_2046);
or U5999 (N_5999,N_3737,N_3031);
nand U6000 (N_6000,N_4017,N_5396);
nor U6001 (N_6001,N_4586,N_5145);
xnor U6002 (N_6002,N_4453,N_5244);
xnor U6003 (N_6003,N_5406,N_5685);
and U6004 (N_6004,N_5848,N_4170);
nand U6005 (N_6005,N_4472,N_4108);
xor U6006 (N_6006,N_5492,N_5797);
and U6007 (N_6007,N_4531,N_4340);
xnor U6008 (N_6008,N_4518,N_4358);
nor U6009 (N_6009,N_5552,N_4977);
and U6010 (N_6010,N_5462,N_5193);
xor U6011 (N_6011,N_4437,N_5968);
xnor U6012 (N_6012,N_5743,N_5773);
nand U6013 (N_6013,N_4339,N_5306);
nand U6014 (N_6014,N_5975,N_5718);
and U6015 (N_6015,N_4448,N_4193);
xnor U6016 (N_6016,N_4069,N_4766);
nor U6017 (N_6017,N_5764,N_5084);
xnor U6018 (N_6018,N_4635,N_4229);
xor U6019 (N_6019,N_5576,N_5699);
xnor U6020 (N_6020,N_4738,N_5088);
nand U6021 (N_6021,N_5816,N_4960);
and U6022 (N_6022,N_5787,N_5133);
or U6023 (N_6023,N_5961,N_5886);
and U6024 (N_6024,N_5606,N_4125);
nand U6025 (N_6025,N_5521,N_5143);
or U6026 (N_6026,N_5809,N_4596);
or U6027 (N_6027,N_4407,N_4562);
xor U6028 (N_6028,N_4782,N_5611);
nand U6029 (N_6029,N_4174,N_5030);
xnor U6030 (N_6030,N_4443,N_4599);
or U6031 (N_6031,N_5982,N_5784);
and U6032 (N_6032,N_4754,N_4941);
nor U6033 (N_6033,N_4616,N_5638);
xnor U6034 (N_6034,N_5615,N_5609);
or U6035 (N_6035,N_5694,N_4888);
and U6036 (N_6036,N_4232,N_4601);
nor U6037 (N_6037,N_4580,N_5264);
nor U6038 (N_6038,N_5379,N_4008);
and U6039 (N_6039,N_5367,N_5496);
and U6040 (N_6040,N_5342,N_5977);
or U6041 (N_6041,N_4481,N_4820);
and U6042 (N_6042,N_4041,N_5880);
and U6043 (N_6043,N_4228,N_5417);
and U6044 (N_6044,N_5094,N_4707);
nand U6045 (N_6045,N_5063,N_5973);
nor U6046 (N_6046,N_5838,N_5112);
xnor U6047 (N_6047,N_4483,N_4692);
xor U6048 (N_6048,N_4508,N_4050);
nand U6049 (N_6049,N_4563,N_5987);
nor U6050 (N_6050,N_4642,N_4414);
and U6051 (N_6051,N_5435,N_5043);
nor U6052 (N_6052,N_5467,N_4280);
and U6053 (N_6053,N_4433,N_4020);
and U6054 (N_6054,N_4882,N_4138);
or U6055 (N_6055,N_4537,N_5085);
nor U6056 (N_6056,N_5051,N_5136);
and U6057 (N_6057,N_5339,N_4704);
or U6058 (N_6058,N_5921,N_4348);
nor U6059 (N_6059,N_5994,N_4729);
or U6060 (N_6060,N_5454,N_4083);
or U6061 (N_6061,N_4762,N_5983);
and U6062 (N_6062,N_5356,N_5795);
nor U6063 (N_6063,N_4587,N_5197);
nor U6064 (N_6064,N_4583,N_5794);
nand U6065 (N_6065,N_5905,N_5759);
and U6066 (N_6066,N_4551,N_5411);
nand U6067 (N_6067,N_5668,N_4651);
or U6068 (N_6068,N_5338,N_5506);
and U6069 (N_6069,N_5767,N_4718);
nand U6070 (N_6070,N_5404,N_5386);
and U6071 (N_6071,N_4637,N_4968);
xnor U6072 (N_6072,N_5431,N_5632);
or U6073 (N_6073,N_5045,N_4474);
and U6074 (N_6074,N_4926,N_4073);
nor U6075 (N_6075,N_4102,N_4917);
xnor U6076 (N_6076,N_4655,N_4239);
or U6077 (N_6077,N_5590,N_5532);
or U6078 (N_6078,N_4479,N_5439);
xnor U6079 (N_6079,N_5579,N_5562);
nand U6080 (N_6080,N_5159,N_5249);
nor U6081 (N_6081,N_5783,N_5240);
or U6082 (N_6082,N_5068,N_5670);
nand U6083 (N_6083,N_5660,N_4177);
or U6084 (N_6084,N_4316,N_4090);
xnor U6085 (N_6085,N_5190,N_4952);
or U6086 (N_6086,N_5275,N_4935);
nand U6087 (N_6087,N_5090,N_4029);
nand U6088 (N_6088,N_5598,N_4459);
nand U6089 (N_6089,N_5107,N_5007);
nor U6090 (N_6090,N_5814,N_5432);
nor U6091 (N_6091,N_5387,N_4507);
nor U6092 (N_6092,N_4263,N_4597);
nor U6093 (N_6093,N_4221,N_4406);
and U6094 (N_6094,N_5969,N_5132);
and U6095 (N_6095,N_4304,N_4311);
nor U6096 (N_6096,N_4319,N_4772);
nand U6097 (N_6097,N_5669,N_4268);
and U6098 (N_6098,N_5257,N_4317);
nand U6099 (N_6099,N_4874,N_5942);
nand U6100 (N_6100,N_4261,N_5503);
and U6101 (N_6101,N_4465,N_4609);
and U6102 (N_6102,N_5763,N_5577);
nor U6103 (N_6103,N_4990,N_5057);
nor U6104 (N_6104,N_5839,N_4135);
xnor U6105 (N_6105,N_5989,N_5673);
and U6106 (N_6106,N_5175,N_5074);
nand U6107 (N_6107,N_5913,N_5617);
nor U6108 (N_6108,N_4717,N_5313);
nor U6109 (N_6109,N_5375,N_5681);
xnor U6110 (N_6110,N_4653,N_5399);
nor U6111 (N_6111,N_5164,N_4997);
and U6112 (N_6112,N_4643,N_4678);
or U6113 (N_6113,N_4375,N_4845);
or U6114 (N_6114,N_5587,N_4591);
xnor U6115 (N_6115,N_5285,N_5185);
nand U6116 (N_6116,N_4030,N_4321);
nor U6117 (N_6117,N_5878,N_5234);
nor U6118 (N_6118,N_4190,N_4656);
nand U6119 (N_6119,N_5952,N_4902);
and U6120 (N_6120,N_4638,N_5186);
xnor U6121 (N_6121,N_4257,N_5545);
xor U6122 (N_6122,N_4702,N_4983);
xor U6123 (N_6123,N_4611,N_5173);
nand U6124 (N_6124,N_4040,N_5362);
xnor U6125 (N_6125,N_4359,N_5600);
nand U6126 (N_6126,N_4514,N_4402);
or U6127 (N_6127,N_5607,N_5753);
and U6128 (N_6128,N_4211,N_5591);
or U6129 (N_6129,N_4734,N_4786);
nor U6130 (N_6130,N_4565,N_4958);
xor U6131 (N_6131,N_4356,N_4788);
xor U6132 (N_6132,N_4370,N_5875);
or U6133 (N_6133,N_4844,N_5093);
xor U6134 (N_6134,N_5550,N_5570);
nand U6135 (N_6135,N_5887,N_4490);
xor U6136 (N_6136,N_4632,N_4592);
and U6137 (N_6137,N_4763,N_4188);
nor U6138 (N_6138,N_5423,N_5873);
nand U6139 (N_6139,N_4781,N_4964);
xor U6140 (N_6140,N_5831,N_4155);
or U6141 (N_6141,N_4376,N_4540);
nand U6142 (N_6142,N_5383,N_4818);
and U6143 (N_6143,N_5381,N_5553);
xnor U6144 (N_6144,N_4708,N_4213);
or U6145 (N_6145,N_4975,N_4898);
xor U6146 (N_6146,N_5341,N_5170);
and U6147 (N_6147,N_5284,N_4242);
or U6148 (N_6148,N_5360,N_4741);
xnor U6149 (N_6149,N_5021,N_4189);
or U6150 (N_6150,N_4314,N_5283);
and U6151 (N_6151,N_4233,N_4525);
or U6152 (N_6152,N_4528,N_4372);
or U6153 (N_6153,N_5626,N_5774);
nor U6154 (N_6154,N_5896,N_5274);
and U6155 (N_6155,N_5042,N_4423);
and U6156 (N_6156,N_5930,N_4066);
nand U6157 (N_6157,N_5091,N_4532);
or U6158 (N_6158,N_5298,N_4392);
xnor U6159 (N_6159,N_4595,N_4342);
xor U6160 (N_6160,N_5566,N_5533);
nand U6161 (N_6161,N_4365,N_5189);
nor U6162 (N_6162,N_4493,N_5675);
or U6163 (N_6163,N_4470,N_4825);
xnor U6164 (N_6164,N_5709,N_4993);
or U6165 (N_6165,N_5209,N_5554);
nand U6166 (N_6166,N_5080,N_5293);
nor U6167 (N_6167,N_4087,N_4761);
nor U6168 (N_6168,N_5378,N_5509);
xor U6169 (N_6169,N_5567,N_4224);
or U6170 (N_6170,N_5461,N_4619);
and U6171 (N_6171,N_5314,N_4962);
nand U6172 (N_6172,N_5882,N_4061);
or U6173 (N_6173,N_4693,N_4856);
xor U6174 (N_6174,N_4059,N_4737);
or U6175 (N_6175,N_5004,N_5020);
nand U6176 (N_6176,N_4462,N_4288);
xor U6177 (N_6177,N_4759,N_4456);
or U6178 (N_6178,N_5203,N_5087);
nor U6179 (N_6179,N_5790,N_5912);
nor U6180 (N_6180,N_4581,N_5345);
nor U6181 (N_6181,N_4113,N_5872);
and U6182 (N_6182,N_5624,N_5012);
or U6183 (N_6183,N_4769,N_4875);
nand U6184 (N_6184,N_5546,N_4054);
xor U6185 (N_6185,N_5154,N_4412);
nand U6186 (N_6186,N_5494,N_5514);
or U6187 (N_6187,N_4184,N_4294);
nand U6188 (N_6188,N_5484,N_4223);
xor U6189 (N_6189,N_4285,N_5149);
nand U6190 (N_6190,N_4355,N_5748);
nand U6191 (N_6191,N_5648,N_5499);
nor U6192 (N_6192,N_5118,N_4389);
or U6193 (N_6193,N_5829,N_4833);
nor U6194 (N_6194,N_4264,N_4515);
xnor U6195 (N_6195,N_4298,N_5963);
or U6196 (N_6196,N_5200,N_5967);
nand U6197 (N_6197,N_5822,N_4696);
nor U6198 (N_6198,N_4201,N_4855);
or U6199 (N_6199,N_5206,N_4038);
and U6200 (N_6200,N_4689,N_5895);
or U6201 (N_6201,N_4327,N_4885);
nor U6202 (N_6202,N_4196,N_4700);
xor U6203 (N_6203,N_4909,N_5789);
or U6204 (N_6204,N_4300,N_4396);
or U6205 (N_6205,N_4731,N_4839);
nor U6206 (N_6206,N_5443,N_4053);
nor U6207 (N_6207,N_4683,N_4149);
nand U6208 (N_6208,N_5129,N_5151);
or U6209 (N_6209,N_5254,N_5015);
nand U6210 (N_6210,N_4222,N_5013);
xor U6211 (N_6211,N_4215,N_5819);
and U6212 (N_6212,N_4042,N_4273);
or U6213 (N_6213,N_5978,N_4710);
xor U6214 (N_6214,N_4886,N_4867);
xor U6215 (N_6215,N_5358,N_5294);
nor U6216 (N_6216,N_4585,N_5637);
and U6217 (N_6217,N_5608,N_4668);
and U6218 (N_6218,N_4085,N_5198);
or U6219 (N_6219,N_5561,N_5531);
nand U6220 (N_6220,N_5265,N_5371);
nor U6221 (N_6221,N_4722,N_4837);
or U6222 (N_6222,N_5455,N_5517);
nor U6223 (N_6223,N_5256,N_5440);
and U6224 (N_6224,N_5120,N_5044);
and U6225 (N_6225,N_4594,N_4129);
and U6226 (N_6226,N_4219,N_4203);
or U6227 (N_6227,N_4901,N_4549);
nor U6228 (N_6228,N_5717,N_4492);
and U6229 (N_6229,N_5067,N_5177);
nand U6230 (N_6230,N_5065,N_4613);
xor U6231 (N_6231,N_4614,N_5248);
nor U6232 (N_6232,N_5459,N_5957);
xor U6233 (N_6233,N_4571,N_4714);
xnor U6234 (N_6234,N_5890,N_5772);
nor U6235 (N_6235,N_5923,N_4932);
and U6236 (N_6236,N_4675,N_4842);
xor U6237 (N_6237,N_5158,N_4659);
or U6238 (N_6238,N_4561,N_5216);
or U6239 (N_6239,N_4081,N_4096);
or U6240 (N_6240,N_4421,N_4512);
or U6241 (N_6241,N_4780,N_4186);
xor U6242 (N_6242,N_5938,N_4095);
or U6243 (N_6243,N_4621,N_4441);
or U6244 (N_6244,N_4172,N_5380);
nand U6245 (N_6245,N_5661,N_5867);
nor U6246 (N_6246,N_5179,N_4380);
or U6247 (N_6247,N_5869,N_5102);
and U6248 (N_6248,N_4629,N_5434);
xnor U6249 (N_6249,N_5903,N_5123);
xor U6250 (N_6250,N_5291,N_5866);
or U6251 (N_6251,N_4516,N_4915);
or U6252 (N_6252,N_5894,N_4454);
nor U6253 (N_6253,N_5762,N_5215);
nand U6254 (N_6254,N_5394,N_5370);
nor U6255 (N_6255,N_4214,N_5842);
nand U6256 (N_6256,N_4176,N_5452);
nand U6257 (N_6257,N_4485,N_5061);
and U6258 (N_6258,N_4123,N_5422);
xor U6259 (N_6259,N_4419,N_4422);
or U6260 (N_6260,N_4234,N_5477);
nor U6261 (N_6261,N_5640,N_4226);
nor U6262 (N_6262,N_5560,N_4179);
or U6263 (N_6263,N_5204,N_5498);
nor U6264 (N_6264,N_4691,N_5263);
and U6265 (N_6265,N_4078,N_4953);
and U6266 (N_6266,N_4497,N_4727);
nand U6267 (N_6267,N_4130,N_4310);
nor U6268 (N_6268,N_5747,N_5416);
nor U6269 (N_6269,N_4178,N_5377);
and U6270 (N_6270,N_4084,N_4436);
xnor U6271 (N_6271,N_4256,N_4897);
and U6272 (N_6272,N_5858,N_5098);
xnor U6273 (N_6273,N_4502,N_4185);
xnor U6274 (N_6274,N_5804,N_5701);
nor U6275 (N_6275,N_4559,N_4289);
nand U6276 (N_6276,N_5733,N_5720);
xnor U6277 (N_6277,N_4164,N_5156);
or U6278 (N_6278,N_4891,N_4027);
nand U6279 (N_6279,N_5475,N_5635);
xor U6280 (N_6280,N_4954,N_5742);
nor U6281 (N_6281,N_4980,N_5744);
xnor U6282 (N_6282,N_5716,N_5403);
nor U6283 (N_6283,N_4354,N_4079);
and U6284 (N_6284,N_5205,N_5910);
xnor U6285 (N_6285,N_5280,N_4344);
nand U6286 (N_6286,N_4449,N_4850);
nand U6287 (N_6287,N_4331,N_4431);
and U6288 (N_6288,N_4631,N_4022);
and U6289 (N_6289,N_4854,N_5349);
and U6290 (N_6290,N_4435,N_5137);
xnor U6291 (N_6291,N_5654,N_4978);
nand U6292 (N_6292,N_4959,N_4357);
nand U6293 (N_6293,N_5703,N_5740);
and U6294 (N_6294,N_5334,N_4267);
xnor U6295 (N_6295,N_4471,N_4630);
xnor U6296 (N_6296,N_4403,N_4163);
xnor U6297 (N_6297,N_4663,N_4914);
xnor U6298 (N_6298,N_4152,N_4482);
xnor U6299 (N_6299,N_4701,N_5620);
nor U6300 (N_6300,N_4641,N_4677);
xnor U6301 (N_6301,N_5397,N_4945);
nor U6302 (N_6302,N_4576,N_4005);
nor U6303 (N_6303,N_4814,N_5575);
and U6304 (N_6304,N_5388,N_5233);
nand U6305 (N_6305,N_5052,N_5262);
nand U6306 (N_6306,N_5147,N_4796);
nor U6307 (N_6307,N_4947,N_5195);
xnor U6308 (N_6308,N_5971,N_4416);
nor U6309 (N_6309,N_5428,N_5395);
nor U6310 (N_6310,N_4447,N_5708);
nor U6311 (N_6311,N_4023,N_5005);
xnor U6312 (N_6312,N_4044,N_5039);
or U6313 (N_6313,N_4259,N_5464);
nor U6314 (N_6314,N_5092,N_4861);
or U6315 (N_6315,N_4503,N_5491);
or U6316 (N_6316,N_4265,N_4627);
nand U6317 (N_6317,N_4037,N_5523);
or U6318 (N_6318,N_4341,N_4031);
nand U6319 (N_6319,N_4523,N_4793);
xor U6320 (N_6320,N_5542,N_4863);
nand U6321 (N_6321,N_4021,N_4409);
or U6322 (N_6322,N_5857,N_4120);
nand U6323 (N_6323,N_4753,N_4058);
or U6324 (N_6324,N_4672,N_4987);
and U6325 (N_6325,N_5781,N_5501);
nor U6326 (N_6326,N_5557,N_5730);
and U6327 (N_6327,N_5304,N_4805);
nor U6328 (N_6328,N_4840,N_5722);
nor U6329 (N_6329,N_4200,N_4127);
nand U6330 (N_6330,N_4981,N_5374);
nor U6331 (N_6331,N_5097,N_4440);
nand U6332 (N_6332,N_4929,N_4816);
and U6333 (N_6333,N_5519,N_4679);
nand U6334 (N_6334,N_4415,N_4100);
nand U6335 (N_6335,N_5138,N_5691);
or U6336 (N_6336,N_5172,N_4399);
nand U6337 (N_6337,N_5704,N_5213);
or U6338 (N_6338,N_5146,N_5954);
xor U6339 (N_6339,N_5686,N_4395);
nand U6340 (N_6340,N_4829,N_5430);
and U6341 (N_6341,N_4007,N_5828);
nand U6342 (N_6342,N_5639,N_5934);
xor U6343 (N_6343,N_4122,N_5758);
nand U6344 (N_6344,N_5802,N_4445);
and U6345 (N_6345,N_4556,N_4794);
or U6346 (N_6346,N_4045,N_4384);
or U6347 (N_6347,N_5746,N_4905);
and U6348 (N_6348,N_5415,N_4735);
xor U6349 (N_6349,N_5096,N_4799);
nand U6350 (N_6350,N_4430,N_5832);
xor U6351 (N_6351,N_4171,N_4494);
and U6352 (N_6352,N_4943,N_5674);
xnor U6353 (N_6353,N_4404,N_5425);
nor U6354 (N_6354,N_4862,N_4016);
nand U6355 (N_6355,N_5086,N_5424);
or U6356 (N_6356,N_4831,N_5937);
nand U6357 (N_6357,N_4963,N_4276);
and U6358 (N_6358,N_5518,N_5047);
or U6359 (N_6359,N_5925,N_4938);
xor U6360 (N_6360,N_4104,N_5695);
and U6361 (N_6361,N_4115,N_5226);
xnor U6362 (N_6362,N_5529,N_4382);
or U6363 (N_6363,N_5166,N_5115);
nor U6364 (N_6364,N_4535,N_4721);
and U6365 (N_6365,N_5153,N_4739);
nor U6366 (N_6366,N_5270,N_5319);
xnor U6367 (N_6367,N_5845,N_4032);
nor U6368 (N_6368,N_4680,N_4669);
xor U6369 (N_6369,N_5228,N_4665);
or U6370 (N_6370,N_5757,N_4896);
and U6371 (N_6371,N_4051,N_5142);
or U6372 (N_6372,N_4003,N_4524);
xnor U6373 (N_6373,N_5391,N_5230);
xnor U6374 (N_6374,N_4610,N_5619);
and U6375 (N_6375,N_5412,N_5656);
xnor U6376 (N_6376,N_5444,N_4381);
nand U6377 (N_6377,N_5785,N_4697);
or U6378 (N_6378,N_4520,N_4334);
or U6379 (N_6379,N_4779,N_5864);
and U6380 (N_6380,N_4136,N_4306);
and U6381 (N_6381,N_4690,N_4057);
xor U6382 (N_6382,N_4230,N_4746);
nor U6383 (N_6383,N_4385,N_4284);
xnor U6384 (N_6384,N_4588,N_4579);
or U6385 (N_6385,N_5548,N_5032);
and U6386 (N_6386,N_4967,N_5644);
nor U6387 (N_6387,N_4168,N_5196);
and U6388 (N_6388,N_5486,N_4957);
xnor U6389 (N_6389,N_5534,N_5465);
nor U6390 (N_6390,N_4335,N_4730);
or U6391 (N_6391,N_5229,N_4132);
nand U6392 (N_6392,N_5980,N_5485);
nor U6393 (N_6393,N_5581,N_5410);
and U6394 (N_6394,N_4574,N_5705);
nor U6395 (N_6395,N_5267,N_5595);
xor U6396 (N_6396,N_4353,N_5456);
nand U6397 (N_6397,N_4881,N_5161);
or U6398 (N_6398,N_5109,N_5859);
xnor U6399 (N_6399,N_4103,N_4789);
or U6400 (N_6400,N_4785,N_5614);
and U6401 (N_6401,N_5682,N_5008);
and U6402 (N_6402,N_5944,N_5917);
xor U6403 (N_6403,N_5460,N_5604);
nor U6404 (N_6404,N_4511,N_4329);
or U6405 (N_6405,N_5458,N_4147);
nand U6406 (N_6406,N_5354,N_5336);
and U6407 (N_6407,N_4343,N_5310);
and U6408 (N_6408,N_5837,N_4519);
nor U6409 (N_6409,N_4795,N_5843);
xor U6410 (N_6410,N_5002,N_5128);
nand U6411 (N_6411,N_5208,N_5515);
xnor U6412 (N_6412,N_4347,N_4501);
xnor U6413 (N_6413,N_5337,N_4777);
and U6414 (N_6414,N_5243,N_4352);
nor U6415 (N_6415,N_4169,N_5194);
and U6416 (N_6416,N_5165,N_4877);
or U6417 (N_6417,N_5277,N_4255);
and U6418 (N_6418,N_5418,N_4612);
and U6419 (N_6419,N_4434,N_5066);
nor U6420 (N_6420,N_4913,N_5986);
or U6421 (N_6421,N_5322,N_5863);
xor U6422 (N_6422,N_4950,N_5992);
nor U6423 (N_6423,N_5698,N_4151);
and U6424 (N_6424,N_5621,N_5714);
nand U6425 (N_6425,N_4815,N_5140);
and U6426 (N_6426,N_5076,N_4890);
or U6427 (N_6427,N_4278,N_5888);
xnor U6428 (N_6428,N_5466,N_5827);
or U6429 (N_6429,N_5945,N_4760);
xnor U6430 (N_6430,N_5688,N_4768);
xnor U6431 (N_6431,N_4984,N_5551);
xor U6432 (N_6432,N_5152,N_4249);
nor U6433 (N_6433,N_4802,N_4603);
nand U6434 (N_6434,N_5897,N_4112);
nand U6435 (N_6435,N_5825,N_4645);
and U6436 (N_6436,N_4198,N_5413);
or U6437 (N_6437,N_4145,N_5777);
or U6438 (N_6438,N_5979,N_5671);
and U6439 (N_6439,N_4602,N_4819);
and U6440 (N_6440,N_4332,N_4667);
nand U6441 (N_6441,N_4870,N_5778);
and U6442 (N_6442,N_5811,N_5125);
and U6443 (N_6443,N_5780,N_4615);
xor U6444 (N_6444,N_4397,N_4371);
or U6445 (N_6445,N_5580,N_5988);
nor U6446 (N_6446,N_4828,N_4661);
nand U6447 (N_6447,N_4049,N_5290);
nor U6448 (N_6448,N_5183,N_5317);
nand U6449 (N_6449,N_4992,N_4640);
nand U6450 (N_6450,N_4608,N_4438);
nand U6451 (N_6451,N_5770,N_5592);
nand U6452 (N_6452,N_4047,N_4142);
xnor U6453 (N_6453,N_5959,N_4251);
and U6454 (N_6454,N_4141,N_5003);
or U6455 (N_6455,N_5993,N_4748);
or U6456 (N_6456,N_5719,N_5148);
or U6457 (N_6457,N_4350,N_5715);
or U6458 (N_6458,N_4187,N_4099);
xnor U6459 (N_6459,N_4408,N_5081);
nand U6460 (N_6460,N_5421,N_5711);
xnor U6461 (N_6461,N_4705,N_4270);
and U6462 (N_6462,N_4832,N_4817);
or U6463 (N_6463,N_5525,N_5582);
nor U6464 (N_6464,N_4166,N_5232);
nor U6465 (N_6465,N_5631,N_5818);
nor U6466 (N_6466,N_4773,N_4019);
and U6467 (N_6467,N_4074,N_5224);
nand U6468 (N_6468,N_5260,N_5414);
or U6469 (N_6469,N_4383,N_5732);
nor U6470 (N_6470,N_5451,N_5041);
or U6471 (N_6471,N_5768,N_4067);
xor U6472 (N_6472,N_4377,N_5144);
and U6473 (N_6473,N_5070,N_5801);
nand U6474 (N_6474,N_5726,N_4568);
or U6475 (N_6475,N_5393,N_5850);
and U6476 (N_6476,N_5854,N_4797);
and U6477 (N_6477,N_4143,N_4312);
xnor U6478 (N_6478,N_5347,N_4401);
and U6479 (N_6479,N_4900,N_5181);
nand U6480 (N_6480,N_5479,N_4110);
or U6481 (N_6481,N_5998,N_5218);
and U6482 (N_6482,N_5258,N_4046);
and U6483 (N_6483,N_5390,N_4254);
and U6484 (N_6484,N_4724,N_5756);
or U6485 (N_6485,N_4468,N_5469);
and U6486 (N_6486,N_5255,N_4903);
or U6487 (N_6487,N_5939,N_4320);
nor U6488 (N_6488,N_5572,N_5027);
and U6489 (N_6489,N_4617,N_5006);
or U6490 (N_6490,N_4148,N_5331);
nor U6491 (N_6491,N_4369,N_5713);
nor U6492 (N_6492,N_5078,N_5947);
xor U6493 (N_6493,N_5019,N_4965);
xnor U6494 (N_6494,N_4391,N_4589);
and U6495 (N_6495,N_5826,N_4644);
or U6496 (N_6496,N_5853,N_4486);
nor U6497 (N_6497,N_4813,N_5736);
and U6498 (N_6498,N_5468,N_5680);
nand U6499 (N_6499,N_4106,N_5010);
nand U6500 (N_6500,N_5540,N_4043);
and U6501 (N_6501,N_4681,N_5940);
nor U6502 (N_6502,N_4564,N_4553);
or U6503 (N_6503,N_4252,N_4217);
nand U6504 (N_6504,N_5252,N_5953);
and U6505 (N_6505,N_4158,N_4787);
nand U6506 (N_6506,N_4670,N_4558);
nor U6507 (N_6507,N_5892,N_5936);
nand U6508 (N_6508,N_5364,N_5478);
nand U6509 (N_6509,N_5502,N_4849);
nand U6510 (N_6510,N_4566,N_4250);
xnor U6511 (N_6511,N_4624,N_5900);
xor U6512 (N_6512,N_5559,N_5752);
and U6513 (N_6513,N_4743,N_5805);
and U6514 (N_6514,N_4117,N_5739);
or U6515 (N_6515,N_5798,N_4366);
or U6516 (N_6516,N_4378,N_4363);
nor U6517 (N_6517,N_4134,N_4093);
nand U6518 (N_6518,N_5326,N_5201);
or U6519 (N_6519,N_5271,N_5327);
and U6520 (N_6520,N_4048,N_4277);
or U6521 (N_6521,N_5634,N_4495);
nand U6522 (N_6522,N_5225,N_4544);
and U6523 (N_6523,N_5211,N_5751);
or U6524 (N_6524,N_4025,N_4056);
xnor U6525 (N_6525,N_4181,N_4361);
and U6526 (N_6526,N_5605,N_4985);
xor U6527 (N_6527,N_4970,N_5578);
or U6528 (N_6528,N_4764,N_4065);
nand U6529 (N_6529,N_5035,N_4418);
or U6530 (N_6530,N_5779,N_4400);
nor U6531 (N_6531,N_4694,N_4246);
nand U6532 (N_6532,N_4002,N_4534);
nand U6533 (N_6533,N_5659,N_4077);
nand U6534 (N_6534,N_5647,N_4633);
and U6535 (N_6535,N_4209,N_4427);
nor U6536 (N_6536,N_5569,N_4126);
xnor U6537 (N_6537,N_5909,N_5001);
nand U6538 (N_6538,N_4346,N_5034);
and U6539 (N_6539,N_5966,N_5239);
nand U6540 (N_6540,N_5919,N_4650);
and U6541 (N_6541,N_4039,N_5309);
nor U6542 (N_6542,N_4951,N_4774);
nand U6543 (N_6543,N_4996,N_5769);
nor U6544 (N_6544,N_4824,N_4218);
xor U6545 (N_6545,N_4530,N_4212);
and U6546 (N_6546,N_4550,N_4274);
and U6547 (N_6547,N_4322,N_4974);
nor U6548 (N_6548,N_4823,N_4572);
xor U6549 (N_6549,N_5946,N_5100);
or U6550 (N_6550,N_4119,N_4070);
nor U6551 (N_6551,N_4918,N_4351);
nor U6552 (N_6552,N_5941,N_4308);
nand U6553 (N_6553,N_4387,N_4527);
or U6554 (N_6554,N_5666,N_5613);
nor U6555 (N_6555,N_4736,N_4725);
xor U6556 (N_6556,N_4808,N_5212);
and U6557 (N_6557,N_5792,N_4554);
and U6558 (N_6558,N_4210,N_4182);
nor U6559 (N_6559,N_5622,N_4660);
or U6560 (N_6560,N_5684,N_5602);
or U6561 (N_6561,N_4539,N_5028);
nand U6562 (N_6562,N_4521,N_4933);
xnor U6563 (N_6563,N_5530,N_4349);
xnor U6564 (N_6564,N_5055,N_5861);
xnor U6565 (N_6565,N_4167,N_5250);
nand U6566 (N_6566,N_4208,N_4719);
nand U6567 (N_6567,N_4139,N_4860);
nand U6568 (N_6568,N_4192,N_5970);
xor U6569 (N_6569,N_4060,N_5507);
nand U6570 (N_6570,N_4428,N_4548);
xnor U6571 (N_6571,N_4429,N_4648);
nor U6572 (N_6572,N_5840,N_5541);
nor U6573 (N_6573,N_5246,N_5131);
and U6574 (N_6574,N_5453,N_4751);
nor U6575 (N_6575,N_5806,N_4411);
xor U6576 (N_6576,N_4634,N_4688);
and U6577 (N_6577,N_5723,N_5297);
or U6578 (N_6578,N_4557,N_5236);
nand U6579 (N_6579,N_4712,N_5048);
or U6580 (N_6580,N_5889,N_4000);
or U6581 (N_6581,N_4466,N_5932);
and U6582 (N_6582,N_5497,N_4750);
xnor U6583 (N_6583,N_4988,N_4205);
xnor U6584 (N_6584,N_4153,N_4745);
nor U6585 (N_6585,N_5543,N_4811);
xor U6586 (N_6586,N_5106,N_4150);
nand U6587 (N_6587,N_5821,N_5130);
and U6588 (N_6588,N_4180,N_4865);
nor U6589 (N_6589,N_5544,N_5369);
xor U6590 (N_6590,N_5050,N_4538);
or U6591 (N_6591,N_5108,N_4128);
nor U6592 (N_6592,N_5299,N_5964);
or U6593 (N_6593,N_4241,N_4034);
nand U6594 (N_6594,N_5392,N_5556);
nor U6595 (N_6595,N_5628,N_5121);
or U6596 (N_6596,N_4920,N_5301);
or U6597 (N_6597,N_5365,N_5558);
xor U6598 (N_6598,N_4699,N_5184);
nor U6599 (N_6599,N_4258,N_4244);
or U6600 (N_6600,N_4857,N_5918);
or U6601 (N_6601,N_5536,N_5276);
xor U6602 (N_6602,N_5351,N_4846);
nor U6603 (N_6603,N_5401,N_5646);
nand U6604 (N_6604,N_5101,N_5343);
and U6605 (N_6605,N_5860,N_5064);
nand U6606 (N_6606,N_5564,N_5796);
xor U6607 (N_6607,N_4028,N_5653);
and U6608 (N_6608,N_5655,N_4577);
xor U6609 (N_6609,N_5881,N_5902);
nand U6610 (N_6610,N_4204,N_4243);
or U6611 (N_6611,N_4101,N_5651);
and U6612 (N_6612,N_4080,N_4732);
xor U6613 (N_6613,N_4197,N_4830);
or U6614 (N_6614,N_5357,N_5124);
nor U6615 (N_6615,N_5436,N_4806);
and U6616 (N_6616,N_5813,N_5815);
nand U6617 (N_6617,N_5315,N_4923);
or U6618 (N_6618,N_4292,N_4636);
nand U6619 (N_6619,N_4272,N_5217);
or U6620 (N_6620,N_4904,N_4976);
nor U6621 (N_6621,N_5965,N_5463);
nor U6622 (N_6622,N_4925,N_5000);
and U6623 (N_6623,N_5053,N_4851);
or U6624 (N_6624,N_5474,N_4927);
and U6625 (N_6625,N_4055,N_5584);
nand U6626 (N_6626,N_4140,N_4937);
or U6627 (N_6627,N_5278,N_5366);
nand U6628 (N_6628,N_5191,N_4812);
xnor U6629 (N_6629,N_5835,N_5329);
xnor U6630 (N_6630,N_5836,N_5678);
xnor U6631 (N_6631,N_5915,N_5029);
nor U6632 (N_6632,N_5775,N_5738);
or U6633 (N_6633,N_5931,N_5596);
xor U6634 (N_6634,N_4942,N_5504);
xnor U6635 (N_6635,N_4216,N_4307);
nand U6636 (N_6636,N_4868,N_5171);
or U6637 (N_6637,N_4299,N_5908);
xor U6638 (N_6638,N_5022,N_4500);
nand U6639 (N_6639,N_5237,N_5493);
nand U6640 (N_6640,N_4006,N_4338);
xnor U6641 (N_6641,N_4605,N_5470);
or U6642 (N_6642,N_4859,N_5728);
and U6643 (N_6643,N_5851,N_5450);
and U6644 (N_6644,N_4749,N_4157);
and U6645 (N_6645,N_5024,N_4510);
nor U6646 (N_6646,N_4253,N_4248);
nor U6647 (N_6647,N_5712,N_5117);
xor U6648 (N_6648,N_5817,N_5856);
and U6649 (N_6649,N_5995,N_5725);
and U6650 (N_6650,N_5402,N_5841);
and U6651 (N_6651,N_4676,N_4720);
or U6652 (N_6652,N_5104,N_4469);
nand U6653 (N_6653,N_4309,N_5238);
or U6654 (N_6654,N_5630,N_4068);
and U6655 (N_6655,N_5480,N_5162);
xor U6656 (N_6656,N_4791,N_4607);
or U6657 (N_6657,N_5141,N_5526);
nor U6658 (N_6658,N_4287,N_4426);
and U6659 (N_6659,N_5429,N_5563);
xor U6660 (N_6660,N_5793,N_5420);
or U6661 (N_6661,N_4790,N_4908);
or U6662 (N_6662,N_5981,N_5259);
nand U6663 (N_6663,N_5231,N_5134);
nor U6664 (N_6664,N_5202,N_4262);
or U6665 (N_6665,N_4302,N_4247);
xnor U6666 (N_6666,N_5568,N_5266);
nor U6667 (N_6667,N_5192,N_5235);
or U6668 (N_6668,N_5038,N_5332);
nor U6669 (N_6669,N_4160,N_5261);
xor U6670 (N_6670,N_5707,N_4011);
and U6671 (N_6671,N_5105,N_4698);
nor U6672 (N_6672,N_4852,N_5333);
nor U6673 (N_6673,N_4360,N_5601);
nand U6674 (N_6674,N_5014,N_5033);
nand U6675 (N_6675,N_5160,N_4133);
nand U6676 (N_6676,N_4111,N_5555);
nand U6677 (N_6677,N_4755,N_5885);
nor U6678 (N_6678,N_4803,N_4575);
or U6679 (N_6679,N_5991,N_5683);
and U6680 (N_6680,N_5904,N_5207);
and U6681 (N_6681,N_4345,N_5652);
nand U6682 (N_6682,N_5056,N_4740);
or U6683 (N_6683,N_5693,N_4089);
nand U6684 (N_6684,N_5312,N_5483);
nand U6685 (N_6685,N_5549,N_4420);
and U6686 (N_6686,N_5139,N_5589);
nor U6687 (N_6687,N_5510,N_5812);
nand U6688 (N_6688,N_5924,N_4144);
or U6689 (N_6689,N_5667,N_5448);
nor U6690 (N_6690,N_5537,N_4159);
or U6691 (N_6691,N_4961,N_5956);
xnor U6692 (N_6692,N_5382,N_4014);
nand U6693 (N_6693,N_4162,N_5157);
and U6694 (N_6694,N_4183,N_5490);
nand U6695 (N_6695,N_4063,N_5222);
nor U6696 (N_6696,N_4892,N_5099);
and U6697 (N_6697,N_4315,N_4658);
nand U6698 (N_6698,N_4386,N_4956);
and U6699 (N_6699,N_4245,N_4477);
or U6700 (N_6700,N_5612,N_4673);
and U6701 (N_6701,N_4035,N_5241);
or U6702 (N_6702,N_5922,N_4026);
or U6703 (N_6703,N_5999,N_4505);
nor U6704 (N_6704,N_5352,N_4484);
nor U6705 (N_6705,N_4622,N_5597);
nand U6706 (N_6706,N_4394,N_4807);
or U6707 (N_6707,N_4509,N_4879);
xor U6708 (N_6708,N_4628,N_4944);
nand U6709 (N_6709,N_4646,N_5023);
and U6710 (N_6710,N_5363,N_4517);
xnor U6711 (N_6711,N_4783,N_5176);
nand U6712 (N_6712,N_4569,N_5672);
or U6713 (N_6713,N_4973,N_4955);
xor U6714 (N_6714,N_5482,N_5724);
nor U6715 (N_6715,N_5323,N_4600);
xor U6716 (N_6716,N_5495,N_4086);
xnor U6717 (N_6717,N_4467,N_5389);
nand U6718 (N_6718,N_5223,N_5122);
nor U6719 (N_6719,N_4018,N_5627);
or U6720 (N_6720,N_5408,N_4281);
nand U6721 (N_6721,N_5016,N_5017);
nor U6722 (N_6722,N_5985,N_5799);
nand U6723 (N_6723,N_4297,N_5665);
xor U6724 (N_6724,N_5847,N_5167);
and U6725 (N_6725,N_4652,N_4841);
or U6726 (N_6726,N_4671,N_5618);
nand U6727 (N_6727,N_5928,N_5119);
and U6728 (N_6728,N_5511,N_5512);
nand U6729 (N_6729,N_4013,N_5662);
nor U6730 (N_6730,N_5163,N_5846);
or U6731 (N_6731,N_5700,N_4552);
nand U6732 (N_6732,N_4271,N_4491);
or U6733 (N_6733,N_5155,N_4809);
nor U6734 (N_6734,N_5588,N_4442);
nand U6735 (N_6735,N_5083,N_5227);
nand U6736 (N_6736,N_5346,N_5025);
and U6737 (N_6737,N_4071,N_4094);
or U6738 (N_6738,N_5488,N_5737);
and U6739 (N_6739,N_5676,N_5344);
nor U6740 (N_6740,N_5089,N_4598);
nand U6741 (N_6741,N_4275,N_5874);
or U6742 (N_6742,N_5547,N_5335);
nand U6743 (N_6743,N_4425,N_5891);
nor U6744 (N_6744,N_4895,N_4971);
nand U6745 (N_6745,N_4578,N_4733);
xnor U6746 (N_6746,N_5407,N_5692);
nand U6747 (N_6747,N_4792,N_4206);
nor U6748 (N_6748,N_4478,N_4883);
and U6749 (N_6749,N_5040,N_5282);
nor U6750 (N_6750,N_5075,N_5073);
xnor U6751 (N_6751,N_5800,N_4869);
nand U6752 (N_6752,N_4463,N_5308);
xnor U6753 (N_6753,N_4364,N_5295);
nand U6754 (N_6754,N_4325,N_5750);
xor U6755 (N_6755,N_4894,N_5049);
nand U6756 (N_6756,N_5113,N_5727);
nand U6757 (N_6757,N_5760,N_5318);
nand U6758 (N_6758,N_4716,N_5471);
xor U6759 (N_6759,N_5210,N_5583);
nor U6760 (N_6760,N_5870,N_5616);
nor U6761 (N_6761,N_4473,N_4301);
nor U6762 (N_6762,N_4744,N_5221);
or U6763 (N_6763,N_4328,N_4541);
nand U6764 (N_6764,N_4367,N_5696);
xor U6765 (N_6765,N_4647,N_5990);
or U6766 (N_6766,N_4283,N_4124);
nand U6767 (N_6767,N_5935,N_4506);
nor U6768 (N_6768,N_4237,N_5955);
and U6769 (N_6769,N_5058,N_4620);
nor U6770 (N_6770,N_5437,N_4489);
or U6771 (N_6771,N_4337,N_4880);
xnor U6772 (N_6772,N_5060,N_5522);
or U6773 (N_6773,N_4584,N_5302);
nor U6774 (N_6774,N_4991,N_4618);
or U6775 (N_6775,N_5449,N_5916);
nor U6776 (N_6776,N_5031,N_5731);
xor U6777 (N_6777,N_5062,N_4684);
nor U6778 (N_6778,N_5997,N_5735);
nand U6779 (N_6779,N_5962,N_4723);
and U6780 (N_6780,N_4388,N_5059);
or U6781 (N_6781,N_4362,N_4398);
and U6782 (N_6782,N_4853,N_5405);
nor U6783 (N_6783,N_5710,N_5340);
nand U6784 (N_6784,N_5807,N_4154);
nor U6785 (N_6785,N_5330,N_5893);
xnor U6786 (N_6786,N_5927,N_5741);
or U6787 (N_6787,N_4109,N_5321);
or U6788 (N_6788,N_4015,N_5761);
nor U6789 (N_6789,N_4413,N_4513);
nand U6790 (N_6790,N_5528,N_5328);
nor U6791 (N_6791,N_4199,N_4871);
nand U6792 (N_6792,N_5273,N_5219);
and U6793 (N_6793,N_4800,N_5110);
nand U6794 (N_6794,N_4747,N_4098);
xor U6795 (N_6795,N_5865,N_5348);
nand U6796 (N_6796,N_4269,N_5242);
nand U6797 (N_6797,N_4207,N_4582);
nand U6798 (N_6798,N_5911,N_5324);
and U6799 (N_6799,N_4405,N_5054);
nor U6800 (N_6800,N_4626,N_5585);
xnor U6801 (N_6801,N_4836,N_4775);
nand U6802 (N_6802,N_4457,N_4930);
nor U6803 (N_6803,N_5500,N_4822);
and U6804 (N_6804,N_5481,N_5573);
and U6805 (N_6805,N_4336,N_4165);
nand U6806 (N_6806,N_5879,N_4156);
xnor U6807 (N_6807,N_4887,N_5920);
nor U6808 (N_6808,N_5251,N_5641);
and U6809 (N_6809,N_5303,N_5855);
or U6810 (N_6810,N_5755,N_4662);
nor U6811 (N_6811,N_4533,N_5766);
xnor U6812 (N_6812,N_5359,N_4266);
xor U6813 (N_6813,N_5272,N_4948);
or U6814 (N_6814,N_4279,N_5996);
nor U6815 (N_6815,N_4912,N_4810);
or U6816 (N_6816,N_5446,N_4333);
nor U6817 (N_6817,N_5245,N_4220);
nand U6818 (N_6818,N_4460,N_4480);
and U6819 (N_6819,N_4161,N_4590);
xnor U6820 (N_6820,N_5565,N_5288);
xnor U6821 (N_6821,N_5907,N_4893);
and U6822 (N_6822,N_4009,N_5072);
nor U6823 (N_6823,N_5788,N_4864);
or U6824 (N_6824,N_5754,N_4848);
or U6825 (N_6825,N_5178,N_5508);
and U6826 (N_6826,N_4560,N_4075);
nor U6827 (N_6827,N_5409,N_4703);
and U6828 (N_6828,N_5135,N_4709);
and U6829 (N_6829,N_4326,N_5948);
xor U6830 (N_6830,N_5636,N_5174);
or U6831 (N_6831,N_5095,N_4452);
and U6832 (N_6832,N_4231,N_5026);
xnor U6833 (N_6833,N_4776,N_4062);
nand U6834 (N_6834,N_4374,N_4934);
nor U6835 (N_6835,N_5765,N_5877);
nand U6836 (N_6836,N_4695,N_5269);
xor U6837 (N_6837,N_4173,N_5833);
nor U6838 (N_6838,N_4567,N_5535);
xor U6839 (N_6839,N_4330,N_5823);
xnor U6840 (N_6840,N_4756,N_4238);
and U6841 (N_6841,N_5943,N_5689);
and U6842 (N_6842,N_4546,N_4131);
nand U6843 (N_6843,N_4227,N_5901);
or U6844 (N_6844,N_4911,N_4866);
nand U6845 (N_6845,N_5289,N_4543);
xnor U6846 (N_6846,N_4604,N_4889);
or U6847 (N_6847,N_5657,N_4835);
nor U6848 (N_6848,N_4593,N_4936);
and U6849 (N_6849,N_5871,N_5629);
and U6850 (N_6850,N_5214,N_4969);
nand U6851 (N_6851,N_5745,N_4116);
nor U6852 (N_6852,N_5296,N_4827);
and U6853 (N_6853,N_4107,N_5513);
and U6854 (N_6854,N_4235,N_4092);
and U6855 (N_6855,N_4765,N_4012);
nand U6856 (N_6856,N_5603,N_5782);
and U6857 (N_6857,N_5623,N_5505);
xnor U6858 (N_6858,N_5771,N_5679);
and U6859 (N_6859,N_5253,N_5111);
or U6860 (N_6860,N_4455,N_4393);
nand U6861 (N_6861,N_4982,N_5824);
and U6862 (N_6862,N_5958,N_4488);
and U6863 (N_6863,N_5960,N_5524);
and U6864 (N_6864,N_5126,N_4225);
or U6865 (N_6865,N_5292,N_5687);
nor U6866 (N_6866,N_5011,N_5457);
and U6867 (N_6867,N_4202,N_4994);
and U6868 (N_6868,N_5376,N_4379);
xor U6869 (N_6869,N_4884,N_5844);
xnor U6870 (N_6870,N_5169,N_5372);
nor U6871 (N_6871,N_4052,N_4674);
nor U6872 (N_6872,N_4838,N_4522);
xor U6873 (N_6873,N_5883,N_4946);
or U6874 (N_6874,N_4555,N_4878);
xor U6875 (N_6875,N_5188,N_5187);
xnor U6876 (N_6876,N_5933,N_4303);
and U6877 (N_6877,N_4033,N_5447);
xor U6878 (N_6878,N_5972,N_5642);
nor U6879 (N_6879,N_5664,N_5926);
and U6880 (N_6880,N_4715,N_5082);
nor U6881 (N_6881,N_4072,N_4922);
and U6882 (N_6882,N_4949,N_5729);
xor U6883 (N_6883,N_5079,N_5373);
nand U6884 (N_6884,N_4105,N_4036);
nor U6885 (N_6885,N_5906,N_4010);
or U6886 (N_6886,N_5353,N_4175);
nand U6887 (N_6887,N_5445,N_5114);
nor U6888 (N_6888,N_4476,N_5974);
or U6889 (N_6889,N_4410,N_5810);
or U6890 (N_6890,N_5180,N_4771);
nand U6891 (N_6891,N_4024,N_4450);
nand U6892 (N_6892,N_4498,N_4236);
nor U6893 (N_6893,N_4798,N_4432);
nor U6894 (N_6894,N_5868,N_5116);
and U6895 (N_6895,N_5384,N_4742);
xnor U6896 (N_6896,N_4821,N_4282);
or U6897 (N_6897,N_5527,N_4940);
xnor U6898 (N_6898,N_4475,N_4417);
nand U6899 (N_6899,N_5697,N_4770);
nand U6900 (N_6900,N_4137,N_5476);
xor U6901 (N_6901,N_4623,N_5898);
or U6902 (N_6902,N_5834,N_4114);
and U6903 (N_6903,N_4784,N_4191);
xnor U6904 (N_6904,N_5574,N_4487);
nand U6905 (N_6905,N_4999,N_5803);
nand U6906 (N_6906,N_5037,N_4570);
xnor U6907 (N_6907,N_4757,N_5571);
nor U6908 (N_6908,N_5951,N_4654);
and U6909 (N_6909,N_5441,N_4291);
nor U6910 (N_6910,N_5046,N_4064);
and U6911 (N_6911,N_4664,N_5316);
nand U6912 (N_6912,N_4542,N_4995);
or U6913 (N_6913,N_4972,N_5984);
nor U6914 (N_6914,N_5018,N_5300);
xnor U6915 (N_6915,N_4318,N_4121);
xor U6916 (N_6916,N_5538,N_4464);
nor U6917 (N_6917,N_4872,N_4685);
and U6918 (N_6918,N_5852,N_5199);
nand U6919 (N_6919,N_5586,N_4966);
or U6920 (N_6920,N_5220,N_5643);
or U6921 (N_6921,N_5721,N_5127);
or U6922 (N_6922,N_5438,N_5929);
xor U6923 (N_6923,N_4082,N_5658);
or U6924 (N_6924,N_4686,N_5168);
or U6925 (N_6925,N_4323,N_5305);
and U6926 (N_6926,N_4293,N_5650);
nand U6927 (N_6927,N_5287,N_5976);
nor U6928 (N_6928,N_4924,N_5398);
xnor U6929 (N_6929,N_5649,N_5884);
nor U6930 (N_6930,N_5914,N_4536);
xor U6931 (N_6931,N_4666,N_4313);
or U6932 (N_6932,N_5433,N_4858);
nor U6933 (N_6933,N_4146,N_5268);
and U6934 (N_6934,N_4899,N_4713);
nor U6935 (N_6935,N_4496,N_5663);
and U6936 (N_6936,N_5830,N_4295);
and U6937 (N_6937,N_5281,N_5385);
or U6938 (N_6938,N_4451,N_4916);
xnor U6939 (N_6939,N_4998,N_4986);
or U6940 (N_6940,N_4290,N_4910);
and U6941 (N_6941,N_4439,N_5808);
or U6942 (N_6942,N_5876,N_5355);
xnor U6943 (N_6943,N_5520,N_4657);
xnor U6944 (N_6944,N_4305,N_4921);
and U6945 (N_6945,N_5400,N_5820);
nand U6946 (N_6946,N_5593,N_4876);
and U6947 (N_6947,N_4919,N_5594);
nand U6948 (N_6948,N_5368,N_5036);
nand U6949 (N_6949,N_4778,N_5516);
nor U6950 (N_6950,N_5702,N_4989);
or U6951 (N_6951,N_4001,N_5247);
nor U6952 (N_6952,N_4979,N_4091);
and U6953 (N_6953,N_5786,N_4373);
or U6954 (N_6954,N_5677,N_4804);
and U6955 (N_6955,N_4625,N_4928);
and U6956 (N_6956,N_4728,N_4529);
nand U6957 (N_6957,N_4390,N_5862);
and U6958 (N_6958,N_4834,N_5633);
or U6959 (N_6959,N_4458,N_5307);
nand U6960 (N_6960,N_5426,N_5150);
xor U6961 (N_6961,N_5625,N_4873);
and U6962 (N_6962,N_5286,N_5473);
nand U6963 (N_6963,N_4194,N_4424);
nor U6964 (N_6964,N_5690,N_5009);
and U6965 (N_6965,N_5749,N_5071);
nor U6966 (N_6966,N_5472,N_5610);
and U6967 (N_6967,N_5489,N_4682);
and U6968 (N_6968,N_4649,N_4118);
and U6969 (N_6969,N_5706,N_4843);
nor U6970 (N_6970,N_4296,N_4504);
nand U6971 (N_6971,N_4706,N_4639);
nand U6972 (N_6972,N_4906,N_4939);
xor U6973 (N_6973,N_5325,N_4767);
xnor U6974 (N_6974,N_4286,N_4260);
nor U6975 (N_6975,N_5487,N_5950);
nand U6976 (N_6976,N_5077,N_5320);
xor U6977 (N_6977,N_5419,N_5849);
nand U6978 (N_6978,N_4826,N_4687);
nor U6979 (N_6979,N_4195,N_4499);
and U6980 (N_6980,N_5645,N_5599);
xnor U6981 (N_6981,N_4097,N_5791);
or U6982 (N_6982,N_4240,N_4931);
nand U6983 (N_6983,N_5427,N_5350);
xor U6984 (N_6984,N_5734,N_4461);
or U6985 (N_6985,N_5539,N_5103);
and U6986 (N_6986,N_5182,N_4907);
xnor U6987 (N_6987,N_4004,N_4711);
nand U6988 (N_6988,N_5442,N_5899);
xnor U6989 (N_6989,N_4088,N_4752);
nand U6990 (N_6990,N_4076,N_4726);
and U6991 (N_6991,N_4526,N_5361);
or U6992 (N_6992,N_4446,N_4758);
xnor U6993 (N_6993,N_5776,N_4444);
or U6994 (N_6994,N_4847,N_4547);
nor U6995 (N_6995,N_4545,N_4324);
nor U6996 (N_6996,N_5279,N_4606);
or U6997 (N_6997,N_4573,N_5069);
nor U6998 (N_6998,N_4368,N_4801);
xor U6999 (N_6999,N_5311,N_5949);
xor U7000 (N_7000,N_4800,N_5594);
xnor U7001 (N_7001,N_5942,N_4970);
and U7002 (N_7002,N_4933,N_4024);
nor U7003 (N_7003,N_5647,N_5619);
xor U7004 (N_7004,N_5745,N_5324);
xor U7005 (N_7005,N_5439,N_5491);
nor U7006 (N_7006,N_5169,N_5507);
nand U7007 (N_7007,N_5028,N_5591);
nor U7008 (N_7008,N_4619,N_4945);
nor U7009 (N_7009,N_4018,N_5923);
nor U7010 (N_7010,N_4832,N_4702);
xor U7011 (N_7011,N_4190,N_5494);
nand U7012 (N_7012,N_5601,N_5113);
nor U7013 (N_7013,N_4057,N_4663);
xor U7014 (N_7014,N_4992,N_4893);
and U7015 (N_7015,N_4869,N_5779);
and U7016 (N_7016,N_4691,N_5419);
or U7017 (N_7017,N_5383,N_4015);
or U7018 (N_7018,N_5389,N_5142);
and U7019 (N_7019,N_4946,N_4190);
nor U7020 (N_7020,N_5949,N_5069);
nand U7021 (N_7021,N_4502,N_4235);
nor U7022 (N_7022,N_5598,N_5548);
or U7023 (N_7023,N_5810,N_5504);
xnor U7024 (N_7024,N_5710,N_4297);
and U7025 (N_7025,N_5488,N_5345);
or U7026 (N_7026,N_5588,N_4509);
nand U7027 (N_7027,N_4915,N_4919);
or U7028 (N_7028,N_5115,N_4319);
and U7029 (N_7029,N_5783,N_5060);
xor U7030 (N_7030,N_4732,N_4688);
xnor U7031 (N_7031,N_5639,N_4599);
nand U7032 (N_7032,N_4076,N_4870);
or U7033 (N_7033,N_5672,N_5412);
and U7034 (N_7034,N_4508,N_5072);
nor U7035 (N_7035,N_4235,N_5239);
xnor U7036 (N_7036,N_4948,N_5688);
nand U7037 (N_7037,N_4054,N_4021);
or U7038 (N_7038,N_4622,N_4476);
and U7039 (N_7039,N_4589,N_4475);
and U7040 (N_7040,N_4309,N_4901);
xnor U7041 (N_7041,N_5828,N_4032);
xor U7042 (N_7042,N_5641,N_5421);
xnor U7043 (N_7043,N_4564,N_5099);
or U7044 (N_7044,N_5155,N_4318);
nor U7045 (N_7045,N_5033,N_5626);
or U7046 (N_7046,N_5136,N_5986);
nor U7047 (N_7047,N_4118,N_5861);
and U7048 (N_7048,N_5943,N_4633);
xnor U7049 (N_7049,N_5021,N_5273);
and U7050 (N_7050,N_4066,N_5538);
and U7051 (N_7051,N_5476,N_4835);
and U7052 (N_7052,N_5093,N_5667);
or U7053 (N_7053,N_4313,N_4445);
nor U7054 (N_7054,N_4261,N_5428);
nand U7055 (N_7055,N_4566,N_5831);
nor U7056 (N_7056,N_4940,N_5209);
nor U7057 (N_7057,N_4345,N_5904);
and U7058 (N_7058,N_4192,N_5292);
xnor U7059 (N_7059,N_4090,N_4257);
or U7060 (N_7060,N_5326,N_4651);
and U7061 (N_7061,N_5480,N_4291);
xor U7062 (N_7062,N_5806,N_5054);
or U7063 (N_7063,N_4606,N_4752);
or U7064 (N_7064,N_5600,N_4788);
or U7065 (N_7065,N_4069,N_5519);
and U7066 (N_7066,N_4001,N_4889);
and U7067 (N_7067,N_4706,N_5313);
nor U7068 (N_7068,N_5042,N_4986);
nand U7069 (N_7069,N_4943,N_4012);
or U7070 (N_7070,N_4956,N_4890);
nand U7071 (N_7071,N_4726,N_4179);
nand U7072 (N_7072,N_5993,N_4550);
nand U7073 (N_7073,N_4492,N_4268);
nand U7074 (N_7074,N_4597,N_5289);
nand U7075 (N_7075,N_4200,N_4911);
nand U7076 (N_7076,N_4540,N_5196);
nand U7077 (N_7077,N_4271,N_4102);
and U7078 (N_7078,N_5509,N_4600);
nor U7079 (N_7079,N_4468,N_5712);
nand U7080 (N_7080,N_5785,N_5938);
or U7081 (N_7081,N_5311,N_5337);
nor U7082 (N_7082,N_4117,N_5085);
and U7083 (N_7083,N_5375,N_5632);
and U7084 (N_7084,N_5889,N_4097);
nor U7085 (N_7085,N_4804,N_4732);
and U7086 (N_7086,N_5708,N_5659);
or U7087 (N_7087,N_5023,N_4193);
nor U7088 (N_7088,N_5885,N_5235);
and U7089 (N_7089,N_5842,N_5318);
and U7090 (N_7090,N_4695,N_5698);
xor U7091 (N_7091,N_5037,N_4160);
nand U7092 (N_7092,N_5309,N_5349);
or U7093 (N_7093,N_5639,N_4848);
xnor U7094 (N_7094,N_4574,N_5876);
or U7095 (N_7095,N_4264,N_5086);
xor U7096 (N_7096,N_4988,N_4926);
xor U7097 (N_7097,N_4297,N_4629);
nor U7098 (N_7098,N_5732,N_4074);
xor U7099 (N_7099,N_5393,N_4631);
xor U7100 (N_7100,N_4378,N_4719);
nand U7101 (N_7101,N_4743,N_5021);
or U7102 (N_7102,N_5138,N_5412);
and U7103 (N_7103,N_4355,N_5315);
nand U7104 (N_7104,N_4985,N_5687);
nand U7105 (N_7105,N_5091,N_4812);
nor U7106 (N_7106,N_4174,N_5410);
nor U7107 (N_7107,N_5225,N_4290);
nand U7108 (N_7108,N_4717,N_4959);
nor U7109 (N_7109,N_4825,N_5717);
or U7110 (N_7110,N_5393,N_4307);
or U7111 (N_7111,N_4432,N_4491);
or U7112 (N_7112,N_4348,N_4208);
nor U7113 (N_7113,N_4793,N_4279);
xor U7114 (N_7114,N_4819,N_4001);
xor U7115 (N_7115,N_5410,N_5983);
nor U7116 (N_7116,N_4257,N_4053);
or U7117 (N_7117,N_5361,N_4392);
or U7118 (N_7118,N_5420,N_5113);
and U7119 (N_7119,N_4145,N_4069);
nor U7120 (N_7120,N_4316,N_5382);
and U7121 (N_7121,N_5853,N_5757);
nand U7122 (N_7122,N_4981,N_4495);
or U7123 (N_7123,N_4459,N_4660);
or U7124 (N_7124,N_4866,N_4033);
nand U7125 (N_7125,N_4500,N_5615);
xor U7126 (N_7126,N_5180,N_4306);
and U7127 (N_7127,N_4996,N_4544);
xor U7128 (N_7128,N_5964,N_5763);
nor U7129 (N_7129,N_5803,N_5560);
and U7130 (N_7130,N_5536,N_5398);
or U7131 (N_7131,N_5755,N_4251);
nand U7132 (N_7132,N_5221,N_5476);
and U7133 (N_7133,N_5688,N_5318);
nor U7134 (N_7134,N_5184,N_4431);
nor U7135 (N_7135,N_4260,N_5734);
xnor U7136 (N_7136,N_4392,N_4170);
and U7137 (N_7137,N_4220,N_4539);
and U7138 (N_7138,N_5518,N_5832);
nor U7139 (N_7139,N_4673,N_4897);
or U7140 (N_7140,N_4988,N_5632);
xnor U7141 (N_7141,N_5695,N_4015);
xnor U7142 (N_7142,N_4119,N_4567);
and U7143 (N_7143,N_5398,N_4267);
and U7144 (N_7144,N_4627,N_5601);
and U7145 (N_7145,N_4411,N_4254);
nand U7146 (N_7146,N_4799,N_4332);
xnor U7147 (N_7147,N_4325,N_4994);
nand U7148 (N_7148,N_4168,N_5139);
nor U7149 (N_7149,N_5971,N_4279);
xor U7150 (N_7150,N_5783,N_4054);
xnor U7151 (N_7151,N_4223,N_5040);
nand U7152 (N_7152,N_4780,N_4415);
or U7153 (N_7153,N_4058,N_4807);
xor U7154 (N_7154,N_4665,N_5833);
or U7155 (N_7155,N_5700,N_5431);
or U7156 (N_7156,N_4066,N_4576);
and U7157 (N_7157,N_4425,N_4581);
xnor U7158 (N_7158,N_5844,N_5496);
nand U7159 (N_7159,N_5182,N_4269);
nand U7160 (N_7160,N_4936,N_5956);
or U7161 (N_7161,N_5972,N_5098);
or U7162 (N_7162,N_4497,N_5647);
or U7163 (N_7163,N_4775,N_4081);
or U7164 (N_7164,N_5802,N_4715);
nand U7165 (N_7165,N_5563,N_4565);
nand U7166 (N_7166,N_5577,N_5181);
nor U7167 (N_7167,N_5154,N_4827);
or U7168 (N_7168,N_4501,N_4091);
nor U7169 (N_7169,N_4982,N_4170);
nor U7170 (N_7170,N_4498,N_4564);
xor U7171 (N_7171,N_5296,N_4162);
or U7172 (N_7172,N_4932,N_4174);
or U7173 (N_7173,N_5867,N_5663);
xnor U7174 (N_7174,N_5861,N_5296);
nand U7175 (N_7175,N_4970,N_4918);
xnor U7176 (N_7176,N_4765,N_5214);
and U7177 (N_7177,N_4002,N_5548);
nand U7178 (N_7178,N_4178,N_5057);
nor U7179 (N_7179,N_4714,N_4176);
nor U7180 (N_7180,N_4674,N_5646);
nand U7181 (N_7181,N_5202,N_4115);
or U7182 (N_7182,N_4151,N_5388);
nand U7183 (N_7183,N_4209,N_4031);
or U7184 (N_7184,N_4428,N_5623);
xnor U7185 (N_7185,N_5344,N_5346);
xnor U7186 (N_7186,N_5106,N_5673);
xnor U7187 (N_7187,N_5383,N_5130);
or U7188 (N_7188,N_4862,N_5617);
xnor U7189 (N_7189,N_4917,N_4232);
xnor U7190 (N_7190,N_4748,N_4380);
or U7191 (N_7191,N_4512,N_4632);
nor U7192 (N_7192,N_4777,N_5226);
or U7193 (N_7193,N_5089,N_4930);
nand U7194 (N_7194,N_5700,N_5615);
nor U7195 (N_7195,N_4435,N_4487);
nor U7196 (N_7196,N_5505,N_4578);
xnor U7197 (N_7197,N_5211,N_5277);
xnor U7198 (N_7198,N_5386,N_5506);
nand U7199 (N_7199,N_5136,N_4955);
and U7200 (N_7200,N_4100,N_5002);
or U7201 (N_7201,N_5654,N_5254);
nand U7202 (N_7202,N_4115,N_4031);
or U7203 (N_7203,N_4711,N_4892);
and U7204 (N_7204,N_4667,N_4177);
and U7205 (N_7205,N_4859,N_5773);
and U7206 (N_7206,N_4408,N_4690);
nor U7207 (N_7207,N_5557,N_4634);
xnor U7208 (N_7208,N_4435,N_4511);
or U7209 (N_7209,N_5095,N_4456);
and U7210 (N_7210,N_5652,N_4364);
and U7211 (N_7211,N_5963,N_4296);
nor U7212 (N_7212,N_4610,N_5708);
nor U7213 (N_7213,N_5255,N_5002);
nor U7214 (N_7214,N_5073,N_4375);
nand U7215 (N_7215,N_4378,N_5570);
and U7216 (N_7216,N_4413,N_5642);
nor U7217 (N_7217,N_4704,N_4442);
and U7218 (N_7218,N_4962,N_4356);
nand U7219 (N_7219,N_4118,N_5658);
and U7220 (N_7220,N_4905,N_5680);
xor U7221 (N_7221,N_5780,N_4782);
xor U7222 (N_7222,N_5963,N_4360);
or U7223 (N_7223,N_4472,N_5223);
xor U7224 (N_7224,N_5395,N_5331);
nor U7225 (N_7225,N_4584,N_4386);
xnor U7226 (N_7226,N_5230,N_4661);
xnor U7227 (N_7227,N_5970,N_5815);
nor U7228 (N_7228,N_4853,N_5411);
xor U7229 (N_7229,N_5883,N_5767);
xnor U7230 (N_7230,N_5375,N_5733);
nand U7231 (N_7231,N_4686,N_5951);
xor U7232 (N_7232,N_4885,N_4581);
nor U7233 (N_7233,N_5888,N_5424);
xor U7234 (N_7234,N_5054,N_5234);
xor U7235 (N_7235,N_4348,N_4138);
xor U7236 (N_7236,N_4589,N_4180);
and U7237 (N_7237,N_4752,N_5974);
xnor U7238 (N_7238,N_5801,N_5034);
xnor U7239 (N_7239,N_4504,N_5772);
nand U7240 (N_7240,N_4939,N_5213);
or U7241 (N_7241,N_4367,N_4311);
or U7242 (N_7242,N_4497,N_5778);
and U7243 (N_7243,N_5692,N_5919);
or U7244 (N_7244,N_4540,N_5289);
and U7245 (N_7245,N_5315,N_5570);
and U7246 (N_7246,N_5591,N_5366);
nor U7247 (N_7247,N_4268,N_4560);
nand U7248 (N_7248,N_5031,N_4856);
nor U7249 (N_7249,N_5775,N_4418);
and U7250 (N_7250,N_5568,N_5822);
nand U7251 (N_7251,N_4599,N_5533);
nor U7252 (N_7252,N_4819,N_4532);
or U7253 (N_7253,N_4907,N_4683);
xnor U7254 (N_7254,N_5315,N_4836);
and U7255 (N_7255,N_5645,N_4128);
or U7256 (N_7256,N_5147,N_4720);
xor U7257 (N_7257,N_5696,N_5744);
xnor U7258 (N_7258,N_4764,N_4680);
and U7259 (N_7259,N_4109,N_5221);
nor U7260 (N_7260,N_5829,N_4568);
and U7261 (N_7261,N_4844,N_5433);
nor U7262 (N_7262,N_4492,N_4344);
nand U7263 (N_7263,N_5142,N_5847);
and U7264 (N_7264,N_4569,N_5990);
xnor U7265 (N_7265,N_5041,N_5086);
nand U7266 (N_7266,N_5773,N_5432);
nor U7267 (N_7267,N_4091,N_5784);
and U7268 (N_7268,N_5122,N_4199);
xor U7269 (N_7269,N_5867,N_5242);
or U7270 (N_7270,N_5384,N_4537);
xnor U7271 (N_7271,N_4789,N_5921);
and U7272 (N_7272,N_4685,N_4791);
xnor U7273 (N_7273,N_5788,N_5723);
xnor U7274 (N_7274,N_4765,N_5821);
or U7275 (N_7275,N_5264,N_4140);
or U7276 (N_7276,N_4452,N_5183);
nor U7277 (N_7277,N_4155,N_4658);
and U7278 (N_7278,N_5764,N_4143);
and U7279 (N_7279,N_5836,N_4441);
and U7280 (N_7280,N_4577,N_5276);
nand U7281 (N_7281,N_5123,N_5265);
and U7282 (N_7282,N_4102,N_5032);
or U7283 (N_7283,N_4177,N_5220);
nor U7284 (N_7284,N_4661,N_5429);
and U7285 (N_7285,N_4213,N_5665);
nand U7286 (N_7286,N_5591,N_5889);
and U7287 (N_7287,N_4633,N_4133);
or U7288 (N_7288,N_5361,N_5340);
and U7289 (N_7289,N_5382,N_4624);
nor U7290 (N_7290,N_4464,N_5960);
nand U7291 (N_7291,N_5337,N_5510);
or U7292 (N_7292,N_5695,N_4985);
and U7293 (N_7293,N_4539,N_5003);
nor U7294 (N_7294,N_5797,N_4338);
nand U7295 (N_7295,N_5919,N_4116);
xor U7296 (N_7296,N_4450,N_5183);
nand U7297 (N_7297,N_5914,N_5890);
nor U7298 (N_7298,N_5630,N_5876);
nand U7299 (N_7299,N_5028,N_5399);
and U7300 (N_7300,N_5804,N_5889);
nor U7301 (N_7301,N_5642,N_5438);
nand U7302 (N_7302,N_5910,N_5138);
nor U7303 (N_7303,N_5752,N_5797);
nor U7304 (N_7304,N_4606,N_4184);
or U7305 (N_7305,N_5715,N_4647);
and U7306 (N_7306,N_4716,N_4879);
nand U7307 (N_7307,N_5568,N_5552);
or U7308 (N_7308,N_5700,N_5157);
xnor U7309 (N_7309,N_4708,N_5752);
nand U7310 (N_7310,N_4104,N_5394);
xnor U7311 (N_7311,N_4200,N_4066);
nor U7312 (N_7312,N_5816,N_5487);
nor U7313 (N_7313,N_5066,N_4195);
nor U7314 (N_7314,N_4294,N_4533);
nand U7315 (N_7315,N_5221,N_4330);
and U7316 (N_7316,N_5507,N_4383);
nor U7317 (N_7317,N_5748,N_4001);
or U7318 (N_7318,N_5299,N_4553);
xnor U7319 (N_7319,N_5779,N_4652);
or U7320 (N_7320,N_4678,N_5879);
xor U7321 (N_7321,N_4309,N_4382);
nand U7322 (N_7322,N_5290,N_4710);
and U7323 (N_7323,N_4158,N_5843);
nand U7324 (N_7324,N_5673,N_5399);
nor U7325 (N_7325,N_5161,N_5163);
or U7326 (N_7326,N_5445,N_5775);
xor U7327 (N_7327,N_4613,N_4576);
or U7328 (N_7328,N_4172,N_4446);
nor U7329 (N_7329,N_5630,N_5827);
nand U7330 (N_7330,N_5873,N_5343);
and U7331 (N_7331,N_4964,N_4960);
nand U7332 (N_7332,N_5983,N_4708);
nor U7333 (N_7333,N_4170,N_5490);
nor U7334 (N_7334,N_4886,N_4861);
nand U7335 (N_7335,N_5846,N_4652);
and U7336 (N_7336,N_4707,N_5113);
or U7337 (N_7337,N_5585,N_5045);
nand U7338 (N_7338,N_4460,N_4169);
xnor U7339 (N_7339,N_4858,N_4558);
xnor U7340 (N_7340,N_5607,N_5858);
xor U7341 (N_7341,N_4034,N_4425);
and U7342 (N_7342,N_4875,N_5075);
xnor U7343 (N_7343,N_5214,N_4835);
nand U7344 (N_7344,N_5907,N_4832);
or U7345 (N_7345,N_4845,N_5813);
nor U7346 (N_7346,N_5660,N_5804);
and U7347 (N_7347,N_5064,N_5677);
xor U7348 (N_7348,N_4696,N_5073);
nand U7349 (N_7349,N_5496,N_4424);
nand U7350 (N_7350,N_5024,N_4439);
xor U7351 (N_7351,N_5135,N_5587);
xnor U7352 (N_7352,N_4078,N_5947);
nor U7353 (N_7353,N_4778,N_5798);
nand U7354 (N_7354,N_5242,N_5597);
nor U7355 (N_7355,N_5896,N_4617);
nor U7356 (N_7356,N_5065,N_5559);
or U7357 (N_7357,N_5946,N_5806);
nor U7358 (N_7358,N_5234,N_4312);
nor U7359 (N_7359,N_5543,N_5709);
or U7360 (N_7360,N_4420,N_5014);
and U7361 (N_7361,N_4633,N_4488);
nor U7362 (N_7362,N_4895,N_5339);
xnor U7363 (N_7363,N_4305,N_4247);
and U7364 (N_7364,N_5217,N_5725);
or U7365 (N_7365,N_4524,N_5152);
xor U7366 (N_7366,N_5892,N_5412);
and U7367 (N_7367,N_4769,N_5178);
xnor U7368 (N_7368,N_4996,N_4173);
xnor U7369 (N_7369,N_5331,N_4069);
nand U7370 (N_7370,N_5205,N_4043);
and U7371 (N_7371,N_4573,N_4114);
xor U7372 (N_7372,N_5908,N_4727);
nand U7373 (N_7373,N_5270,N_4128);
nor U7374 (N_7374,N_4187,N_4205);
nand U7375 (N_7375,N_4315,N_5501);
xnor U7376 (N_7376,N_5807,N_4161);
and U7377 (N_7377,N_5134,N_4379);
xnor U7378 (N_7378,N_5303,N_5176);
nand U7379 (N_7379,N_5705,N_5724);
and U7380 (N_7380,N_4044,N_4811);
or U7381 (N_7381,N_4036,N_5278);
xor U7382 (N_7382,N_5738,N_5115);
nor U7383 (N_7383,N_5258,N_5819);
or U7384 (N_7384,N_5737,N_4792);
nor U7385 (N_7385,N_4489,N_5591);
nor U7386 (N_7386,N_5671,N_4512);
xnor U7387 (N_7387,N_5428,N_5377);
or U7388 (N_7388,N_4593,N_4694);
xnor U7389 (N_7389,N_4102,N_4800);
or U7390 (N_7390,N_4959,N_4506);
nor U7391 (N_7391,N_5285,N_4302);
or U7392 (N_7392,N_5444,N_5676);
nor U7393 (N_7393,N_4084,N_4122);
nor U7394 (N_7394,N_4901,N_4933);
nand U7395 (N_7395,N_5498,N_4836);
nand U7396 (N_7396,N_4159,N_5855);
or U7397 (N_7397,N_4227,N_5355);
or U7398 (N_7398,N_5267,N_5618);
or U7399 (N_7399,N_4237,N_4953);
xor U7400 (N_7400,N_4590,N_5915);
xor U7401 (N_7401,N_4061,N_5829);
nor U7402 (N_7402,N_4253,N_4063);
xnor U7403 (N_7403,N_4266,N_4666);
nand U7404 (N_7404,N_4960,N_5314);
nor U7405 (N_7405,N_5460,N_5511);
and U7406 (N_7406,N_5350,N_4957);
xnor U7407 (N_7407,N_5706,N_4065);
nand U7408 (N_7408,N_4208,N_4633);
nand U7409 (N_7409,N_5929,N_4209);
or U7410 (N_7410,N_5340,N_4134);
or U7411 (N_7411,N_5433,N_4923);
or U7412 (N_7412,N_4372,N_5848);
and U7413 (N_7413,N_4228,N_4150);
and U7414 (N_7414,N_5570,N_4482);
xor U7415 (N_7415,N_4760,N_4613);
and U7416 (N_7416,N_5622,N_4024);
and U7417 (N_7417,N_5634,N_5267);
nand U7418 (N_7418,N_5460,N_5499);
xnor U7419 (N_7419,N_4050,N_5092);
and U7420 (N_7420,N_5918,N_4090);
nand U7421 (N_7421,N_4901,N_5834);
and U7422 (N_7422,N_5212,N_4411);
nor U7423 (N_7423,N_4723,N_4379);
and U7424 (N_7424,N_4505,N_5352);
nand U7425 (N_7425,N_4961,N_5864);
and U7426 (N_7426,N_4833,N_5274);
nand U7427 (N_7427,N_5938,N_4754);
nand U7428 (N_7428,N_4491,N_5994);
nor U7429 (N_7429,N_5236,N_4634);
or U7430 (N_7430,N_4903,N_5022);
and U7431 (N_7431,N_5015,N_5208);
nor U7432 (N_7432,N_4496,N_4102);
or U7433 (N_7433,N_5126,N_5399);
or U7434 (N_7434,N_4014,N_5212);
nand U7435 (N_7435,N_4462,N_5237);
nor U7436 (N_7436,N_4939,N_4538);
nand U7437 (N_7437,N_4663,N_5365);
xnor U7438 (N_7438,N_4744,N_5000);
and U7439 (N_7439,N_5839,N_4809);
or U7440 (N_7440,N_5109,N_4368);
xnor U7441 (N_7441,N_4133,N_5556);
and U7442 (N_7442,N_4619,N_5302);
nor U7443 (N_7443,N_5846,N_4461);
or U7444 (N_7444,N_4896,N_5922);
or U7445 (N_7445,N_4578,N_5635);
nor U7446 (N_7446,N_5733,N_5735);
nor U7447 (N_7447,N_4628,N_4228);
xnor U7448 (N_7448,N_5254,N_5583);
xor U7449 (N_7449,N_4715,N_4051);
xor U7450 (N_7450,N_4864,N_4485);
or U7451 (N_7451,N_5157,N_5741);
nor U7452 (N_7452,N_4557,N_4791);
xnor U7453 (N_7453,N_5507,N_5123);
or U7454 (N_7454,N_4122,N_4967);
nor U7455 (N_7455,N_5423,N_5352);
xnor U7456 (N_7456,N_4258,N_4590);
nand U7457 (N_7457,N_4853,N_5604);
xor U7458 (N_7458,N_4274,N_4199);
nor U7459 (N_7459,N_5086,N_4066);
and U7460 (N_7460,N_5734,N_5039);
xor U7461 (N_7461,N_4934,N_5776);
or U7462 (N_7462,N_4742,N_5002);
or U7463 (N_7463,N_5358,N_4425);
xor U7464 (N_7464,N_4856,N_5440);
nand U7465 (N_7465,N_4035,N_5637);
xor U7466 (N_7466,N_5682,N_5207);
or U7467 (N_7467,N_5855,N_5783);
and U7468 (N_7468,N_5882,N_5759);
nor U7469 (N_7469,N_5439,N_5928);
or U7470 (N_7470,N_4547,N_5167);
and U7471 (N_7471,N_5589,N_4164);
xor U7472 (N_7472,N_4473,N_4806);
nor U7473 (N_7473,N_5520,N_4486);
and U7474 (N_7474,N_5632,N_5519);
and U7475 (N_7475,N_5797,N_5678);
and U7476 (N_7476,N_5874,N_4372);
or U7477 (N_7477,N_5110,N_4354);
nand U7478 (N_7478,N_4393,N_4499);
nor U7479 (N_7479,N_4126,N_5325);
nor U7480 (N_7480,N_5024,N_5648);
and U7481 (N_7481,N_5114,N_5866);
nand U7482 (N_7482,N_5860,N_5997);
nand U7483 (N_7483,N_5021,N_5717);
nand U7484 (N_7484,N_5672,N_4682);
or U7485 (N_7485,N_5372,N_5887);
nand U7486 (N_7486,N_4396,N_4124);
and U7487 (N_7487,N_5542,N_5915);
nor U7488 (N_7488,N_5190,N_4787);
xor U7489 (N_7489,N_4084,N_4687);
nor U7490 (N_7490,N_5638,N_5618);
or U7491 (N_7491,N_4155,N_4326);
and U7492 (N_7492,N_4132,N_4446);
nand U7493 (N_7493,N_4716,N_5325);
and U7494 (N_7494,N_4262,N_5635);
nor U7495 (N_7495,N_5204,N_4912);
xnor U7496 (N_7496,N_5912,N_5155);
nand U7497 (N_7497,N_4507,N_4752);
nor U7498 (N_7498,N_4259,N_5567);
or U7499 (N_7499,N_4263,N_5040);
or U7500 (N_7500,N_4891,N_4821);
or U7501 (N_7501,N_4142,N_5677);
or U7502 (N_7502,N_5783,N_4845);
or U7503 (N_7503,N_5270,N_5095);
or U7504 (N_7504,N_4986,N_5432);
nand U7505 (N_7505,N_5841,N_4584);
nand U7506 (N_7506,N_4660,N_5732);
nor U7507 (N_7507,N_5956,N_4343);
xnor U7508 (N_7508,N_4392,N_5532);
xor U7509 (N_7509,N_4637,N_4783);
nor U7510 (N_7510,N_4024,N_4473);
xor U7511 (N_7511,N_5982,N_4409);
nor U7512 (N_7512,N_4583,N_5194);
and U7513 (N_7513,N_5493,N_4156);
or U7514 (N_7514,N_5941,N_4006);
or U7515 (N_7515,N_5455,N_5298);
nor U7516 (N_7516,N_5021,N_4301);
nor U7517 (N_7517,N_5604,N_4435);
nor U7518 (N_7518,N_5944,N_5419);
xnor U7519 (N_7519,N_5843,N_4313);
nand U7520 (N_7520,N_4942,N_4908);
nor U7521 (N_7521,N_4667,N_5719);
nand U7522 (N_7522,N_4400,N_5959);
xor U7523 (N_7523,N_4627,N_5449);
and U7524 (N_7524,N_5796,N_5340);
xnor U7525 (N_7525,N_5058,N_5438);
and U7526 (N_7526,N_4558,N_5366);
and U7527 (N_7527,N_5889,N_5405);
nand U7528 (N_7528,N_4420,N_4761);
or U7529 (N_7529,N_4787,N_5046);
and U7530 (N_7530,N_5492,N_4852);
nor U7531 (N_7531,N_4730,N_4301);
or U7532 (N_7532,N_5524,N_5089);
and U7533 (N_7533,N_4278,N_5076);
or U7534 (N_7534,N_4936,N_4364);
xnor U7535 (N_7535,N_4359,N_5482);
nor U7536 (N_7536,N_4399,N_4167);
or U7537 (N_7537,N_4342,N_4249);
nand U7538 (N_7538,N_5270,N_4432);
nand U7539 (N_7539,N_5696,N_4360);
or U7540 (N_7540,N_4553,N_5950);
xor U7541 (N_7541,N_4749,N_4814);
xnor U7542 (N_7542,N_5042,N_5230);
xnor U7543 (N_7543,N_4232,N_4632);
xnor U7544 (N_7544,N_5590,N_4128);
nand U7545 (N_7545,N_4295,N_4774);
nor U7546 (N_7546,N_5024,N_4563);
nand U7547 (N_7547,N_4879,N_5975);
and U7548 (N_7548,N_5747,N_4019);
and U7549 (N_7549,N_4489,N_5255);
nand U7550 (N_7550,N_4343,N_4574);
nand U7551 (N_7551,N_4387,N_4893);
and U7552 (N_7552,N_5045,N_4203);
and U7553 (N_7553,N_5749,N_5195);
nor U7554 (N_7554,N_4369,N_5115);
nand U7555 (N_7555,N_4187,N_4175);
nand U7556 (N_7556,N_5242,N_4215);
and U7557 (N_7557,N_4939,N_4607);
and U7558 (N_7558,N_5846,N_5003);
nand U7559 (N_7559,N_4756,N_4516);
nor U7560 (N_7560,N_4488,N_5038);
or U7561 (N_7561,N_5037,N_4449);
nand U7562 (N_7562,N_5586,N_4961);
nand U7563 (N_7563,N_4626,N_5461);
xor U7564 (N_7564,N_5297,N_4072);
and U7565 (N_7565,N_5163,N_5495);
or U7566 (N_7566,N_5948,N_5514);
xor U7567 (N_7567,N_4232,N_4040);
xor U7568 (N_7568,N_5096,N_4463);
and U7569 (N_7569,N_5815,N_5626);
and U7570 (N_7570,N_5574,N_5493);
nor U7571 (N_7571,N_4328,N_5109);
xnor U7572 (N_7572,N_4624,N_5001);
nor U7573 (N_7573,N_5681,N_5953);
nand U7574 (N_7574,N_5841,N_4637);
nor U7575 (N_7575,N_5295,N_4437);
or U7576 (N_7576,N_4688,N_4528);
nand U7577 (N_7577,N_4877,N_5900);
xnor U7578 (N_7578,N_4551,N_5423);
nor U7579 (N_7579,N_5786,N_4862);
nand U7580 (N_7580,N_4906,N_5367);
xor U7581 (N_7581,N_4526,N_4006);
nand U7582 (N_7582,N_5977,N_4908);
nand U7583 (N_7583,N_5977,N_5714);
and U7584 (N_7584,N_5310,N_4678);
nor U7585 (N_7585,N_4582,N_4547);
nor U7586 (N_7586,N_5836,N_5647);
nand U7587 (N_7587,N_4354,N_5211);
xnor U7588 (N_7588,N_5812,N_4799);
xnor U7589 (N_7589,N_4274,N_5856);
xnor U7590 (N_7590,N_5411,N_4586);
xnor U7591 (N_7591,N_4879,N_4753);
nor U7592 (N_7592,N_5434,N_4840);
nand U7593 (N_7593,N_5186,N_5386);
nand U7594 (N_7594,N_4443,N_5069);
and U7595 (N_7595,N_4477,N_5230);
and U7596 (N_7596,N_4052,N_4139);
or U7597 (N_7597,N_5507,N_4304);
and U7598 (N_7598,N_5260,N_4021);
nor U7599 (N_7599,N_4472,N_5749);
and U7600 (N_7600,N_4090,N_5446);
or U7601 (N_7601,N_5348,N_5926);
xor U7602 (N_7602,N_5996,N_4403);
xor U7603 (N_7603,N_5875,N_5397);
or U7604 (N_7604,N_4767,N_5124);
nor U7605 (N_7605,N_4434,N_5838);
or U7606 (N_7606,N_4458,N_5766);
or U7607 (N_7607,N_4819,N_4296);
xor U7608 (N_7608,N_4089,N_5015);
or U7609 (N_7609,N_4944,N_5092);
xnor U7610 (N_7610,N_5018,N_4848);
xor U7611 (N_7611,N_5624,N_4124);
xnor U7612 (N_7612,N_4953,N_4123);
xor U7613 (N_7613,N_5925,N_5006);
nand U7614 (N_7614,N_4299,N_5631);
and U7615 (N_7615,N_4533,N_4519);
xnor U7616 (N_7616,N_4101,N_4047);
or U7617 (N_7617,N_5089,N_5752);
nor U7618 (N_7618,N_5796,N_4124);
nand U7619 (N_7619,N_4023,N_4922);
or U7620 (N_7620,N_5654,N_4263);
or U7621 (N_7621,N_4572,N_5529);
nand U7622 (N_7622,N_5160,N_5321);
nand U7623 (N_7623,N_4389,N_4221);
nand U7624 (N_7624,N_5234,N_5302);
nor U7625 (N_7625,N_5535,N_5243);
nand U7626 (N_7626,N_4210,N_5520);
or U7627 (N_7627,N_4420,N_5905);
nand U7628 (N_7628,N_4342,N_4040);
nor U7629 (N_7629,N_5257,N_4004);
and U7630 (N_7630,N_4699,N_5222);
nor U7631 (N_7631,N_4812,N_4231);
xnor U7632 (N_7632,N_5739,N_5395);
xnor U7633 (N_7633,N_5391,N_4434);
or U7634 (N_7634,N_5971,N_4254);
nand U7635 (N_7635,N_5212,N_4560);
or U7636 (N_7636,N_5144,N_5092);
nor U7637 (N_7637,N_4247,N_5139);
and U7638 (N_7638,N_5708,N_4877);
or U7639 (N_7639,N_5598,N_4563);
xor U7640 (N_7640,N_4275,N_4981);
nand U7641 (N_7641,N_4831,N_5518);
nand U7642 (N_7642,N_4822,N_5882);
or U7643 (N_7643,N_5407,N_4523);
nand U7644 (N_7644,N_5273,N_5956);
and U7645 (N_7645,N_4700,N_5428);
nand U7646 (N_7646,N_5762,N_4083);
and U7647 (N_7647,N_5181,N_5000);
or U7648 (N_7648,N_5575,N_5116);
nand U7649 (N_7649,N_5869,N_4635);
xor U7650 (N_7650,N_4401,N_5400);
or U7651 (N_7651,N_5084,N_5731);
and U7652 (N_7652,N_5825,N_4161);
and U7653 (N_7653,N_5964,N_4773);
xor U7654 (N_7654,N_4630,N_4074);
nor U7655 (N_7655,N_5573,N_5010);
or U7656 (N_7656,N_4791,N_4088);
or U7657 (N_7657,N_5692,N_5606);
nand U7658 (N_7658,N_4049,N_4107);
nand U7659 (N_7659,N_4304,N_5241);
or U7660 (N_7660,N_4091,N_5149);
nor U7661 (N_7661,N_4664,N_5157);
xnor U7662 (N_7662,N_5100,N_4189);
nor U7663 (N_7663,N_4264,N_5431);
or U7664 (N_7664,N_4485,N_5453);
or U7665 (N_7665,N_4460,N_4240);
nor U7666 (N_7666,N_5102,N_5514);
nor U7667 (N_7667,N_4677,N_4918);
or U7668 (N_7668,N_4429,N_4271);
xnor U7669 (N_7669,N_5160,N_4115);
or U7670 (N_7670,N_4827,N_5110);
nor U7671 (N_7671,N_5578,N_4208);
xor U7672 (N_7672,N_5396,N_5269);
nand U7673 (N_7673,N_5030,N_4013);
xor U7674 (N_7674,N_4368,N_4308);
nand U7675 (N_7675,N_5715,N_5740);
and U7676 (N_7676,N_5902,N_4949);
or U7677 (N_7677,N_4254,N_5627);
and U7678 (N_7678,N_4540,N_4674);
nand U7679 (N_7679,N_5404,N_4157);
nand U7680 (N_7680,N_4845,N_4522);
xnor U7681 (N_7681,N_4857,N_4567);
and U7682 (N_7682,N_4457,N_4824);
and U7683 (N_7683,N_5500,N_4530);
nand U7684 (N_7684,N_4103,N_5977);
or U7685 (N_7685,N_4543,N_4411);
nor U7686 (N_7686,N_4567,N_5975);
and U7687 (N_7687,N_5641,N_4113);
nor U7688 (N_7688,N_4898,N_5974);
xnor U7689 (N_7689,N_5906,N_5004);
xor U7690 (N_7690,N_4651,N_4671);
nand U7691 (N_7691,N_5019,N_4436);
xor U7692 (N_7692,N_5152,N_4130);
or U7693 (N_7693,N_5362,N_5518);
and U7694 (N_7694,N_5907,N_5335);
xnor U7695 (N_7695,N_5426,N_4727);
nand U7696 (N_7696,N_5463,N_4330);
nor U7697 (N_7697,N_4291,N_5640);
nand U7698 (N_7698,N_5817,N_5457);
nor U7699 (N_7699,N_4336,N_4075);
or U7700 (N_7700,N_4206,N_4643);
nand U7701 (N_7701,N_4217,N_4168);
nor U7702 (N_7702,N_5340,N_4895);
xnor U7703 (N_7703,N_5001,N_5618);
xor U7704 (N_7704,N_4783,N_5849);
or U7705 (N_7705,N_4499,N_4017);
and U7706 (N_7706,N_4002,N_4735);
nor U7707 (N_7707,N_5607,N_4383);
nand U7708 (N_7708,N_5256,N_5963);
xnor U7709 (N_7709,N_4376,N_5969);
nand U7710 (N_7710,N_5509,N_5817);
or U7711 (N_7711,N_5611,N_5121);
nand U7712 (N_7712,N_5246,N_4750);
nor U7713 (N_7713,N_4702,N_5701);
and U7714 (N_7714,N_4522,N_5704);
and U7715 (N_7715,N_5409,N_5877);
and U7716 (N_7716,N_4621,N_5617);
nor U7717 (N_7717,N_4183,N_4629);
and U7718 (N_7718,N_4344,N_4276);
or U7719 (N_7719,N_4496,N_4420);
nand U7720 (N_7720,N_5218,N_5623);
xor U7721 (N_7721,N_5938,N_4638);
and U7722 (N_7722,N_4415,N_4760);
and U7723 (N_7723,N_4806,N_4454);
and U7724 (N_7724,N_4878,N_5840);
and U7725 (N_7725,N_5207,N_5420);
xnor U7726 (N_7726,N_5631,N_4790);
and U7727 (N_7727,N_5445,N_5813);
or U7728 (N_7728,N_5373,N_4587);
xnor U7729 (N_7729,N_4771,N_4473);
nor U7730 (N_7730,N_5705,N_5092);
nor U7731 (N_7731,N_4037,N_4511);
and U7732 (N_7732,N_5744,N_5142);
nand U7733 (N_7733,N_4881,N_4590);
or U7734 (N_7734,N_5654,N_5475);
or U7735 (N_7735,N_4848,N_5281);
or U7736 (N_7736,N_5105,N_5115);
nand U7737 (N_7737,N_4742,N_4068);
and U7738 (N_7738,N_4130,N_5725);
nand U7739 (N_7739,N_4665,N_5103);
xor U7740 (N_7740,N_4579,N_5561);
nand U7741 (N_7741,N_4121,N_4030);
or U7742 (N_7742,N_5940,N_5993);
or U7743 (N_7743,N_4701,N_5211);
nor U7744 (N_7744,N_5775,N_5572);
or U7745 (N_7745,N_5297,N_4996);
or U7746 (N_7746,N_5467,N_4680);
xnor U7747 (N_7747,N_4266,N_4920);
nor U7748 (N_7748,N_4607,N_5314);
or U7749 (N_7749,N_4522,N_5767);
nand U7750 (N_7750,N_4515,N_5217);
and U7751 (N_7751,N_4179,N_5185);
nor U7752 (N_7752,N_4948,N_5430);
and U7753 (N_7753,N_5596,N_4067);
or U7754 (N_7754,N_5149,N_5492);
nor U7755 (N_7755,N_4897,N_5914);
or U7756 (N_7756,N_5296,N_5242);
nor U7757 (N_7757,N_4187,N_4888);
nor U7758 (N_7758,N_5042,N_5923);
or U7759 (N_7759,N_5504,N_4739);
xnor U7760 (N_7760,N_5861,N_5917);
or U7761 (N_7761,N_5114,N_4524);
and U7762 (N_7762,N_5393,N_4762);
xnor U7763 (N_7763,N_5040,N_5858);
and U7764 (N_7764,N_5027,N_4200);
or U7765 (N_7765,N_5456,N_4583);
nor U7766 (N_7766,N_5222,N_5655);
nor U7767 (N_7767,N_5044,N_5701);
xor U7768 (N_7768,N_4632,N_4445);
nor U7769 (N_7769,N_4039,N_5864);
nor U7770 (N_7770,N_4074,N_4411);
xnor U7771 (N_7771,N_5171,N_4255);
or U7772 (N_7772,N_5530,N_5615);
nor U7773 (N_7773,N_5477,N_4455);
xor U7774 (N_7774,N_5908,N_4871);
nand U7775 (N_7775,N_4053,N_5221);
nand U7776 (N_7776,N_5717,N_5800);
and U7777 (N_7777,N_5053,N_4636);
or U7778 (N_7778,N_4921,N_5451);
xor U7779 (N_7779,N_5379,N_4181);
and U7780 (N_7780,N_4487,N_4285);
and U7781 (N_7781,N_4327,N_5459);
xor U7782 (N_7782,N_5886,N_5275);
nor U7783 (N_7783,N_4997,N_5356);
or U7784 (N_7784,N_5205,N_4728);
nand U7785 (N_7785,N_5399,N_5994);
and U7786 (N_7786,N_5173,N_4125);
or U7787 (N_7787,N_4880,N_4553);
and U7788 (N_7788,N_4673,N_4245);
and U7789 (N_7789,N_4938,N_4221);
or U7790 (N_7790,N_4517,N_5402);
or U7791 (N_7791,N_5989,N_5835);
nor U7792 (N_7792,N_4551,N_4747);
and U7793 (N_7793,N_4165,N_5696);
xnor U7794 (N_7794,N_4975,N_4932);
and U7795 (N_7795,N_5043,N_5690);
or U7796 (N_7796,N_4559,N_5948);
xor U7797 (N_7797,N_4929,N_4804);
nor U7798 (N_7798,N_5008,N_4076);
nand U7799 (N_7799,N_5935,N_4903);
nor U7800 (N_7800,N_4851,N_4062);
or U7801 (N_7801,N_4496,N_4401);
or U7802 (N_7802,N_4929,N_4547);
nand U7803 (N_7803,N_5067,N_5003);
nand U7804 (N_7804,N_5362,N_4329);
xnor U7805 (N_7805,N_5440,N_4076);
xor U7806 (N_7806,N_4963,N_5566);
or U7807 (N_7807,N_5456,N_4837);
or U7808 (N_7808,N_4294,N_5556);
and U7809 (N_7809,N_4723,N_4134);
and U7810 (N_7810,N_5541,N_5533);
or U7811 (N_7811,N_4620,N_5656);
xnor U7812 (N_7812,N_5561,N_4661);
or U7813 (N_7813,N_4719,N_5229);
nand U7814 (N_7814,N_5212,N_5026);
and U7815 (N_7815,N_4971,N_4055);
nor U7816 (N_7816,N_5762,N_4739);
xor U7817 (N_7817,N_4050,N_4284);
nor U7818 (N_7818,N_4471,N_5984);
xor U7819 (N_7819,N_4713,N_5363);
xor U7820 (N_7820,N_4721,N_4093);
and U7821 (N_7821,N_5056,N_5748);
or U7822 (N_7822,N_4299,N_4346);
nand U7823 (N_7823,N_4394,N_5289);
and U7824 (N_7824,N_4634,N_5106);
or U7825 (N_7825,N_4715,N_4351);
nor U7826 (N_7826,N_4422,N_5703);
xnor U7827 (N_7827,N_4995,N_4449);
and U7828 (N_7828,N_5514,N_4155);
nand U7829 (N_7829,N_5233,N_5534);
or U7830 (N_7830,N_4568,N_4075);
nor U7831 (N_7831,N_4683,N_5490);
and U7832 (N_7832,N_4071,N_5148);
and U7833 (N_7833,N_5460,N_5899);
or U7834 (N_7834,N_5741,N_4384);
nand U7835 (N_7835,N_5136,N_4785);
nor U7836 (N_7836,N_5652,N_5869);
xnor U7837 (N_7837,N_5446,N_4221);
or U7838 (N_7838,N_4986,N_5618);
xnor U7839 (N_7839,N_5475,N_4873);
or U7840 (N_7840,N_5063,N_4250);
and U7841 (N_7841,N_5250,N_4356);
nor U7842 (N_7842,N_4997,N_5941);
xnor U7843 (N_7843,N_5360,N_5187);
nor U7844 (N_7844,N_5184,N_4880);
and U7845 (N_7845,N_4902,N_4349);
or U7846 (N_7846,N_5098,N_5914);
nor U7847 (N_7847,N_4269,N_4429);
and U7848 (N_7848,N_5735,N_4471);
nand U7849 (N_7849,N_4767,N_4643);
or U7850 (N_7850,N_4750,N_5391);
xor U7851 (N_7851,N_5264,N_4418);
xor U7852 (N_7852,N_4046,N_4831);
and U7853 (N_7853,N_4519,N_4574);
xor U7854 (N_7854,N_5691,N_5417);
and U7855 (N_7855,N_5924,N_4258);
nand U7856 (N_7856,N_5001,N_5333);
xnor U7857 (N_7857,N_5141,N_5683);
xor U7858 (N_7858,N_4588,N_4838);
nand U7859 (N_7859,N_5811,N_4660);
nand U7860 (N_7860,N_5608,N_5941);
nand U7861 (N_7861,N_4853,N_5085);
nor U7862 (N_7862,N_5481,N_4280);
nand U7863 (N_7863,N_5904,N_5791);
nand U7864 (N_7864,N_4068,N_4440);
and U7865 (N_7865,N_4693,N_5067);
and U7866 (N_7866,N_5981,N_4744);
nand U7867 (N_7867,N_5496,N_4862);
xor U7868 (N_7868,N_5929,N_5780);
xnor U7869 (N_7869,N_4102,N_5570);
xnor U7870 (N_7870,N_4403,N_4573);
nor U7871 (N_7871,N_5627,N_4052);
and U7872 (N_7872,N_4117,N_5163);
nand U7873 (N_7873,N_5419,N_4195);
or U7874 (N_7874,N_4361,N_4816);
nand U7875 (N_7875,N_4972,N_4776);
nand U7876 (N_7876,N_4255,N_5023);
and U7877 (N_7877,N_4637,N_5106);
xor U7878 (N_7878,N_5759,N_4826);
nor U7879 (N_7879,N_5158,N_4827);
nor U7880 (N_7880,N_4923,N_4126);
or U7881 (N_7881,N_5607,N_5766);
or U7882 (N_7882,N_4167,N_5875);
and U7883 (N_7883,N_4181,N_4964);
and U7884 (N_7884,N_4061,N_5393);
nor U7885 (N_7885,N_4281,N_4844);
xor U7886 (N_7886,N_4998,N_4466);
and U7887 (N_7887,N_5960,N_4689);
or U7888 (N_7888,N_5541,N_5198);
nand U7889 (N_7889,N_5458,N_5878);
nand U7890 (N_7890,N_5479,N_5446);
xor U7891 (N_7891,N_5513,N_4424);
xor U7892 (N_7892,N_5035,N_4095);
or U7893 (N_7893,N_4695,N_5975);
and U7894 (N_7894,N_4622,N_4813);
nor U7895 (N_7895,N_5796,N_5003);
or U7896 (N_7896,N_5622,N_4193);
nand U7897 (N_7897,N_5898,N_4209);
nor U7898 (N_7898,N_4703,N_4793);
and U7899 (N_7899,N_5190,N_4953);
and U7900 (N_7900,N_4436,N_4379);
nand U7901 (N_7901,N_5609,N_4110);
nor U7902 (N_7902,N_4525,N_5349);
or U7903 (N_7903,N_4510,N_4480);
or U7904 (N_7904,N_4043,N_5396);
and U7905 (N_7905,N_4793,N_5480);
and U7906 (N_7906,N_5451,N_5704);
nand U7907 (N_7907,N_4647,N_5488);
nand U7908 (N_7908,N_5211,N_5288);
or U7909 (N_7909,N_4801,N_5128);
and U7910 (N_7910,N_5391,N_4223);
nor U7911 (N_7911,N_5540,N_4587);
and U7912 (N_7912,N_5282,N_4391);
and U7913 (N_7913,N_4304,N_4431);
xor U7914 (N_7914,N_5758,N_5433);
xor U7915 (N_7915,N_4986,N_5724);
nor U7916 (N_7916,N_4507,N_5039);
nor U7917 (N_7917,N_4425,N_5823);
xnor U7918 (N_7918,N_5469,N_4749);
xor U7919 (N_7919,N_5375,N_5609);
or U7920 (N_7920,N_4211,N_5608);
nand U7921 (N_7921,N_5714,N_5217);
and U7922 (N_7922,N_4060,N_4652);
or U7923 (N_7923,N_4712,N_4001);
nand U7924 (N_7924,N_4507,N_4923);
nand U7925 (N_7925,N_4579,N_5165);
and U7926 (N_7926,N_4409,N_4618);
xnor U7927 (N_7927,N_4050,N_4224);
nor U7928 (N_7928,N_4283,N_4295);
xor U7929 (N_7929,N_4035,N_4100);
or U7930 (N_7930,N_5652,N_5246);
nand U7931 (N_7931,N_5192,N_4407);
xor U7932 (N_7932,N_5920,N_5906);
xor U7933 (N_7933,N_5529,N_5456);
or U7934 (N_7934,N_5147,N_4216);
nor U7935 (N_7935,N_4113,N_4993);
nand U7936 (N_7936,N_4752,N_5188);
nand U7937 (N_7937,N_4065,N_4070);
and U7938 (N_7938,N_4518,N_5311);
or U7939 (N_7939,N_5999,N_4310);
and U7940 (N_7940,N_4714,N_4281);
xnor U7941 (N_7941,N_5536,N_5333);
xnor U7942 (N_7942,N_4136,N_5494);
xor U7943 (N_7943,N_5582,N_4198);
nand U7944 (N_7944,N_5115,N_5266);
xnor U7945 (N_7945,N_5783,N_5475);
xor U7946 (N_7946,N_5725,N_4307);
nand U7947 (N_7947,N_5329,N_4224);
nor U7948 (N_7948,N_5924,N_5592);
nand U7949 (N_7949,N_4451,N_4431);
xor U7950 (N_7950,N_5077,N_4530);
or U7951 (N_7951,N_5051,N_5318);
nand U7952 (N_7952,N_5824,N_5140);
xor U7953 (N_7953,N_5312,N_5727);
nand U7954 (N_7954,N_4074,N_5443);
or U7955 (N_7955,N_4578,N_5675);
xor U7956 (N_7956,N_4286,N_5771);
and U7957 (N_7957,N_4116,N_4545);
nor U7958 (N_7958,N_5311,N_4339);
or U7959 (N_7959,N_5852,N_4437);
nand U7960 (N_7960,N_4943,N_4142);
nand U7961 (N_7961,N_4886,N_4245);
and U7962 (N_7962,N_4177,N_4704);
nor U7963 (N_7963,N_5393,N_5580);
or U7964 (N_7964,N_4343,N_5846);
nor U7965 (N_7965,N_5835,N_5817);
and U7966 (N_7966,N_4259,N_4142);
xor U7967 (N_7967,N_5237,N_4593);
or U7968 (N_7968,N_5274,N_5767);
nand U7969 (N_7969,N_4279,N_5955);
and U7970 (N_7970,N_5368,N_4671);
nand U7971 (N_7971,N_4703,N_4140);
or U7972 (N_7972,N_4138,N_4629);
and U7973 (N_7973,N_4050,N_4009);
nand U7974 (N_7974,N_5353,N_5231);
or U7975 (N_7975,N_4558,N_5835);
nand U7976 (N_7976,N_5450,N_4929);
nor U7977 (N_7977,N_4632,N_5478);
nor U7978 (N_7978,N_5870,N_4921);
and U7979 (N_7979,N_4737,N_4954);
nand U7980 (N_7980,N_5432,N_5279);
and U7981 (N_7981,N_4325,N_4701);
nor U7982 (N_7982,N_4423,N_4267);
and U7983 (N_7983,N_4257,N_4395);
nand U7984 (N_7984,N_5339,N_4681);
nand U7985 (N_7985,N_4558,N_5238);
xor U7986 (N_7986,N_4360,N_5533);
or U7987 (N_7987,N_5206,N_5881);
nor U7988 (N_7988,N_4634,N_4135);
and U7989 (N_7989,N_4989,N_4547);
nor U7990 (N_7990,N_5810,N_5652);
and U7991 (N_7991,N_4101,N_5636);
and U7992 (N_7992,N_5925,N_5935);
or U7993 (N_7993,N_4977,N_4690);
nand U7994 (N_7994,N_4609,N_5745);
xnor U7995 (N_7995,N_4325,N_5298);
nand U7996 (N_7996,N_5633,N_4860);
or U7997 (N_7997,N_5001,N_4495);
nor U7998 (N_7998,N_4571,N_4676);
xnor U7999 (N_7999,N_4031,N_4050);
nand U8000 (N_8000,N_7318,N_7915);
nand U8001 (N_8001,N_7303,N_7940);
and U8002 (N_8002,N_7863,N_6961);
or U8003 (N_8003,N_7828,N_7161);
nand U8004 (N_8004,N_6241,N_7596);
nor U8005 (N_8005,N_6713,N_7108);
xnor U8006 (N_8006,N_7075,N_7930);
or U8007 (N_8007,N_6670,N_7539);
nand U8008 (N_8008,N_6821,N_6279);
and U8009 (N_8009,N_7740,N_6493);
xnor U8010 (N_8010,N_6283,N_6980);
nor U8011 (N_8011,N_7272,N_6846);
xor U8012 (N_8012,N_7483,N_6917);
and U8013 (N_8013,N_6574,N_6571);
nor U8014 (N_8014,N_6415,N_7455);
and U8015 (N_8015,N_6428,N_7273);
nand U8016 (N_8016,N_6792,N_7908);
or U8017 (N_8017,N_7301,N_6944);
nand U8018 (N_8018,N_6263,N_7632);
and U8019 (N_8019,N_7566,N_6752);
nand U8020 (N_8020,N_7046,N_6437);
and U8021 (N_8021,N_7495,N_7124);
or U8022 (N_8022,N_6839,N_6921);
nand U8023 (N_8023,N_6854,N_7487);
nor U8024 (N_8024,N_7992,N_6856);
nand U8025 (N_8025,N_7575,N_7742);
nand U8026 (N_8026,N_7793,N_7997);
and U8027 (N_8027,N_7942,N_7041);
and U8028 (N_8028,N_7984,N_7486);
or U8029 (N_8029,N_7673,N_6001);
and U8030 (N_8030,N_7594,N_7088);
or U8031 (N_8031,N_6138,N_6629);
nor U8032 (N_8032,N_6442,N_7344);
nand U8033 (N_8033,N_6047,N_6294);
or U8034 (N_8034,N_6297,N_7474);
nor U8035 (N_8035,N_6551,N_7284);
nand U8036 (N_8036,N_6278,N_6050);
nor U8037 (N_8037,N_7432,N_6897);
or U8038 (N_8038,N_6410,N_6749);
nand U8039 (N_8039,N_7751,N_6417);
and U8040 (N_8040,N_6421,N_6561);
and U8041 (N_8041,N_6740,N_7674);
nand U8042 (N_8042,N_7343,N_6105);
and U8043 (N_8043,N_6676,N_7228);
nand U8044 (N_8044,N_6034,N_7456);
or U8045 (N_8045,N_6125,N_7978);
or U8046 (N_8046,N_7694,N_7248);
or U8047 (N_8047,N_6120,N_6024);
nand U8048 (N_8048,N_7559,N_7346);
nand U8049 (N_8049,N_7219,N_6965);
nor U8050 (N_8050,N_7961,N_7900);
or U8051 (N_8051,N_6890,N_7720);
and U8052 (N_8052,N_7563,N_6804);
or U8053 (N_8053,N_6218,N_6943);
xnor U8054 (N_8054,N_6336,N_7047);
and U8055 (N_8055,N_6150,N_6128);
nand U8056 (N_8056,N_7147,N_7542);
xor U8057 (N_8057,N_6175,N_7711);
nor U8058 (N_8058,N_7240,N_7198);
nor U8059 (N_8059,N_7689,N_7618);
nor U8060 (N_8060,N_6626,N_7239);
and U8061 (N_8061,N_7823,N_7431);
and U8062 (N_8062,N_7347,N_6790);
nor U8063 (N_8063,N_6778,N_6510);
and U8064 (N_8064,N_6580,N_7119);
or U8065 (N_8065,N_7599,N_7924);
nor U8066 (N_8066,N_7561,N_7913);
or U8067 (N_8067,N_7579,N_7173);
or U8068 (N_8068,N_6553,N_6027);
or U8069 (N_8069,N_6562,N_7317);
or U8070 (N_8070,N_7496,N_6738);
nor U8071 (N_8071,N_7033,N_7274);
nand U8072 (N_8072,N_7769,N_7645);
or U8073 (N_8073,N_7378,N_7236);
or U8074 (N_8074,N_6525,N_6793);
or U8075 (N_8075,N_7926,N_6158);
nand U8076 (N_8076,N_7578,N_7507);
xnor U8077 (N_8077,N_7049,N_7857);
xnor U8078 (N_8078,N_6775,N_7960);
nand U8079 (N_8079,N_6457,N_7146);
or U8080 (N_8080,N_7759,N_6837);
or U8081 (N_8081,N_6518,N_6806);
or U8082 (N_8082,N_6545,N_7730);
xnor U8083 (N_8083,N_7061,N_6686);
xor U8084 (N_8084,N_7326,N_7194);
nand U8085 (N_8085,N_6989,N_6824);
nor U8086 (N_8086,N_7149,N_7439);
and U8087 (N_8087,N_7941,N_6005);
or U8088 (N_8088,N_6329,N_7741);
nor U8089 (N_8089,N_7083,N_6311);
nand U8090 (N_8090,N_6645,N_6883);
nand U8091 (N_8091,N_6986,N_6231);
nand U8092 (N_8092,N_6134,N_7567);
or U8093 (N_8093,N_6119,N_7520);
and U8094 (N_8094,N_7830,N_7148);
xor U8095 (N_8095,N_7949,N_7081);
or U8096 (N_8096,N_7381,N_6305);
nor U8097 (N_8097,N_6282,N_7154);
or U8098 (N_8098,N_6472,N_7766);
nor U8099 (N_8099,N_6333,N_6742);
nand U8100 (N_8100,N_6028,N_6527);
nor U8101 (N_8101,N_6835,N_7386);
nand U8102 (N_8102,N_7158,N_6404);
xnor U8103 (N_8103,N_7145,N_7609);
nor U8104 (N_8104,N_7979,N_7846);
nand U8105 (N_8105,N_7505,N_6974);
and U8106 (N_8106,N_7899,N_6253);
nor U8107 (N_8107,N_6289,N_7062);
nand U8108 (N_8108,N_6164,N_6530);
nor U8109 (N_8109,N_6478,N_6464);
and U8110 (N_8110,N_7509,N_7195);
xnor U8111 (N_8111,N_7706,N_6217);
nand U8112 (N_8112,N_6092,N_6782);
or U8113 (N_8113,N_7529,N_7393);
nand U8114 (N_8114,N_6032,N_7245);
nand U8115 (N_8115,N_6157,N_7137);
or U8116 (N_8116,N_6358,N_6007);
and U8117 (N_8117,N_6176,N_7739);
or U8118 (N_8118,N_7349,N_7351);
and U8119 (N_8119,N_7664,N_6045);
nand U8120 (N_8120,N_6697,N_6950);
and U8121 (N_8121,N_6129,N_6747);
or U8122 (N_8122,N_7150,N_7933);
nand U8123 (N_8123,N_6744,N_7438);
and U8124 (N_8124,N_7196,N_6998);
and U8125 (N_8125,N_6221,N_6165);
nand U8126 (N_8126,N_7805,N_7078);
nor U8127 (N_8127,N_7867,N_7768);
nor U8128 (N_8128,N_6549,N_6113);
nand U8129 (N_8129,N_6768,N_6363);
or U8130 (N_8130,N_7527,N_7192);
xor U8131 (N_8131,N_6242,N_6148);
nor U8132 (N_8132,N_6145,N_6287);
or U8133 (N_8133,N_7868,N_6108);
xnor U8134 (N_8134,N_7528,N_7855);
or U8135 (N_8135,N_7259,N_6813);
or U8136 (N_8136,N_7564,N_6817);
or U8137 (N_8137,N_6632,N_6750);
nor U8138 (N_8138,N_6262,N_6056);
and U8139 (N_8139,N_7110,N_6465);
or U8140 (N_8140,N_7523,N_7948);
and U8141 (N_8141,N_6834,N_6444);
nand U8142 (N_8142,N_7494,N_7947);
nor U8143 (N_8143,N_7329,N_7657);
and U8144 (N_8144,N_6992,N_6192);
xnor U8145 (N_8145,N_6570,N_6754);
xnor U8146 (N_8146,N_6907,N_6521);
xnor U8147 (N_8147,N_7889,N_6402);
and U8148 (N_8148,N_6416,N_7633);
nor U8149 (N_8149,N_6062,N_7059);
or U8150 (N_8150,N_6162,N_6963);
nand U8151 (N_8151,N_6709,N_7186);
or U8152 (N_8152,N_6631,N_7652);
nor U8153 (N_8153,N_7371,N_7927);
or U8154 (N_8154,N_7953,N_6433);
and U8155 (N_8155,N_6331,N_6181);
or U8156 (N_8156,N_6894,N_6985);
and U8157 (N_8157,N_6436,N_7576);
and U8158 (N_8158,N_7157,N_7403);
and U8159 (N_8159,N_7525,N_6653);
or U8160 (N_8160,N_6213,N_7521);
xnor U8161 (N_8161,N_7121,N_6296);
and U8162 (N_8162,N_6703,N_6334);
and U8163 (N_8163,N_6797,N_6885);
xor U8164 (N_8164,N_6006,N_7190);
nor U8165 (N_8165,N_6597,N_7454);
or U8166 (N_8166,N_7399,N_7018);
xnor U8167 (N_8167,N_7373,N_6042);
nand U8168 (N_8168,N_7015,N_6630);
and U8169 (N_8169,N_6168,N_7697);
nand U8170 (N_8170,N_7723,N_6224);
and U8171 (N_8171,N_6893,N_6348);
and U8172 (N_8172,N_6452,N_6802);
or U8173 (N_8173,N_6903,N_6516);
and U8174 (N_8174,N_6277,N_7458);
nand U8175 (N_8175,N_7925,N_6724);
or U8176 (N_8176,N_6850,N_7315);
xnor U8177 (N_8177,N_6151,N_6678);
xnor U8178 (N_8178,N_7334,N_7208);
or U8179 (N_8179,N_6316,N_7125);
and U8180 (N_8180,N_6867,N_6648);
and U8181 (N_8181,N_6857,N_6957);
xor U8182 (N_8182,N_6714,N_6236);
or U8183 (N_8183,N_7874,N_6968);
nand U8184 (N_8184,N_6863,N_6689);
nand U8185 (N_8185,N_6400,N_7389);
nor U8186 (N_8186,N_7881,N_7612);
xnor U8187 (N_8187,N_6187,N_7355);
and U8188 (N_8188,N_6508,N_6734);
nand U8189 (N_8189,N_7701,N_6576);
or U8190 (N_8190,N_6865,N_7824);
xor U8191 (N_8191,N_7477,N_7009);
nand U8192 (N_8192,N_7002,N_7096);
xor U8193 (N_8193,N_6216,N_6814);
nor U8194 (N_8194,N_6399,N_7115);
or U8195 (N_8195,N_7524,N_7917);
nor U8196 (N_8196,N_7985,N_6051);
and U8197 (N_8197,N_7503,N_6984);
xnor U8198 (N_8198,N_6431,N_7242);
or U8199 (N_8199,N_7490,N_6506);
nor U8200 (N_8200,N_7698,N_7310);
xnor U8201 (N_8201,N_7314,N_6052);
and U8202 (N_8202,N_7591,N_7847);
nand U8203 (N_8203,N_7462,N_7790);
nand U8204 (N_8204,N_6945,N_6731);
or U8205 (N_8205,N_7400,N_6847);
nor U8206 (N_8206,N_6445,N_6873);
and U8207 (N_8207,N_6876,N_7815);
nand U8208 (N_8208,N_7181,N_6939);
and U8209 (N_8209,N_6702,N_6357);
and U8210 (N_8210,N_7593,N_6591);
nand U8211 (N_8211,N_7852,N_6351);
nand U8212 (N_8212,N_7595,N_7784);
nor U8213 (N_8213,N_6239,N_6326);
and U8214 (N_8214,N_7728,N_6567);
nor U8215 (N_8215,N_6841,N_7773);
nor U8216 (N_8216,N_6153,N_6684);
or U8217 (N_8217,N_6378,N_7257);
and U8218 (N_8218,N_6668,N_7508);
nand U8219 (N_8219,N_7057,N_7144);
or U8220 (N_8220,N_6665,N_6388);
or U8221 (N_8221,N_6203,N_6065);
or U8222 (N_8222,N_6615,N_7030);
nor U8223 (N_8223,N_7692,N_6906);
nand U8224 (N_8224,N_6441,N_6579);
nand U8225 (N_8225,N_7991,N_6913);
xnor U8226 (N_8226,N_7166,N_6757);
and U8227 (N_8227,N_6016,N_6741);
and U8228 (N_8228,N_7936,N_7643);
nand U8229 (N_8229,N_6341,N_6805);
and U8230 (N_8230,N_6206,N_7986);
and U8231 (N_8231,N_7020,N_6095);
nor U8232 (N_8232,N_7325,N_6584);
xnor U8233 (N_8233,N_7649,N_6967);
nand U8234 (N_8234,N_6932,N_7835);
or U8235 (N_8235,N_6067,N_7699);
nand U8236 (N_8236,N_6819,N_7557);
nor U8237 (N_8237,N_6526,N_6878);
nand U8238 (N_8238,N_6722,N_7972);
xor U8239 (N_8239,N_7390,N_7656);
and U8240 (N_8240,N_6711,N_6461);
nor U8241 (N_8241,N_6405,N_6572);
nor U8242 (N_8242,N_7909,N_7820);
and U8243 (N_8243,N_7928,N_7234);
xor U8244 (N_8244,N_6550,N_7043);
nor U8245 (N_8245,N_6240,N_7029);
nand U8246 (N_8246,N_6735,N_7762);
or U8247 (N_8247,N_7313,N_6466);
or U8248 (N_8248,N_6910,N_6385);
nand U8249 (N_8249,N_7089,N_6086);
nand U8250 (N_8250,N_7770,N_7911);
xnor U8251 (N_8251,N_6599,N_7869);
xor U8252 (N_8252,N_7258,N_7353);
nand U8253 (N_8253,N_7538,N_7263);
and U8254 (N_8254,N_6022,N_6650);
and U8255 (N_8255,N_7405,N_6302);
or U8256 (N_8256,N_6126,N_6091);
nor U8257 (N_8257,N_7001,N_6866);
nor U8258 (N_8258,N_7266,N_7159);
nor U8259 (N_8259,N_7114,N_6657);
or U8260 (N_8260,N_6487,N_7058);
xnor U8261 (N_8261,N_7348,N_6017);
xnor U8262 (N_8262,N_7129,N_6332);
nand U8263 (N_8263,N_6081,N_7806);
xnor U8264 (N_8264,N_6268,N_7705);
nand U8265 (N_8265,N_7401,N_6557);
and U8266 (N_8266,N_6877,N_6513);
xor U8267 (N_8267,N_6271,N_7411);
xor U8268 (N_8268,N_7444,N_6829);
nand U8269 (N_8269,N_6952,N_6620);
or U8270 (N_8270,N_6902,N_6142);
xnor U8271 (N_8271,N_7920,N_6468);
nand U8272 (N_8272,N_6233,N_6769);
nand U8273 (N_8273,N_7415,N_7918);
and U8274 (N_8274,N_6563,N_6089);
nand U8275 (N_8275,N_7466,N_7316);
nand U8276 (N_8276,N_6060,N_7796);
or U8277 (N_8277,N_6777,N_7324);
xor U8278 (N_8278,N_7101,N_7333);
xnor U8279 (N_8279,N_7533,N_7134);
xor U8280 (N_8280,N_7844,N_6654);
and U8281 (N_8281,N_7327,N_6088);
or U8282 (N_8282,N_7998,N_6238);
xnor U8283 (N_8283,N_7890,N_7668);
nor U8284 (N_8284,N_7260,N_7535);
or U8285 (N_8285,N_6672,N_6083);
xnor U8286 (N_8286,N_6215,N_7719);
nor U8287 (N_8287,N_6141,N_7048);
nor U8288 (N_8288,N_7878,N_7369);
nand U8289 (N_8289,N_6785,N_6803);
nand U8290 (N_8290,N_7204,N_7461);
nor U8291 (N_8291,N_6717,N_7756);
nand U8292 (N_8292,N_6315,N_6080);
or U8293 (N_8293,N_7504,N_6337);
or U8294 (N_8294,N_6692,N_7850);
and U8295 (N_8295,N_6170,N_6664);
xnor U8296 (N_8296,N_7307,N_7956);
nor U8297 (N_8297,N_6783,N_6604);
xnor U8298 (N_8298,N_6760,N_7975);
or U8299 (N_8299,N_7265,N_7989);
and U8300 (N_8300,N_6130,N_6755);
nand U8301 (N_8301,N_7385,N_6313);
or U8302 (N_8302,N_6174,N_7357);
nand U8303 (N_8303,N_7638,N_6977);
nor U8304 (N_8304,N_7299,N_6344);
nand U8305 (N_8305,N_7397,N_7826);
xor U8306 (N_8306,N_6403,N_6275);
and U8307 (N_8307,N_6761,N_6798);
nand U8308 (N_8308,N_7546,N_7330);
nor U8309 (N_8309,N_7544,N_6122);
nor U8310 (N_8310,N_6031,N_7782);
and U8311 (N_8311,N_7210,N_7870);
or U8312 (N_8312,N_6661,N_6690);
nand U8313 (N_8313,N_7996,N_6391);
nor U8314 (N_8314,N_6260,N_6662);
nor U8315 (N_8315,N_7537,N_6166);
and U8316 (N_8316,N_7893,N_6160);
nand U8317 (N_8317,N_6926,N_7218);
nor U8318 (N_8318,N_7269,N_6698);
and U8319 (N_8319,N_6172,N_7302);
or U8320 (N_8320,N_7498,N_6109);
or U8321 (N_8321,N_6049,N_6087);
or U8322 (N_8322,N_7064,N_7808);
and U8323 (N_8323,N_7262,N_7787);
or U8324 (N_8324,N_6383,N_6851);
nand U8325 (N_8325,N_7969,N_7099);
xnor U8326 (N_8326,N_6439,N_7843);
nand U8327 (N_8327,N_7216,N_6446);
and U8328 (N_8328,N_6077,N_6243);
nand U8329 (N_8329,N_6780,N_7296);
xor U8330 (N_8330,N_6801,N_6414);
xnor U8331 (N_8331,N_6053,N_6840);
or U8332 (N_8332,N_6842,N_6295);
or U8333 (N_8333,N_6976,N_6640);
nand U8334 (N_8334,N_7182,N_7799);
nor U8335 (N_8335,N_6618,N_6528);
xnor U8336 (N_8336,N_6343,N_7073);
or U8337 (N_8337,N_6966,N_6246);
xor U8338 (N_8338,N_7631,N_6021);
or U8339 (N_8339,N_7515,N_7209);
or U8340 (N_8340,N_6019,N_7905);
and U8341 (N_8341,N_7623,N_7577);
xnor U8342 (N_8342,N_7338,N_6889);
nand U8343 (N_8343,N_6636,N_6960);
and U8344 (N_8344,N_7514,N_6727);
nand U8345 (N_8345,N_7885,N_7054);
or U8346 (N_8346,N_7188,N_6467);
or U8347 (N_8347,N_6486,N_6208);
xnor U8348 (N_8348,N_6407,N_7988);
nand U8349 (N_8349,N_7737,N_7902);
xor U8350 (N_8350,N_6425,N_7713);
nand U8351 (N_8351,N_6492,N_7876);
nor U8352 (N_8352,N_7873,N_7382);
xnor U8353 (N_8353,N_7050,N_7285);
and U8354 (N_8354,N_6905,N_7422);
nor U8355 (N_8355,N_7388,N_6836);
nor U8356 (N_8356,N_7798,N_7027);
nand U8357 (N_8357,N_7249,N_6258);
or U8358 (N_8358,N_6578,N_6322);
nor U8359 (N_8359,N_7819,N_7128);
and U8360 (N_8360,N_7748,N_7007);
nor U8361 (N_8361,N_6361,N_7446);
and U8362 (N_8362,N_6002,N_6951);
xor U8363 (N_8363,N_6788,N_7380);
nand U8364 (N_8364,N_7571,N_6147);
nor U8365 (N_8365,N_6641,N_6773);
xor U8366 (N_8366,N_6651,N_7907);
xor U8367 (N_8367,N_6912,N_7959);
or U8368 (N_8368,N_7809,N_7028);
nand U8369 (N_8369,N_7880,N_6306);
and U8370 (N_8370,N_7560,N_6990);
and U8371 (N_8371,N_7410,N_6882);
nand U8372 (N_8372,N_6003,N_6230);
xnor U8373 (N_8373,N_6325,N_6568);
and U8374 (N_8374,N_6420,N_7116);
and U8375 (N_8375,N_7034,N_6879);
nor U8376 (N_8376,N_6642,N_7207);
xor U8377 (N_8377,N_6144,N_7085);
nor U8378 (N_8378,N_6064,N_6541);
nor U8379 (N_8379,N_6888,N_6303);
nor U8380 (N_8380,N_6794,N_7214);
nand U8381 (N_8381,N_7647,N_7232);
and U8382 (N_8382,N_6456,N_6368);
xor U8383 (N_8383,N_7513,N_7200);
nand U8384 (N_8384,N_6340,N_7662);
nor U8385 (N_8385,N_6059,N_6533);
and U8386 (N_8386,N_6234,N_7681);
or U8387 (N_8387,N_6408,N_7251);
nand U8388 (N_8388,N_6390,N_6936);
xnor U8389 (N_8389,N_7279,N_6892);
nand U8390 (N_8390,N_6029,N_7375);
nor U8391 (N_8391,N_7725,N_6292);
and U8392 (N_8392,N_7871,N_7614);
xor U8393 (N_8393,N_7293,N_6276);
xnor U8394 (N_8394,N_6581,N_6762);
xor U8395 (N_8395,N_6135,N_7939);
or U8396 (N_8396,N_6307,N_6078);
nand U8397 (N_8397,N_7982,N_7825);
xor U8398 (N_8398,N_7532,N_7669);
or U8399 (N_8399,N_6843,N_6443);
nand U8400 (N_8400,N_6281,N_6502);
nor U8401 (N_8401,N_7500,N_6143);
or U8402 (N_8402,N_7688,N_7914);
nor U8403 (N_8403,N_7882,N_7331);
nor U8404 (N_8404,N_7063,N_6666);
and U8405 (N_8405,N_6891,N_7761);
xnor U8406 (N_8406,N_7076,N_6765);
nand U8407 (N_8407,N_6860,N_6715);
xnor U8408 (N_8408,N_7923,N_6647);
or U8409 (N_8409,N_6247,N_6071);
or U8410 (N_8410,N_7836,N_7686);
nand U8411 (N_8411,N_6023,N_6084);
xnor U8412 (N_8412,N_7441,N_7903);
and U8413 (N_8413,N_7056,N_6061);
xnor U8414 (N_8414,N_7789,N_7225);
nand U8415 (N_8415,N_6532,N_6511);
or U8416 (N_8416,N_6124,N_7090);
nand U8417 (N_8417,N_6531,N_6729);
or U8418 (N_8418,N_6623,N_6373);
xor U8419 (N_8419,N_7901,N_7765);
xor U8420 (N_8420,N_6638,N_7543);
and U8421 (N_8421,N_7603,N_6044);
or U8422 (N_8422,N_7690,N_6352);
nor U8423 (N_8423,N_7526,N_7139);
or U8424 (N_8424,N_7460,N_7019);
xor U8425 (N_8425,N_7394,N_7039);
nor U8426 (N_8426,N_7764,N_7729);
xor U8427 (N_8427,N_6188,N_7341);
xnor U8428 (N_8428,N_7220,N_7493);
and U8429 (N_8429,N_6245,N_7700);
nand U8430 (N_8430,N_7592,N_7555);
nor U8431 (N_8431,N_7687,N_7111);
nor U8432 (N_8432,N_7103,N_7797);
nor U8433 (N_8433,N_6479,N_6367);
nor U8434 (N_8434,N_6041,N_7754);
nand U8435 (N_8435,N_6475,N_7345);
xor U8436 (N_8436,N_6288,N_7123);
nor U8437 (N_8437,N_6335,N_7837);
nor U8438 (N_8438,N_6110,N_6809);
and U8439 (N_8439,N_6540,N_6759);
xnor U8440 (N_8440,N_7981,N_6595);
xnor U8441 (N_8441,N_7280,N_7255);
xor U8442 (N_8442,N_7661,N_7724);
and U8443 (N_8443,N_6687,N_6252);
nand U8444 (N_8444,N_6489,N_6736);
and U8445 (N_8445,N_6074,N_7842);
or U8446 (N_8446,N_7359,N_7177);
or U8447 (N_8447,N_6434,N_7191);
and U8448 (N_8448,N_6947,N_7010);
and U8449 (N_8449,N_6159,N_6321);
and U8450 (N_8450,N_7223,N_7884);
nor U8451 (N_8451,N_7800,N_7420);
xnor U8452 (N_8452,N_6046,N_6560);
xor U8453 (N_8453,N_6725,N_6701);
or U8454 (N_8454,N_6462,N_7202);
and U8455 (N_8455,N_7977,N_6732);
xnor U8456 (N_8456,N_7672,N_7448);
or U8457 (N_8457,N_7004,N_6911);
nand U8458 (N_8458,N_6432,N_7601);
or U8459 (N_8459,N_7140,N_6721);
nor U8460 (N_8460,N_6555,N_6063);
and U8461 (N_8461,N_7426,N_6152);
xnor U8462 (N_8462,N_7747,N_7957);
or U8463 (N_8463,N_7423,N_7624);
nand U8464 (N_8464,N_7215,N_6035);
or U8465 (N_8465,N_6106,N_7340);
and U8466 (N_8466,N_7051,N_6808);
and U8467 (N_8467,N_7172,N_7021);
and U8468 (N_8468,N_7135,N_7752);
and U8469 (N_8469,N_6619,N_6094);
and U8470 (N_8470,N_6938,N_6828);
xor U8471 (N_8471,N_7339,N_6609);
and U8472 (N_8472,N_6248,N_7628);
or U8473 (N_8473,N_7095,N_7617);
nor U8474 (N_8474,N_7642,N_7944);
nor U8475 (N_8475,N_7696,N_7608);
nand U8476 (N_8476,N_7952,N_7464);
xor U8477 (N_8477,N_6293,N_7625);
and U8478 (N_8478,N_6696,N_6566);
and U8479 (N_8479,N_7562,N_6232);
nand U8480 (N_8480,N_7286,N_7112);
or U8481 (N_8481,N_6499,N_7987);
nor U8482 (N_8482,N_7803,N_7120);
nor U8483 (N_8483,N_6683,N_6658);
and U8484 (N_8484,N_7100,N_6012);
or U8485 (N_8485,N_6132,N_6509);
and U8486 (N_8486,N_6256,N_7463);
and U8487 (N_8487,N_6112,N_7206);
xnor U8488 (N_8488,N_7008,N_6688);
and U8489 (N_8489,N_7547,N_6259);
and U8490 (N_8490,N_7467,N_6830);
or U8491 (N_8491,N_7292,N_6946);
and U8492 (N_8492,N_7968,N_7726);
or U8493 (N_8493,N_6393,N_7113);
xnor U8494 (N_8494,N_7413,N_7127);
xnor U8495 (N_8495,N_6085,N_7781);
nor U8496 (N_8496,N_6719,N_7680);
xnor U8497 (N_8497,N_6386,N_7983);
nand U8498 (N_8498,N_6995,N_6987);
and U8499 (N_8499,N_7832,N_6018);
or U8500 (N_8500,N_6708,N_7716);
and U8501 (N_8501,N_7067,N_6534);
nor U8502 (N_8502,N_6916,N_7685);
and U8503 (N_8503,N_6667,N_6999);
or U8504 (N_8504,N_7501,N_6497);
nand U8505 (N_8505,N_7621,N_7606);
xnor U8506 (N_8506,N_6072,N_6048);
nor U8507 (N_8507,N_7276,N_7077);
or U8508 (N_8508,N_7006,N_6169);
nand U8509 (N_8509,N_7241,N_6707);
or U8510 (N_8510,N_6370,N_6376);
nor U8511 (N_8511,N_7875,N_6073);
and U8512 (N_8512,N_6544,N_7185);
nor U8513 (N_8513,N_6177,N_7678);
nor U8514 (N_8514,N_7270,N_6369);
or U8515 (N_8515,N_6483,N_6543);
nand U8516 (N_8516,N_7966,N_6723);
nand U8517 (N_8517,N_6875,N_7552);
nand U8518 (N_8518,N_7641,N_6603);
nand U8519 (N_8519,N_6249,N_6342);
nand U8520 (N_8520,N_7118,N_6409);
nor U8521 (N_8521,N_7169,N_6222);
nor U8522 (N_8522,N_6624,N_7497);
xor U8523 (N_8523,N_6058,N_7646);
nand U8524 (N_8524,N_7582,N_6438);
and U8525 (N_8525,N_7531,N_7679);
or U8526 (N_8526,N_7473,N_6384);
nand U8527 (N_8527,N_6927,N_6225);
nor U8528 (N_8528,N_7457,N_6140);
or U8529 (N_8529,N_7677,N_6396);
xnor U8530 (N_8530,N_6310,N_7160);
nand U8531 (N_8531,N_7419,N_6776);
and U8532 (N_8532,N_6269,N_6101);
and U8533 (N_8533,N_7153,N_6627);
nand U8534 (N_8534,N_6887,N_6955);
nor U8535 (N_8535,N_7356,N_7743);
nor U8536 (N_8536,N_6899,N_6154);
and U8537 (N_8537,N_6931,N_6745);
nor U8538 (N_8538,N_6107,N_6193);
xnor U8539 (N_8539,N_6201,N_6605);
and U8540 (N_8540,N_6831,N_6339);
or U8541 (N_8541,N_6845,N_7328);
or U8542 (N_8542,N_6975,N_6227);
nand U8543 (N_8543,N_6395,N_7271);
nand U8544 (N_8544,N_7946,N_6593);
and U8545 (N_8545,N_7398,N_7201);
or U8546 (N_8546,N_6637,N_6300);
xor U8547 (N_8547,N_7091,N_7634);
xnor U8548 (N_8548,N_6855,N_7636);
or U8549 (N_8549,N_6592,N_7243);
nor U8550 (N_8550,N_7187,N_6184);
or U8551 (N_8551,N_7440,N_6942);
and U8552 (N_8552,N_7447,N_7087);
nand U8553 (N_8553,N_6180,N_7916);
and U8554 (N_8554,N_6535,N_6418);
and U8555 (N_8555,N_6054,N_6104);
nand U8556 (N_8556,N_7407,N_6274);
nor U8557 (N_8557,N_6720,N_6660);
nand U8558 (N_8558,N_6484,N_7906);
and U8559 (N_8559,N_6382,N_6111);
nand U8560 (N_8560,N_6377,N_6312);
and U8561 (N_8561,N_6784,N_7282);
nand U8562 (N_8562,N_7335,N_6996);
nand U8563 (N_8563,N_7583,N_6807);
and U8564 (N_8564,N_6387,N_7675);
nand U8565 (N_8565,N_6204,N_7237);
and U8566 (N_8566,N_7471,N_6874);
nor U8567 (N_8567,N_7084,N_7605);
nor U8568 (N_8568,N_7630,N_6503);
or U8569 (N_8569,N_7267,N_6304);
and U8570 (N_8570,N_7492,N_6674);
xnor U8571 (N_8571,N_7502,N_7336);
nand U8572 (N_8572,N_7465,N_6800);
xor U8573 (N_8573,N_6398,N_6766);
nand U8574 (N_8574,N_7306,N_6614);
nand U8575 (N_8575,N_7810,N_6748);
or U8576 (N_8576,N_7749,N_7040);
and U8577 (N_8577,N_6827,N_7037);
xnor U8578 (N_8578,N_6490,N_6354);
xor U8579 (N_8579,N_7165,N_7435);
and U8580 (N_8580,N_7235,N_6822);
xnor U8581 (N_8581,N_6149,N_7731);
nor U8582 (N_8582,N_6940,N_6770);
or U8583 (N_8583,N_6301,N_7626);
nand U8584 (N_8584,N_7767,N_7291);
nand U8585 (N_8585,N_6458,N_6504);
nand U8586 (N_8586,N_6552,N_6190);
or U8587 (N_8587,N_7470,N_6789);
and U8588 (N_8588,N_7607,N_7409);
nand U8589 (N_8589,N_7478,N_7052);
nand U8590 (N_8590,N_7660,N_7012);
or U8591 (N_8591,N_6474,N_6324);
nor U8592 (N_8592,N_6833,N_7963);
xnor U8593 (N_8593,N_7199,N_7155);
nand U8594 (N_8594,N_6838,N_7418);
or U8595 (N_8595,N_6459,N_7246);
and U8596 (N_8596,N_6898,N_6070);
and U8597 (N_8597,N_6481,N_7580);
nand U8598 (N_8598,N_6435,N_7910);
nor U8599 (N_8599,N_6505,N_6036);
and U8600 (N_8600,N_7289,N_7629);
or U8601 (N_8601,N_7221,N_6114);
and U8602 (N_8602,N_6849,N_6699);
or U8603 (N_8603,N_7229,N_7588);
nor U8604 (N_8604,N_7733,N_7060);
and U8605 (N_8605,N_6196,N_7590);
or U8606 (N_8606,N_7813,N_7704);
and U8607 (N_8607,N_6392,N_6918);
xnor U8608 (N_8608,N_6694,N_7468);
or U8609 (N_8609,N_6539,N_7708);
nor U8610 (N_8610,N_6189,N_6753);
and U8611 (N_8611,N_6779,N_6937);
nor U8612 (N_8612,N_7042,N_6596);
or U8613 (N_8613,N_6451,N_6038);
or U8614 (N_8614,N_6825,N_7757);
xnor U8615 (N_8615,N_6772,N_6209);
and U8616 (N_8616,N_7841,N_6096);
and U8617 (N_8617,N_6482,N_7429);
nor U8618 (N_8618,N_6934,N_6097);
nand U8619 (N_8619,N_6102,N_6205);
xor U8620 (N_8620,N_6285,N_6496);
or U8621 (N_8621,N_7587,N_6677);
nand U8622 (N_8622,N_6251,N_6575);
nor U8623 (N_8623,N_7834,N_6969);
nand U8624 (N_8624,N_7802,N_6537);
and U8625 (N_8625,N_7620,N_7156);
nand U8626 (N_8626,N_6349,N_6673);
nor U8627 (N_8627,N_6909,N_6167);
nand U8628 (N_8628,N_7550,N_7812);
xor U8629 (N_8629,N_7107,N_7517);
or U8630 (N_8630,N_7055,N_7999);
nor U8631 (N_8631,N_7203,N_7211);
nand U8632 (N_8632,N_7141,N_6832);
nand U8633 (N_8633,N_6235,N_6298);
xnor U8634 (N_8634,N_7639,N_6818);
and U8635 (N_8635,N_7976,N_7071);
xor U8636 (N_8636,N_7000,N_7162);
xor U8637 (N_8637,N_6639,N_7995);
and U8638 (N_8638,N_7442,N_6622);
or U8639 (N_8639,N_7025,N_7654);
xor U8640 (N_8640,N_7569,N_7412);
xor U8641 (N_8641,N_6020,N_7970);
xor U8642 (N_8642,N_6372,N_7321);
nor U8643 (N_8643,N_7732,N_7945);
or U8644 (N_8644,N_6450,N_6728);
or U8645 (N_8645,N_7264,N_7253);
xnor U8646 (N_8646,N_7358,N_7712);
or U8647 (N_8647,N_7707,N_7102);
nor U8648 (N_8648,N_7453,N_6194);
and U8649 (N_8649,N_6237,N_7031);
or U8650 (N_8650,N_7604,N_7919);
or U8651 (N_8651,N_6314,N_7428);
nor U8652 (N_8652,N_6146,N_6449);
xor U8653 (N_8653,N_7152,N_6223);
nand U8654 (N_8654,N_7032,N_6191);
nor U8655 (N_8655,N_6994,N_7510);
nor U8656 (N_8656,N_7943,N_7193);
and U8657 (N_8657,N_7231,N_6774);
nand U8658 (N_8658,N_6704,N_6959);
xor U8659 (N_8659,N_7014,N_7540);
nand U8660 (N_8660,N_6473,N_6270);
nor U8661 (N_8661,N_6371,N_6971);
nor U8662 (N_8662,N_7791,N_7597);
xnor U8663 (N_8663,N_7300,N_7671);
and U8664 (N_8664,N_6956,N_7635);
and U8665 (N_8665,N_7776,N_6925);
or U8666 (N_8666,N_6116,N_7268);
nand U8667 (N_8667,N_6261,N_7763);
nor U8668 (N_8668,N_6810,N_7779);
nand U8669 (N_8669,N_7003,N_6954);
nand U8670 (N_8670,N_6663,N_7383);
xor U8671 (N_8671,N_7534,N_7433);
or U8672 (N_8672,N_7573,N_6123);
and U8673 (N_8673,N_7488,N_7178);
and U8674 (N_8674,N_7074,N_7322);
nand U8675 (N_8675,N_6601,N_6869);
xor U8676 (N_8676,N_7132,N_6212);
xnor U8677 (N_8677,N_6010,N_6796);
xnor U8678 (N_8678,N_7658,N_6360);
nand U8679 (N_8679,N_6941,N_7602);
nor U8680 (N_8680,N_7117,N_6374);
and U8681 (N_8681,N_7305,N_6338);
or U8682 (N_8682,N_7840,N_6476);
nand U8683 (N_8683,N_7892,N_7912);
and U8684 (N_8684,N_7512,N_7650);
or U8685 (N_8685,N_6015,N_6935);
nor U8686 (N_8686,N_7247,N_6908);
or U8687 (N_8687,N_6055,N_6470);
nor U8688 (N_8688,N_6726,N_6182);
and U8689 (N_8689,N_7097,N_7971);
xor U8690 (N_8690,N_6397,N_7176);
xor U8691 (N_8691,N_6455,N_6895);
and U8692 (N_8692,N_6066,N_6621);
nor U8693 (N_8693,N_6634,N_7958);
xnor U8694 (N_8694,N_6610,N_6680);
nand U8695 (N_8695,N_7424,N_6930);
and U8696 (N_8696,N_6214,N_6861);
and U8697 (N_8697,N_6904,N_7684);
xnor U8698 (N_8698,N_7829,N_6635);
xnor U8699 (N_8699,N_7586,N_6355);
nand U8700 (N_8700,N_6426,N_6973);
and U8701 (N_8701,N_6272,N_7072);
xor U8702 (N_8702,N_7168,N_6075);
nor U8703 (N_8703,N_7205,N_6671);
nor U8704 (N_8704,N_7370,N_6254);
nor U8705 (N_8705,N_7665,N_7715);
and U8706 (N_8706,N_7862,N_6009);
nor U8707 (N_8707,N_6914,N_6308);
nand U8708 (N_8708,N_7136,N_7298);
nand U8709 (N_8709,N_6291,N_6118);
or U8710 (N_8710,N_6617,N_7792);
xnor U8711 (N_8711,N_7469,N_7482);
or U8712 (N_8712,N_6198,N_6121);
xnor U8713 (N_8713,N_6423,N_6183);
or U8714 (N_8714,N_6323,N_7024);
nor U8715 (N_8715,N_6364,N_7702);
nand U8716 (N_8716,N_7794,N_7691);
xor U8717 (N_8717,N_7352,N_6613);
or U8718 (N_8718,N_7774,N_7891);
or U8719 (N_8719,N_6577,N_7536);
or U8720 (N_8720,N_7408,N_6522);
or U8721 (N_8721,N_7833,N_7736);
nand U8722 (N_8722,N_7549,N_6565);
nand U8723 (N_8723,N_7954,N_7804);
nand U8724 (N_8724,N_6286,N_7616);
and U8725 (N_8725,N_6853,N_7721);
nand U8726 (N_8726,N_6786,N_6583);
or U8727 (N_8727,N_7290,N_6430);
nand U8728 (N_8728,N_6795,N_6547);
nand U8729 (N_8729,N_7045,N_6844);
and U8730 (N_8730,N_6043,N_7142);
or U8731 (N_8731,N_6679,N_7859);
nor U8732 (N_8732,N_6319,N_6030);
and U8733 (N_8733,N_7277,N_7133);
nor U8734 (N_8734,N_6685,N_6488);
or U8735 (N_8735,N_7973,N_7250);
xnor U8736 (N_8736,N_6716,N_7682);
or U8737 (N_8737,N_7556,N_6406);
nand U8738 (N_8738,N_7430,N_7479);
or U8739 (N_8739,N_7189,N_6356);
nand U8740 (N_8740,N_7437,N_6359);
and U8741 (N_8741,N_7934,N_6394);
xor U8742 (N_8742,N_7342,N_6880);
or U8743 (N_8743,N_7755,N_6767);
xnor U8744 (N_8744,N_7443,N_6988);
nor U8745 (N_8745,N_7853,N_6014);
and U8746 (N_8746,N_6548,N_6607);
and U8747 (N_8747,N_7865,N_7745);
nand U8748 (N_8748,N_7572,N_7667);
nor U8749 (N_8749,N_6712,N_6718);
and U8750 (N_8750,N_7417,N_6962);
and U8751 (N_8751,N_7637,N_7485);
xor U8752 (N_8752,N_7974,N_6743);
xor U8753 (N_8753,N_6546,N_6764);
or U8754 (N_8754,N_7450,N_7511);
nand U8755 (N_8755,N_6099,N_6919);
nor U8756 (N_8756,N_7817,N_7894);
xnor U8757 (N_8757,N_6381,N_6013);
xor U8758 (N_8758,N_7811,N_7287);
nor U8759 (N_8759,N_6155,N_7238);
or U8760 (N_8760,N_6280,N_7551);
and U8761 (N_8761,N_6453,N_7822);
and U8762 (N_8762,N_7860,N_7778);
nand U8763 (N_8763,N_7275,N_7644);
and U8764 (N_8764,N_6471,N_6556);
and U8765 (N_8765,N_6520,N_6008);
xor U8766 (N_8766,N_7163,N_7312);
or U8767 (N_8767,N_7693,N_6185);
or U8768 (N_8768,N_6257,N_7184);
nor U8769 (N_8769,N_7640,N_7230);
nor U8770 (N_8770,N_7395,N_6655);
and U8771 (N_8771,N_7922,N_6244);
xor U8772 (N_8772,N_7777,N_7750);
nor U8773 (N_8773,N_6758,N_7746);
xnor U8774 (N_8774,N_7807,N_7013);
or U8775 (N_8775,N_7093,N_7518);
nor U8776 (N_8776,N_6079,N_7735);
xor U8777 (N_8777,N_7783,N_7887);
or U8778 (N_8778,N_7854,N_7760);
xor U8779 (N_8779,N_6695,N_7421);
xnor U8780 (N_8780,N_7788,N_6494);
or U8781 (N_8781,N_7427,N_6037);
or U8782 (N_8782,N_6958,N_6900);
nor U8783 (N_8783,N_7839,N_6156);
xnor U8784 (N_8784,N_6542,N_7297);
nand U8785 (N_8785,N_7244,N_7354);
or U8786 (N_8786,N_6864,N_6737);
xnor U8787 (N_8787,N_7131,N_6380);
or U8788 (N_8788,N_6691,N_7709);
and U8789 (N_8789,N_7472,N_7082);
nand U8790 (N_8790,N_6589,N_7655);
nand U8791 (N_8791,N_6137,N_6068);
nor U8792 (N_8792,N_7795,N_6922);
nor U8793 (N_8793,N_7506,N_7332);
nand U8794 (N_8794,N_6082,N_6594);
nand U8795 (N_8795,N_7683,N_7217);
xnor U8796 (N_8796,N_6127,N_6710);
and U8797 (N_8797,N_7079,N_7574);
or U8798 (N_8798,N_7886,N_6163);
and U8799 (N_8799,N_6210,N_7106);
nor U8800 (N_8800,N_6573,N_6705);
xor U8801 (N_8801,N_6858,N_6179);
nand U8802 (N_8802,N_6327,N_6317);
or U8803 (N_8803,N_7717,N_7589);
xnor U8804 (N_8804,N_7130,N_6480);
and U8805 (N_8805,N_7848,N_7391);
and U8806 (N_8806,N_7283,N_6812);
xnor U8807 (N_8807,N_6979,N_7921);
nand U8808 (N_8808,N_6848,N_6362);
or U8809 (N_8809,N_6602,N_6375);
nor U8810 (N_8810,N_7714,N_7558);
xnor U8811 (N_8811,N_6991,N_7366);
nand U8812 (N_8812,N_7362,N_6350);
and U8813 (N_8813,N_7718,N_7522);
nand U8814 (N_8814,N_7167,N_6815);
or U8815 (N_8815,N_6949,N_6982);
and U8816 (N_8816,N_6345,N_7967);
and U8817 (N_8817,N_7035,N_7449);
or U8818 (N_8818,N_7935,N_6463);
xnor U8819 (N_8819,N_7785,N_7396);
xnor U8820 (N_8820,N_7387,N_6559);
xor U8821 (N_8821,N_7425,N_6098);
and U8822 (N_8822,N_6554,N_6675);
and U8823 (N_8823,N_6920,N_6507);
and U8824 (N_8824,N_6413,N_6649);
xor U8825 (N_8825,N_7179,N_6948);
xor U8826 (N_8826,N_7827,N_7931);
and U8827 (N_8827,N_7722,N_6347);
nor U8828 (N_8828,N_7951,N_6186);
and U8829 (N_8829,N_7615,N_6739);
nor U8830 (N_8830,N_7281,N_6131);
xor U8831 (N_8831,N_7519,N_6564);
or U8832 (N_8832,N_6090,N_7005);
xor U8833 (N_8833,N_6040,N_7098);
nor U8834 (N_8834,N_7068,N_7738);
nand U8835 (N_8835,N_7350,N_7904);
xor U8836 (N_8836,N_7814,N_6820);
xor U8837 (N_8837,N_6771,N_6625);
nand U8838 (N_8838,N_7222,N_6477);
xnor U8839 (N_8839,N_6669,N_6981);
xor U8840 (N_8840,N_7541,N_6964);
nand U8841 (N_8841,N_6515,N_7105);
nor U8842 (N_8842,N_6255,N_7452);
nand U8843 (N_8843,N_7663,N_7295);
and U8844 (N_8844,N_6787,N_6799);
xor U8845 (N_8845,N_6076,N_6264);
nor U8846 (N_8846,N_7445,N_6517);
nor U8847 (N_8847,N_7143,N_7212);
and U8848 (N_8848,N_7771,N_6868);
nand U8849 (N_8849,N_6353,N_6448);
and U8850 (N_8850,N_6422,N_7252);
nand U8851 (N_8851,N_7288,N_7962);
xor U8852 (N_8852,N_7197,N_7780);
nand U8853 (N_8853,N_6460,N_7065);
nor U8854 (N_8854,N_7937,N_7367);
or U8855 (N_8855,N_6440,N_7772);
or U8856 (N_8856,N_7016,N_7753);
nand U8857 (N_8857,N_7304,N_7598);
xnor U8858 (N_8858,N_7775,N_6953);
nand U8859 (N_8859,N_7416,N_7585);
nor U8860 (N_8860,N_7319,N_6265);
and U8861 (N_8861,N_6454,N_6859);
or U8862 (N_8862,N_7053,N_7744);
nand U8863 (N_8863,N_6585,N_7294);
xnor U8864 (N_8864,N_6318,N_6250);
nor U8865 (N_8865,N_7092,N_7109);
nand U8866 (N_8866,N_6659,N_7233);
or U8867 (N_8867,N_6781,N_7648);
nor U8868 (N_8868,N_6972,N_7360);
nor U8869 (N_8869,N_6823,N_7964);
nor U8870 (N_8870,N_7786,N_6495);
or U8871 (N_8871,N_6519,N_7402);
xor U8872 (N_8872,N_7581,N_7320);
and U8873 (N_8873,N_7363,N_7311);
nand U8874 (N_8874,N_6173,N_7610);
nand U8875 (N_8875,N_7851,N_6646);
xnor U8876 (N_8876,N_7026,N_7611);
or U8877 (N_8877,N_6226,N_7858);
nor U8878 (N_8878,N_6901,N_6195);
nor U8879 (N_8879,N_6025,N_6491);
xor U8880 (N_8880,N_7877,N_7368);
and U8881 (N_8881,N_6993,N_7861);
xnor U8882 (N_8882,N_7727,N_6267);
nor U8883 (N_8883,N_7011,N_7436);
or U8884 (N_8884,N_6498,N_7554);
and U8885 (N_8885,N_6529,N_7364);
nor U8886 (N_8886,N_7022,N_7126);
nand U8887 (N_8887,N_6485,N_6612);
nand U8888 (N_8888,N_7406,N_7570);
and U8889 (N_8889,N_6197,N_7017);
nand U8890 (N_8890,N_7170,N_7404);
nand U8891 (N_8891,N_7066,N_7069);
nor U8892 (N_8892,N_7666,N_7379);
nor U8893 (N_8893,N_6026,N_6524);
or U8894 (N_8894,N_6273,N_6523);
nor U8895 (N_8895,N_6039,N_7337);
xnor U8896 (N_8896,N_6401,N_6284);
nor U8897 (N_8897,N_7653,N_7323);
nor U8898 (N_8898,N_7480,N_6590);
nand U8899 (N_8899,N_6366,N_6299);
and U8900 (N_8900,N_7703,N_7710);
xor U8901 (N_8901,N_7568,N_6582);
xnor U8902 (N_8902,N_6057,N_7104);
nand U8903 (N_8903,N_7414,N_7651);
and U8904 (N_8904,N_6652,N_7932);
nor U8905 (N_8905,N_6136,N_7183);
and U8906 (N_8906,N_7080,N_6569);
and U8907 (N_8907,N_7038,N_6791);
and U8908 (N_8908,N_7530,N_6586);
xnor U8909 (N_8909,N_7094,N_6811);
or U8910 (N_8910,N_6816,N_6328);
nor U8911 (N_8911,N_7256,N_7929);
and U8912 (N_8912,N_7872,N_7174);
nor U8913 (N_8913,N_6746,N_6706);
or U8914 (N_8914,N_7821,N_6644);
nand U8915 (N_8915,N_7499,N_6093);
or U8916 (N_8916,N_7484,N_6117);
nor U8917 (N_8917,N_7384,N_6266);
or U8918 (N_8918,N_6929,N_6600);
nand U8919 (N_8919,N_7164,N_7965);
or U8920 (N_8920,N_6219,N_6886);
xor U8921 (N_8921,N_7023,N_6536);
nand U8922 (N_8922,N_7676,N_7036);
xor U8923 (N_8923,N_6424,N_6419);
and U8924 (N_8924,N_6103,N_7627);
nand U8925 (N_8925,N_7613,N_7619);
nor U8926 (N_8926,N_7372,N_7553);
and U8927 (N_8927,N_7888,N_6763);
xnor U8928 (N_8928,N_6133,N_7864);
xor U8929 (N_8929,N_6733,N_7122);
and U8930 (N_8930,N_6656,N_6643);
and U8931 (N_8931,N_6870,N_7950);
nor U8932 (N_8932,N_6538,N_7622);
xnor U8933 (N_8933,N_7879,N_6756);
nor U8934 (N_8934,N_6200,N_7895);
nor U8935 (N_8935,N_7734,N_7376);
xnor U8936 (N_8936,N_6100,N_6000);
and U8937 (N_8937,N_7308,N_7309);
and U8938 (N_8938,N_6320,N_6228);
nand U8939 (N_8939,N_6862,N_7938);
nand U8940 (N_8940,N_6633,N_7224);
or U8941 (N_8941,N_6161,N_6730);
nor U8942 (N_8942,N_7491,N_7993);
nand U8943 (N_8943,N_6852,N_7451);
and U8944 (N_8944,N_7545,N_7831);
nand U8945 (N_8945,N_7459,N_6933);
xnor U8946 (N_8946,N_7565,N_7898);
xor U8947 (N_8947,N_6611,N_6826);
nor U8948 (N_8948,N_6069,N_6004);
nand U8949 (N_8949,N_7516,N_6970);
nand U8950 (N_8950,N_7883,N_6923);
or U8951 (N_8951,N_7481,N_6587);
or U8952 (N_8952,N_7365,N_6011);
xnor U8953 (N_8953,N_6628,N_6220);
nand U8954 (N_8954,N_6412,N_6211);
or U8955 (N_8955,N_6501,N_7434);
and U8956 (N_8956,N_6202,N_6872);
nor U8957 (N_8957,N_6290,N_6500);
nand U8958 (N_8958,N_6171,N_7600);
or U8959 (N_8959,N_7138,N_7845);
nor U8960 (N_8960,N_6330,N_7849);
xnor U8961 (N_8961,N_7818,N_6379);
xor U8962 (N_8962,N_7489,N_7086);
and U8963 (N_8963,N_6751,N_7070);
nor U8964 (N_8964,N_7475,N_6447);
and U8965 (N_8965,N_7213,N_7758);
nor U8966 (N_8966,N_7838,N_7278);
nand U8967 (N_8967,N_6178,N_7175);
xor U8968 (N_8968,N_7584,N_6346);
and U8969 (N_8969,N_6427,N_6309);
xnor U8970 (N_8970,N_6682,N_6115);
nor U8971 (N_8971,N_7180,N_7801);
and U8972 (N_8972,N_6139,N_7990);
or U8973 (N_8973,N_7866,N_7254);
or U8974 (N_8974,N_7227,N_6207);
and U8975 (N_8975,N_6700,N_6616);
nor U8976 (N_8976,N_7659,N_6608);
xnor U8977 (N_8977,N_6915,N_7361);
nor U8978 (N_8978,N_6978,N_7816);
and U8979 (N_8979,N_6598,N_7392);
and U8980 (N_8980,N_7044,N_6681);
xnor U8981 (N_8981,N_6928,N_6881);
nor U8982 (N_8982,N_7994,N_6469);
xor U8983 (N_8983,N_6514,N_6693);
xor U8984 (N_8984,N_6512,N_6411);
nor U8985 (N_8985,N_6997,N_7548);
and U8986 (N_8986,N_7377,N_6429);
or U8987 (N_8987,N_6924,N_7171);
xnor U8988 (N_8988,N_7856,N_6558);
nand U8989 (N_8989,N_6896,N_7695);
xor U8990 (N_8990,N_7897,N_7980);
or U8991 (N_8991,N_6229,N_6588);
xor U8992 (N_8992,N_6199,N_7476);
and U8993 (N_8993,N_6365,N_7896);
or U8994 (N_8994,N_7955,N_7151);
nor U8995 (N_8995,N_6389,N_6884);
xnor U8996 (N_8996,N_7374,N_7226);
and U8997 (N_8997,N_6033,N_6983);
and U8998 (N_8998,N_7261,N_6606);
xor U8999 (N_8999,N_7670,N_6871);
and U9000 (N_9000,N_7974,N_6735);
xor U9001 (N_9001,N_6426,N_6831);
nor U9002 (N_9002,N_7645,N_7940);
nor U9003 (N_9003,N_7837,N_7955);
xnor U9004 (N_9004,N_7282,N_7920);
nand U9005 (N_9005,N_7742,N_7183);
xor U9006 (N_9006,N_7470,N_6925);
nand U9007 (N_9007,N_7042,N_7610);
xor U9008 (N_9008,N_6468,N_7409);
and U9009 (N_9009,N_7993,N_6250);
or U9010 (N_9010,N_6568,N_7678);
and U9011 (N_9011,N_6536,N_7987);
nand U9012 (N_9012,N_6970,N_7330);
xnor U9013 (N_9013,N_6370,N_7276);
nand U9014 (N_9014,N_6243,N_7661);
nor U9015 (N_9015,N_7559,N_7549);
nand U9016 (N_9016,N_7297,N_7957);
nand U9017 (N_9017,N_7913,N_7655);
or U9018 (N_9018,N_6285,N_7505);
and U9019 (N_9019,N_6215,N_7347);
nor U9020 (N_9020,N_6458,N_7646);
xnor U9021 (N_9021,N_7234,N_7632);
and U9022 (N_9022,N_6389,N_7806);
xor U9023 (N_9023,N_7071,N_6138);
nand U9024 (N_9024,N_7441,N_7512);
xor U9025 (N_9025,N_7824,N_7459);
nor U9026 (N_9026,N_7005,N_6341);
and U9027 (N_9027,N_6552,N_7814);
or U9028 (N_9028,N_6403,N_7514);
or U9029 (N_9029,N_6496,N_6516);
xor U9030 (N_9030,N_7601,N_7707);
nand U9031 (N_9031,N_6019,N_6488);
nor U9032 (N_9032,N_6644,N_7226);
and U9033 (N_9033,N_6130,N_7179);
nor U9034 (N_9034,N_6338,N_7828);
nor U9035 (N_9035,N_7414,N_7275);
nor U9036 (N_9036,N_6144,N_7426);
and U9037 (N_9037,N_6694,N_6354);
nor U9038 (N_9038,N_6853,N_6182);
and U9039 (N_9039,N_7217,N_7803);
nand U9040 (N_9040,N_7242,N_6280);
nand U9041 (N_9041,N_7844,N_7574);
and U9042 (N_9042,N_6061,N_6016);
and U9043 (N_9043,N_6036,N_6942);
and U9044 (N_9044,N_7736,N_7771);
nor U9045 (N_9045,N_7043,N_6072);
or U9046 (N_9046,N_6446,N_6483);
or U9047 (N_9047,N_7656,N_6203);
nor U9048 (N_9048,N_6611,N_6957);
or U9049 (N_9049,N_7600,N_7250);
or U9050 (N_9050,N_6421,N_6446);
and U9051 (N_9051,N_7246,N_6938);
xnor U9052 (N_9052,N_6917,N_6880);
and U9053 (N_9053,N_6436,N_7821);
nand U9054 (N_9054,N_6970,N_7834);
xnor U9055 (N_9055,N_7318,N_7050);
and U9056 (N_9056,N_6770,N_7963);
xnor U9057 (N_9057,N_6227,N_7398);
nand U9058 (N_9058,N_6223,N_7394);
xor U9059 (N_9059,N_7156,N_7196);
nand U9060 (N_9060,N_6967,N_6088);
nor U9061 (N_9061,N_7739,N_7442);
nand U9062 (N_9062,N_7628,N_6719);
xnor U9063 (N_9063,N_6266,N_7014);
nand U9064 (N_9064,N_6894,N_6794);
and U9065 (N_9065,N_7830,N_6717);
nor U9066 (N_9066,N_6650,N_6209);
and U9067 (N_9067,N_6752,N_7036);
nand U9068 (N_9068,N_6086,N_6567);
nand U9069 (N_9069,N_6741,N_7400);
xnor U9070 (N_9070,N_7715,N_6285);
and U9071 (N_9071,N_7795,N_7729);
nand U9072 (N_9072,N_7852,N_6439);
nor U9073 (N_9073,N_6983,N_6699);
xor U9074 (N_9074,N_6331,N_6161);
and U9075 (N_9075,N_6458,N_6116);
nor U9076 (N_9076,N_6662,N_6683);
or U9077 (N_9077,N_6162,N_6998);
and U9078 (N_9078,N_6798,N_7636);
and U9079 (N_9079,N_6057,N_6679);
and U9080 (N_9080,N_7117,N_7107);
or U9081 (N_9081,N_7608,N_6459);
and U9082 (N_9082,N_6370,N_6927);
xor U9083 (N_9083,N_6841,N_7110);
nor U9084 (N_9084,N_6582,N_6675);
or U9085 (N_9085,N_7772,N_7854);
nand U9086 (N_9086,N_7350,N_7735);
or U9087 (N_9087,N_6162,N_7027);
xnor U9088 (N_9088,N_7392,N_6319);
and U9089 (N_9089,N_6698,N_7592);
nor U9090 (N_9090,N_6068,N_6545);
and U9091 (N_9091,N_7848,N_6660);
xnor U9092 (N_9092,N_6259,N_7873);
xor U9093 (N_9093,N_6341,N_6356);
nor U9094 (N_9094,N_6928,N_6598);
or U9095 (N_9095,N_6604,N_6076);
nand U9096 (N_9096,N_6974,N_6926);
xor U9097 (N_9097,N_6692,N_6832);
nor U9098 (N_9098,N_7751,N_7283);
xnor U9099 (N_9099,N_7268,N_6675);
or U9100 (N_9100,N_7725,N_7612);
or U9101 (N_9101,N_6246,N_6800);
xnor U9102 (N_9102,N_6258,N_7253);
and U9103 (N_9103,N_6406,N_6095);
or U9104 (N_9104,N_6344,N_7021);
and U9105 (N_9105,N_6001,N_7181);
or U9106 (N_9106,N_7899,N_7440);
or U9107 (N_9107,N_6527,N_6036);
nor U9108 (N_9108,N_6732,N_6044);
or U9109 (N_9109,N_7505,N_6078);
and U9110 (N_9110,N_7957,N_6282);
nor U9111 (N_9111,N_7808,N_7679);
and U9112 (N_9112,N_6567,N_7223);
or U9113 (N_9113,N_7460,N_6701);
xor U9114 (N_9114,N_7199,N_6945);
nand U9115 (N_9115,N_6297,N_6543);
xor U9116 (N_9116,N_7353,N_7144);
nor U9117 (N_9117,N_6499,N_6708);
and U9118 (N_9118,N_6052,N_7841);
nand U9119 (N_9119,N_7675,N_7459);
and U9120 (N_9120,N_7222,N_7190);
or U9121 (N_9121,N_7953,N_6364);
and U9122 (N_9122,N_6993,N_6431);
xor U9123 (N_9123,N_7589,N_6521);
or U9124 (N_9124,N_6629,N_7673);
or U9125 (N_9125,N_6493,N_7490);
or U9126 (N_9126,N_6581,N_6831);
nor U9127 (N_9127,N_7881,N_6912);
nor U9128 (N_9128,N_6595,N_6307);
nand U9129 (N_9129,N_7948,N_7898);
xnor U9130 (N_9130,N_6529,N_6841);
nor U9131 (N_9131,N_6972,N_6642);
nand U9132 (N_9132,N_6786,N_6133);
xor U9133 (N_9133,N_6136,N_6877);
xor U9134 (N_9134,N_6164,N_7832);
nand U9135 (N_9135,N_6751,N_6985);
nor U9136 (N_9136,N_6806,N_7236);
or U9137 (N_9137,N_7352,N_6338);
nor U9138 (N_9138,N_6669,N_7927);
nor U9139 (N_9139,N_7211,N_7305);
nor U9140 (N_9140,N_6383,N_6945);
nor U9141 (N_9141,N_6552,N_6023);
nand U9142 (N_9142,N_6361,N_7476);
nand U9143 (N_9143,N_7821,N_6484);
and U9144 (N_9144,N_6929,N_6568);
nand U9145 (N_9145,N_7484,N_7550);
nor U9146 (N_9146,N_7689,N_6868);
or U9147 (N_9147,N_7279,N_7043);
nand U9148 (N_9148,N_6088,N_6629);
xor U9149 (N_9149,N_6777,N_6961);
and U9150 (N_9150,N_6262,N_6639);
xnor U9151 (N_9151,N_7744,N_6413);
or U9152 (N_9152,N_7405,N_7468);
nand U9153 (N_9153,N_6151,N_6754);
xor U9154 (N_9154,N_6092,N_6375);
xor U9155 (N_9155,N_6695,N_6188);
nand U9156 (N_9156,N_7489,N_7617);
or U9157 (N_9157,N_6950,N_6706);
and U9158 (N_9158,N_6128,N_7322);
xor U9159 (N_9159,N_7205,N_6738);
nand U9160 (N_9160,N_7250,N_6046);
or U9161 (N_9161,N_6774,N_7532);
xor U9162 (N_9162,N_7742,N_7803);
xor U9163 (N_9163,N_6508,N_7207);
nand U9164 (N_9164,N_7509,N_7649);
nor U9165 (N_9165,N_7301,N_7199);
nor U9166 (N_9166,N_7927,N_6286);
and U9167 (N_9167,N_6848,N_6031);
nand U9168 (N_9168,N_6441,N_7518);
nand U9169 (N_9169,N_7646,N_7199);
and U9170 (N_9170,N_7426,N_7483);
and U9171 (N_9171,N_6198,N_7876);
and U9172 (N_9172,N_7993,N_7100);
nor U9173 (N_9173,N_6513,N_7597);
xnor U9174 (N_9174,N_6337,N_6586);
nor U9175 (N_9175,N_6232,N_7827);
nand U9176 (N_9176,N_7522,N_7763);
nand U9177 (N_9177,N_7452,N_6005);
or U9178 (N_9178,N_6357,N_6537);
or U9179 (N_9179,N_6317,N_7370);
and U9180 (N_9180,N_7851,N_6200);
nor U9181 (N_9181,N_6440,N_6703);
or U9182 (N_9182,N_6554,N_7429);
or U9183 (N_9183,N_6345,N_6205);
nor U9184 (N_9184,N_7782,N_6313);
nor U9185 (N_9185,N_7441,N_7465);
xnor U9186 (N_9186,N_7694,N_7679);
nand U9187 (N_9187,N_6573,N_7483);
and U9188 (N_9188,N_7025,N_6077);
nand U9189 (N_9189,N_6541,N_6687);
xnor U9190 (N_9190,N_7705,N_7898);
nand U9191 (N_9191,N_7241,N_7978);
or U9192 (N_9192,N_7496,N_7782);
and U9193 (N_9193,N_7600,N_6795);
xor U9194 (N_9194,N_6103,N_6344);
xor U9195 (N_9195,N_7614,N_7551);
xor U9196 (N_9196,N_6404,N_6096);
and U9197 (N_9197,N_6057,N_6204);
nand U9198 (N_9198,N_6499,N_6992);
nand U9199 (N_9199,N_7579,N_7297);
xnor U9200 (N_9200,N_6484,N_7203);
nand U9201 (N_9201,N_7369,N_7001);
nor U9202 (N_9202,N_6672,N_7309);
and U9203 (N_9203,N_7524,N_7617);
and U9204 (N_9204,N_7144,N_6556);
nand U9205 (N_9205,N_7521,N_6532);
or U9206 (N_9206,N_6932,N_6570);
nor U9207 (N_9207,N_6272,N_6842);
nor U9208 (N_9208,N_7196,N_7151);
or U9209 (N_9209,N_7206,N_7754);
xor U9210 (N_9210,N_6491,N_7999);
xor U9211 (N_9211,N_6780,N_6216);
and U9212 (N_9212,N_6250,N_6296);
and U9213 (N_9213,N_6705,N_7030);
xor U9214 (N_9214,N_7542,N_7685);
and U9215 (N_9215,N_7471,N_6950);
and U9216 (N_9216,N_7159,N_6752);
and U9217 (N_9217,N_6328,N_7829);
and U9218 (N_9218,N_6582,N_6443);
or U9219 (N_9219,N_6911,N_7239);
and U9220 (N_9220,N_7515,N_6015);
and U9221 (N_9221,N_6850,N_7326);
or U9222 (N_9222,N_6807,N_6867);
nand U9223 (N_9223,N_7870,N_6996);
nand U9224 (N_9224,N_7046,N_6285);
and U9225 (N_9225,N_7049,N_6253);
xor U9226 (N_9226,N_7317,N_7291);
and U9227 (N_9227,N_6340,N_7772);
nand U9228 (N_9228,N_6489,N_6237);
nand U9229 (N_9229,N_6179,N_6581);
xnor U9230 (N_9230,N_6749,N_6215);
xor U9231 (N_9231,N_7201,N_7048);
and U9232 (N_9232,N_6214,N_6468);
xnor U9233 (N_9233,N_6633,N_7616);
or U9234 (N_9234,N_6276,N_6524);
nor U9235 (N_9235,N_7634,N_6643);
xnor U9236 (N_9236,N_7781,N_6229);
nor U9237 (N_9237,N_6342,N_7357);
nor U9238 (N_9238,N_6051,N_6985);
xnor U9239 (N_9239,N_6024,N_7845);
nand U9240 (N_9240,N_7996,N_7918);
and U9241 (N_9241,N_7834,N_6311);
nor U9242 (N_9242,N_6052,N_7513);
nand U9243 (N_9243,N_6914,N_7552);
nand U9244 (N_9244,N_7455,N_6023);
or U9245 (N_9245,N_7741,N_7215);
or U9246 (N_9246,N_7798,N_7970);
nor U9247 (N_9247,N_7216,N_7353);
nand U9248 (N_9248,N_7256,N_7141);
nor U9249 (N_9249,N_6397,N_6514);
nand U9250 (N_9250,N_7531,N_6196);
nor U9251 (N_9251,N_6623,N_6948);
xnor U9252 (N_9252,N_7122,N_6732);
or U9253 (N_9253,N_7314,N_6266);
or U9254 (N_9254,N_6261,N_7592);
nand U9255 (N_9255,N_7526,N_7421);
and U9256 (N_9256,N_6503,N_7137);
or U9257 (N_9257,N_7725,N_7722);
nor U9258 (N_9258,N_6753,N_7629);
nand U9259 (N_9259,N_6421,N_7538);
nor U9260 (N_9260,N_7215,N_7253);
and U9261 (N_9261,N_6022,N_7620);
or U9262 (N_9262,N_6871,N_7312);
and U9263 (N_9263,N_6276,N_7386);
or U9264 (N_9264,N_7457,N_7551);
nor U9265 (N_9265,N_7618,N_6669);
and U9266 (N_9266,N_6158,N_7272);
xnor U9267 (N_9267,N_7289,N_6694);
or U9268 (N_9268,N_7374,N_7739);
xnor U9269 (N_9269,N_7968,N_7649);
xnor U9270 (N_9270,N_6388,N_7813);
and U9271 (N_9271,N_6560,N_6780);
or U9272 (N_9272,N_6137,N_7511);
nand U9273 (N_9273,N_7746,N_6163);
xor U9274 (N_9274,N_7657,N_6059);
xor U9275 (N_9275,N_6194,N_7415);
or U9276 (N_9276,N_6265,N_6982);
and U9277 (N_9277,N_6623,N_7430);
nand U9278 (N_9278,N_7196,N_6948);
or U9279 (N_9279,N_7058,N_6175);
nor U9280 (N_9280,N_6613,N_6222);
nor U9281 (N_9281,N_6083,N_7408);
and U9282 (N_9282,N_6510,N_6118);
nand U9283 (N_9283,N_7599,N_6091);
nand U9284 (N_9284,N_6961,N_6290);
nor U9285 (N_9285,N_7931,N_7789);
nor U9286 (N_9286,N_7523,N_6846);
or U9287 (N_9287,N_7458,N_7453);
or U9288 (N_9288,N_7373,N_6608);
or U9289 (N_9289,N_7838,N_7716);
and U9290 (N_9290,N_6865,N_6928);
nand U9291 (N_9291,N_6199,N_7558);
and U9292 (N_9292,N_7670,N_6764);
xnor U9293 (N_9293,N_6267,N_6842);
or U9294 (N_9294,N_7411,N_6455);
or U9295 (N_9295,N_7999,N_7896);
xnor U9296 (N_9296,N_7135,N_6848);
or U9297 (N_9297,N_7568,N_6794);
xor U9298 (N_9298,N_6186,N_7683);
or U9299 (N_9299,N_7208,N_6656);
and U9300 (N_9300,N_7695,N_6997);
or U9301 (N_9301,N_7880,N_7122);
or U9302 (N_9302,N_6931,N_6121);
nor U9303 (N_9303,N_6845,N_6412);
and U9304 (N_9304,N_6652,N_7054);
or U9305 (N_9305,N_6958,N_7604);
nor U9306 (N_9306,N_6537,N_6745);
nor U9307 (N_9307,N_7154,N_7824);
xor U9308 (N_9308,N_6307,N_7873);
or U9309 (N_9309,N_6884,N_7726);
xnor U9310 (N_9310,N_7466,N_7581);
or U9311 (N_9311,N_6306,N_6546);
or U9312 (N_9312,N_6539,N_7287);
and U9313 (N_9313,N_7936,N_7285);
and U9314 (N_9314,N_7698,N_6838);
or U9315 (N_9315,N_6022,N_6940);
nand U9316 (N_9316,N_6383,N_6720);
nor U9317 (N_9317,N_7130,N_7089);
or U9318 (N_9318,N_6391,N_6096);
or U9319 (N_9319,N_6597,N_7396);
nand U9320 (N_9320,N_6629,N_7883);
xnor U9321 (N_9321,N_6493,N_7726);
nor U9322 (N_9322,N_7103,N_7415);
nor U9323 (N_9323,N_6704,N_7514);
nand U9324 (N_9324,N_6757,N_6792);
nand U9325 (N_9325,N_6332,N_6580);
xnor U9326 (N_9326,N_6354,N_6402);
nand U9327 (N_9327,N_6772,N_6351);
nand U9328 (N_9328,N_6723,N_6965);
or U9329 (N_9329,N_7255,N_7006);
nor U9330 (N_9330,N_7781,N_7442);
nand U9331 (N_9331,N_6760,N_7779);
or U9332 (N_9332,N_7596,N_6258);
nor U9333 (N_9333,N_7325,N_6722);
and U9334 (N_9334,N_7695,N_6726);
and U9335 (N_9335,N_6542,N_7525);
xnor U9336 (N_9336,N_6412,N_6385);
nor U9337 (N_9337,N_7290,N_7797);
nor U9338 (N_9338,N_7882,N_7040);
or U9339 (N_9339,N_6578,N_7675);
nand U9340 (N_9340,N_6657,N_6356);
and U9341 (N_9341,N_7616,N_6652);
or U9342 (N_9342,N_7560,N_7175);
xor U9343 (N_9343,N_6439,N_7471);
or U9344 (N_9344,N_7328,N_7255);
xor U9345 (N_9345,N_6619,N_7581);
xor U9346 (N_9346,N_7486,N_7390);
nand U9347 (N_9347,N_7718,N_6357);
nand U9348 (N_9348,N_6581,N_7350);
and U9349 (N_9349,N_6954,N_7439);
xor U9350 (N_9350,N_7792,N_6278);
nor U9351 (N_9351,N_6359,N_7965);
nand U9352 (N_9352,N_7754,N_7479);
xnor U9353 (N_9353,N_7132,N_7304);
and U9354 (N_9354,N_7091,N_7386);
nor U9355 (N_9355,N_6452,N_6144);
xnor U9356 (N_9356,N_7462,N_6545);
nor U9357 (N_9357,N_7815,N_7540);
xor U9358 (N_9358,N_6676,N_6579);
xor U9359 (N_9359,N_7225,N_7127);
nand U9360 (N_9360,N_7643,N_6082);
nor U9361 (N_9361,N_6271,N_6375);
or U9362 (N_9362,N_6704,N_7046);
and U9363 (N_9363,N_6041,N_6046);
nand U9364 (N_9364,N_6249,N_6667);
nor U9365 (N_9365,N_7370,N_7340);
xnor U9366 (N_9366,N_6106,N_7250);
or U9367 (N_9367,N_7116,N_6538);
nor U9368 (N_9368,N_7006,N_7176);
nor U9369 (N_9369,N_6707,N_6032);
xor U9370 (N_9370,N_6775,N_7694);
or U9371 (N_9371,N_6548,N_7748);
nor U9372 (N_9372,N_6608,N_6440);
xor U9373 (N_9373,N_7491,N_7537);
and U9374 (N_9374,N_7949,N_6242);
nor U9375 (N_9375,N_6344,N_6852);
or U9376 (N_9376,N_7006,N_7132);
nand U9377 (N_9377,N_6416,N_6927);
nand U9378 (N_9378,N_6470,N_6729);
nor U9379 (N_9379,N_7463,N_7548);
and U9380 (N_9380,N_6982,N_6590);
or U9381 (N_9381,N_6739,N_6191);
xnor U9382 (N_9382,N_6490,N_6826);
and U9383 (N_9383,N_7233,N_7801);
nand U9384 (N_9384,N_6983,N_6480);
or U9385 (N_9385,N_7668,N_6230);
nor U9386 (N_9386,N_6626,N_6031);
xnor U9387 (N_9387,N_6291,N_7084);
nor U9388 (N_9388,N_7189,N_6294);
nand U9389 (N_9389,N_6701,N_7819);
nand U9390 (N_9390,N_6110,N_6272);
xor U9391 (N_9391,N_6879,N_7774);
nand U9392 (N_9392,N_6145,N_7108);
nor U9393 (N_9393,N_6242,N_6682);
xnor U9394 (N_9394,N_7000,N_7115);
or U9395 (N_9395,N_6339,N_6727);
nand U9396 (N_9396,N_6137,N_6947);
nand U9397 (N_9397,N_6059,N_6757);
nor U9398 (N_9398,N_7034,N_6753);
xor U9399 (N_9399,N_7770,N_6868);
xor U9400 (N_9400,N_6613,N_7720);
xor U9401 (N_9401,N_6544,N_7158);
nand U9402 (N_9402,N_7340,N_6995);
nand U9403 (N_9403,N_7296,N_7371);
and U9404 (N_9404,N_6992,N_6343);
nor U9405 (N_9405,N_6557,N_7657);
xnor U9406 (N_9406,N_7378,N_7588);
nand U9407 (N_9407,N_6773,N_6531);
or U9408 (N_9408,N_7604,N_6962);
and U9409 (N_9409,N_6267,N_7118);
nor U9410 (N_9410,N_7754,N_7844);
and U9411 (N_9411,N_6908,N_6230);
and U9412 (N_9412,N_6822,N_6542);
nor U9413 (N_9413,N_7357,N_6486);
nor U9414 (N_9414,N_7644,N_7224);
nor U9415 (N_9415,N_6671,N_6539);
xor U9416 (N_9416,N_7352,N_6589);
nor U9417 (N_9417,N_7850,N_6092);
nor U9418 (N_9418,N_6997,N_7371);
and U9419 (N_9419,N_6386,N_6546);
or U9420 (N_9420,N_6851,N_7214);
or U9421 (N_9421,N_7925,N_6965);
and U9422 (N_9422,N_7863,N_6453);
nor U9423 (N_9423,N_7863,N_7597);
nand U9424 (N_9424,N_7139,N_7398);
nor U9425 (N_9425,N_6821,N_7555);
nor U9426 (N_9426,N_6373,N_7973);
and U9427 (N_9427,N_6627,N_6540);
nand U9428 (N_9428,N_6386,N_6503);
or U9429 (N_9429,N_6522,N_6689);
nor U9430 (N_9430,N_7614,N_7576);
and U9431 (N_9431,N_6860,N_7061);
xor U9432 (N_9432,N_7551,N_7932);
nor U9433 (N_9433,N_6655,N_7304);
or U9434 (N_9434,N_6221,N_7207);
nor U9435 (N_9435,N_6362,N_6382);
and U9436 (N_9436,N_7693,N_6689);
xnor U9437 (N_9437,N_6804,N_6712);
or U9438 (N_9438,N_6412,N_6230);
or U9439 (N_9439,N_7697,N_7023);
nor U9440 (N_9440,N_6087,N_7541);
or U9441 (N_9441,N_6785,N_6462);
and U9442 (N_9442,N_6370,N_7555);
nand U9443 (N_9443,N_7320,N_7442);
xnor U9444 (N_9444,N_6177,N_6396);
or U9445 (N_9445,N_6673,N_7922);
and U9446 (N_9446,N_6765,N_7996);
and U9447 (N_9447,N_6464,N_6303);
or U9448 (N_9448,N_7377,N_6683);
xnor U9449 (N_9449,N_6332,N_6084);
nor U9450 (N_9450,N_6206,N_6165);
or U9451 (N_9451,N_7958,N_6255);
xnor U9452 (N_9452,N_7374,N_6884);
and U9453 (N_9453,N_7763,N_7090);
and U9454 (N_9454,N_7212,N_7285);
nor U9455 (N_9455,N_6553,N_6716);
xor U9456 (N_9456,N_6277,N_7545);
and U9457 (N_9457,N_6439,N_7137);
nor U9458 (N_9458,N_6465,N_7085);
and U9459 (N_9459,N_7836,N_6593);
xor U9460 (N_9460,N_7035,N_7578);
xor U9461 (N_9461,N_6031,N_7863);
nand U9462 (N_9462,N_6195,N_7244);
nor U9463 (N_9463,N_7578,N_7980);
xnor U9464 (N_9464,N_7419,N_7790);
nand U9465 (N_9465,N_6162,N_7148);
xnor U9466 (N_9466,N_6436,N_6903);
xnor U9467 (N_9467,N_7494,N_7781);
or U9468 (N_9468,N_6503,N_6249);
nor U9469 (N_9469,N_7419,N_6246);
nor U9470 (N_9470,N_7618,N_6668);
nor U9471 (N_9471,N_7400,N_6019);
and U9472 (N_9472,N_7305,N_7361);
nor U9473 (N_9473,N_7092,N_7921);
and U9474 (N_9474,N_7856,N_6174);
and U9475 (N_9475,N_7558,N_7823);
nand U9476 (N_9476,N_7280,N_6638);
nor U9477 (N_9477,N_6044,N_6261);
nor U9478 (N_9478,N_7161,N_7142);
nor U9479 (N_9479,N_6321,N_7931);
nand U9480 (N_9480,N_6092,N_7480);
xnor U9481 (N_9481,N_7879,N_6358);
nor U9482 (N_9482,N_6239,N_6608);
and U9483 (N_9483,N_6849,N_7754);
xor U9484 (N_9484,N_6567,N_6259);
and U9485 (N_9485,N_7036,N_6915);
nor U9486 (N_9486,N_6963,N_7591);
xor U9487 (N_9487,N_6412,N_6055);
nor U9488 (N_9488,N_6367,N_7160);
and U9489 (N_9489,N_6440,N_7192);
and U9490 (N_9490,N_7565,N_7497);
nand U9491 (N_9491,N_7391,N_6282);
and U9492 (N_9492,N_6387,N_6666);
nand U9493 (N_9493,N_6675,N_7027);
and U9494 (N_9494,N_7275,N_6884);
nand U9495 (N_9495,N_7412,N_7293);
nor U9496 (N_9496,N_7983,N_7736);
or U9497 (N_9497,N_7318,N_7964);
xnor U9498 (N_9498,N_6422,N_7974);
or U9499 (N_9499,N_6388,N_7088);
nor U9500 (N_9500,N_7317,N_6441);
or U9501 (N_9501,N_6909,N_6998);
and U9502 (N_9502,N_6188,N_7668);
nand U9503 (N_9503,N_7491,N_7602);
xor U9504 (N_9504,N_6250,N_6263);
nor U9505 (N_9505,N_7642,N_6186);
and U9506 (N_9506,N_7470,N_7843);
nor U9507 (N_9507,N_7083,N_6301);
nand U9508 (N_9508,N_6652,N_6539);
nor U9509 (N_9509,N_7438,N_7790);
and U9510 (N_9510,N_7590,N_6056);
or U9511 (N_9511,N_7667,N_7473);
xor U9512 (N_9512,N_6778,N_6192);
nand U9513 (N_9513,N_7847,N_7799);
xnor U9514 (N_9514,N_6795,N_7321);
xnor U9515 (N_9515,N_6793,N_7424);
or U9516 (N_9516,N_7758,N_7753);
or U9517 (N_9517,N_7995,N_6633);
or U9518 (N_9518,N_6884,N_6939);
nand U9519 (N_9519,N_7344,N_7540);
or U9520 (N_9520,N_6731,N_6801);
nor U9521 (N_9521,N_7984,N_6136);
or U9522 (N_9522,N_6990,N_7850);
and U9523 (N_9523,N_6547,N_6024);
nor U9524 (N_9524,N_6635,N_6398);
or U9525 (N_9525,N_7912,N_6368);
xnor U9526 (N_9526,N_6276,N_7552);
or U9527 (N_9527,N_7374,N_7404);
or U9528 (N_9528,N_7818,N_6354);
and U9529 (N_9529,N_7623,N_6028);
or U9530 (N_9530,N_6282,N_7555);
or U9531 (N_9531,N_6443,N_7067);
nand U9532 (N_9532,N_7876,N_7977);
nand U9533 (N_9533,N_7620,N_6173);
or U9534 (N_9534,N_7577,N_6783);
nand U9535 (N_9535,N_7143,N_7025);
and U9536 (N_9536,N_7892,N_6971);
xnor U9537 (N_9537,N_7970,N_6705);
or U9538 (N_9538,N_6458,N_7216);
or U9539 (N_9539,N_6533,N_6236);
nand U9540 (N_9540,N_7000,N_7900);
or U9541 (N_9541,N_7472,N_6816);
and U9542 (N_9542,N_6975,N_6007);
nand U9543 (N_9543,N_6536,N_6341);
xnor U9544 (N_9544,N_7797,N_7534);
and U9545 (N_9545,N_7872,N_6108);
nor U9546 (N_9546,N_7730,N_6559);
nor U9547 (N_9547,N_6862,N_6890);
nand U9548 (N_9548,N_7813,N_7848);
nand U9549 (N_9549,N_6707,N_7070);
and U9550 (N_9550,N_7026,N_7059);
nor U9551 (N_9551,N_6954,N_6193);
or U9552 (N_9552,N_7839,N_6774);
and U9553 (N_9553,N_7217,N_6743);
xnor U9554 (N_9554,N_7085,N_7366);
and U9555 (N_9555,N_6531,N_7985);
or U9556 (N_9556,N_7231,N_7154);
and U9557 (N_9557,N_6605,N_6153);
nor U9558 (N_9558,N_6197,N_7233);
or U9559 (N_9559,N_7569,N_7173);
and U9560 (N_9560,N_6351,N_6403);
and U9561 (N_9561,N_6377,N_6559);
nand U9562 (N_9562,N_6926,N_6288);
xor U9563 (N_9563,N_6287,N_7060);
nor U9564 (N_9564,N_6550,N_6336);
xnor U9565 (N_9565,N_6654,N_6229);
nor U9566 (N_9566,N_7341,N_6264);
nor U9567 (N_9567,N_7396,N_6018);
xor U9568 (N_9568,N_7754,N_6019);
or U9569 (N_9569,N_6230,N_7478);
or U9570 (N_9570,N_6496,N_7380);
and U9571 (N_9571,N_6930,N_6689);
and U9572 (N_9572,N_6957,N_6940);
and U9573 (N_9573,N_6883,N_6673);
or U9574 (N_9574,N_7368,N_6532);
nand U9575 (N_9575,N_7378,N_6240);
xnor U9576 (N_9576,N_6250,N_7832);
or U9577 (N_9577,N_6025,N_6143);
or U9578 (N_9578,N_6675,N_7413);
nand U9579 (N_9579,N_6098,N_6092);
and U9580 (N_9580,N_7915,N_7225);
or U9581 (N_9581,N_7630,N_6207);
and U9582 (N_9582,N_7278,N_6431);
and U9583 (N_9583,N_7122,N_6458);
xor U9584 (N_9584,N_6968,N_7881);
xor U9585 (N_9585,N_6670,N_6751);
nand U9586 (N_9586,N_7630,N_7654);
xor U9587 (N_9587,N_7988,N_6796);
and U9588 (N_9588,N_6489,N_7015);
xnor U9589 (N_9589,N_7623,N_7179);
nor U9590 (N_9590,N_6883,N_7882);
or U9591 (N_9591,N_6783,N_6137);
xnor U9592 (N_9592,N_6798,N_6620);
nor U9593 (N_9593,N_6488,N_7160);
and U9594 (N_9594,N_6461,N_7598);
nand U9595 (N_9595,N_6474,N_7305);
xor U9596 (N_9596,N_6823,N_7669);
or U9597 (N_9597,N_6696,N_7025);
nor U9598 (N_9598,N_6837,N_6653);
nand U9599 (N_9599,N_6877,N_6399);
nor U9600 (N_9600,N_7149,N_7655);
nand U9601 (N_9601,N_6778,N_6080);
nor U9602 (N_9602,N_6666,N_6483);
xnor U9603 (N_9603,N_6778,N_6407);
nor U9604 (N_9604,N_7742,N_7410);
xnor U9605 (N_9605,N_6896,N_7025);
nor U9606 (N_9606,N_6898,N_6517);
or U9607 (N_9607,N_6541,N_7645);
xor U9608 (N_9608,N_6464,N_6058);
nor U9609 (N_9609,N_7075,N_7320);
nor U9610 (N_9610,N_6900,N_6288);
xnor U9611 (N_9611,N_6054,N_7258);
xnor U9612 (N_9612,N_6065,N_7998);
or U9613 (N_9613,N_6835,N_6233);
and U9614 (N_9614,N_6668,N_6573);
and U9615 (N_9615,N_6202,N_6843);
xnor U9616 (N_9616,N_6685,N_6305);
xor U9617 (N_9617,N_7117,N_6655);
nor U9618 (N_9618,N_7246,N_7870);
or U9619 (N_9619,N_6346,N_6759);
and U9620 (N_9620,N_7983,N_6033);
or U9621 (N_9621,N_7013,N_6873);
xnor U9622 (N_9622,N_6833,N_6721);
nand U9623 (N_9623,N_7393,N_6527);
nand U9624 (N_9624,N_6452,N_6988);
nor U9625 (N_9625,N_7558,N_7605);
and U9626 (N_9626,N_6060,N_7733);
nand U9627 (N_9627,N_7196,N_6523);
nor U9628 (N_9628,N_6657,N_6714);
nor U9629 (N_9629,N_7214,N_6039);
and U9630 (N_9630,N_7482,N_7180);
xor U9631 (N_9631,N_7428,N_7754);
nand U9632 (N_9632,N_7195,N_7874);
or U9633 (N_9633,N_7969,N_7628);
nor U9634 (N_9634,N_6459,N_7923);
xnor U9635 (N_9635,N_6425,N_7516);
nand U9636 (N_9636,N_6517,N_6238);
xnor U9637 (N_9637,N_6542,N_7564);
xnor U9638 (N_9638,N_7409,N_6045);
nand U9639 (N_9639,N_7790,N_6608);
or U9640 (N_9640,N_7994,N_7860);
and U9641 (N_9641,N_7921,N_7265);
nand U9642 (N_9642,N_6615,N_6909);
xor U9643 (N_9643,N_7576,N_7620);
nand U9644 (N_9644,N_7250,N_7704);
and U9645 (N_9645,N_6312,N_7063);
and U9646 (N_9646,N_7276,N_7157);
nor U9647 (N_9647,N_7689,N_6394);
nand U9648 (N_9648,N_6552,N_7372);
nor U9649 (N_9649,N_6013,N_6191);
or U9650 (N_9650,N_7270,N_7415);
xor U9651 (N_9651,N_6143,N_6687);
xnor U9652 (N_9652,N_7742,N_6851);
xor U9653 (N_9653,N_6240,N_7530);
and U9654 (N_9654,N_7062,N_6381);
nor U9655 (N_9655,N_7041,N_7938);
xor U9656 (N_9656,N_7621,N_6432);
nor U9657 (N_9657,N_6569,N_7866);
nand U9658 (N_9658,N_7806,N_7415);
xnor U9659 (N_9659,N_7626,N_7696);
xnor U9660 (N_9660,N_7956,N_7137);
nor U9661 (N_9661,N_7778,N_6219);
and U9662 (N_9662,N_6758,N_7130);
or U9663 (N_9663,N_6304,N_6260);
nand U9664 (N_9664,N_7367,N_6704);
nor U9665 (N_9665,N_6496,N_6818);
nor U9666 (N_9666,N_7096,N_7435);
nand U9667 (N_9667,N_7286,N_7836);
xnor U9668 (N_9668,N_6961,N_7534);
or U9669 (N_9669,N_7204,N_7426);
or U9670 (N_9670,N_6256,N_7923);
nand U9671 (N_9671,N_7018,N_7236);
or U9672 (N_9672,N_6912,N_6024);
nand U9673 (N_9673,N_7960,N_7704);
nor U9674 (N_9674,N_7015,N_7335);
or U9675 (N_9675,N_6895,N_7265);
or U9676 (N_9676,N_6407,N_7836);
and U9677 (N_9677,N_6762,N_6368);
nor U9678 (N_9678,N_6855,N_6002);
nand U9679 (N_9679,N_7642,N_7315);
nor U9680 (N_9680,N_7784,N_7453);
nor U9681 (N_9681,N_7332,N_7030);
nand U9682 (N_9682,N_6892,N_7911);
nor U9683 (N_9683,N_6231,N_7477);
nor U9684 (N_9684,N_6794,N_7168);
and U9685 (N_9685,N_6810,N_7889);
nand U9686 (N_9686,N_6615,N_7119);
nor U9687 (N_9687,N_6478,N_7963);
nand U9688 (N_9688,N_7326,N_7211);
nor U9689 (N_9689,N_7888,N_6636);
or U9690 (N_9690,N_7766,N_7534);
xor U9691 (N_9691,N_6250,N_6646);
nor U9692 (N_9692,N_7217,N_6586);
nand U9693 (N_9693,N_7481,N_6079);
or U9694 (N_9694,N_6773,N_7702);
nand U9695 (N_9695,N_7212,N_7695);
and U9696 (N_9696,N_7579,N_6791);
or U9697 (N_9697,N_7888,N_6194);
nand U9698 (N_9698,N_7048,N_6983);
and U9699 (N_9699,N_7569,N_7856);
nand U9700 (N_9700,N_6322,N_6353);
and U9701 (N_9701,N_7925,N_7707);
nor U9702 (N_9702,N_7894,N_6979);
or U9703 (N_9703,N_6336,N_7307);
or U9704 (N_9704,N_7671,N_7976);
nand U9705 (N_9705,N_7395,N_6810);
xor U9706 (N_9706,N_6712,N_7813);
nand U9707 (N_9707,N_6818,N_7693);
or U9708 (N_9708,N_7485,N_6385);
nor U9709 (N_9709,N_6557,N_7443);
nor U9710 (N_9710,N_6400,N_7495);
xnor U9711 (N_9711,N_6103,N_7984);
and U9712 (N_9712,N_6376,N_6830);
nand U9713 (N_9713,N_6988,N_6694);
nand U9714 (N_9714,N_7597,N_6324);
xor U9715 (N_9715,N_7959,N_7447);
or U9716 (N_9716,N_6105,N_7456);
xnor U9717 (N_9717,N_6184,N_6577);
nor U9718 (N_9718,N_6377,N_7855);
nor U9719 (N_9719,N_6533,N_6035);
xnor U9720 (N_9720,N_7907,N_6654);
nor U9721 (N_9721,N_6411,N_6030);
and U9722 (N_9722,N_7076,N_7221);
nor U9723 (N_9723,N_6786,N_6207);
or U9724 (N_9724,N_7634,N_6684);
nor U9725 (N_9725,N_6147,N_7357);
and U9726 (N_9726,N_6277,N_7800);
and U9727 (N_9727,N_6601,N_6256);
nand U9728 (N_9728,N_7762,N_7417);
or U9729 (N_9729,N_7161,N_7482);
xor U9730 (N_9730,N_6493,N_6754);
xnor U9731 (N_9731,N_6023,N_6088);
or U9732 (N_9732,N_6838,N_6715);
or U9733 (N_9733,N_6175,N_6937);
and U9734 (N_9734,N_7645,N_6103);
or U9735 (N_9735,N_6843,N_6627);
xor U9736 (N_9736,N_6241,N_7747);
nor U9737 (N_9737,N_7807,N_6957);
nor U9738 (N_9738,N_6252,N_6960);
nand U9739 (N_9739,N_7140,N_7161);
nand U9740 (N_9740,N_7871,N_7757);
or U9741 (N_9741,N_6150,N_6408);
nor U9742 (N_9742,N_7145,N_7710);
or U9743 (N_9743,N_6372,N_6024);
nand U9744 (N_9744,N_6683,N_6042);
or U9745 (N_9745,N_6900,N_7245);
nand U9746 (N_9746,N_7568,N_6226);
nor U9747 (N_9747,N_7455,N_6885);
xor U9748 (N_9748,N_7010,N_6691);
nor U9749 (N_9749,N_6713,N_7204);
and U9750 (N_9750,N_6164,N_6256);
or U9751 (N_9751,N_7371,N_7981);
nor U9752 (N_9752,N_6643,N_6724);
xor U9753 (N_9753,N_7264,N_7610);
nor U9754 (N_9754,N_7737,N_6635);
nor U9755 (N_9755,N_6371,N_6328);
and U9756 (N_9756,N_7690,N_7855);
nor U9757 (N_9757,N_6488,N_7881);
or U9758 (N_9758,N_7626,N_6487);
nor U9759 (N_9759,N_6256,N_7600);
nor U9760 (N_9760,N_6555,N_6931);
or U9761 (N_9761,N_7388,N_6267);
or U9762 (N_9762,N_6152,N_7522);
and U9763 (N_9763,N_6755,N_7332);
xnor U9764 (N_9764,N_7556,N_6947);
and U9765 (N_9765,N_7605,N_7560);
xor U9766 (N_9766,N_7329,N_7815);
and U9767 (N_9767,N_7662,N_6392);
nand U9768 (N_9768,N_7334,N_7100);
and U9769 (N_9769,N_6431,N_6949);
xnor U9770 (N_9770,N_7987,N_7658);
and U9771 (N_9771,N_7046,N_7032);
or U9772 (N_9772,N_7628,N_6265);
nand U9773 (N_9773,N_7364,N_6167);
and U9774 (N_9774,N_6144,N_7070);
xor U9775 (N_9775,N_6757,N_6273);
nor U9776 (N_9776,N_6822,N_7208);
and U9777 (N_9777,N_6189,N_7860);
and U9778 (N_9778,N_6722,N_7019);
and U9779 (N_9779,N_7330,N_6114);
xnor U9780 (N_9780,N_7341,N_6199);
xor U9781 (N_9781,N_7796,N_6517);
xnor U9782 (N_9782,N_7829,N_6981);
nand U9783 (N_9783,N_7241,N_7478);
xnor U9784 (N_9784,N_7315,N_7078);
and U9785 (N_9785,N_7879,N_7583);
xor U9786 (N_9786,N_6930,N_6760);
or U9787 (N_9787,N_7206,N_7312);
or U9788 (N_9788,N_6628,N_6200);
nor U9789 (N_9789,N_6201,N_7827);
or U9790 (N_9790,N_7587,N_7599);
nor U9791 (N_9791,N_6775,N_7635);
and U9792 (N_9792,N_6761,N_7582);
and U9793 (N_9793,N_7838,N_7516);
nor U9794 (N_9794,N_6524,N_6206);
and U9795 (N_9795,N_6520,N_6917);
and U9796 (N_9796,N_6861,N_6591);
nor U9797 (N_9797,N_6938,N_7484);
nand U9798 (N_9798,N_6339,N_7917);
nand U9799 (N_9799,N_6633,N_6315);
and U9800 (N_9800,N_7572,N_6412);
nand U9801 (N_9801,N_7250,N_7692);
and U9802 (N_9802,N_7587,N_6638);
nand U9803 (N_9803,N_7031,N_6051);
and U9804 (N_9804,N_7424,N_7386);
nand U9805 (N_9805,N_7621,N_7989);
and U9806 (N_9806,N_6401,N_7524);
or U9807 (N_9807,N_7020,N_7996);
xor U9808 (N_9808,N_6188,N_7051);
and U9809 (N_9809,N_6426,N_6039);
nand U9810 (N_9810,N_6117,N_6643);
nor U9811 (N_9811,N_6693,N_6890);
and U9812 (N_9812,N_6892,N_7071);
or U9813 (N_9813,N_7735,N_7782);
or U9814 (N_9814,N_6463,N_6725);
or U9815 (N_9815,N_7899,N_7692);
nand U9816 (N_9816,N_7522,N_6138);
xnor U9817 (N_9817,N_7224,N_7449);
xnor U9818 (N_9818,N_6584,N_6713);
nor U9819 (N_9819,N_7669,N_7605);
and U9820 (N_9820,N_6540,N_7396);
nand U9821 (N_9821,N_6309,N_6203);
and U9822 (N_9822,N_6762,N_7027);
xnor U9823 (N_9823,N_7631,N_7195);
or U9824 (N_9824,N_6758,N_6229);
nor U9825 (N_9825,N_6895,N_7778);
nor U9826 (N_9826,N_6068,N_7284);
or U9827 (N_9827,N_6117,N_7791);
nand U9828 (N_9828,N_7581,N_6889);
nor U9829 (N_9829,N_7633,N_6575);
nor U9830 (N_9830,N_7139,N_7966);
or U9831 (N_9831,N_6636,N_6522);
nand U9832 (N_9832,N_6021,N_6763);
xnor U9833 (N_9833,N_7243,N_7590);
or U9834 (N_9834,N_7957,N_6293);
nor U9835 (N_9835,N_7812,N_6676);
xor U9836 (N_9836,N_7792,N_7545);
xor U9837 (N_9837,N_6592,N_7583);
xor U9838 (N_9838,N_6261,N_6414);
xnor U9839 (N_9839,N_6128,N_6386);
nor U9840 (N_9840,N_6942,N_7994);
xnor U9841 (N_9841,N_7179,N_7319);
xor U9842 (N_9842,N_6922,N_6964);
nor U9843 (N_9843,N_7649,N_7717);
nor U9844 (N_9844,N_6028,N_7507);
nand U9845 (N_9845,N_7034,N_6140);
nor U9846 (N_9846,N_6444,N_7573);
xor U9847 (N_9847,N_6474,N_7619);
nand U9848 (N_9848,N_7639,N_6813);
nor U9849 (N_9849,N_6206,N_6716);
and U9850 (N_9850,N_7426,N_7031);
nand U9851 (N_9851,N_7950,N_7492);
nand U9852 (N_9852,N_7813,N_7472);
xor U9853 (N_9853,N_6292,N_7332);
nor U9854 (N_9854,N_7429,N_7147);
or U9855 (N_9855,N_7700,N_7031);
and U9856 (N_9856,N_7167,N_7209);
nand U9857 (N_9857,N_6884,N_6414);
nand U9858 (N_9858,N_6035,N_6369);
xor U9859 (N_9859,N_6118,N_7690);
nand U9860 (N_9860,N_6187,N_7047);
nand U9861 (N_9861,N_6854,N_7543);
and U9862 (N_9862,N_6770,N_6548);
and U9863 (N_9863,N_7776,N_6383);
and U9864 (N_9864,N_7887,N_7001);
nand U9865 (N_9865,N_7503,N_6479);
nand U9866 (N_9866,N_6775,N_7753);
nor U9867 (N_9867,N_7831,N_7457);
or U9868 (N_9868,N_6671,N_6902);
nor U9869 (N_9869,N_7862,N_6042);
nand U9870 (N_9870,N_7039,N_6055);
nor U9871 (N_9871,N_7169,N_7084);
xnor U9872 (N_9872,N_6496,N_7752);
nor U9873 (N_9873,N_7540,N_6870);
xor U9874 (N_9874,N_7737,N_7077);
nor U9875 (N_9875,N_6722,N_7182);
or U9876 (N_9876,N_7843,N_6244);
and U9877 (N_9877,N_6888,N_7113);
xor U9878 (N_9878,N_7204,N_7275);
nor U9879 (N_9879,N_6169,N_6515);
xor U9880 (N_9880,N_7836,N_6845);
nor U9881 (N_9881,N_7547,N_7561);
and U9882 (N_9882,N_7414,N_6969);
and U9883 (N_9883,N_7055,N_6122);
nand U9884 (N_9884,N_7143,N_7426);
nor U9885 (N_9885,N_7173,N_7431);
nor U9886 (N_9886,N_6726,N_6560);
nor U9887 (N_9887,N_6343,N_6454);
or U9888 (N_9888,N_7487,N_7925);
xnor U9889 (N_9889,N_7932,N_6169);
xnor U9890 (N_9890,N_7192,N_7212);
and U9891 (N_9891,N_7637,N_6737);
and U9892 (N_9892,N_6342,N_7141);
or U9893 (N_9893,N_7674,N_7163);
or U9894 (N_9894,N_7732,N_7109);
nand U9895 (N_9895,N_7981,N_6456);
and U9896 (N_9896,N_6690,N_7016);
nand U9897 (N_9897,N_7191,N_6889);
or U9898 (N_9898,N_7841,N_7880);
xor U9899 (N_9899,N_7613,N_7835);
xor U9900 (N_9900,N_6132,N_6645);
or U9901 (N_9901,N_6623,N_6711);
nor U9902 (N_9902,N_7673,N_7224);
nand U9903 (N_9903,N_6359,N_7195);
or U9904 (N_9904,N_6067,N_6897);
and U9905 (N_9905,N_6383,N_7658);
nand U9906 (N_9906,N_7374,N_7587);
and U9907 (N_9907,N_6280,N_7995);
and U9908 (N_9908,N_7236,N_7212);
nand U9909 (N_9909,N_7522,N_6730);
or U9910 (N_9910,N_7960,N_7839);
nor U9911 (N_9911,N_7991,N_6483);
or U9912 (N_9912,N_6561,N_6356);
and U9913 (N_9913,N_7844,N_6134);
or U9914 (N_9914,N_6578,N_7728);
and U9915 (N_9915,N_7978,N_6166);
and U9916 (N_9916,N_6275,N_7886);
nand U9917 (N_9917,N_6565,N_7461);
xnor U9918 (N_9918,N_7779,N_6950);
nor U9919 (N_9919,N_6950,N_6889);
and U9920 (N_9920,N_6182,N_7528);
xnor U9921 (N_9921,N_7058,N_6182);
or U9922 (N_9922,N_7566,N_7523);
and U9923 (N_9923,N_7042,N_6129);
nand U9924 (N_9924,N_7323,N_7100);
nand U9925 (N_9925,N_7133,N_6746);
xor U9926 (N_9926,N_7613,N_7927);
or U9927 (N_9927,N_7448,N_7002);
or U9928 (N_9928,N_6308,N_7197);
and U9929 (N_9929,N_7742,N_6445);
xnor U9930 (N_9930,N_7275,N_7792);
and U9931 (N_9931,N_6625,N_6107);
nor U9932 (N_9932,N_7743,N_6056);
and U9933 (N_9933,N_6109,N_7653);
nand U9934 (N_9934,N_6773,N_6739);
nor U9935 (N_9935,N_7300,N_6851);
xor U9936 (N_9936,N_6669,N_7882);
nand U9937 (N_9937,N_6185,N_7981);
or U9938 (N_9938,N_7598,N_7036);
xnor U9939 (N_9939,N_6935,N_6221);
or U9940 (N_9940,N_6457,N_6128);
and U9941 (N_9941,N_7194,N_6304);
nor U9942 (N_9942,N_7499,N_7445);
nor U9943 (N_9943,N_6129,N_6694);
xnor U9944 (N_9944,N_6954,N_6467);
or U9945 (N_9945,N_7776,N_6340);
xor U9946 (N_9946,N_7101,N_7726);
xor U9947 (N_9947,N_6045,N_7395);
nor U9948 (N_9948,N_6052,N_7131);
xor U9949 (N_9949,N_7480,N_6062);
nand U9950 (N_9950,N_6521,N_7343);
nand U9951 (N_9951,N_6790,N_6063);
or U9952 (N_9952,N_6652,N_7719);
and U9953 (N_9953,N_6927,N_7540);
nand U9954 (N_9954,N_6897,N_7676);
or U9955 (N_9955,N_6667,N_7080);
xor U9956 (N_9956,N_6357,N_6160);
or U9957 (N_9957,N_6676,N_6569);
nor U9958 (N_9958,N_6044,N_7403);
or U9959 (N_9959,N_6740,N_7717);
and U9960 (N_9960,N_6082,N_7772);
xnor U9961 (N_9961,N_6826,N_7732);
or U9962 (N_9962,N_6740,N_6144);
or U9963 (N_9963,N_6706,N_6551);
nor U9964 (N_9964,N_7102,N_6497);
nor U9965 (N_9965,N_7451,N_6695);
nor U9966 (N_9966,N_6923,N_7327);
and U9967 (N_9967,N_6776,N_7397);
nor U9968 (N_9968,N_6550,N_6972);
or U9969 (N_9969,N_7144,N_6951);
xor U9970 (N_9970,N_7952,N_6754);
nand U9971 (N_9971,N_6992,N_7474);
nor U9972 (N_9972,N_7169,N_7290);
xnor U9973 (N_9973,N_6026,N_7277);
and U9974 (N_9974,N_7987,N_6119);
or U9975 (N_9975,N_7392,N_6421);
nand U9976 (N_9976,N_7342,N_6496);
or U9977 (N_9977,N_6787,N_7807);
nand U9978 (N_9978,N_6485,N_6742);
xor U9979 (N_9979,N_7326,N_7547);
nor U9980 (N_9980,N_7315,N_6312);
nand U9981 (N_9981,N_6850,N_7201);
or U9982 (N_9982,N_7314,N_6669);
and U9983 (N_9983,N_6562,N_6748);
xor U9984 (N_9984,N_7982,N_7161);
and U9985 (N_9985,N_6599,N_7776);
nor U9986 (N_9986,N_6051,N_6692);
nor U9987 (N_9987,N_6807,N_7593);
xnor U9988 (N_9988,N_7248,N_6837);
xor U9989 (N_9989,N_7277,N_7663);
xnor U9990 (N_9990,N_6595,N_7684);
nand U9991 (N_9991,N_6013,N_7505);
nor U9992 (N_9992,N_6959,N_6679);
and U9993 (N_9993,N_6658,N_7627);
and U9994 (N_9994,N_6969,N_6599);
xor U9995 (N_9995,N_7040,N_6017);
xor U9996 (N_9996,N_6235,N_7921);
or U9997 (N_9997,N_6625,N_7272);
nand U9998 (N_9998,N_7066,N_6003);
and U9999 (N_9999,N_6026,N_6092);
nand U10000 (N_10000,N_8407,N_9463);
nand U10001 (N_10001,N_9763,N_8959);
or U10002 (N_10002,N_8426,N_9148);
and U10003 (N_10003,N_8304,N_9978);
and U10004 (N_10004,N_9854,N_8374);
nor U10005 (N_10005,N_9368,N_8370);
nand U10006 (N_10006,N_9813,N_9259);
nor U10007 (N_10007,N_8845,N_9779);
xnor U10008 (N_10008,N_9161,N_9401);
or U10009 (N_10009,N_9611,N_9270);
nand U10010 (N_10010,N_8296,N_8583);
and U10011 (N_10011,N_9659,N_9150);
xnor U10012 (N_10012,N_8377,N_8473);
and U10013 (N_10013,N_8770,N_9921);
xor U10014 (N_10014,N_9929,N_9363);
xnor U10015 (N_10015,N_9308,N_9636);
nor U10016 (N_10016,N_8405,N_9907);
or U10017 (N_10017,N_8223,N_8855);
and U10018 (N_10018,N_8506,N_9496);
or U10019 (N_10019,N_9880,N_8432);
xor U10020 (N_10020,N_8086,N_8019);
and U10021 (N_10021,N_9169,N_9371);
or U10022 (N_10022,N_8962,N_9361);
or U10023 (N_10023,N_8725,N_9153);
nor U10024 (N_10024,N_9803,N_9831);
nand U10025 (N_10025,N_8309,N_9777);
and U10026 (N_10026,N_8616,N_9588);
nand U10027 (N_10027,N_8918,N_8105);
nor U10028 (N_10028,N_8665,N_8668);
or U10029 (N_10029,N_8498,N_9589);
or U10030 (N_10030,N_8993,N_9677);
xnor U10031 (N_10031,N_8122,N_9132);
and U10032 (N_10032,N_8253,N_8630);
nor U10033 (N_10033,N_8631,N_9290);
xnor U10034 (N_10034,N_8521,N_8948);
or U10035 (N_10035,N_8698,N_8767);
nor U10036 (N_10036,N_9489,N_8600);
nand U10037 (N_10037,N_8230,N_8531);
and U10038 (N_10038,N_8522,N_8797);
and U10039 (N_10039,N_8452,N_8284);
nor U10040 (N_10040,N_9580,N_8115);
nand U10041 (N_10041,N_8205,N_9322);
or U10042 (N_10042,N_8999,N_8656);
nand U10043 (N_10043,N_8158,N_8933);
nand U10044 (N_10044,N_9772,N_8879);
or U10045 (N_10045,N_9435,N_9151);
nand U10046 (N_10046,N_9491,N_8662);
nor U10047 (N_10047,N_8641,N_8977);
and U10048 (N_10048,N_9296,N_9941);
or U10049 (N_10049,N_8460,N_8132);
nand U10050 (N_10050,N_8661,N_8308);
and U10051 (N_10051,N_9547,N_9556);
nand U10052 (N_10052,N_8741,N_9681);
nor U10053 (N_10053,N_9657,N_9615);
xor U10054 (N_10054,N_9874,N_9468);
xnor U10055 (N_10055,N_8495,N_9952);
nand U10056 (N_10056,N_8821,N_8333);
xnor U10057 (N_10057,N_9718,N_9538);
or U10058 (N_10058,N_9914,N_9469);
nand U10059 (N_10059,N_8776,N_9833);
or U10060 (N_10060,N_8275,N_9273);
nand U10061 (N_10061,N_8591,N_9931);
nor U10062 (N_10062,N_9386,N_8929);
nor U10063 (N_10063,N_9550,N_9184);
nor U10064 (N_10064,N_9356,N_8049);
or U10065 (N_10065,N_8010,N_9258);
or U10066 (N_10066,N_8120,N_8366);
or U10067 (N_10067,N_8623,N_8087);
nor U10068 (N_10068,N_9506,N_9108);
nand U10069 (N_10069,N_8260,N_8097);
nor U10070 (N_10070,N_8624,N_9725);
nor U10071 (N_10071,N_8898,N_8337);
xor U10072 (N_10072,N_9440,N_8839);
and U10073 (N_10073,N_8637,N_9924);
nand U10074 (N_10074,N_8615,N_9284);
and U10075 (N_10075,N_8173,N_9050);
xor U10076 (N_10076,N_9853,N_9080);
nor U10077 (N_10077,N_9011,N_9487);
nand U10078 (N_10078,N_8981,N_8055);
nor U10079 (N_10079,N_9965,N_9970);
nor U10080 (N_10080,N_8729,N_9243);
nand U10081 (N_10081,N_8081,N_9790);
xnor U10082 (N_10082,N_8576,N_8501);
or U10083 (N_10083,N_8082,N_9445);
xnor U10084 (N_10084,N_8970,N_9774);
and U10085 (N_10085,N_9093,N_9382);
nand U10086 (N_10086,N_9137,N_8372);
xnor U10087 (N_10087,N_8730,N_9622);
nand U10088 (N_10088,N_9141,N_8266);
and U10089 (N_10089,N_9343,N_8660);
nand U10090 (N_10090,N_9688,N_9647);
nor U10091 (N_10091,N_9254,N_9497);
nand U10092 (N_10092,N_9005,N_8563);
nor U10093 (N_10093,N_8357,N_8453);
nand U10094 (N_10094,N_8575,N_9094);
xor U10095 (N_10095,N_9825,N_8772);
xor U10096 (N_10096,N_8713,N_9748);
and U10097 (N_10097,N_9620,N_9616);
or U10098 (N_10098,N_9626,N_8386);
and U10099 (N_10099,N_9376,N_8995);
nor U10100 (N_10100,N_8645,N_9239);
nor U10101 (N_10101,N_8565,N_9134);
nor U10102 (N_10102,N_8611,N_8709);
or U10103 (N_10103,N_8718,N_8472);
and U10104 (N_10104,N_8973,N_9302);
nor U10105 (N_10105,N_8860,N_8315);
or U10106 (N_10106,N_9052,N_9808);
or U10107 (N_10107,N_9089,N_9895);
or U10108 (N_10108,N_8449,N_8066);
or U10109 (N_10109,N_9127,N_9158);
and U10110 (N_10110,N_8877,N_9063);
and U10111 (N_10111,N_8510,N_9384);
and U10112 (N_10112,N_8540,N_8701);
or U10113 (N_10113,N_9707,N_8146);
or U10114 (N_10114,N_8383,N_9083);
nor U10115 (N_10115,N_8674,N_8279);
xor U10116 (N_10116,N_9960,N_9160);
nor U10117 (N_10117,N_8378,N_9652);
or U10118 (N_10118,N_8423,N_9848);
nor U10119 (N_10119,N_9564,N_9680);
and U10120 (N_10120,N_8569,N_8924);
nand U10121 (N_10121,N_9872,N_8737);
xnor U10122 (N_10122,N_8803,N_8037);
and U10123 (N_10123,N_8069,N_8939);
nand U10124 (N_10124,N_9128,N_8829);
and U10125 (N_10125,N_9663,N_9199);
nand U10126 (N_10126,N_9757,N_9003);
nand U10127 (N_10127,N_8654,N_9282);
nor U10128 (N_10128,N_8567,N_9219);
or U10129 (N_10129,N_9536,N_8707);
xnor U10130 (N_10130,N_8710,N_8912);
nand U10131 (N_10131,N_9608,N_8966);
or U10132 (N_10132,N_9344,N_9812);
nand U10133 (N_10133,N_9403,N_8195);
nand U10134 (N_10134,N_8610,N_9909);
nor U10135 (N_10135,N_9216,N_9561);
or U10136 (N_10136,N_8858,N_8189);
nand U10137 (N_10137,N_9665,N_8721);
and U10138 (N_10138,N_8893,N_9274);
and U10139 (N_10139,N_8834,N_8258);
xnor U10140 (N_10140,N_9495,N_8218);
and U10141 (N_10141,N_8448,N_8468);
xor U10142 (N_10142,N_8492,N_8633);
nor U10143 (N_10143,N_9662,N_8853);
xor U10144 (N_10144,N_8989,N_8910);
nand U10145 (N_10145,N_9694,N_9037);
nand U10146 (N_10146,N_8997,N_9028);
and U10147 (N_10147,N_9143,N_9939);
and U10148 (N_10148,N_8926,N_8067);
and U10149 (N_10149,N_8722,N_9181);
nor U10150 (N_10150,N_8290,N_8738);
nor U10151 (N_10151,N_8881,N_8325);
nor U10152 (N_10152,N_9845,N_8482);
xnor U10153 (N_10153,N_8469,N_8620);
nor U10154 (N_10154,N_9464,N_9780);
nand U10155 (N_10155,N_8850,N_8470);
or U10156 (N_10156,N_9072,N_8270);
nor U10157 (N_10157,N_8208,N_9533);
nand U10158 (N_10158,N_9627,N_9773);
nand U10159 (N_10159,N_9612,N_8647);
and U10160 (N_10160,N_8231,N_9634);
or U10161 (N_10161,N_9610,N_8140);
xor U10162 (N_10162,N_8534,N_8344);
or U10163 (N_10163,N_9568,N_8638);
or U10164 (N_10164,N_9856,N_8272);
or U10165 (N_10165,N_9458,N_8245);
nand U10166 (N_10166,N_9508,N_9018);
nor U10167 (N_10167,N_8161,N_9316);
or U10168 (N_10168,N_9949,N_8382);
or U10169 (N_10169,N_9815,N_8593);
or U10170 (N_10170,N_9044,N_8006);
and U10171 (N_10171,N_9753,N_8694);
and U10172 (N_10172,N_9022,N_9360);
nor U10173 (N_10173,N_8237,N_9849);
nand U10174 (N_10174,N_9117,N_8833);
and U10175 (N_10175,N_8676,N_9473);
nor U10176 (N_10176,N_8794,N_8091);
xnor U10177 (N_10177,N_9041,N_8009);
and U10178 (N_10178,N_8868,N_9521);
and U10179 (N_10179,N_9514,N_9999);
xor U10180 (N_10180,N_8792,N_9175);
nand U10181 (N_10181,N_8040,N_9706);
and U10182 (N_10182,N_8972,N_9786);
nand U10183 (N_10183,N_9074,N_9043);
or U10184 (N_10184,N_9498,N_9756);
and U10185 (N_10185,N_9852,N_9947);
nand U10186 (N_10186,N_9244,N_8490);
or U10187 (N_10187,N_9472,N_8273);
and U10188 (N_10188,N_9743,N_9250);
or U10189 (N_10189,N_9972,N_8340);
nor U10190 (N_10190,N_8675,N_9606);
and U10191 (N_10191,N_8542,N_9925);
and U10192 (N_10192,N_9233,N_8288);
nand U10193 (N_10193,N_9112,N_9144);
and U10194 (N_10194,N_9251,N_8181);
nand U10195 (N_10195,N_8935,N_8271);
nor U10196 (N_10196,N_8937,N_8311);
or U10197 (N_10197,N_9574,N_9915);
nor U10198 (N_10198,N_8658,N_8994);
or U10199 (N_10199,N_9271,N_9715);
nor U10200 (N_10200,N_8119,N_9846);
xnor U10201 (N_10201,N_9213,N_8026);
or U10202 (N_10202,N_9370,N_9884);
nor U10203 (N_10203,N_8815,N_8047);
and U10204 (N_10204,N_9323,N_9224);
nand U10205 (N_10205,N_9422,N_9217);
nor U10206 (N_10206,N_8265,N_9090);
nor U10207 (N_10207,N_9406,N_9327);
xor U10208 (N_10208,N_8058,N_8920);
and U10209 (N_10209,N_9099,N_8338);
nor U10210 (N_10210,N_9412,N_8439);
xnor U10211 (N_10211,N_9352,N_9512);
xnor U10212 (N_10212,N_8095,N_9367);
and U10213 (N_10213,N_8945,N_9670);
nor U10214 (N_10214,N_8419,N_8692);
nand U10215 (N_10215,N_8403,N_8018);
xor U10216 (N_10216,N_9045,N_9122);
and U10217 (N_10217,N_8734,N_9317);
and U10218 (N_10218,N_9110,N_8391);
nor U10219 (N_10219,N_9300,N_8336);
nand U10220 (N_10220,N_8030,N_9246);
xor U10221 (N_10221,N_9193,N_8950);
nor U10222 (N_10222,N_8528,N_9858);
xnor U10223 (N_10223,N_9085,N_9792);
nor U10224 (N_10224,N_9565,N_9782);
xnor U10225 (N_10225,N_8762,N_8418);
xor U10226 (N_10226,N_9971,N_8594);
and U10227 (N_10227,N_8609,N_8346);
nand U10228 (N_10228,N_8437,N_9188);
xor U10229 (N_10229,N_8795,N_8201);
nor U10230 (N_10230,N_8785,N_8033);
and U10231 (N_10231,N_8278,N_8800);
nand U10232 (N_10232,N_8276,N_8389);
and U10233 (N_10233,N_8180,N_8988);
and U10234 (N_10234,N_8072,N_9225);
xnor U10235 (N_10235,N_9378,N_8628);
xnor U10236 (N_10236,N_9346,N_8282);
and U10237 (N_10237,N_9525,N_8960);
nor U10238 (N_10238,N_8001,N_8663);
or U10239 (N_10239,N_8753,N_9056);
and U10240 (N_10240,N_9645,N_8043);
or U10241 (N_10241,N_9220,N_8552);
nor U10242 (N_10242,N_9866,N_9211);
and U10243 (N_10243,N_9221,N_8683);
nand U10244 (N_10244,N_8487,N_8404);
xor U10245 (N_10245,N_9791,N_9030);
xnor U10246 (N_10246,N_8252,N_9278);
or U10247 (N_10247,N_8297,N_9338);
nor U10248 (N_10248,N_8783,N_8758);
and U10249 (N_10249,N_8537,N_9180);
or U10250 (N_10250,N_9391,N_9326);
nand U10251 (N_10251,N_9119,N_8664);
and U10252 (N_10252,N_8232,N_8518);
or U10253 (N_10253,N_8690,N_9457);
xnor U10254 (N_10254,N_9399,N_8556);
and U10255 (N_10255,N_9519,N_9493);
xor U10256 (N_10256,N_8728,N_8618);
nand U10257 (N_10257,N_8882,N_8209);
nand U10258 (N_10258,N_8817,N_8176);
nor U10259 (N_10259,N_8614,N_9172);
xor U10260 (N_10260,N_9750,N_9329);
and U10261 (N_10261,N_9294,N_9903);
xor U10262 (N_10262,N_9269,N_8923);
nand U10263 (N_10263,N_8318,N_8570);
or U10264 (N_10264,N_8568,N_9276);
and U10265 (N_10265,N_9967,N_8847);
nor U10266 (N_10266,N_8027,N_9920);
nand U10267 (N_10267,N_9751,N_8184);
or U10268 (N_10268,N_8394,N_8375);
nand U10269 (N_10269,N_8339,N_9766);
nor U10270 (N_10270,N_9804,N_8213);
nor U10271 (N_10271,N_9655,N_8678);
nand U10272 (N_10272,N_9686,N_9484);
xor U10273 (N_10273,N_9097,N_9770);
or U10274 (N_10274,N_8233,N_8524);
nor U10275 (N_10275,N_9827,N_9631);
nand U10276 (N_10276,N_8739,N_8379);
nor U10277 (N_10277,N_8077,N_9460);
nor U10278 (N_10278,N_9973,N_9073);
or U10279 (N_10279,N_9047,N_8306);
nor U10280 (N_10280,N_9765,N_8327);
or U10281 (N_10281,N_9524,N_9544);
or U10282 (N_10282,N_8113,N_8254);
and U10283 (N_10283,N_8416,N_9196);
and U10284 (N_10284,N_8836,N_9732);
or U10285 (N_10285,N_8480,N_9877);
and U10286 (N_10286,N_9078,N_8462);
nor U10287 (N_10287,N_8969,N_9828);
xor U10288 (N_10288,N_8194,N_9761);
or U10289 (N_10289,N_8559,N_8842);
and U10290 (N_10290,N_9930,N_8951);
nor U10291 (N_10291,N_9335,N_9345);
or U10292 (N_10292,N_9964,N_8869);
or U10293 (N_10293,N_8399,N_9426);
xor U10294 (N_10294,N_9836,N_9191);
nor U10295 (N_10295,N_9850,N_8771);
or U10296 (N_10296,N_9795,N_9847);
xnor U10297 (N_10297,N_9746,N_9229);
nor U10298 (N_10298,N_8479,N_9842);
nand U10299 (N_10299,N_8151,N_9424);
and U10300 (N_10300,N_9505,N_9515);
or U10301 (N_10301,N_8578,N_8560);
or U10302 (N_10302,N_9559,N_9373);
and U10303 (N_10303,N_9374,N_9528);
nor U10304 (N_10304,N_9883,N_9265);
nand U10305 (N_10305,N_9310,N_9025);
nand U10306 (N_10306,N_8174,N_8813);
xnor U10307 (N_10307,N_9891,N_9860);
nand U10308 (N_10308,N_8515,N_8451);
xor U10309 (N_10309,N_9992,N_9466);
xnor U10310 (N_10310,N_8886,N_9987);
or U10311 (N_10311,N_9502,N_8247);
nand U10312 (N_10312,N_8261,N_8790);
and U10313 (N_10313,N_8241,N_8466);
xor U10314 (N_10314,N_8427,N_9055);
xnor U10315 (N_10315,N_8581,N_9332);
and U10316 (N_10316,N_9724,N_8435);
xor U10317 (N_10317,N_8597,N_8070);
or U10318 (N_10318,N_9560,N_9837);
nor U10319 (N_10319,N_8588,N_8411);
or U10320 (N_10320,N_8085,N_9876);
and U10321 (N_10321,N_9597,N_9867);
and U10322 (N_10322,N_8301,N_8878);
xor U10323 (N_10323,N_8234,N_9079);
xnor U10324 (N_10324,N_9318,N_9297);
and U10325 (N_10325,N_8827,N_8635);
nand U10326 (N_10326,N_9535,N_8526);
and U10327 (N_10327,N_9618,N_8643);
and U10328 (N_10328,N_8554,N_8687);
nor U10329 (N_10329,N_8443,N_8903);
and U10330 (N_10330,N_8135,N_8511);
and U10331 (N_10331,N_8857,N_8704);
or U10332 (N_10332,N_9632,N_8627);
or U10333 (N_10333,N_8250,N_9054);
and U10334 (N_10334,N_9709,N_8814);
xor U10335 (N_10335,N_8916,N_8777);
nor U10336 (N_10336,N_9811,N_8291);
nand U10337 (N_10337,N_9393,N_8329);
nor U10338 (N_10338,N_8582,N_9307);
nand U10339 (N_10339,N_8513,N_9537);
or U10340 (N_10340,N_9938,N_9552);
or U10341 (N_10341,N_9764,N_9584);
nor U10342 (N_10342,N_9542,N_9567);
and U10343 (N_10343,N_8185,N_9288);
nor U10344 (N_10344,N_9526,N_8793);
xnor U10345 (N_10345,N_9592,N_8984);
or U10346 (N_10346,N_8360,N_8889);
or U10347 (N_10347,N_8280,N_8242);
or U10348 (N_10348,N_9948,N_9065);
or U10349 (N_10349,N_9985,N_9660);
xor U10350 (N_10350,N_9576,N_9113);
nand U10351 (N_10351,N_9260,N_8596);
xor U10352 (N_10352,N_9864,N_8310);
nand U10353 (N_10353,N_8170,N_8356);
and U10354 (N_10354,N_8429,N_8369);
xnor U10355 (N_10355,N_9404,N_8128);
nand U10356 (N_10356,N_9824,N_9979);
nand U10357 (N_10357,N_9299,N_9805);
nand U10358 (N_10358,N_9479,N_9477);
or U10359 (N_10359,N_9628,N_8961);
nor U10360 (N_10360,N_9135,N_8430);
nor U10361 (N_10361,N_8157,N_8021);
nor U10362 (N_10362,N_8186,N_8034);
xnor U10363 (N_10363,N_9263,N_9014);
nand U10364 (N_10364,N_8564,N_8222);
and U10365 (N_10365,N_9111,N_8155);
nor U10366 (N_10366,N_8450,N_9951);
or U10367 (N_10367,N_8684,N_9165);
nand U10368 (N_10368,N_9630,N_8905);
or U10369 (N_10369,N_9607,N_9136);
nand U10370 (N_10370,N_8198,N_9103);
xnor U10371 (N_10371,N_9739,N_9983);
nand U10372 (N_10372,N_9204,N_8975);
or U10373 (N_10373,N_9336,N_9142);
or U10374 (N_10374,N_8782,N_9449);
nand U10375 (N_10375,N_8523,N_8384);
nand U10376 (N_10376,N_9741,N_9486);
xnor U10377 (N_10377,N_9637,N_8688);
and U10378 (N_10378,N_8530,N_9434);
and U10379 (N_10379,N_8459,N_9400);
nor U10380 (N_10380,N_9916,N_9405);
nand U10381 (N_10381,N_9747,N_9591);
and U10382 (N_10382,N_8870,N_9784);
nor U10383 (N_10383,N_8517,N_8715);
or U10384 (N_10384,N_9185,N_9086);
or U10385 (N_10385,N_8805,N_8062);
and U10386 (N_10386,N_9830,N_8786);
nor U10387 (N_10387,N_8917,N_8612);
nor U10388 (N_10388,N_8685,N_9075);
or U10389 (N_10389,N_8371,N_9430);
nor U10390 (N_10390,N_8228,N_8111);
nor U10391 (N_10391,N_8401,N_8166);
or U10392 (N_10392,N_8285,N_8798);
xnor U10393 (N_10393,N_8976,N_9116);
nand U10394 (N_10394,N_8352,N_8073);
nor U10395 (N_10395,N_8235,N_8619);
xor U10396 (N_10396,N_8368,N_9775);
nor U10397 (N_10397,N_9762,N_9928);
nor U10398 (N_10398,N_8035,N_8532);
xor U10399 (N_10399,N_8063,N_9015);
nor U10400 (N_10400,N_9459,N_9549);
xor U10401 (N_10401,N_8395,N_8670);
nand U10402 (N_10402,N_9887,N_9974);
nand U10403 (N_10403,N_8896,N_8749);
nand U10404 (N_10404,N_9602,N_9010);
or U10405 (N_10405,N_8673,N_9726);
xnor U10406 (N_10406,N_8884,N_8003);
nor U10407 (N_10407,N_8461,N_8101);
or U10408 (N_10408,N_9397,N_8548);
nand U10409 (N_10409,N_8457,N_8529);
nor U10410 (N_10410,N_9878,N_8367);
xnor U10411 (N_10411,N_8109,N_8312);
nor U10412 (N_10412,N_9901,N_9354);
nand U10413 (N_10413,N_9742,N_9413);
or U10414 (N_10414,N_9333,N_8714);
nand U10415 (N_10415,N_9593,N_8483);
nand U10416 (N_10416,N_9034,N_8053);
nor U10417 (N_10417,N_8023,N_8179);
xnor U10418 (N_10418,N_9328,N_8139);
xnor U10419 (N_10419,N_9410,N_8544);
nand U10420 (N_10420,N_9183,N_9714);
and U10421 (N_10421,N_9996,N_9863);
nor U10422 (N_10422,N_8986,N_8032);
nand U10423 (N_10423,N_9668,N_8212);
nand U10424 (N_10424,N_9409,N_9155);
xnor U10425 (N_10425,N_8543,N_9717);
and U10426 (N_10426,N_9759,N_8440);
nor U10427 (N_10427,N_9671,N_8657);
xnor U10428 (N_10428,N_9927,N_8491);
or U10429 (N_10429,N_9087,N_9981);
and U10430 (N_10430,N_8446,N_8240);
or U10431 (N_10431,N_8425,N_8351);
and U10432 (N_10432,N_9039,N_9699);
xnor U10433 (N_10433,N_8550,N_9242);
and U10434 (N_10434,N_8331,N_9095);
and U10435 (N_10435,N_9334,N_8041);
nor U10436 (N_10436,N_9625,N_9088);
nand U10437 (N_10437,N_9076,N_8696);
and U10438 (N_10438,N_9214,N_8160);
and U10439 (N_10439,N_8020,N_8823);
and U10440 (N_10440,N_8693,N_9955);
and U10441 (N_10441,N_9685,N_8595);
or U10442 (N_10442,N_8355,N_8298);
nand U10443 (N_10443,N_9913,N_9289);
or U10444 (N_10444,N_9053,N_8586);
nor U10445 (N_10445,N_8703,N_9942);
nor U10446 (N_10446,N_9383,N_9541);
xor U10447 (N_10447,N_8178,N_8484);
xnor U10448 (N_10448,N_9461,N_9737);
nor U10449 (N_10449,N_8096,N_8551);
nand U10450 (N_10450,N_8971,N_9059);
and U10451 (N_10451,N_9474,N_8188);
xor U10452 (N_10452,N_8334,N_9963);
xor U10453 (N_10453,N_8804,N_9862);
xor U10454 (N_10454,N_8478,N_9871);
nand U10455 (N_10455,N_9557,N_9977);
xor U10456 (N_10456,N_8732,N_9994);
xnor U10457 (N_10457,N_9342,N_8458);
nand U10458 (N_10458,N_9569,N_8150);
xor U10459 (N_10459,N_8979,N_9446);
and U10460 (N_10460,N_9868,N_9562);
or U10461 (N_10461,N_9480,N_9279);
nand U10462 (N_10462,N_8810,N_8863);
or U10463 (N_10463,N_8811,N_9358);
nand U10464 (N_10464,N_8302,N_9396);
xnor U10465 (N_10465,N_9917,N_9692);
or U10466 (N_10466,N_9070,N_9411);
or U10467 (N_10467,N_9377,N_9922);
xor U10468 (N_10468,N_9869,N_9285);
and U10469 (N_10469,N_8434,N_8016);
nand U10470 (N_10470,N_8689,N_8604);
and U10471 (N_10471,N_9684,N_8779);
xor U10472 (N_10472,N_9234,N_8267);
or U10473 (N_10473,N_8536,N_9106);
and U10474 (N_10474,N_8801,N_9171);
nor U10475 (N_10475,N_9066,N_9966);
nor U10476 (N_10476,N_9036,N_8126);
nand U10477 (N_10477,N_8078,N_9101);
nand U10478 (N_10478,N_9031,N_9320);
nand U10479 (N_10479,N_8885,N_9800);
xnor U10480 (N_10480,N_9157,N_9232);
nor U10481 (N_10481,N_8071,N_8013);
and U10482 (N_10482,N_8717,N_9207);
or U10483 (N_10483,N_9545,N_9247);
nand U10484 (N_10484,N_8719,N_9531);
and U10485 (N_10485,N_8930,N_8328);
and U10486 (N_10486,N_8044,N_9267);
nand U10487 (N_10487,N_9357,N_8682);
nor U10488 (N_10488,N_8765,N_9355);
xor U10489 (N_10489,N_8625,N_8332);
and U10490 (N_10490,N_8843,N_9933);
and U10491 (N_10491,N_8224,N_9482);
xnor U10492 (N_10492,N_8104,N_9266);
nor U10493 (N_10493,N_8752,N_9313);
nand U10494 (N_10494,N_9991,N_9209);
xnor U10495 (N_10495,N_8477,N_9575);
or U10496 (N_10496,N_9534,N_8909);
and U10497 (N_10497,N_8216,N_9324);
nand U10498 (N_10498,N_9281,N_8154);
nand U10499 (N_10499,N_9203,N_8946);
xnor U10500 (N_10500,N_9305,N_9566);
xnor U10501 (N_10501,N_8538,N_8629);
or U10502 (N_10502,N_9154,N_8778);
nor U10503 (N_10503,N_8187,N_8299);
nor U10504 (N_10504,N_9583,N_8726);
or U10505 (N_10505,N_9236,N_8464);
or U10506 (N_10506,N_9231,N_8901);
nor U10507 (N_10507,N_9644,N_9176);
nand U10508 (N_10508,N_9619,N_8156);
nor U10509 (N_10509,N_9801,N_8215);
and U10510 (N_10510,N_9295,N_8121);
nor U10511 (N_10511,N_8206,N_9820);
and U10512 (N_10512,N_8130,N_9441);
and U10513 (N_10513,N_8114,N_9235);
nand U10514 (N_10514,N_9767,N_9168);
or U10515 (N_10515,N_8042,N_8784);
and U10516 (N_10516,N_8447,N_8396);
nand U10517 (N_10517,N_8052,N_8880);
nor U10518 (N_10518,N_8390,N_9904);
xnor U10519 (N_10519,N_8431,N_9926);
nor U10520 (N_10520,N_8118,N_8846);
and U10521 (N_10521,N_8277,N_9421);
nand U10522 (N_10522,N_9245,N_9339);
nor U10523 (N_10523,N_8193,N_8031);
or U10524 (N_10524,N_8789,N_8539);
nor U10525 (N_10525,N_9009,N_8519);
xnor U10526 (N_10526,N_9959,N_8321);
xor U10527 (N_10527,N_8764,N_8968);
and U10528 (N_10528,N_9023,N_9797);
and U10529 (N_10529,N_8816,N_8392);
and U10530 (N_10530,N_9776,N_9013);
or U10531 (N_10531,N_8475,N_9624);
nor U10532 (N_10532,N_8949,N_8171);
xnor U10533 (N_10533,N_8942,N_8955);
nor U10534 (N_10534,N_9582,N_9590);
xor U10535 (N_10535,N_8134,N_8486);
and U10536 (N_10536,N_8133,N_8402);
or U10537 (N_10537,N_8421,N_9268);
xnor U10538 (N_10538,N_8899,N_9198);
and U10539 (N_10539,N_8292,N_9178);
nand U10540 (N_10540,N_8471,N_9802);
and U10541 (N_10541,N_9192,N_9851);
nor U10542 (N_10542,N_8561,N_9008);
or U10543 (N_10543,N_8756,N_8711);
and U10544 (N_10544,N_9120,N_9572);
xnor U10545 (N_10545,N_9130,N_8246);
and U10546 (N_10546,N_8196,N_8617);
nand U10547 (N_10547,N_8967,N_9595);
nand U10548 (N_10548,N_8388,N_8463);
or U10549 (N_10549,N_9398,N_8385);
xnor U10550 (N_10550,N_9040,N_9527);
nand U10551 (N_10551,N_9810,N_8603);
nand U10552 (N_10552,N_8553,N_9696);
nor U10553 (N_10553,N_9897,N_9123);
xnor U10554 (N_10554,N_9483,N_8705);
xor U10555 (N_10555,N_9799,N_9453);
or U10556 (N_10556,N_8566,N_9190);
nand U10557 (N_10557,N_9359,N_8520);
and U10558 (N_10558,N_9348,N_9470);
nor U10559 (N_10559,N_8965,N_9456);
or U10560 (N_10560,N_9443,N_9280);
or U10561 (N_10561,N_9661,N_8397);
xnor U10562 (N_10562,N_9744,N_9911);
nor U10563 (N_10563,N_8757,N_8621);
nor U10564 (N_10564,N_9675,N_8607);
nand U10565 (N_10565,N_8788,N_8436);
nor U10566 (N_10566,N_8642,N_8225);
nor U10567 (N_10567,N_9029,N_9511);
nand U10568 (N_10568,N_9771,N_8514);
and U10569 (N_10569,N_9730,N_9923);
nand U10570 (N_10570,N_9425,N_9980);
or U10571 (N_10571,N_8787,N_8326);
xnor U10572 (N_10572,N_8851,N_8874);
xnor U10573 (N_10573,N_8956,N_9609);
or U10574 (N_10574,N_9641,N_9530);
nor U10575 (N_10575,N_9740,N_9369);
nand U10576 (N_10576,N_9691,N_9814);
nand U10577 (N_10577,N_9096,N_9201);
nand U10578 (N_10578,N_8902,N_8985);
nand U10579 (N_10579,N_8313,N_8287);
xnor U10580 (N_10580,N_8283,N_8364);
xor U10581 (N_10581,N_9304,N_9760);
nand U10582 (N_10582,N_8735,N_9754);
nand U10583 (N_10583,N_8613,N_9447);
or U10584 (N_10584,N_8598,N_8653);
nor U10585 (N_10585,N_8289,N_9807);
nand U10586 (N_10586,N_8512,N_8183);
nor U10587 (N_10587,N_8263,N_9380);
nor U10588 (N_10588,N_9021,N_8084);
or U10589 (N_10589,N_9529,N_9614);
and U10590 (N_10590,N_9450,N_8695);
xnor U10591 (N_10591,N_8830,N_8866);
nand U10592 (N_10592,N_8017,N_9001);
nand U10593 (N_10593,N_9573,N_8921);
nand U10594 (N_10594,N_9778,N_9414);
nand U10595 (N_10595,N_8697,N_9613);
xnor U10596 (N_10596,N_9653,N_9841);
nor U10597 (N_10597,N_9210,N_8089);
or U10598 (N_10598,N_8555,N_8589);
xor U10599 (N_10599,N_8137,N_8632);
nand U10600 (N_10600,N_8932,N_9131);
nand U10601 (N_10601,N_8864,N_8143);
xor U10602 (N_10602,N_9432,N_8796);
or U10603 (N_10603,N_8648,N_9603);
nand U10604 (N_10604,N_8415,N_9989);
xor U10605 (N_10605,N_8541,N_8507);
nor U10606 (N_10606,N_8493,N_9272);
xor U10607 (N_10607,N_9716,N_9164);
nand U10608 (N_10608,N_8269,N_9712);
or U10609 (N_10609,N_9954,N_9843);
xnor U10610 (N_10610,N_9667,N_9027);
or U10611 (N_10611,N_9553,N_8579);
or U10612 (N_10612,N_9452,N_9071);
xnor U10613 (N_10613,N_9787,N_8907);
nor U10614 (N_10614,N_8400,N_8991);
nand U10615 (N_10615,N_8671,N_9387);
or U10616 (N_10616,N_9252,N_8229);
xnor U10617 (N_10617,N_8039,N_8761);
or U10618 (N_10618,N_9016,N_8264);
or U10619 (N_10619,N_8941,N_8412);
xnor U10620 (N_10620,N_8669,N_8755);
nor U10621 (N_10621,N_8259,N_8666);
xnor U10622 (N_10622,N_8686,N_8094);
and U10623 (N_10623,N_8505,N_9540);
nand U10624 (N_10624,N_9291,N_9438);
or U10625 (N_10625,N_9738,N_8343);
nand U10626 (N_10626,N_9674,N_8774);
or U10627 (N_10627,N_8074,N_8872);
and U10628 (N_10628,N_9222,N_8065);
nor U10629 (N_10629,N_8826,N_9621);
xor U10630 (N_10630,N_9394,N_9976);
xor U10631 (N_10631,N_9682,N_9577);
xor U10632 (N_10632,N_9431,N_8572);
and U10633 (N_10633,N_9501,N_9783);
and U10634 (N_10634,N_8509,N_9253);
nand U10635 (N_10635,N_9205,N_9121);
xnor U10636 (N_10636,N_8751,N_9509);
or U10637 (N_10637,N_8100,N_9264);
and U10638 (N_10638,N_8585,N_9875);
or U10639 (N_10639,N_9385,N_8210);
or U10640 (N_10640,N_9145,N_9042);
or U10641 (N_10641,N_8943,N_8424);
nor U10642 (N_10642,N_8467,N_8828);
or U10643 (N_10643,N_8142,N_8387);
nand U10644 (N_10644,N_9839,N_8147);
and U10645 (N_10645,N_9309,N_8908);
and U10646 (N_10646,N_9428,N_9713);
or U10647 (N_10647,N_8489,N_8763);
and U10648 (N_10648,N_8873,N_9669);
xnor U10649 (N_10649,N_9351,N_9912);
nor U10650 (N_10650,N_8983,N_9492);
xor U10651 (N_10651,N_9115,N_9892);
and U10652 (N_10652,N_9152,N_9857);
xnor U10653 (N_10653,N_9656,N_9091);
or U10654 (N_10654,N_9140,N_8848);
and U10655 (N_10655,N_8736,N_8652);
or U10656 (N_10656,N_9303,N_9173);
nand U10657 (N_10657,N_8599,N_8859);
or U10658 (N_10658,N_8349,N_9364);
nor U10659 (N_10659,N_8117,N_8906);
xor U10660 (N_10660,N_8200,N_9170);
or U10661 (N_10661,N_8982,N_9488);
or U10662 (N_10662,N_9956,N_9934);
or U10663 (N_10663,N_8347,N_8079);
or U10664 (N_10664,N_8980,N_8199);
and U10665 (N_10665,N_8649,N_8293);
nand U10666 (N_10666,N_8954,N_8838);
nor U10667 (N_10667,N_9648,N_8996);
or U10668 (N_10668,N_8769,N_9633);
xor U10669 (N_10669,N_9451,N_9720);
xor U10670 (N_10670,N_9733,N_8303);
nor U10671 (N_10671,N_9639,N_9024);
and U10672 (N_10672,N_8172,N_9816);
nor U10673 (N_10673,N_9490,N_8672);
xnor U10674 (N_10674,N_8894,N_8116);
xor U10675 (N_10675,N_8164,N_8820);
or U10676 (N_10676,N_8606,N_9311);
nand U10677 (N_10677,N_8677,N_9548);
xor U10678 (N_10678,N_8897,N_9212);
nor U10679 (N_10679,N_8354,N_8634);
and U10680 (N_10680,N_8365,N_9353);
and U10681 (N_10681,N_9068,N_8626);
nor U10682 (N_10682,N_9084,N_8005);
or U10683 (N_10683,N_9082,N_9437);
nor U10684 (N_10684,N_8822,N_9420);
or U10685 (N_10685,N_8244,N_9186);
xor U10686 (N_10686,N_8255,N_9894);
nand U10687 (N_10687,N_9126,N_9019);
nor U10688 (N_10688,N_9167,N_9395);
nand U10689 (N_10689,N_9256,N_9520);
and U10690 (N_10690,N_9649,N_9064);
xor U10691 (N_10691,N_8876,N_8348);
nand U10692 (N_10692,N_9932,N_8474);
xor U10693 (N_10693,N_8780,N_8438);
xor U10694 (N_10694,N_8274,N_9982);
or U10695 (N_10695,N_8175,N_9330);
nand U10696 (N_10696,N_8558,N_9885);
nor U10697 (N_10697,N_8502,N_8974);
nand U10698 (N_10698,N_9984,N_9642);
and U10699 (N_10699,N_9882,N_8716);
and U10700 (N_10700,N_9240,N_9163);
nand U10701 (N_10701,N_9026,N_8129);
or U10702 (N_10702,N_9475,N_8887);
and U10703 (N_10703,N_9703,N_9228);
or U10704 (N_10704,N_8655,N_8028);
xor U10705 (N_10705,N_9873,N_9215);
nor U10706 (N_10706,N_8211,N_9896);
and U10707 (N_10707,N_9372,N_8428);
or U10708 (N_10708,N_9835,N_8500);
and U10709 (N_10709,N_8636,N_8928);
and U10710 (N_10710,N_9325,N_8102);
xor U10711 (N_10711,N_9672,N_8808);
or U10712 (N_10712,N_9579,N_9898);
nor U10713 (N_10713,N_9206,N_9337);
nor U10714 (N_10714,N_9563,N_8840);
nor U10715 (N_10715,N_8720,N_9004);
xnor U10716 (N_10716,N_8317,N_9809);
and U10717 (N_10717,N_8825,N_8900);
nor U10718 (N_10718,N_9238,N_8410);
nand U10719 (N_10719,N_8527,N_9109);
nor U10720 (N_10720,N_8099,N_8862);
and U10721 (N_10721,N_8064,N_8465);
or U10722 (N_10722,N_8802,N_8243);
nand U10723 (N_10723,N_8281,N_8008);
or U10724 (N_10724,N_9179,N_9935);
or U10725 (N_10725,N_9950,N_8987);
and U10726 (N_10726,N_9331,N_9366);
nand U10727 (N_10727,N_9789,N_8699);
nand U10728 (N_10728,N_9494,N_8362);
nand U10729 (N_10729,N_9693,N_9362);
or U10730 (N_10730,N_8051,N_9507);
and U10731 (N_10731,N_8083,N_9187);
xor U10732 (N_10732,N_9587,N_9476);
xnor U10733 (N_10733,N_8915,N_9518);
xor U10734 (N_10734,N_9598,N_9953);
nand U10735 (N_10735,N_8499,N_9051);
and U10736 (N_10736,N_9283,N_8192);
and U10737 (N_10737,N_8587,N_8644);
or U10738 (N_10738,N_9417,N_9658);
xor U10739 (N_10739,N_9844,N_8110);
xnor U10740 (N_10740,N_9555,N_8503);
nand U10741 (N_10741,N_9944,N_8220);
nor U10742 (N_10742,N_9998,N_8045);
nand U10743 (N_10743,N_8927,N_9182);
xnor U10744 (N_10744,N_9439,N_8197);
nor U10745 (N_10745,N_8373,N_9666);
xor U10746 (N_10746,N_9448,N_8835);
nor U10747 (N_10747,N_8890,N_8867);
nand U10748 (N_10748,N_9341,N_8481);
xnor U10749 (N_10749,N_9255,N_9689);
or U10750 (N_10750,N_9262,N_8056);
nand U10751 (N_10751,N_8141,N_8214);
and U10752 (N_10752,N_9781,N_8590);
nor U10753 (N_10753,N_8733,N_8766);
xor U10754 (N_10754,N_9275,N_8496);
nand U10755 (N_10755,N_9000,N_9822);
nand U10756 (N_10756,N_9687,N_9708);
nor U10757 (N_10757,N_8691,N_8262);
and U10758 (N_10758,N_9710,N_8667);
nor U10759 (N_10759,N_9350,N_9241);
and U10760 (N_10760,N_9946,N_9105);
nor U10761 (N_10761,N_8380,N_9166);
and U10762 (N_10762,N_8852,N_9943);
nor U10763 (N_10763,N_9020,N_9174);
nor U10764 (N_10764,N_8345,N_9695);
nor U10765 (N_10765,N_8750,N_8724);
or U10766 (N_10766,N_9319,N_9650);
or U10767 (N_10767,N_8592,N_8549);
and U10768 (N_10768,N_9292,N_9230);
or U10769 (N_10769,N_8535,N_9504);
or U10770 (N_10770,N_8025,N_9061);
nand U10771 (N_10771,N_9237,N_8745);
xnor U10772 (N_10772,N_8895,N_9594);
or U10773 (N_10773,N_9937,N_8075);
and U10774 (N_10774,N_9129,N_8934);
xnor U10775 (N_10775,N_9060,N_8408);
or U10776 (N_10776,N_9226,N_8014);
nor U10777 (N_10777,N_8207,N_8050);
xor U10778 (N_10778,N_8057,N_8012);
nand U10779 (N_10779,N_9755,N_8919);
and U10780 (N_10780,N_9436,N_9698);
nand U10781 (N_10781,N_9375,N_8153);
xnor U10782 (N_10782,N_8650,N_8219);
nand U10783 (N_10783,N_9793,N_8409);
nor U10784 (N_10784,N_9919,N_9736);
xor U10785 (N_10785,N_9908,N_8007);
xnor U10786 (N_10786,N_8573,N_8746);
nand U10787 (N_10787,N_8307,N_9419);
xnor U10788 (N_10788,N_8891,N_9500);
nand U10789 (N_10789,N_8168,N_9643);
xor U10790 (N_10790,N_8844,N_8547);
or U10791 (N_10791,N_8011,N_9349);
and U10792 (N_10792,N_9711,N_9081);
or U10793 (N_10793,N_9257,N_9392);
nor U10794 (N_10794,N_9697,N_9118);
xor U10795 (N_10795,N_8000,N_9905);
or U10796 (N_10796,N_8314,N_9752);
or U10797 (N_10797,N_8913,N_9002);
nand U10798 (N_10798,N_8545,N_8883);
nor U10799 (N_10799,N_9705,N_8871);
xnor U10800 (N_10800,N_8319,N_9993);
and U10801 (N_10801,N_8107,N_9033);
and U10802 (N_10802,N_8454,N_9551);
and U10803 (N_10803,N_9418,N_8680);
nand U10804 (N_10804,N_8316,N_9865);
nand U10805 (N_10805,N_8217,N_9312);
xor U10806 (N_10806,N_8236,N_9635);
nor U10807 (N_10807,N_9676,N_8162);
or U10808 (N_10808,N_9988,N_9147);
and U10809 (N_10809,N_8601,N_9416);
nor U10810 (N_10810,N_8727,N_9900);
xnor U10811 (N_10811,N_9306,N_8088);
nor U10812 (N_10812,N_9881,N_9859);
and U10813 (N_10813,N_9286,N_9581);
xnor U10814 (N_10814,N_9067,N_8914);
nor U10815 (N_10815,N_9758,N_8577);
and U10816 (N_10816,N_9679,N_9745);
or U10817 (N_10817,N_9638,N_8068);
or U10818 (N_10818,N_9961,N_8422);
nor U10819 (N_10819,N_8268,N_9886);
nand U10820 (N_10820,N_8190,N_8203);
nand U10821 (N_10821,N_9007,N_8061);
nand U10822 (N_10822,N_9046,N_8998);
nand U10823 (N_10823,N_9057,N_8702);
nand U10824 (N_10824,N_9124,N_9879);
xor U10825 (N_10825,N_9077,N_9314);
and U10826 (N_10826,N_9683,N_9402);
nand U10827 (N_10827,N_8226,N_9197);
xor U10828 (N_10828,N_8957,N_9600);
or U10829 (N_10829,N_8832,N_8022);
and U10830 (N_10830,N_8127,N_8940);
nand U10831 (N_10831,N_8093,N_8305);
nor U10832 (N_10832,N_9585,N_8004);
and U10833 (N_10833,N_9571,N_8238);
nand U10834 (N_10834,N_8054,N_8455);
nor U10835 (N_10835,N_9049,N_8952);
nor U10836 (N_10836,N_9539,N_8740);
nor U10837 (N_10837,N_8163,N_8865);
xnor U10838 (N_10838,N_9510,N_8742);
xnor U10839 (N_10839,N_9817,N_8090);
or U10840 (N_10840,N_8546,N_8256);
nand U10841 (N_10841,N_9975,N_8931);
and U10842 (N_10842,N_8300,N_8138);
nand U10843 (N_10843,N_8456,N_8131);
nor U10844 (N_10844,N_9218,N_8679);
or U10845 (N_10845,N_8892,N_9454);
and U10846 (N_10846,N_8106,N_8476);
or U10847 (N_10847,N_9321,N_8169);
and U10848 (N_10848,N_9829,N_8406);
nor U10849 (N_10849,N_9995,N_8706);
and U10850 (N_10850,N_9098,N_8182);
nand U10851 (N_10851,N_8125,N_9893);
nor U10852 (N_10852,N_8508,N_9728);
nand U10853 (N_10853,N_8992,N_9570);
xor U10854 (N_10854,N_8177,N_8791);
nand U10855 (N_10855,N_9177,N_8080);
nand U10856 (N_10856,N_8202,N_9826);
nand U10857 (N_10857,N_9467,N_8831);
nand U10858 (N_10858,N_9365,N_9902);
and U10859 (N_10859,N_9499,N_9200);
nand U10860 (N_10860,N_9818,N_9223);
or U10861 (N_10861,N_9890,N_8342);
nor U10862 (N_10862,N_9069,N_9444);
or U10863 (N_10863,N_8708,N_8525);
nor U10864 (N_10864,N_8361,N_9623);
xor U10865 (N_10865,N_9700,N_8239);
and U10866 (N_10866,N_8775,N_9516);
nand U10867 (N_10867,N_9546,N_9227);
nand U10868 (N_10868,N_8562,N_9690);
xor U10869 (N_10869,N_8002,N_8651);
xnor U10870 (N_10870,N_9503,N_8605);
xor U10871 (N_10871,N_8191,N_8904);
nand U10872 (N_10872,N_8112,N_8249);
nand U10873 (N_10873,N_9596,N_8809);
or U10874 (N_10874,N_9731,N_9277);
and U10875 (N_10875,N_9471,N_9455);
xnor U10876 (N_10876,N_8849,N_8248);
nor U10877 (N_10877,N_9586,N_9133);
xnor U10878 (N_10878,N_9298,N_8420);
xor U10879 (N_10879,N_8584,N_9940);
xor U10880 (N_10880,N_9062,N_8149);
and U10881 (N_10881,N_8754,N_9423);
nand U10882 (N_10882,N_9798,N_8024);
and U10883 (N_10883,N_9702,N_8781);
xor U10884 (N_10884,N_9195,N_9604);
xor U10885 (N_10885,N_8108,N_8145);
nand U10886 (N_10886,N_9485,N_9640);
nor U10887 (N_10887,N_9617,N_8124);
nand U10888 (N_10888,N_9017,N_9840);
nor U10889 (N_10889,N_9945,N_8159);
and U10890 (N_10890,N_8167,N_9629);
xnor U10891 (N_10891,N_9729,N_8046);
and U10892 (N_10892,N_9823,N_8295);
and U10893 (N_10893,N_9532,N_9433);
nand U10894 (N_10894,N_9701,N_8799);
or U10895 (N_10895,N_8557,N_9601);
and U10896 (N_10896,N_9139,N_8875);
and U10897 (N_10897,N_9721,N_8944);
nand U10898 (N_10898,N_8060,N_9855);
or U10899 (N_10899,N_8257,N_8744);
and U10900 (N_10900,N_9114,N_9107);
nor U10901 (N_10901,N_9517,N_8743);
and U10902 (N_10902,N_9202,N_9719);
and U10903 (N_10903,N_9735,N_8417);
xnor U10904 (N_10904,N_9958,N_8712);
xor U10905 (N_10905,N_8824,N_9806);
xnor U10906 (N_10906,N_9678,N_8433);
or U10907 (N_10907,N_8807,N_9389);
nand U10908 (N_10908,N_9962,N_8494);
xor U10909 (N_10909,N_8076,N_8123);
and U10910 (N_10910,N_8445,N_9646);
nand U10911 (N_10911,N_8856,N_9722);
xor U10912 (N_10912,N_8294,N_8098);
and U10913 (N_10913,N_9768,N_9249);
nand U10914 (N_10914,N_9788,N_9146);
nor U10915 (N_10915,N_8571,N_9340);
xnor U10916 (N_10916,N_8700,N_8978);
nand U10917 (N_10917,N_8504,N_8759);
nand U10918 (N_10918,N_8760,N_8330);
and U10919 (N_10919,N_9819,N_9605);
and U10920 (N_10920,N_8646,N_8516);
or U10921 (N_10921,N_8837,N_8768);
or U10922 (N_10922,N_9156,N_8812);
and U10923 (N_10923,N_8488,N_9162);
nor U10924 (N_10924,N_9870,N_9429);
and U10925 (N_10925,N_9769,N_9554);
xnor U10926 (N_10926,N_9315,N_9032);
xnor U10927 (N_10927,N_9861,N_9293);
nor U10928 (N_10928,N_8964,N_8038);
nor U10929 (N_10929,N_9208,N_9664);
xor U10930 (N_10930,N_9159,N_8165);
nand U10931 (N_10931,N_8911,N_9379);
nor U10932 (N_10932,N_8938,N_8922);
nor U10933 (N_10933,N_9442,N_8353);
nor U10934 (N_10934,N_8227,N_9189);
or U10935 (N_10935,N_8322,N_8398);
nand U10936 (N_10936,N_9513,N_9936);
nand U10937 (N_10937,N_9138,N_8747);
xor U10938 (N_10938,N_9481,N_8818);
or U10939 (N_10939,N_8136,N_9301);
nand U10940 (N_10940,N_9785,N_9899);
or U10941 (N_10941,N_9102,N_9006);
nor U10942 (N_10942,N_8048,N_8444);
xnor U10943 (N_10943,N_8103,N_8413);
nor U10944 (N_10944,N_9888,N_8144);
and U10945 (N_10945,N_8497,N_8602);
or U10946 (N_10946,N_9796,N_8221);
xor U10947 (N_10947,N_8748,N_8723);
xnor U10948 (N_10948,N_8819,N_9058);
nand U10949 (N_10949,N_8622,N_8320);
xnor U10950 (N_10950,N_9578,N_9035);
or U10951 (N_10951,N_8963,N_9388);
nor U10952 (N_10952,N_8148,N_8414);
nand U10953 (N_10953,N_9543,N_9407);
nand U10954 (N_10954,N_8251,N_8888);
xor U10955 (N_10955,N_9012,N_9149);
nand U10956 (N_10956,N_9794,N_9465);
and U10957 (N_10957,N_8363,N_9654);
and U10958 (N_10958,N_8393,N_9427);
xor U10959 (N_10959,N_9523,N_9651);
xnor U10960 (N_10960,N_9104,N_9478);
or U10961 (N_10961,N_8323,N_9990);
xnor U10962 (N_10962,N_9834,N_9968);
xor U10963 (N_10963,N_8358,N_8861);
xnor U10964 (N_10964,N_8731,N_9969);
nor U10965 (N_10965,N_9287,N_8947);
and U10966 (N_10966,N_9194,N_8485);
nand U10967 (N_10967,N_9415,N_9910);
xor U10968 (N_10968,N_8681,N_8204);
or U10969 (N_10969,N_8341,N_8990);
nor U10970 (N_10970,N_9986,N_8659);
or U10971 (N_10971,N_9390,N_9838);
and U10972 (N_10972,N_8854,N_8639);
nor U10973 (N_10973,N_9248,N_8335);
nor U10974 (N_10974,N_8381,N_9048);
nor U10975 (N_10975,N_9038,N_8441);
nand U10976 (N_10976,N_8092,N_8533);
xnor U10977 (N_10977,N_9832,N_8958);
or U10978 (N_10978,N_9727,N_9522);
xor U10979 (N_10979,N_9918,N_8936);
and U10980 (N_10980,N_8324,N_8925);
xor U10981 (N_10981,N_9261,N_9957);
nand U10982 (N_10982,N_8806,N_9408);
nand U10983 (N_10983,N_8773,N_8350);
nor U10984 (N_10984,N_9673,N_9599);
nor U10985 (N_10985,N_9906,N_8152);
xor U10986 (N_10986,N_8841,N_9889);
nand U10987 (N_10987,N_9997,N_8036);
nand U10988 (N_10988,N_9092,N_8608);
nor U10989 (N_10989,N_8442,N_8376);
nor U10990 (N_10990,N_9462,N_8015);
nor U10991 (N_10991,N_9704,N_9347);
xnor U10992 (N_10992,N_9749,N_8059);
or U10993 (N_10993,N_8359,N_9100);
xor U10994 (N_10994,N_9734,N_8580);
or U10995 (N_10995,N_8640,N_8286);
xnor U10996 (N_10996,N_9723,N_9821);
xor U10997 (N_10997,N_9381,N_8029);
nand U10998 (N_10998,N_9558,N_9125);
nor U10999 (N_10999,N_8953,N_8574);
xor U11000 (N_11000,N_9886,N_9535);
and U11001 (N_11001,N_8524,N_9869);
and U11002 (N_11002,N_8495,N_8283);
xor U11003 (N_11003,N_8855,N_8346);
or U11004 (N_11004,N_9815,N_8676);
and U11005 (N_11005,N_9538,N_8711);
nor U11006 (N_11006,N_8341,N_9709);
or U11007 (N_11007,N_9713,N_8619);
nor U11008 (N_11008,N_8355,N_9406);
xnor U11009 (N_11009,N_8267,N_8720);
nand U11010 (N_11010,N_8743,N_9123);
xnor U11011 (N_11011,N_8143,N_8094);
nand U11012 (N_11012,N_8580,N_8709);
xnor U11013 (N_11013,N_9015,N_9470);
nor U11014 (N_11014,N_8440,N_8047);
xor U11015 (N_11015,N_8442,N_9886);
nor U11016 (N_11016,N_9215,N_9214);
and U11017 (N_11017,N_8014,N_8646);
xnor U11018 (N_11018,N_8411,N_8048);
and U11019 (N_11019,N_9037,N_9804);
or U11020 (N_11020,N_9294,N_8129);
xnor U11021 (N_11021,N_8551,N_9735);
nand U11022 (N_11022,N_8392,N_9358);
and U11023 (N_11023,N_8629,N_9409);
and U11024 (N_11024,N_8843,N_9436);
and U11025 (N_11025,N_8783,N_8206);
nand U11026 (N_11026,N_8220,N_9425);
nor U11027 (N_11027,N_9853,N_8527);
nand U11028 (N_11028,N_9488,N_9557);
or U11029 (N_11029,N_8480,N_8664);
nor U11030 (N_11030,N_9688,N_8871);
or U11031 (N_11031,N_8979,N_8363);
nor U11032 (N_11032,N_8163,N_8665);
nand U11033 (N_11033,N_8104,N_8771);
nand U11034 (N_11034,N_8176,N_8731);
or U11035 (N_11035,N_9407,N_8458);
xor U11036 (N_11036,N_9148,N_8954);
xnor U11037 (N_11037,N_9324,N_8147);
nand U11038 (N_11038,N_9627,N_8772);
nand U11039 (N_11039,N_8372,N_9265);
nor U11040 (N_11040,N_8276,N_8134);
xnor U11041 (N_11041,N_8081,N_9016);
xor U11042 (N_11042,N_8293,N_9543);
xor U11043 (N_11043,N_9139,N_9599);
nand U11044 (N_11044,N_9118,N_8825);
xor U11045 (N_11045,N_8154,N_9233);
and U11046 (N_11046,N_8167,N_8947);
nor U11047 (N_11047,N_9314,N_8219);
xnor U11048 (N_11048,N_9068,N_8274);
nor U11049 (N_11049,N_9970,N_8941);
or U11050 (N_11050,N_9146,N_9570);
or U11051 (N_11051,N_9458,N_9060);
and U11052 (N_11052,N_9531,N_9443);
nor U11053 (N_11053,N_8990,N_8580);
or U11054 (N_11054,N_8533,N_8353);
nand U11055 (N_11055,N_8408,N_8153);
xnor U11056 (N_11056,N_9892,N_8228);
nand U11057 (N_11057,N_9579,N_9445);
xor U11058 (N_11058,N_9921,N_9195);
and U11059 (N_11059,N_9692,N_8606);
or U11060 (N_11060,N_8045,N_9319);
nand U11061 (N_11061,N_9378,N_9521);
or U11062 (N_11062,N_8957,N_8944);
nor U11063 (N_11063,N_9972,N_8650);
xnor U11064 (N_11064,N_9718,N_9842);
nand U11065 (N_11065,N_8036,N_9326);
nand U11066 (N_11066,N_9867,N_8246);
nor U11067 (N_11067,N_8246,N_9269);
nand U11068 (N_11068,N_9635,N_9652);
nor U11069 (N_11069,N_9751,N_8890);
or U11070 (N_11070,N_9125,N_8949);
and U11071 (N_11071,N_8607,N_8704);
nor U11072 (N_11072,N_9594,N_9086);
xor U11073 (N_11073,N_8223,N_9795);
or U11074 (N_11074,N_9028,N_8849);
or U11075 (N_11075,N_8970,N_8648);
nor U11076 (N_11076,N_9935,N_9663);
and U11077 (N_11077,N_9246,N_9255);
or U11078 (N_11078,N_8491,N_8141);
nand U11079 (N_11079,N_9341,N_8689);
nand U11080 (N_11080,N_9429,N_9292);
nor U11081 (N_11081,N_8141,N_8339);
and U11082 (N_11082,N_9493,N_9195);
or U11083 (N_11083,N_8026,N_9460);
or U11084 (N_11084,N_9296,N_9332);
and U11085 (N_11085,N_8070,N_8327);
or U11086 (N_11086,N_8061,N_8872);
and U11087 (N_11087,N_9538,N_8664);
or U11088 (N_11088,N_9008,N_8567);
or U11089 (N_11089,N_8692,N_8967);
or U11090 (N_11090,N_9990,N_8377);
nand U11091 (N_11091,N_9399,N_9723);
nand U11092 (N_11092,N_9726,N_9376);
nand U11093 (N_11093,N_9744,N_8831);
nand U11094 (N_11094,N_9582,N_9166);
or U11095 (N_11095,N_9293,N_9929);
nor U11096 (N_11096,N_8644,N_9486);
nor U11097 (N_11097,N_9315,N_9418);
nor U11098 (N_11098,N_8151,N_9604);
and U11099 (N_11099,N_8941,N_8543);
xnor U11100 (N_11100,N_9136,N_9030);
nand U11101 (N_11101,N_9140,N_9847);
nor U11102 (N_11102,N_8569,N_8051);
xor U11103 (N_11103,N_8825,N_8030);
nor U11104 (N_11104,N_9127,N_9199);
or U11105 (N_11105,N_9636,N_9655);
xnor U11106 (N_11106,N_8064,N_8111);
nand U11107 (N_11107,N_8893,N_9418);
or U11108 (N_11108,N_9036,N_8280);
nand U11109 (N_11109,N_9909,N_9424);
nor U11110 (N_11110,N_9974,N_8364);
or U11111 (N_11111,N_9420,N_8412);
nand U11112 (N_11112,N_8318,N_9218);
or U11113 (N_11113,N_8233,N_9032);
and U11114 (N_11114,N_9988,N_8621);
nand U11115 (N_11115,N_9697,N_8096);
or U11116 (N_11116,N_8911,N_9052);
xor U11117 (N_11117,N_9652,N_8092);
or U11118 (N_11118,N_9388,N_9948);
and U11119 (N_11119,N_8874,N_8200);
or U11120 (N_11120,N_8659,N_8743);
and U11121 (N_11121,N_9953,N_9956);
and U11122 (N_11122,N_8984,N_8752);
nand U11123 (N_11123,N_8376,N_9914);
nor U11124 (N_11124,N_8723,N_8406);
xnor U11125 (N_11125,N_8644,N_9463);
and U11126 (N_11126,N_8694,N_9830);
xnor U11127 (N_11127,N_8646,N_8766);
xnor U11128 (N_11128,N_8092,N_9452);
xnor U11129 (N_11129,N_9459,N_8832);
or U11130 (N_11130,N_8696,N_9282);
and U11131 (N_11131,N_8687,N_9075);
or U11132 (N_11132,N_9242,N_9683);
xnor U11133 (N_11133,N_8030,N_9440);
or U11134 (N_11134,N_9965,N_8595);
xor U11135 (N_11135,N_8340,N_9012);
nor U11136 (N_11136,N_8595,N_9856);
nand U11137 (N_11137,N_9101,N_9377);
xnor U11138 (N_11138,N_9332,N_8895);
and U11139 (N_11139,N_9228,N_9586);
or U11140 (N_11140,N_8754,N_8686);
and U11141 (N_11141,N_8866,N_9902);
xor U11142 (N_11142,N_9177,N_8625);
or U11143 (N_11143,N_9449,N_8746);
or U11144 (N_11144,N_8809,N_9410);
nand U11145 (N_11145,N_9677,N_9929);
nand U11146 (N_11146,N_9726,N_8432);
nor U11147 (N_11147,N_9723,N_9772);
nor U11148 (N_11148,N_9112,N_8500);
nand U11149 (N_11149,N_8295,N_9473);
and U11150 (N_11150,N_8869,N_9328);
and U11151 (N_11151,N_9768,N_9673);
or U11152 (N_11152,N_9447,N_9981);
xor U11153 (N_11153,N_8537,N_8056);
nor U11154 (N_11154,N_9769,N_9543);
and U11155 (N_11155,N_8633,N_9427);
or U11156 (N_11156,N_8669,N_9763);
and U11157 (N_11157,N_8340,N_9581);
xor U11158 (N_11158,N_9828,N_9605);
or U11159 (N_11159,N_9987,N_8373);
and U11160 (N_11160,N_8547,N_9812);
xor U11161 (N_11161,N_9519,N_8373);
nand U11162 (N_11162,N_8769,N_9636);
xnor U11163 (N_11163,N_9185,N_8815);
xnor U11164 (N_11164,N_8860,N_9553);
or U11165 (N_11165,N_9077,N_9385);
or U11166 (N_11166,N_9071,N_8129);
nand U11167 (N_11167,N_8490,N_8667);
xor U11168 (N_11168,N_9489,N_8276);
nor U11169 (N_11169,N_8598,N_8813);
nor U11170 (N_11170,N_9470,N_8656);
nor U11171 (N_11171,N_9511,N_8757);
or U11172 (N_11172,N_8360,N_8297);
xnor U11173 (N_11173,N_9214,N_8516);
and U11174 (N_11174,N_8669,N_8668);
or U11175 (N_11175,N_8056,N_8194);
xor U11176 (N_11176,N_9421,N_9027);
xor U11177 (N_11177,N_9774,N_8459);
nor U11178 (N_11178,N_8380,N_9452);
xnor U11179 (N_11179,N_9307,N_8004);
nor U11180 (N_11180,N_8235,N_9200);
xor U11181 (N_11181,N_9611,N_9905);
nor U11182 (N_11182,N_8710,N_8670);
xor U11183 (N_11183,N_9144,N_9060);
or U11184 (N_11184,N_9687,N_9099);
and U11185 (N_11185,N_8206,N_9443);
and U11186 (N_11186,N_9802,N_8943);
nor U11187 (N_11187,N_8547,N_8356);
nand U11188 (N_11188,N_9329,N_8619);
xor U11189 (N_11189,N_9613,N_8519);
xor U11190 (N_11190,N_8921,N_8505);
and U11191 (N_11191,N_9563,N_9805);
and U11192 (N_11192,N_9071,N_8220);
nor U11193 (N_11193,N_8807,N_8664);
and U11194 (N_11194,N_9297,N_9394);
nor U11195 (N_11195,N_8242,N_9693);
and U11196 (N_11196,N_9543,N_9356);
and U11197 (N_11197,N_8437,N_8587);
xor U11198 (N_11198,N_8004,N_8183);
or U11199 (N_11199,N_9719,N_8837);
or U11200 (N_11200,N_8198,N_9853);
or U11201 (N_11201,N_9645,N_8061);
nor U11202 (N_11202,N_8620,N_9997);
or U11203 (N_11203,N_9596,N_8283);
nand U11204 (N_11204,N_8380,N_9135);
xnor U11205 (N_11205,N_8944,N_8909);
nand U11206 (N_11206,N_9779,N_9524);
nand U11207 (N_11207,N_9106,N_8541);
xnor U11208 (N_11208,N_9516,N_9204);
nor U11209 (N_11209,N_8850,N_9084);
nand U11210 (N_11210,N_9285,N_9843);
and U11211 (N_11211,N_9751,N_9197);
nor U11212 (N_11212,N_9219,N_9518);
xnor U11213 (N_11213,N_8567,N_8297);
nor U11214 (N_11214,N_8349,N_9701);
nor U11215 (N_11215,N_9909,N_8139);
nand U11216 (N_11216,N_8389,N_9420);
xor U11217 (N_11217,N_9468,N_9238);
and U11218 (N_11218,N_9591,N_8629);
nand U11219 (N_11219,N_8314,N_8585);
nand U11220 (N_11220,N_9626,N_9538);
nand U11221 (N_11221,N_8692,N_9338);
xor U11222 (N_11222,N_8601,N_9875);
xnor U11223 (N_11223,N_9314,N_9587);
nand U11224 (N_11224,N_9894,N_9135);
nand U11225 (N_11225,N_8199,N_9424);
and U11226 (N_11226,N_9859,N_8962);
xnor U11227 (N_11227,N_9786,N_8973);
or U11228 (N_11228,N_8119,N_8897);
nand U11229 (N_11229,N_8925,N_8785);
and U11230 (N_11230,N_9453,N_8184);
and U11231 (N_11231,N_8395,N_9837);
nand U11232 (N_11232,N_8191,N_9060);
nand U11233 (N_11233,N_8321,N_8355);
and U11234 (N_11234,N_8565,N_8538);
xnor U11235 (N_11235,N_9963,N_9302);
nor U11236 (N_11236,N_9294,N_8173);
nor U11237 (N_11237,N_9624,N_8555);
and U11238 (N_11238,N_9839,N_8891);
and U11239 (N_11239,N_9326,N_9578);
xor U11240 (N_11240,N_8372,N_8003);
or U11241 (N_11241,N_8477,N_9103);
or U11242 (N_11242,N_9720,N_9797);
nand U11243 (N_11243,N_8634,N_8590);
nor U11244 (N_11244,N_8312,N_8353);
nand U11245 (N_11245,N_9657,N_8571);
nor U11246 (N_11246,N_8911,N_8295);
xor U11247 (N_11247,N_8699,N_9862);
nand U11248 (N_11248,N_9433,N_9603);
xnor U11249 (N_11249,N_9528,N_8088);
or U11250 (N_11250,N_9612,N_8362);
xor U11251 (N_11251,N_9362,N_9626);
or U11252 (N_11252,N_8279,N_9736);
and U11253 (N_11253,N_9122,N_8912);
nand U11254 (N_11254,N_9166,N_9397);
nor U11255 (N_11255,N_8132,N_8860);
nand U11256 (N_11256,N_8483,N_9329);
or U11257 (N_11257,N_9032,N_9558);
nor U11258 (N_11258,N_9844,N_9441);
or U11259 (N_11259,N_9364,N_9245);
or U11260 (N_11260,N_9455,N_8000);
xor U11261 (N_11261,N_8313,N_8852);
nor U11262 (N_11262,N_9678,N_8476);
xnor U11263 (N_11263,N_9485,N_8285);
xnor U11264 (N_11264,N_9649,N_9435);
or U11265 (N_11265,N_9543,N_9588);
and U11266 (N_11266,N_9268,N_8522);
xor U11267 (N_11267,N_9933,N_9358);
nor U11268 (N_11268,N_8135,N_9486);
or U11269 (N_11269,N_8393,N_9019);
nand U11270 (N_11270,N_9810,N_9947);
xor U11271 (N_11271,N_8920,N_8307);
xnor U11272 (N_11272,N_8211,N_8958);
xor U11273 (N_11273,N_9084,N_9587);
or U11274 (N_11274,N_8029,N_9873);
or U11275 (N_11275,N_8118,N_9808);
and U11276 (N_11276,N_8272,N_8943);
and U11277 (N_11277,N_9024,N_8140);
nand U11278 (N_11278,N_9679,N_9912);
xor U11279 (N_11279,N_9921,N_8717);
nor U11280 (N_11280,N_8946,N_8036);
nor U11281 (N_11281,N_9282,N_9570);
and U11282 (N_11282,N_9278,N_9475);
nor U11283 (N_11283,N_9240,N_8887);
nor U11284 (N_11284,N_8223,N_9313);
xor U11285 (N_11285,N_9355,N_8037);
nand U11286 (N_11286,N_9652,N_9934);
and U11287 (N_11287,N_8741,N_8093);
xor U11288 (N_11288,N_9800,N_9497);
nand U11289 (N_11289,N_8811,N_9528);
nor U11290 (N_11290,N_8347,N_9006);
nand U11291 (N_11291,N_9467,N_8107);
xor U11292 (N_11292,N_9264,N_8037);
xnor U11293 (N_11293,N_8269,N_8868);
nand U11294 (N_11294,N_8151,N_9328);
nand U11295 (N_11295,N_9411,N_8870);
and U11296 (N_11296,N_9627,N_9706);
and U11297 (N_11297,N_8246,N_9178);
xor U11298 (N_11298,N_8574,N_9404);
nand U11299 (N_11299,N_9238,N_9195);
or U11300 (N_11300,N_9950,N_8717);
or U11301 (N_11301,N_8829,N_8961);
xnor U11302 (N_11302,N_9909,N_8732);
nor U11303 (N_11303,N_8292,N_9069);
nor U11304 (N_11304,N_9736,N_9737);
nor U11305 (N_11305,N_9015,N_8648);
nor U11306 (N_11306,N_8493,N_9448);
nand U11307 (N_11307,N_8064,N_9908);
xor U11308 (N_11308,N_9713,N_8109);
xor U11309 (N_11309,N_8507,N_9734);
nand U11310 (N_11310,N_8436,N_9745);
nor U11311 (N_11311,N_9146,N_9525);
or U11312 (N_11312,N_8302,N_9170);
nand U11313 (N_11313,N_9152,N_9598);
and U11314 (N_11314,N_9415,N_9994);
or U11315 (N_11315,N_8673,N_9349);
or U11316 (N_11316,N_8541,N_9895);
or U11317 (N_11317,N_9530,N_8145);
nor U11318 (N_11318,N_9879,N_9471);
nor U11319 (N_11319,N_9644,N_8658);
and U11320 (N_11320,N_9113,N_9660);
or U11321 (N_11321,N_9795,N_9528);
nor U11322 (N_11322,N_8777,N_9341);
nand U11323 (N_11323,N_9274,N_8925);
nand U11324 (N_11324,N_9052,N_9093);
nor U11325 (N_11325,N_8839,N_8728);
or U11326 (N_11326,N_8125,N_8458);
nor U11327 (N_11327,N_8505,N_8648);
nor U11328 (N_11328,N_9037,N_9882);
nor U11329 (N_11329,N_9494,N_8469);
and U11330 (N_11330,N_8263,N_8404);
or U11331 (N_11331,N_9295,N_8891);
or U11332 (N_11332,N_9692,N_8969);
xnor U11333 (N_11333,N_9308,N_8891);
nor U11334 (N_11334,N_8024,N_8469);
and U11335 (N_11335,N_9240,N_8403);
and U11336 (N_11336,N_9971,N_8701);
nor U11337 (N_11337,N_9585,N_9222);
or U11338 (N_11338,N_8559,N_9487);
and U11339 (N_11339,N_8096,N_8499);
nor U11340 (N_11340,N_9743,N_8224);
nand U11341 (N_11341,N_9736,N_8223);
or U11342 (N_11342,N_9176,N_9616);
or U11343 (N_11343,N_9452,N_9424);
and U11344 (N_11344,N_8022,N_8043);
and U11345 (N_11345,N_8461,N_8174);
nand U11346 (N_11346,N_8221,N_8363);
and U11347 (N_11347,N_8998,N_9191);
and U11348 (N_11348,N_8430,N_8219);
nor U11349 (N_11349,N_9830,N_9709);
or U11350 (N_11350,N_9807,N_8593);
nand U11351 (N_11351,N_9390,N_9553);
nor U11352 (N_11352,N_9318,N_8368);
nor U11353 (N_11353,N_9184,N_9555);
or U11354 (N_11354,N_8687,N_9275);
nor U11355 (N_11355,N_9743,N_8841);
nand U11356 (N_11356,N_9001,N_8266);
nor U11357 (N_11357,N_8034,N_9948);
and U11358 (N_11358,N_8685,N_8678);
or U11359 (N_11359,N_9972,N_9694);
nand U11360 (N_11360,N_8396,N_9310);
nand U11361 (N_11361,N_8285,N_9103);
xnor U11362 (N_11362,N_8212,N_8575);
xnor U11363 (N_11363,N_8921,N_8626);
or U11364 (N_11364,N_9496,N_8930);
nand U11365 (N_11365,N_9846,N_8557);
nor U11366 (N_11366,N_8481,N_9713);
or U11367 (N_11367,N_9434,N_9126);
and U11368 (N_11368,N_8853,N_8929);
xnor U11369 (N_11369,N_9640,N_8707);
or U11370 (N_11370,N_8026,N_9842);
xnor U11371 (N_11371,N_8843,N_9672);
and U11372 (N_11372,N_9323,N_8682);
or U11373 (N_11373,N_8392,N_9970);
xor U11374 (N_11374,N_9043,N_8941);
nand U11375 (N_11375,N_9981,N_8421);
nand U11376 (N_11376,N_8267,N_8740);
nand U11377 (N_11377,N_9074,N_8721);
xor U11378 (N_11378,N_9800,N_8528);
nor U11379 (N_11379,N_9298,N_8704);
nand U11380 (N_11380,N_8141,N_9436);
nand U11381 (N_11381,N_9550,N_9206);
or U11382 (N_11382,N_9428,N_8816);
nand U11383 (N_11383,N_9744,N_8527);
nor U11384 (N_11384,N_9849,N_9682);
or U11385 (N_11385,N_8002,N_9564);
or U11386 (N_11386,N_9866,N_9961);
and U11387 (N_11387,N_9874,N_8651);
nand U11388 (N_11388,N_9395,N_8792);
nor U11389 (N_11389,N_9647,N_8617);
and U11390 (N_11390,N_8694,N_8501);
and U11391 (N_11391,N_8284,N_9615);
and U11392 (N_11392,N_9441,N_9989);
nand U11393 (N_11393,N_9297,N_9781);
and U11394 (N_11394,N_8240,N_8438);
nand U11395 (N_11395,N_9995,N_9962);
and U11396 (N_11396,N_8014,N_8289);
or U11397 (N_11397,N_9738,N_9427);
or U11398 (N_11398,N_8018,N_9483);
nand U11399 (N_11399,N_9282,N_9056);
and U11400 (N_11400,N_9479,N_8146);
xnor U11401 (N_11401,N_9126,N_9332);
or U11402 (N_11402,N_8835,N_9966);
nand U11403 (N_11403,N_8433,N_9227);
nand U11404 (N_11404,N_8418,N_9369);
nand U11405 (N_11405,N_8797,N_8385);
and U11406 (N_11406,N_9248,N_9809);
nor U11407 (N_11407,N_9042,N_9317);
nand U11408 (N_11408,N_9036,N_8400);
nand U11409 (N_11409,N_8734,N_9310);
nand U11410 (N_11410,N_9560,N_8543);
and U11411 (N_11411,N_9279,N_8836);
nand U11412 (N_11412,N_9723,N_8517);
and U11413 (N_11413,N_9424,N_8386);
nand U11414 (N_11414,N_8809,N_8419);
or U11415 (N_11415,N_8871,N_8685);
xor U11416 (N_11416,N_9332,N_9214);
nand U11417 (N_11417,N_9488,N_9201);
or U11418 (N_11418,N_8295,N_8060);
nand U11419 (N_11419,N_8210,N_9538);
xor U11420 (N_11420,N_8992,N_8218);
nand U11421 (N_11421,N_8358,N_9304);
nor U11422 (N_11422,N_8024,N_8510);
nor U11423 (N_11423,N_8862,N_9082);
and U11424 (N_11424,N_8384,N_9046);
or U11425 (N_11425,N_9497,N_8399);
nor U11426 (N_11426,N_8255,N_9034);
and U11427 (N_11427,N_8697,N_9210);
nor U11428 (N_11428,N_9432,N_8559);
nor U11429 (N_11429,N_9797,N_8416);
or U11430 (N_11430,N_9729,N_8891);
and U11431 (N_11431,N_9811,N_9567);
xor U11432 (N_11432,N_9926,N_9139);
nor U11433 (N_11433,N_9651,N_8833);
and U11434 (N_11434,N_9530,N_9320);
or U11435 (N_11435,N_9661,N_8847);
nand U11436 (N_11436,N_8046,N_9375);
and U11437 (N_11437,N_9690,N_9148);
nor U11438 (N_11438,N_8059,N_9595);
and U11439 (N_11439,N_8871,N_9576);
xnor U11440 (N_11440,N_8508,N_9129);
xnor U11441 (N_11441,N_8750,N_9231);
nand U11442 (N_11442,N_8800,N_8138);
and U11443 (N_11443,N_9992,N_9760);
xor U11444 (N_11444,N_9313,N_9669);
nor U11445 (N_11445,N_9829,N_9692);
nor U11446 (N_11446,N_9600,N_9312);
nand U11447 (N_11447,N_8590,N_8791);
or U11448 (N_11448,N_8228,N_9865);
and U11449 (N_11449,N_8869,N_9335);
or U11450 (N_11450,N_9364,N_8015);
and U11451 (N_11451,N_9563,N_9304);
nand U11452 (N_11452,N_8787,N_9591);
nand U11453 (N_11453,N_8283,N_9153);
xor U11454 (N_11454,N_8435,N_9561);
nand U11455 (N_11455,N_9663,N_8077);
and U11456 (N_11456,N_9455,N_9820);
or U11457 (N_11457,N_9110,N_8865);
xnor U11458 (N_11458,N_9420,N_9117);
nor U11459 (N_11459,N_8087,N_8705);
nor U11460 (N_11460,N_9916,N_8007);
or U11461 (N_11461,N_9740,N_8266);
or U11462 (N_11462,N_9782,N_8143);
nand U11463 (N_11463,N_8361,N_9956);
nand U11464 (N_11464,N_9471,N_9396);
nor U11465 (N_11465,N_8173,N_9904);
xor U11466 (N_11466,N_8165,N_9931);
and U11467 (N_11467,N_9517,N_8620);
nand U11468 (N_11468,N_9374,N_9249);
nand U11469 (N_11469,N_9752,N_9233);
nand U11470 (N_11470,N_9540,N_8137);
and U11471 (N_11471,N_8574,N_8428);
nand U11472 (N_11472,N_8973,N_8246);
or U11473 (N_11473,N_9771,N_8524);
nand U11474 (N_11474,N_8221,N_9382);
nor U11475 (N_11475,N_8650,N_8634);
nor U11476 (N_11476,N_9699,N_9852);
xnor U11477 (N_11477,N_8957,N_8054);
and U11478 (N_11478,N_9673,N_8449);
nor U11479 (N_11479,N_8906,N_8419);
xor U11480 (N_11480,N_9626,N_8276);
nand U11481 (N_11481,N_8021,N_8668);
nor U11482 (N_11482,N_9591,N_9779);
or U11483 (N_11483,N_8798,N_8708);
or U11484 (N_11484,N_9629,N_8904);
and U11485 (N_11485,N_8599,N_8823);
xnor U11486 (N_11486,N_8965,N_8563);
and U11487 (N_11487,N_9026,N_9494);
and U11488 (N_11488,N_9975,N_8612);
nor U11489 (N_11489,N_8681,N_9135);
nand U11490 (N_11490,N_8927,N_9224);
or U11491 (N_11491,N_8312,N_8359);
and U11492 (N_11492,N_9154,N_9182);
or U11493 (N_11493,N_8840,N_9212);
or U11494 (N_11494,N_9109,N_9546);
nor U11495 (N_11495,N_9543,N_9135);
nor U11496 (N_11496,N_8517,N_9404);
and U11497 (N_11497,N_9596,N_8852);
nor U11498 (N_11498,N_9648,N_8330);
and U11499 (N_11499,N_8789,N_9692);
nand U11500 (N_11500,N_8805,N_9506);
and U11501 (N_11501,N_9099,N_9544);
nand U11502 (N_11502,N_9434,N_8072);
nor U11503 (N_11503,N_9308,N_9379);
xor U11504 (N_11504,N_9990,N_8108);
or U11505 (N_11505,N_8584,N_9042);
or U11506 (N_11506,N_8068,N_8111);
nand U11507 (N_11507,N_9934,N_9953);
nand U11508 (N_11508,N_8109,N_9179);
xnor U11509 (N_11509,N_8542,N_9278);
and U11510 (N_11510,N_8068,N_9602);
or U11511 (N_11511,N_9351,N_9821);
xor U11512 (N_11512,N_9503,N_9054);
nand U11513 (N_11513,N_8232,N_9389);
nand U11514 (N_11514,N_9392,N_9769);
xor U11515 (N_11515,N_9268,N_9050);
and U11516 (N_11516,N_9765,N_8100);
xnor U11517 (N_11517,N_8598,N_8679);
nand U11518 (N_11518,N_9546,N_9149);
xnor U11519 (N_11519,N_9355,N_8643);
xor U11520 (N_11520,N_8480,N_9646);
or U11521 (N_11521,N_8879,N_9982);
nor U11522 (N_11522,N_8495,N_9816);
nand U11523 (N_11523,N_8077,N_9247);
nand U11524 (N_11524,N_8149,N_8827);
nand U11525 (N_11525,N_9762,N_9623);
nand U11526 (N_11526,N_9778,N_8894);
nor U11527 (N_11527,N_8181,N_8058);
and U11528 (N_11528,N_9938,N_9257);
nor U11529 (N_11529,N_8417,N_9148);
nand U11530 (N_11530,N_9245,N_8298);
or U11531 (N_11531,N_8664,N_8522);
xnor U11532 (N_11532,N_9874,N_8464);
or U11533 (N_11533,N_8151,N_8264);
nor U11534 (N_11534,N_8741,N_8470);
and U11535 (N_11535,N_9217,N_9847);
or U11536 (N_11536,N_9162,N_8106);
and U11537 (N_11537,N_9045,N_9146);
xor U11538 (N_11538,N_9023,N_9397);
nor U11539 (N_11539,N_9054,N_8227);
nand U11540 (N_11540,N_8407,N_9332);
nor U11541 (N_11541,N_8980,N_8080);
xnor U11542 (N_11542,N_8509,N_9590);
nor U11543 (N_11543,N_9050,N_8945);
nand U11544 (N_11544,N_9349,N_9315);
or U11545 (N_11545,N_9226,N_9215);
nand U11546 (N_11546,N_9005,N_8024);
nand U11547 (N_11547,N_9239,N_9987);
or U11548 (N_11548,N_8663,N_8397);
nor U11549 (N_11549,N_8155,N_8485);
xor U11550 (N_11550,N_8605,N_8851);
and U11551 (N_11551,N_9638,N_8631);
and U11552 (N_11552,N_9853,N_9949);
nand U11553 (N_11553,N_8393,N_9702);
xor U11554 (N_11554,N_9313,N_8340);
nor U11555 (N_11555,N_9168,N_9655);
nor U11556 (N_11556,N_8794,N_8045);
xor U11557 (N_11557,N_8705,N_8111);
nand U11558 (N_11558,N_9692,N_9018);
nor U11559 (N_11559,N_8338,N_9648);
nand U11560 (N_11560,N_9766,N_8583);
nor U11561 (N_11561,N_8861,N_9125);
xnor U11562 (N_11562,N_9997,N_9216);
or U11563 (N_11563,N_8857,N_8779);
and U11564 (N_11564,N_9103,N_9413);
nor U11565 (N_11565,N_8006,N_8170);
nor U11566 (N_11566,N_8891,N_9167);
xnor U11567 (N_11567,N_8148,N_8378);
nand U11568 (N_11568,N_9131,N_8827);
xor U11569 (N_11569,N_9070,N_9569);
nand U11570 (N_11570,N_9091,N_9147);
nand U11571 (N_11571,N_8827,N_8613);
or U11572 (N_11572,N_9339,N_9470);
nor U11573 (N_11573,N_8056,N_8240);
nor U11574 (N_11574,N_9662,N_8316);
or U11575 (N_11575,N_8517,N_8381);
or U11576 (N_11576,N_9442,N_9965);
xor U11577 (N_11577,N_9080,N_9319);
nor U11578 (N_11578,N_8860,N_9887);
or U11579 (N_11579,N_9312,N_8248);
or U11580 (N_11580,N_8158,N_9648);
xnor U11581 (N_11581,N_9808,N_8680);
nor U11582 (N_11582,N_9199,N_9751);
nand U11583 (N_11583,N_9194,N_9749);
nand U11584 (N_11584,N_8358,N_8664);
nand U11585 (N_11585,N_9140,N_8959);
nand U11586 (N_11586,N_8654,N_9252);
nand U11587 (N_11587,N_9747,N_8792);
or U11588 (N_11588,N_9449,N_9458);
xnor U11589 (N_11589,N_9902,N_8324);
xor U11590 (N_11590,N_8232,N_8637);
or U11591 (N_11591,N_8589,N_9614);
nand U11592 (N_11592,N_8181,N_9257);
xor U11593 (N_11593,N_9611,N_9478);
and U11594 (N_11594,N_8542,N_8238);
nor U11595 (N_11595,N_9244,N_8525);
or U11596 (N_11596,N_8033,N_9944);
or U11597 (N_11597,N_9822,N_9638);
nor U11598 (N_11598,N_9032,N_8412);
xnor U11599 (N_11599,N_9958,N_8929);
nand U11600 (N_11600,N_8910,N_8671);
nor U11601 (N_11601,N_8525,N_8041);
xnor U11602 (N_11602,N_8496,N_9878);
nor U11603 (N_11603,N_9285,N_8617);
xor U11604 (N_11604,N_9082,N_8860);
nor U11605 (N_11605,N_8047,N_9593);
nand U11606 (N_11606,N_9604,N_9387);
xnor U11607 (N_11607,N_9028,N_8298);
and U11608 (N_11608,N_9437,N_8055);
nand U11609 (N_11609,N_9700,N_8783);
or U11610 (N_11610,N_9911,N_9661);
or U11611 (N_11611,N_8849,N_8584);
nand U11612 (N_11612,N_8175,N_8395);
nor U11613 (N_11613,N_8751,N_9000);
nand U11614 (N_11614,N_8288,N_9961);
and U11615 (N_11615,N_9365,N_8800);
xnor U11616 (N_11616,N_8727,N_9379);
xor U11617 (N_11617,N_9692,N_8631);
nand U11618 (N_11618,N_9768,N_8939);
xor U11619 (N_11619,N_8184,N_9587);
and U11620 (N_11620,N_8369,N_9912);
nor U11621 (N_11621,N_9578,N_9331);
and U11622 (N_11622,N_8717,N_9112);
or U11623 (N_11623,N_9539,N_9710);
and U11624 (N_11624,N_9331,N_8169);
nand U11625 (N_11625,N_9094,N_9480);
or U11626 (N_11626,N_8699,N_8070);
xnor U11627 (N_11627,N_9447,N_9167);
nor U11628 (N_11628,N_9588,N_8330);
or U11629 (N_11629,N_8893,N_9268);
and U11630 (N_11630,N_9880,N_8780);
nand U11631 (N_11631,N_8604,N_8893);
and U11632 (N_11632,N_9693,N_9350);
xnor U11633 (N_11633,N_8701,N_8287);
nor U11634 (N_11634,N_9599,N_9721);
xnor U11635 (N_11635,N_9157,N_8357);
xor U11636 (N_11636,N_9708,N_9344);
or U11637 (N_11637,N_9165,N_9984);
nand U11638 (N_11638,N_9584,N_8648);
and U11639 (N_11639,N_8279,N_9742);
xor U11640 (N_11640,N_9331,N_8293);
nor U11641 (N_11641,N_8686,N_9044);
or U11642 (N_11642,N_8465,N_8058);
nand U11643 (N_11643,N_8532,N_9751);
xnor U11644 (N_11644,N_8388,N_8239);
xnor U11645 (N_11645,N_8611,N_9470);
nand U11646 (N_11646,N_8079,N_9855);
and U11647 (N_11647,N_9127,N_9021);
nand U11648 (N_11648,N_9766,N_9215);
nand U11649 (N_11649,N_8439,N_8127);
xor U11650 (N_11650,N_9447,N_9098);
and U11651 (N_11651,N_8432,N_9540);
xor U11652 (N_11652,N_9633,N_9693);
xnor U11653 (N_11653,N_8280,N_8808);
nor U11654 (N_11654,N_8182,N_9558);
nand U11655 (N_11655,N_8664,N_9145);
xnor U11656 (N_11656,N_9320,N_8419);
xor U11657 (N_11657,N_9985,N_9266);
or U11658 (N_11658,N_9227,N_8188);
and U11659 (N_11659,N_9536,N_8693);
nand U11660 (N_11660,N_9634,N_8041);
and U11661 (N_11661,N_8089,N_9653);
xor U11662 (N_11662,N_8411,N_8700);
or U11663 (N_11663,N_9648,N_8588);
or U11664 (N_11664,N_9596,N_9755);
nand U11665 (N_11665,N_8071,N_8576);
nor U11666 (N_11666,N_9562,N_9206);
and U11667 (N_11667,N_9190,N_8204);
nand U11668 (N_11668,N_9689,N_9443);
and U11669 (N_11669,N_9746,N_8769);
nor U11670 (N_11670,N_8562,N_9039);
or U11671 (N_11671,N_8023,N_9316);
and U11672 (N_11672,N_9182,N_8993);
or U11673 (N_11673,N_9764,N_8791);
nand U11674 (N_11674,N_9698,N_8070);
or U11675 (N_11675,N_9635,N_9928);
nor U11676 (N_11676,N_8706,N_9630);
xnor U11677 (N_11677,N_8634,N_8178);
or U11678 (N_11678,N_9965,N_8399);
nor U11679 (N_11679,N_8986,N_9205);
xnor U11680 (N_11680,N_9414,N_8402);
nand U11681 (N_11681,N_9720,N_8774);
nor U11682 (N_11682,N_9502,N_8083);
nand U11683 (N_11683,N_9655,N_8274);
nand U11684 (N_11684,N_9999,N_9766);
xnor U11685 (N_11685,N_9779,N_9681);
or U11686 (N_11686,N_9811,N_8177);
nor U11687 (N_11687,N_9772,N_8969);
or U11688 (N_11688,N_8963,N_8144);
xnor U11689 (N_11689,N_8613,N_8394);
nor U11690 (N_11690,N_8881,N_8463);
or U11691 (N_11691,N_9272,N_9131);
and U11692 (N_11692,N_9091,N_9149);
nand U11693 (N_11693,N_9867,N_8804);
xor U11694 (N_11694,N_8243,N_8612);
and U11695 (N_11695,N_9320,N_8702);
nand U11696 (N_11696,N_8621,N_9386);
xor U11697 (N_11697,N_9880,N_8028);
xnor U11698 (N_11698,N_9643,N_8334);
xnor U11699 (N_11699,N_8810,N_8929);
xnor U11700 (N_11700,N_9380,N_9236);
and U11701 (N_11701,N_9161,N_8194);
or U11702 (N_11702,N_9668,N_8573);
nor U11703 (N_11703,N_9259,N_9706);
nand U11704 (N_11704,N_9725,N_9386);
or U11705 (N_11705,N_9831,N_8421);
xor U11706 (N_11706,N_8957,N_9426);
nor U11707 (N_11707,N_9215,N_9820);
nor U11708 (N_11708,N_9894,N_9544);
nand U11709 (N_11709,N_8713,N_9135);
or U11710 (N_11710,N_8495,N_9688);
and U11711 (N_11711,N_8476,N_9346);
or U11712 (N_11712,N_9866,N_8148);
and U11713 (N_11713,N_9023,N_9084);
or U11714 (N_11714,N_8683,N_9406);
or U11715 (N_11715,N_9478,N_8218);
xor U11716 (N_11716,N_8209,N_8338);
xor U11717 (N_11717,N_8781,N_8110);
and U11718 (N_11718,N_8643,N_9025);
nand U11719 (N_11719,N_8887,N_8098);
or U11720 (N_11720,N_9447,N_9285);
and U11721 (N_11721,N_9408,N_8918);
and U11722 (N_11722,N_8735,N_9824);
xor U11723 (N_11723,N_8080,N_8968);
xnor U11724 (N_11724,N_8905,N_8560);
nand U11725 (N_11725,N_9982,N_9582);
nor U11726 (N_11726,N_8304,N_8925);
or U11727 (N_11727,N_9781,N_8528);
or U11728 (N_11728,N_9285,N_8342);
nand U11729 (N_11729,N_8905,N_8849);
nor U11730 (N_11730,N_9092,N_9100);
nor U11731 (N_11731,N_8945,N_9424);
and U11732 (N_11732,N_8796,N_8960);
or U11733 (N_11733,N_8919,N_9343);
and U11734 (N_11734,N_8943,N_9623);
xor U11735 (N_11735,N_8148,N_8735);
or U11736 (N_11736,N_8748,N_9895);
nand U11737 (N_11737,N_9538,N_9196);
or U11738 (N_11738,N_9316,N_9761);
or U11739 (N_11739,N_8477,N_8411);
nand U11740 (N_11740,N_8217,N_8053);
xnor U11741 (N_11741,N_9782,N_8592);
nand U11742 (N_11742,N_8864,N_9164);
and U11743 (N_11743,N_8278,N_8017);
or U11744 (N_11744,N_8318,N_8719);
nor U11745 (N_11745,N_9411,N_8123);
or U11746 (N_11746,N_8381,N_9833);
and U11747 (N_11747,N_9012,N_9022);
or U11748 (N_11748,N_9524,N_8672);
and U11749 (N_11749,N_9376,N_9275);
nand U11750 (N_11750,N_8283,N_9598);
nor U11751 (N_11751,N_9659,N_9663);
nand U11752 (N_11752,N_9350,N_9931);
nand U11753 (N_11753,N_8688,N_8704);
nand U11754 (N_11754,N_8803,N_9802);
or U11755 (N_11755,N_9881,N_9048);
and U11756 (N_11756,N_8570,N_9831);
or U11757 (N_11757,N_8207,N_9370);
or U11758 (N_11758,N_9304,N_8759);
nand U11759 (N_11759,N_8817,N_9437);
xnor U11760 (N_11760,N_8451,N_8580);
nand U11761 (N_11761,N_9598,N_8060);
xor U11762 (N_11762,N_8686,N_8938);
or U11763 (N_11763,N_9528,N_9112);
nand U11764 (N_11764,N_9352,N_9423);
xnor U11765 (N_11765,N_8976,N_9194);
nor U11766 (N_11766,N_9475,N_8847);
or U11767 (N_11767,N_8988,N_9924);
or U11768 (N_11768,N_9876,N_9558);
nor U11769 (N_11769,N_8582,N_8783);
or U11770 (N_11770,N_8529,N_9765);
nand U11771 (N_11771,N_9012,N_8658);
or U11772 (N_11772,N_9469,N_9101);
or U11773 (N_11773,N_8864,N_8273);
or U11774 (N_11774,N_9204,N_9769);
xnor U11775 (N_11775,N_8205,N_8916);
nor U11776 (N_11776,N_9027,N_8304);
xnor U11777 (N_11777,N_9762,N_8310);
nand U11778 (N_11778,N_8663,N_9505);
or U11779 (N_11779,N_8438,N_8006);
or U11780 (N_11780,N_9134,N_9797);
or U11781 (N_11781,N_8524,N_9016);
nand U11782 (N_11782,N_9096,N_9480);
nor U11783 (N_11783,N_9568,N_9878);
nor U11784 (N_11784,N_8107,N_8298);
and U11785 (N_11785,N_8954,N_8217);
nand U11786 (N_11786,N_8943,N_9790);
xor U11787 (N_11787,N_8462,N_9524);
xnor U11788 (N_11788,N_8228,N_8187);
nor U11789 (N_11789,N_9847,N_9984);
nor U11790 (N_11790,N_9299,N_8859);
or U11791 (N_11791,N_9667,N_8827);
nor U11792 (N_11792,N_8230,N_9423);
and U11793 (N_11793,N_9958,N_9767);
or U11794 (N_11794,N_8252,N_9888);
nor U11795 (N_11795,N_9168,N_9059);
and U11796 (N_11796,N_8257,N_9809);
nor U11797 (N_11797,N_9528,N_9580);
nand U11798 (N_11798,N_8461,N_9471);
nand U11799 (N_11799,N_8626,N_9110);
or U11800 (N_11800,N_9779,N_8159);
nand U11801 (N_11801,N_8183,N_9058);
and U11802 (N_11802,N_9170,N_8130);
xnor U11803 (N_11803,N_8200,N_8528);
nand U11804 (N_11804,N_8059,N_9661);
nor U11805 (N_11805,N_8594,N_8507);
nand U11806 (N_11806,N_8599,N_9682);
xnor U11807 (N_11807,N_8925,N_9863);
xnor U11808 (N_11808,N_9598,N_8912);
or U11809 (N_11809,N_8227,N_8442);
nor U11810 (N_11810,N_9891,N_8022);
xnor U11811 (N_11811,N_8491,N_8416);
xor U11812 (N_11812,N_9602,N_9983);
and U11813 (N_11813,N_9947,N_8657);
nor U11814 (N_11814,N_9228,N_9819);
nor U11815 (N_11815,N_9822,N_9015);
or U11816 (N_11816,N_8518,N_9894);
xnor U11817 (N_11817,N_8426,N_9602);
or U11818 (N_11818,N_8165,N_8970);
xor U11819 (N_11819,N_9896,N_8581);
xor U11820 (N_11820,N_9271,N_8882);
or U11821 (N_11821,N_9996,N_9341);
or U11822 (N_11822,N_8277,N_9936);
xor U11823 (N_11823,N_9945,N_9330);
xnor U11824 (N_11824,N_9241,N_9634);
nand U11825 (N_11825,N_8317,N_9164);
nand U11826 (N_11826,N_9755,N_8504);
and U11827 (N_11827,N_8229,N_9889);
and U11828 (N_11828,N_9981,N_8838);
or U11829 (N_11829,N_9342,N_8837);
nor U11830 (N_11830,N_9528,N_9951);
nand U11831 (N_11831,N_9629,N_8099);
nand U11832 (N_11832,N_8997,N_9810);
xor U11833 (N_11833,N_9996,N_8750);
nor U11834 (N_11834,N_9700,N_8042);
xnor U11835 (N_11835,N_9198,N_8262);
nor U11836 (N_11836,N_9981,N_9950);
and U11837 (N_11837,N_8686,N_8275);
and U11838 (N_11838,N_9769,N_8149);
nand U11839 (N_11839,N_9094,N_9261);
nand U11840 (N_11840,N_9868,N_8949);
xnor U11841 (N_11841,N_8055,N_8703);
xor U11842 (N_11842,N_9930,N_9652);
xor U11843 (N_11843,N_9738,N_8873);
and U11844 (N_11844,N_9670,N_8944);
xnor U11845 (N_11845,N_8059,N_9023);
xor U11846 (N_11846,N_8107,N_8994);
xnor U11847 (N_11847,N_9733,N_9667);
and U11848 (N_11848,N_8062,N_9919);
and U11849 (N_11849,N_8645,N_8380);
nand U11850 (N_11850,N_9334,N_8851);
or U11851 (N_11851,N_9732,N_9778);
nand U11852 (N_11852,N_9539,N_9507);
xnor U11853 (N_11853,N_9457,N_9593);
nand U11854 (N_11854,N_9588,N_9937);
xor U11855 (N_11855,N_8244,N_9288);
nand U11856 (N_11856,N_9529,N_9576);
nor U11857 (N_11857,N_8436,N_8387);
and U11858 (N_11858,N_8463,N_8916);
nand U11859 (N_11859,N_8020,N_9452);
nand U11860 (N_11860,N_8142,N_8959);
xor U11861 (N_11861,N_8717,N_9203);
and U11862 (N_11862,N_9261,N_8557);
and U11863 (N_11863,N_9601,N_9807);
nand U11864 (N_11864,N_9546,N_9439);
and U11865 (N_11865,N_9285,N_9358);
nor U11866 (N_11866,N_9073,N_9900);
or U11867 (N_11867,N_8682,N_9759);
xor U11868 (N_11868,N_9079,N_9841);
or U11869 (N_11869,N_8873,N_8627);
and U11870 (N_11870,N_9623,N_8344);
nor U11871 (N_11871,N_8137,N_9793);
nand U11872 (N_11872,N_9208,N_9680);
nor U11873 (N_11873,N_8693,N_9463);
nand U11874 (N_11874,N_8933,N_8766);
nand U11875 (N_11875,N_9014,N_8376);
and U11876 (N_11876,N_9413,N_8942);
nand U11877 (N_11877,N_9789,N_9003);
and U11878 (N_11878,N_8136,N_9877);
nor U11879 (N_11879,N_8506,N_9964);
xnor U11880 (N_11880,N_9809,N_9883);
nand U11881 (N_11881,N_8135,N_9459);
xnor U11882 (N_11882,N_9178,N_9523);
nand U11883 (N_11883,N_9633,N_8187);
or U11884 (N_11884,N_8993,N_8832);
nor U11885 (N_11885,N_8492,N_8690);
and U11886 (N_11886,N_8593,N_9136);
or U11887 (N_11887,N_8300,N_9626);
or U11888 (N_11888,N_9650,N_9107);
nor U11889 (N_11889,N_9136,N_8657);
nand U11890 (N_11890,N_9723,N_8068);
nand U11891 (N_11891,N_8160,N_9570);
nor U11892 (N_11892,N_8161,N_9541);
and U11893 (N_11893,N_8923,N_8095);
and U11894 (N_11894,N_8416,N_9224);
xor U11895 (N_11895,N_9077,N_8096);
or U11896 (N_11896,N_8494,N_9640);
nor U11897 (N_11897,N_9852,N_8852);
nor U11898 (N_11898,N_9804,N_9725);
nand U11899 (N_11899,N_8307,N_8084);
xor U11900 (N_11900,N_9315,N_8787);
nor U11901 (N_11901,N_8207,N_9545);
and U11902 (N_11902,N_9695,N_8034);
nand U11903 (N_11903,N_9127,N_8032);
xor U11904 (N_11904,N_9981,N_9686);
or U11905 (N_11905,N_8632,N_8659);
nand U11906 (N_11906,N_9874,N_8458);
or U11907 (N_11907,N_8419,N_8530);
nor U11908 (N_11908,N_9433,N_8589);
and U11909 (N_11909,N_8330,N_9769);
xor U11910 (N_11910,N_8924,N_8267);
and U11911 (N_11911,N_8485,N_9925);
xor U11912 (N_11912,N_9586,N_8703);
nand U11913 (N_11913,N_8292,N_8109);
nor U11914 (N_11914,N_8718,N_8372);
nand U11915 (N_11915,N_8638,N_8632);
and U11916 (N_11916,N_9230,N_8698);
or U11917 (N_11917,N_8396,N_9712);
xnor U11918 (N_11918,N_9059,N_9090);
nor U11919 (N_11919,N_9351,N_9108);
xnor U11920 (N_11920,N_9679,N_9924);
nor U11921 (N_11921,N_8154,N_9092);
or U11922 (N_11922,N_9420,N_8661);
or U11923 (N_11923,N_9137,N_9956);
or U11924 (N_11924,N_9701,N_8892);
xor U11925 (N_11925,N_8666,N_9119);
or U11926 (N_11926,N_9384,N_9908);
or U11927 (N_11927,N_9819,N_8896);
xor U11928 (N_11928,N_8611,N_9151);
nor U11929 (N_11929,N_8130,N_9393);
or U11930 (N_11930,N_9879,N_9035);
xnor U11931 (N_11931,N_8837,N_9119);
xnor U11932 (N_11932,N_9197,N_8815);
and U11933 (N_11933,N_9277,N_8955);
xor U11934 (N_11934,N_9876,N_9653);
and U11935 (N_11935,N_8977,N_9011);
and U11936 (N_11936,N_8250,N_8406);
xnor U11937 (N_11937,N_9490,N_9649);
or U11938 (N_11938,N_9335,N_8696);
and U11939 (N_11939,N_9332,N_9362);
nor U11940 (N_11940,N_8530,N_9924);
or U11941 (N_11941,N_9974,N_9382);
nor U11942 (N_11942,N_8424,N_9165);
nor U11943 (N_11943,N_9192,N_9923);
xnor U11944 (N_11944,N_8885,N_9038);
or U11945 (N_11945,N_8106,N_8281);
and U11946 (N_11946,N_9233,N_9212);
xor U11947 (N_11947,N_8074,N_9285);
nor U11948 (N_11948,N_8711,N_9584);
nor U11949 (N_11949,N_8894,N_8252);
nor U11950 (N_11950,N_8547,N_9328);
xor U11951 (N_11951,N_8966,N_8783);
and U11952 (N_11952,N_9069,N_9883);
xor U11953 (N_11953,N_9237,N_8628);
or U11954 (N_11954,N_9698,N_8687);
and U11955 (N_11955,N_9803,N_9710);
or U11956 (N_11956,N_9507,N_9184);
or U11957 (N_11957,N_8407,N_8249);
or U11958 (N_11958,N_9253,N_8515);
xnor U11959 (N_11959,N_9053,N_9945);
nand U11960 (N_11960,N_9145,N_9846);
nor U11961 (N_11961,N_8006,N_9863);
or U11962 (N_11962,N_8326,N_9672);
nand U11963 (N_11963,N_9092,N_8968);
or U11964 (N_11964,N_8004,N_8134);
and U11965 (N_11965,N_9743,N_9216);
nand U11966 (N_11966,N_8538,N_8285);
nand U11967 (N_11967,N_9573,N_9857);
nor U11968 (N_11968,N_9261,N_9018);
and U11969 (N_11969,N_9358,N_8366);
nor U11970 (N_11970,N_9992,N_9675);
and U11971 (N_11971,N_9087,N_9780);
nor U11972 (N_11972,N_9487,N_8498);
nand U11973 (N_11973,N_8583,N_8095);
nand U11974 (N_11974,N_9032,N_9459);
nand U11975 (N_11975,N_9267,N_9758);
or U11976 (N_11976,N_8980,N_9087);
xor U11977 (N_11977,N_8238,N_8794);
and U11978 (N_11978,N_8235,N_9362);
nor U11979 (N_11979,N_9709,N_9817);
xnor U11980 (N_11980,N_8073,N_9668);
xor U11981 (N_11981,N_9243,N_9235);
and U11982 (N_11982,N_8587,N_9269);
or U11983 (N_11983,N_8336,N_8182);
and U11984 (N_11984,N_9090,N_9666);
nor U11985 (N_11985,N_9413,N_8293);
nor U11986 (N_11986,N_9591,N_8565);
nor U11987 (N_11987,N_8693,N_8518);
and U11988 (N_11988,N_8558,N_9258);
nand U11989 (N_11989,N_9306,N_8856);
xor U11990 (N_11990,N_8127,N_9148);
nand U11991 (N_11991,N_9903,N_9262);
xnor U11992 (N_11992,N_9161,N_9224);
nand U11993 (N_11993,N_9662,N_9528);
xnor U11994 (N_11994,N_8510,N_9983);
nor U11995 (N_11995,N_8142,N_9098);
nand U11996 (N_11996,N_9883,N_9970);
xor U11997 (N_11997,N_8311,N_9635);
and U11998 (N_11998,N_8571,N_8171);
nand U11999 (N_11999,N_8263,N_8946);
and U12000 (N_12000,N_10843,N_10348);
nor U12001 (N_12001,N_11789,N_11664);
or U12002 (N_12002,N_11464,N_10753);
nand U12003 (N_12003,N_11764,N_11395);
nand U12004 (N_12004,N_10349,N_10723);
nor U12005 (N_12005,N_10690,N_10022);
and U12006 (N_12006,N_11746,N_10368);
nor U12007 (N_12007,N_11966,N_11648);
nand U12008 (N_12008,N_11305,N_10315);
nor U12009 (N_12009,N_11117,N_10018);
and U12010 (N_12010,N_11227,N_11673);
nand U12011 (N_12011,N_10037,N_10304);
or U12012 (N_12012,N_10489,N_11425);
or U12013 (N_12013,N_10780,N_11466);
and U12014 (N_12014,N_10943,N_11178);
nor U12015 (N_12015,N_11758,N_11420);
and U12016 (N_12016,N_10718,N_11377);
nor U12017 (N_12017,N_11027,N_10034);
or U12018 (N_12018,N_10934,N_11209);
xnor U12019 (N_12019,N_10076,N_11110);
nand U12020 (N_12020,N_11916,N_10777);
nor U12021 (N_12021,N_10886,N_11855);
xor U12022 (N_12022,N_11347,N_10142);
nor U12023 (N_12023,N_10906,N_11287);
and U12024 (N_12024,N_10385,N_11109);
or U12025 (N_12025,N_11546,N_10169);
xor U12026 (N_12026,N_10448,N_11279);
xor U12027 (N_12027,N_10439,N_10722);
and U12028 (N_12028,N_10631,N_11460);
nand U12029 (N_12029,N_11190,N_11358);
or U12030 (N_12030,N_10061,N_10975);
nor U12031 (N_12031,N_10774,N_11840);
xor U12032 (N_12032,N_10325,N_11261);
xor U12033 (N_12033,N_11747,N_11543);
xor U12034 (N_12034,N_11427,N_11432);
nor U12035 (N_12035,N_10426,N_11226);
or U12036 (N_12036,N_11839,N_10027);
and U12037 (N_12037,N_11353,N_10532);
or U12038 (N_12038,N_11208,N_11384);
nand U12039 (N_12039,N_11069,N_10819);
nor U12040 (N_12040,N_11875,N_11731);
or U12041 (N_12041,N_11535,N_11539);
xnor U12042 (N_12042,N_10612,N_11797);
nor U12043 (N_12043,N_10458,N_11307);
and U12044 (N_12044,N_11179,N_10566);
or U12045 (N_12045,N_10624,N_10845);
and U12046 (N_12046,N_11965,N_11807);
nor U12047 (N_12047,N_11046,N_11575);
xor U12048 (N_12048,N_11336,N_10903);
nand U12049 (N_12049,N_10860,N_11195);
or U12050 (N_12050,N_10374,N_11224);
or U12051 (N_12051,N_10643,N_10912);
nor U12052 (N_12052,N_10996,N_10447);
xnor U12053 (N_12053,N_11055,N_11578);
and U12054 (N_12054,N_11762,N_10545);
nor U12055 (N_12055,N_11104,N_11620);
or U12056 (N_12056,N_11102,N_10776);
nand U12057 (N_12057,N_10237,N_10367);
or U12058 (N_12058,N_11262,N_11035);
nand U12059 (N_12059,N_10540,N_11662);
or U12060 (N_12060,N_10987,N_10789);
xnor U12061 (N_12061,N_10883,N_10657);
and U12062 (N_12062,N_11342,N_10562);
and U12063 (N_12063,N_10381,N_11599);
nor U12064 (N_12064,N_10699,N_11145);
or U12065 (N_12065,N_11832,N_11201);
nor U12066 (N_12066,N_11130,N_11625);
nand U12067 (N_12067,N_11785,N_11008);
nand U12068 (N_12068,N_10294,N_11710);
or U12069 (N_12069,N_11865,N_10069);
xor U12070 (N_12070,N_11422,N_11619);
nor U12071 (N_12071,N_10927,N_11489);
and U12072 (N_12072,N_11142,N_10878);
nand U12073 (N_12073,N_11180,N_10415);
xnor U12074 (N_12074,N_10316,N_10354);
or U12075 (N_12075,N_10627,N_11253);
or U12076 (N_12076,N_11589,N_11565);
and U12077 (N_12077,N_11717,N_10908);
nor U12078 (N_12078,N_11940,N_10118);
nor U12079 (N_12079,N_11309,N_11094);
and U12080 (N_12080,N_10762,N_11900);
and U12081 (N_12081,N_11150,N_10885);
nor U12082 (N_12082,N_10497,N_11500);
nor U12083 (N_12083,N_11666,N_11756);
nand U12084 (N_12084,N_11729,N_10937);
or U12085 (N_12085,N_10495,N_10010);
and U12086 (N_12086,N_10500,N_10117);
nor U12087 (N_12087,N_10088,N_11860);
xor U12088 (N_12088,N_10710,N_10605);
nand U12089 (N_12089,N_10375,N_11609);
and U12090 (N_12090,N_11517,N_10477);
xor U12091 (N_12091,N_11655,N_11293);
and U12092 (N_12092,N_11853,N_10282);
or U12093 (N_12093,N_11282,N_11001);
nand U12094 (N_12094,N_11159,N_11817);
xnor U12095 (N_12095,N_10429,N_11786);
xor U12096 (N_12096,N_11868,N_10583);
and U12097 (N_12097,N_10632,N_10530);
and U12098 (N_12098,N_11448,N_10758);
or U12099 (N_12099,N_11087,N_11996);
nand U12100 (N_12100,N_10979,N_10697);
and U12101 (N_12101,N_10863,N_11158);
nand U12102 (N_12102,N_11049,N_10582);
nor U12103 (N_12103,N_11725,N_11127);
and U12104 (N_12104,N_10298,N_11401);
nand U12105 (N_12105,N_10038,N_10152);
xor U12106 (N_12106,N_11879,N_11375);
nand U12107 (N_12107,N_11041,N_11635);
or U12108 (N_12108,N_10479,N_11498);
xnor U12109 (N_12109,N_10411,N_10848);
and U12110 (N_12110,N_11140,N_10748);
and U12111 (N_12111,N_11101,N_11885);
or U12112 (N_12112,N_10097,N_11902);
nor U12113 (N_12113,N_10503,N_10330);
nor U12114 (N_12114,N_10572,N_10200);
nor U12115 (N_12115,N_10740,N_10214);
nor U12116 (N_12116,N_11289,N_11246);
nor U12117 (N_12117,N_10279,N_11769);
xnor U12118 (N_12118,N_11939,N_10935);
or U12119 (N_12119,N_11590,N_11230);
nand U12120 (N_12120,N_10311,N_10441);
nor U12121 (N_12121,N_10161,N_10916);
nor U12122 (N_12122,N_10160,N_10766);
and U12123 (N_12123,N_11311,N_10114);
xor U12124 (N_12124,N_10955,N_10059);
nor U12125 (N_12125,N_10179,N_11251);
nor U12126 (N_12126,N_10534,N_10427);
nand U12127 (N_12127,N_11737,N_11985);
or U12128 (N_12128,N_10588,N_10004);
or U12129 (N_12129,N_10666,N_10094);
nor U12130 (N_12130,N_11653,N_10194);
nand U12131 (N_12131,N_11412,N_10086);
nand U12132 (N_12132,N_11429,N_10615);
xor U12133 (N_12133,N_10983,N_10980);
nor U12134 (N_12134,N_10757,N_11438);
nand U12135 (N_12135,N_10750,N_10393);
xor U12136 (N_12136,N_11470,N_11728);
nor U12137 (N_12137,N_11125,N_11632);
and U12138 (N_12138,N_11880,N_10058);
and U12139 (N_12139,N_10767,N_10982);
nor U12140 (N_12140,N_10190,N_11273);
xor U12141 (N_12141,N_10695,N_11611);
and U12142 (N_12142,N_10444,N_11167);
xor U12143 (N_12143,N_11095,N_11318);
xnor U12144 (N_12144,N_10351,N_11556);
xnor U12145 (N_12145,N_11265,N_10029);
or U12146 (N_12146,N_10749,N_11838);
and U12147 (N_12147,N_10063,N_11415);
nor U12148 (N_12148,N_10577,N_11114);
xor U12149 (N_12149,N_10339,N_10023);
xnor U12150 (N_12150,N_11480,N_10905);
xnor U12151 (N_12151,N_10866,N_11410);
nand U12152 (N_12152,N_10981,N_11275);
nand U12153 (N_12153,N_11269,N_11942);
xor U12154 (N_12154,N_10779,N_10896);
xnor U12155 (N_12155,N_10528,N_11783);
or U12156 (N_12156,N_10678,N_10910);
and U12157 (N_12157,N_10614,N_10265);
nand U12158 (N_12158,N_11058,N_11613);
nor U12159 (N_12159,N_11630,N_10681);
and U12160 (N_12160,N_11315,N_11568);
nor U12161 (N_12161,N_10775,N_10150);
nor U12162 (N_12162,N_10842,N_10652);
xor U12163 (N_12163,N_11726,N_11695);
nand U12164 (N_12164,N_10628,N_10144);
or U12165 (N_12165,N_11544,N_10128);
nand U12166 (N_12166,N_10240,N_10801);
or U12167 (N_12167,N_10956,N_10637);
xnor U12168 (N_12168,N_10806,N_10419);
nor U12169 (N_12169,N_10388,N_11848);
nor U12170 (N_12170,N_11022,N_11426);
xnor U12171 (N_12171,N_10278,N_11514);
nor U12172 (N_12172,N_11864,N_11258);
or U12173 (N_12173,N_10920,N_11862);
or U12174 (N_12174,N_10884,N_11332);
nor U12175 (N_12175,N_11207,N_11247);
nand U12176 (N_12176,N_10317,N_10131);
nand U12177 (N_12177,N_10539,N_11782);
and U12178 (N_12178,N_11337,N_11955);
or U12179 (N_12179,N_10186,N_11435);
or U12180 (N_12180,N_11943,N_10998);
and U12181 (N_12181,N_11536,N_11937);
xor U12182 (N_12182,N_11820,N_10377);
or U12183 (N_12183,N_11692,N_11340);
and U12184 (N_12184,N_10705,N_10341);
or U12185 (N_12185,N_10591,N_11928);
or U12186 (N_12186,N_11799,N_10711);
nor U12187 (N_12187,N_11255,N_11172);
and U12188 (N_12188,N_10786,N_11971);
and U12189 (N_12189,N_10234,N_10736);
nor U12190 (N_12190,N_10424,N_11123);
and U12191 (N_12191,N_10111,N_10251);
and U12192 (N_12192,N_11161,N_10665);
nor U12193 (N_12193,N_10549,N_10850);
nor U12194 (N_12194,N_10266,N_11335);
and U12195 (N_12195,N_10033,N_11457);
or U12196 (N_12196,N_11453,N_10084);
xnor U12197 (N_12197,N_10735,N_10891);
xnor U12198 (N_12198,N_11886,N_10832);
or U12199 (N_12199,N_10554,N_11947);
nand U12200 (N_12200,N_11693,N_10276);
nor U12201 (N_12201,N_11199,N_10668);
or U12202 (N_12202,N_10536,N_10602);
nor U12203 (N_12203,N_11491,N_11750);
nor U12204 (N_12204,N_11711,N_10049);
and U12205 (N_12205,N_11948,N_11310);
nor U12206 (N_12206,N_11702,N_10133);
xnor U12207 (N_12207,N_11564,N_10918);
nand U12208 (N_12208,N_11829,N_11461);
xnor U12209 (N_12209,N_10565,N_10456);
xnor U12210 (N_12210,N_10683,N_10544);
or U12211 (N_12211,N_11152,N_11021);
nand U12212 (N_12212,N_11897,N_11134);
nor U12213 (N_12213,N_11512,N_11112);
nand U12214 (N_12214,N_11592,N_11248);
nand U12215 (N_12215,N_10202,N_10391);
xnor U12216 (N_12216,N_11739,N_11507);
nor U12217 (N_12217,N_11964,N_11346);
xnor U12218 (N_12218,N_11509,N_11588);
xnor U12219 (N_12219,N_11321,N_11014);
nor U12220 (N_12220,N_10725,N_11276);
nor U12221 (N_12221,N_11373,N_10993);
nor U12222 (N_12222,N_10679,N_11171);
nand U12223 (N_12223,N_10764,N_11793);
nand U12224 (N_12224,N_10480,N_10012);
or U12225 (N_12225,N_10106,N_10510);
xnor U12226 (N_12226,N_11534,N_10299);
or U12227 (N_12227,N_10007,N_11268);
nand U12228 (N_12228,N_11608,N_10992);
or U12229 (N_12229,N_11042,N_11944);
xnor U12230 (N_12230,N_11424,N_10809);
xor U12231 (N_12231,N_11052,N_11039);
xor U12232 (N_12232,N_10066,N_10134);
or U12233 (N_12233,N_11601,N_10384);
and U12234 (N_12234,N_10941,N_11791);
and U12235 (N_12235,N_10598,N_10292);
or U12236 (N_12236,N_10263,N_11800);
and U12237 (N_12237,N_10873,N_10702);
or U12238 (N_12238,N_10446,N_10407);
nor U12239 (N_12239,N_10387,N_11437);
nand U12240 (N_12240,N_11774,N_11122);
or U12241 (N_12241,N_10694,N_10994);
and U12242 (N_12242,N_11621,N_11249);
nor U12243 (N_12243,N_10283,N_10726);
or U12244 (N_12244,N_10345,N_11407);
nand U12245 (N_12245,N_11932,N_11124);
and U12246 (N_12246,N_11802,N_10932);
xor U12247 (N_12247,N_11175,N_11174);
xor U12248 (N_12248,N_11079,N_10470);
nor U12249 (N_12249,N_10971,N_11409);
xnor U12250 (N_12250,N_11364,N_10457);
nand U12251 (N_12251,N_10701,N_11166);
xor U12252 (N_12252,N_10921,N_11765);
nand U12253 (N_12253,N_10737,N_10019);
xnor U12254 (N_12254,N_11075,N_10636);
nor U12255 (N_12255,N_11478,N_11618);
or U12256 (N_12256,N_11736,N_11640);
or U12257 (N_12257,N_10296,N_10225);
or U12258 (N_12258,N_11149,N_10645);
xor U12259 (N_12259,N_11492,N_11983);
nand U12260 (N_12260,N_10101,N_11413);
nor U12261 (N_12261,N_10442,N_10914);
nor U12262 (N_12262,N_11675,N_10228);
xor U12263 (N_12263,N_11077,N_11417);
xnor U12264 (N_12264,N_11542,N_10693);
xor U12265 (N_12265,N_10406,N_10314);
xnor U12266 (N_12266,N_11271,N_10449);
or U12267 (N_12267,N_10923,N_10210);
or U12268 (N_12268,N_10610,N_10356);
and U12269 (N_12269,N_10744,N_11604);
xor U12270 (N_12270,N_11157,N_10287);
nand U12271 (N_12271,N_11627,N_10051);
nor U12272 (N_12272,N_10015,N_10733);
xnor U12273 (N_12273,N_10352,N_10378);
nor U12274 (N_12274,N_11560,N_11391);
xnor U12275 (N_12275,N_11936,N_10856);
nor U12276 (N_12276,N_11724,N_11007);
and U12277 (N_12277,N_11363,N_10344);
and U12278 (N_12278,N_10793,N_11020);
and U12279 (N_12279,N_11775,N_11925);
nand U12280 (N_12280,N_11892,N_11629);
and U12281 (N_12281,N_10862,N_10826);
or U12282 (N_12282,N_11354,N_10521);
nor U12283 (N_12283,N_10222,N_11091);
and U12284 (N_12284,N_11779,N_10432);
nor U12285 (N_12285,N_10574,N_11397);
or U12286 (N_12286,N_11128,N_11582);
xor U12287 (N_12287,N_11106,N_11286);
and U12288 (N_12288,N_10601,N_10464);
nand U12289 (N_12289,N_10350,N_10644);
and U12290 (N_12290,N_11994,N_10973);
nand U12291 (N_12291,N_10204,N_10274);
or U12292 (N_12292,N_10443,N_11463);
nor U12293 (N_12293,N_10014,N_10291);
and U12294 (N_12294,N_10846,N_11096);
nand U12295 (N_12295,N_10707,N_10663);
and U12296 (N_12296,N_11033,N_10492);
or U12297 (N_12297,N_10176,N_11869);
or U12298 (N_12298,N_10413,N_11844);
and U12299 (N_12299,N_10796,N_10782);
nand U12300 (N_12300,N_11953,N_11369);
nor U12301 (N_12301,N_11767,N_10229);
or U12302 (N_12302,N_11168,N_10656);
and U12303 (N_12303,N_10974,N_10110);
nor U12304 (N_12304,N_10513,N_10940);
nor U12305 (N_12305,N_11242,N_10970);
and U12306 (N_12306,N_10039,N_11245);
xnor U12307 (N_12307,N_11169,N_11277);
nand U12308 (N_12308,N_11177,N_11366);
or U12309 (N_12309,N_10535,N_10165);
nor U12310 (N_12310,N_10332,N_11532);
xnor U12311 (N_12311,N_11691,N_11283);
xnor U12312 (N_12312,N_10425,N_11189);
xnor U12313 (N_12313,N_10180,N_10095);
xor U12314 (N_12314,N_10437,N_10370);
nand U12315 (N_12315,N_10901,N_10585);
xor U12316 (N_12316,N_10512,N_10538);
nand U12317 (N_12317,N_11907,N_11383);
xnor U12318 (N_12318,N_11399,N_10136);
xor U12319 (N_12319,N_11083,N_10504);
or U12320 (N_12320,N_11144,N_10248);
nand U12321 (N_12321,N_11495,N_10396);
nand U12322 (N_12322,N_11626,N_10098);
or U12323 (N_12323,N_11525,N_10221);
nor U12324 (N_12324,N_10171,N_10831);
nand U12325 (N_12325,N_11388,N_10147);
xor U12326 (N_12326,N_11721,N_10343);
and U12327 (N_12327,N_11334,N_10999);
nand U12328 (N_12328,N_11333,N_11576);
nand U12329 (N_12329,N_10360,N_11981);
nand U12330 (N_12330,N_11993,N_11233);
or U12331 (N_12331,N_11951,N_10989);
or U12332 (N_12332,N_10765,N_11659);
xnor U12333 (N_12333,N_10103,N_11538);
or U12334 (N_12334,N_10670,N_11610);
nand U12335 (N_12335,N_10060,N_10508);
and U12336 (N_12336,N_10686,N_11098);
xor U12337 (N_12337,N_11115,N_10361);
nand U12338 (N_12338,N_11784,N_11636);
nor U12339 (N_12339,N_11408,N_10564);
and U12340 (N_12340,N_10647,N_11813);
xnor U12341 (N_12341,N_10295,N_10099);
nor U12342 (N_12342,N_10235,N_11181);
nand U12343 (N_12343,N_10042,N_11074);
or U12344 (N_12344,N_10900,N_11234);
or U12345 (N_12345,N_10719,N_10342);
and U12346 (N_12346,N_11794,N_11452);
nand U12347 (N_12347,N_11605,N_10875);
or U12348 (N_12348,N_10650,N_10195);
nor U12349 (N_12349,N_11763,N_10309);
or U12350 (N_12350,N_10919,N_11028);
or U12351 (N_12351,N_11920,N_10347);
nand U12352 (N_12352,N_10435,N_10249);
nand U12353 (N_12353,N_11024,N_10575);
or U12354 (N_12354,N_10269,N_11441);
xnor U12355 (N_12355,N_11281,N_10082);
nor U12356 (N_12356,N_11476,N_10423);
and U12357 (N_12357,N_11773,N_11066);
and U12358 (N_12358,N_11958,N_10825);
and U12359 (N_12359,N_11097,N_11136);
nor U12360 (N_12360,N_11863,N_11210);
and U12361 (N_12361,N_10984,N_11715);
nor U12362 (N_12362,N_11776,N_11531);
or U12363 (N_12363,N_10524,N_11989);
nand U12364 (N_12364,N_10728,N_10531);
xor U12365 (N_12365,N_10972,N_11393);
or U12366 (N_12366,N_10593,N_10865);
nor U12367 (N_12367,N_11694,N_10041);
or U12368 (N_12368,N_11898,N_11707);
nor U12369 (N_12369,N_10493,N_10043);
and U12370 (N_12370,N_10026,N_11639);
xor U12371 (N_12371,N_11176,N_11795);
and U12372 (N_12372,N_11946,N_10658);
xnor U12373 (N_12373,N_11557,N_10882);
nand U12374 (N_12374,N_11978,N_10902);
and U12375 (N_12375,N_10380,N_10915);
xnor U12376 (N_12376,N_11396,N_10466);
nor U12377 (N_12377,N_11467,N_11705);
xor U12378 (N_12378,N_10416,N_11871);
nor U12379 (N_12379,N_10673,N_11219);
nand U12380 (N_12380,N_11186,N_10175);
nand U12381 (N_12381,N_10810,N_11945);
nand U12382 (N_12382,N_11753,N_10199);
xor U12383 (N_12383,N_10125,N_11634);
and U12384 (N_12384,N_11792,N_10233);
and U12385 (N_12385,N_10870,N_10603);
nand U12386 (N_12386,N_11019,N_10166);
nand U12387 (N_12387,N_11043,N_10849);
nand U12388 (N_12388,N_11206,N_11191);
nand U12389 (N_12389,N_10680,N_11063);
and U12390 (N_12390,N_10818,N_10243);
xor U12391 (N_12391,N_11571,N_11780);
nand U12392 (N_12392,N_10463,N_10035);
nand U12393 (N_12393,N_10164,N_11676);
nand U12394 (N_12394,N_11003,N_11405);
nor U12395 (N_12395,N_11727,N_10067);
or U12396 (N_12396,N_10167,N_10293);
nor U12397 (N_12397,N_11644,N_11749);
nor U12398 (N_12398,N_10410,N_10484);
and U12399 (N_12399,N_11433,N_10080);
nor U12400 (N_12400,N_11320,N_10815);
xor U12401 (N_12401,N_11895,N_10720);
xnor U12402 (N_12402,N_10966,N_11845);
and U12403 (N_12403,N_11990,N_10467);
or U12404 (N_12404,N_11883,N_11714);
nor U12405 (N_12405,N_11641,N_11411);
xor U12406 (N_12406,N_10674,N_11952);
or U12407 (N_12407,N_11456,N_11600);
nor U12408 (N_12408,N_11528,N_10646);
or U12409 (N_12409,N_11672,N_10817);
xnor U12410 (N_12410,N_10820,N_10717);
xor U12411 (N_12411,N_10879,N_11006);
or U12412 (N_12412,N_11980,N_11530);
or U12413 (N_12413,N_10568,N_10253);
and U12414 (N_12414,N_11451,N_11235);
or U12415 (N_12415,N_11704,N_11935);
and U12416 (N_12416,N_10578,N_11103);
xor U12417 (N_12417,N_10091,N_10433);
nand U12418 (N_12418,N_10799,N_10145);
or U12419 (N_12419,N_11891,N_11882);
and U12420 (N_12420,N_10267,N_11482);
or U12421 (N_12421,N_11541,N_10877);
nand U12422 (N_12422,N_11645,N_11257);
nand U12423 (N_12423,N_10092,N_11593);
nand U12424 (N_12424,N_10548,N_11876);
nor U12425 (N_12425,N_10397,N_11473);
or U12426 (N_12426,N_11919,N_10157);
and U12427 (N_12427,N_11468,N_11365);
or U12428 (N_12428,N_11051,N_11893);
nor U12429 (N_12429,N_11483,N_10048);
nand U12430 (N_12430,N_10773,N_10077);
nand U12431 (N_12431,N_11830,N_11011);
xor U12432 (N_12432,N_11216,N_10430);
nand U12433 (N_12433,N_10861,N_10153);
or U12434 (N_12434,N_11558,N_10006);
nor U12435 (N_12435,N_11047,N_11595);
xor U12436 (N_12436,N_11434,N_11905);
or U12437 (N_12437,N_10949,N_11976);
xnor U12438 (N_12438,N_11402,N_11651);
or U12439 (N_12439,N_10013,N_11280);
nor U12440 (N_12440,N_11352,N_10338);
nor U12441 (N_12441,N_10068,N_10622);
nor U12442 (N_12442,N_10741,N_11836);
xnor U12443 (N_12443,N_11914,N_11044);
nand U12444 (N_12444,N_11894,N_10021);
nor U12445 (N_12445,N_10533,N_11183);
or U12446 (N_12446,N_10478,N_10995);
and U12447 (N_12447,N_10428,N_10008);
xnor U12448 (N_12448,N_11505,N_11961);
and U12449 (N_12449,N_11067,N_11445);
or U12450 (N_12450,N_10206,N_10555);
and U12451 (N_12451,N_10085,N_10151);
nor U12452 (N_12452,N_11744,N_10191);
nor U12453 (N_12453,N_10698,N_10633);
xor U12454 (N_12454,N_11968,N_10703);
or U12455 (N_12455,N_10626,N_10302);
xnor U12456 (N_12456,N_10005,N_11013);
or U12457 (N_12457,N_11995,N_11888);
and U12458 (N_12458,N_11004,N_11970);
or U12459 (N_12459,N_11959,N_10219);
and U12460 (N_12460,N_11718,N_10706);
or U12461 (N_12461,N_11585,N_11931);
or U12462 (N_12462,N_11223,N_10499);
nand U12463 (N_12463,N_10337,N_10911);
xor U12464 (N_12464,N_11072,N_11684);
and U12465 (N_12465,N_10178,N_10207);
nor U12466 (N_12466,N_11548,N_10065);
or U12467 (N_12467,N_10881,N_10813);
and U12468 (N_12468,N_10855,N_11518);
nor U12469 (N_12469,N_10149,N_10392);
nor U12470 (N_12470,N_11475,N_10840);
nand U12471 (N_12471,N_11658,N_10730);
or U12472 (N_12472,N_10032,N_10198);
and U12473 (N_12473,N_10262,N_10551);
nor U12474 (N_12474,N_11455,N_11814);
and U12475 (N_12475,N_10455,N_11062);
xor U12476 (N_12476,N_11678,N_10600);
nor U12477 (N_12477,N_10917,N_10571);
xnor U12478 (N_12478,N_11120,N_11351);
and U12479 (N_12479,N_11513,N_10496);
xnor U12480 (N_12480,N_10841,N_11740);
nand U12481 (N_12481,N_10899,N_10787);
or U12482 (N_12482,N_10215,N_11587);
or U12483 (N_12483,N_11924,N_11992);
or U12484 (N_12484,N_11225,N_10183);
and U12485 (N_12485,N_11870,N_10898);
nand U12486 (N_12486,N_10890,N_10141);
and U12487 (N_12487,N_11819,N_10682);
and U12488 (N_12488,N_11143,N_11348);
or U12489 (N_12489,N_10137,N_11584);
nor U12490 (N_12490,N_10320,N_11759);
and U12491 (N_12491,N_11573,N_10322);
or U12492 (N_12492,N_10327,N_11387);
or U12493 (N_12493,N_10258,N_11508);
nand U12494 (N_12494,N_10020,N_11849);
or U12495 (N_12495,N_10404,N_10978);
or U12496 (N_12496,N_10708,N_11722);
or U12497 (N_12497,N_10514,N_10254);
nor U12498 (N_12498,N_10727,N_10691);
xnor U12499 (N_12499,N_10520,N_11059);
or U12500 (N_12500,N_11465,N_10802);
nand U12501 (N_12501,N_10220,N_11825);
nand U12502 (N_12502,N_10724,N_10481);
and U12503 (N_12503,N_10791,N_11757);
or U12504 (N_12504,N_11679,N_11745);
and U12505 (N_12505,N_10421,N_10434);
nand U12506 (N_12506,N_10768,N_10828);
nand U12507 (N_12507,N_11766,N_11668);
nand U12508 (N_12508,N_10700,N_11867);
and U12509 (N_12509,N_11743,N_11633);
xor U12510 (N_12510,N_11126,N_10642);
or U12511 (N_12511,N_11598,N_10606);
or U12512 (N_12512,N_10071,N_11349);
and U12513 (N_12513,N_11316,N_11100);
xnor U12514 (N_12514,N_11121,N_11669);
nand U12515 (N_12515,N_11419,N_11555);
xnor U12516 (N_12516,N_11787,N_11567);
xor U12517 (N_12517,N_10651,N_10880);
or U12518 (N_12518,N_11471,N_11086);
xor U12519 (N_12519,N_11772,N_10968);
xor U12520 (N_12520,N_11856,N_11156);
or U12521 (N_12521,N_10121,N_10326);
nor U12522 (N_12522,N_11918,N_11547);
nand U12523 (N_12523,N_10963,N_10162);
or U12524 (N_12524,N_11654,N_11973);
and U12525 (N_12525,N_10123,N_11663);
xor U12526 (N_12526,N_10055,N_10864);
xnor U12527 (N_12527,N_11030,N_11141);
xor U12528 (N_12528,N_11972,N_11846);
and U12529 (N_12529,N_10420,N_11360);
and U12530 (N_12530,N_11606,N_11322);
or U12531 (N_12531,N_10155,N_10382);
and U12532 (N_12532,N_11416,N_10759);
or U12533 (N_12533,N_10851,N_11295);
nand U12534 (N_12534,N_10662,N_10868);
nand U12535 (N_12535,N_10129,N_10648);
or U12536 (N_12536,N_10579,N_11355);
nor U12537 (N_12537,N_11515,N_10261);
nand U12538 (N_12538,N_11237,N_11760);
and U12539 (N_12539,N_10743,N_10729);
or U12540 (N_12540,N_10445,N_10053);
and U12541 (N_12541,N_11550,N_10372);
nor U12542 (N_12542,N_10239,N_11956);
xnor U12543 (N_12543,N_10188,N_11828);
nor U12544 (N_12544,N_10140,N_11447);
nand U12545 (N_12545,N_11708,N_11977);
and U12546 (N_12546,N_11449,N_10189);
nor U12547 (N_12547,N_10894,N_10784);
xnor U12548 (N_12548,N_11960,N_10364);
nor U12549 (N_12549,N_11496,N_11071);
and U12550 (N_12550,N_10509,N_11450);
xor U12551 (N_12551,N_11080,N_10218);
and U12552 (N_12552,N_10550,N_10769);
xor U12553 (N_12553,N_11572,N_10079);
xnor U12554 (N_12554,N_10224,N_10529);
xnor U12555 (N_12555,N_11023,N_10816);
or U12556 (N_12556,N_10135,N_11327);
xnor U12557 (N_12557,N_10552,N_11000);
or U12558 (N_12558,N_11537,N_10839);
or U12559 (N_12559,N_10057,N_10822);
and U12560 (N_12560,N_11881,N_10389);
nor U12561 (N_12561,N_11154,N_10259);
and U12562 (N_12562,N_11479,N_11801);
xor U12563 (N_12563,N_10398,N_10526);
nor U12564 (N_12564,N_11921,N_10515);
nand U12565 (N_12565,N_10611,N_11038);
xnor U12566 (N_12566,N_10373,N_10704);
or U12567 (N_12567,N_10939,N_11697);
nand U12568 (N_12568,N_10976,N_10830);
nand U12569 (N_12569,N_10286,N_10379);
and U12570 (N_12570,N_10072,N_10472);
nand U12571 (N_12571,N_11328,N_10560);
and U12572 (N_12572,N_11809,N_11371);
xor U12573 (N_12573,N_10469,N_11957);
and U12574 (N_12574,N_11719,N_10738);
and U12575 (N_12575,N_10542,N_10277);
xor U12576 (N_12576,N_11815,N_10944);
nor U12577 (N_12577,N_11529,N_10607);
or U12578 (N_12578,N_10000,N_11188);
or U12579 (N_12579,N_10096,N_11222);
xnor U12580 (N_12580,N_10438,N_10867);
and U12581 (N_12581,N_10561,N_11398);
nand U12582 (N_12582,N_11341,N_10567);
xor U12583 (N_12583,N_11665,N_10002);
nand U12584 (N_12584,N_10771,N_10025);
xor U12585 (N_12585,N_11442,N_10482);
nand U12586 (N_12586,N_11070,N_11788);
or U12587 (N_12587,N_11562,N_11054);
nor U12588 (N_12588,N_11696,N_11381);
nor U12589 (N_12589,N_11804,N_10328);
xor U12590 (N_12590,N_10359,N_11812);
nand U12591 (N_12591,N_10604,N_11748);
nand U12592 (N_12592,N_10838,N_10197);
nand U12593 (N_12593,N_10897,N_11701);
and U12594 (N_12594,N_11490,N_10146);
or U12595 (N_12595,N_10331,N_10203);
or U12596 (N_12596,N_10403,N_11771);
nand U12597 (N_12597,N_10300,N_10412);
or U12598 (N_12598,N_10924,N_10358);
or U12599 (N_12599,N_11581,N_10461);
nand U12600 (N_12600,N_11263,N_11612);
and U12601 (N_12601,N_11854,N_11709);
xnor U12602 (N_12602,N_11314,N_11912);
nor U12603 (N_12603,N_11526,N_10310);
nand U12604 (N_12604,N_10709,N_11139);
xor U12605 (N_12605,N_11284,N_11085);
or U12606 (N_12606,N_11768,N_10772);
and U12607 (N_12607,N_10355,N_10115);
or U12608 (N_12608,N_11833,N_11643);
or U12609 (N_12609,N_10193,N_11484);
or U12610 (N_12610,N_11851,N_11850);
and U12611 (N_12611,N_11076,N_10127);
nand U12612 (N_12612,N_10742,N_10516);
or U12613 (N_12613,N_11504,N_10790);
nand U12614 (N_12614,N_10511,N_10858);
nand U12615 (N_12615,N_10618,N_11950);
nand U12616 (N_12616,N_10307,N_10132);
xor U12617 (N_12617,N_11217,N_10454);
nor U12618 (N_12618,N_11974,N_11382);
nor U12619 (N_12619,N_10671,N_11738);
nor U12620 (N_12620,N_11842,N_10045);
and U12621 (N_12621,N_11204,N_10570);
and U12622 (N_12622,N_10460,N_11908);
and U12623 (N_12623,N_10090,N_11138);
xor U12624 (N_12624,N_10785,N_11674);
or U12625 (N_12625,N_10363,N_11323);
or U12626 (N_12626,N_10313,N_11133);
nor U12627 (N_12627,N_10369,N_10609);
nand U12628 (N_12628,N_11198,N_10599);
xnor U12629 (N_12629,N_11847,N_10431);
nor U12630 (N_12630,N_11680,N_11624);
xor U12631 (N_12631,N_10659,N_10946);
nor U12632 (N_12632,N_10245,N_11390);
xor U12633 (N_12633,N_10957,N_10948);
and U12634 (N_12634,N_11808,N_11155);
and U12635 (N_12635,N_10319,N_11212);
xor U12636 (N_12636,N_11521,N_11681);
nor U12637 (N_12637,N_11927,N_11660);
and U12638 (N_12638,N_11754,N_10172);
nand U12639 (N_12639,N_10256,N_11324);
xnor U12640 (N_12640,N_10953,N_10547);
and U12641 (N_12641,N_10230,N_11615);
and U12642 (N_12642,N_11093,N_10223);
and U12643 (N_12643,N_11887,N_10073);
or U12644 (N_12644,N_11304,N_11229);
nand U12645 (N_12645,N_11687,N_10408);
and U12646 (N_12646,N_10312,N_11215);
or U12647 (N_12647,N_10409,N_10046);
or U12648 (N_12648,N_11690,N_11999);
nor U12649 (N_12649,N_10712,N_11319);
nor U12650 (N_12650,N_11469,N_11646);
nand U12651 (N_12651,N_10505,N_11200);
nand U12652 (N_12652,N_10143,N_10062);
xor U12653 (N_12653,N_10272,N_10158);
xnor U12654 (N_12654,N_10543,N_11010);
and U12655 (N_12655,N_11065,N_11026);
xnor U12656 (N_12656,N_10405,N_10664);
nand U12657 (N_12657,N_11137,N_10483);
or U12658 (N_12658,N_11583,N_10933);
nor U12659 (N_12659,N_10625,N_11594);
nor U12660 (N_12660,N_11841,N_10244);
and U12661 (N_12661,N_10044,N_11078);
nand U12662 (N_12662,N_10620,N_11474);
nor U12663 (N_12663,N_10336,N_10205);
or U12664 (N_12664,N_11523,N_10093);
nor U12665 (N_12665,N_10402,N_10211);
nand U12666 (N_12666,N_10807,N_10187);
or U12667 (N_12667,N_11308,N_11913);
nand U12668 (N_12668,N_10485,N_11511);
and U12669 (N_12669,N_10945,N_10788);
nor U12670 (N_12670,N_11803,N_10714);
or U12671 (N_12671,N_11359,N_11081);
and U12672 (N_12672,N_10333,N_11628);
or U12673 (N_12673,N_10792,N_10490);
nor U12674 (N_12674,N_10696,N_11540);
nand U12675 (N_12675,N_11911,N_11938);
and U12676 (N_12676,N_11256,N_10926);
nor U12677 (N_12677,N_10623,N_10488);
or U12678 (N_12678,N_11732,N_11376);
and U12679 (N_12679,N_11053,N_10986);
and U12680 (N_12680,N_10024,N_10453);
and U12681 (N_12681,N_11713,N_10054);
and U12682 (N_12682,N_11826,N_10231);
xnor U12683 (N_12683,N_10522,N_10306);
or U12684 (N_12684,N_10030,N_10685);
nor U12685 (N_12685,N_11250,N_10653);
nand U12686 (N_12686,N_10318,N_10836);
xnor U12687 (N_12687,N_11811,N_11683);
nand U12688 (N_12688,N_10321,N_10834);
nand U12689 (N_12689,N_11221,N_11356);
nand U12690 (N_12690,N_11821,N_11616);
nand U12691 (N_12691,N_11462,N_10105);
nor U12692 (N_12692,N_11031,N_10334);
nor U12693 (N_12693,N_10227,N_10452);
nand U12694 (N_12694,N_11165,N_11487);
xor U12695 (N_12695,N_11147,N_11494);
or U12696 (N_12696,N_10163,N_11901);
nand U12697 (N_12697,N_11874,N_10487);
or U12698 (N_12698,N_11481,N_11670);
xor U12699 (N_12699,N_11073,N_10553);
or U12700 (N_12700,N_11761,N_10078);
and U12701 (N_12701,N_11278,N_11712);
nor U12702 (N_12702,N_10289,N_10357);
nor U12703 (N_12703,N_10675,N_11264);
and U12704 (N_12704,N_10346,N_11423);
or U12705 (N_12705,N_11056,N_10386);
or U12706 (N_12706,N_11671,N_11299);
nor U12707 (N_12707,N_11119,N_11566);
nand U12708 (N_12708,N_11686,N_10783);
xor U12709 (N_12709,N_11338,N_11859);
xnor U12710 (N_12710,N_10009,N_11822);
xor U12711 (N_12711,N_10216,N_10473);
or U12712 (N_12712,N_11443,N_10518);
nor U12713 (N_12713,N_10541,N_10692);
and U12714 (N_12714,N_11151,N_10506);
xnor U12715 (N_12715,N_10246,N_11372);
nand U12716 (N_12716,N_10931,N_10854);
or U12717 (N_12717,N_10936,N_10112);
nand U12718 (N_12718,N_10770,N_10122);
nor U12719 (N_12719,N_10573,N_10661);
and U12720 (N_12720,N_10688,N_11400);
xnor U12721 (N_12721,N_11113,N_10011);
nor U12722 (N_12722,N_11752,N_11503);
xor U12723 (N_12723,N_11781,N_10303);
and U12724 (N_12724,N_10803,N_11446);
nor U12725 (N_12725,N_10997,N_10590);
and U12726 (N_12726,N_11910,N_11904);
xor U12727 (N_12727,N_10950,N_11755);
nand U12728 (N_12728,N_11975,N_10595);
nor U12729 (N_12729,N_11404,N_10148);
or U12730 (N_12730,N_11406,N_10264);
or U12731 (N_12731,N_11906,N_11330);
nand U12732 (N_12732,N_11915,N_10958);
and U12733 (N_12733,N_11300,N_11368);
or U12734 (N_12734,N_10250,N_11831);
nand U12735 (N_12735,N_10558,N_11638);
xnor U12736 (N_12736,N_11267,N_10462);
nand U12737 (N_12737,N_11131,N_10752);
nor U12738 (N_12738,N_10847,N_10938);
or U12739 (N_12739,N_11602,N_10798);
and U12740 (N_12740,N_11184,N_10763);
nor U12741 (N_12741,N_11969,N_10113);
xor U12742 (N_12742,N_11477,N_10281);
nand U12743 (N_12743,N_11213,N_10174);
nand U12744 (N_12744,N_10667,N_10965);
or U12745 (N_12745,N_11431,N_10108);
nor U12746 (N_12746,N_10829,N_10734);
nor U12747 (N_12747,N_11667,N_10507);
nand U12748 (N_12748,N_11533,N_11649);
nor U12749 (N_12749,N_11259,N_10465);
xnor U12750 (N_12750,N_11301,N_10892);
and U12751 (N_12751,N_11703,N_10761);
xnor U12752 (N_12752,N_11734,N_11984);
and U12753 (N_12753,N_10468,N_10959);
nand U12754 (N_12754,N_10960,N_10498);
or U12755 (N_12755,N_11878,N_11012);
and U12756 (N_12756,N_11933,N_11962);
xnor U12757 (N_12757,N_10977,N_11770);
nor U12758 (N_12758,N_10275,N_11266);
or U12759 (N_12759,N_10857,N_11285);
and U12760 (N_12760,N_11890,N_11506);
nor U12761 (N_12761,N_11326,N_11650);
and U12762 (N_12762,N_10592,N_11563);
or U12763 (N_12763,N_10040,N_10217);
or U12764 (N_12764,N_11088,N_11561);
nor U12765 (N_12765,N_11459,N_11294);
xor U12766 (N_12766,N_10621,N_10089);
nor U12767 (N_12767,N_11378,N_11034);
and U12768 (N_12768,N_10754,N_11923);
xor U12769 (N_12769,N_10436,N_10888);
nand U12770 (N_12770,N_11877,N_11105);
nand U12771 (N_12771,N_10260,N_11231);
nor U12772 (N_12772,N_11025,N_10001);
or U12773 (N_12773,N_10800,N_11810);
xor U12774 (N_12774,N_11723,N_11861);
xor U12775 (N_12775,N_10241,N_11930);
or U12776 (N_12776,N_11274,N_10301);
or U12777 (N_12777,N_11045,N_11068);
or U12778 (N_12778,N_10399,N_11577);
nand U12779 (N_12779,N_11260,N_10247);
xor U12780 (N_12780,N_11843,N_11163);
xnor U12781 (N_12781,N_10546,N_11552);
nand U12782 (N_12782,N_10739,N_10654);
and U12783 (N_12783,N_11084,N_11818);
nor U12784 (N_12784,N_11241,N_10185);
xor U12785 (N_12785,N_11032,N_11889);
nor U12786 (N_12786,N_11949,N_11806);
xor U12787 (N_12787,N_10804,N_10104);
xnor U12788 (N_12788,N_10951,N_10721);
nor U12789 (N_12789,N_11858,N_10942);
xnor U12790 (N_12790,N_10569,N_11357);
and U12791 (N_12791,N_10794,N_10440);
xor U12792 (N_12792,N_10284,N_11343);
and U12793 (N_12793,N_11834,N_11185);
and U12794 (N_12794,N_11607,N_10676);
nand U12795 (N_12795,N_10471,N_11436);
or U12796 (N_12796,N_10797,N_11689);
nand U12797 (N_12797,N_11380,N_10871);
or U12798 (N_12798,N_10922,N_11685);
or U12799 (N_12799,N_10576,N_11997);
or U12800 (N_12800,N_11720,N_10589);
nand U12801 (N_12801,N_10003,N_10451);
or U12802 (N_12802,N_11485,N_11586);
or U12803 (N_12803,N_11545,N_10559);
nand U12804 (N_12804,N_10476,N_10760);
or U12805 (N_12805,N_10689,N_11614);
or U12806 (N_12806,N_11472,N_10329);
nand U12807 (N_12807,N_11370,N_11292);
or U12808 (N_12808,N_10597,N_11187);
nand U12809 (N_12809,N_10212,N_10811);
nor U12810 (N_12810,N_11270,N_11306);
or U12811 (N_12811,N_11118,N_10418);
or U12812 (N_12812,N_11929,N_11192);
nor U12813 (N_12813,N_11700,N_11297);
and U12814 (N_12814,N_11519,N_11580);
xnor U12815 (N_12815,N_11884,N_10844);
nand U12816 (N_12816,N_10201,N_11656);
nand U12817 (N_12817,N_10308,N_11497);
or U12818 (N_12818,N_10017,N_10168);
nor U12819 (N_12819,N_10952,N_11569);
xnor U12820 (N_12820,N_10833,N_11116);
and U12821 (N_12821,N_10616,N_11735);
nor U12822 (N_12822,N_10859,N_11403);
xnor U12823 (N_12823,N_10365,N_10124);
xnor U12824 (N_12824,N_11232,N_10109);
and U12825 (N_12825,N_11244,N_10119);
and U12826 (N_12826,N_11029,N_11524);
and U12827 (N_12827,N_11164,N_10102);
xor U12828 (N_12828,N_11903,N_10638);
xor U12829 (N_12829,N_10297,N_10395);
xnor U12830 (N_12830,N_11657,N_10120);
and U12831 (N_12831,N_11389,N_10893);
xnor U12832 (N_12832,N_11228,N_10414);
nor U12833 (N_12833,N_11182,N_11196);
nand U12834 (N_12834,N_11899,N_10967);
xnor U12835 (N_12835,N_11254,N_10517);
and U12836 (N_12836,N_11173,N_10138);
xor U12837 (N_12837,N_10954,N_10837);
nor U12838 (N_12838,N_11967,N_10047);
and U12839 (N_12839,N_10422,N_10629);
or U12840 (N_12840,N_10236,N_10641);
and U12841 (N_12841,N_11998,N_10081);
xor U12842 (N_12842,N_11016,N_11873);
nand U12843 (N_12843,N_10087,N_10181);
nand U12844 (N_12844,N_11963,N_10170);
nor U12845 (N_12845,N_10288,N_11385);
and U12846 (N_12846,N_10745,N_11979);
nor U12847 (N_12847,N_10580,N_10417);
nand U12848 (N_12848,N_10961,N_11428);
nor U12849 (N_12849,N_11742,N_11288);
xnor U12850 (N_12850,N_10985,N_10812);
and U12851 (N_12851,N_10824,N_11730);
nor U12852 (N_12852,N_11991,N_10581);
nand U12853 (N_12853,N_11510,N_11617);
nor U12854 (N_12854,N_10713,N_11502);
nor U12855 (N_12855,N_11805,N_10756);
or U12856 (N_12856,N_11239,N_10630);
nor U12857 (N_12857,N_10887,N_11089);
or U12858 (N_12858,N_11922,N_11345);
and U12859 (N_12859,N_10677,N_10556);
xnor U12860 (N_12860,N_11061,N_11699);
nand U12861 (N_12861,N_11238,N_11677);
nor U12862 (N_12862,N_11444,N_10557);
nand U12863 (N_12863,N_10687,N_10486);
nor U12864 (N_12864,N_10527,N_10028);
or U12865 (N_12865,N_11559,N_11272);
nand U12866 (N_12866,N_11367,N_11099);
and U12867 (N_12867,N_10177,N_11303);
and U12868 (N_12868,N_10192,N_11499);
xnor U12869 (N_12869,N_10182,N_10889);
xnor U12870 (N_12870,N_10525,N_10853);
xnor U12871 (N_12871,N_11623,N_10660);
xnor U12872 (N_12872,N_10684,N_11252);
xor U12873 (N_12873,N_10947,N_11092);
nor U12874 (N_12874,N_11778,N_11193);
or U12875 (N_12875,N_11486,N_10990);
xnor U12876 (N_12876,N_10991,N_11866);
or U12877 (N_12877,N_11362,N_10126);
xnor U12878 (N_12878,N_10383,N_11982);
nor U12879 (N_12879,N_10587,N_11597);
nor U12880 (N_12880,N_11009,N_10586);
nand U12881 (N_12881,N_10617,N_11374);
or U12882 (N_12882,N_11203,N_10613);
or U12883 (N_12883,N_10340,N_10751);
nor U12884 (N_12884,N_11934,N_10909);
or U12885 (N_12885,N_10805,N_10390);
or U12886 (N_12886,N_10929,N_11160);
and U12887 (N_12887,N_11111,N_11135);
and U12888 (N_12888,N_11146,N_11603);
nor U12889 (N_12889,N_11941,N_10226);
nand U12890 (N_12890,N_11458,N_10285);
nand U12891 (N_12891,N_10156,N_11835);
nand U12892 (N_12892,N_10872,N_11339);
or U12893 (N_12893,N_11796,N_10502);
nand U12894 (N_12894,N_10808,N_10962);
nor U12895 (N_12895,N_10778,N_11170);
and U12896 (N_12896,N_11211,N_10394);
nor U12897 (N_12897,N_11002,N_11108);
nor U12898 (N_12898,N_10074,N_10116);
nand U12899 (N_12899,N_11148,N_11236);
or U12900 (N_12900,N_10459,N_10672);
nor U12901 (N_12901,N_11516,N_11090);
nor U12902 (N_12902,N_11777,N_10083);
nor U12903 (N_12903,N_11050,N_11872);
nand U12904 (N_12904,N_11790,N_10634);
and U12905 (N_12905,N_11909,N_10852);
xnor U12906 (N_12906,N_11197,N_10746);
and U12907 (N_12907,N_11688,N_10130);
xnor U12908 (N_12908,N_11954,N_11647);
xnor U12909 (N_12909,N_11852,N_10257);
or U12910 (N_12910,N_10640,N_10290);
xor U12911 (N_12911,N_10070,N_10252);
nand U12912 (N_12912,N_11394,N_10064);
or U12913 (N_12913,N_11733,N_10731);
and U12914 (N_12914,N_10052,N_10715);
nand U12915 (N_12915,N_11418,N_10649);
nand U12916 (N_12916,N_10173,N_11917);
or U12917 (N_12917,N_10474,N_10619);
or U12918 (N_12918,N_11857,N_10494);
nor U12919 (N_12919,N_10716,N_10904);
nor U12920 (N_12920,N_11652,N_10376);
and U12921 (N_12921,N_10242,N_10747);
nor U12922 (N_12922,N_10523,N_11060);
nor U12923 (N_12923,N_11005,N_11243);
nor U12924 (N_12924,N_11816,N_11291);
xnor U12925 (N_12925,N_10669,N_10491);
and U12926 (N_12926,N_11386,N_11240);
xnor U12927 (N_12927,N_11214,N_11827);
xor U12928 (N_12928,N_10056,N_10400);
or U12929 (N_12929,N_10501,N_11574);
xnor U12930 (N_12930,N_11716,N_11329);
nor U12931 (N_12931,N_11986,N_10139);
and U12932 (N_12932,N_10869,N_10608);
and U12933 (N_12933,N_10323,N_10635);
xnor U12934 (N_12934,N_10075,N_10655);
or U12935 (N_12935,N_11312,N_10969);
nor U12936 (N_12936,N_11549,N_10874);
xor U12937 (N_12937,N_11824,N_11325);
nand U12938 (N_12938,N_10100,N_11896);
or U12939 (N_12939,N_10305,N_11162);
xnor U12940 (N_12940,N_10821,N_11064);
nor U12941 (N_12941,N_10988,N_11132);
nand U12942 (N_12942,N_11661,N_11344);
nor U12943 (N_12943,N_11591,N_11798);
and U12944 (N_12944,N_11302,N_11823);
nor U12945 (N_12945,N_10232,N_11202);
or U12946 (N_12946,N_11596,N_10827);
or U12947 (N_12947,N_10401,N_11218);
nor U12948 (N_12948,N_11082,N_11493);
xnor U12949 (N_12949,N_10876,N_11205);
or U12950 (N_12950,N_10184,N_10036);
and U12951 (N_12951,N_10154,N_11642);
nand U12952 (N_12952,N_11036,N_11751);
xor U12953 (N_12953,N_10270,N_10209);
nand U12954 (N_12954,N_11554,N_10273);
xnor U12955 (N_12955,N_11622,N_11579);
or U12956 (N_12956,N_11698,N_10519);
nor U12957 (N_12957,N_10324,N_11057);
or U12958 (N_12958,N_11926,N_10814);
nor U12959 (N_12959,N_10964,N_11350);
nand U12960 (N_12960,N_11421,N_11331);
or U12961 (N_12961,N_10639,N_11392);
nand U12962 (N_12962,N_10930,N_11015);
and U12963 (N_12963,N_11522,N_11040);
nor U12964 (N_12964,N_10255,N_11631);
nand U12965 (N_12965,N_10781,N_10475);
and U12966 (N_12966,N_11313,N_10213);
xnor U12967 (N_12967,N_11527,N_11018);
or U12968 (N_12968,N_10371,N_10755);
nand U12969 (N_12969,N_10107,N_11637);
nor U12970 (N_12970,N_11987,N_10584);
nor U12971 (N_12971,N_11317,N_10913);
or U12972 (N_12972,N_11194,N_11153);
xnor U12973 (N_12973,N_10835,N_11454);
nand U12974 (N_12974,N_10795,N_11553);
nor U12975 (N_12975,N_11048,N_11520);
or U12976 (N_12976,N_10594,N_10362);
or U12977 (N_12977,N_11706,N_10280);
or U12978 (N_12978,N_10159,N_11439);
and U12979 (N_12979,N_11837,N_10335);
or U12980 (N_12980,N_10238,N_10925);
nor U12981 (N_12981,N_10450,N_11296);
and U12982 (N_12982,N_11488,N_11107);
or U12983 (N_12983,N_10050,N_11298);
and U12984 (N_12984,N_10596,N_11017);
and U12985 (N_12985,N_10271,N_11501);
nand U12986 (N_12986,N_11570,N_11741);
xnor U12987 (N_12987,N_10895,N_10353);
nor U12988 (N_12988,N_10563,N_10732);
nor U12989 (N_12989,N_10537,N_10016);
nor U12990 (N_12990,N_10366,N_10196);
xor U12991 (N_12991,N_11290,N_10907);
or U12992 (N_12992,N_10928,N_11682);
xnor U12993 (N_12993,N_11379,N_10823);
and U12994 (N_12994,N_11361,N_11037);
or U12995 (N_12995,N_11551,N_11414);
nand U12996 (N_12996,N_10208,N_11129);
or U12997 (N_12997,N_11430,N_11440);
or U12998 (N_12998,N_10031,N_10268);
and U12999 (N_12999,N_11220,N_11988);
or U13000 (N_13000,N_11290,N_11011);
xor U13001 (N_13001,N_10893,N_10319);
or U13002 (N_13002,N_10557,N_10201);
and U13003 (N_13003,N_10049,N_10775);
or U13004 (N_13004,N_10017,N_10704);
xor U13005 (N_13005,N_11938,N_10441);
or U13006 (N_13006,N_10986,N_11049);
nand U13007 (N_13007,N_11405,N_11410);
nor U13008 (N_13008,N_11099,N_10583);
nor U13009 (N_13009,N_10059,N_10068);
and U13010 (N_13010,N_10159,N_11502);
and U13011 (N_13011,N_11363,N_11868);
nor U13012 (N_13012,N_11510,N_10346);
and U13013 (N_13013,N_11955,N_11636);
nor U13014 (N_13014,N_11392,N_11194);
and U13015 (N_13015,N_11294,N_10668);
nor U13016 (N_13016,N_11758,N_11928);
xor U13017 (N_13017,N_10024,N_11524);
and U13018 (N_13018,N_10373,N_11762);
or U13019 (N_13019,N_10471,N_11452);
or U13020 (N_13020,N_11172,N_11178);
nor U13021 (N_13021,N_11656,N_11746);
or U13022 (N_13022,N_10878,N_10309);
nand U13023 (N_13023,N_11364,N_11564);
and U13024 (N_13024,N_11059,N_11151);
nand U13025 (N_13025,N_10478,N_11763);
and U13026 (N_13026,N_10887,N_11909);
nand U13027 (N_13027,N_10598,N_10961);
and U13028 (N_13028,N_11800,N_11146);
or U13029 (N_13029,N_11854,N_11899);
and U13030 (N_13030,N_10861,N_11372);
nand U13031 (N_13031,N_11418,N_10173);
nand U13032 (N_13032,N_10705,N_10454);
xor U13033 (N_13033,N_11221,N_10127);
or U13034 (N_13034,N_10172,N_11934);
or U13035 (N_13035,N_11583,N_10692);
or U13036 (N_13036,N_11962,N_10566);
nand U13037 (N_13037,N_10005,N_10407);
and U13038 (N_13038,N_10925,N_10004);
nor U13039 (N_13039,N_11315,N_11274);
or U13040 (N_13040,N_10358,N_10350);
nand U13041 (N_13041,N_10730,N_10735);
or U13042 (N_13042,N_11075,N_11555);
nor U13043 (N_13043,N_11004,N_10234);
nand U13044 (N_13044,N_11105,N_11917);
and U13045 (N_13045,N_11392,N_10081);
and U13046 (N_13046,N_11452,N_11349);
nand U13047 (N_13047,N_10621,N_10288);
xnor U13048 (N_13048,N_11970,N_11060);
nor U13049 (N_13049,N_11668,N_11048);
or U13050 (N_13050,N_11289,N_10532);
nor U13051 (N_13051,N_11646,N_10696);
nor U13052 (N_13052,N_10362,N_10592);
nor U13053 (N_13053,N_11632,N_10523);
nand U13054 (N_13054,N_10492,N_11773);
or U13055 (N_13055,N_10944,N_11069);
and U13056 (N_13056,N_10884,N_10167);
and U13057 (N_13057,N_10048,N_10126);
and U13058 (N_13058,N_10246,N_10680);
xnor U13059 (N_13059,N_11234,N_10330);
nor U13060 (N_13060,N_11965,N_11441);
and U13061 (N_13061,N_10785,N_10986);
and U13062 (N_13062,N_11904,N_11562);
nor U13063 (N_13063,N_10734,N_10145);
nand U13064 (N_13064,N_11957,N_11490);
or U13065 (N_13065,N_10533,N_11120);
or U13066 (N_13066,N_10839,N_10247);
xnor U13067 (N_13067,N_10951,N_10654);
or U13068 (N_13068,N_10106,N_10530);
and U13069 (N_13069,N_11560,N_10613);
and U13070 (N_13070,N_10054,N_11799);
or U13071 (N_13071,N_11614,N_11713);
nor U13072 (N_13072,N_11238,N_11161);
and U13073 (N_13073,N_11605,N_11061);
nand U13074 (N_13074,N_11262,N_10570);
nand U13075 (N_13075,N_10123,N_11155);
and U13076 (N_13076,N_10443,N_11979);
nand U13077 (N_13077,N_10487,N_10270);
and U13078 (N_13078,N_10279,N_10009);
nor U13079 (N_13079,N_10245,N_11364);
nand U13080 (N_13080,N_10143,N_10126);
nor U13081 (N_13081,N_10504,N_11252);
xor U13082 (N_13082,N_10772,N_11633);
nand U13083 (N_13083,N_11044,N_11120);
nor U13084 (N_13084,N_10542,N_11565);
nor U13085 (N_13085,N_10246,N_11024);
nand U13086 (N_13086,N_11652,N_11411);
nor U13087 (N_13087,N_10967,N_11750);
xnor U13088 (N_13088,N_10908,N_10749);
xnor U13089 (N_13089,N_10535,N_11472);
and U13090 (N_13090,N_10717,N_11465);
nand U13091 (N_13091,N_11982,N_11943);
or U13092 (N_13092,N_11156,N_10388);
and U13093 (N_13093,N_10877,N_10225);
nand U13094 (N_13094,N_11458,N_10513);
or U13095 (N_13095,N_11207,N_10886);
xnor U13096 (N_13096,N_10408,N_11750);
nand U13097 (N_13097,N_10707,N_10749);
nand U13098 (N_13098,N_10111,N_10887);
or U13099 (N_13099,N_10946,N_11156);
xor U13100 (N_13100,N_11910,N_11528);
nor U13101 (N_13101,N_10599,N_11044);
and U13102 (N_13102,N_10052,N_10502);
xnor U13103 (N_13103,N_11995,N_10243);
or U13104 (N_13104,N_10902,N_10527);
nand U13105 (N_13105,N_11865,N_11170);
nand U13106 (N_13106,N_11098,N_10632);
xor U13107 (N_13107,N_10505,N_11332);
nand U13108 (N_13108,N_11262,N_11755);
or U13109 (N_13109,N_10190,N_11567);
and U13110 (N_13110,N_10419,N_10563);
nor U13111 (N_13111,N_10773,N_10672);
nand U13112 (N_13112,N_10777,N_10631);
or U13113 (N_13113,N_10248,N_11544);
xnor U13114 (N_13114,N_11197,N_10711);
and U13115 (N_13115,N_10122,N_10081);
nand U13116 (N_13116,N_11237,N_10247);
or U13117 (N_13117,N_11088,N_10472);
or U13118 (N_13118,N_11385,N_10700);
nor U13119 (N_13119,N_11095,N_11264);
nand U13120 (N_13120,N_11269,N_11624);
nand U13121 (N_13121,N_10864,N_11391);
nand U13122 (N_13122,N_11608,N_11275);
xnor U13123 (N_13123,N_11225,N_11774);
xnor U13124 (N_13124,N_10264,N_10013);
or U13125 (N_13125,N_10352,N_11373);
or U13126 (N_13126,N_10578,N_11806);
and U13127 (N_13127,N_11270,N_11124);
xor U13128 (N_13128,N_10160,N_10637);
nor U13129 (N_13129,N_10257,N_11289);
nor U13130 (N_13130,N_10780,N_10461);
nor U13131 (N_13131,N_10393,N_11191);
and U13132 (N_13132,N_11562,N_11980);
nand U13133 (N_13133,N_10042,N_10772);
xor U13134 (N_13134,N_11436,N_10434);
nand U13135 (N_13135,N_11026,N_10644);
or U13136 (N_13136,N_11451,N_11301);
nand U13137 (N_13137,N_11278,N_10447);
and U13138 (N_13138,N_11710,N_11395);
nand U13139 (N_13139,N_10388,N_10465);
xnor U13140 (N_13140,N_10499,N_10645);
or U13141 (N_13141,N_10779,N_10624);
nand U13142 (N_13142,N_10415,N_10103);
nand U13143 (N_13143,N_10603,N_10679);
or U13144 (N_13144,N_11813,N_11437);
nand U13145 (N_13145,N_11462,N_10184);
nand U13146 (N_13146,N_11444,N_11668);
or U13147 (N_13147,N_10815,N_10047);
and U13148 (N_13148,N_10890,N_11582);
xnor U13149 (N_13149,N_10865,N_10081);
or U13150 (N_13150,N_10524,N_10668);
or U13151 (N_13151,N_11898,N_10798);
or U13152 (N_13152,N_11154,N_11971);
and U13153 (N_13153,N_10904,N_10665);
nand U13154 (N_13154,N_11496,N_11732);
or U13155 (N_13155,N_11375,N_11871);
nand U13156 (N_13156,N_11594,N_10125);
and U13157 (N_13157,N_11327,N_10762);
or U13158 (N_13158,N_10382,N_11595);
or U13159 (N_13159,N_10143,N_10899);
and U13160 (N_13160,N_11930,N_11288);
nand U13161 (N_13161,N_10871,N_10140);
xor U13162 (N_13162,N_11003,N_11214);
nand U13163 (N_13163,N_10185,N_10311);
nor U13164 (N_13164,N_11069,N_10520);
and U13165 (N_13165,N_11548,N_10996);
nor U13166 (N_13166,N_10679,N_10021);
nand U13167 (N_13167,N_11616,N_10753);
nand U13168 (N_13168,N_10444,N_10666);
and U13169 (N_13169,N_11766,N_11875);
nor U13170 (N_13170,N_10977,N_11717);
or U13171 (N_13171,N_11648,N_11365);
nor U13172 (N_13172,N_11589,N_11745);
xnor U13173 (N_13173,N_11027,N_10743);
and U13174 (N_13174,N_11825,N_10077);
nor U13175 (N_13175,N_11932,N_10259);
nor U13176 (N_13176,N_10929,N_10928);
xnor U13177 (N_13177,N_11180,N_10891);
xor U13178 (N_13178,N_10629,N_11518);
nor U13179 (N_13179,N_10431,N_11750);
or U13180 (N_13180,N_11253,N_11570);
or U13181 (N_13181,N_10723,N_10257);
or U13182 (N_13182,N_10062,N_11148);
nor U13183 (N_13183,N_10759,N_10510);
nand U13184 (N_13184,N_10101,N_11084);
or U13185 (N_13185,N_10082,N_11737);
nand U13186 (N_13186,N_10681,N_11039);
nor U13187 (N_13187,N_11242,N_11515);
and U13188 (N_13188,N_10096,N_10910);
nand U13189 (N_13189,N_10720,N_10267);
nand U13190 (N_13190,N_10684,N_11636);
nor U13191 (N_13191,N_10318,N_11252);
xor U13192 (N_13192,N_11249,N_10799);
nand U13193 (N_13193,N_10519,N_11137);
and U13194 (N_13194,N_11186,N_11835);
nand U13195 (N_13195,N_10178,N_10342);
and U13196 (N_13196,N_11318,N_10327);
nor U13197 (N_13197,N_11070,N_10255);
and U13198 (N_13198,N_10999,N_10934);
xnor U13199 (N_13199,N_11919,N_11204);
nor U13200 (N_13200,N_11043,N_10856);
or U13201 (N_13201,N_10570,N_10719);
and U13202 (N_13202,N_10317,N_11011);
nand U13203 (N_13203,N_11801,N_10475);
and U13204 (N_13204,N_10368,N_10460);
or U13205 (N_13205,N_10257,N_11243);
or U13206 (N_13206,N_10210,N_10635);
and U13207 (N_13207,N_10570,N_11489);
and U13208 (N_13208,N_11584,N_10709);
or U13209 (N_13209,N_10199,N_10511);
or U13210 (N_13210,N_11017,N_11427);
xnor U13211 (N_13211,N_11743,N_10130);
nand U13212 (N_13212,N_11834,N_10617);
nor U13213 (N_13213,N_11079,N_10478);
nand U13214 (N_13214,N_11302,N_11729);
or U13215 (N_13215,N_11494,N_10077);
nand U13216 (N_13216,N_11429,N_11554);
and U13217 (N_13217,N_11209,N_10758);
nor U13218 (N_13218,N_11368,N_10304);
and U13219 (N_13219,N_10499,N_11665);
and U13220 (N_13220,N_11985,N_11756);
xnor U13221 (N_13221,N_10732,N_10741);
or U13222 (N_13222,N_11646,N_10279);
or U13223 (N_13223,N_11262,N_10400);
nor U13224 (N_13224,N_10169,N_10175);
nand U13225 (N_13225,N_11760,N_11033);
or U13226 (N_13226,N_10997,N_11855);
or U13227 (N_13227,N_11203,N_11834);
xnor U13228 (N_13228,N_11190,N_11763);
xor U13229 (N_13229,N_10293,N_11341);
and U13230 (N_13230,N_11936,N_10605);
and U13231 (N_13231,N_10432,N_10271);
xor U13232 (N_13232,N_10202,N_11799);
xnor U13233 (N_13233,N_10239,N_11338);
nand U13234 (N_13234,N_10120,N_11248);
xor U13235 (N_13235,N_11361,N_10092);
or U13236 (N_13236,N_11344,N_10727);
and U13237 (N_13237,N_11749,N_11555);
nand U13238 (N_13238,N_10530,N_10725);
or U13239 (N_13239,N_10899,N_11410);
nand U13240 (N_13240,N_10786,N_10199);
nor U13241 (N_13241,N_11218,N_11849);
and U13242 (N_13242,N_10687,N_10476);
and U13243 (N_13243,N_10405,N_10117);
xor U13244 (N_13244,N_11838,N_10557);
nor U13245 (N_13245,N_11626,N_10770);
or U13246 (N_13246,N_10237,N_11041);
nand U13247 (N_13247,N_11680,N_11222);
nand U13248 (N_13248,N_10636,N_11716);
or U13249 (N_13249,N_11010,N_11033);
nor U13250 (N_13250,N_10859,N_11785);
nand U13251 (N_13251,N_11501,N_11437);
nor U13252 (N_13252,N_10323,N_11145);
nand U13253 (N_13253,N_11137,N_11264);
or U13254 (N_13254,N_11455,N_11457);
xor U13255 (N_13255,N_10852,N_11881);
or U13256 (N_13256,N_11655,N_10400);
nand U13257 (N_13257,N_10343,N_10254);
and U13258 (N_13258,N_11850,N_11376);
and U13259 (N_13259,N_11623,N_10952);
xnor U13260 (N_13260,N_10992,N_10473);
nor U13261 (N_13261,N_10057,N_11409);
or U13262 (N_13262,N_11805,N_11877);
nand U13263 (N_13263,N_11182,N_10502);
and U13264 (N_13264,N_11471,N_10763);
nor U13265 (N_13265,N_10570,N_11926);
and U13266 (N_13266,N_10932,N_11960);
and U13267 (N_13267,N_11307,N_10437);
nor U13268 (N_13268,N_11363,N_11128);
and U13269 (N_13269,N_11039,N_11896);
nand U13270 (N_13270,N_10340,N_10649);
and U13271 (N_13271,N_10257,N_10543);
or U13272 (N_13272,N_10450,N_11668);
and U13273 (N_13273,N_11415,N_10475);
xnor U13274 (N_13274,N_11279,N_11164);
and U13275 (N_13275,N_10552,N_10213);
xor U13276 (N_13276,N_11899,N_10674);
and U13277 (N_13277,N_10146,N_10813);
and U13278 (N_13278,N_10378,N_10737);
and U13279 (N_13279,N_11947,N_10420);
xor U13280 (N_13280,N_10292,N_11665);
and U13281 (N_13281,N_11116,N_11698);
and U13282 (N_13282,N_10679,N_10633);
and U13283 (N_13283,N_11225,N_11187);
or U13284 (N_13284,N_11386,N_11676);
and U13285 (N_13285,N_10156,N_11901);
nand U13286 (N_13286,N_11970,N_10896);
nand U13287 (N_13287,N_10672,N_11982);
and U13288 (N_13288,N_11252,N_11109);
or U13289 (N_13289,N_11172,N_11746);
xnor U13290 (N_13290,N_11754,N_10065);
xor U13291 (N_13291,N_11407,N_10982);
or U13292 (N_13292,N_11068,N_11482);
xor U13293 (N_13293,N_10623,N_10060);
nor U13294 (N_13294,N_10994,N_11501);
xnor U13295 (N_13295,N_11620,N_10812);
or U13296 (N_13296,N_11022,N_10845);
or U13297 (N_13297,N_10200,N_10815);
nor U13298 (N_13298,N_11131,N_10697);
nor U13299 (N_13299,N_11436,N_10454);
or U13300 (N_13300,N_10557,N_11907);
and U13301 (N_13301,N_11185,N_11846);
nand U13302 (N_13302,N_11745,N_10544);
nor U13303 (N_13303,N_11399,N_10660);
nand U13304 (N_13304,N_11217,N_11587);
nand U13305 (N_13305,N_11041,N_11047);
or U13306 (N_13306,N_10241,N_11875);
and U13307 (N_13307,N_10329,N_10125);
xnor U13308 (N_13308,N_10822,N_10831);
and U13309 (N_13309,N_11225,N_10405);
and U13310 (N_13310,N_11414,N_11780);
nand U13311 (N_13311,N_11368,N_11174);
nand U13312 (N_13312,N_10805,N_11697);
nor U13313 (N_13313,N_11752,N_10147);
nand U13314 (N_13314,N_10886,N_11339);
nor U13315 (N_13315,N_10468,N_11193);
nand U13316 (N_13316,N_10219,N_10653);
xnor U13317 (N_13317,N_10531,N_10802);
and U13318 (N_13318,N_11519,N_11711);
or U13319 (N_13319,N_11998,N_10863);
xor U13320 (N_13320,N_10762,N_11490);
nor U13321 (N_13321,N_11834,N_11871);
nor U13322 (N_13322,N_10399,N_10035);
or U13323 (N_13323,N_11507,N_11249);
nor U13324 (N_13324,N_11630,N_10627);
nand U13325 (N_13325,N_10972,N_10758);
nor U13326 (N_13326,N_11131,N_11578);
or U13327 (N_13327,N_10952,N_10042);
xnor U13328 (N_13328,N_10479,N_11111);
nand U13329 (N_13329,N_11095,N_11844);
nand U13330 (N_13330,N_11529,N_11814);
or U13331 (N_13331,N_10270,N_11512);
xnor U13332 (N_13332,N_10170,N_11587);
and U13333 (N_13333,N_10406,N_11513);
or U13334 (N_13334,N_10142,N_11544);
and U13335 (N_13335,N_10459,N_10915);
and U13336 (N_13336,N_11383,N_10663);
or U13337 (N_13337,N_10832,N_11520);
nand U13338 (N_13338,N_11900,N_10254);
or U13339 (N_13339,N_10885,N_11974);
and U13340 (N_13340,N_10412,N_11782);
xor U13341 (N_13341,N_11282,N_11414);
and U13342 (N_13342,N_11344,N_10885);
and U13343 (N_13343,N_10247,N_11670);
nor U13344 (N_13344,N_10193,N_10560);
or U13345 (N_13345,N_11377,N_10407);
nand U13346 (N_13346,N_10635,N_11981);
or U13347 (N_13347,N_10965,N_10070);
xnor U13348 (N_13348,N_10792,N_11902);
xor U13349 (N_13349,N_10674,N_11113);
and U13350 (N_13350,N_11579,N_10873);
nor U13351 (N_13351,N_10307,N_11017);
xnor U13352 (N_13352,N_10924,N_11298);
or U13353 (N_13353,N_10921,N_11541);
xnor U13354 (N_13354,N_10380,N_11981);
nor U13355 (N_13355,N_10043,N_10781);
nand U13356 (N_13356,N_11729,N_11756);
nand U13357 (N_13357,N_11081,N_10429);
nand U13358 (N_13358,N_11636,N_11643);
or U13359 (N_13359,N_11856,N_10525);
or U13360 (N_13360,N_10670,N_11236);
nand U13361 (N_13361,N_11898,N_10092);
nor U13362 (N_13362,N_10961,N_10217);
or U13363 (N_13363,N_11746,N_11435);
xor U13364 (N_13364,N_11117,N_11996);
and U13365 (N_13365,N_11264,N_10218);
or U13366 (N_13366,N_10062,N_11688);
and U13367 (N_13367,N_11186,N_10706);
or U13368 (N_13368,N_10182,N_11759);
nand U13369 (N_13369,N_10899,N_11809);
or U13370 (N_13370,N_10030,N_10636);
and U13371 (N_13371,N_10120,N_10108);
or U13372 (N_13372,N_11570,N_10534);
or U13373 (N_13373,N_11557,N_10015);
nand U13374 (N_13374,N_10367,N_11805);
xnor U13375 (N_13375,N_11617,N_10068);
xnor U13376 (N_13376,N_10998,N_10885);
nand U13377 (N_13377,N_11705,N_11150);
xnor U13378 (N_13378,N_11894,N_10281);
nor U13379 (N_13379,N_11972,N_11145);
nand U13380 (N_13380,N_11458,N_11076);
xor U13381 (N_13381,N_10021,N_11221);
or U13382 (N_13382,N_11308,N_11773);
xor U13383 (N_13383,N_11988,N_11331);
xor U13384 (N_13384,N_11935,N_10186);
nor U13385 (N_13385,N_10113,N_11473);
nand U13386 (N_13386,N_11984,N_11469);
and U13387 (N_13387,N_11847,N_11401);
or U13388 (N_13388,N_11208,N_11337);
or U13389 (N_13389,N_11592,N_10300);
or U13390 (N_13390,N_11484,N_11338);
and U13391 (N_13391,N_11249,N_11240);
or U13392 (N_13392,N_10876,N_11308);
nand U13393 (N_13393,N_11066,N_11708);
nor U13394 (N_13394,N_11153,N_11833);
nor U13395 (N_13395,N_10037,N_10758);
or U13396 (N_13396,N_11130,N_11452);
nor U13397 (N_13397,N_11006,N_11509);
xor U13398 (N_13398,N_10823,N_10498);
and U13399 (N_13399,N_11503,N_10988);
nor U13400 (N_13400,N_11749,N_11588);
or U13401 (N_13401,N_11684,N_10264);
xor U13402 (N_13402,N_11337,N_10057);
nand U13403 (N_13403,N_10888,N_10906);
and U13404 (N_13404,N_10104,N_11885);
nand U13405 (N_13405,N_10012,N_10410);
nor U13406 (N_13406,N_10805,N_10339);
xnor U13407 (N_13407,N_10656,N_10771);
xnor U13408 (N_13408,N_11776,N_10928);
or U13409 (N_13409,N_11165,N_11761);
or U13410 (N_13410,N_10796,N_11315);
and U13411 (N_13411,N_11318,N_11877);
xor U13412 (N_13412,N_11496,N_10809);
and U13413 (N_13413,N_10417,N_10627);
or U13414 (N_13414,N_11710,N_10202);
xor U13415 (N_13415,N_11868,N_10769);
nor U13416 (N_13416,N_11854,N_11963);
xnor U13417 (N_13417,N_10424,N_10341);
nand U13418 (N_13418,N_10218,N_10697);
nor U13419 (N_13419,N_10222,N_11365);
and U13420 (N_13420,N_10910,N_10487);
or U13421 (N_13421,N_10542,N_10694);
nand U13422 (N_13422,N_11132,N_11165);
or U13423 (N_13423,N_11821,N_11680);
nand U13424 (N_13424,N_10861,N_11166);
and U13425 (N_13425,N_10436,N_10200);
nor U13426 (N_13426,N_11006,N_11578);
or U13427 (N_13427,N_10727,N_10867);
xnor U13428 (N_13428,N_11036,N_11013);
xor U13429 (N_13429,N_10862,N_10155);
nor U13430 (N_13430,N_10701,N_11880);
xor U13431 (N_13431,N_11164,N_11595);
nand U13432 (N_13432,N_11951,N_11702);
or U13433 (N_13433,N_11856,N_10995);
nand U13434 (N_13434,N_10714,N_11094);
or U13435 (N_13435,N_11163,N_11219);
or U13436 (N_13436,N_10782,N_10133);
nor U13437 (N_13437,N_11499,N_11431);
nand U13438 (N_13438,N_10709,N_11247);
and U13439 (N_13439,N_10043,N_10475);
nor U13440 (N_13440,N_10070,N_10261);
nand U13441 (N_13441,N_11020,N_11812);
xnor U13442 (N_13442,N_11505,N_10061);
and U13443 (N_13443,N_10254,N_10367);
nor U13444 (N_13444,N_10441,N_10470);
nand U13445 (N_13445,N_11023,N_11155);
or U13446 (N_13446,N_11501,N_11513);
nand U13447 (N_13447,N_10936,N_11332);
nand U13448 (N_13448,N_10771,N_11079);
xor U13449 (N_13449,N_11733,N_10346);
nand U13450 (N_13450,N_10391,N_10390);
nor U13451 (N_13451,N_10156,N_11775);
xnor U13452 (N_13452,N_11970,N_11917);
xnor U13453 (N_13453,N_10409,N_10441);
or U13454 (N_13454,N_10430,N_11931);
and U13455 (N_13455,N_11145,N_10602);
nor U13456 (N_13456,N_11508,N_10186);
and U13457 (N_13457,N_11404,N_10481);
nand U13458 (N_13458,N_11950,N_10457);
xor U13459 (N_13459,N_11305,N_11181);
xor U13460 (N_13460,N_11828,N_10301);
xnor U13461 (N_13461,N_10437,N_11086);
and U13462 (N_13462,N_11689,N_11264);
xnor U13463 (N_13463,N_11197,N_10629);
nand U13464 (N_13464,N_10060,N_11459);
and U13465 (N_13465,N_10504,N_11747);
nor U13466 (N_13466,N_11216,N_10879);
nor U13467 (N_13467,N_11357,N_11048);
nand U13468 (N_13468,N_10784,N_11953);
xnor U13469 (N_13469,N_11372,N_11406);
nor U13470 (N_13470,N_11894,N_10135);
nand U13471 (N_13471,N_11365,N_11122);
nor U13472 (N_13472,N_11065,N_11337);
xnor U13473 (N_13473,N_11588,N_10710);
nand U13474 (N_13474,N_11647,N_11061);
nand U13475 (N_13475,N_11117,N_10435);
nor U13476 (N_13476,N_11690,N_10272);
xnor U13477 (N_13477,N_11441,N_10642);
and U13478 (N_13478,N_11563,N_11215);
and U13479 (N_13479,N_10491,N_10438);
xor U13480 (N_13480,N_10730,N_10948);
or U13481 (N_13481,N_11159,N_10050);
nand U13482 (N_13482,N_10649,N_10096);
xnor U13483 (N_13483,N_11243,N_11568);
xnor U13484 (N_13484,N_11799,N_10392);
or U13485 (N_13485,N_10409,N_10832);
or U13486 (N_13486,N_11196,N_10298);
xnor U13487 (N_13487,N_11722,N_11705);
xnor U13488 (N_13488,N_10250,N_11366);
xor U13489 (N_13489,N_10498,N_10451);
nand U13490 (N_13490,N_11156,N_11643);
and U13491 (N_13491,N_10041,N_11260);
nor U13492 (N_13492,N_10875,N_10961);
and U13493 (N_13493,N_11136,N_10488);
or U13494 (N_13494,N_10600,N_10029);
or U13495 (N_13495,N_10999,N_10751);
nor U13496 (N_13496,N_10407,N_10001);
nand U13497 (N_13497,N_10727,N_11609);
xor U13498 (N_13498,N_10184,N_11439);
or U13499 (N_13499,N_10560,N_11046);
nor U13500 (N_13500,N_11274,N_11145);
and U13501 (N_13501,N_11137,N_11155);
nor U13502 (N_13502,N_11727,N_11759);
nor U13503 (N_13503,N_11895,N_11113);
nand U13504 (N_13504,N_10379,N_11115);
xor U13505 (N_13505,N_11564,N_10393);
xor U13506 (N_13506,N_10187,N_10761);
nor U13507 (N_13507,N_11722,N_10795);
nand U13508 (N_13508,N_10148,N_11322);
xnor U13509 (N_13509,N_10460,N_10091);
nor U13510 (N_13510,N_11332,N_10969);
nand U13511 (N_13511,N_10867,N_11180);
nand U13512 (N_13512,N_10198,N_11092);
xnor U13513 (N_13513,N_11714,N_11637);
nand U13514 (N_13514,N_10980,N_11391);
nand U13515 (N_13515,N_10911,N_10464);
xnor U13516 (N_13516,N_10818,N_11434);
or U13517 (N_13517,N_11483,N_10417);
nor U13518 (N_13518,N_10597,N_11584);
or U13519 (N_13519,N_11133,N_10807);
nand U13520 (N_13520,N_10471,N_10093);
and U13521 (N_13521,N_11952,N_10852);
and U13522 (N_13522,N_11140,N_11575);
and U13523 (N_13523,N_11647,N_11012);
or U13524 (N_13524,N_11393,N_10135);
or U13525 (N_13525,N_10941,N_10466);
xnor U13526 (N_13526,N_10964,N_11953);
and U13527 (N_13527,N_11609,N_10021);
xnor U13528 (N_13528,N_10456,N_10954);
xor U13529 (N_13529,N_10299,N_10186);
nor U13530 (N_13530,N_10191,N_10832);
or U13531 (N_13531,N_10219,N_10026);
nor U13532 (N_13532,N_10504,N_10722);
nor U13533 (N_13533,N_11772,N_10517);
and U13534 (N_13534,N_10625,N_10697);
nor U13535 (N_13535,N_10514,N_10849);
and U13536 (N_13536,N_10891,N_11883);
and U13537 (N_13537,N_11399,N_11864);
nor U13538 (N_13538,N_10755,N_11702);
nand U13539 (N_13539,N_10517,N_11204);
nand U13540 (N_13540,N_10827,N_10763);
nand U13541 (N_13541,N_11050,N_10593);
nand U13542 (N_13542,N_11676,N_11520);
xor U13543 (N_13543,N_11126,N_10700);
or U13544 (N_13544,N_11899,N_11465);
nor U13545 (N_13545,N_11060,N_11514);
or U13546 (N_13546,N_11307,N_10885);
nor U13547 (N_13547,N_11888,N_11303);
and U13548 (N_13548,N_11799,N_10461);
or U13549 (N_13549,N_11589,N_10393);
and U13550 (N_13550,N_11818,N_11995);
nor U13551 (N_13551,N_11962,N_11231);
xor U13552 (N_13552,N_10070,N_10577);
nor U13553 (N_13553,N_10701,N_10579);
nand U13554 (N_13554,N_10080,N_11000);
or U13555 (N_13555,N_10767,N_10783);
xor U13556 (N_13556,N_10093,N_10078);
nor U13557 (N_13557,N_10924,N_10451);
or U13558 (N_13558,N_10822,N_11263);
xnor U13559 (N_13559,N_11386,N_10010);
nand U13560 (N_13560,N_11606,N_10241);
nand U13561 (N_13561,N_11835,N_11018);
and U13562 (N_13562,N_10831,N_10600);
xnor U13563 (N_13563,N_11900,N_10630);
or U13564 (N_13564,N_10039,N_11367);
and U13565 (N_13565,N_10022,N_10060);
nor U13566 (N_13566,N_10210,N_11937);
nor U13567 (N_13567,N_10748,N_10184);
xor U13568 (N_13568,N_10764,N_10332);
or U13569 (N_13569,N_10045,N_10485);
and U13570 (N_13570,N_10824,N_11049);
or U13571 (N_13571,N_11641,N_11682);
and U13572 (N_13572,N_10181,N_11398);
or U13573 (N_13573,N_10677,N_11371);
nand U13574 (N_13574,N_10597,N_10945);
or U13575 (N_13575,N_11210,N_10101);
nor U13576 (N_13576,N_11662,N_11087);
and U13577 (N_13577,N_10460,N_11748);
or U13578 (N_13578,N_10499,N_10202);
nor U13579 (N_13579,N_10654,N_11603);
nand U13580 (N_13580,N_10063,N_10483);
nand U13581 (N_13581,N_11296,N_11938);
nand U13582 (N_13582,N_10544,N_11384);
and U13583 (N_13583,N_11748,N_11628);
xnor U13584 (N_13584,N_11081,N_11028);
xnor U13585 (N_13585,N_11607,N_11378);
and U13586 (N_13586,N_11478,N_11419);
nand U13587 (N_13587,N_11905,N_11704);
nand U13588 (N_13588,N_10305,N_11568);
nand U13589 (N_13589,N_10953,N_10454);
and U13590 (N_13590,N_11774,N_11055);
nor U13591 (N_13591,N_11399,N_11957);
and U13592 (N_13592,N_10100,N_11071);
nor U13593 (N_13593,N_10972,N_10134);
nor U13594 (N_13594,N_11869,N_10484);
xnor U13595 (N_13595,N_10925,N_11685);
and U13596 (N_13596,N_11414,N_10977);
or U13597 (N_13597,N_11499,N_11700);
and U13598 (N_13598,N_11010,N_10995);
xor U13599 (N_13599,N_11434,N_11406);
and U13600 (N_13600,N_10223,N_11573);
nor U13601 (N_13601,N_10204,N_11067);
and U13602 (N_13602,N_11100,N_11186);
and U13603 (N_13603,N_10843,N_11550);
xor U13604 (N_13604,N_10188,N_11830);
nand U13605 (N_13605,N_11886,N_10891);
or U13606 (N_13606,N_11208,N_10332);
xnor U13607 (N_13607,N_10591,N_10045);
xor U13608 (N_13608,N_10644,N_10661);
and U13609 (N_13609,N_10599,N_10493);
nand U13610 (N_13610,N_11716,N_11241);
nor U13611 (N_13611,N_11437,N_11634);
nand U13612 (N_13612,N_11237,N_10319);
xnor U13613 (N_13613,N_11348,N_10895);
and U13614 (N_13614,N_11491,N_10150);
xor U13615 (N_13615,N_10029,N_11508);
nand U13616 (N_13616,N_11272,N_11164);
or U13617 (N_13617,N_10386,N_11469);
and U13618 (N_13618,N_11167,N_11510);
nand U13619 (N_13619,N_10176,N_10181);
nand U13620 (N_13620,N_11317,N_11231);
nor U13621 (N_13621,N_11153,N_10933);
or U13622 (N_13622,N_11151,N_10639);
xnor U13623 (N_13623,N_10260,N_10488);
nor U13624 (N_13624,N_11582,N_10101);
nor U13625 (N_13625,N_11791,N_10482);
nand U13626 (N_13626,N_10340,N_10262);
or U13627 (N_13627,N_11282,N_10039);
nand U13628 (N_13628,N_11544,N_10951);
nand U13629 (N_13629,N_10118,N_11611);
nor U13630 (N_13630,N_10867,N_11128);
nand U13631 (N_13631,N_11138,N_11438);
or U13632 (N_13632,N_11815,N_11629);
and U13633 (N_13633,N_11644,N_10188);
xnor U13634 (N_13634,N_10234,N_10559);
and U13635 (N_13635,N_11056,N_10983);
and U13636 (N_13636,N_10476,N_10507);
xnor U13637 (N_13637,N_10955,N_11884);
and U13638 (N_13638,N_10179,N_11415);
nor U13639 (N_13639,N_10510,N_10729);
nand U13640 (N_13640,N_10765,N_10856);
xor U13641 (N_13641,N_10442,N_10057);
and U13642 (N_13642,N_10452,N_10245);
and U13643 (N_13643,N_11243,N_10749);
xor U13644 (N_13644,N_11799,N_10855);
nor U13645 (N_13645,N_11742,N_10181);
nor U13646 (N_13646,N_11153,N_10551);
or U13647 (N_13647,N_11204,N_11625);
xnor U13648 (N_13648,N_11966,N_10797);
or U13649 (N_13649,N_10250,N_10429);
nor U13650 (N_13650,N_11815,N_11417);
and U13651 (N_13651,N_10051,N_10122);
or U13652 (N_13652,N_11750,N_10811);
xor U13653 (N_13653,N_10436,N_10831);
and U13654 (N_13654,N_10057,N_11084);
or U13655 (N_13655,N_10308,N_10930);
nand U13656 (N_13656,N_11552,N_11134);
nor U13657 (N_13657,N_11906,N_11666);
xor U13658 (N_13658,N_11657,N_11556);
nor U13659 (N_13659,N_11356,N_11526);
or U13660 (N_13660,N_10874,N_11658);
nor U13661 (N_13661,N_10884,N_11036);
or U13662 (N_13662,N_10311,N_11090);
nand U13663 (N_13663,N_10253,N_10800);
or U13664 (N_13664,N_11216,N_10385);
and U13665 (N_13665,N_11620,N_10737);
nor U13666 (N_13666,N_10364,N_10436);
xnor U13667 (N_13667,N_11667,N_10581);
and U13668 (N_13668,N_11170,N_10362);
or U13669 (N_13669,N_10221,N_10965);
nand U13670 (N_13670,N_10413,N_11541);
nand U13671 (N_13671,N_11799,N_11598);
xor U13672 (N_13672,N_11938,N_10154);
or U13673 (N_13673,N_11869,N_10375);
and U13674 (N_13674,N_10645,N_11044);
nor U13675 (N_13675,N_11459,N_11021);
nor U13676 (N_13676,N_10025,N_11897);
and U13677 (N_13677,N_10513,N_10284);
nor U13678 (N_13678,N_10282,N_10162);
or U13679 (N_13679,N_11600,N_11234);
xor U13680 (N_13680,N_11601,N_10249);
nor U13681 (N_13681,N_10646,N_10206);
nor U13682 (N_13682,N_10381,N_11505);
or U13683 (N_13683,N_10952,N_10144);
and U13684 (N_13684,N_11018,N_11349);
xor U13685 (N_13685,N_11803,N_11012);
and U13686 (N_13686,N_11908,N_10984);
and U13687 (N_13687,N_10220,N_10173);
nor U13688 (N_13688,N_11579,N_10901);
xnor U13689 (N_13689,N_10267,N_10282);
nand U13690 (N_13690,N_11419,N_10195);
and U13691 (N_13691,N_10991,N_11756);
and U13692 (N_13692,N_10773,N_10491);
and U13693 (N_13693,N_10683,N_11425);
or U13694 (N_13694,N_11950,N_10381);
and U13695 (N_13695,N_11843,N_11911);
nand U13696 (N_13696,N_10115,N_11721);
nor U13697 (N_13697,N_10328,N_10542);
or U13698 (N_13698,N_10986,N_11780);
or U13699 (N_13699,N_11030,N_11885);
and U13700 (N_13700,N_10892,N_11036);
and U13701 (N_13701,N_10833,N_10677);
xnor U13702 (N_13702,N_11437,N_10625);
nor U13703 (N_13703,N_11212,N_10080);
nand U13704 (N_13704,N_10942,N_11541);
xnor U13705 (N_13705,N_10467,N_11941);
xor U13706 (N_13706,N_10996,N_11646);
nand U13707 (N_13707,N_11314,N_10530);
xnor U13708 (N_13708,N_11174,N_10261);
xor U13709 (N_13709,N_10803,N_10482);
and U13710 (N_13710,N_10527,N_11981);
and U13711 (N_13711,N_11338,N_11481);
and U13712 (N_13712,N_10585,N_11604);
or U13713 (N_13713,N_10637,N_11199);
or U13714 (N_13714,N_11158,N_10873);
and U13715 (N_13715,N_11602,N_11479);
xnor U13716 (N_13716,N_10320,N_10724);
nand U13717 (N_13717,N_11887,N_11096);
nand U13718 (N_13718,N_10299,N_10348);
or U13719 (N_13719,N_11057,N_10143);
and U13720 (N_13720,N_11365,N_10082);
nand U13721 (N_13721,N_11222,N_11876);
nand U13722 (N_13722,N_10598,N_11597);
xnor U13723 (N_13723,N_11489,N_11622);
nand U13724 (N_13724,N_11822,N_10659);
nand U13725 (N_13725,N_10297,N_11562);
and U13726 (N_13726,N_10797,N_10683);
nor U13727 (N_13727,N_11406,N_10832);
and U13728 (N_13728,N_11515,N_10492);
nand U13729 (N_13729,N_11281,N_11046);
xnor U13730 (N_13730,N_10715,N_10098);
or U13731 (N_13731,N_10643,N_11744);
or U13732 (N_13732,N_11451,N_10657);
nand U13733 (N_13733,N_10856,N_10178);
or U13734 (N_13734,N_10745,N_11218);
xor U13735 (N_13735,N_10054,N_10093);
or U13736 (N_13736,N_11161,N_10839);
and U13737 (N_13737,N_11747,N_11390);
and U13738 (N_13738,N_11753,N_11219);
or U13739 (N_13739,N_11789,N_11036);
nor U13740 (N_13740,N_11840,N_10639);
or U13741 (N_13741,N_10434,N_10164);
or U13742 (N_13742,N_10111,N_10815);
nor U13743 (N_13743,N_11700,N_10931);
xor U13744 (N_13744,N_10439,N_10248);
nand U13745 (N_13745,N_10701,N_11930);
or U13746 (N_13746,N_11589,N_11526);
nor U13747 (N_13747,N_10695,N_11703);
nand U13748 (N_13748,N_11563,N_11164);
nand U13749 (N_13749,N_10101,N_10540);
nand U13750 (N_13750,N_11771,N_11754);
or U13751 (N_13751,N_10559,N_10778);
xor U13752 (N_13752,N_11749,N_10260);
xor U13753 (N_13753,N_11336,N_10771);
nand U13754 (N_13754,N_10707,N_10251);
or U13755 (N_13755,N_11789,N_11974);
and U13756 (N_13756,N_11174,N_10566);
nand U13757 (N_13757,N_10349,N_10606);
or U13758 (N_13758,N_11437,N_10228);
and U13759 (N_13759,N_10943,N_10434);
nand U13760 (N_13760,N_11015,N_10442);
xnor U13761 (N_13761,N_10902,N_10758);
nand U13762 (N_13762,N_11637,N_11372);
xnor U13763 (N_13763,N_10992,N_11599);
xor U13764 (N_13764,N_10301,N_10672);
or U13765 (N_13765,N_10895,N_11723);
or U13766 (N_13766,N_11787,N_11565);
and U13767 (N_13767,N_11182,N_11672);
or U13768 (N_13768,N_10886,N_10854);
nor U13769 (N_13769,N_11437,N_11457);
and U13770 (N_13770,N_10635,N_10534);
and U13771 (N_13771,N_11529,N_10217);
or U13772 (N_13772,N_10357,N_11399);
or U13773 (N_13773,N_11979,N_10734);
nor U13774 (N_13774,N_10441,N_10755);
or U13775 (N_13775,N_10734,N_10411);
or U13776 (N_13776,N_11639,N_11064);
nand U13777 (N_13777,N_11628,N_11741);
xor U13778 (N_13778,N_10631,N_10188);
and U13779 (N_13779,N_11732,N_11151);
xnor U13780 (N_13780,N_10475,N_10549);
or U13781 (N_13781,N_11323,N_11075);
nor U13782 (N_13782,N_11289,N_10357);
or U13783 (N_13783,N_11698,N_10031);
nor U13784 (N_13784,N_10200,N_10362);
or U13785 (N_13785,N_11931,N_11505);
nand U13786 (N_13786,N_11809,N_11713);
or U13787 (N_13787,N_10167,N_11523);
nand U13788 (N_13788,N_11427,N_11960);
or U13789 (N_13789,N_10701,N_11918);
or U13790 (N_13790,N_11492,N_11903);
or U13791 (N_13791,N_11955,N_10154);
xnor U13792 (N_13792,N_10778,N_10290);
xnor U13793 (N_13793,N_10878,N_10480);
nor U13794 (N_13794,N_11650,N_10213);
nand U13795 (N_13795,N_10205,N_11709);
nor U13796 (N_13796,N_11266,N_10464);
and U13797 (N_13797,N_10802,N_10357);
nand U13798 (N_13798,N_10649,N_10760);
xnor U13799 (N_13799,N_10197,N_10881);
nand U13800 (N_13800,N_10831,N_11945);
or U13801 (N_13801,N_10829,N_10718);
nor U13802 (N_13802,N_10909,N_10541);
and U13803 (N_13803,N_11305,N_11642);
nor U13804 (N_13804,N_10598,N_10204);
xnor U13805 (N_13805,N_11376,N_11219);
nand U13806 (N_13806,N_10125,N_10580);
or U13807 (N_13807,N_11280,N_11905);
and U13808 (N_13808,N_11848,N_10014);
or U13809 (N_13809,N_10017,N_10221);
nand U13810 (N_13810,N_10674,N_11008);
nand U13811 (N_13811,N_10625,N_11214);
xnor U13812 (N_13812,N_10014,N_10971);
xor U13813 (N_13813,N_10832,N_11135);
or U13814 (N_13814,N_11369,N_10962);
or U13815 (N_13815,N_11320,N_11954);
nand U13816 (N_13816,N_11473,N_11246);
or U13817 (N_13817,N_11244,N_10883);
xor U13818 (N_13818,N_10185,N_10765);
nor U13819 (N_13819,N_10442,N_10487);
xnor U13820 (N_13820,N_10689,N_10062);
nand U13821 (N_13821,N_10864,N_11369);
or U13822 (N_13822,N_10101,N_10623);
and U13823 (N_13823,N_11367,N_10775);
or U13824 (N_13824,N_11399,N_10879);
xnor U13825 (N_13825,N_11405,N_11624);
nor U13826 (N_13826,N_11385,N_10129);
and U13827 (N_13827,N_11048,N_10096);
nand U13828 (N_13828,N_11931,N_11854);
nand U13829 (N_13829,N_11716,N_11923);
nor U13830 (N_13830,N_10985,N_10388);
and U13831 (N_13831,N_10812,N_10999);
or U13832 (N_13832,N_11391,N_10914);
nor U13833 (N_13833,N_11301,N_11956);
and U13834 (N_13834,N_11012,N_10677);
or U13835 (N_13835,N_11180,N_10912);
and U13836 (N_13836,N_10211,N_11918);
xnor U13837 (N_13837,N_11223,N_11585);
xnor U13838 (N_13838,N_11769,N_10284);
nand U13839 (N_13839,N_10790,N_10424);
xor U13840 (N_13840,N_10532,N_11433);
xor U13841 (N_13841,N_10643,N_11761);
nand U13842 (N_13842,N_10894,N_10799);
nand U13843 (N_13843,N_10061,N_11008);
or U13844 (N_13844,N_10609,N_11237);
nand U13845 (N_13845,N_11324,N_10244);
and U13846 (N_13846,N_10445,N_11097);
and U13847 (N_13847,N_11728,N_11419);
nor U13848 (N_13848,N_10215,N_10028);
or U13849 (N_13849,N_10904,N_11242);
nor U13850 (N_13850,N_10369,N_11462);
nand U13851 (N_13851,N_10786,N_11501);
nand U13852 (N_13852,N_11686,N_10417);
nand U13853 (N_13853,N_10001,N_10095);
nor U13854 (N_13854,N_10259,N_11101);
and U13855 (N_13855,N_11262,N_11594);
and U13856 (N_13856,N_11309,N_10694);
xnor U13857 (N_13857,N_11402,N_11597);
nand U13858 (N_13858,N_10688,N_11431);
nor U13859 (N_13859,N_10038,N_10977);
or U13860 (N_13860,N_11761,N_11461);
xnor U13861 (N_13861,N_11639,N_10656);
and U13862 (N_13862,N_11890,N_10564);
or U13863 (N_13863,N_10749,N_10262);
or U13864 (N_13864,N_10250,N_10770);
and U13865 (N_13865,N_10481,N_11702);
and U13866 (N_13866,N_11002,N_11597);
xnor U13867 (N_13867,N_10178,N_10009);
nand U13868 (N_13868,N_10053,N_10231);
nand U13869 (N_13869,N_10140,N_10146);
and U13870 (N_13870,N_11387,N_11999);
xnor U13871 (N_13871,N_11795,N_11478);
or U13872 (N_13872,N_11422,N_10169);
and U13873 (N_13873,N_11857,N_11091);
nand U13874 (N_13874,N_10958,N_11689);
nor U13875 (N_13875,N_10378,N_10137);
and U13876 (N_13876,N_11593,N_10339);
and U13877 (N_13877,N_11351,N_10104);
nand U13878 (N_13878,N_10260,N_11499);
and U13879 (N_13879,N_10537,N_11375);
nand U13880 (N_13880,N_11311,N_11617);
nand U13881 (N_13881,N_10188,N_11490);
nor U13882 (N_13882,N_10277,N_10955);
nand U13883 (N_13883,N_11092,N_11512);
nand U13884 (N_13884,N_11512,N_11509);
and U13885 (N_13885,N_10394,N_11283);
xor U13886 (N_13886,N_11646,N_10305);
nor U13887 (N_13887,N_10584,N_11060);
nand U13888 (N_13888,N_11175,N_10683);
nor U13889 (N_13889,N_10039,N_11179);
and U13890 (N_13890,N_11376,N_11063);
and U13891 (N_13891,N_10244,N_10582);
and U13892 (N_13892,N_10018,N_11199);
nor U13893 (N_13893,N_10419,N_10835);
nor U13894 (N_13894,N_11322,N_11290);
nand U13895 (N_13895,N_10067,N_11583);
xnor U13896 (N_13896,N_10818,N_11274);
and U13897 (N_13897,N_10104,N_10715);
xnor U13898 (N_13898,N_11538,N_11324);
and U13899 (N_13899,N_11868,N_10611);
and U13900 (N_13900,N_10785,N_10453);
or U13901 (N_13901,N_10127,N_10593);
xor U13902 (N_13902,N_10509,N_10257);
nand U13903 (N_13903,N_11315,N_11358);
or U13904 (N_13904,N_10894,N_11512);
nand U13905 (N_13905,N_11885,N_10172);
nor U13906 (N_13906,N_10418,N_11334);
nand U13907 (N_13907,N_11117,N_11982);
and U13908 (N_13908,N_10685,N_10508);
xor U13909 (N_13909,N_11796,N_10183);
xnor U13910 (N_13910,N_11674,N_10961);
or U13911 (N_13911,N_11838,N_10209);
xnor U13912 (N_13912,N_11151,N_10855);
or U13913 (N_13913,N_10066,N_11128);
and U13914 (N_13914,N_11379,N_10889);
nor U13915 (N_13915,N_11701,N_10695);
or U13916 (N_13916,N_11999,N_10660);
nor U13917 (N_13917,N_11908,N_11050);
nor U13918 (N_13918,N_11536,N_10613);
and U13919 (N_13919,N_11666,N_10780);
nand U13920 (N_13920,N_10047,N_10248);
xnor U13921 (N_13921,N_10730,N_11361);
nor U13922 (N_13922,N_10740,N_10359);
and U13923 (N_13923,N_10729,N_10057);
xor U13924 (N_13924,N_10186,N_11194);
and U13925 (N_13925,N_10462,N_10626);
or U13926 (N_13926,N_11695,N_11852);
and U13927 (N_13927,N_10740,N_10699);
or U13928 (N_13928,N_11860,N_10395);
or U13929 (N_13929,N_10907,N_10093);
nand U13930 (N_13930,N_11108,N_10583);
or U13931 (N_13931,N_10090,N_11475);
xnor U13932 (N_13932,N_10122,N_11773);
and U13933 (N_13933,N_11644,N_11158);
nor U13934 (N_13934,N_10406,N_11632);
and U13935 (N_13935,N_10405,N_11944);
xor U13936 (N_13936,N_11220,N_10059);
nand U13937 (N_13937,N_10606,N_10192);
or U13938 (N_13938,N_10874,N_10727);
nand U13939 (N_13939,N_10357,N_10808);
or U13940 (N_13940,N_11719,N_11139);
and U13941 (N_13941,N_11792,N_11655);
nor U13942 (N_13942,N_11018,N_10392);
nand U13943 (N_13943,N_10450,N_11746);
nand U13944 (N_13944,N_10709,N_10870);
nand U13945 (N_13945,N_10934,N_11562);
nor U13946 (N_13946,N_10170,N_10599);
nor U13947 (N_13947,N_11799,N_11362);
nand U13948 (N_13948,N_11940,N_10945);
nor U13949 (N_13949,N_11178,N_11134);
or U13950 (N_13950,N_11246,N_11795);
xnor U13951 (N_13951,N_11904,N_10506);
and U13952 (N_13952,N_11206,N_11689);
or U13953 (N_13953,N_10475,N_11361);
nor U13954 (N_13954,N_11093,N_11143);
or U13955 (N_13955,N_11068,N_10127);
xor U13956 (N_13956,N_11190,N_11863);
nand U13957 (N_13957,N_10781,N_10523);
or U13958 (N_13958,N_11098,N_11211);
or U13959 (N_13959,N_11379,N_11055);
nand U13960 (N_13960,N_10666,N_11033);
nor U13961 (N_13961,N_11200,N_10934);
nand U13962 (N_13962,N_10719,N_11307);
nand U13963 (N_13963,N_11063,N_11183);
and U13964 (N_13964,N_10649,N_11132);
and U13965 (N_13965,N_11544,N_10363);
nor U13966 (N_13966,N_11451,N_10012);
nand U13967 (N_13967,N_10189,N_10399);
nand U13968 (N_13968,N_11560,N_10401);
and U13969 (N_13969,N_10377,N_11717);
nor U13970 (N_13970,N_10414,N_10641);
or U13971 (N_13971,N_11738,N_11267);
nor U13972 (N_13972,N_10981,N_11728);
or U13973 (N_13973,N_11703,N_10460);
nor U13974 (N_13974,N_10887,N_10924);
or U13975 (N_13975,N_11364,N_10569);
and U13976 (N_13976,N_11211,N_11898);
or U13977 (N_13977,N_10781,N_10459);
nor U13978 (N_13978,N_11311,N_10814);
xor U13979 (N_13979,N_11392,N_11951);
or U13980 (N_13980,N_10945,N_11192);
or U13981 (N_13981,N_11234,N_10727);
or U13982 (N_13982,N_11439,N_10019);
nand U13983 (N_13983,N_10444,N_10299);
or U13984 (N_13984,N_11345,N_10477);
xnor U13985 (N_13985,N_11310,N_10540);
nor U13986 (N_13986,N_10232,N_11435);
nor U13987 (N_13987,N_11632,N_11006);
nand U13988 (N_13988,N_10582,N_10278);
or U13989 (N_13989,N_10277,N_11454);
and U13990 (N_13990,N_10760,N_10563);
or U13991 (N_13991,N_11271,N_11467);
or U13992 (N_13992,N_11471,N_10454);
nand U13993 (N_13993,N_10521,N_10455);
or U13994 (N_13994,N_10136,N_11298);
or U13995 (N_13995,N_10689,N_10026);
nand U13996 (N_13996,N_10284,N_10676);
and U13997 (N_13997,N_11517,N_10567);
or U13998 (N_13998,N_10725,N_11975);
nor U13999 (N_13999,N_10156,N_10990);
or U14000 (N_14000,N_12649,N_12120);
or U14001 (N_14001,N_13106,N_13961);
nand U14002 (N_14002,N_12848,N_12043);
and U14003 (N_14003,N_12521,N_13341);
and U14004 (N_14004,N_12886,N_13173);
nand U14005 (N_14005,N_13814,N_12740);
or U14006 (N_14006,N_13286,N_13216);
xor U14007 (N_14007,N_12842,N_12541);
nor U14008 (N_14008,N_12709,N_12760);
xor U14009 (N_14009,N_13801,N_12482);
and U14010 (N_14010,N_12939,N_12602);
or U14011 (N_14011,N_12802,N_13530);
nand U14012 (N_14012,N_13969,N_13573);
nor U14013 (N_14013,N_13137,N_12394);
xnor U14014 (N_14014,N_12009,N_13214);
or U14015 (N_14015,N_12417,N_12107);
xor U14016 (N_14016,N_13670,N_13939);
xor U14017 (N_14017,N_13118,N_12458);
nor U14018 (N_14018,N_13056,N_13498);
nand U14019 (N_14019,N_13015,N_12500);
nand U14020 (N_14020,N_13626,N_12858);
nor U14021 (N_14021,N_12092,N_13171);
xor U14022 (N_14022,N_13743,N_12762);
or U14023 (N_14023,N_13692,N_12337);
and U14024 (N_14024,N_13955,N_12201);
nand U14025 (N_14025,N_12030,N_13684);
xnor U14026 (N_14026,N_12272,N_13985);
and U14027 (N_14027,N_13160,N_13889);
nor U14028 (N_14028,N_12639,N_12416);
and U14029 (N_14029,N_13415,N_13459);
nor U14030 (N_14030,N_12090,N_12140);
nand U14031 (N_14031,N_13510,N_12651);
and U14032 (N_14032,N_12827,N_12733);
xor U14033 (N_14033,N_12642,N_12840);
nand U14034 (N_14034,N_13629,N_13943);
or U14035 (N_14035,N_13824,N_13759);
or U14036 (N_14036,N_12369,N_13721);
nor U14037 (N_14037,N_13536,N_12803);
or U14038 (N_14038,N_13613,N_12495);
or U14039 (N_14039,N_13226,N_13689);
nand U14040 (N_14040,N_12245,N_12062);
xnor U14041 (N_14041,N_12446,N_13622);
or U14042 (N_14042,N_12868,N_13618);
xnor U14043 (N_14043,N_12817,N_12242);
or U14044 (N_14044,N_12470,N_13896);
nor U14045 (N_14045,N_13616,N_12979);
nor U14046 (N_14046,N_13558,N_13997);
and U14047 (N_14047,N_13846,N_12240);
or U14048 (N_14048,N_12927,N_12695);
nand U14049 (N_14049,N_13877,N_13856);
nand U14050 (N_14050,N_13931,N_13747);
nor U14051 (N_14051,N_12266,N_12471);
and U14052 (N_14052,N_13075,N_12662);
or U14053 (N_14053,N_12932,N_13835);
nor U14054 (N_14054,N_12924,N_12605);
xor U14055 (N_14055,N_12752,N_13054);
and U14056 (N_14056,N_13456,N_12040);
nand U14057 (N_14057,N_13474,N_12857);
xnor U14058 (N_14058,N_12851,N_12819);
and U14059 (N_14059,N_12168,N_12945);
or U14060 (N_14060,N_12061,N_12428);
nand U14061 (N_14061,N_13537,N_12192);
nor U14062 (N_14062,N_12688,N_12034);
or U14063 (N_14063,N_12408,N_12431);
or U14064 (N_14064,N_12419,N_12370);
nand U14065 (N_14065,N_13947,N_12130);
nor U14066 (N_14066,N_12320,N_13087);
or U14067 (N_14067,N_13201,N_12308);
or U14068 (N_14068,N_13076,N_12133);
and U14069 (N_14069,N_13957,N_13664);
xor U14070 (N_14070,N_12248,N_13061);
nand U14071 (N_14071,N_12583,N_12769);
nor U14072 (N_14072,N_13051,N_12497);
xnor U14073 (N_14073,N_12005,N_12493);
nor U14074 (N_14074,N_13387,N_13722);
and U14075 (N_14075,N_13928,N_12582);
xnor U14076 (N_14076,N_13332,N_13239);
nand U14077 (N_14077,N_12850,N_13577);
nor U14078 (N_14078,N_13775,N_13384);
nand U14079 (N_14079,N_13275,N_12671);
and U14080 (N_14080,N_12862,N_12866);
nand U14081 (N_14081,N_13739,N_12341);
nand U14082 (N_14082,N_12676,N_12435);
or U14083 (N_14083,N_13965,N_12164);
and U14084 (N_14084,N_13042,N_12813);
xor U14085 (N_14085,N_12852,N_13150);
or U14086 (N_14086,N_12312,N_12514);
xor U14087 (N_14087,N_12230,N_12468);
and U14088 (N_14088,N_12641,N_13967);
xnor U14089 (N_14089,N_12534,N_13126);
nand U14090 (N_14090,N_12089,N_13322);
nand U14091 (N_14091,N_13529,N_13060);
and U14092 (N_14092,N_12678,N_13110);
nand U14093 (N_14093,N_13027,N_12053);
and U14094 (N_14094,N_12954,N_12158);
or U14095 (N_14095,N_13477,N_13608);
nand U14096 (N_14096,N_13603,N_12413);
or U14097 (N_14097,N_13755,N_13496);
and U14098 (N_14098,N_12776,N_13047);
xor U14099 (N_14099,N_12455,N_13463);
nand U14100 (N_14100,N_12871,N_12375);
nor U14101 (N_14101,N_12667,N_12247);
or U14102 (N_14102,N_13866,N_13794);
xnor U14103 (N_14103,N_12045,N_13554);
nor U14104 (N_14104,N_12761,N_12047);
nor U14105 (N_14105,N_13521,N_12473);
and U14106 (N_14106,N_12981,N_13964);
and U14107 (N_14107,N_13590,N_13585);
nor U14108 (N_14108,N_12481,N_12820);
nand U14109 (N_14109,N_12147,N_13687);
and U14110 (N_14110,N_13612,N_12966);
nand U14111 (N_14111,N_12665,N_12148);
or U14112 (N_14112,N_13854,N_12211);
or U14113 (N_14113,N_12755,N_13649);
nand U14114 (N_14114,N_12388,N_12054);
nand U14115 (N_14115,N_12313,N_12552);
and U14116 (N_14116,N_12303,N_12281);
or U14117 (N_14117,N_12474,N_12747);
or U14118 (N_14118,N_13409,N_13881);
and U14119 (N_14119,N_12238,N_13340);
or U14120 (N_14120,N_12759,N_13669);
or U14121 (N_14121,N_13401,N_12773);
nand U14122 (N_14122,N_13520,N_13424);
xor U14123 (N_14123,N_13000,N_12186);
xor U14124 (N_14124,N_13502,N_13458);
xnor U14125 (N_14125,N_12578,N_12619);
nor U14126 (N_14126,N_13567,N_13806);
xor U14127 (N_14127,N_13091,N_12128);
nand U14128 (N_14128,N_13419,N_12905);
or U14129 (N_14129,N_13812,N_13528);
and U14130 (N_14130,N_12443,N_12208);
or U14131 (N_14131,N_13238,N_13615);
nor U14132 (N_14132,N_12854,N_12483);
and U14133 (N_14133,N_12228,N_13919);
or U14134 (N_14134,N_13768,N_12929);
and U14135 (N_14135,N_12793,N_12088);
nor U14136 (N_14136,N_13240,N_13952);
nand U14137 (N_14137,N_13548,N_12356);
and U14138 (N_14138,N_13431,N_13503);
or U14139 (N_14139,N_13904,N_12178);
or U14140 (N_14140,N_12690,N_12318);
nand U14141 (N_14141,N_12745,N_12349);
and U14142 (N_14142,N_12643,N_13819);
and U14143 (N_14143,N_13145,N_13190);
nand U14144 (N_14144,N_13080,N_13674);
nand U14145 (N_14145,N_13542,N_13705);
or U14146 (N_14146,N_13349,N_13380);
or U14147 (N_14147,N_13465,N_13187);
nor U14148 (N_14148,N_13915,N_12906);
nand U14149 (N_14149,N_12588,N_12718);
nor U14150 (N_14150,N_12908,N_13823);
and U14151 (N_14151,N_12461,N_12306);
nor U14152 (N_14152,N_12898,N_13324);
xnor U14153 (N_14153,N_13559,N_12996);
xor U14154 (N_14154,N_13072,N_12644);
xor U14155 (N_14155,N_12738,N_13936);
and U14156 (N_14156,N_13049,N_13423);
nor U14157 (N_14157,N_12322,N_12933);
and U14158 (N_14158,N_13836,N_13888);
or U14159 (N_14159,N_13641,N_12594);
nand U14160 (N_14160,N_12623,N_12251);
or U14161 (N_14161,N_12372,N_12576);
or U14162 (N_14162,N_12239,N_12877);
xor U14163 (N_14163,N_12606,N_13647);
nand U14164 (N_14164,N_13840,N_12300);
nand U14165 (N_14165,N_13976,N_12050);
and U14166 (N_14166,N_12173,N_13245);
xor U14167 (N_14167,N_12319,N_13081);
nor U14168 (N_14168,N_13271,N_13399);
or U14169 (N_14169,N_13476,N_13725);
nand U14170 (N_14170,N_12544,N_13645);
and U14171 (N_14171,N_12525,N_13307);
or U14172 (N_14172,N_12693,N_13442);
xor U14173 (N_14173,N_13086,N_13916);
nor U14174 (N_14174,N_13105,N_12444);
nand U14175 (N_14175,N_13313,N_12125);
or U14176 (N_14176,N_12859,N_12406);
nor U14177 (N_14177,N_13138,N_12340);
or U14178 (N_14178,N_13561,N_12007);
or U14179 (N_14179,N_12590,N_13578);
nor U14180 (N_14180,N_12343,N_12124);
or U14181 (N_14181,N_13695,N_13233);
nor U14182 (N_14182,N_12922,N_12687);
nand U14183 (N_14183,N_12589,N_13795);
and U14184 (N_14184,N_12450,N_12279);
or U14185 (N_14185,N_13259,N_12316);
xor U14186 (N_14186,N_13815,N_12537);
nand U14187 (N_14187,N_13164,N_12785);
or U14188 (N_14188,N_13129,N_13323);
or U14189 (N_14189,N_13434,N_13495);
or U14190 (N_14190,N_12824,N_13998);
xnor U14191 (N_14191,N_12392,N_13139);
or U14192 (N_14192,N_12305,N_13291);
or U14193 (N_14193,N_13913,N_13490);
xnor U14194 (N_14194,N_13041,N_12065);
or U14195 (N_14195,N_12104,N_13223);
xnor U14196 (N_14196,N_13925,N_13436);
nand U14197 (N_14197,N_13777,N_13065);
xnor U14198 (N_14198,N_12293,N_12520);
and U14199 (N_14199,N_13330,N_12501);
and U14200 (N_14200,N_13607,N_12599);
xor U14201 (N_14201,N_12256,N_13974);
nand U14202 (N_14202,N_13445,N_13638);
nand U14203 (N_14203,N_12015,N_12867);
xnor U14204 (N_14204,N_13175,N_13547);
nor U14205 (N_14205,N_12309,N_13365);
and U14206 (N_14206,N_13698,N_12921);
nand U14207 (N_14207,N_13588,N_13774);
xor U14208 (N_14208,N_12713,N_12162);
and U14209 (N_14209,N_13518,N_13215);
nand U14210 (N_14210,N_13780,N_12351);
and U14211 (N_14211,N_12097,N_13412);
or U14212 (N_14212,N_13299,N_13954);
and U14213 (N_14213,N_13809,N_13269);
xor U14214 (N_14214,N_13335,N_13370);
or U14215 (N_14215,N_12553,N_12347);
xnor U14216 (N_14216,N_12629,N_12911);
nand U14217 (N_14217,N_12951,N_13486);
or U14218 (N_14218,N_13772,N_12696);
or U14219 (N_14219,N_13543,N_13873);
and U14220 (N_14220,N_13298,N_12839);
and U14221 (N_14221,N_12568,N_13910);
nand U14222 (N_14222,N_13879,N_13994);
or U14223 (N_14223,N_13374,N_12847);
and U14224 (N_14224,N_12020,N_12650);
or U14225 (N_14225,N_13480,N_12071);
nand U14226 (N_14226,N_13094,N_13439);
nand U14227 (N_14227,N_12398,N_13099);
nand U14228 (N_14228,N_12253,N_13733);
and U14229 (N_14229,N_13200,N_13350);
xor U14230 (N_14230,N_12581,N_12961);
nor U14231 (N_14231,N_13485,N_12000);
nand U14232 (N_14232,N_13630,N_12113);
and U14233 (N_14233,N_12625,N_13760);
xor U14234 (N_14234,N_12660,N_12724);
nor U14235 (N_14235,N_13966,N_12818);
nand U14236 (N_14236,N_13932,N_12060);
nand U14237 (N_14237,N_12899,N_12485);
and U14238 (N_14238,N_12390,N_13037);
xnor U14239 (N_14239,N_13659,N_13123);
and U14240 (N_14240,N_12756,N_13472);
xor U14241 (N_14241,N_13662,N_12519);
xnor U14242 (N_14242,N_13753,N_13198);
nand U14243 (N_14243,N_12527,N_12902);
and U14244 (N_14244,N_13539,N_13451);
xor U14245 (N_14245,N_12700,N_13863);
nor U14246 (N_14246,N_12325,N_13709);
xnor U14247 (N_14247,N_12551,N_12466);
and U14248 (N_14248,N_13209,N_13508);
nand U14249 (N_14249,N_12214,N_13688);
nand U14250 (N_14250,N_12442,N_12571);
nor U14251 (N_14251,N_13610,N_13851);
or U14252 (N_14252,N_12975,N_12462);
nor U14253 (N_14253,N_12365,N_12310);
and U14254 (N_14254,N_13277,N_13992);
xnor U14255 (N_14255,N_13852,N_13107);
and U14256 (N_14256,N_12901,N_12704);
and U14257 (N_14257,N_13842,N_13410);
nand U14258 (N_14258,N_12560,N_13191);
xor U14259 (N_14259,N_13923,N_12679);
nand U14260 (N_14260,N_12804,N_12286);
xor U14261 (N_14261,N_13611,N_12895);
or U14262 (N_14262,N_12295,N_13908);
or U14263 (N_14263,N_13716,N_12670);
nand U14264 (N_14264,N_13734,N_13584);
nand U14265 (N_14265,N_13276,N_13407);
and U14266 (N_14266,N_13433,N_12993);
or U14267 (N_14267,N_13749,N_13386);
or U14268 (N_14268,N_12692,N_12331);
xnor U14269 (N_14269,N_12056,N_12283);
or U14270 (N_14270,N_13926,N_13135);
nor U14271 (N_14271,N_13295,N_13728);
nand U14272 (N_14272,N_12064,N_13235);
or U14273 (N_14273,N_12430,N_13142);
or U14274 (N_14274,N_13726,N_13229);
and U14275 (N_14275,N_12685,N_13044);
nor U14276 (N_14276,N_12216,N_13596);
xor U14277 (N_14277,N_12779,N_12978);
xnor U14278 (N_14278,N_13132,N_12913);
nand U14279 (N_14279,N_13951,N_13345);
nand U14280 (N_14280,N_12159,N_13461);
or U14281 (N_14281,N_12965,N_13673);
xor U14282 (N_14282,N_12962,N_13564);
or U14283 (N_14283,N_12114,N_12539);
nand U14284 (N_14284,N_12093,N_12983);
or U14285 (N_14285,N_13064,N_13179);
nor U14286 (N_14286,N_12952,N_12875);
and U14287 (N_14287,N_13421,N_13392);
nor U14288 (N_14288,N_12410,N_13297);
nor U14289 (N_14289,N_13406,N_12845);
and U14290 (N_14290,N_12421,N_13071);
or U14291 (N_14291,N_13222,N_13019);
or U14292 (N_14292,N_12066,N_12480);
or U14293 (N_14293,N_12658,N_13720);
or U14294 (N_14294,N_12476,N_13898);
nand U14295 (N_14295,N_12330,N_12972);
xnor U14296 (N_14296,N_12035,N_13282);
and U14297 (N_14297,N_13002,N_12735);
xnor U14298 (N_14298,N_13601,N_12275);
or U14299 (N_14299,N_13515,N_13319);
and U14300 (N_14300,N_12730,N_13111);
nor U14301 (N_14301,N_12668,N_13327);
and U14302 (N_14302,N_13970,N_13804);
nand U14303 (N_14303,N_13635,N_13422);
or U14304 (N_14304,N_13217,N_13752);
or U14305 (N_14305,N_13162,N_12765);
and U14306 (N_14306,N_13029,N_13632);
or U14307 (N_14307,N_12167,N_12105);
xor U14308 (N_14308,N_12255,N_13792);
nor U14309 (N_14309,N_13012,N_12563);
nand U14310 (N_14310,N_13304,N_13468);
or U14311 (N_14311,N_13991,N_13252);
and U14312 (N_14312,N_12049,N_12812);
or U14313 (N_14313,N_12076,N_12073);
xor U14314 (N_14314,N_12094,N_13121);
and U14315 (N_14315,N_13545,N_13154);
or U14316 (N_14316,N_12108,N_12452);
and U14317 (N_14317,N_12948,N_12223);
xor U14318 (N_14318,N_13575,N_12106);
nand U14319 (N_14319,N_13911,N_13152);
or U14320 (N_14320,N_13972,N_12411);
and U14321 (N_14321,N_13599,N_13131);
or U14322 (N_14322,N_13742,N_13724);
xnor U14323 (N_14323,N_13225,N_13651);
nand U14324 (N_14324,N_12134,N_13156);
xor U14325 (N_14325,N_12736,N_12327);
or U14326 (N_14326,N_12456,N_12420);
nor U14327 (N_14327,N_12226,N_12418);
nand U14328 (N_14328,N_12155,N_12666);
and U14329 (N_14329,N_13292,N_12002);
and U14330 (N_14330,N_12467,N_12753);
nor U14331 (N_14331,N_13837,N_12973);
or U14332 (N_14332,N_13874,N_12004);
and U14333 (N_14333,N_12930,N_12522);
and U14334 (N_14334,N_13628,N_12652);
xnor U14335 (N_14335,N_13803,N_13623);
nor U14336 (N_14336,N_12722,N_12373);
and U14337 (N_14337,N_12870,N_13924);
and U14338 (N_14338,N_12259,N_13268);
nand U14339 (N_14339,N_13074,N_13540);
or U14340 (N_14340,N_12654,N_13023);
or U14341 (N_14341,N_13427,N_12119);
and U14342 (N_14342,N_12987,N_13203);
or U14343 (N_14343,N_13978,N_12741);
nand U14344 (N_14344,N_12160,N_13580);
nand U14345 (N_14345,N_12032,N_12788);
nor U14346 (N_14346,N_12326,N_12919);
and U14347 (N_14347,N_12021,N_12821);
and U14348 (N_14348,N_12669,N_13813);
and U14349 (N_14349,N_13713,N_13982);
or U14350 (N_14350,N_12250,N_12379);
nand U14351 (N_14351,N_13859,N_13971);
and U14352 (N_14352,N_12604,N_13241);
or U14353 (N_14353,N_13507,N_12451);
or U14354 (N_14354,N_12241,N_13642);
nand U14355 (N_14355,N_12109,N_13557);
or U14356 (N_14356,N_13115,N_13098);
xnor U14357 (N_14357,N_12796,N_13050);
nand U14358 (N_14358,N_13796,N_13211);
xor U14359 (N_14359,N_12491,N_13650);
xor U14360 (N_14360,N_12346,N_12194);
or U14361 (N_14361,N_13586,N_13085);
nor U14362 (N_14362,N_13184,N_12013);
and U14363 (N_14363,N_12511,N_12082);
nand U14364 (N_14364,N_12081,N_13244);
and U14365 (N_14365,N_12332,N_13127);
and U14366 (N_14366,N_13784,N_12424);
nand U14367 (N_14367,N_13597,N_13331);
nor U14368 (N_14368,N_13999,N_13668);
xor U14369 (N_14369,N_12145,N_12403);
nor U14370 (N_14370,N_13619,N_12206);
nand U14371 (N_14371,N_12797,N_12663);
nor U14372 (N_14372,N_12529,N_13799);
or U14373 (N_14373,N_13761,N_12396);
xor U14374 (N_14374,N_13769,N_12548);
xor U14375 (N_14375,N_13306,N_13736);
xor U14376 (N_14376,N_12810,N_13989);
nand U14377 (N_14377,N_12798,N_13026);
nand U14378 (N_14378,N_13302,N_12748);
or U14379 (N_14379,N_12041,N_12976);
xor U14380 (N_14380,N_13254,N_13308);
nor U14381 (N_14381,N_12187,N_12790);
and U14382 (N_14382,N_12878,N_12823);
nor U14383 (N_14383,N_12661,N_12448);
nand U14384 (N_14384,N_12907,N_13287);
nand U14385 (N_14385,N_12277,N_12433);
nand U14386 (N_14386,N_13416,N_13776);
or U14387 (N_14387,N_13188,N_13555);
nor U14388 (N_14388,N_13544,N_12807);
nand U14389 (N_14389,N_12874,N_12195);
xor U14390 (N_14390,N_13155,N_13614);
or U14391 (N_14391,N_12737,N_12397);
or U14392 (N_14392,N_12533,N_12103);
xnor U14393 (N_14393,N_13828,N_13918);
nor U14394 (N_14394,N_13031,N_13165);
nor U14395 (N_14395,N_12982,N_12405);
or U14396 (N_14396,N_13182,N_12564);
and U14397 (N_14397,N_13046,N_13646);
or U14398 (N_14398,N_12774,N_12570);
or U14399 (N_14399,N_13832,N_12352);
or U14400 (N_14400,N_12731,N_12296);
and U14401 (N_14401,N_12361,N_13260);
nand U14402 (N_14402,N_13210,N_13605);
nor U14403 (N_14403,N_12787,N_13730);
nand U14404 (N_14404,N_12946,N_12717);
or U14405 (N_14405,N_13283,N_13218);
xnor U14406 (N_14406,N_13653,N_12699);
nor U14407 (N_14407,N_12573,N_12229);
xnor U14408 (N_14408,N_12152,N_12014);
xnor U14409 (N_14409,N_13893,N_12287);
nand U14410 (N_14410,N_13849,N_12083);
nand U14411 (N_14411,N_13378,N_13945);
or U14412 (N_14412,N_12706,N_13021);
and U14413 (N_14413,N_13870,N_12540);
or U14414 (N_14414,N_13983,N_13746);
nor U14415 (N_14415,N_13839,N_13426);
xor U14416 (N_14416,N_13617,N_12989);
xnor U14417 (N_14417,N_12879,N_13853);
xor U14418 (N_14418,N_13694,N_12958);
and U14419 (N_14419,N_13883,N_12267);
or U14420 (N_14420,N_12855,N_12550);
nor U14421 (N_14421,N_13379,N_13574);
and U14422 (N_14422,N_12472,N_13073);
or U14423 (N_14423,N_12243,N_12236);
nand U14424 (N_14424,N_12301,N_12626);
nor U14425 (N_14425,N_12486,N_13572);
nand U14426 (N_14426,N_12861,N_12338);
xor U14427 (N_14427,N_13373,N_13243);
or U14428 (N_14428,N_12115,N_12044);
nor U14429 (N_14429,N_12630,N_13811);
and U14430 (N_14430,N_12401,N_13320);
nand U14431 (N_14431,N_12118,N_13643);
nand U14432 (N_14432,N_13360,N_13903);
nand U14433 (N_14433,N_13258,N_13741);
and U14434 (N_14434,N_12531,N_12555);
nor U14435 (N_14435,N_13062,N_13827);
or U14436 (N_14436,N_12575,N_13602);
xnor U14437 (N_14437,N_13942,N_12077);
or U14438 (N_14438,N_12136,N_13718);
xor U14439 (N_14439,N_12172,N_12117);
nand U14440 (N_14440,N_13337,N_12734);
nor U14441 (N_14441,N_13533,N_13489);
nor U14442 (N_14442,N_13334,N_13764);
nor U14443 (N_14443,N_13861,N_12637);
and U14444 (N_14444,N_13354,N_12789);
nand U14445 (N_14445,N_13375,N_13822);
nand U14446 (N_14446,N_12684,N_12648);
and U14447 (N_14447,N_12366,N_13563);
or U14448 (N_14448,N_12767,N_12628);
and U14449 (N_14449,N_12615,N_13467);
xnor U14450 (N_14450,N_13083,N_13512);
and U14451 (N_14451,N_12903,N_12012);
nand U14452 (N_14452,N_12166,N_12387);
xor U14453 (N_14453,N_12068,N_12768);
and U14454 (N_14454,N_13070,N_12404);
nand U14455 (N_14455,N_12900,N_12121);
and U14456 (N_14456,N_13587,N_13147);
and U14457 (N_14457,N_12607,N_13478);
xnor U14458 (N_14458,N_13686,N_12188);
and U14459 (N_14459,N_13862,N_12333);
nor U14460 (N_14460,N_13569,N_13591);
or U14461 (N_14461,N_12196,N_12725);
nor U14462 (N_14462,N_12059,N_13285);
or U14463 (N_14463,N_12139,N_12783);
and U14464 (N_14464,N_12191,N_13312);
xnor U14465 (N_14465,N_13680,N_13977);
xnor U14466 (N_14466,N_13473,N_12273);
xnor U14467 (N_14467,N_13634,N_12890);
nor U14468 (N_14468,N_12940,N_12750);
nor U14469 (N_14469,N_13927,N_13033);
and U14470 (N_14470,N_12834,N_13600);
xor U14471 (N_14471,N_13036,N_13788);
and U14472 (N_14472,N_12008,N_12227);
nor U14473 (N_14473,N_12910,N_12942);
or U14474 (N_14474,N_12509,N_12438);
nor U14475 (N_14475,N_12042,N_13956);
xnor U14476 (N_14476,N_13579,N_13882);
nor U14477 (N_14477,N_13711,N_13273);
nand U14478 (N_14478,N_13114,N_12632);
nor U14479 (N_14479,N_12806,N_13385);
and U14480 (N_14480,N_13592,N_12585);
nand U14481 (N_14481,N_12697,N_13935);
and U14482 (N_14482,N_12686,N_13336);
or U14483 (N_14483,N_13797,N_13946);
or U14484 (N_14484,N_12393,N_13782);
or U14485 (N_14485,N_12749,N_13493);
or U14486 (N_14486,N_13937,N_13344);
and U14487 (N_14487,N_12367,N_13805);
xor U14488 (N_14488,N_13348,N_13250);
nand U14489 (N_14489,N_13063,N_12084);
nand U14490 (N_14490,N_12538,N_12532);
or U14491 (N_14491,N_12453,N_13356);
and U14492 (N_14492,N_12381,N_13606);
and U14493 (N_14493,N_13017,N_13527);
nand U14494 (N_14494,N_12364,N_12934);
nand U14495 (N_14495,N_13040,N_13719);
nand U14496 (N_14496,N_13194,N_13134);
nor U14497 (N_14497,N_13737,N_12865);
nand U14498 (N_14498,N_12881,N_13161);
nand U14499 (N_14499,N_13693,N_12197);
xor U14500 (N_14500,N_12781,N_13690);
nand U14501 (N_14501,N_12825,N_13255);
or U14502 (N_14502,N_12317,N_12204);
or U14503 (N_14503,N_12307,N_13003);
nor U14504 (N_14504,N_13857,N_12153);
nand U14505 (N_14505,N_13594,N_12218);
xnor U14506 (N_14506,N_13363,N_13627);
or U14507 (N_14507,N_13487,N_13583);
or U14508 (N_14508,N_12677,N_12869);
or U14509 (N_14509,N_12572,N_13949);
and U14510 (N_14510,N_13466,N_12489);
xor U14511 (N_14511,N_13876,N_13878);
and U14512 (N_14512,N_13895,N_12732);
nand U14513 (N_14513,N_12828,N_13314);
or U14514 (N_14514,N_12627,N_12328);
or U14515 (N_14515,N_12199,N_13035);
nand U14516 (N_14516,N_12673,N_12918);
nor U14517 (N_14517,N_12098,N_13248);
nand U14518 (N_14518,N_13220,N_12284);
nor U14519 (N_14519,N_13231,N_12885);
nor U14520 (N_14520,N_13082,N_12095);
and U14521 (N_14521,N_12617,N_12502);
nand U14522 (N_14522,N_12914,N_12131);
and U14523 (N_14523,N_12778,N_13025);
nand U14524 (N_14524,N_13671,N_12888);
xor U14525 (N_14525,N_13745,N_13499);
xnor U14526 (N_14526,N_12503,N_12180);
xor U14527 (N_14527,N_12138,N_12546);
nor U14528 (N_14528,N_13206,N_13868);
or U14529 (N_14529,N_12031,N_13408);
nor U14530 (N_14530,N_12782,N_13010);
or U14531 (N_14531,N_12833,N_13428);
or U14532 (N_14532,N_12549,N_13552);
nand U14533 (N_14533,N_13701,N_13168);
nand U14534 (N_14534,N_12892,N_12079);
or U14535 (N_14535,N_13084,N_13352);
nor U14536 (N_14536,N_12512,N_13435);
nand U14537 (N_14537,N_12383,N_13368);
or U14538 (N_14538,N_13169,N_12183);
nor U14539 (N_14539,N_13395,N_12184);
xnor U14540 (N_14540,N_12708,N_13202);
and U14541 (N_14541,N_13289,N_12955);
or U14542 (N_14542,N_13186,N_12947);
xnor U14543 (N_14543,N_12758,N_13855);
nor U14544 (N_14544,N_12610,N_12382);
or U14545 (N_14545,N_12574,N_13020);
or U14546 (N_14546,N_13128,N_13704);
xor U14547 (N_14547,N_12252,N_13933);
nor U14548 (N_14548,N_12436,N_12634);
xor U14549 (N_14549,N_13310,N_13143);
or U14550 (N_14550,N_12355,N_12786);
and U14551 (N_14551,N_12872,N_12179);
xor U14552 (N_14552,N_12498,N_13549);
or U14553 (N_14553,N_13800,N_13818);
or U14554 (N_14554,N_12335,N_12915);
xnor U14555 (N_14555,N_13364,N_12176);
and U14556 (N_14556,N_13667,N_13270);
xor U14557 (N_14557,N_13714,N_13024);
xnor U14558 (N_14558,N_13938,N_13479);
xor U14559 (N_14559,N_13383,N_12526);
xnor U14560 (N_14560,N_12321,N_13183);
and U14561 (N_14561,N_13325,N_12175);
and U14562 (N_14562,N_12800,N_12920);
or U14563 (N_14563,N_12377,N_13712);
xnor U14564 (N_14564,N_13078,N_12635);
and U14565 (N_14565,N_13462,N_12350);
and U14566 (N_14566,N_12809,N_12883);
xnor U14567 (N_14567,N_12799,N_13867);
xnor U14568 (N_14568,N_13798,N_13717);
and U14569 (N_14569,N_13117,N_13506);
nand U14570 (N_14570,N_12507,N_13771);
nand U14571 (N_14571,N_12757,N_13192);
or U14572 (N_14572,N_13962,N_13766);
and U14573 (N_14573,N_12716,N_12297);
or U14574 (N_14574,N_12754,N_12051);
or U14575 (N_14575,N_13281,N_13525);
and U14576 (N_14576,N_13140,N_13864);
and U14577 (N_14577,N_12944,N_13727);
xnor U14578 (N_14578,N_13052,N_12067);
and U14579 (N_14579,N_13494,N_13326);
or U14580 (N_14580,N_12510,N_12096);
nor U14581 (N_14581,N_13232,N_12990);
xor U14582 (N_14582,N_12215,N_12763);
xor U14583 (N_14583,N_13683,N_12659);
nand U14584 (N_14584,N_13816,N_12579);
nand U14585 (N_14585,N_12202,N_13279);
xnor U14586 (N_14586,N_13089,N_12477);
nor U14587 (N_14587,N_13001,N_12189);
or U14588 (N_14588,N_13751,N_12791);
or U14589 (N_14589,N_12530,N_13300);
nor U14590 (N_14590,N_13589,N_13095);
nor U14591 (N_14591,N_12425,N_12298);
nor U14592 (N_14592,N_12161,N_13940);
and U14593 (N_14593,N_13030,N_13892);
xnor U14594 (N_14594,N_12876,N_12329);
or U14595 (N_14595,N_13361,N_12235);
or U14596 (N_14596,N_13754,N_12033);
nor U14597 (N_14597,N_13894,N_12423);
nand U14598 (N_14598,N_13691,N_12407);
nor U14599 (N_14599,N_13660,N_13675);
nand U14600 (N_14600,N_13700,N_12943);
xor U14601 (N_14601,N_12516,N_13055);
nand U14602 (N_14602,N_12282,N_13224);
xor U14603 (N_14603,N_13909,N_12395);
nor U14604 (N_14604,N_12101,N_13566);
nand U14605 (N_14605,N_12728,N_13256);
nor U14606 (N_14606,N_13517,N_12566);
nor U14607 (N_14607,N_12909,N_13672);
nor U14608 (N_14608,N_13820,N_13347);
nor U14609 (N_14609,N_12505,N_13912);
and U14610 (N_14610,N_13261,N_12655);
nor U14611 (N_14611,N_12640,N_13457);
or U14612 (N_14612,N_12624,N_13393);
xor U14613 (N_14613,N_13130,N_13390);
nand U14614 (N_14614,N_13362,N_13090);
and U14615 (N_14615,N_12440,N_12811);
or U14616 (N_14616,N_13891,N_12938);
xnor U14617 (N_14617,N_13656,N_12400);
and U14618 (N_14618,N_12841,N_12746);
and U14619 (N_14619,N_12036,N_13438);
nor U14620 (N_14620,N_13262,N_12265);
and U14621 (N_14621,N_12249,N_12132);
xnor U14622 (N_14622,N_12949,N_13397);
nor U14623 (N_14623,N_12710,N_13034);
xor U14624 (N_14624,N_13413,N_12638);
nor U14625 (N_14625,N_13550,N_12702);
and U14626 (N_14626,N_12339,N_12344);
or U14627 (N_14627,N_12441,N_13011);
xnor U14628 (N_14628,N_13185,N_13405);
or U14629 (N_14629,N_13221,N_12058);
xnor U14630 (N_14630,N_13620,N_13731);
nor U14631 (N_14631,N_12234,N_12646);
nor U14632 (N_14632,N_12151,N_12645);
and U14633 (N_14633,N_12302,N_12985);
nor U14634 (N_14634,N_12142,N_13346);
nor U14635 (N_14635,N_12986,N_13914);
and U14636 (N_14636,N_13885,N_13920);
xnor U14637 (N_14637,N_13979,N_12620);
xor U14638 (N_14638,N_12657,N_12099);
nor U14639 (N_14639,N_12837,N_13501);
nand U14640 (N_14640,N_13167,N_13018);
xnor U14641 (N_14641,N_13471,N_13236);
or U14642 (N_14642,N_13865,N_13100);
nor U14643 (N_14643,N_13988,N_13633);
and U14644 (N_14644,N_12931,N_13833);
xnor U14645 (N_14645,N_13699,N_12729);
xnor U14646 (N_14646,N_12998,N_12792);
nor U14647 (N_14647,N_13355,N_12856);
xnor U14648 (N_14648,N_13560,N_12680);
nor U14649 (N_14649,N_13987,N_12360);
and U14650 (N_14650,N_13391,N_12742);
nand U14651 (N_14651,N_12714,N_13959);
xor U14652 (N_14652,N_13290,N_13343);
xor U14653 (N_14653,N_12743,N_12011);
and U14654 (N_14654,N_13163,N_12006);
xor U14655 (N_14655,N_13593,N_12672);
nand U14656 (N_14656,N_12126,N_12304);
or U14657 (N_14657,N_12488,N_13196);
and U14658 (N_14658,N_12621,N_13980);
and U14659 (N_14659,N_13516,N_12830);
xnor U14660 (N_14660,N_13257,N_13884);
xor U14661 (N_14661,N_13568,N_13102);
nor U14662 (N_14662,N_12916,N_12535);
and U14663 (N_14663,N_13204,N_12912);
or U14664 (N_14664,N_13316,N_13120);
or U14665 (N_14665,N_13595,N_12936);
nor U14666 (N_14666,N_12554,N_13381);
and U14667 (N_14667,N_12542,N_13661);
nand U14668 (N_14668,N_13016,N_13522);
nand U14669 (N_14669,N_13789,N_13875);
nor U14670 (N_14670,N_13990,N_12691);
and U14671 (N_14671,N_13901,N_12917);
or U14672 (N_14672,N_13708,N_12891);
nor U14673 (N_14673,N_13958,N_12977);
or U14674 (N_14674,N_13723,N_13443);
nor U14675 (N_14675,N_13318,N_13382);
and U14676 (N_14676,N_12795,N_12558);
nor U14677 (N_14677,N_12721,N_13103);
nor U14678 (N_14678,N_12508,N_13144);
nor U14679 (N_14679,N_12023,N_12225);
nand U14680 (N_14680,N_13872,N_12289);
and U14681 (N_14681,N_13570,N_12720);
or U14682 (N_14682,N_12263,N_13750);
nand U14683 (N_14683,N_13059,N_12210);
nand U14684 (N_14684,N_12941,N_12018);
nor U14685 (N_14685,N_12490,N_12597);
or U14686 (N_14686,N_12603,N_13237);
xnor U14687 (N_14687,N_13781,N_13367);
nor U14688 (N_14688,N_12376,N_13097);
and U14689 (N_14689,N_13763,N_13008);
and U14690 (N_14690,N_12739,N_12601);
nand U14691 (N_14691,N_13009,N_12950);
xor U14692 (N_14692,N_12280,N_13571);
nand U14693 (N_14693,N_12523,N_12496);
and U14694 (N_14694,N_13500,N_13133);
xor U14695 (N_14695,N_13732,N_12016);
xor U14696 (N_14696,N_13174,N_12292);
xor U14697 (N_14697,N_12999,N_12592);
or U14698 (N_14698,N_12291,N_12141);
or U14699 (N_14699,N_12971,N_12386);
nand U14700 (N_14700,N_12726,N_13677);
and U14701 (N_14701,N_13902,N_12478);
nand U14702 (N_14702,N_13598,N_12299);
nor U14703 (N_14703,N_13230,N_12027);
nand U14704 (N_14704,N_13821,N_12294);
and U14705 (N_14705,N_13624,N_12371);
or U14706 (N_14706,N_13265,N_12561);
xnor U14707 (N_14707,N_12969,N_12780);
and U14708 (N_14708,N_12244,N_13484);
nand U14709 (N_14709,N_12233,N_13411);
and U14710 (N_14710,N_12359,N_13897);
or U14711 (N_14711,N_13715,N_13066);
nor U14712 (N_14712,N_12213,N_13351);
or U14713 (N_14713,N_13249,N_12037);
nand U14714 (N_14714,N_13511,N_12681);
xnor U14715 (N_14715,N_13278,N_13141);
xnor U14716 (N_14716,N_12715,N_13665);
nor U14717 (N_14717,N_13305,N_12463);
nand U14718 (N_14718,N_13838,N_12135);
or U14719 (N_14719,N_12518,N_13475);
nor U14720 (N_14720,N_13359,N_13841);
xor U14721 (N_14721,N_13565,N_12209);
or U14722 (N_14722,N_12380,N_13470);
and U14723 (N_14723,N_13513,N_13786);
xnor U14724 (N_14724,N_12384,N_12577);
nand U14725 (N_14725,N_12469,N_13829);
xnor U14726 (N_14726,N_12698,N_12038);
or U14727 (N_14727,N_13639,N_12559);
and U14728 (N_14728,N_13272,N_12254);
xnor U14729 (N_14729,N_13284,N_13984);
xor U14730 (N_14730,N_12712,N_13358);
nor U14731 (N_14731,N_13039,N_13398);
nand U14732 (N_14732,N_13464,N_13696);
nor U14733 (N_14733,N_13871,N_13826);
xor U14734 (N_14734,N_12111,N_13043);
nand U14735 (N_14735,N_13482,N_12935);
nor U14736 (N_14736,N_12426,N_12290);
or U14737 (N_14737,N_13644,N_13122);
and U14738 (N_14738,N_12409,N_13779);
and U14739 (N_14739,N_12271,N_13905);
and U14740 (N_14740,N_13817,N_12353);
xor U14741 (N_14741,N_12207,N_12631);
xnor U14742 (N_14742,N_12402,N_12072);
xnor U14743 (N_14743,N_13850,N_13453);
xor U14744 (N_14744,N_12464,N_12853);
nand U14745 (N_14745,N_13157,N_13625);
or U14746 (N_14746,N_13679,N_12169);
or U14747 (N_14747,N_12960,N_13890);
nand U14748 (N_14748,N_13038,N_12766);
and U14749 (N_14749,N_13553,N_13729);
nand U14750 (N_14750,N_12001,N_12222);
or U14751 (N_14751,N_13783,N_13440);
nor U14752 (N_14752,N_12070,N_13930);
nand U14753 (N_14753,N_13844,N_12689);
or U14754 (N_14754,N_12957,N_12956);
nand U14755 (N_14755,N_13296,N_12459);
nand U14756 (N_14756,N_12843,N_12220);
or U14757 (N_14757,N_13953,N_13551);
nand U14758 (N_14758,N_12288,N_12653);
or U14759 (N_14759,N_13420,N_12063);
xnor U14760 (N_14760,N_13005,N_13756);
nand U14761 (N_14761,N_12028,N_13013);
and U14762 (N_14762,N_12224,N_12844);
nor U14763 (N_14763,N_12612,N_12026);
or U14764 (N_14764,N_13636,N_12719);
xor U14765 (N_14765,N_12024,N_13267);
xnor U14766 (N_14766,N_12633,N_13088);
and U14767 (N_14767,N_12897,N_13069);
xnor U14768 (N_14768,N_13685,N_13514);
xnor U14769 (N_14769,N_12046,N_13096);
nor U14770 (N_14770,N_12591,N_12814);
nor U14771 (N_14771,N_13710,N_12595);
xnor U14772 (N_14772,N_12143,N_13178);
nor U14773 (N_14773,N_12494,N_13032);
xnor U14774 (N_14774,N_12723,N_13648);
nand U14775 (N_14775,N_13417,N_12880);
nand U14776 (N_14776,N_12057,N_12334);
and U14777 (N_14777,N_12744,N_13830);
and U14778 (N_14778,N_13197,N_13993);
or U14779 (N_14779,N_12751,N_13077);
and U14780 (N_14780,N_12517,N_13880);
nor U14781 (N_14781,N_12772,N_13113);
nor U14782 (N_14782,N_12270,N_12080);
nand U14783 (N_14783,N_12988,N_13251);
or U14784 (N_14784,N_12593,N_12893);
xnor U14785 (N_14785,N_12991,N_13372);
or U14786 (N_14786,N_13125,N_12378);
and U14787 (N_14787,N_12150,N_13227);
nand U14788 (N_14788,N_13253,N_12039);
xnor U14789 (N_14789,N_13303,N_12524);
or U14790 (N_14790,N_13758,N_12029);
nor U14791 (N_14791,N_12110,N_13452);
xor U14792 (N_14792,N_12596,N_13329);
and U14793 (N_14793,N_13917,N_13455);
nand U14794 (N_14794,N_13654,N_13681);
xnor U14795 (N_14795,N_13481,N_13948);
and U14796 (N_14796,N_12826,N_12181);
nand U14797 (N_14797,N_12177,N_13981);
nor U14798 (N_14798,N_13315,N_12565);
nor U14799 (N_14799,N_13153,N_12260);
nor U14800 (N_14800,N_13793,N_13582);
xnor U14801 (N_14801,N_12664,N_12219);
nor U14802 (N_14802,N_12232,N_13429);
nand U14803 (N_14803,N_13609,N_13447);
nor U14804 (N_14804,N_13843,N_12953);
nor U14805 (N_14805,N_13941,N_13621);
xnor U14806 (N_14806,N_13787,N_13400);
or U14807 (N_14807,N_12163,N_13491);
xor U14808 (N_14808,N_13524,N_13228);
xor U14809 (N_14809,N_12904,N_13488);
nand U14810 (N_14810,N_13509,N_12261);
nor U14811 (N_14811,N_13007,N_12445);
or U14812 (N_14812,N_12703,N_13177);
nor U14813 (N_14813,N_13022,N_13604);
or U14814 (N_14814,N_12925,N_13492);
nor U14815 (N_14815,N_13556,N_13280);
and U14816 (N_14816,N_13425,N_13151);
xor U14817 (N_14817,N_13309,N_12622);
nor U14818 (N_14818,N_12616,N_12285);
nand U14819 (N_14819,N_13234,N_12562);
nor U14820 (N_14820,N_12368,N_13311);
nor U14821 (N_14821,N_13791,N_12984);
nand U14822 (N_14822,N_13834,N_13389);
and U14823 (N_14823,N_13048,N_12357);
nand U14824 (N_14824,N_12970,N_12129);
and U14825 (N_14825,N_12432,N_12314);
or U14826 (N_14826,N_13166,N_13531);
nand U14827 (N_14827,N_13907,N_13808);
or U14828 (N_14828,N_12217,N_12479);
nand U14829 (N_14829,N_13657,N_12315);
nand U14830 (N_14830,N_12831,N_12048);
and U14831 (N_14831,N_12543,N_12091);
and U14832 (N_14832,N_13944,N_12203);
xnor U14833 (N_14833,N_12995,N_13195);
and U14834 (N_14834,N_13450,N_12580);
xnor U14835 (N_14835,N_12454,N_12873);
nand U14836 (N_14836,N_12269,N_12701);
or U14837 (N_14837,N_13274,N_13454);
xnor U14838 (N_14838,N_13172,N_13353);
and U14839 (N_14839,N_13666,N_13193);
nor U14840 (N_14840,N_12967,N_13676);
and U14841 (N_14841,N_12515,N_12484);
nand U14842 (N_14842,N_13678,N_12074);
and U14843 (N_14843,N_13176,N_13294);
xor U14844 (N_14844,N_13469,N_12816);
xnor U14845 (N_14845,N_12075,N_13929);
nor U14846 (N_14846,N_12808,N_12707);
xnor U14847 (N_14847,N_12959,N_13785);
and U14848 (N_14848,N_12156,N_13158);
nor U14849 (N_14849,N_12727,N_13067);
nand U14850 (N_14850,N_12087,N_13170);
or U14851 (N_14851,N_12504,N_12598);
xnor U14852 (N_14852,N_12078,N_12586);
or U14853 (N_14853,N_13869,N_12569);
or U14854 (N_14854,N_12429,N_13053);
xnor U14855 (N_14855,N_12584,N_12613);
xor U14856 (N_14856,N_12182,N_12846);
nor U14857 (N_14857,N_12711,N_13212);
or U14858 (N_14858,N_13181,N_12427);
nor U14859 (N_14859,N_12887,N_12487);
nor U14860 (N_14860,N_13887,N_12122);
and U14861 (N_14861,N_12964,N_13321);
nand U14862 (N_14862,N_12968,N_13847);
or U14863 (N_14863,N_13339,N_13921);
nand U14864 (N_14864,N_13986,N_12513);
or U14865 (N_14865,N_13748,N_12889);
and U14866 (N_14866,N_12449,N_13109);
nor U14867 (N_14867,N_12447,N_12149);
nand U14868 (N_14868,N_12771,N_13207);
nor U14869 (N_14869,N_12278,N_13006);
and U14870 (N_14870,N_13706,N_12980);
nand U14871 (N_14871,N_12439,N_12205);
and U14872 (N_14872,N_13333,N_13404);
nor U14873 (N_14873,N_12146,N_12414);
xnor U14874 (N_14874,N_13004,N_12614);
xor U14875 (N_14875,N_12055,N_12465);
nand U14876 (N_14876,N_12545,N_12896);
xor U14877 (N_14877,N_12237,N_12069);
nor U14878 (N_14878,N_13652,N_12587);
nor U14879 (N_14879,N_13448,N_13860);
and U14880 (N_14880,N_12102,N_13414);
and U14881 (N_14881,N_13963,N_12832);
nand U14882 (N_14882,N_13922,N_12611);
or U14883 (N_14883,N_12262,N_12674);
nor U14884 (N_14884,N_13658,N_13112);
nand U14885 (N_14885,N_13697,N_12608);
nor U14886 (N_14886,N_12770,N_12835);
xnor U14887 (N_14887,N_12258,N_13079);
and U14888 (N_14888,N_13058,N_12116);
or U14889 (N_14889,N_12025,N_13403);
nand U14890 (N_14890,N_13328,N_12085);
nor U14891 (N_14891,N_12600,N_13845);
or U14892 (N_14892,N_12412,N_13376);
and U14893 (N_14893,N_13703,N_13663);
nor U14894 (N_14894,N_13702,N_13968);
nand U14895 (N_14895,N_12884,N_12264);
and U14896 (N_14896,N_13535,N_13108);
or U14897 (N_14897,N_12894,N_13906);
xor U14898 (N_14898,N_12144,N_13159);
xor U14899 (N_14899,N_13858,N_13317);
or U14900 (N_14900,N_13483,N_12992);
nor U14901 (N_14901,N_13116,N_13523);
nand U14902 (N_14902,N_12682,N_12694);
nand U14903 (N_14903,N_12475,N_12127);
nor U14904 (N_14904,N_12165,N_12198);
nor U14905 (N_14905,N_12185,N_13205);
nand U14906 (N_14906,N_12193,N_12838);
xnor U14907 (N_14907,N_12212,N_12137);
and U14908 (N_14908,N_12123,N_13149);
or U14909 (N_14909,N_12374,N_13767);
nor U14910 (N_14910,N_13960,N_12864);
and U14911 (N_14911,N_12974,N_13430);
or U14912 (N_14912,N_13934,N_12997);
nor U14913 (N_14913,N_13301,N_12112);
xnor U14914 (N_14914,N_13377,N_13092);
xnor U14915 (N_14915,N_13146,N_12860);
nor U14916 (N_14916,N_13057,N_13655);
nand U14917 (N_14917,N_12536,N_13810);
and U14918 (N_14918,N_12274,N_13825);
nor U14919 (N_14919,N_13357,N_13637);
or U14920 (N_14920,N_12805,N_13640);
xor U14921 (N_14921,N_13246,N_12022);
or U14922 (N_14922,N_13790,N_13449);
xnor U14923 (N_14923,N_13505,N_12557);
xor U14924 (N_14924,N_13263,N_13242);
xor U14925 (N_14925,N_12415,N_12434);
nor U14926 (N_14926,N_12764,N_13562);
nand U14927 (N_14927,N_12246,N_12963);
or U14928 (N_14928,N_12157,N_13581);
xnor U14929 (N_14929,N_12354,N_12348);
xor U14930 (N_14930,N_12257,N_13995);
nand U14931 (N_14931,N_12528,N_13180);
nand U14932 (N_14932,N_13189,N_13119);
and U14933 (N_14933,N_13293,N_13757);
nor U14934 (N_14934,N_12556,N_13342);
or U14935 (N_14935,N_12174,N_13534);
nor U14936 (N_14936,N_13504,N_13199);
nand U14937 (N_14937,N_13437,N_12342);
nand U14938 (N_14938,N_13831,N_13802);
nor U14939 (N_14939,N_13148,N_12928);
or U14940 (N_14940,N_13104,N_12086);
and U14941 (N_14941,N_13773,N_12389);
nand U14942 (N_14942,N_13532,N_12636);
or U14943 (N_14943,N_13541,N_12399);
or U14944 (N_14944,N_12100,N_12362);
nor U14945 (N_14945,N_13213,N_13444);
xnor U14946 (N_14946,N_12492,N_13735);
nor U14947 (N_14947,N_13848,N_12358);
or U14948 (N_14948,N_13682,N_12336);
nor U14949 (N_14949,N_12324,N_13093);
xor U14950 (N_14950,N_12609,N_12506);
xnor U14951 (N_14951,N_13744,N_12457);
nand U14952 (N_14952,N_12882,N_12019);
nor U14953 (N_14953,N_13266,N_12437);
nand U14954 (N_14954,N_12221,N_12547);
nand U14955 (N_14955,N_13369,N_12849);
and U14956 (N_14956,N_12052,N_13446);
and U14957 (N_14957,N_12801,N_13366);
xnor U14958 (N_14958,N_12683,N_12863);
or U14959 (N_14959,N_12618,N_13028);
xor U14960 (N_14960,N_12994,N_13738);
nor U14961 (N_14961,N_12231,N_13219);
nor U14962 (N_14962,N_13288,N_12391);
and U14963 (N_14963,N_12171,N_13886);
and U14964 (N_14964,N_12017,N_13497);
xnor U14965 (N_14965,N_12815,N_12777);
xor U14966 (N_14966,N_13975,N_13418);
and U14967 (N_14967,N_12311,N_13900);
or U14968 (N_14968,N_13740,N_13338);
nand U14969 (N_14969,N_13101,N_13432);
xnor U14970 (N_14970,N_12003,N_13538);
and U14971 (N_14971,N_13631,N_12784);
or U14972 (N_14972,N_12363,N_13950);
nand U14973 (N_14973,N_12268,N_13807);
and U14974 (N_14974,N_12345,N_12010);
xnor U14975 (N_14975,N_12499,N_13546);
xor U14976 (N_14976,N_12926,N_13068);
nor U14977 (N_14977,N_12647,N_13045);
nor U14978 (N_14978,N_13388,N_13394);
xor U14979 (N_14979,N_12794,N_12323);
nand U14980 (N_14980,N_13526,N_12675);
or U14981 (N_14981,N_12276,N_12656);
nand U14982 (N_14982,N_13124,N_12775);
or U14983 (N_14983,N_13996,N_13778);
and U14984 (N_14984,N_13371,N_13441);
nor U14985 (N_14985,N_12460,N_13136);
xor U14986 (N_14986,N_12154,N_12836);
or U14987 (N_14987,N_13264,N_13765);
nor U14988 (N_14988,N_12170,N_13014);
nand U14989 (N_14989,N_13519,N_13770);
nor U14990 (N_14990,N_13208,N_12567);
nor U14991 (N_14991,N_13402,N_12385);
nor U14992 (N_14992,N_13576,N_13460);
xnor U14993 (N_14993,N_12705,N_12200);
xnor U14994 (N_14994,N_12190,N_13396);
and U14995 (N_14995,N_12829,N_13762);
xnor U14996 (N_14996,N_13707,N_12422);
or U14997 (N_14997,N_13899,N_13247);
xor U14998 (N_14998,N_13973,N_12822);
nand U14999 (N_14999,N_12937,N_12923);
or U15000 (N_15000,N_12595,N_13441);
nor U15001 (N_15001,N_13472,N_12287);
and U15002 (N_15002,N_13722,N_13474);
and U15003 (N_15003,N_12346,N_12204);
nand U15004 (N_15004,N_12747,N_12375);
and U15005 (N_15005,N_13058,N_12491);
and U15006 (N_15006,N_13021,N_13655);
nand U15007 (N_15007,N_12343,N_12318);
nand U15008 (N_15008,N_13836,N_12964);
xnor U15009 (N_15009,N_12309,N_13886);
nand U15010 (N_15010,N_12316,N_12403);
and U15011 (N_15011,N_13102,N_13319);
nand U15012 (N_15012,N_12992,N_12846);
nor U15013 (N_15013,N_13040,N_13621);
nor U15014 (N_15014,N_13023,N_13382);
xnor U15015 (N_15015,N_13059,N_13655);
or U15016 (N_15016,N_13802,N_12911);
and U15017 (N_15017,N_13321,N_13560);
or U15018 (N_15018,N_13133,N_13049);
and U15019 (N_15019,N_13564,N_12771);
and U15020 (N_15020,N_13423,N_13274);
or U15021 (N_15021,N_13040,N_13205);
and U15022 (N_15022,N_12752,N_13148);
or U15023 (N_15023,N_13935,N_13478);
and U15024 (N_15024,N_12455,N_12498);
nor U15025 (N_15025,N_12196,N_12088);
nor U15026 (N_15026,N_13922,N_13962);
nor U15027 (N_15027,N_12727,N_12186);
or U15028 (N_15028,N_12251,N_13056);
xor U15029 (N_15029,N_13567,N_12381);
xor U15030 (N_15030,N_12229,N_13655);
xor U15031 (N_15031,N_13537,N_12955);
nand U15032 (N_15032,N_13704,N_13584);
or U15033 (N_15033,N_12483,N_13762);
nor U15034 (N_15034,N_12807,N_12440);
or U15035 (N_15035,N_13444,N_13657);
or U15036 (N_15036,N_12681,N_12019);
and U15037 (N_15037,N_13348,N_12816);
xnor U15038 (N_15038,N_12842,N_12088);
nor U15039 (N_15039,N_12579,N_13423);
nand U15040 (N_15040,N_12901,N_13692);
nand U15041 (N_15041,N_13995,N_13281);
or U15042 (N_15042,N_12954,N_13261);
nor U15043 (N_15043,N_13242,N_12786);
xor U15044 (N_15044,N_13590,N_12747);
nor U15045 (N_15045,N_13263,N_13566);
and U15046 (N_15046,N_13686,N_12562);
or U15047 (N_15047,N_12815,N_13929);
and U15048 (N_15048,N_13435,N_12704);
and U15049 (N_15049,N_13981,N_12923);
and U15050 (N_15050,N_13587,N_12609);
nor U15051 (N_15051,N_12707,N_13517);
nor U15052 (N_15052,N_13802,N_12269);
and U15053 (N_15053,N_13507,N_12528);
nor U15054 (N_15054,N_13110,N_12675);
and U15055 (N_15055,N_12353,N_12841);
xnor U15056 (N_15056,N_13360,N_12496);
and U15057 (N_15057,N_13890,N_12214);
nand U15058 (N_15058,N_12022,N_13241);
or U15059 (N_15059,N_13969,N_12969);
or U15060 (N_15060,N_13758,N_13167);
nand U15061 (N_15061,N_13989,N_12244);
xor U15062 (N_15062,N_12938,N_13213);
and U15063 (N_15063,N_12318,N_13840);
or U15064 (N_15064,N_12599,N_12437);
or U15065 (N_15065,N_13998,N_13718);
or U15066 (N_15066,N_12907,N_12124);
and U15067 (N_15067,N_12288,N_13562);
nor U15068 (N_15068,N_12088,N_12687);
nor U15069 (N_15069,N_12553,N_12779);
xnor U15070 (N_15070,N_12397,N_12592);
xnor U15071 (N_15071,N_12153,N_12218);
nand U15072 (N_15072,N_13377,N_12401);
nand U15073 (N_15073,N_12621,N_13792);
or U15074 (N_15074,N_13536,N_13129);
nor U15075 (N_15075,N_12626,N_12958);
nand U15076 (N_15076,N_13476,N_12647);
xnor U15077 (N_15077,N_13846,N_12915);
nand U15078 (N_15078,N_12329,N_13675);
xor U15079 (N_15079,N_13601,N_13670);
or U15080 (N_15080,N_12803,N_12842);
xnor U15081 (N_15081,N_13027,N_12825);
xnor U15082 (N_15082,N_12906,N_12469);
nand U15083 (N_15083,N_12215,N_13361);
nand U15084 (N_15084,N_12027,N_12401);
xnor U15085 (N_15085,N_12410,N_12196);
and U15086 (N_15086,N_13922,N_12883);
or U15087 (N_15087,N_12006,N_13100);
nor U15088 (N_15088,N_12122,N_12144);
xnor U15089 (N_15089,N_12700,N_12765);
nor U15090 (N_15090,N_12988,N_12120);
nor U15091 (N_15091,N_12466,N_12484);
nor U15092 (N_15092,N_13126,N_12340);
xor U15093 (N_15093,N_12852,N_12828);
xor U15094 (N_15094,N_12087,N_12421);
xor U15095 (N_15095,N_13742,N_13259);
and U15096 (N_15096,N_12217,N_13379);
nor U15097 (N_15097,N_12426,N_13737);
nor U15098 (N_15098,N_12237,N_13278);
or U15099 (N_15099,N_13840,N_12493);
or U15100 (N_15100,N_13634,N_13887);
xnor U15101 (N_15101,N_12777,N_13074);
nor U15102 (N_15102,N_13259,N_13664);
or U15103 (N_15103,N_12528,N_12868);
nor U15104 (N_15104,N_12480,N_13771);
or U15105 (N_15105,N_13957,N_12565);
or U15106 (N_15106,N_12259,N_13703);
or U15107 (N_15107,N_12960,N_12062);
xor U15108 (N_15108,N_13809,N_12419);
and U15109 (N_15109,N_13124,N_13105);
xor U15110 (N_15110,N_13568,N_13454);
nand U15111 (N_15111,N_13277,N_13127);
nand U15112 (N_15112,N_12251,N_12901);
nor U15113 (N_15113,N_12710,N_13821);
nor U15114 (N_15114,N_13885,N_12946);
and U15115 (N_15115,N_12432,N_13025);
nand U15116 (N_15116,N_13464,N_13943);
or U15117 (N_15117,N_12688,N_12798);
nor U15118 (N_15118,N_12855,N_13394);
and U15119 (N_15119,N_12824,N_12594);
nor U15120 (N_15120,N_13168,N_12807);
nor U15121 (N_15121,N_13585,N_12661);
nor U15122 (N_15122,N_12634,N_12321);
xor U15123 (N_15123,N_12898,N_12005);
xnor U15124 (N_15124,N_13887,N_13378);
nand U15125 (N_15125,N_12949,N_12875);
and U15126 (N_15126,N_12417,N_13288);
or U15127 (N_15127,N_13709,N_12843);
xnor U15128 (N_15128,N_12295,N_12227);
nand U15129 (N_15129,N_12326,N_13065);
or U15130 (N_15130,N_12842,N_12110);
nor U15131 (N_15131,N_13390,N_13074);
nand U15132 (N_15132,N_12502,N_12998);
nand U15133 (N_15133,N_13578,N_12083);
and U15134 (N_15134,N_12183,N_12172);
or U15135 (N_15135,N_13990,N_12690);
nand U15136 (N_15136,N_12772,N_12594);
or U15137 (N_15137,N_12677,N_12270);
or U15138 (N_15138,N_13901,N_13543);
nand U15139 (N_15139,N_13361,N_12332);
nand U15140 (N_15140,N_13790,N_13880);
nor U15141 (N_15141,N_13934,N_13845);
xnor U15142 (N_15142,N_12839,N_13074);
nor U15143 (N_15143,N_13266,N_13783);
nand U15144 (N_15144,N_13453,N_12957);
nand U15145 (N_15145,N_13877,N_12630);
xor U15146 (N_15146,N_13532,N_12053);
nand U15147 (N_15147,N_13814,N_12240);
nor U15148 (N_15148,N_12813,N_13098);
nand U15149 (N_15149,N_12515,N_12747);
and U15150 (N_15150,N_12673,N_13923);
or U15151 (N_15151,N_12834,N_13018);
or U15152 (N_15152,N_12433,N_13391);
nand U15153 (N_15153,N_12894,N_13497);
and U15154 (N_15154,N_13255,N_13699);
nor U15155 (N_15155,N_13841,N_12481);
and U15156 (N_15156,N_13948,N_12795);
or U15157 (N_15157,N_13828,N_13072);
nor U15158 (N_15158,N_13381,N_13974);
and U15159 (N_15159,N_13908,N_12815);
nor U15160 (N_15160,N_12254,N_13611);
nand U15161 (N_15161,N_13381,N_12627);
nand U15162 (N_15162,N_13530,N_13412);
xor U15163 (N_15163,N_13384,N_12663);
or U15164 (N_15164,N_13612,N_13358);
nand U15165 (N_15165,N_12790,N_13715);
xnor U15166 (N_15166,N_12502,N_12958);
and U15167 (N_15167,N_12564,N_12094);
and U15168 (N_15168,N_13053,N_12015);
xor U15169 (N_15169,N_13282,N_13644);
and U15170 (N_15170,N_12440,N_13803);
nor U15171 (N_15171,N_12935,N_12400);
nor U15172 (N_15172,N_13930,N_13300);
nand U15173 (N_15173,N_12034,N_13615);
xor U15174 (N_15174,N_12702,N_13277);
and U15175 (N_15175,N_12127,N_12193);
and U15176 (N_15176,N_13360,N_12809);
or U15177 (N_15177,N_12092,N_12949);
xnor U15178 (N_15178,N_12196,N_12447);
nand U15179 (N_15179,N_13950,N_12957);
xor U15180 (N_15180,N_12227,N_13950);
nand U15181 (N_15181,N_13449,N_13358);
and U15182 (N_15182,N_13406,N_13467);
and U15183 (N_15183,N_13741,N_12227);
nand U15184 (N_15184,N_13036,N_12454);
xor U15185 (N_15185,N_12836,N_12910);
nand U15186 (N_15186,N_13943,N_13555);
nor U15187 (N_15187,N_13602,N_12941);
nand U15188 (N_15188,N_12547,N_12828);
and U15189 (N_15189,N_13504,N_12421);
nand U15190 (N_15190,N_12063,N_13029);
nand U15191 (N_15191,N_13284,N_12362);
and U15192 (N_15192,N_12125,N_12075);
nand U15193 (N_15193,N_13489,N_13740);
xnor U15194 (N_15194,N_12867,N_13945);
xnor U15195 (N_15195,N_12781,N_12690);
and U15196 (N_15196,N_13290,N_13110);
xnor U15197 (N_15197,N_13122,N_13785);
and U15198 (N_15198,N_13131,N_13337);
or U15199 (N_15199,N_13558,N_12426);
nand U15200 (N_15200,N_13078,N_13538);
nor U15201 (N_15201,N_12800,N_13605);
nor U15202 (N_15202,N_13696,N_13098);
and U15203 (N_15203,N_13860,N_13012);
nor U15204 (N_15204,N_13475,N_12127);
nand U15205 (N_15205,N_12508,N_13579);
nand U15206 (N_15206,N_12680,N_12062);
and U15207 (N_15207,N_13665,N_13317);
xnor U15208 (N_15208,N_12476,N_12846);
nand U15209 (N_15209,N_13143,N_12318);
nand U15210 (N_15210,N_12149,N_12595);
or U15211 (N_15211,N_12128,N_12260);
and U15212 (N_15212,N_13401,N_13515);
or U15213 (N_15213,N_13831,N_12800);
and U15214 (N_15214,N_12652,N_13683);
nand U15215 (N_15215,N_12024,N_12585);
nand U15216 (N_15216,N_13548,N_12212);
xnor U15217 (N_15217,N_13280,N_13933);
or U15218 (N_15218,N_13011,N_13861);
nor U15219 (N_15219,N_13907,N_12102);
nor U15220 (N_15220,N_13700,N_13243);
xnor U15221 (N_15221,N_13717,N_12637);
or U15222 (N_15222,N_12022,N_12137);
nand U15223 (N_15223,N_12733,N_12288);
and U15224 (N_15224,N_13711,N_12577);
or U15225 (N_15225,N_13701,N_12106);
xnor U15226 (N_15226,N_12149,N_12862);
and U15227 (N_15227,N_12170,N_13077);
and U15228 (N_15228,N_12648,N_13131);
xor U15229 (N_15229,N_12262,N_12673);
and U15230 (N_15230,N_12688,N_12358);
nor U15231 (N_15231,N_12854,N_13224);
or U15232 (N_15232,N_12147,N_13035);
nor U15233 (N_15233,N_13153,N_13853);
nand U15234 (N_15234,N_13071,N_13802);
or U15235 (N_15235,N_13431,N_13567);
and U15236 (N_15236,N_13469,N_12898);
nand U15237 (N_15237,N_12167,N_13878);
xnor U15238 (N_15238,N_13176,N_13137);
nand U15239 (N_15239,N_12769,N_12787);
nor U15240 (N_15240,N_12691,N_12043);
or U15241 (N_15241,N_12869,N_12098);
nand U15242 (N_15242,N_13084,N_12948);
xor U15243 (N_15243,N_13275,N_13898);
nand U15244 (N_15244,N_12646,N_12521);
nand U15245 (N_15245,N_13124,N_12800);
or U15246 (N_15246,N_12949,N_12918);
xnor U15247 (N_15247,N_12031,N_13675);
and U15248 (N_15248,N_12802,N_12769);
and U15249 (N_15249,N_13740,N_12261);
or U15250 (N_15250,N_12625,N_13980);
nand U15251 (N_15251,N_12968,N_13416);
and U15252 (N_15252,N_13327,N_13141);
xor U15253 (N_15253,N_12618,N_12515);
nor U15254 (N_15254,N_12613,N_12704);
and U15255 (N_15255,N_13364,N_13410);
and U15256 (N_15256,N_12536,N_13743);
and U15257 (N_15257,N_12150,N_12997);
nor U15258 (N_15258,N_12887,N_13808);
xnor U15259 (N_15259,N_13943,N_13319);
nand U15260 (N_15260,N_12711,N_12984);
xor U15261 (N_15261,N_13034,N_12861);
nand U15262 (N_15262,N_12517,N_12979);
nor U15263 (N_15263,N_12993,N_12976);
nand U15264 (N_15264,N_13639,N_12288);
xnor U15265 (N_15265,N_13922,N_12793);
nand U15266 (N_15266,N_13675,N_13407);
or U15267 (N_15267,N_12669,N_12026);
and U15268 (N_15268,N_13078,N_12074);
nand U15269 (N_15269,N_12438,N_12673);
xor U15270 (N_15270,N_12973,N_13437);
xor U15271 (N_15271,N_13053,N_13278);
nand U15272 (N_15272,N_13878,N_13360);
and U15273 (N_15273,N_12822,N_13168);
nand U15274 (N_15274,N_13536,N_12863);
nand U15275 (N_15275,N_13049,N_13088);
nand U15276 (N_15276,N_12648,N_12203);
or U15277 (N_15277,N_12442,N_13601);
and U15278 (N_15278,N_12402,N_13686);
xnor U15279 (N_15279,N_12631,N_12864);
nor U15280 (N_15280,N_13968,N_13784);
nor U15281 (N_15281,N_13669,N_12764);
nand U15282 (N_15282,N_13909,N_13721);
xor U15283 (N_15283,N_13165,N_13218);
xor U15284 (N_15284,N_12413,N_13599);
and U15285 (N_15285,N_13134,N_13740);
nor U15286 (N_15286,N_12143,N_13060);
nor U15287 (N_15287,N_12462,N_12840);
nor U15288 (N_15288,N_13118,N_12098);
xnor U15289 (N_15289,N_12688,N_13189);
nand U15290 (N_15290,N_13042,N_13872);
and U15291 (N_15291,N_12071,N_13665);
nor U15292 (N_15292,N_13574,N_12162);
and U15293 (N_15293,N_13624,N_12563);
xnor U15294 (N_15294,N_13369,N_12936);
or U15295 (N_15295,N_12940,N_12072);
or U15296 (N_15296,N_12685,N_12364);
nor U15297 (N_15297,N_12029,N_12936);
or U15298 (N_15298,N_12524,N_13675);
nor U15299 (N_15299,N_12178,N_13527);
nand U15300 (N_15300,N_12158,N_13848);
nand U15301 (N_15301,N_13253,N_13680);
or U15302 (N_15302,N_13945,N_13183);
nor U15303 (N_15303,N_12054,N_13425);
nor U15304 (N_15304,N_12060,N_13029);
or U15305 (N_15305,N_13994,N_12031);
nand U15306 (N_15306,N_13817,N_12056);
or U15307 (N_15307,N_12859,N_13559);
nor U15308 (N_15308,N_13281,N_12747);
xnor U15309 (N_15309,N_13523,N_12357);
or U15310 (N_15310,N_13905,N_13043);
nor U15311 (N_15311,N_12350,N_12842);
nand U15312 (N_15312,N_13518,N_13158);
nand U15313 (N_15313,N_12928,N_13229);
nand U15314 (N_15314,N_13945,N_12673);
nand U15315 (N_15315,N_12121,N_12341);
and U15316 (N_15316,N_13979,N_13075);
or U15317 (N_15317,N_13489,N_13179);
and U15318 (N_15318,N_12816,N_13315);
or U15319 (N_15319,N_13383,N_13216);
nand U15320 (N_15320,N_13779,N_12061);
or U15321 (N_15321,N_12179,N_12739);
nand U15322 (N_15322,N_12708,N_13024);
nand U15323 (N_15323,N_12023,N_13462);
xnor U15324 (N_15324,N_12101,N_13698);
and U15325 (N_15325,N_12684,N_12125);
nand U15326 (N_15326,N_12338,N_13268);
or U15327 (N_15327,N_12440,N_12097);
xnor U15328 (N_15328,N_13923,N_13418);
xnor U15329 (N_15329,N_13620,N_13890);
or U15330 (N_15330,N_12396,N_12065);
nand U15331 (N_15331,N_12680,N_12957);
or U15332 (N_15332,N_12783,N_12869);
xnor U15333 (N_15333,N_12672,N_13306);
and U15334 (N_15334,N_12261,N_12031);
nand U15335 (N_15335,N_13838,N_12078);
and U15336 (N_15336,N_12132,N_13855);
xor U15337 (N_15337,N_12924,N_13115);
and U15338 (N_15338,N_12184,N_13392);
or U15339 (N_15339,N_13883,N_12436);
nor U15340 (N_15340,N_12093,N_12197);
or U15341 (N_15341,N_13878,N_12598);
xnor U15342 (N_15342,N_12258,N_13318);
nand U15343 (N_15343,N_13539,N_13996);
and U15344 (N_15344,N_12018,N_12861);
xor U15345 (N_15345,N_13021,N_12230);
nor U15346 (N_15346,N_12800,N_12554);
xor U15347 (N_15347,N_12584,N_13638);
xor U15348 (N_15348,N_12436,N_13653);
and U15349 (N_15349,N_13996,N_13999);
and U15350 (N_15350,N_13516,N_12642);
or U15351 (N_15351,N_13472,N_12699);
and U15352 (N_15352,N_13869,N_13094);
nand U15353 (N_15353,N_13024,N_12886);
and U15354 (N_15354,N_12567,N_12419);
nor U15355 (N_15355,N_13238,N_13224);
or U15356 (N_15356,N_13038,N_13795);
or U15357 (N_15357,N_13603,N_13081);
nor U15358 (N_15358,N_12591,N_13982);
or U15359 (N_15359,N_12245,N_12969);
or U15360 (N_15360,N_12179,N_12343);
or U15361 (N_15361,N_12458,N_12431);
nor U15362 (N_15362,N_12463,N_12694);
and U15363 (N_15363,N_13796,N_12687);
nand U15364 (N_15364,N_12093,N_13804);
nand U15365 (N_15365,N_12241,N_12941);
xor U15366 (N_15366,N_13982,N_13342);
xor U15367 (N_15367,N_12052,N_12164);
nor U15368 (N_15368,N_12482,N_13235);
and U15369 (N_15369,N_13782,N_12598);
nor U15370 (N_15370,N_12979,N_13590);
or U15371 (N_15371,N_12468,N_12073);
xor U15372 (N_15372,N_12128,N_12343);
xor U15373 (N_15373,N_12759,N_13785);
nor U15374 (N_15374,N_13402,N_13613);
or U15375 (N_15375,N_12849,N_12533);
or U15376 (N_15376,N_13885,N_12532);
nor U15377 (N_15377,N_12060,N_13851);
xor U15378 (N_15378,N_12654,N_13646);
xor U15379 (N_15379,N_13085,N_13609);
and U15380 (N_15380,N_13717,N_13642);
and U15381 (N_15381,N_12503,N_12518);
nand U15382 (N_15382,N_12032,N_12936);
or U15383 (N_15383,N_12587,N_12913);
and U15384 (N_15384,N_13317,N_13642);
nand U15385 (N_15385,N_13647,N_12285);
nand U15386 (N_15386,N_12521,N_13924);
and U15387 (N_15387,N_13925,N_13525);
and U15388 (N_15388,N_12414,N_13299);
nand U15389 (N_15389,N_12105,N_13386);
nor U15390 (N_15390,N_12872,N_13134);
xor U15391 (N_15391,N_12917,N_12406);
and U15392 (N_15392,N_12101,N_12167);
nor U15393 (N_15393,N_12297,N_13333);
xnor U15394 (N_15394,N_13867,N_12272);
nor U15395 (N_15395,N_12603,N_13234);
nand U15396 (N_15396,N_13264,N_13192);
xor U15397 (N_15397,N_12194,N_13192);
and U15398 (N_15398,N_13709,N_12930);
nand U15399 (N_15399,N_12447,N_12783);
nand U15400 (N_15400,N_13732,N_13854);
nand U15401 (N_15401,N_12192,N_12403);
nand U15402 (N_15402,N_13743,N_12680);
and U15403 (N_15403,N_13431,N_12396);
and U15404 (N_15404,N_12549,N_13516);
or U15405 (N_15405,N_13219,N_13503);
xor U15406 (N_15406,N_12432,N_12678);
xor U15407 (N_15407,N_13690,N_12270);
nor U15408 (N_15408,N_13704,N_13303);
and U15409 (N_15409,N_13687,N_12036);
xnor U15410 (N_15410,N_12050,N_13610);
nand U15411 (N_15411,N_13045,N_12980);
nor U15412 (N_15412,N_13992,N_12137);
and U15413 (N_15413,N_12493,N_13463);
nor U15414 (N_15414,N_13406,N_12604);
nor U15415 (N_15415,N_13794,N_12587);
nor U15416 (N_15416,N_13554,N_12395);
nor U15417 (N_15417,N_13630,N_13785);
nor U15418 (N_15418,N_12826,N_12535);
or U15419 (N_15419,N_12991,N_12641);
xor U15420 (N_15420,N_13350,N_12666);
or U15421 (N_15421,N_13619,N_13839);
or U15422 (N_15422,N_13712,N_13073);
and U15423 (N_15423,N_13596,N_12394);
nand U15424 (N_15424,N_12705,N_13625);
and U15425 (N_15425,N_12461,N_13431);
nand U15426 (N_15426,N_13545,N_13065);
xnor U15427 (N_15427,N_13442,N_13491);
and U15428 (N_15428,N_12125,N_12379);
and U15429 (N_15429,N_12988,N_12881);
nor U15430 (N_15430,N_12730,N_12788);
xor U15431 (N_15431,N_12116,N_13538);
and U15432 (N_15432,N_12456,N_12538);
or U15433 (N_15433,N_13192,N_13642);
or U15434 (N_15434,N_12318,N_13919);
and U15435 (N_15435,N_13745,N_13862);
nand U15436 (N_15436,N_13249,N_12982);
nor U15437 (N_15437,N_12957,N_12972);
nor U15438 (N_15438,N_12960,N_12842);
and U15439 (N_15439,N_12549,N_13113);
nor U15440 (N_15440,N_13989,N_13406);
nand U15441 (N_15441,N_13784,N_12370);
or U15442 (N_15442,N_13178,N_13265);
nand U15443 (N_15443,N_12297,N_13479);
nor U15444 (N_15444,N_13380,N_13814);
xnor U15445 (N_15445,N_12823,N_13398);
and U15446 (N_15446,N_13227,N_13202);
or U15447 (N_15447,N_12919,N_13616);
or U15448 (N_15448,N_12592,N_12506);
nand U15449 (N_15449,N_13049,N_13163);
nand U15450 (N_15450,N_12336,N_13263);
nor U15451 (N_15451,N_13812,N_13462);
and U15452 (N_15452,N_13115,N_12817);
and U15453 (N_15453,N_12265,N_12704);
nor U15454 (N_15454,N_12910,N_13567);
or U15455 (N_15455,N_13196,N_13205);
or U15456 (N_15456,N_13657,N_12623);
nand U15457 (N_15457,N_13536,N_12306);
or U15458 (N_15458,N_12860,N_12890);
or U15459 (N_15459,N_13017,N_12499);
nand U15460 (N_15460,N_13322,N_13106);
nor U15461 (N_15461,N_12710,N_12298);
or U15462 (N_15462,N_12444,N_12206);
xor U15463 (N_15463,N_12328,N_12356);
or U15464 (N_15464,N_12726,N_13207);
or U15465 (N_15465,N_12541,N_13142);
nand U15466 (N_15466,N_12253,N_13350);
nand U15467 (N_15467,N_12482,N_13260);
nand U15468 (N_15468,N_12882,N_13680);
and U15469 (N_15469,N_13937,N_12865);
and U15470 (N_15470,N_12765,N_13111);
or U15471 (N_15471,N_13287,N_12176);
xnor U15472 (N_15472,N_13006,N_13145);
nand U15473 (N_15473,N_12047,N_12114);
nor U15474 (N_15474,N_13615,N_12242);
nor U15475 (N_15475,N_12782,N_13407);
or U15476 (N_15476,N_12462,N_13357);
nor U15477 (N_15477,N_13758,N_13636);
nor U15478 (N_15478,N_13098,N_12521);
or U15479 (N_15479,N_13550,N_12936);
or U15480 (N_15480,N_13417,N_13913);
nand U15481 (N_15481,N_12381,N_13207);
nand U15482 (N_15482,N_13914,N_12902);
or U15483 (N_15483,N_13019,N_13527);
or U15484 (N_15484,N_12682,N_12118);
xor U15485 (N_15485,N_13321,N_13122);
or U15486 (N_15486,N_13828,N_12462);
xnor U15487 (N_15487,N_13989,N_13773);
or U15488 (N_15488,N_12983,N_13768);
and U15489 (N_15489,N_13604,N_12379);
nor U15490 (N_15490,N_12742,N_12732);
and U15491 (N_15491,N_13795,N_12403);
or U15492 (N_15492,N_12559,N_13682);
nor U15493 (N_15493,N_12575,N_13883);
nand U15494 (N_15494,N_13126,N_12201);
and U15495 (N_15495,N_12752,N_12462);
xor U15496 (N_15496,N_12443,N_12832);
and U15497 (N_15497,N_12510,N_12072);
and U15498 (N_15498,N_12416,N_12789);
and U15499 (N_15499,N_13561,N_13747);
xor U15500 (N_15500,N_12298,N_13889);
nand U15501 (N_15501,N_13601,N_13298);
and U15502 (N_15502,N_12593,N_12943);
xor U15503 (N_15503,N_13658,N_12871);
nor U15504 (N_15504,N_13401,N_13203);
or U15505 (N_15505,N_12312,N_12271);
nor U15506 (N_15506,N_12866,N_12333);
nand U15507 (N_15507,N_12588,N_13862);
xnor U15508 (N_15508,N_13631,N_12610);
nor U15509 (N_15509,N_12274,N_12430);
and U15510 (N_15510,N_13949,N_12211);
xor U15511 (N_15511,N_13783,N_13686);
xnor U15512 (N_15512,N_13407,N_13523);
nor U15513 (N_15513,N_12613,N_12952);
and U15514 (N_15514,N_13601,N_13198);
nand U15515 (N_15515,N_12977,N_12825);
or U15516 (N_15516,N_12225,N_13844);
xor U15517 (N_15517,N_12162,N_12185);
and U15518 (N_15518,N_13968,N_12047);
and U15519 (N_15519,N_12519,N_13181);
nor U15520 (N_15520,N_13583,N_12579);
nor U15521 (N_15521,N_13331,N_13934);
nor U15522 (N_15522,N_13032,N_12208);
xor U15523 (N_15523,N_13011,N_13666);
xnor U15524 (N_15524,N_13149,N_12897);
or U15525 (N_15525,N_12745,N_12966);
or U15526 (N_15526,N_13126,N_12628);
and U15527 (N_15527,N_13019,N_12741);
and U15528 (N_15528,N_12372,N_12530);
nor U15529 (N_15529,N_13324,N_12670);
nor U15530 (N_15530,N_12270,N_13859);
nor U15531 (N_15531,N_12907,N_12309);
or U15532 (N_15532,N_12233,N_12345);
and U15533 (N_15533,N_13278,N_12601);
or U15534 (N_15534,N_13450,N_13552);
nor U15535 (N_15535,N_12943,N_13269);
xor U15536 (N_15536,N_12207,N_12487);
nor U15537 (N_15537,N_13179,N_13610);
nor U15538 (N_15538,N_12328,N_13852);
nand U15539 (N_15539,N_12753,N_12091);
and U15540 (N_15540,N_13016,N_12630);
nand U15541 (N_15541,N_12978,N_12283);
or U15542 (N_15542,N_13127,N_12767);
nor U15543 (N_15543,N_13606,N_13829);
nand U15544 (N_15544,N_12613,N_13323);
xnor U15545 (N_15545,N_13208,N_13026);
nand U15546 (N_15546,N_13359,N_13373);
or U15547 (N_15547,N_13839,N_12376);
and U15548 (N_15548,N_12907,N_13347);
nor U15549 (N_15549,N_13754,N_12024);
or U15550 (N_15550,N_12596,N_13138);
nor U15551 (N_15551,N_13078,N_13308);
nor U15552 (N_15552,N_12644,N_13216);
xor U15553 (N_15553,N_12556,N_12016);
xnor U15554 (N_15554,N_12214,N_13843);
nand U15555 (N_15555,N_13522,N_12891);
xnor U15556 (N_15556,N_12400,N_13398);
nor U15557 (N_15557,N_13960,N_12607);
and U15558 (N_15558,N_12422,N_12593);
nor U15559 (N_15559,N_12403,N_12901);
xor U15560 (N_15560,N_12187,N_13451);
or U15561 (N_15561,N_12484,N_13819);
nor U15562 (N_15562,N_13064,N_12300);
or U15563 (N_15563,N_12032,N_12469);
nand U15564 (N_15564,N_13656,N_12194);
xor U15565 (N_15565,N_13249,N_13579);
xor U15566 (N_15566,N_12749,N_13861);
nand U15567 (N_15567,N_13103,N_13677);
nand U15568 (N_15568,N_13393,N_13389);
nand U15569 (N_15569,N_12377,N_13099);
or U15570 (N_15570,N_12335,N_12694);
nand U15571 (N_15571,N_13248,N_13595);
nor U15572 (N_15572,N_12413,N_13209);
nor U15573 (N_15573,N_13748,N_13798);
nor U15574 (N_15574,N_12985,N_13496);
nor U15575 (N_15575,N_13588,N_12173);
or U15576 (N_15576,N_13868,N_12613);
and U15577 (N_15577,N_13078,N_12792);
xnor U15578 (N_15578,N_12929,N_13295);
or U15579 (N_15579,N_12916,N_12325);
xor U15580 (N_15580,N_12053,N_12273);
xnor U15581 (N_15581,N_13895,N_12754);
or U15582 (N_15582,N_13231,N_12094);
or U15583 (N_15583,N_12953,N_13886);
nor U15584 (N_15584,N_12917,N_13922);
and U15585 (N_15585,N_12434,N_12245);
xor U15586 (N_15586,N_12287,N_12693);
nor U15587 (N_15587,N_12551,N_12229);
and U15588 (N_15588,N_12638,N_13623);
nand U15589 (N_15589,N_12832,N_13784);
or U15590 (N_15590,N_13909,N_13341);
nor U15591 (N_15591,N_12845,N_12117);
or U15592 (N_15592,N_12285,N_12975);
nor U15593 (N_15593,N_13333,N_13316);
xnor U15594 (N_15594,N_12743,N_13714);
nand U15595 (N_15595,N_12330,N_12931);
and U15596 (N_15596,N_13452,N_13100);
nor U15597 (N_15597,N_12394,N_13460);
and U15598 (N_15598,N_13112,N_13028);
nor U15599 (N_15599,N_13251,N_12174);
nor U15600 (N_15600,N_12700,N_12362);
and U15601 (N_15601,N_12869,N_13659);
nand U15602 (N_15602,N_13949,N_13161);
nor U15603 (N_15603,N_12985,N_12214);
xor U15604 (N_15604,N_13391,N_12871);
nor U15605 (N_15605,N_12819,N_12041);
or U15606 (N_15606,N_13548,N_13921);
nand U15607 (N_15607,N_12446,N_12742);
nor U15608 (N_15608,N_13699,N_12006);
nor U15609 (N_15609,N_13283,N_12885);
nand U15610 (N_15610,N_13452,N_12876);
and U15611 (N_15611,N_12852,N_12513);
nand U15612 (N_15612,N_13470,N_13729);
nor U15613 (N_15613,N_13066,N_13691);
and U15614 (N_15614,N_12113,N_13311);
xor U15615 (N_15615,N_13548,N_13193);
and U15616 (N_15616,N_13663,N_13376);
nand U15617 (N_15617,N_12675,N_13970);
and U15618 (N_15618,N_12477,N_13199);
and U15619 (N_15619,N_12051,N_12675);
xnor U15620 (N_15620,N_12729,N_12798);
nor U15621 (N_15621,N_12671,N_13587);
xnor U15622 (N_15622,N_13186,N_13296);
nand U15623 (N_15623,N_12293,N_12402);
and U15624 (N_15624,N_12822,N_12433);
xnor U15625 (N_15625,N_13953,N_13366);
xnor U15626 (N_15626,N_13327,N_13484);
xnor U15627 (N_15627,N_13426,N_12464);
or U15628 (N_15628,N_13046,N_13585);
nand U15629 (N_15629,N_12234,N_13524);
nor U15630 (N_15630,N_12411,N_12038);
and U15631 (N_15631,N_12866,N_12372);
xnor U15632 (N_15632,N_13823,N_12473);
nand U15633 (N_15633,N_13247,N_13149);
xor U15634 (N_15634,N_12975,N_13101);
nand U15635 (N_15635,N_12340,N_13826);
nand U15636 (N_15636,N_13102,N_13751);
xor U15637 (N_15637,N_12121,N_13265);
or U15638 (N_15638,N_13135,N_13399);
or U15639 (N_15639,N_12013,N_12332);
nor U15640 (N_15640,N_12613,N_13418);
nor U15641 (N_15641,N_13072,N_13399);
nor U15642 (N_15642,N_12080,N_13480);
nand U15643 (N_15643,N_13005,N_13539);
or U15644 (N_15644,N_13399,N_12902);
xnor U15645 (N_15645,N_12483,N_13075);
xor U15646 (N_15646,N_12521,N_12168);
nand U15647 (N_15647,N_13636,N_13865);
xnor U15648 (N_15648,N_13275,N_12644);
xnor U15649 (N_15649,N_13108,N_12676);
nor U15650 (N_15650,N_12182,N_12767);
and U15651 (N_15651,N_13794,N_13348);
and U15652 (N_15652,N_13215,N_13659);
nand U15653 (N_15653,N_12992,N_12112);
nand U15654 (N_15654,N_12173,N_13134);
xor U15655 (N_15655,N_12680,N_12987);
or U15656 (N_15656,N_12028,N_13707);
nand U15657 (N_15657,N_13036,N_13052);
and U15658 (N_15658,N_13135,N_13107);
and U15659 (N_15659,N_13712,N_13600);
nand U15660 (N_15660,N_13914,N_12201);
nand U15661 (N_15661,N_12382,N_12939);
nor U15662 (N_15662,N_12216,N_12613);
nor U15663 (N_15663,N_12215,N_12552);
or U15664 (N_15664,N_13383,N_13657);
nor U15665 (N_15665,N_12054,N_13435);
xnor U15666 (N_15666,N_12770,N_13738);
and U15667 (N_15667,N_13420,N_13576);
or U15668 (N_15668,N_12708,N_13549);
or U15669 (N_15669,N_13502,N_12201);
and U15670 (N_15670,N_13610,N_13746);
nand U15671 (N_15671,N_12459,N_12777);
nand U15672 (N_15672,N_13229,N_12930);
nor U15673 (N_15673,N_13156,N_12444);
nand U15674 (N_15674,N_13912,N_12097);
or U15675 (N_15675,N_12433,N_13972);
or U15676 (N_15676,N_13994,N_12392);
nand U15677 (N_15677,N_12533,N_13532);
or U15678 (N_15678,N_13066,N_12411);
or U15679 (N_15679,N_13107,N_12346);
or U15680 (N_15680,N_13254,N_13430);
or U15681 (N_15681,N_12126,N_12944);
xor U15682 (N_15682,N_12837,N_12804);
xnor U15683 (N_15683,N_13768,N_13540);
or U15684 (N_15684,N_13600,N_13764);
xnor U15685 (N_15685,N_13805,N_12105);
nor U15686 (N_15686,N_12875,N_12573);
xor U15687 (N_15687,N_12035,N_13726);
nand U15688 (N_15688,N_13309,N_12180);
or U15689 (N_15689,N_13825,N_13511);
nand U15690 (N_15690,N_12408,N_12550);
xnor U15691 (N_15691,N_13350,N_12374);
and U15692 (N_15692,N_13007,N_13125);
nand U15693 (N_15693,N_12254,N_12287);
or U15694 (N_15694,N_13133,N_13452);
nand U15695 (N_15695,N_12000,N_12830);
nand U15696 (N_15696,N_13443,N_13050);
nor U15697 (N_15697,N_13744,N_13575);
nor U15698 (N_15698,N_13978,N_13057);
nor U15699 (N_15699,N_12148,N_12757);
and U15700 (N_15700,N_12340,N_12392);
and U15701 (N_15701,N_13028,N_13832);
xor U15702 (N_15702,N_12352,N_13415);
nor U15703 (N_15703,N_13796,N_12117);
nor U15704 (N_15704,N_12892,N_13974);
nor U15705 (N_15705,N_12548,N_13751);
nor U15706 (N_15706,N_13206,N_12544);
nor U15707 (N_15707,N_12171,N_12202);
or U15708 (N_15708,N_12508,N_12593);
or U15709 (N_15709,N_13499,N_13903);
nand U15710 (N_15710,N_13655,N_13005);
xnor U15711 (N_15711,N_13943,N_12811);
nor U15712 (N_15712,N_12462,N_12711);
nand U15713 (N_15713,N_12339,N_12436);
nand U15714 (N_15714,N_12754,N_12307);
or U15715 (N_15715,N_12871,N_12182);
xnor U15716 (N_15716,N_12560,N_13616);
nand U15717 (N_15717,N_13510,N_12083);
nand U15718 (N_15718,N_13881,N_12619);
and U15719 (N_15719,N_12096,N_12341);
and U15720 (N_15720,N_12702,N_13582);
nand U15721 (N_15721,N_12372,N_12504);
or U15722 (N_15722,N_13499,N_12775);
xor U15723 (N_15723,N_13858,N_13035);
nor U15724 (N_15724,N_13388,N_13055);
nand U15725 (N_15725,N_12192,N_12286);
nor U15726 (N_15726,N_13547,N_12184);
nor U15727 (N_15727,N_13754,N_12020);
nor U15728 (N_15728,N_13971,N_13350);
nand U15729 (N_15729,N_12741,N_13818);
nand U15730 (N_15730,N_12089,N_12905);
xor U15731 (N_15731,N_13812,N_13323);
nor U15732 (N_15732,N_13281,N_12180);
or U15733 (N_15733,N_12914,N_12527);
xnor U15734 (N_15734,N_13260,N_13497);
nand U15735 (N_15735,N_12920,N_12189);
nor U15736 (N_15736,N_13079,N_13907);
and U15737 (N_15737,N_13165,N_12139);
xor U15738 (N_15738,N_12618,N_12824);
xnor U15739 (N_15739,N_13579,N_12923);
nand U15740 (N_15740,N_12412,N_13037);
nor U15741 (N_15741,N_13154,N_13707);
xor U15742 (N_15742,N_13673,N_12307);
xor U15743 (N_15743,N_13666,N_12228);
or U15744 (N_15744,N_12204,N_12434);
nor U15745 (N_15745,N_13205,N_12479);
xnor U15746 (N_15746,N_12470,N_13027);
nand U15747 (N_15747,N_13423,N_13421);
xor U15748 (N_15748,N_13783,N_13256);
or U15749 (N_15749,N_13348,N_13264);
xnor U15750 (N_15750,N_12621,N_12036);
nand U15751 (N_15751,N_12689,N_13805);
or U15752 (N_15752,N_12993,N_13061);
and U15753 (N_15753,N_13418,N_13872);
nand U15754 (N_15754,N_13021,N_12769);
xnor U15755 (N_15755,N_13487,N_13871);
xor U15756 (N_15756,N_12413,N_12281);
nand U15757 (N_15757,N_13393,N_12170);
and U15758 (N_15758,N_13262,N_12659);
xnor U15759 (N_15759,N_13126,N_13292);
nor U15760 (N_15760,N_13563,N_12537);
or U15761 (N_15761,N_12639,N_12116);
xor U15762 (N_15762,N_12694,N_13991);
or U15763 (N_15763,N_13617,N_12538);
nor U15764 (N_15764,N_13302,N_12059);
nand U15765 (N_15765,N_12532,N_13671);
or U15766 (N_15766,N_13495,N_12734);
and U15767 (N_15767,N_12437,N_12228);
or U15768 (N_15768,N_13624,N_12343);
and U15769 (N_15769,N_13221,N_13393);
or U15770 (N_15770,N_13128,N_13136);
and U15771 (N_15771,N_12582,N_12957);
or U15772 (N_15772,N_12194,N_12309);
nor U15773 (N_15773,N_13511,N_13089);
or U15774 (N_15774,N_13632,N_12339);
nand U15775 (N_15775,N_13442,N_13118);
and U15776 (N_15776,N_13013,N_12700);
nor U15777 (N_15777,N_12114,N_13706);
or U15778 (N_15778,N_13482,N_13407);
and U15779 (N_15779,N_12833,N_13187);
or U15780 (N_15780,N_12249,N_13862);
nor U15781 (N_15781,N_12469,N_12157);
xnor U15782 (N_15782,N_13562,N_13581);
and U15783 (N_15783,N_12340,N_13493);
nand U15784 (N_15784,N_13595,N_13095);
xnor U15785 (N_15785,N_13940,N_12476);
xor U15786 (N_15786,N_12840,N_12573);
nand U15787 (N_15787,N_13390,N_13076);
or U15788 (N_15788,N_12994,N_12698);
nand U15789 (N_15789,N_13778,N_12989);
xnor U15790 (N_15790,N_12279,N_12201);
xor U15791 (N_15791,N_13627,N_12141);
nand U15792 (N_15792,N_13434,N_13408);
and U15793 (N_15793,N_13299,N_13911);
nor U15794 (N_15794,N_12112,N_12451);
and U15795 (N_15795,N_13126,N_13775);
nand U15796 (N_15796,N_12153,N_12361);
nor U15797 (N_15797,N_12354,N_12537);
and U15798 (N_15798,N_12053,N_13661);
xnor U15799 (N_15799,N_12293,N_12837);
nor U15800 (N_15800,N_12991,N_12939);
or U15801 (N_15801,N_12660,N_13349);
nor U15802 (N_15802,N_13578,N_13600);
nand U15803 (N_15803,N_13813,N_12489);
and U15804 (N_15804,N_12940,N_13270);
nand U15805 (N_15805,N_13586,N_13101);
or U15806 (N_15806,N_13886,N_12221);
or U15807 (N_15807,N_12163,N_13543);
and U15808 (N_15808,N_12434,N_12298);
nand U15809 (N_15809,N_13322,N_12731);
nand U15810 (N_15810,N_13047,N_13116);
nor U15811 (N_15811,N_13676,N_13792);
nand U15812 (N_15812,N_12505,N_13290);
nor U15813 (N_15813,N_12777,N_12566);
or U15814 (N_15814,N_12023,N_12657);
nand U15815 (N_15815,N_12079,N_13966);
nor U15816 (N_15816,N_12088,N_13691);
or U15817 (N_15817,N_13473,N_13200);
nor U15818 (N_15818,N_13121,N_12848);
nor U15819 (N_15819,N_13507,N_13516);
or U15820 (N_15820,N_12012,N_12694);
or U15821 (N_15821,N_12582,N_12257);
nor U15822 (N_15822,N_12058,N_13309);
nor U15823 (N_15823,N_13247,N_13981);
and U15824 (N_15824,N_12505,N_12543);
xnor U15825 (N_15825,N_13409,N_12613);
and U15826 (N_15826,N_12280,N_13321);
or U15827 (N_15827,N_12214,N_13443);
and U15828 (N_15828,N_13367,N_12750);
and U15829 (N_15829,N_12472,N_12559);
nand U15830 (N_15830,N_13000,N_13133);
nor U15831 (N_15831,N_12648,N_13912);
nand U15832 (N_15832,N_12422,N_12920);
nor U15833 (N_15833,N_12282,N_13297);
and U15834 (N_15834,N_13579,N_12698);
nand U15835 (N_15835,N_12928,N_13217);
and U15836 (N_15836,N_12195,N_13607);
xor U15837 (N_15837,N_13164,N_13300);
nand U15838 (N_15838,N_12032,N_13300);
and U15839 (N_15839,N_13738,N_13547);
nor U15840 (N_15840,N_12047,N_12589);
or U15841 (N_15841,N_12548,N_13154);
xnor U15842 (N_15842,N_13979,N_12885);
or U15843 (N_15843,N_13808,N_12293);
nor U15844 (N_15844,N_13564,N_12804);
xor U15845 (N_15845,N_13769,N_13050);
and U15846 (N_15846,N_12339,N_12864);
xor U15847 (N_15847,N_13327,N_12003);
xnor U15848 (N_15848,N_13522,N_13565);
nor U15849 (N_15849,N_13056,N_12427);
nand U15850 (N_15850,N_12598,N_12809);
nand U15851 (N_15851,N_12656,N_12382);
nor U15852 (N_15852,N_13096,N_12451);
nand U15853 (N_15853,N_13773,N_13461);
nand U15854 (N_15854,N_12689,N_13682);
nor U15855 (N_15855,N_12321,N_12282);
nor U15856 (N_15856,N_12191,N_12653);
xor U15857 (N_15857,N_13233,N_13038);
nand U15858 (N_15858,N_13889,N_13310);
or U15859 (N_15859,N_12361,N_12047);
and U15860 (N_15860,N_13768,N_12229);
xnor U15861 (N_15861,N_13796,N_13583);
or U15862 (N_15862,N_13580,N_13135);
xnor U15863 (N_15863,N_12598,N_13968);
or U15864 (N_15864,N_12630,N_13323);
nand U15865 (N_15865,N_12164,N_13092);
and U15866 (N_15866,N_12624,N_13497);
and U15867 (N_15867,N_12947,N_12615);
nor U15868 (N_15868,N_12564,N_13322);
or U15869 (N_15869,N_12672,N_13213);
nand U15870 (N_15870,N_12653,N_12309);
and U15871 (N_15871,N_13860,N_12013);
nand U15872 (N_15872,N_12301,N_13990);
nor U15873 (N_15873,N_13498,N_12984);
xor U15874 (N_15874,N_13998,N_13124);
nand U15875 (N_15875,N_12295,N_12688);
nand U15876 (N_15876,N_13506,N_13449);
nand U15877 (N_15877,N_12682,N_13884);
or U15878 (N_15878,N_13150,N_13283);
and U15879 (N_15879,N_12138,N_12205);
or U15880 (N_15880,N_12931,N_13634);
nand U15881 (N_15881,N_12151,N_13143);
nand U15882 (N_15882,N_12215,N_13298);
and U15883 (N_15883,N_12754,N_12003);
nand U15884 (N_15884,N_12199,N_13181);
nor U15885 (N_15885,N_12948,N_13617);
xor U15886 (N_15886,N_13714,N_12086);
nor U15887 (N_15887,N_13802,N_13381);
xor U15888 (N_15888,N_13402,N_12056);
nand U15889 (N_15889,N_12361,N_12159);
and U15890 (N_15890,N_12068,N_13456);
and U15891 (N_15891,N_13871,N_12247);
nand U15892 (N_15892,N_12057,N_12042);
nand U15893 (N_15893,N_12317,N_12381);
nand U15894 (N_15894,N_12956,N_12838);
xor U15895 (N_15895,N_12187,N_12959);
and U15896 (N_15896,N_13425,N_12114);
and U15897 (N_15897,N_13991,N_12168);
or U15898 (N_15898,N_12921,N_13785);
nor U15899 (N_15899,N_13228,N_12861);
nand U15900 (N_15900,N_13944,N_13328);
xnor U15901 (N_15901,N_12320,N_13276);
or U15902 (N_15902,N_12739,N_13479);
xor U15903 (N_15903,N_13749,N_12301);
or U15904 (N_15904,N_12113,N_13954);
nor U15905 (N_15905,N_13387,N_13219);
or U15906 (N_15906,N_13171,N_12840);
nor U15907 (N_15907,N_13340,N_12027);
nand U15908 (N_15908,N_13208,N_13173);
and U15909 (N_15909,N_13445,N_13528);
nand U15910 (N_15910,N_13305,N_13471);
and U15911 (N_15911,N_13342,N_12622);
xor U15912 (N_15912,N_13960,N_12851);
and U15913 (N_15913,N_12293,N_12905);
and U15914 (N_15914,N_13073,N_13133);
xnor U15915 (N_15915,N_13159,N_12966);
nor U15916 (N_15916,N_13857,N_13584);
xnor U15917 (N_15917,N_13785,N_13305);
and U15918 (N_15918,N_12392,N_13942);
nand U15919 (N_15919,N_12751,N_13358);
xnor U15920 (N_15920,N_12154,N_12572);
or U15921 (N_15921,N_12386,N_13401);
nor U15922 (N_15922,N_13513,N_12678);
or U15923 (N_15923,N_13653,N_12051);
nand U15924 (N_15924,N_12915,N_13607);
nand U15925 (N_15925,N_12251,N_12060);
or U15926 (N_15926,N_12482,N_13612);
xor U15927 (N_15927,N_13876,N_13678);
nor U15928 (N_15928,N_12359,N_13393);
and U15929 (N_15929,N_12687,N_12553);
or U15930 (N_15930,N_12275,N_13477);
or U15931 (N_15931,N_13046,N_12052);
nor U15932 (N_15932,N_12957,N_13896);
and U15933 (N_15933,N_13018,N_13737);
and U15934 (N_15934,N_12078,N_13345);
nand U15935 (N_15935,N_12302,N_13881);
nor U15936 (N_15936,N_13121,N_13306);
nor U15937 (N_15937,N_12700,N_12554);
xnor U15938 (N_15938,N_13209,N_13577);
xor U15939 (N_15939,N_13965,N_12850);
and U15940 (N_15940,N_12834,N_12332);
or U15941 (N_15941,N_12600,N_13482);
xnor U15942 (N_15942,N_12348,N_13058);
or U15943 (N_15943,N_12861,N_12431);
and U15944 (N_15944,N_12243,N_12629);
and U15945 (N_15945,N_12670,N_12648);
xor U15946 (N_15946,N_12682,N_13973);
nand U15947 (N_15947,N_13948,N_12217);
xnor U15948 (N_15948,N_13118,N_13052);
nand U15949 (N_15949,N_12064,N_12456);
or U15950 (N_15950,N_13455,N_12114);
or U15951 (N_15951,N_12007,N_12763);
xor U15952 (N_15952,N_12595,N_12859);
nand U15953 (N_15953,N_12551,N_13087);
or U15954 (N_15954,N_13200,N_13755);
and U15955 (N_15955,N_12022,N_12794);
nand U15956 (N_15956,N_13827,N_12139);
or U15957 (N_15957,N_13128,N_12500);
nand U15958 (N_15958,N_12567,N_13977);
nand U15959 (N_15959,N_13772,N_13223);
nand U15960 (N_15960,N_12365,N_13246);
xnor U15961 (N_15961,N_13019,N_13538);
and U15962 (N_15962,N_12417,N_13397);
nand U15963 (N_15963,N_13942,N_12985);
and U15964 (N_15964,N_13808,N_12051);
nor U15965 (N_15965,N_13839,N_13263);
nor U15966 (N_15966,N_13675,N_12965);
nand U15967 (N_15967,N_12931,N_13569);
or U15968 (N_15968,N_12231,N_13706);
xnor U15969 (N_15969,N_13138,N_12824);
nand U15970 (N_15970,N_13245,N_13164);
xnor U15971 (N_15971,N_13569,N_12317);
nand U15972 (N_15972,N_13033,N_13238);
xor U15973 (N_15973,N_13322,N_12562);
nor U15974 (N_15974,N_12015,N_12218);
nand U15975 (N_15975,N_12576,N_12373);
or U15976 (N_15976,N_12192,N_12970);
or U15977 (N_15977,N_13242,N_13517);
nand U15978 (N_15978,N_12240,N_13509);
nand U15979 (N_15979,N_13638,N_12794);
and U15980 (N_15980,N_12980,N_12146);
or U15981 (N_15981,N_13726,N_13457);
or U15982 (N_15982,N_13017,N_12021);
nor U15983 (N_15983,N_12728,N_12706);
nor U15984 (N_15984,N_12712,N_12582);
xor U15985 (N_15985,N_12731,N_12846);
or U15986 (N_15986,N_12737,N_13807);
nor U15987 (N_15987,N_13451,N_12424);
or U15988 (N_15988,N_13361,N_12271);
xor U15989 (N_15989,N_12044,N_12900);
or U15990 (N_15990,N_12372,N_13319);
and U15991 (N_15991,N_13650,N_12187);
nor U15992 (N_15992,N_12718,N_13498);
and U15993 (N_15993,N_12996,N_12586);
xnor U15994 (N_15994,N_12226,N_12550);
and U15995 (N_15995,N_13887,N_13449);
or U15996 (N_15996,N_12480,N_12894);
nand U15997 (N_15997,N_12356,N_13393);
nand U15998 (N_15998,N_13498,N_12245);
nor U15999 (N_15999,N_12464,N_13402);
and U16000 (N_16000,N_14438,N_15169);
xnor U16001 (N_16001,N_14238,N_14807);
nor U16002 (N_16002,N_14595,N_15778);
or U16003 (N_16003,N_15777,N_14952);
or U16004 (N_16004,N_14070,N_15592);
xor U16005 (N_16005,N_15679,N_14944);
or U16006 (N_16006,N_15109,N_15611);
or U16007 (N_16007,N_15924,N_15906);
and U16008 (N_16008,N_14061,N_15087);
nand U16009 (N_16009,N_14092,N_15500);
nand U16010 (N_16010,N_14085,N_15655);
or U16011 (N_16011,N_14527,N_14310);
nor U16012 (N_16012,N_14491,N_15352);
xor U16013 (N_16013,N_15652,N_15260);
nor U16014 (N_16014,N_15470,N_15650);
nand U16015 (N_16015,N_14671,N_15519);
xnor U16016 (N_16016,N_15090,N_14300);
and U16017 (N_16017,N_14764,N_15971);
xor U16018 (N_16018,N_15189,N_14689);
and U16019 (N_16019,N_15581,N_14261);
xor U16020 (N_16020,N_14776,N_14584);
xnor U16021 (N_16021,N_15337,N_15226);
nor U16022 (N_16022,N_14477,N_14251);
nor U16023 (N_16023,N_14763,N_15736);
nand U16024 (N_16024,N_15615,N_15153);
xor U16025 (N_16025,N_14194,N_15217);
or U16026 (N_16026,N_15218,N_14857);
or U16027 (N_16027,N_15911,N_15469);
or U16028 (N_16028,N_14606,N_15474);
and U16029 (N_16029,N_15496,N_14225);
and U16030 (N_16030,N_14531,N_15741);
or U16031 (N_16031,N_15306,N_14228);
xor U16032 (N_16032,N_14521,N_15892);
and U16033 (N_16033,N_15468,N_14887);
or U16034 (N_16034,N_15794,N_14710);
nand U16035 (N_16035,N_14983,N_15312);
and U16036 (N_16036,N_15871,N_14945);
xor U16037 (N_16037,N_14016,N_15811);
xnor U16038 (N_16038,N_15970,N_15098);
and U16039 (N_16039,N_14824,N_14991);
and U16040 (N_16040,N_14965,N_14856);
xor U16041 (N_16041,N_14153,N_14898);
nor U16042 (N_16042,N_15877,N_15332);
and U16043 (N_16043,N_15840,N_15094);
xor U16044 (N_16044,N_15585,N_14948);
nand U16045 (N_16045,N_14314,N_15651);
xor U16046 (N_16046,N_14534,N_14392);
and U16047 (N_16047,N_15683,N_14455);
or U16048 (N_16048,N_14968,N_14620);
nor U16049 (N_16049,N_15073,N_14789);
and U16050 (N_16050,N_14974,N_14291);
nor U16051 (N_16051,N_14217,N_14648);
nand U16052 (N_16052,N_15605,N_15026);
nand U16053 (N_16053,N_14193,N_14575);
nand U16054 (N_16054,N_14494,N_15543);
nand U16055 (N_16055,N_15419,N_14600);
or U16056 (N_16056,N_15542,N_15300);
and U16057 (N_16057,N_15873,N_14698);
nand U16058 (N_16058,N_14843,N_14057);
xor U16059 (N_16059,N_15205,N_14564);
nor U16060 (N_16060,N_14877,N_15015);
xnor U16061 (N_16061,N_14652,N_14559);
xor U16062 (N_16062,N_14592,N_15345);
nand U16063 (N_16063,N_14331,N_15942);
nand U16064 (N_16064,N_14554,N_15059);
and U16065 (N_16065,N_15768,N_14541);
or U16066 (N_16066,N_14465,N_14956);
nor U16067 (N_16067,N_14400,N_15621);
nor U16068 (N_16068,N_14267,N_15351);
or U16069 (N_16069,N_15359,N_14608);
nand U16070 (N_16070,N_15939,N_15759);
or U16071 (N_16071,N_15647,N_14731);
nand U16072 (N_16072,N_14551,N_15412);
nand U16073 (N_16073,N_15480,N_15701);
and U16074 (N_16074,N_15068,N_14044);
nor U16075 (N_16075,N_15163,N_14256);
nor U16076 (N_16076,N_15734,N_15688);
or U16077 (N_16077,N_15950,N_14986);
xnor U16078 (N_16078,N_15624,N_14495);
and U16079 (N_16079,N_15917,N_14663);
or U16080 (N_16080,N_15162,N_14177);
nor U16081 (N_16081,N_14389,N_15275);
or U16082 (N_16082,N_15618,N_15744);
nand U16083 (N_16083,N_15416,N_15267);
nand U16084 (N_16084,N_14703,N_15154);
nand U16085 (N_16085,N_14448,N_14647);
nand U16086 (N_16086,N_15274,N_15856);
nand U16087 (N_16087,N_14315,N_14918);
nor U16088 (N_16088,N_15248,N_14246);
and U16089 (N_16089,N_14988,N_15381);
nor U16090 (N_16090,N_14481,N_14659);
nor U16091 (N_16091,N_15635,N_15425);
or U16092 (N_16092,N_15780,N_15482);
and U16093 (N_16093,N_15358,N_15414);
nor U16094 (N_16094,N_15232,N_15121);
xor U16095 (N_16095,N_14621,N_15423);
nor U16096 (N_16096,N_15545,N_14169);
nor U16097 (N_16097,N_15727,N_14915);
or U16098 (N_16098,N_15712,N_15437);
and U16099 (N_16099,N_15531,N_14394);
nand U16100 (N_16100,N_15057,N_15161);
nand U16101 (N_16101,N_14462,N_15724);
nor U16102 (N_16102,N_14355,N_14733);
and U16103 (N_16103,N_14650,N_14087);
and U16104 (N_16104,N_15401,N_15338);
nor U16105 (N_16105,N_14207,N_15674);
nand U16106 (N_16106,N_15321,N_15852);
nand U16107 (N_16107,N_15051,N_15328);
xnor U16108 (N_16108,N_14978,N_14697);
nand U16109 (N_16109,N_14399,N_15739);
xnor U16110 (N_16110,N_15032,N_14667);
nand U16111 (N_16111,N_14132,N_15834);
xnor U16112 (N_16112,N_14961,N_15822);
nand U16113 (N_16113,N_14295,N_15965);
nand U16114 (N_16114,N_15999,N_14138);
and U16115 (N_16115,N_15870,N_14955);
nor U16116 (N_16116,N_14290,N_15932);
or U16117 (N_16117,N_14405,N_14017);
and U16118 (N_16118,N_14249,N_15014);
or U16119 (N_16119,N_14736,N_15633);
and U16120 (N_16120,N_15012,N_15748);
xnor U16121 (N_16121,N_14076,N_15272);
or U16122 (N_16122,N_14230,N_14591);
xnor U16123 (N_16123,N_15879,N_15540);
nor U16124 (N_16124,N_14363,N_15361);
and U16125 (N_16125,N_15796,N_15456);
nor U16126 (N_16126,N_15910,N_14082);
nor U16127 (N_16127,N_14084,N_14641);
or U16128 (N_16128,N_14243,N_15681);
or U16129 (N_16129,N_14189,N_14094);
xor U16130 (N_16130,N_14938,N_15536);
and U16131 (N_16131,N_14254,N_14599);
and U16132 (N_16132,N_14456,N_14135);
nor U16133 (N_16133,N_14274,N_14432);
and U16134 (N_16134,N_15256,N_14439);
and U16135 (N_16135,N_15080,N_15640);
nor U16136 (N_16136,N_14859,N_14739);
nand U16137 (N_16137,N_15622,N_15983);
nand U16138 (N_16138,N_15367,N_15630);
and U16139 (N_16139,N_15296,N_15704);
and U16140 (N_16140,N_15065,N_15603);
and U16141 (N_16141,N_14014,N_15411);
and U16142 (N_16142,N_15063,N_15926);
or U16143 (N_16143,N_15703,N_14939);
and U16144 (N_16144,N_15956,N_14008);
or U16145 (N_16145,N_15067,N_15718);
xor U16146 (N_16146,N_14007,N_15857);
xor U16147 (N_16147,N_14519,N_14645);
or U16148 (N_16148,N_14990,N_15092);
or U16149 (N_16149,N_14120,N_15392);
or U16150 (N_16150,N_14700,N_14572);
xnor U16151 (N_16151,N_14513,N_15571);
xnor U16152 (N_16152,N_15476,N_15442);
xnor U16153 (N_16153,N_14660,N_15225);
or U16154 (N_16154,N_15707,N_14340);
nand U16155 (N_16155,N_14910,N_14335);
and U16156 (N_16156,N_14470,N_14875);
nand U16157 (N_16157,N_15071,N_14505);
nand U16158 (N_16158,N_15935,N_14619);
nor U16159 (N_16159,N_15667,N_14508);
and U16160 (N_16160,N_14374,N_15731);
nor U16161 (N_16161,N_14878,N_15875);
xor U16162 (N_16162,N_14587,N_15363);
xor U16163 (N_16163,N_15504,N_15390);
or U16164 (N_16164,N_14269,N_14270);
and U16165 (N_16165,N_15963,N_15379);
or U16166 (N_16166,N_15064,N_15758);
or U16167 (N_16167,N_14283,N_15675);
nand U16168 (N_16168,N_15610,N_15058);
nor U16169 (N_16169,N_15607,N_14576);
and U16170 (N_16170,N_15116,N_15659);
or U16171 (N_16171,N_14742,N_14760);
nor U16172 (N_16172,N_14123,N_15544);
and U16173 (N_16173,N_14743,N_14024);
nor U16174 (N_16174,N_14629,N_15548);
and U16175 (N_16175,N_15502,N_15207);
or U16176 (N_16176,N_15334,N_14571);
nand U16177 (N_16177,N_15881,N_14717);
xnor U16178 (N_16178,N_14560,N_15961);
xor U16179 (N_16179,N_15353,N_14906);
xnor U16180 (N_16180,N_15402,N_15564);
and U16181 (N_16181,N_14771,N_15042);
nand U16182 (N_16182,N_15027,N_15342);
and U16183 (N_16183,N_15993,N_14239);
or U16184 (N_16184,N_15103,N_15937);
xor U16185 (N_16185,N_15096,N_15899);
xor U16186 (N_16186,N_14210,N_14449);
or U16187 (N_16187,N_14370,N_15649);
nand U16188 (N_16188,N_15770,N_14036);
or U16189 (N_16189,N_14000,N_15427);
nor U16190 (N_16190,N_14369,N_15959);
or U16191 (N_16191,N_14478,N_15355);
and U16192 (N_16192,N_14826,N_14860);
xnor U16193 (N_16193,N_15966,N_15553);
and U16194 (N_16194,N_14607,N_15938);
nor U16195 (N_16195,N_14218,N_15575);
or U16196 (N_16196,N_15754,N_15897);
xnor U16197 (N_16197,N_14488,N_14737);
xor U16198 (N_16198,N_15830,N_15805);
nand U16199 (N_16199,N_14330,N_15717);
nand U16200 (N_16200,N_15900,N_15927);
xnor U16201 (N_16201,N_14065,N_14053);
nand U16202 (N_16202,N_15286,N_14015);
nor U16203 (N_16203,N_15185,N_15998);
nand U16204 (N_16204,N_15273,N_14440);
xnor U16205 (N_16205,N_15224,N_14640);
and U16206 (N_16206,N_14281,N_14287);
nand U16207 (N_16207,N_15577,N_15011);
nand U16208 (N_16208,N_15580,N_15319);
nand U16209 (N_16209,N_14302,N_15197);
nand U16210 (N_16210,N_15645,N_14474);
or U16211 (N_16211,N_15453,N_14905);
nand U16212 (N_16212,N_15271,N_14435);
nand U16213 (N_16213,N_14711,N_14581);
nor U16214 (N_16214,N_15643,N_14954);
or U16215 (N_16215,N_14540,N_14496);
nor U16216 (N_16216,N_14598,N_15831);
and U16217 (N_16217,N_14543,N_15559);
or U16218 (N_16218,N_15085,N_15141);
and U16219 (N_16219,N_15955,N_14402);
and U16220 (N_16220,N_15343,N_14917);
or U16221 (N_16221,N_15046,N_15409);
xnor U16222 (N_16222,N_15658,N_15820);
and U16223 (N_16223,N_14786,N_15590);
xor U16224 (N_16224,N_14473,N_15044);
or U16225 (N_16225,N_15295,N_15054);
xnor U16226 (N_16226,N_15293,N_15018);
and U16227 (N_16227,N_14761,N_15627);
nor U16228 (N_16228,N_14196,N_15378);
xnor U16229 (N_16229,N_14770,N_14732);
nand U16230 (N_16230,N_15019,N_15920);
xor U16231 (N_16231,N_15428,N_15804);
nand U16232 (N_16232,N_15093,N_14908);
and U16233 (N_16233,N_14755,N_15960);
or U16234 (N_16234,N_14212,N_14959);
nand U16235 (N_16235,N_15006,N_15002);
or U16236 (N_16236,N_15866,N_14814);
xor U16237 (N_16237,N_14104,N_15130);
nor U16238 (N_16238,N_14977,N_14025);
and U16239 (N_16239,N_14268,N_14767);
nor U16240 (N_16240,N_14923,N_15750);
or U16241 (N_16241,N_15843,N_14371);
nand U16242 (N_16242,N_14951,N_14561);
xor U16243 (N_16243,N_14326,N_14021);
and U16244 (N_16244,N_14806,N_14117);
xnor U16245 (N_16245,N_15538,N_15994);
nor U16246 (N_16246,N_14886,N_14289);
nand U16247 (N_16247,N_14683,N_15311);
xor U16248 (N_16248,N_14034,N_14837);
nand U16249 (N_16249,N_14907,N_14900);
and U16250 (N_16250,N_14458,N_15576);
nor U16251 (N_16251,N_15166,N_14811);
nand U16252 (N_16252,N_14817,N_14553);
xnor U16253 (N_16253,N_14026,N_14067);
or U16254 (N_16254,N_15240,N_15516);
nand U16255 (N_16255,N_14976,N_14752);
xor U16256 (N_16256,N_15765,N_14188);
nand U16257 (N_16257,N_15336,N_15007);
or U16258 (N_16258,N_15714,N_15431);
and U16259 (N_16259,N_14597,N_14216);
xnor U16260 (N_16260,N_14115,N_14921);
nand U16261 (N_16261,N_15746,N_14728);
nor U16262 (N_16262,N_14029,N_14863);
or U16263 (N_16263,N_15565,N_14497);
or U16264 (N_16264,N_15833,N_15716);
xor U16265 (N_16265,N_15394,N_15405);
or U16266 (N_16266,N_14181,N_14866);
nand U16267 (N_16267,N_15572,N_14294);
or U16268 (N_16268,N_14143,N_14799);
and U16269 (N_16269,N_15666,N_15033);
or U16270 (N_16270,N_15255,N_15061);
or U16271 (N_16271,N_14902,N_15030);
xor U16272 (N_16272,N_14680,N_15634);
nor U16273 (N_16273,N_14825,N_14932);
and U16274 (N_16274,N_14804,N_15884);
nand U16275 (N_16275,N_15299,N_14089);
xnor U16276 (N_16276,N_15689,N_15948);
nor U16277 (N_16277,N_15612,N_14631);
nand U16278 (N_16278,N_15458,N_14338);
and U16279 (N_16279,N_15609,N_15056);
and U16280 (N_16280,N_15546,N_14174);
and U16281 (N_16281,N_14694,N_15368);
nand U16282 (N_16282,N_14077,N_15113);
nand U16283 (N_16283,N_14293,N_14499);
xor U16284 (N_16284,N_14844,N_14199);
or U16285 (N_16285,N_15028,N_14219);
nand U16286 (N_16286,N_14846,N_14872);
xor U16287 (N_16287,N_14782,N_14422);
or U16288 (N_16288,N_15172,N_14260);
nor U16289 (N_16289,N_14151,N_14202);
xnor U16290 (N_16290,N_14420,N_15975);
and U16291 (N_16291,N_15354,N_15931);
xnor U16292 (N_16292,N_14333,N_15620);
nor U16293 (N_16293,N_15479,N_14232);
xor U16294 (N_16294,N_15554,N_15824);
xnor U16295 (N_16295,N_14276,N_14453);
and U16296 (N_16296,N_14937,N_14266);
xor U16297 (N_16297,N_14913,N_15880);
nor U16298 (N_16298,N_14914,N_14653);
or U16299 (N_16299,N_14768,N_15287);
and U16300 (N_16300,N_14288,N_14022);
xnor U16301 (N_16301,N_15426,N_14766);
nor U16302 (N_16302,N_15761,N_15471);
and U16303 (N_16303,N_14351,N_14836);
or U16304 (N_16304,N_15159,N_14842);
nand U16305 (N_16305,N_15639,N_14769);
or U16306 (N_16306,N_15219,N_15753);
nand U16307 (N_16307,N_14103,N_14615);
xor U16308 (N_16308,N_15529,N_15115);
or U16309 (N_16309,N_14433,N_14633);
and U16310 (N_16310,N_14383,N_15896);
xnor U16311 (N_16311,N_14055,N_14108);
and U16312 (N_16312,N_14729,N_14040);
and U16313 (N_16313,N_14626,N_14975);
nor U16314 (N_16314,N_15292,N_15922);
nand U16315 (N_16315,N_15827,N_14275);
and U16316 (N_16316,N_14450,N_14662);
nor U16317 (N_16317,N_14144,N_15430);
nand U16318 (N_16318,N_15081,N_15454);
and U16319 (N_16319,N_15636,N_15493);
xnor U16320 (N_16320,N_14911,N_15472);
xnor U16321 (N_16321,N_15140,N_14931);
and U16322 (N_16322,N_15783,N_14614);
and U16323 (N_16323,N_14655,N_15752);
or U16324 (N_16324,N_15608,N_15258);
nand U16325 (N_16325,N_14447,N_15791);
nor U16326 (N_16326,N_14419,N_15563);
and U16327 (N_16327,N_14198,N_14401);
nand U16328 (N_16328,N_14573,N_15503);
nor U16329 (N_16329,N_14444,N_15766);
nand U16330 (N_16330,N_14539,N_14727);
and U16331 (N_16331,N_15281,N_15771);
and U16332 (N_16332,N_15957,N_15000);
or U16333 (N_16333,N_14979,N_14498);
and U16334 (N_16334,N_15370,N_14642);
nand U16335 (N_16335,N_14110,N_14095);
nand U16336 (N_16336,N_15194,N_14895);
xnor U16337 (N_16337,N_14052,N_15558);
xnor U16338 (N_16338,N_15829,N_14738);
nor U16339 (N_16339,N_14482,N_15747);
xor U16340 (N_16340,N_15672,N_15541);
xnor U16341 (N_16341,N_14154,N_14899);
and U16342 (N_16342,N_14639,N_14841);
or U16343 (N_16343,N_14759,N_15013);
and U16344 (N_16344,N_14884,N_14503);
nand U16345 (N_16345,N_15216,N_14118);
nor U16346 (N_16346,N_14791,N_14066);
nand U16347 (N_16347,N_14031,N_15097);
or U16348 (N_16348,N_14244,N_15127);
or U16349 (N_16349,N_14590,N_14721);
nor U16350 (N_16350,N_14226,N_14828);
nand U16351 (N_16351,N_14970,N_14183);
and U16352 (N_16352,N_15726,N_15719);
or U16353 (N_16353,N_14972,N_15798);
and U16354 (N_16354,N_15117,N_15821);
nand U16355 (N_16355,N_14708,N_14876);
or U16356 (N_16356,N_14083,N_15534);
nand U16357 (N_16357,N_14427,N_15720);
and U16358 (N_16358,N_14492,N_14039);
or U16359 (N_16359,N_14953,N_15797);
or U16360 (N_16360,N_15763,N_14585);
or U16361 (N_16361,N_15532,N_15158);
xnor U16362 (N_16362,N_15322,N_15291);
xnor U16363 (N_16363,N_14546,N_15452);
nand U16364 (N_16364,N_14041,N_14681);
xnor U16365 (N_16365,N_15816,N_14547);
nor U16366 (N_16366,N_15555,N_14201);
nor U16367 (N_16367,N_15523,N_14670);
nor U16368 (N_16368,N_15987,N_14715);
xnor U16369 (N_16369,N_14853,N_14012);
nor U16370 (N_16370,N_14957,N_14725);
nor U16371 (N_16371,N_14549,N_14509);
and U16372 (N_16372,N_15526,N_14033);
nor U16373 (N_16373,N_14054,N_15799);
or U16374 (N_16374,N_14718,N_15415);
or U16375 (N_16375,N_14308,N_14479);
nor U16376 (N_16376,N_14064,N_15953);
nor U16377 (N_16377,N_15732,N_14685);
and U16378 (N_16378,N_14090,N_14442);
nand U16379 (N_16379,N_14272,N_14168);
nor U16380 (N_16380,N_14726,N_14709);
nor U16381 (N_16381,N_15586,N_14386);
nor U16382 (N_16382,N_15290,N_14296);
nand U16383 (N_16383,N_15661,N_15108);
xor U16384 (N_16384,N_14320,N_15396);
nor U16385 (N_16385,N_15330,N_14045);
and U16386 (N_16386,N_14765,N_15992);
nand U16387 (N_16387,N_15515,N_15035);
or U16388 (N_16388,N_14920,N_15835);
xnor U16389 (N_16389,N_15270,N_15421);
xor U16390 (N_16390,N_15184,N_14963);
xor U16391 (N_16391,N_15076,N_15233);
or U16392 (N_16392,N_14529,N_14839);
xnor U16393 (N_16393,N_15024,N_15253);
or U16394 (N_16394,N_14037,N_14312);
or U16395 (N_16395,N_14942,N_15118);
nand U16396 (N_16396,N_14062,N_14705);
xor U16397 (N_16397,N_15213,N_15933);
nor U16398 (N_16398,N_15851,N_14368);
nor U16399 (N_16399,N_14879,N_15190);
nor U16400 (N_16400,N_14426,N_14517);
nor U16401 (N_16401,N_15512,N_14880);
nor U16402 (N_16402,N_14992,N_15022);
or U16403 (N_16403,N_14617,N_14416);
nor U16404 (N_16404,N_14851,N_15560);
or U16405 (N_16405,N_14903,N_15340);
nor U16406 (N_16406,N_15786,N_15946);
xnor U16407 (N_16407,N_15393,N_14236);
and U16408 (N_16408,N_15303,N_15745);
nand U16409 (N_16409,N_14993,N_14332);
xnor U16410 (N_16410,N_14930,N_15702);
xnor U16411 (N_16411,N_15613,N_14486);
or U16412 (N_16412,N_14167,N_14441);
xor U16413 (N_16413,N_15451,N_15008);
nor U16414 (N_16414,N_15883,N_15305);
or U16415 (N_16415,N_15878,N_14885);
and U16416 (N_16416,N_15201,N_15671);
nand U16417 (N_16417,N_15461,N_14396);
and U16418 (N_16418,N_15004,N_15242);
xor U16419 (N_16419,N_14306,N_15606);
nor U16420 (N_16420,N_15574,N_14632);
xnor U16421 (N_16421,N_15079,N_14612);
nor U16422 (N_16422,N_15823,N_15849);
xor U16423 (N_16423,N_14313,N_14861);
xnor U16424 (N_16424,N_15773,N_14317);
xor U16425 (N_16425,N_15254,N_15914);
nand U16426 (N_16426,N_14801,N_14203);
or U16427 (N_16427,N_14073,N_14934);
nand U16428 (N_16428,N_14748,N_15517);
nor U16429 (N_16429,N_14460,N_15637);
xnor U16430 (N_16430,N_15069,N_14746);
or U16431 (N_16431,N_15890,N_14162);
or U16432 (N_16432,N_14278,N_14137);
or U16433 (N_16433,N_14596,N_15980);
xor U16434 (N_16434,N_14686,N_14195);
nor U16435 (N_16435,N_14161,N_15737);
or U16436 (N_16436,N_14344,N_15694);
nor U16437 (N_16437,N_14179,N_15733);
nor U16438 (N_16438,N_15530,N_15440);
xor U16439 (N_16439,N_14941,N_14343);
nor U16440 (N_16440,N_15302,N_14637);
nand U16441 (N_16441,N_15148,N_14809);
nand U16442 (N_16442,N_15839,N_14381);
and U16443 (N_16443,N_14305,N_14068);
nand U16444 (N_16444,N_14613,N_14247);
and U16445 (N_16445,N_15095,N_14004);
xor U16446 (N_16446,N_15101,N_15335);
nand U16447 (N_16447,N_15297,N_14520);
nor U16448 (N_16448,N_14373,N_14971);
nor U16449 (N_16449,N_15528,N_15863);
xnor U16450 (N_16450,N_14157,N_14538);
nor U16451 (N_16451,N_15350,N_14901);
and U16452 (N_16452,N_15749,N_15447);
xnor U16453 (N_16453,N_14960,N_14578);
nand U16454 (N_16454,N_15868,N_14661);
nand U16455 (N_16455,N_15601,N_15170);
and U16456 (N_16456,N_15133,N_14156);
or U16457 (N_16457,N_15844,N_14778);
and U16458 (N_16458,N_14796,N_15903);
xnor U16459 (N_16459,N_14235,N_14241);
xor U16460 (N_16460,N_15860,N_15484);
nand U16461 (N_16461,N_14248,N_15916);
nor U16462 (N_16462,N_14060,N_15331);
xor U16463 (N_16463,N_15584,N_14186);
nor U16464 (N_16464,N_14468,N_14208);
and U16465 (N_16465,N_15664,N_15874);
xnor U16466 (N_16466,N_14506,N_15762);
nor U16467 (N_16467,N_15188,N_14904);
or U16468 (N_16468,N_14601,N_14020);
or U16469 (N_16469,N_15438,N_15083);
nor U16470 (N_16470,N_15323,N_15245);
or U16471 (N_16471,N_14795,N_15969);
xnor U16472 (N_16472,N_15236,N_14712);
xnor U16473 (N_16473,N_14081,N_15356);
nand U16474 (N_16474,N_15991,N_15524);
or U16475 (N_16475,N_15176,N_15173);
and U16476 (N_16476,N_15373,N_14802);
nand U16477 (N_16477,N_15325,N_15930);
nor U16478 (N_16478,N_15537,N_15889);
xor U16479 (N_16479,N_15589,N_14471);
nor U16480 (N_16480,N_15498,N_14178);
and U16481 (N_16481,N_15481,N_14562);
xor U16482 (N_16482,N_15697,N_14229);
or U16483 (N_16483,N_15962,N_14329);
nand U16484 (N_16484,N_15155,N_15923);
or U16485 (N_16485,N_15143,N_14750);
xor U16486 (N_16486,N_14056,N_14740);
and U16487 (N_16487,N_14365,N_14443);
and U16488 (N_16488,N_14522,N_15049);
xnor U16489 (N_16489,N_14451,N_15348);
xor U16490 (N_16490,N_15138,N_15055);
xor U16491 (N_16491,N_15790,N_14676);
nor U16492 (N_16492,N_14526,N_15106);
nand U16493 (N_16493,N_14382,N_14150);
nor U16494 (N_16494,N_15776,N_14867);
or U16495 (N_16495,N_15550,N_15964);
nand U16496 (N_16496,N_15787,N_14530);
or U16497 (N_16497,N_15149,N_14935);
nor U16498 (N_16498,N_15417,N_15867);
xnor U16499 (N_16499,N_15486,N_15713);
and U16500 (N_16500,N_15317,N_14500);
xor U16501 (N_16501,N_15501,N_15886);
nor U16502 (N_16502,N_14466,N_14030);
nor U16503 (N_16503,N_15673,N_15365);
nand U16504 (N_16504,N_15641,N_14088);
nand U16505 (N_16505,N_14490,N_15380);
nor U16506 (N_16506,N_15246,N_15204);
and U16507 (N_16507,N_15507,N_15105);
nor U16508 (N_16508,N_15465,N_15156);
nand U16509 (N_16509,N_14558,N_14051);
xnor U16510 (N_16510,N_14475,N_14175);
xor U16511 (N_16511,N_15743,N_14618);
or U16512 (N_16512,N_14398,N_14038);
and U16513 (N_16513,N_15395,N_15110);
or U16514 (N_16514,N_15132,N_15842);
xnor U16515 (N_16515,N_15066,N_14140);
nor U16516 (N_16516,N_15339,N_15135);
nor U16517 (N_16517,N_15757,N_14518);
nor U16518 (N_16518,N_15146,N_14385);
xor U16519 (N_16519,N_15509,N_14569);
xnor U16520 (N_16520,N_14924,N_14155);
xnor U16521 (N_16521,N_14469,N_14797);
nand U16522 (N_16522,N_14644,N_14950);
nor U16523 (N_16523,N_14234,N_14744);
or U16524 (N_16524,N_15539,N_14311);
nor U16525 (N_16525,N_14749,N_14545);
nor U16526 (N_16526,N_15264,N_14820);
nor U16527 (N_16527,N_14724,N_14656);
xor U16528 (N_16528,N_14100,N_14042);
nor U16529 (N_16529,N_15375,N_14158);
nand U16530 (N_16530,N_15594,N_14322);
and U16531 (N_16531,N_14130,N_14893);
nand U16532 (N_16532,N_15628,N_14136);
xor U16533 (N_16533,N_15177,N_15855);
xnor U16534 (N_16534,N_14318,N_15187);
nor U16535 (N_16535,N_14048,N_15239);
and U16536 (N_16536,N_14783,N_14428);
and U16537 (N_16537,N_14605,N_15439);
nor U16538 (N_16538,N_15632,N_14695);
and U16539 (N_16539,N_15145,N_15040);
nor U16540 (N_16540,N_14299,N_15485);
nand U16541 (N_16541,N_15052,N_15846);
and U16542 (N_16542,N_15220,N_15795);
xnor U16543 (N_16543,N_14128,N_14745);
and U16544 (N_16544,N_14069,N_15711);
and U16545 (N_16545,N_14696,N_14831);
xor U16546 (N_16546,N_14962,N_15789);
or U16547 (N_16547,N_15898,N_15385);
or U16548 (N_16548,N_14404,N_14616);
xor U16549 (N_16549,N_14211,N_15785);
nand U16550 (N_16550,N_15832,N_15656);
nor U16551 (N_16551,N_14909,N_14565);
xnor U16552 (N_16552,N_14429,N_14995);
nor U16553 (N_16553,N_14714,N_15915);
and U16554 (N_16554,N_15648,N_14304);
and U16555 (N_16555,N_14634,N_14342);
or U16556 (N_16556,N_15075,N_15284);
xnor U16557 (N_16557,N_15619,N_15668);
nor U16558 (N_16558,N_14690,N_14532);
nand U16559 (N_16559,N_15089,N_14536);
and U16560 (N_16560,N_14049,N_15782);
and U16561 (N_16561,N_15048,N_15403);
and U16562 (N_16562,N_15237,N_15693);
nand U16563 (N_16563,N_14032,N_14704);
nor U16564 (N_16564,N_15151,N_14145);
nand U16565 (N_16565,N_14139,N_14301);
nor U16566 (N_16566,N_14947,N_14414);
nand U16567 (N_16567,N_14431,N_15644);
nand U16568 (N_16568,N_15617,N_15326);
and U16569 (N_16569,N_15828,N_15588);
or U16570 (N_16570,N_15706,N_14346);
xor U16571 (N_16571,N_15696,N_14542);
nand U16572 (N_16572,N_14929,N_14604);
xor U16573 (N_16573,N_14699,N_15912);
nor U16574 (N_16574,N_15781,N_15690);
nor U16575 (N_16575,N_15372,N_14933);
nor U16576 (N_16576,N_15979,N_14417);
xnor U16577 (N_16577,N_15371,N_14756);
nor U16578 (N_16578,N_14013,N_15837);
nor U16579 (N_16579,N_15045,N_14116);
and U16580 (N_16580,N_14949,N_14713);
xor U16581 (N_16581,N_15985,N_15397);
and U16582 (N_16582,N_14125,N_14222);
or U16583 (N_16583,N_15277,N_14537);
xor U16584 (N_16584,N_15017,N_14325);
nand U16585 (N_16585,N_15025,N_14829);
nand U16586 (N_16586,N_15769,N_15244);
nand U16587 (N_16587,N_15573,N_14446);
xor U16588 (N_16588,N_15010,N_14058);
xor U16589 (N_16589,N_14982,N_15945);
nor U16590 (N_16590,N_15060,N_15142);
xnor U16591 (N_16591,N_14926,N_15623);
or U16592 (N_16592,N_15891,N_15990);
nand U16593 (N_16593,N_14425,N_15386);
or U16594 (N_16594,N_14579,N_14485);
or U16595 (N_16595,N_14362,N_15200);
and U16596 (N_16596,N_14354,N_15131);
nand U16597 (N_16597,N_14206,N_15266);
nor U16598 (N_16598,N_14946,N_15413);
and U16599 (N_16599,N_14327,N_15308);
or U16600 (N_16600,N_14421,N_15525);
nor U16601 (N_16601,N_15626,N_15947);
nor U16602 (N_16602,N_14515,N_15663);
or U16603 (N_16603,N_15228,N_14091);
or U16604 (N_16604,N_14258,N_14191);
nor U16605 (N_16605,N_14847,N_14324);
and U16606 (N_16606,N_15788,N_14121);
nor U16607 (N_16607,N_15968,N_15865);
or U16608 (N_16608,N_15784,N_15708);
nor U16609 (N_16609,N_14735,N_14262);
nor U16610 (N_16610,N_15099,N_14566);
nor U16611 (N_16611,N_15949,N_15209);
and U16612 (N_16612,N_14664,N_15175);
or U16613 (N_16613,N_15112,N_15494);
nor U16614 (N_16614,N_15180,N_15477);
and U16615 (N_16615,N_14775,N_14307);
and U16616 (N_16616,N_14205,N_14334);
or U16617 (N_16617,N_15203,N_15557);
and U16618 (N_16618,N_15001,N_15329);
or U16619 (N_16619,N_14556,N_15511);
and U16620 (N_16620,N_15806,N_14464);
or U16621 (N_16621,N_15241,N_15347);
xor U16622 (N_16622,N_14454,N_15301);
xnor U16623 (N_16623,N_14003,N_14674);
and U16624 (N_16624,N_15041,N_15178);
nor U16625 (N_16625,N_14544,N_15808);
nor U16626 (N_16626,N_14122,N_14411);
and U16627 (N_16627,N_15404,N_15122);
nand U16628 (N_16628,N_15801,N_15850);
and U16629 (N_16629,N_14784,N_14883);
or U16630 (N_16630,N_15384,N_15756);
and U16631 (N_16631,N_14570,N_14163);
or U16632 (N_16632,N_14722,N_14927);
or U16633 (N_16633,N_15597,N_15196);
nor U16634 (N_16634,N_14668,N_14434);
and U16635 (N_16635,N_14577,N_15918);
or U16636 (N_16636,N_15441,N_15362);
and U16637 (N_16637,N_14119,N_15072);
nand U16638 (N_16638,N_14651,N_14366);
nor U16639 (N_16639,N_15104,N_15377);
nor U16640 (N_16640,N_14423,N_15518);
or U16641 (N_16641,N_14146,N_15520);
xor U16642 (N_16642,N_15685,N_15872);
or U16643 (N_16643,N_15313,N_14849);
nand U16644 (N_16644,N_14723,N_14430);
or U16645 (N_16645,N_15646,N_15206);
nand U16646 (N_16646,N_15802,N_14666);
and U16647 (N_16647,N_14827,N_15705);
or U16648 (N_16648,N_14574,N_14582);
and U16649 (N_16649,N_15760,N_15406);
and U16650 (N_16650,N_14336,N_15893);
and U16651 (N_16651,N_14981,N_14046);
and U16652 (N_16652,N_14213,N_14510);
xnor U16653 (N_16653,N_15819,N_15445);
and U16654 (N_16654,N_15029,N_14758);
or U16655 (N_16655,N_14535,N_14567);
nand U16656 (N_16656,N_15210,N_14476);
nor U16657 (N_16657,N_15229,N_15876);
nand U16658 (N_16658,N_15152,N_14372);
xor U16659 (N_16659,N_15021,N_14649);
nand U16660 (N_16660,N_14245,N_14989);
xor U16661 (N_16661,N_15126,N_14943);
xnor U16662 (N_16662,N_14461,N_15136);
nand U16663 (N_16663,N_15315,N_14376);
nand U16664 (N_16664,N_15547,N_14487);
nor U16665 (N_16665,N_14502,N_15324);
or U16666 (N_16666,N_14098,N_14360);
or U16667 (N_16667,N_15450,N_14380);
nor U16668 (N_16668,N_15629,N_15989);
nand U16669 (N_16669,N_14242,N_14928);
or U16670 (N_16670,N_15977,N_14684);
or U16671 (N_16671,N_14028,N_14353);
and U16672 (N_16672,N_14316,N_14716);
nor U16673 (N_16673,N_15952,N_14273);
or U16674 (N_16674,N_15457,N_14457);
nor U16675 (N_16675,N_15813,N_15909);
nor U16676 (N_16676,N_15552,N_15344);
and U16677 (N_16677,N_14215,N_15742);
or U16678 (N_16678,N_15692,N_14757);
and U16679 (N_16679,N_15958,N_15227);
nand U16680 (N_16680,N_14832,N_14821);
nor U16681 (N_16681,N_15139,N_14164);
or U16682 (N_16682,N_14852,N_15399);
or U16683 (N_16683,N_14730,N_14171);
or U16684 (N_16684,N_15815,N_14277);
or U16685 (N_16685,N_14912,N_14265);
nor U16686 (N_16686,N_14610,N_15578);
nand U16687 (N_16687,N_15091,N_15684);
and U16688 (N_16688,N_15566,N_15463);
or U16689 (N_16689,N_14204,N_15114);
xor U16690 (N_16690,N_14808,N_15967);
and U16691 (N_16691,N_15374,N_15709);
xor U16692 (N_16692,N_14964,N_15662);
or U16693 (N_16693,N_15279,N_15549);
nand U16694 (N_16694,N_15077,N_14395);
nor U16695 (N_16695,N_15826,N_15818);
nor U16696 (N_16696,N_15680,N_15280);
or U16697 (N_16697,N_14657,N_14378);
xor U16698 (N_16698,N_14794,N_15464);
and U16699 (N_16699,N_15179,N_14793);
xnor U16700 (N_16700,N_15513,N_15252);
nand U16701 (N_16701,N_14557,N_14868);
and U16702 (N_16702,N_15941,N_14999);
nand U16703 (N_16703,N_14958,N_14452);
or U16704 (N_16704,N_15888,N_15288);
or U16705 (N_16705,N_14658,N_15848);
and U16706 (N_16706,N_15665,N_15023);
xnor U16707 (N_16707,N_14890,N_15310);
and U16708 (N_16708,N_14609,N_14359);
nand U16709 (N_16709,N_15568,N_14285);
or U16710 (N_16710,N_15186,N_14747);
or U16711 (N_16711,N_14093,N_15729);
nor U16712 (N_16712,N_14005,N_15120);
nor U16713 (N_16713,N_15304,N_14638);
nor U16714 (N_16714,N_15653,N_15625);
nor U16715 (N_16715,N_15100,N_14822);
nor U16716 (N_16716,N_14840,N_14341);
nand U16717 (N_16717,N_15369,N_15111);
xor U16718 (N_16718,N_15247,N_14321);
nor U16719 (N_16719,N_14413,N_15614);
or U16720 (N_16720,N_15212,N_14691);
and U16721 (N_16721,N_14504,N_14319);
xor U16722 (N_16722,N_14114,N_14071);
xor U16723 (N_16723,N_15215,N_14436);
and U16724 (N_16724,N_15487,N_14966);
or U16725 (N_16725,N_14984,N_15676);
and U16726 (N_16726,N_15869,N_14862);
nor U16727 (N_16727,N_15424,N_15074);
xor U16728 (N_16728,N_15198,N_14101);
and U16729 (N_16729,N_14160,N_15462);
nor U16730 (N_16730,N_14501,N_14525);
nand U16731 (N_16731,N_15533,N_15853);
nand U16732 (N_16732,N_15919,N_15521);
xnor U16733 (N_16733,N_14568,N_14390);
nor U16734 (N_16734,N_15309,N_15506);
or U16735 (N_16735,N_15974,N_15388);
and U16736 (N_16736,N_14264,N_14550);
xor U16737 (N_16737,N_15984,N_15429);
and U16738 (N_16738,N_15157,N_15020);
or U16739 (N_16739,N_14969,N_14009);
nor U16740 (N_16740,N_14643,N_14480);
nand U16741 (N_16741,N_15642,N_15208);
and U16742 (N_16742,N_14611,N_15660);
nor U16743 (N_16743,N_14922,N_15887);
nor U16744 (N_16744,N_14253,N_15738);
nor U16745 (N_16745,N_15710,N_14096);
or U16746 (N_16746,N_15183,N_14896);
or U16747 (N_16747,N_14850,N_15807);
nor U16748 (N_16748,N_15638,N_14985);
nor U16749 (N_16749,N_15202,N_15483);
and U16750 (N_16750,N_15591,N_14309);
or U16751 (N_16751,N_14339,N_14019);
nand U16752 (N_16752,N_15257,N_15191);
nand U16753 (N_16753,N_14864,N_14833);
xor U16754 (N_16754,N_15398,N_14563);
xnor U16755 (N_16755,N_14377,N_14773);
xor U16756 (N_16756,N_14682,N_15473);
and U16757 (N_16757,N_15475,N_15003);
or U16758 (N_16758,N_15432,N_14916);
and U16759 (N_16759,N_15570,N_15408);
and U16760 (N_16760,N_14142,N_14445);
nand U16761 (N_16761,N_15034,N_15722);
xnor U16762 (N_16762,N_14925,N_15124);
and U16763 (N_16763,N_14693,N_14816);
and U16764 (N_16764,N_14001,N_15243);
and U16765 (N_16765,N_15812,N_14589);
xnor U16766 (N_16766,N_15972,N_15981);
nand U16767 (N_16767,N_14463,N_15211);
or U16768 (N_16768,N_14780,N_14762);
and U16769 (N_16769,N_15174,N_15978);
or U16770 (N_16770,N_15901,N_15443);
nor U16771 (N_16771,N_14815,N_14484);
and U16772 (N_16772,N_15740,N_15600);
nor U16773 (N_16773,N_14751,N_14410);
xor U16774 (N_16774,N_14255,N_15814);
nand U16775 (N_16775,N_14080,N_14298);
and U16776 (N_16776,N_14707,N_15448);
nor U16777 (N_16777,N_15583,N_15687);
nand U16778 (N_16778,N_15005,N_15366);
nor U16779 (N_16779,N_14112,N_15341);
nor U16780 (N_16780,N_14865,N_14010);
nor U16781 (N_16781,N_14364,N_14552);
or U16782 (N_16782,N_15376,N_14357);
or U16783 (N_16783,N_15490,N_14675);
nand U16784 (N_16784,N_15436,N_15755);
nor U16785 (N_16785,N_15973,N_14516);
or U16786 (N_16786,N_14018,N_15466);
or U16787 (N_16787,N_14176,N_15327);
nor U16788 (N_16788,N_14111,N_14753);
nand U16789 (N_16789,N_14412,N_14665);
and U16790 (N_16790,N_14734,N_14361);
nand U16791 (N_16791,N_15165,N_15908);
nor U16792 (N_16792,N_15764,N_15593);
or U16793 (N_16793,N_14512,N_14078);
and U16794 (N_16794,N_15861,N_15551);
nand U16795 (N_16795,N_14580,N_14102);
nor U16796 (N_16796,N_14790,N_15195);
nor U16797 (N_16797,N_14672,N_14063);
or U16798 (N_16798,N_14124,N_15449);
xnor U16799 (N_16799,N_14845,N_15383);
nand U16800 (N_16800,N_15269,N_15595);
xnor U16801 (N_16801,N_14075,N_15954);
or U16802 (N_16802,N_15859,N_15682);
nand U16803 (N_16803,N_14514,N_15895);
xor U16804 (N_16804,N_15669,N_15357);
nand U16805 (N_16805,N_14810,N_15460);
nor U16806 (N_16806,N_14375,N_14187);
nand U16807 (N_16807,N_14002,N_15825);
and U16808 (N_16808,N_15678,N_14940);
xor U16809 (N_16809,N_14358,N_15182);
xor U16810 (N_16810,N_15510,N_15772);
or U16811 (N_16811,N_14622,N_15508);
xnor U16812 (N_16812,N_15039,N_15199);
or U16813 (N_16813,N_14688,N_15598);
nand U16814 (N_16814,N_14472,N_14059);
and U16815 (N_16815,N_14097,N_14348);
or U16816 (N_16816,N_14192,N_15561);
nor U16817 (N_16817,N_14720,N_15940);
nor U16818 (N_16818,N_14777,N_15996);
xnor U16819 (N_16819,N_14891,N_14209);
xor U16820 (N_16820,N_14528,N_14678);
or U16821 (N_16821,N_15986,N_14692);
nor U16822 (N_16822,N_15444,N_15150);
or U16823 (N_16823,N_15459,N_15902);
xor U16824 (N_16824,N_14043,N_14646);
and U16825 (N_16825,N_15767,N_15389);
nor U16826 (N_16826,N_14874,N_14224);
nand U16827 (N_16827,N_14818,N_14533);
nor U16828 (N_16828,N_15387,N_14892);
nand U16829 (N_16829,N_14263,N_14855);
or U16830 (N_16830,N_15522,N_15251);
xor U16831 (N_16831,N_15943,N_14337);
nand U16832 (N_16832,N_14424,N_14805);
and U16833 (N_16833,N_15282,N_15699);
nor U16834 (N_16834,N_15434,N_14099);
or U16835 (N_16835,N_14197,N_15144);
or U16836 (N_16836,N_15193,N_15928);
nor U16837 (N_16837,N_14129,N_14835);
nand U16838 (N_16838,N_15082,N_15314);
nor U16839 (N_16839,N_15320,N_14677);
nor U16840 (N_16840,N_14967,N_14823);
and U16841 (N_16841,N_15037,N_14408);
or U16842 (N_16842,N_14147,N_15858);
and U16843 (N_16843,N_15488,N_15137);
xnor U16844 (N_16844,N_14871,N_14996);
nand U16845 (N_16845,N_15499,N_14586);
nand U16846 (N_16846,N_15491,N_15587);
nand U16847 (N_16847,N_14220,N_14107);
nor U16848 (N_16848,N_15433,N_15168);
nor U16849 (N_16849,N_15318,N_14237);
and U16850 (N_16850,N_14593,N_15882);
or U16851 (N_16851,N_14279,N_15084);
nor U16852 (N_16852,N_15360,N_15230);
or U16853 (N_16853,N_14006,N_14190);
nor U16854 (N_16854,N_15988,N_15774);
nor U16855 (N_16855,N_15907,N_14848);
and U16856 (N_16856,N_14507,N_14182);
nor U16857 (N_16857,N_14406,N_15864);
nand U16858 (N_16858,N_14303,N_15800);
nor U16859 (N_16859,N_14393,N_15435);
nor U16860 (N_16860,N_15078,N_14200);
xnor U16861 (N_16861,N_14603,N_14583);
nor U16862 (N_16862,N_14280,N_14636);
nand U16863 (N_16863,N_15294,N_15929);
or U16864 (N_16864,N_14706,N_14994);
or U16865 (N_16865,N_15936,N_14936);
or U16866 (N_16866,N_14741,N_15925);
or U16867 (N_16867,N_14998,N_15803);
xor U16868 (N_16868,N_14830,N_14800);
xnor U16869 (N_16869,N_15809,N_15995);
nand U16870 (N_16870,N_15599,N_15349);
or U16871 (N_16871,N_15125,N_15728);
nand U16872 (N_16872,N_15686,N_15249);
nand U16873 (N_16873,N_14679,N_14701);
and U16874 (N_16874,N_15921,N_14798);
and U16875 (N_16875,N_15751,N_14919);
xor U16876 (N_16876,N_15631,N_14602);
or U16877 (N_16877,N_14109,N_15263);
and U16878 (N_16878,N_15562,N_14838);
or U16879 (N_16879,N_14409,N_15841);
nor U16880 (N_16880,N_14350,N_15223);
and U16881 (N_16881,N_14403,N_14050);
xnor U16882 (N_16882,N_14286,N_15467);
nor U16883 (N_16883,N_15527,N_14397);
nor U16884 (N_16884,N_15810,N_15944);
or U16885 (N_16885,N_14259,N_15285);
and U16886 (N_16886,N_15298,N_14131);
and U16887 (N_16887,N_15181,N_14407);
or U16888 (N_16888,N_14134,N_15894);
nand U16889 (N_16889,N_14148,N_15262);
xor U16890 (N_16890,N_14625,N_14997);
xor U16891 (N_16891,N_14881,N_15038);
nor U16892 (N_16892,N_15725,N_14511);
or U16893 (N_16893,N_15775,N_14282);
and U16894 (N_16894,N_15053,N_14113);
nand U16895 (N_16895,N_14214,N_14391);
nand U16896 (N_16896,N_15129,N_14352);
and U16897 (N_16897,N_14787,N_15160);
nor U16898 (N_16898,N_14774,N_14271);
nor U16899 (N_16899,N_15579,N_15420);
nor U16900 (N_16900,N_14870,N_15535);
nor U16901 (N_16901,N_14106,N_15164);
or U16902 (N_16902,N_14973,N_15905);
or U16903 (N_16903,N_15250,N_14882);
nor U16904 (N_16904,N_14126,N_15817);
xnor U16905 (N_16905,N_14788,N_14387);
or U16906 (N_16906,N_15495,N_14673);
nand U16907 (N_16907,N_15723,N_15489);
and U16908 (N_16908,N_15997,N_14223);
and U16909 (N_16909,N_15316,N_14047);
and U16910 (N_16910,N_15422,N_15654);
or U16911 (N_16911,N_14493,N_15009);
or U16912 (N_16912,N_15779,N_15222);
nand U16913 (N_16913,N_15904,N_15102);
nand U16914 (N_16914,N_14772,N_14384);
nor U16915 (N_16915,N_15845,N_14779);
or U16916 (N_16916,N_14897,N_15410);
nor U16917 (N_16917,N_15214,N_14347);
xor U16918 (N_16918,N_14630,N_15698);
xnor U16919 (N_16919,N_14172,N_15086);
or U16920 (N_16920,N_14328,N_15497);
or U16921 (N_16921,N_14011,N_14803);
nand U16922 (N_16922,N_14086,N_15047);
and U16923 (N_16923,N_14221,N_15569);
nor U16924 (N_16924,N_14719,N_15128);
and U16925 (N_16925,N_14834,N_15677);
or U16926 (N_16926,N_14594,N_15171);
nand U16927 (N_16927,N_15657,N_14133);
or U16928 (N_16928,N_14257,N_15147);
nor U16929 (N_16929,N_14813,N_15221);
and U16930 (N_16930,N_15582,N_14027);
nor U16931 (N_16931,N_14980,N_15616);
nand U16932 (N_16932,N_14467,N_15192);
nor U16933 (N_16933,N_15307,N_15730);
xnor U16934 (N_16934,N_14233,N_15715);
xnor U16935 (N_16935,N_15847,N_14623);
nand U16936 (N_16936,N_15885,N_15982);
and U16937 (N_16937,N_14165,N_15167);
nor U16938 (N_16938,N_15346,N_15455);
and U16939 (N_16939,N_15596,N_15735);
xor U16940 (N_16940,N_14669,N_14074);
or U16941 (N_16941,N_15976,N_14785);
nand U16942 (N_16942,N_15602,N_15792);
and U16943 (N_16943,N_15231,N_15107);
xnor U16944 (N_16944,N_14180,N_14869);
nand U16945 (N_16945,N_14792,N_14873);
nand U16946 (N_16946,N_15391,N_15276);
nor U16947 (N_16947,N_14754,N_14240);
nand U16948 (N_16948,N_14323,N_15604);
and U16949 (N_16949,N_14888,N_15119);
nor U16950 (N_16950,N_15050,N_14588);
or U16951 (N_16951,N_14367,N_15670);
xnor U16952 (N_16952,N_14548,N_15333);
nand U16953 (N_16953,N_14079,N_15838);
or U16954 (N_16954,N_14987,N_14170);
nor U16955 (N_16955,N_14889,N_15265);
and U16956 (N_16956,N_15088,N_14349);
or U16957 (N_16957,N_14687,N_14185);
xor U16958 (N_16958,N_14523,N_15062);
nand U16959 (N_16959,N_15407,N_14173);
xnor U16960 (N_16960,N_14345,N_14231);
and U16961 (N_16961,N_15478,N_14297);
or U16962 (N_16962,N_15268,N_14035);
and U16963 (N_16963,N_14166,N_14149);
and U16964 (N_16964,N_15123,N_14483);
and U16965 (N_16965,N_15556,N_15492);
nand U16966 (N_16966,N_14819,N_14284);
nand U16967 (N_16967,N_15235,N_14141);
and U16968 (N_16968,N_15913,N_14388);
nand U16969 (N_16969,N_15934,N_15016);
xor U16970 (N_16970,N_15278,N_15446);
or U16971 (N_16971,N_14356,N_15700);
xor U16972 (N_16972,N_15134,N_14379);
and U16973 (N_16973,N_14635,N_14894);
or U16974 (N_16974,N_15043,N_14415);
nand U16975 (N_16975,N_15070,N_14252);
nor U16976 (N_16976,N_15721,N_14524);
or U16977 (N_16977,N_14152,N_15951);
or U16978 (N_16978,N_15031,N_14437);
xnor U16979 (N_16979,N_15854,N_15418);
nand U16980 (N_16980,N_14858,N_14105);
xor U16981 (N_16981,N_14628,N_15238);
nand U16982 (N_16982,N_15836,N_15234);
xor U16983 (N_16983,N_14781,N_14459);
and U16984 (N_16984,N_15691,N_14159);
or U16985 (N_16985,N_14654,N_14702);
nand U16986 (N_16986,N_15695,N_15505);
nor U16987 (N_16987,N_15514,N_14627);
or U16988 (N_16988,N_14854,N_14812);
and U16989 (N_16989,N_15400,N_14489);
or U16990 (N_16990,N_15793,N_15259);
and U16991 (N_16991,N_14023,N_14072);
nand U16992 (N_16992,N_14292,N_14184);
xor U16993 (N_16993,N_15382,N_15289);
xor U16994 (N_16994,N_14555,N_15036);
nor U16995 (N_16995,N_15261,N_15283);
or U16996 (N_16996,N_15567,N_15364);
nand U16997 (N_16997,N_15862,N_14418);
and U16998 (N_16998,N_14127,N_14227);
nor U16999 (N_16999,N_14250,N_14624);
xnor U17000 (N_17000,N_14633,N_14298);
and U17001 (N_17001,N_15226,N_14717);
and U17002 (N_17002,N_15439,N_14578);
nand U17003 (N_17003,N_15010,N_15252);
nor U17004 (N_17004,N_14154,N_15576);
nand U17005 (N_17005,N_15771,N_15129);
nor U17006 (N_17006,N_14156,N_15237);
and U17007 (N_17007,N_14202,N_15070);
nor U17008 (N_17008,N_15364,N_15808);
or U17009 (N_17009,N_15895,N_14498);
or U17010 (N_17010,N_14938,N_14216);
or U17011 (N_17011,N_15211,N_14641);
nor U17012 (N_17012,N_15229,N_15094);
or U17013 (N_17013,N_15918,N_14969);
nand U17014 (N_17014,N_14848,N_15010);
nor U17015 (N_17015,N_14029,N_14073);
nand U17016 (N_17016,N_14628,N_15836);
or U17017 (N_17017,N_14154,N_15477);
and U17018 (N_17018,N_15699,N_14107);
nand U17019 (N_17019,N_15906,N_14416);
or U17020 (N_17020,N_15278,N_14705);
nor U17021 (N_17021,N_15973,N_14806);
xnor U17022 (N_17022,N_14828,N_14587);
and U17023 (N_17023,N_14035,N_15561);
or U17024 (N_17024,N_15567,N_15379);
and U17025 (N_17025,N_15133,N_15946);
and U17026 (N_17026,N_15502,N_14618);
xor U17027 (N_17027,N_15424,N_15062);
and U17028 (N_17028,N_15208,N_15352);
xnor U17029 (N_17029,N_14448,N_15511);
nand U17030 (N_17030,N_15731,N_14148);
nand U17031 (N_17031,N_15889,N_14492);
and U17032 (N_17032,N_14380,N_15905);
xor U17033 (N_17033,N_15693,N_15671);
nor U17034 (N_17034,N_14414,N_15903);
or U17035 (N_17035,N_14849,N_14794);
or U17036 (N_17036,N_14496,N_15220);
nand U17037 (N_17037,N_14538,N_15442);
and U17038 (N_17038,N_14070,N_14922);
xnor U17039 (N_17039,N_15417,N_15025);
nand U17040 (N_17040,N_14052,N_14308);
nand U17041 (N_17041,N_14583,N_15195);
nand U17042 (N_17042,N_14428,N_15489);
nor U17043 (N_17043,N_14369,N_15637);
and U17044 (N_17044,N_14449,N_15113);
xnor U17045 (N_17045,N_14117,N_14481);
nor U17046 (N_17046,N_15735,N_15876);
xor U17047 (N_17047,N_14939,N_15990);
nor U17048 (N_17048,N_14299,N_15165);
and U17049 (N_17049,N_14711,N_15293);
nor U17050 (N_17050,N_15777,N_14899);
nor U17051 (N_17051,N_15379,N_15508);
nor U17052 (N_17052,N_15006,N_15355);
or U17053 (N_17053,N_15006,N_15191);
or U17054 (N_17054,N_14398,N_14570);
and U17055 (N_17055,N_14441,N_15064);
and U17056 (N_17056,N_15354,N_15985);
xnor U17057 (N_17057,N_15693,N_15889);
and U17058 (N_17058,N_14210,N_14822);
nor U17059 (N_17059,N_14999,N_14716);
and U17060 (N_17060,N_15874,N_14007);
or U17061 (N_17061,N_14247,N_14480);
nand U17062 (N_17062,N_15761,N_14853);
and U17063 (N_17063,N_14523,N_14940);
xnor U17064 (N_17064,N_15243,N_15259);
nor U17065 (N_17065,N_14006,N_15789);
or U17066 (N_17066,N_14352,N_14445);
or U17067 (N_17067,N_15820,N_14592);
nor U17068 (N_17068,N_14037,N_15067);
xnor U17069 (N_17069,N_15620,N_14692);
nor U17070 (N_17070,N_14288,N_15125);
or U17071 (N_17071,N_14107,N_14274);
xor U17072 (N_17072,N_14912,N_14664);
nor U17073 (N_17073,N_15360,N_15341);
nand U17074 (N_17074,N_14446,N_14807);
xor U17075 (N_17075,N_14597,N_15541);
xnor U17076 (N_17076,N_15210,N_14597);
and U17077 (N_17077,N_14803,N_14652);
nand U17078 (N_17078,N_15096,N_14389);
and U17079 (N_17079,N_15441,N_14859);
and U17080 (N_17080,N_15118,N_14920);
xor U17081 (N_17081,N_15517,N_15267);
nor U17082 (N_17082,N_15619,N_15840);
xor U17083 (N_17083,N_15249,N_14592);
nand U17084 (N_17084,N_14437,N_14118);
or U17085 (N_17085,N_14434,N_14013);
or U17086 (N_17086,N_15426,N_14053);
nand U17087 (N_17087,N_15243,N_15393);
or U17088 (N_17088,N_15206,N_15242);
and U17089 (N_17089,N_14773,N_14928);
nor U17090 (N_17090,N_14875,N_15881);
nor U17091 (N_17091,N_15294,N_14851);
nor U17092 (N_17092,N_15614,N_14295);
xor U17093 (N_17093,N_15862,N_14941);
nor U17094 (N_17094,N_14265,N_14980);
or U17095 (N_17095,N_14432,N_15453);
and U17096 (N_17096,N_14823,N_15440);
nor U17097 (N_17097,N_15015,N_15320);
and U17098 (N_17098,N_15158,N_15435);
xnor U17099 (N_17099,N_14366,N_15448);
nand U17100 (N_17100,N_14778,N_14271);
or U17101 (N_17101,N_14554,N_14562);
or U17102 (N_17102,N_14836,N_15708);
or U17103 (N_17103,N_14434,N_15830);
or U17104 (N_17104,N_15831,N_15075);
and U17105 (N_17105,N_15795,N_15546);
nor U17106 (N_17106,N_14460,N_14743);
nor U17107 (N_17107,N_15305,N_14649);
nor U17108 (N_17108,N_14612,N_14196);
or U17109 (N_17109,N_15052,N_15053);
and U17110 (N_17110,N_15688,N_14756);
or U17111 (N_17111,N_14146,N_15794);
nor U17112 (N_17112,N_14545,N_15342);
or U17113 (N_17113,N_15006,N_14575);
xor U17114 (N_17114,N_14148,N_14240);
and U17115 (N_17115,N_14490,N_14363);
and U17116 (N_17116,N_15598,N_14411);
nor U17117 (N_17117,N_15360,N_14153);
xnor U17118 (N_17118,N_14253,N_15849);
and U17119 (N_17119,N_15394,N_15262);
or U17120 (N_17120,N_14502,N_14353);
and U17121 (N_17121,N_14835,N_15035);
nor U17122 (N_17122,N_14970,N_15329);
xnor U17123 (N_17123,N_15090,N_14881);
or U17124 (N_17124,N_14658,N_14417);
xor U17125 (N_17125,N_14895,N_14323);
xor U17126 (N_17126,N_14857,N_14541);
or U17127 (N_17127,N_14056,N_14054);
or U17128 (N_17128,N_15529,N_14064);
nor U17129 (N_17129,N_15121,N_15374);
xor U17130 (N_17130,N_15826,N_15871);
nand U17131 (N_17131,N_15890,N_15412);
xnor U17132 (N_17132,N_14747,N_15608);
or U17133 (N_17133,N_15829,N_14204);
nor U17134 (N_17134,N_15452,N_15942);
xor U17135 (N_17135,N_15450,N_15831);
nor U17136 (N_17136,N_14349,N_14975);
nor U17137 (N_17137,N_15380,N_14048);
nor U17138 (N_17138,N_14865,N_15008);
nand U17139 (N_17139,N_15667,N_15882);
or U17140 (N_17140,N_14088,N_14650);
nor U17141 (N_17141,N_15804,N_14880);
nand U17142 (N_17142,N_15816,N_15788);
nor U17143 (N_17143,N_14570,N_15023);
nor U17144 (N_17144,N_15323,N_15582);
and U17145 (N_17145,N_15721,N_14817);
and U17146 (N_17146,N_14314,N_15423);
or U17147 (N_17147,N_14164,N_15357);
nand U17148 (N_17148,N_15729,N_15880);
and U17149 (N_17149,N_15507,N_14347);
and U17150 (N_17150,N_15575,N_14859);
xnor U17151 (N_17151,N_15731,N_14650);
xor U17152 (N_17152,N_15190,N_15291);
or U17153 (N_17153,N_14564,N_15532);
nor U17154 (N_17154,N_14987,N_15947);
nand U17155 (N_17155,N_15072,N_14845);
nand U17156 (N_17156,N_15206,N_14654);
xor U17157 (N_17157,N_15117,N_14969);
nor U17158 (N_17158,N_15023,N_14569);
and U17159 (N_17159,N_15990,N_15705);
xnor U17160 (N_17160,N_14198,N_15585);
or U17161 (N_17161,N_14552,N_14762);
and U17162 (N_17162,N_15297,N_15851);
nor U17163 (N_17163,N_15468,N_15962);
and U17164 (N_17164,N_14966,N_15946);
xnor U17165 (N_17165,N_15455,N_15583);
xor U17166 (N_17166,N_15343,N_14668);
nor U17167 (N_17167,N_15692,N_14723);
and U17168 (N_17168,N_14139,N_15985);
or U17169 (N_17169,N_15461,N_14686);
or U17170 (N_17170,N_14261,N_14024);
or U17171 (N_17171,N_15960,N_15716);
and U17172 (N_17172,N_15971,N_14864);
nand U17173 (N_17173,N_14904,N_15010);
xor U17174 (N_17174,N_15536,N_14224);
and U17175 (N_17175,N_15917,N_15893);
xnor U17176 (N_17176,N_14901,N_15646);
or U17177 (N_17177,N_14057,N_14818);
and U17178 (N_17178,N_14834,N_14406);
or U17179 (N_17179,N_15571,N_15055);
or U17180 (N_17180,N_14779,N_15905);
nor U17181 (N_17181,N_14431,N_15995);
xor U17182 (N_17182,N_14979,N_14308);
nor U17183 (N_17183,N_14112,N_15087);
nor U17184 (N_17184,N_15538,N_15807);
xnor U17185 (N_17185,N_15630,N_15716);
xnor U17186 (N_17186,N_15119,N_15434);
nand U17187 (N_17187,N_14831,N_15822);
or U17188 (N_17188,N_14738,N_14079);
or U17189 (N_17189,N_15562,N_15360);
nor U17190 (N_17190,N_15898,N_15846);
and U17191 (N_17191,N_15819,N_15329);
and U17192 (N_17192,N_15205,N_15306);
nor U17193 (N_17193,N_15475,N_14876);
and U17194 (N_17194,N_14530,N_15056);
nor U17195 (N_17195,N_14700,N_15270);
nand U17196 (N_17196,N_14886,N_14767);
xor U17197 (N_17197,N_15340,N_14132);
xor U17198 (N_17198,N_14466,N_15885);
or U17199 (N_17199,N_15510,N_15384);
nand U17200 (N_17200,N_14513,N_14523);
xnor U17201 (N_17201,N_15215,N_14375);
nand U17202 (N_17202,N_14515,N_15201);
nor U17203 (N_17203,N_15782,N_14771);
or U17204 (N_17204,N_15761,N_14111);
nand U17205 (N_17205,N_14998,N_15842);
or U17206 (N_17206,N_14126,N_15568);
nand U17207 (N_17207,N_14350,N_14404);
nor U17208 (N_17208,N_14257,N_14541);
or U17209 (N_17209,N_14975,N_14016);
or U17210 (N_17210,N_15866,N_15190);
xor U17211 (N_17211,N_14076,N_15147);
nor U17212 (N_17212,N_14349,N_14532);
or U17213 (N_17213,N_14376,N_14278);
and U17214 (N_17214,N_15469,N_15917);
nand U17215 (N_17215,N_14170,N_15759);
nand U17216 (N_17216,N_15968,N_14264);
nand U17217 (N_17217,N_15261,N_14073);
and U17218 (N_17218,N_14124,N_14853);
nand U17219 (N_17219,N_15872,N_14156);
xnor U17220 (N_17220,N_15812,N_14966);
nand U17221 (N_17221,N_15061,N_15849);
or U17222 (N_17222,N_14126,N_15518);
nor U17223 (N_17223,N_15267,N_15374);
and U17224 (N_17224,N_14665,N_15062);
xnor U17225 (N_17225,N_14845,N_15165);
and U17226 (N_17226,N_15487,N_14868);
nor U17227 (N_17227,N_14307,N_15975);
or U17228 (N_17228,N_14379,N_15868);
and U17229 (N_17229,N_15851,N_15445);
nor U17230 (N_17230,N_14315,N_14817);
nand U17231 (N_17231,N_14806,N_15382);
and U17232 (N_17232,N_15779,N_15730);
nor U17233 (N_17233,N_15041,N_15015);
and U17234 (N_17234,N_14548,N_15326);
xor U17235 (N_17235,N_14489,N_15545);
nand U17236 (N_17236,N_14151,N_15079);
and U17237 (N_17237,N_15476,N_14827);
and U17238 (N_17238,N_15863,N_14744);
nor U17239 (N_17239,N_15143,N_14043);
nand U17240 (N_17240,N_14179,N_15069);
or U17241 (N_17241,N_14372,N_14448);
nor U17242 (N_17242,N_15956,N_15419);
or U17243 (N_17243,N_15229,N_15446);
nor U17244 (N_17244,N_15487,N_15613);
nor U17245 (N_17245,N_15893,N_15630);
or U17246 (N_17246,N_15451,N_14076);
nor U17247 (N_17247,N_14812,N_15203);
or U17248 (N_17248,N_14204,N_15555);
nand U17249 (N_17249,N_15189,N_15617);
nand U17250 (N_17250,N_14283,N_14800);
nand U17251 (N_17251,N_15519,N_14042);
xnor U17252 (N_17252,N_14635,N_15490);
or U17253 (N_17253,N_14430,N_15356);
nor U17254 (N_17254,N_14837,N_14161);
and U17255 (N_17255,N_15765,N_15684);
and U17256 (N_17256,N_15694,N_15746);
and U17257 (N_17257,N_14450,N_15260);
nand U17258 (N_17258,N_15305,N_14935);
or U17259 (N_17259,N_15227,N_15159);
nor U17260 (N_17260,N_15740,N_15874);
nand U17261 (N_17261,N_14465,N_14189);
and U17262 (N_17262,N_14239,N_15766);
nand U17263 (N_17263,N_14539,N_15895);
or U17264 (N_17264,N_15711,N_14156);
nor U17265 (N_17265,N_15748,N_14947);
nor U17266 (N_17266,N_14704,N_15741);
nor U17267 (N_17267,N_15656,N_15729);
or U17268 (N_17268,N_15511,N_15414);
or U17269 (N_17269,N_15859,N_15048);
and U17270 (N_17270,N_15299,N_14393);
nor U17271 (N_17271,N_15127,N_14763);
nor U17272 (N_17272,N_14922,N_14372);
nand U17273 (N_17273,N_15882,N_15521);
nor U17274 (N_17274,N_15304,N_14347);
and U17275 (N_17275,N_15706,N_14089);
xnor U17276 (N_17276,N_15177,N_14279);
nor U17277 (N_17277,N_15572,N_14987);
nand U17278 (N_17278,N_15087,N_14685);
nand U17279 (N_17279,N_15614,N_14723);
xor U17280 (N_17280,N_15710,N_15570);
nand U17281 (N_17281,N_14877,N_14774);
xnor U17282 (N_17282,N_14746,N_15773);
nand U17283 (N_17283,N_15358,N_15021);
xor U17284 (N_17284,N_15292,N_15730);
nand U17285 (N_17285,N_14139,N_15754);
nor U17286 (N_17286,N_15548,N_14266);
or U17287 (N_17287,N_15392,N_14098);
xnor U17288 (N_17288,N_14992,N_15440);
or U17289 (N_17289,N_14921,N_15085);
and U17290 (N_17290,N_14596,N_14953);
or U17291 (N_17291,N_15803,N_15006);
and U17292 (N_17292,N_14661,N_15161);
xnor U17293 (N_17293,N_15343,N_15987);
nand U17294 (N_17294,N_15191,N_14097);
or U17295 (N_17295,N_14526,N_15100);
and U17296 (N_17296,N_14250,N_15322);
xnor U17297 (N_17297,N_14416,N_15614);
nor U17298 (N_17298,N_15601,N_15674);
xnor U17299 (N_17299,N_14235,N_14096);
nor U17300 (N_17300,N_15330,N_15900);
or U17301 (N_17301,N_15349,N_14694);
nand U17302 (N_17302,N_14622,N_14532);
xor U17303 (N_17303,N_14282,N_14889);
nand U17304 (N_17304,N_14158,N_15372);
nand U17305 (N_17305,N_14977,N_15677);
or U17306 (N_17306,N_15418,N_14901);
nor U17307 (N_17307,N_14041,N_14566);
nor U17308 (N_17308,N_15241,N_14686);
and U17309 (N_17309,N_14834,N_15976);
nand U17310 (N_17310,N_14343,N_14989);
nor U17311 (N_17311,N_15369,N_14378);
nor U17312 (N_17312,N_15338,N_14311);
xor U17313 (N_17313,N_14685,N_15976);
and U17314 (N_17314,N_14216,N_15656);
xor U17315 (N_17315,N_15949,N_15206);
nand U17316 (N_17316,N_14226,N_14249);
and U17317 (N_17317,N_15329,N_14142);
xor U17318 (N_17318,N_14551,N_15537);
xor U17319 (N_17319,N_15074,N_14882);
and U17320 (N_17320,N_14559,N_15001);
xor U17321 (N_17321,N_15788,N_14663);
xor U17322 (N_17322,N_14977,N_14820);
xor U17323 (N_17323,N_15244,N_15426);
xor U17324 (N_17324,N_15685,N_15335);
or U17325 (N_17325,N_14917,N_14921);
xor U17326 (N_17326,N_15042,N_14664);
nor U17327 (N_17327,N_15040,N_15871);
and U17328 (N_17328,N_14064,N_15032);
nand U17329 (N_17329,N_15842,N_14761);
or U17330 (N_17330,N_15921,N_15515);
nand U17331 (N_17331,N_14656,N_14297);
or U17332 (N_17332,N_14368,N_15531);
xnor U17333 (N_17333,N_15501,N_14760);
or U17334 (N_17334,N_15923,N_15799);
or U17335 (N_17335,N_15324,N_15271);
nor U17336 (N_17336,N_14652,N_14313);
xnor U17337 (N_17337,N_14276,N_15677);
and U17338 (N_17338,N_14881,N_14321);
nand U17339 (N_17339,N_15974,N_14041);
nand U17340 (N_17340,N_14521,N_14819);
nor U17341 (N_17341,N_15986,N_14079);
and U17342 (N_17342,N_15014,N_15295);
and U17343 (N_17343,N_15596,N_14902);
or U17344 (N_17344,N_14326,N_14127);
or U17345 (N_17345,N_15225,N_14246);
xnor U17346 (N_17346,N_14451,N_14537);
nand U17347 (N_17347,N_15511,N_14616);
xnor U17348 (N_17348,N_14324,N_14882);
or U17349 (N_17349,N_15987,N_14056);
or U17350 (N_17350,N_14351,N_14816);
nor U17351 (N_17351,N_14522,N_15918);
nand U17352 (N_17352,N_14783,N_14770);
xnor U17353 (N_17353,N_15645,N_14555);
nor U17354 (N_17354,N_15122,N_15224);
nor U17355 (N_17355,N_14362,N_15408);
nor U17356 (N_17356,N_14976,N_15866);
or U17357 (N_17357,N_14712,N_14606);
and U17358 (N_17358,N_14170,N_15082);
or U17359 (N_17359,N_15330,N_14455);
nand U17360 (N_17360,N_14706,N_15551);
nor U17361 (N_17361,N_15688,N_14115);
and U17362 (N_17362,N_15613,N_14476);
xnor U17363 (N_17363,N_15572,N_14494);
nor U17364 (N_17364,N_14559,N_14057);
or U17365 (N_17365,N_14553,N_14204);
or U17366 (N_17366,N_14561,N_14225);
xnor U17367 (N_17367,N_14598,N_14886);
and U17368 (N_17368,N_15475,N_15978);
xnor U17369 (N_17369,N_14602,N_15795);
nor U17370 (N_17370,N_14887,N_15363);
and U17371 (N_17371,N_14534,N_14120);
xnor U17372 (N_17372,N_15274,N_15922);
or U17373 (N_17373,N_14303,N_14364);
or U17374 (N_17374,N_15060,N_14841);
nor U17375 (N_17375,N_15681,N_14264);
xnor U17376 (N_17376,N_14756,N_15111);
or U17377 (N_17377,N_14574,N_14407);
or U17378 (N_17378,N_15217,N_14175);
xnor U17379 (N_17379,N_14938,N_14456);
nor U17380 (N_17380,N_14384,N_14897);
nand U17381 (N_17381,N_14134,N_14323);
and U17382 (N_17382,N_15034,N_14442);
or U17383 (N_17383,N_14543,N_15191);
or U17384 (N_17384,N_15772,N_15836);
nand U17385 (N_17385,N_15160,N_15235);
nand U17386 (N_17386,N_14067,N_14365);
and U17387 (N_17387,N_14884,N_15871);
and U17388 (N_17388,N_14894,N_15635);
or U17389 (N_17389,N_14113,N_15066);
nand U17390 (N_17390,N_15229,N_14303);
or U17391 (N_17391,N_15917,N_14471);
xor U17392 (N_17392,N_14980,N_15157);
nand U17393 (N_17393,N_15272,N_15099);
xor U17394 (N_17394,N_14895,N_14013);
xnor U17395 (N_17395,N_14666,N_15772);
or U17396 (N_17396,N_15522,N_14414);
nand U17397 (N_17397,N_15123,N_14315);
nor U17398 (N_17398,N_15689,N_15367);
nand U17399 (N_17399,N_15957,N_14652);
or U17400 (N_17400,N_15973,N_14414);
xnor U17401 (N_17401,N_15877,N_14545);
or U17402 (N_17402,N_15950,N_14117);
and U17403 (N_17403,N_15890,N_14021);
or U17404 (N_17404,N_14262,N_15997);
and U17405 (N_17405,N_14215,N_15946);
or U17406 (N_17406,N_15199,N_14515);
nand U17407 (N_17407,N_14365,N_14971);
and U17408 (N_17408,N_14207,N_15153);
nor U17409 (N_17409,N_15185,N_14418);
nor U17410 (N_17410,N_15042,N_14192);
and U17411 (N_17411,N_14619,N_15480);
nor U17412 (N_17412,N_14655,N_14460);
nand U17413 (N_17413,N_15572,N_14018);
nand U17414 (N_17414,N_14338,N_14114);
or U17415 (N_17415,N_15776,N_15796);
and U17416 (N_17416,N_14734,N_14986);
xnor U17417 (N_17417,N_14650,N_15527);
and U17418 (N_17418,N_14461,N_15773);
or U17419 (N_17419,N_15419,N_14179);
or U17420 (N_17420,N_15981,N_15983);
nor U17421 (N_17421,N_15366,N_15746);
nor U17422 (N_17422,N_14321,N_14378);
or U17423 (N_17423,N_14801,N_15556);
or U17424 (N_17424,N_14605,N_14552);
and U17425 (N_17425,N_15298,N_14531);
or U17426 (N_17426,N_15323,N_15468);
and U17427 (N_17427,N_15720,N_15678);
and U17428 (N_17428,N_15477,N_14884);
xor U17429 (N_17429,N_14996,N_14623);
xnor U17430 (N_17430,N_14252,N_14629);
and U17431 (N_17431,N_15029,N_14290);
or U17432 (N_17432,N_15851,N_15761);
nor U17433 (N_17433,N_14085,N_14601);
and U17434 (N_17434,N_15043,N_14841);
xor U17435 (N_17435,N_14341,N_15354);
or U17436 (N_17436,N_14640,N_14206);
or U17437 (N_17437,N_15510,N_14826);
nand U17438 (N_17438,N_14624,N_15555);
nand U17439 (N_17439,N_14283,N_14130);
nand U17440 (N_17440,N_15378,N_15399);
nor U17441 (N_17441,N_15847,N_14457);
nand U17442 (N_17442,N_14491,N_15361);
nor U17443 (N_17443,N_14804,N_15039);
xnor U17444 (N_17444,N_15141,N_14437);
xnor U17445 (N_17445,N_14790,N_14772);
xor U17446 (N_17446,N_15357,N_14047);
nor U17447 (N_17447,N_14683,N_14627);
nand U17448 (N_17448,N_15819,N_14212);
and U17449 (N_17449,N_15883,N_15166);
nand U17450 (N_17450,N_14889,N_15776);
and U17451 (N_17451,N_14353,N_14067);
nand U17452 (N_17452,N_14751,N_14838);
nor U17453 (N_17453,N_15113,N_14160);
nor U17454 (N_17454,N_15312,N_14450);
and U17455 (N_17455,N_14826,N_14502);
and U17456 (N_17456,N_15109,N_14898);
xor U17457 (N_17457,N_15774,N_14116);
or U17458 (N_17458,N_14610,N_14340);
nand U17459 (N_17459,N_14264,N_14603);
or U17460 (N_17460,N_14655,N_15957);
and U17461 (N_17461,N_14763,N_14456);
xnor U17462 (N_17462,N_15036,N_14754);
xor U17463 (N_17463,N_14964,N_14672);
xnor U17464 (N_17464,N_15178,N_15676);
nor U17465 (N_17465,N_14237,N_14842);
nor U17466 (N_17466,N_14601,N_14424);
and U17467 (N_17467,N_15168,N_14116);
and U17468 (N_17468,N_15715,N_14805);
or U17469 (N_17469,N_15574,N_14873);
and U17470 (N_17470,N_15999,N_14966);
nor U17471 (N_17471,N_15716,N_14061);
and U17472 (N_17472,N_14447,N_14848);
and U17473 (N_17473,N_15717,N_14753);
nor U17474 (N_17474,N_14564,N_15735);
nor U17475 (N_17475,N_14623,N_14394);
or U17476 (N_17476,N_14192,N_15281);
nand U17477 (N_17477,N_14049,N_14977);
nand U17478 (N_17478,N_15233,N_14264);
nor U17479 (N_17479,N_14081,N_15450);
xor U17480 (N_17480,N_15898,N_14305);
nand U17481 (N_17481,N_14769,N_14802);
nand U17482 (N_17482,N_15749,N_15984);
nor U17483 (N_17483,N_15690,N_14328);
xnor U17484 (N_17484,N_14157,N_14540);
nor U17485 (N_17485,N_14159,N_14304);
nand U17486 (N_17486,N_14003,N_14801);
or U17487 (N_17487,N_14493,N_15483);
or U17488 (N_17488,N_15394,N_15922);
nand U17489 (N_17489,N_15351,N_15830);
and U17490 (N_17490,N_15113,N_14146);
xnor U17491 (N_17491,N_14119,N_15132);
xor U17492 (N_17492,N_15494,N_15844);
or U17493 (N_17493,N_15867,N_15933);
nand U17494 (N_17494,N_15227,N_14269);
nand U17495 (N_17495,N_14334,N_14927);
nor U17496 (N_17496,N_15550,N_15876);
nand U17497 (N_17497,N_14351,N_14824);
and U17498 (N_17498,N_15517,N_14895);
nor U17499 (N_17499,N_14662,N_15243);
xor U17500 (N_17500,N_15220,N_14731);
nand U17501 (N_17501,N_14767,N_15546);
nand U17502 (N_17502,N_14166,N_15560);
and U17503 (N_17503,N_14657,N_14669);
or U17504 (N_17504,N_14080,N_14650);
and U17505 (N_17505,N_14409,N_14420);
nor U17506 (N_17506,N_15819,N_15663);
and U17507 (N_17507,N_14263,N_14271);
and U17508 (N_17508,N_15275,N_15425);
nor U17509 (N_17509,N_14680,N_15793);
or U17510 (N_17510,N_15260,N_15673);
xor U17511 (N_17511,N_14605,N_15683);
and U17512 (N_17512,N_14357,N_15505);
or U17513 (N_17513,N_15601,N_14904);
or U17514 (N_17514,N_15442,N_15294);
xnor U17515 (N_17515,N_15755,N_14058);
nor U17516 (N_17516,N_15765,N_14908);
nor U17517 (N_17517,N_15228,N_15218);
or U17518 (N_17518,N_15369,N_15883);
or U17519 (N_17519,N_15131,N_14842);
and U17520 (N_17520,N_15534,N_14471);
xor U17521 (N_17521,N_14667,N_14817);
and U17522 (N_17522,N_14328,N_14363);
and U17523 (N_17523,N_15324,N_15756);
xor U17524 (N_17524,N_14076,N_14301);
xnor U17525 (N_17525,N_14157,N_14739);
and U17526 (N_17526,N_15187,N_15081);
or U17527 (N_17527,N_14336,N_14619);
or U17528 (N_17528,N_14753,N_14452);
nand U17529 (N_17529,N_15144,N_14987);
xor U17530 (N_17530,N_15851,N_15867);
and U17531 (N_17531,N_14612,N_14976);
or U17532 (N_17532,N_14960,N_14678);
nor U17533 (N_17533,N_14175,N_14794);
and U17534 (N_17534,N_14982,N_14108);
or U17535 (N_17535,N_15657,N_15079);
nand U17536 (N_17536,N_14470,N_15626);
nand U17537 (N_17537,N_15205,N_14052);
and U17538 (N_17538,N_14189,N_15043);
and U17539 (N_17539,N_14231,N_14762);
nand U17540 (N_17540,N_14001,N_15343);
xor U17541 (N_17541,N_14244,N_15866);
and U17542 (N_17542,N_14895,N_14827);
xor U17543 (N_17543,N_14174,N_14413);
nor U17544 (N_17544,N_15157,N_15387);
nand U17545 (N_17545,N_14478,N_14642);
or U17546 (N_17546,N_14778,N_15394);
or U17547 (N_17547,N_14933,N_14328);
xor U17548 (N_17548,N_14430,N_14244);
xor U17549 (N_17549,N_15278,N_14138);
nor U17550 (N_17550,N_14562,N_15964);
and U17551 (N_17551,N_15981,N_15143);
nand U17552 (N_17552,N_14993,N_14352);
and U17553 (N_17553,N_14505,N_14684);
xnor U17554 (N_17554,N_15791,N_14062);
and U17555 (N_17555,N_14712,N_15515);
or U17556 (N_17556,N_15347,N_14635);
or U17557 (N_17557,N_14301,N_15231);
or U17558 (N_17558,N_14922,N_15535);
and U17559 (N_17559,N_15527,N_14520);
nand U17560 (N_17560,N_14282,N_14965);
and U17561 (N_17561,N_14637,N_15433);
xor U17562 (N_17562,N_14917,N_15283);
or U17563 (N_17563,N_15549,N_15792);
and U17564 (N_17564,N_14125,N_15884);
or U17565 (N_17565,N_15640,N_14961);
and U17566 (N_17566,N_14761,N_14654);
or U17567 (N_17567,N_14007,N_15131);
or U17568 (N_17568,N_15120,N_14419);
nor U17569 (N_17569,N_15669,N_14084);
and U17570 (N_17570,N_14503,N_15234);
xor U17571 (N_17571,N_14429,N_14081);
nand U17572 (N_17572,N_15574,N_15719);
nand U17573 (N_17573,N_15422,N_15306);
nor U17574 (N_17574,N_15950,N_14271);
and U17575 (N_17575,N_15691,N_14125);
nand U17576 (N_17576,N_14705,N_15953);
xnor U17577 (N_17577,N_14691,N_14726);
and U17578 (N_17578,N_15660,N_15108);
and U17579 (N_17579,N_14415,N_15177);
or U17580 (N_17580,N_14986,N_14382);
nand U17581 (N_17581,N_15127,N_15379);
nor U17582 (N_17582,N_15139,N_15817);
nor U17583 (N_17583,N_15841,N_14740);
and U17584 (N_17584,N_14369,N_14725);
and U17585 (N_17585,N_15154,N_14186);
xnor U17586 (N_17586,N_14336,N_15923);
or U17587 (N_17587,N_14293,N_14916);
xor U17588 (N_17588,N_14356,N_15010);
nand U17589 (N_17589,N_15140,N_14242);
or U17590 (N_17590,N_14712,N_15945);
nor U17591 (N_17591,N_14714,N_14640);
or U17592 (N_17592,N_15206,N_14167);
nor U17593 (N_17593,N_14673,N_15015);
nor U17594 (N_17594,N_14337,N_15973);
xor U17595 (N_17595,N_15768,N_15414);
nand U17596 (N_17596,N_14743,N_15545);
and U17597 (N_17597,N_15357,N_14753);
nor U17598 (N_17598,N_14839,N_15899);
and U17599 (N_17599,N_15367,N_15416);
or U17600 (N_17600,N_14207,N_15888);
or U17601 (N_17601,N_15590,N_15016);
nor U17602 (N_17602,N_14522,N_15409);
and U17603 (N_17603,N_14639,N_15787);
and U17604 (N_17604,N_15564,N_14691);
and U17605 (N_17605,N_14856,N_15240);
or U17606 (N_17606,N_14727,N_14299);
nor U17607 (N_17607,N_15806,N_15847);
xnor U17608 (N_17608,N_14721,N_14260);
nand U17609 (N_17609,N_14352,N_15103);
nand U17610 (N_17610,N_14047,N_14101);
xor U17611 (N_17611,N_14897,N_14406);
xnor U17612 (N_17612,N_14496,N_14342);
nor U17613 (N_17613,N_14902,N_14377);
nor U17614 (N_17614,N_14492,N_15694);
or U17615 (N_17615,N_15087,N_14786);
or U17616 (N_17616,N_15563,N_14093);
xor U17617 (N_17617,N_15861,N_15830);
xnor U17618 (N_17618,N_14446,N_14930);
xor U17619 (N_17619,N_15094,N_15388);
and U17620 (N_17620,N_14622,N_14507);
nor U17621 (N_17621,N_15520,N_15985);
nand U17622 (N_17622,N_15538,N_15655);
and U17623 (N_17623,N_15544,N_15792);
or U17624 (N_17624,N_14613,N_14206);
nor U17625 (N_17625,N_15441,N_15220);
xnor U17626 (N_17626,N_14511,N_15201);
and U17627 (N_17627,N_14889,N_15029);
xnor U17628 (N_17628,N_15368,N_14758);
xor U17629 (N_17629,N_14325,N_15911);
or U17630 (N_17630,N_15794,N_15487);
or U17631 (N_17631,N_14975,N_14672);
and U17632 (N_17632,N_15594,N_14307);
or U17633 (N_17633,N_15637,N_14020);
xor U17634 (N_17634,N_14678,N_14299);
and U17635 (N_17635,N_14567,N_15466);
xor U17636 (N_17636,N_14283,N_14471);
and U17637 (N_17637,N_15189,N_14117);
and U17638 (N_17638,N_14371,N_14997);
nor U17639 (N_17639,N_15389,N_15012);
nand U17640 (N_17640,N_15396,N_15774);
nor U17641 (N_17641,N_14346,N_14436);
and U17642 (N_17642,N_15922,N_15122);
and U17643 (N_17643,N_14194,N_15934);
and U17644 (N_17644,N_15184,N_15464);
xor U17645 (N_17645,N_14764,N_15138);
nor U17646 (N_17646,N_15873,N_15493);
nor U17647 (N_17647,N_14817,N_14636);
or U17648 (N_17648,N_15662,N_14237);
or U17649 (N_17649,N_15836,N_14530);
xor U17650 (N_17650,N_14014,N_15903);
nand U17651 (N_17651,N_15485,N_14107);
xnor U17652 (N_17652,N_15497,N_14607);
xnor U17653 (N_17653,N_15398,N_14784);
nand U17654 (N_17654,N_15365,N_14588);
xor U17655 (N_17655,N_15698,N_15381);
nor U17656 (N_17656,N_14500,N_15703);
and U17657 (N_17657,N_15136,N_15880);
and U17658 (N_17658,N_15140,N_15394);
and U17659 (N_17659,N_14145,N_15045);
xnor U17660 (N_17660,N_14092,N_14168);
nand U17661 (N_17661,N_14770,N_15454);
or U17662 (N_17662,N_15328,N_15076);
xnor U17663 (N_17663,N_14328,N_14440);
xor U17664 (N_17664,N_15784,N_14562);
or U17665 (N_17665,N_15870,N_14659);
nor U17666 (N_17666,N_14529,N_14562);
or U17667 (N_17667,N_15563,N_15116);
nor U17668 (N_17668,N_14765,N_14468);
and U17669 (N_17669,N_15899,N_15383);
nand U17670 (N_17670,N_14689,N_14869);
nor U17671 (N_17671,N_15762,N_14087);
and U17672 (N_17672,N_15570,N_14386);
nor U17673 (N_17673,N_14204,N_15797);
or U17674 (N_17674,N_15183,N_14554);
or U17675 (N_17675,N_15206,N_15812);
nor U17676 (N_17676,N_14702,N_14103);
nand U17677 (N_17677,N_14800,N_15691);
xnor U17678 (N_17678,N_15634,N_15314);
and U17679 (N_17679,N_14383,N_14632);
xor U17680 (N_17680,N_15949,N_14589);
nand U17681 (N_17681,N_14719,N_15934);
and U17682 (N_17682,N_14425,N_14083);
nand U17683 (N_17683,N_14328,N_14169);
or U17684 (N_17684,N_15455,N_14103);
xor U17685 (N_17685,N_15677,N_15684);
or U17686 (N_17686,N_14443,N_15289);
xor U17687 (N_17687,N_15315,N_14927);
xor U17688 (N_17688,N_15653,N_15289);
nor U17689 (N_17689,N_15145,N_14169);
nor U17690 (N_17690,N_14430,N_14673);
xor U17691 (N_17691,N_15872,N_14745);
xor U17692 (N_17692,N_15064,N_14471);
and U17693 (N_17693,N_15962,N_14799);
xor U17694 (N_17694,N_14211,N_15178);
and U17695 (N_17695,N_15506,N_14320);
or U17696 (N_17696,N_14659,N_15470);
nor U17697 (N_17697,N_15122,N_15827);
xor U17698 (N_17698,N_14564,N_15867);
and U17699 (N_17699,N_15989,N_14570);
or U17700 (N_17700,N_15972,N_14263);
nand U17701 (N_17701,N_14837,N_15708);
xor U17702 (N_17702,N_15439,N_14724);
or U17703 (N_17703,N_15115,N_15999);
nand U17704 (N_17704,N_15027,N_14565);
nor U17705 (N_17705,N_15111,N_14350);
or U17706 (N_17706,N_14961,N_14372);
or U17707 (N_17707,N_15584,N_15873);
and U17708 (N_17708,N_15141,N_14155);
or U17709 (N_17709,N_15668,N_14109);
xor U17710 (N_17710,N_15346,N_15082);
and U17711 (N_17711,N_15967,N_14937);
and U17712 (N_17712,N_15368,N_14100);
nor U17713 (N_17713,N_14866,N_14997);
xnor U17714 (N_17714,N_14388,N_15631);
nor U17715 (N_17715,N_14178,N_15659);
xnor U17716 (N_17716,N_14156,N_15774);
and U17717 (N_17717,N_14348,N_14614);
xnor U17718 (N_17718,N_15324,N_15143);
xnor U17719 (N_17719,N_14422,N_15237);
nor U17720 (N_17720,N_15205,N_14992);
nor U17721 (N_17721,N_15397,N_14039);
xnor U17722 (N_17722,N_15605,N_15220);
and U17723 (N_17723,N_15690,N_14644);
or U17724 (N_17724,N_15032,N_15002);
or U17725 (N_17725,N_14882,N_14701);
nand U17726 (N_17726,N_14726,N_14543);
nand U17727 (N_17727,N_15805,N_14296);
and U17728 (N_17728,N_14467,N_14081);
nand U17729 (N_17729,N_15800,N_14882);
xor U17730 (N_17730,N_15669,N_14729);
xnor U17731 (N_17731,N_15396,N_15406);
and U17732 (N_17732,N_14554,N_15439);
or U17733 (N_17733,N_14508,N_14021);
nor U17734 (N_17734,N_15123,N_15337);
and U17735 (N_17735,N_14419,N_15490);
nor U17736 (N_17736,N_14794,N_15891);
and U17737 (N_17737,N_14397,N_14267);
nand U17738 (N_17738,N_14450,N_15271);
nor U17739 (N_17739,N_14748,N_15104);
and U17740 (N_17740,N_14915,N_14624);
nor U17741 (N_17741,N_14518,N_14729);
nor U17742 (N_17742,N_14342,N_15586);
nor U17743 (N_17743,N_14315,N_14436);
xor U17744 (N_17744,N_15157,N_15090);
or U17745 (N_17745,N_14906,N_14352);
nor U17746 (N_17746,N_14745,N_14732);
and U17747 (N_17747,N_14274,N_14003);
nand U17748 (N_17748,N_14711,N_14799);
or U17749 (N_17749,N_15787,N_14608);
nand U17750 (N_17750,N_14332,N_15814);
nand U17751 (N_17751,N_15545,N_14854);
or U17752 (N_17752,N_15495,N_14371);
xor U17753 (N_17753,N_15413,N_14527);
and U17754 (N_17754,N_14579,N_15004);
or U17755 (N_17755,N_15586,N_14005);
and U17756 (N_17756,N_15083,N_14847);
nand U17757 (N_17757,N_15000,N_14889);
xnor U17758 (N_17758,N_15041,N_15344);
xnor U17759 (N_17759,N_15281,N_14700);
nand U17760 (N_17760,N_15495,N_14284);
and U17761 (N_17761,N_14366,N_15519);
xor U17762 (N_17762,N_15206,N_15921);
xor U17763 (N_17763,N_14430,N_15431);
xnor U17764 (N_17764,N_14824,N_15320);
or U17765 (N_17765,N_15624,N_15670);
nand U17766 (N_17766,N_14563,N_14312);
nor U17767 (N_17767,N_14544,N_15783);
or U17768 (N_17768,N_14696,N_15050);
xnor U17769 (N_17769,N_15947,N_15771);
nor U17770 (N_17770,N_14196,N_15961);
nand U17771 (N_17771,N_15749,N_14244);
nand U17772 (N_17772,N_15634,N_14392);
nand U17773 (N_17773,N_14598,N_14285);
xnor U17774 (N_17774,N_14372,N_15281);
nand U17775 (N_17775,N_14337,N_14892);
nand U17776 (N_17776,N_14771,N_15135);
or U17777 (N_17777,N_14639,N_14830);
nand U17778 (N_17778,N_15127,N_14508);
xor U17779 (N_17779,N_14217,N_14876);
nor U17780 (N_17780,N_15680,N_15273);
nor U17781 (N_17781,N_14353,N_15325);
or U17782 (N_17782,N_15466,N_15508);
and U17783 (N_17783,N_14618,N_14066);
nand U17784 (N_17784,N_14915,N_15177);
or U17785 (N_17785,N_14382,N_15558);
xnor U17786 (N_17786,N_15146,N_14336);
xor U17787 (N_17787,N_14521,N_14193);
or U17788 (N_17788,N_15197,N_14554);
xnor U17789 (N_17789,N_14212,N_14504);
or U17790 (N_17790,N_15036,N_14396);
or U17791 (N_17791,N_15132,N_14756);
nand U17792 (N_17792,N_15063,N_15475);
nor U17793 (N_17793,N_14744,N_15681);
nor U17794 (N_17794,N_14331,N_14432);
or U17795 (N_17795,N_15451,N_15449);
nor U17796 (N_17796,N_15773,N_14770);
or U17797 (N_17797,N_14644,N_15802);
and U17798 (N_17798,N_15532,N_15661);
nor U17799 (N_17799,N_15082,N_14986);
and U17800 (N_17800,N_15231,N_14870);
nor U17801 (N_17801,N_15742,N_15475);
or U17802 (N_17802,N_15656,N_14376);
nor U17803 (N_17803,N_14925,N_14212);
or U17804 (N_17804,N_14800,N_15172);
nor U17805 (N_17805,N_15518,N_15878);
and U17806 (N_17806,N_15048,N_15012);
xor U17807 (N_17807,N_14654,N_15695);
or U17808 (N_17808,N_14604,N_15316);
and U17809 (N_17809,N_14826,N_14489);
xnor U17810 (N_17810,N_14600,N_15218);
or U17811 (N_17811,N_15181,N_15525);
or U17812 (N_17812,N_14960,N_14304);
or U17813 (N_17813,N_14056,N_14832);
nand U17814 (N_17814,N_14692,N_15095);
nor U17815 (N_17815,N_14776,N_14076);
or U17816 (N_17816,N_15003,N_15638);
nor U17817 (N_17817,N_14723,N_15751);
xor U17818 (N_17818,N_14591,N_14023);
and U17819 (N_17819,N_14176,N_14942);
nand U17820 (N_17820,N_14417,N_15215);
nor U17821 (N_17821,N_15595,N_15270);
or U17822 (N_17822,N_15780,N_15073);
xnor U17823 (N_17823,N_15031,N_15831);
xor U17824 (N_17824,N_14418,N_15614);
nor U17825 (N_17825,N_15180,N_15160);
and U17826 (N_17826,N_15320,N_15592);
nand U17827 (N_17827,N_15749,N_14134);
xnor U17828 (N_17828,N_15040,N_15696);
xor U17829 (N_17829,N_15254,N_15874);
xor U17830 (N_17830,N_14148,N_15914);
and U17831 (N_17831,N_14453,N_15039);
xnor U17832 (N_17832,N_14302,N_14314);
and U17833 (N_17833,N_15104,N_15322);
nor U17834 (N_17834,N_14662,N_14157);
nand U17835 (N_17835,N_15185,N_15671);
and U17836 (N_17836,N_14302,N_15755);
or U17837 (N_17837,N_14319,N_15872);
nand U17838 (N_17838,N_14987,N_14473);
and U17839 (N_17839,N_14966,N_15244);
and U17840 (N_17840,N_15257,N_14413);
and U17841 (N_17841,N_14143,N_15196);
xnor U17842 (N_17842,N_14563,N_15954);
nor U17843 (N_17843,N_14401,N_15959);
nor U17844 (N_17844,N_14983,N_15494);
xnor U17845 (N_17845,N_14520,N_15240);
or U17846 (N_17846,N_14432,N_15322);
or U17847 (N_17847,N_14874,N_14625);
or U17848 (N_17848,N_15858,N_15860);
nor U17849 (N_17849,N_14880,N_15308);
xor U17850 (N_17850,N_15536,N_15344);
and U17851 (N_17851,N_15423,N_15446);
or U17852 (N_17852,N_14699,N_14317);
xnor U17853 (N_17853,N_15452,N_15820);
and U17854 (N_17854,N_15777,N_14210);
xnor U17855 (N_17855,N_14339,N_14927);
nor U17856 (N_17856,N_14556,N_15731);
or U17857 (N_17857,N_14903,N_15335);
nor U17858 (N_17858,N_15569,N_15770);
nor U17859 (N_17859,N_14778,N_14417);
xor U17860 (N_17860,N_15305,N_15828);
or U17861 (N_17861,N_14632,N_15572);
nor U17862 (N_17862,N_15914,N_15762);
xnor U17863 (N_17863,N_14388,N_14463);
nor U17864 (N_17864,N_14413,N_15617);
xnor U17865 (N_17865,N_14337,N_15288);
nor U17866 (N_17866,N_15796,N_15152);
and U17867 (N_17867,N_14614,N_14413);
xnor U17868 (N_17868,N_15198,N_15938);
and U17869 (N_17869,N_14697,N_15410);
nand U17870 (N_17870,N_15863,N_15222);
nand U17871 (N_17871,N_14627,N_15041);
or U17872 (N_17872,N_15792,N_15172);
nand U17873 (N_17873,N_15868,N_14985);
xor U17874 (N_17874,N_14274,N_14539);
nand U17875 (N_17875,N_15357,N_14991);
or U17876 (N_17876,N_15595,N_15941);
or U17877 (N_17877,N_14230,N_15452);
nor U17878 (N_17878,N_15456,N_14554);
xor U17879 (N_17879,N_14266,N_14444);
nand U17880 (N_17880,N_14307,N_14360);
xnor U17881 (N_17881,N_14063,N_15292);
and U17882 (N_17882,N_14395,N_15960);
or U17883 (N_17883,N_14428,N_14926);
nand U17884 (N_17884,N_15182,N_15298);
nor U17885 (N_17885,N_14818,N_14156);
and U17886 (N_17886,N_14844,N_15655);
xnor U17887 (N_17887,N_15838,N_14796);
or U17888 (N_17888,N_15134,N_15370);
and U17889 (N_17889,N_14955,N_15621);
and U17890 (N_17890,N_14599,N_14192);
nand U17891 (N_17891,N_15211,N_15687);
and U17892 (N_17892,N_14137,N_15307);
and U17893 (N_17893,N_14411,N_15102);
nand U17894 (N_17894,N_14804,N_15402);
or U17895 (N_17895,N_15121,N_15481);
nand U17896 (N_17896,N_14500,N_15359);
nor U17897 (N_17897,N_14719,N_15046);
xnor U17898 (N_17898,N_15663,N_14885);
or U17899 (N_17899,N_14455,N_15264);
xnor U17900 (N_17900,N_14366,N_14029);
xor U17901 (N_17901,N_15315,N_14504);
or U17902 (N_17902,N_15069,N_14870);
nor U17903 (N_17903,N_14778,N_14980);
and U17904 (N_17904,N_15455,N_14297);
and U17905 (N_17905,N_15199,N_14314);
xnor U17906 (N_17906,N_14806,N_14338);
xor U17907 (N_17907,N_15733,N_14758);
and U17908 (N_17908,N_14902,N_15128);
or U17909 (N_17909,N_15388,N_14878);
nor U17910 (N_17910,N_14042,N_15858);
or U17911 (N_17911,N_15313,N_14437);
and U17912 (N_17912,N_14766,N_14820);
nand U17913 (N_17913,N_15744,N_14971);
nand U17914 (N_17914,N_14532,N_15638);
and U17915 (N_17915,N_14702,N_14944);
nand U17916 (N_17916,N_15308,N_14078);
nor U17917 (N_17917,N_14469,N_15754);
and U17918 (N_17918,N_14769,N_14413);
nor U17919 (N_17919,N_15877,N_15010);
nor U17920 (N_17920,N_15676,N_14555);
xnor U17921 (N_17921,N_15307,N_14908);
nand U17922 (N_17922,N_15700,N_15071);
and U17923 (N_17923,N_14271,N_15926);
nor U17924 (N_17924,N_15886,N_15604);
or U17925 (N_17925,N_14433,N_14332);
and U17926 (N_17926,N_14596,N_14067);
and U17927 (N_17927,N_15458,N_15393);
nor U17928 (N_17928,N_15073,N_14659);
and U17929 (N_17929,N_14235,N_14366);
xnor U17930 (N_17930,N_15564,N_15466);
nor U17931 (N_17931,N_15317,N_14684);
and U17932 (N_17932,N_14488,N_14740);
and U17933 (N_17933,N_14793,N_14419);
xnor U17934 (N_17934,N_15169,N_15484);
or U17935 (N_17935,N_15214,N_14132);
nand U17936 (N_17936,N_15839,N_14988);
nor U17937 (N_17937,N_14501,N_14429);
nor U17938 (N_17938,N_14032,N_15754);
or U17939 (N_17939,N_14964,N_15711);
nor U17940 (N_17940,N_14209,N_15423);
or U17941 (N_17941,N_15127,N_14743);
nor U17942 (N_17942,N_15930,N_15306);
or U17943 (N_17943,N_14986,N_14362);
or U17944 (N_17944,N_14992,N_14253);
xor U17945 (N_17945,N_14876,N_14228);
and U17946 (N_17946,N_14612,N_14871);
xnor U17947 (N_17947,N_15712,N_15760);
nor U17948 (N_17948,N_14764,N_14264);
nand U17949 (N_17949,N_15290,N_15479);
or U17950 (N_17950,N_15644,N_14907);
nand U17951 (N_17951,N_14604,N_14419);
nand U17952 (N_17952,N_14804,N_14599);
or U17953 (N_17953,N_15318,N_15092);
or U17954 (N_17954,N_14451,N_14217);
nor U17955 (N_17955,N_15750,N_15723);
and U17956 (N_17956,N_15679,N_15338);
nor U17957 (N_17957,N_14151,N_15613);
nand U17958 (N_17958,N_15952,N_14075);
and U17959 (N_17959,N_14140,N_15374);
xnor U17960 (N_17960,N_15186,N_14135);
xor U17961 (N_17961,N_14231,N_14344);
xnor U17962 (N_17962,N_15623,N_14928);
nor U17963 (N_17963,N_14440,N_14260);
or U17964 (N_17964,N_14138,N_15031);
or U17965 (N_17965,N_15334,N_14769);
xor U17966 (N_17966,N_14311,N_15158);
or U17967 (N_17967,N_15161,N_15439);
nor U17968 (N_17968,N_14838,N_15176);
and U17969 (N_17969,N_14281,N_15982);
nand U17970 (N_17970,N_15211,N_15420);
xor U17971 (N_17971,N_14887,N_14178);
xor U17972 (N_17972,N_14995,N_14556);
nand U17973 (N_17973,N_14308,N_15507);
xnor U17974 (N_17974,N_14950,N_15241);
and U17975 (N_17975,N_15786,N_15224);
xor U17976 (N_17976,N_14270,N_14268);
xor U17977 (N_17977,N_14265,N_15611);
xnor U17978 (N_17978,N_15303,N_14535);
or U17979 (N_17979,N_14904,N_14534);
nand U17980 (N_17980,N_14850,N_14896);
or U17981 (N_17981,N_14471,N_15664);
xor U17982 (N_17982,N_14077,N_14611);
and U17983 (N_17983,N_14635,N_14532);
xor U17984 (N_17984,N_15247,N_15884);
or U17985 (N_17985,N_14007,N_15025);
nand U17986 (N_17986,N_14909,N_15824);
or U17987 (N_17987,N_15431,N_15402);
or U17988 (N_17988,N_15108,N_14910);
xor U17989 (N_17989,N_15146,N_15296);
or U17990 (N_17990,N_14600,N_14729);
or U17991 (N_17991,N_15953,N_15781);
or U17992 (N_17992,N_15199,N_15365);
nand U17993 (N_17993,N_14935,N_14323);
nand U17994 (N_17994,N_14227,N_15862);
or U17995 (N_17995,N_15645,N_15264);
or U17996 (N_17996,N_14192,N_15703);
xnor U17997 (N_17997,N_15651,N_15410);
or U17998 (N_17998,N_14385,N_15870);
and U17999 (N_17999,N_14449,N_15222);
xnor U18000 (N_18000,N_16436,N_16762);
nand U18001 (N_18001,N_17777,N_17396);
or U18002 (N_18002,N_16990,N_17940);
nor U18003 (N_18003,N_16405,N_17436);
nor U18004 (N_18004,N_17857,N_16159);
or U18005 (N_18005,N_17805,N_17788);
or U18006 (N_18006,N_17025,N_17644);
and U18007 (N_18007,N_16863,N_17115);
nor U18008 (N_18008,N_16321,N_16134);
xnor U18009 (N_18009,N_17840,N_16169);
nor U18010 (N_18010,N_17884,N_17511);
nand U18011 (N_18011,N_16805,N_16688);
nand U18012 (N_18012,N_16227,N_17889);
and U18013 (N_18013,N_17712,N_16474);
and U18014 (N_18014,N_16322,N_17019);
or U18015 (N_18015,N_17223,N_17070);
xnor U18016 (N_18016,N_17688,N_16555);
or U18017 (N_18017,N_17091,N_17759);
or U18018 (N_18018,N_17819,N_16291);
nand U18019 (N_18019,N_17228,N_16786);
or U18020 (N_18020,N_16437,N_16387);
nor U18021 (N_18021,N_17670,N_16923);
or U18022 (N_18022,N_16293,N_16820);
xor U18023 (N_18023,N_16734,N_17903);
nand U18024 (N_18024,N_17166,N_17835);
and U18025 (N_18025,N_16592,N_16070);
nand U18026 (N_18026,N_16206,N_17135);
nor U18027 (N_18027,N_16010,N_16913);
xnor U18028 (N_18028,N_17462,N_16535);
and U18029 (N_18029,N_17333,N_17660);
and U18030 (N_18030,N_17807,N_17191);
or U18031 (N_18031,N_17230,N_17495);
and U18032 (N_18032,N_16229,N_16720);
or U18033 (N_18033,N_17621,N_17862);
or U18034 (N_18034,N_17939,N_17614);
nand U18035 (N_18035,N_16658,N_16003);
nand U18036 (N_18036,N_16794,N_17211);
and U18037 (N_18037,N_16237,N_17311);
xnor U18038 (N_18038,N_17365,N_16578);
nand U18039 (N_18039,N_17162,N_16957);
and U18040 (N_18040,N_17737,N_16386);
xor U18041 (N_18041,N_17420,N_17180);
nor U18042 (N_18042,N_16438,N_16097);
or U18043 (N_18043,N_16123,N_16701);
nand U18044 (N_18044,N_17957,N_16766);
nor U18045 (N_18045,N_16187,N_17993);
nand U18046 (N_18046,N_17765,N_17848);
and U18047 (N_18047,N_16966,N_17978);
or U18048 (N_18048,N_17685,N_16162);
or U18049 (N_18049,N_17183,N_17446);
and U18050 (N_18050,N_17624,N_16675);
or U18051 (N_18051,N_16171,N_17932);
and U18052 (N_18052,N_16788,N_17547);
or U18053 (N_18053,N_16938,N_16796);
nand U18054 (N_18054,N_17798,N_17813);
or U18055 (N_18055,N_17584,N_16396);
xnor U18056 (N_18056,N_16116,N_17970);
xnor U18057 (N_18057,N_17533,N_16281);
nor U18058 (N_18058,N_16672,N_16248);
nand U18059 (N_18059,N_17770,N_17871);
nor U18060 (N_18060,N_17029,N_17176);
xor U18061 (N_18061,N_16088,N_17042);
xor U18062 (N_18062,N_17640,N_16349);
or U18063 (N_18063,N_16458,N_16409);
nand U18064 (N_18064,N_16414,N_17906);
and U18065 (N_18065,N_16754,N_16965);
xnor U18066 (N_18066,N_16098,N_16582);
nand U18067 (N_18067,N_17052,N_17874);
or U18068 (N_18068,N_16031,N_16566);
nor U18069 (N_18069,N_17910,N_17376);
nor U18070 (N_18070,N_16091,N_16967);
and U18071 (N_18071,N_17307,N_17698);
xnor U18072 (N_18072,N_16308,N_17060);
or U18073 (N_18073,N_17161,N_17847);
and U18074 (N_18074,N_16263,N_16154);
nand U18075 (N_18075,N_17404,N_17157);
nor U18076 (N_18076,N_17449,N_16970);
nand U18077 (N_18077,N_16502,N_16363);
and U18078 (N_18078,N_16935,N_17682);
nor U18079 (N_18079,N_16001,N_17207);
nor U18080 (N_18080,N_17309,N_17145);
xnor U18081 (N_18081,N_17429,N_17124);
xnor U18082 (N_18082,N_17268,N_17753);
nand U18083 (N_18083,N_16225,N_16579);
and U18084 (N_18084,N_17633,N_17796);
and U18085 (N_18085,N_16252,N_17310);
nor U18086 (N_18086,N_17968,N_16201);
and U18087 (N_18087,N_17266,N_16175);
nor U18088 (N_18088,N_16523,N_16122);
and U18089 (N_18089,N_16163,N_17986);
nor U18090 (N_18090,N_16583,N_16121);
or U18091 (N_18091,N_16027,N_17755);
nand U18092 (N_18092,N_16993,N_16849);
xnor U18093 (N_18093,N_17861,N_17590);
or U18094 (N_18094,N_16912,N_17062);
nor U18095 (N_18095,N_16017,N_17817);
nor U18096 (N_18096,N_17540,N_16039);
or U18097 (N_18097,N_16055,N_17959);
or U18098 (N_18098,N_16898,N_17214);
nand U18099 (N_18099,N_17832,N_17087);
nand U18100 (N_18100,N_16499,N_17530);
nor U18101 (N_18101,N_17262,N_17233);
nor U18102 (N_18102,N_17278,N_16310);
nand U18103 (N_18103,N_17041,N_17470);
nor U18104 (N_18104,N_17177,N_16807);
xor U18105 (N_18105,N_17395,N_16595);
xnor U18106 (N_18106,N_17487,N_16011);
and U18107 (N_18107,N_16899,N_17219);
and U18108 (N_18108,N_17438,N_16633);
or U18109 (N_18109,N_17163,N_16197);
nand U18110 (N_18110,N_16369,N_16346);
and U18111 (N_18111,N_16258,N_16576);
nor U18112 (N_18112,N_16265,N_17460);
and U18113 (N_18113,N_16767,N_16973);
and U18114 (N_18114,N_17295,N_17814);
and U18115 (N_18115,N_17601,N_16478);
xnor U18116 (N_18116,N_16932,N_16850);
or U18117 (N_18117,N_16226,N_17471);
nand U18118 (N_18118,N_17631,N_17064);
and U18119 (N_18119,N_16251,N_17238);
or U18120 (N_18120,N_16541,N_16267);
or U18121 (N_18121,N_17342,N_16832);
nor U18122 (N_18122,N_16961,N_16282);
xor U18123 (N_18123,N_16462,N_17141);
nand U18124 (N_18124,N_17224,N_17885);
and U18125 (N_18125,N_17024,N_16096);
nor U18126 (N_18126,N_16273,N_16681);
and U18127 (N_18127,N_16002,N_16545);
or U18128 (N_18128,N_17564,N_16066);
xnor U18129 (N_18129,N_16606,N_16764);
or U18130 (N_18130,N_17764,N_17281);
nand U18131 (N_18131,N_17683,N_16234);
xor U18132 (N_18132,N_17694,N_17469);
nand U18133 (N_18133,N_17121,N_17137);
or U18134 (N_18134,N_17702,N_17156);
nand U18135 (N_18135,N_17269,N_17909);
nor U18136 (N_18136,N_17200,N_16869);
xor U18137 (N_18137,N_16599,N_17732);
xor U18138 (N_18138,N_16848,N_16765);
and U18139 (N_18139,N_17724,N_17567);
nand U18140 (N_18140,N_16909,N_17231);
or U18141 (N_18141,N_17105,N_17627);
or U18142 (N_18142,N_16079,N_17237);
or U18143 (N_18143,N_16433,N_17696);
or U18144 (N_18144,N_17119,N_17594);
nand U18145 (N_18145,N_17865,N_17397);
nand U18146 (N_18146,N_16315,N_17852);
nand U18147 (N_18147,N_17984,N_17506);
and U18148 (N_18148,N_17022,N_17719);
nor U18149 (N_18149,N_16419,N_16657);
nand U18150 (N_18150,N_17808,N_16731);
or U18151 (N_18151,N_17983,N_16507);
or U18152 (N_18152,N_17314,N_17246);
or U18153 (N_18153,N_16926,N_17328);
or U18154 (N_18154,N_16365,N_16275);
nand U18155 (N_18155,N_16558,N_17913);
nand U18156 (N_18156,N_16008,N_17801);
nor U18157 (N_18157,N_16650,N_16646);
nor U18158 (N_18158,N_17632,N_17824);
nand U18159 (N_18159,N_16800,N_16316);
and U18160 (N_18160,N_16485,N_17083);
nand U18161 (N_18161,N_17854,N_16895);
nand U18162 (N_18162,N_17227,N_17418);
and U18163 (N_18163,N_16435,N_16110);
xnor U18164 (N_18164,N_17198,N_16808);
and U18165 (N_18165,N_17665,N_17241);
nor U18166 (N_18166,N_17744,N_16245);
nand U18167 (N_18167,N_16843,N_16751);
nor U18168 (N_18168,N_16306,N_16907);
and U18169 (N_18169,N_17155,N_16540);
or U18170 (N_18170,N_16420,N_17403);
nand U18171 (N_18171,N_17747,N_17629);
nor U18172 (N_18172,N_17958,N_16812);
xor U18173 (N_18173,N_17437,N_17989);
and U18174 (N_18174,N_16454,N_17148);
nand U18175 (N_18175,N_17315,N_17346);
nor U18176 (N_18176,N_17464,N_17040);
xnor U18177 (N_18177,N_16773,N_17351);
or U18178 (N_18178,N_16571,N_17969);
nand U18179 (N_18179,N_17804,N_16689);
and U18180 (N_18180,N_17528,N_17373);
xnor U18181 (N_18181,N_16126,N_17714);
and U18182 (N_18182,N_16586,N_17409);
nor U18183 (N_18183,N_16603,N_16569);
nand U18184 (N_18184,N_16094,N_17305);
or U18185 (N_18185,N_17008,N_16219);
nand U18186 (N_18186,N_16391,N_16030);
and U18187 (N_18187,N_16568,N_16286);
nor U18188 (N_18188,N_17878,N_16718);
nor U18189 (N_18189,N_17662,N_17297);
or U18190 (N_18190,N_17419,N_17456);
and U18191 (N_18191,N_17806,N_16732);
and U18192 (N_18192,N_16573,N_17159);
nand U18193 (N_18193,N_17357,N_17525);
xnor U18194 (N_18194,N_17339,N_17676);
or U18195 (N_18195,N_16194,N_16232);
nor U18196 (N_18196,N_16213,N_17381);
nand U18197 (N_18197,N_16905,N_17941);
nand U18198 (N_18198,N_16500,N_17619);
nand U18199 (N_18199,N_16312,N_16472);
nand U18200 (N_18200,N_17782,N_16294);
or U18201 (N_18201,N_17267,N_16709);
xor U18202 (N_18202,N_16934,N_16401);
xnor U18203 (N_18203,N_17543,N_17317);
xor U18204 (N_18204,N_16262,N_16092);
and U18205 (N_18205,N_17630,N_16906);
or U18206 (N_18206,N_17285,N_17844);
or U18207 (N_18207,N_17868,N_16590);
nor U18208 (N_18208,N_16374,N_16975);
xnor U18209 (N_18209,N_17360,N_17192);
nor U18210 (N_18210,N_17474,N_16285);
and U18211 (N_18211,N_17879,N_17028);
nor U18212 (N_18212,N_17457,N_16461);
xnor U18213 (N_18213,N_16109,N_17208);
nand U18214 (N_18214,N_17050,N_17542);
and U18215 (N_18215,N_17972,N_16519);
or U18216 (N_18216,N_17997,N_17673);
xnor U18217 (N_18217,N_16418,N_16356);
nand U18218 (N_18218,N_16914,N_16609);
or U18219 (N_18219,N_16528,N_17242);
and U18220 (N_18220,N_16944,N_17946);
and U18221 (N_18221,N_17182,N_17501);
nor U18222 (N_18222,N_16803,N_17658);
nor U18223 (N_18223,N_16127,N_17034);
and U18224 (N_18224,N_17738,N_16743);
and U18225 (N_18225,N_17820,N_16133);
nand U18226 (N_18226,N_17664,N_16652);
and U18227 (N_18227,N_16594,N_16928);
or U18228 (N_18228,N_16292,N_16852);
xnor U18229 (N_18229,N_16522,N_17125);
and U18230 (N_18230,N_16342,N_16903);
xor U18231 (N_18231,N_17049,N_16168);
nand U18232 (N_18232,N_16693,N_16793);
or U18233 (N_18233,N_16798,N_17800);
nor U18234 (N_18234,N_17992,N_17341);
xor U18235 (N_18235,N_16212,N_16028);
and U18236 (N_18236,N_17952,N_17810);
or U18237 (N_18237,N_16868,N_17519);
or U18238 (N_18238,N_17850,N_16503);
nor U18239 (N_18239,N_17197,N_17094);
nand U18240 (N_18240,N_16198,N_17802);
nand U18241 (N_18241,N_17385,N_16704);
xnor U18242 (N_18242,N_17065,N_17152);
xnor U18243 (N_18243,N_17170,N_16388);
nand U18244 (N_18244,N_16955,N_17518);
xor U18245 (N_18245,N_17595,N_16880);
and U18246 (N_18246,N_16750,N_16918);
nand U18247 (N_18247,N_16649,N_17510);
nand U18248 (N_18248,N_16196,N_17102);
nor U18249 (N_18249,N_17799,N_16441);
and U18250 (N_18250,N_17608,N_17489);
and U18251 (N_18251,N_16891,N_16685);
nand U18252 (N_18252,N_17054,N_17776);
and U18253 (N_18253,N_16642,N_17006);
nand U18254 (N_18254,N_16986,N_17118);
and U18255 (N_18255,N_17195,N_17549);
xnor U18256 (N_18256,N_17563,N_16301);
or U18257 (N_18257,N_17826,N_17063);
xnor U18258 (N_18258,N_16236,N_16825);
nor U18259 (N_18259,N_16431,N_16644);
xnor U18260 (N_18260,N_17488,N_17911);
and U18261 (N_18261,N_16239,N_17090);
nand U18262 (N_18262,N_16287,N_16640);
nor U18263 (N_18263,N_16819,N_16412);
and U18264 (N_18264,N_17925,N_17966);
nor U18265 (N_18265,N_16288,N_17340);
or U18266 (N_18266,N_16884,N_17888);
or U18267 (N_18267,N_17153,N_17706);
xor U18268 (N_18268,N_16370,N_16543);
nor U18269 (N_18269,N_16982,N_17383);
nor U18270 (N_18270,N_17916,N_17016);
nand U18271 (N_18271,N_17362,N_16785);
nor U18272 (N_18272,N_17828,N_16131);
xor U18273 (N_18273,N_17920,N_17545);
or U18274 (N_18274,N_16814,N_16733);
nand U18275 (N_18275,N_16948,N_16108);
xor U18276 (N_18276,N_17203,N_17407);
nor U18277 (N_18277,N_16656,N_17181);
or U18278 (N_18278,N_17569,N_16980);
nor U18279 (N_18279,N_16679,N_16671);
nand U18280 (N_18280,N_17015,N_16333);
and U18281 (N_18281,N_17654,N_16509);
nor U18282 (N_18282,N_16632,N_17769);
nor U18283 (N_18283,N_17226,N_17494);
xor U18284 (N_18284,N_16997,N_16538);
and U18285 (N_18285,N_16223,N_17412);
nand U18286 (N_18286,N_16337,N_17736);
or U18287 (N_18287,N_17037,N_17723);
nor U18288 (N_18288,N_17215,N_17423);
and U18289 (N_18289,N_16553,N_17821);
nand U18290 (N_18290,N_17922,N_16802);
or U18291 (N_18291,N_17031,N_16466);
and U18292 (N_18292,N_17338,N_17294);
or U18293 (N_18293,N_17604,N_16985);
or U18294 (N_18294,N_16402,N_17277);
xor U18295 (N_18295,N_16491,N_17898);
xor U18296 (N_18296,N_16327,N_16560);
nor U18297 (N_18297,N_16596,N_16591);
and U18298 (N_18298,N_17768,N_16249);
or U18299 (N_18299,N_17308,N_16741);
or U18300 (N_18300,N_17554,N_16371);
nand U18301 (N_18301,N_17445,N_17582);
xnor U18302 (N_18302,N_16775,N_17974);
or U18303 (N_18303,N_16151,N_17739);
nand U18304 (N_18304,N_16083,N_16328);
xor U18305 (N_18305,N_17144,N_17918);
nor U18306 (N_18306,N_17674,N_17875);
nor U18307 (N_18307,N_16887,N_16958);
and U18308 (N_18308,N_17709,N_17822);
and U18309 (N_18309,N_16824,N_16953);
and U18310 (N_18310,N_16790,N_16853);
xnor U18311 (N_18311,N_17692,N_16467);
or U18312 (N_18312,N_16084,N_16639);
nand U18313 (N_18313,N_16866,N_17484);
nand U18314 (N_18314,N_17876,N_17441);
and U18315 (N_18315,N_16900,N_16736);
xnor U18316 (N_18316,N_16470,N_17615);
nor U18317 (N_18317,N_16125,N_17032);
or U18318 (N_18318,N_16574,N_16006);
nand U18319 (N_18319,N_17524,N_17949);
nand U18320 (N_18320,N_17873,N_17477);
nor U18321 (N_18321,N_16902,N_17565);
nor U18322 (N_18322,N_17523,N_17715);
nand U18323 (N_18323,N_16620,N_17526);
xnor U18324 (N_18324,N_16859,N_16460);
nand U18325 (N_18325,N_16300,N_17963);
nor U18326 (N_18326,N_16115,N_17539);
nand U18327 (N_18327,N_16057,N_16145);
nor U18328 (N_18328,N_16564,N_17675);
and U18329 (N_18329,N_17686,N_16886);
xnor U18330 (N_18330,N_16770,N_17815);
or U18331 (N_18331,N_16577,N_17646);
nor U18332 (N_18332,N_17504,N_16314);
nand U18333 (N_18333,N_16231,N_16960);
xor U18334 (N_18334,N_17435,N_16468);
nand U18335 (N_18335,N_16137,N_17842);
nor U18336 (N_18336,N_16015,N_16627);
xnor U18337 (N_18337,N_16214,N_17727);
xor U18338 (N_18338,N_17113,N_16837);
or U18339 (N_18339,N_16394,N_17369);
or U18340 (N_18340,N_17812,N_16284);
and U18341 (N_18341,N_16994,N_16715);
nor U18342 (N_18342,N_16455,N_16525);
and U18343 (N_18343,N_17078,N_17803);
nand U18344 (N_18344,N_16303,N_17379);
or U18345 (N_18345,N_17893,N_17666);
nand U18346 (N_18346,N_16271,N_17047);
and U18347 (N_18347,N_17167,N_17048);
and U18348 (N_18348,N_17058,N_17560);
nand U18349 (N_18349,N_16009,N_16992);
nand U18350 (N_18350,N_16012,N_16457);
nor U18351 (N_18351,N_16411,N_16013);
and U18352 (N_18352,N_17829,N_17264);
nand U18353 (N_18353,N_17741,N_17387);
or U18354 (N_18354,N_17074,N_17790);
nand U18355 (N_18355,N_17240,N_16447);
xor U18356 (N_18356,N_17252,N_16876);
and U18357 (N_18357,N_17718,N_16324);
nand U18358 (N_18358,N_16473,N_17934);
nand U18359 (N_18359,N_16811,N_17274);
or U18360 (N_18360,N_16514,N_16516);
xor U18361 (N_18361,N_17599,N_17372);
nand U18362 (N_18362,N_16052,N_16546);
xnor U18363 (N_18363,N_17845,N_16508);
xnor U18364 (N_18364,N_17864,N_16721);
nand U18365 (N_18365,N_17981,N_16998);
and U18366 (N_18366,N_16730,N_17089);
xnor U18367 (N_18367,N_17475,N_17251);
nand U18368 (N_18368,N_17985,N_17209);
and U18369 (N_18369,N_17575,N_16724);
nand U18370 (N_18370,N_16873,N_16020);
and U18371 (N_18371,N_17072,N_16691);
xor U18372 (N_18372,N_16915,N_16476);
and U18373 (N_18373,N_16243,N_16389);
or U18374 (N_18374,N_16927,N_17760);
or U18375 (N_18375,N_17668,N_17669);
xor U18376 (N_18376,N_17093,N_16554);
and U18377 (N_18377,N_16073,N_17923);
or U18378 (N_18378,N_16618,N_16677);
and U18379 (N_18379,N_17243,N_17010);
or U18380 (N_18380,N_16240,N_17026);
or U18381 (N_18381,N_17443,N_17742);
nand U18382 (N_18382,N_16302,N_16138);
nor U18383 (N_18383,N_17147,N_17610);
or U18384 (N_18384,N_17110,N_17421);
xnor U18385 (N_18385,N_17452,N_17573);
xor U18386 (N_18386,N_16362,N_16836);
nor U18387 (N_18387,N_16102,N_16373);
or U18388 (N_18388,N_16539,N_16061);
and U18389 (N_18389,N_16183,N_16180);
nor U18390 (N_18390,N_17129,N_17516);
nor U18391 (N_18391,N_16497,N_16779);
and U18392 (N_18392,N_16833,N_16729);
nor U18393 (N_18393,N_17336,N_16043);
nand U18394 (N_18394,N_16429,N_17392);
nand U18395 (N_18395,N_16864,N_17576);
nand U18396 (N_18396,N_16524,N_17035);
and U18397 (N_18397,N_17882,N_16581);
or U18398 (N_18398,N_16984,N_16044);
nor U18399 (N_18399,N_17361,N_17391);
xnor U18400 (N_18400,N_17282,N_16233);
and U18401 (N_18401,N_16385,N_16381);
nor U18402 (N_18402,N_17905,N_16593);
or U18403 (N_18403,N_17169,N_17534);
nor U18404 (N_18404,N_17809,N_17345);
or U18405 (N_18405,N_17347,N_17779);
or U18406 (N_18406,N_16075,N_16439);
or U18407 (N_18407,N_16763,N_16746);
nor U18408 (N_18408,N_17432,N_16924);
nand U18409 (N_18409,N_17960,N_17684);
xnor U18410 (N_18410,N_17187,N_17303);
nor U18411 (N_18411,N_16427,N_17825);
and U18412 (N_18412,N_17165,N_17433);
nor U18413 (N_18413,N_17127,N_17935);
nand U18414 (N_18414,N_17117,N_17350);
xor U18415 (N_18415,N_16320,N_16352);
nand U18416 (N_18416,N_17716,N_16921);
nand U18417 (N_18417,N_16246,N_16426);
xor U18418 (N_18418,N_16166,N_17454);
nand U18419 (N_18419,N_16247,N_17831);
and U18420 (N_18420,N_16334,N_16529);
or U18421 (N_18421,N_17912,N_17580);
xnor U18422 (N_18422,N_16339,N_16547);
nor U18423 (N_18423,N_16482,N_16826);
nand U18424 (N_18424,N_16112,N_16158);
xnor U18425 (N_18425,N_16113,N_17971);
nand U18426 (N_18426,N_17174,N_17258);
or U18427 (N_18427,N_16834,N_16963);
and U18428 (N_18428,N_16380,N_17577);
nand U18429 (N_18429,N_17917,N_16655);
or U18430 (N_18430,N_16318,N_16550);
nor U18431 (N_18431,N_17870,N_17261);
and U18432 (N_18432,N_16208,N_16710);
nand U18433 (N_18433,N_17143,N_16047);
nand U18434 (N_18434,N_16890,N_17571);
xor U18435 (N_18435,N_17926,N_16674);
nand U18436 (N_18436,N_16635,N_16256);
and U18437 (N_18437,N_16257,N_17961);
and U18438 (N_18438,N_17908,N_16533);
nor U18439 (N_18439,N_17834,N_16141);
and U18440 (N_18440,N_17617,N_16019);
xor U18441 (N_18441,N_16737,N_16795);
and U18442 (N_18442,N_16492,N_16192);
nor U18443 (N_18443,N_17626,N_16086);
or U18444 (N_18444,N_17408,N_16559);
xor U18445 (N_18445,N_16996,N_17216);
xnor U18446 (N_18446,N_17212,N_17425);
nand U18447 (N_18447,N_17703,N_16597);
and U18448 (N_18448,N_16977,N_17492);
nand U18449 (N_18449,N_17232,N_16952);
xnor U18450 (N_18450,N_16705,N_17559);
nor U18451 (N_18451,N_17111,N_16176);
xnor U18452 (N_18452,N_16959,N_16034);
or U18453 (N_18453,N_16222,N_16615);
nand U18454 (N_18454,N_17607,N_17318);
and U18455 (N_18455,N_16165,N_17532);
or U18456 (N_18456,N_17481,N_17229);
xor U18457 (N_18457,N_16621,N_17355);
and U18458 (N_18458,N_16424,N_16081);
xor U18459 (N_18459,N_17907,N_17273);
or U18460 (N_18460,N_17792,N_16202);
nor U18461 (N_18461,N_16801,N_17793);
xnor U18462 (N_18462,N_17455,N_16442);
or U18463 (N_18463,N_17440,N_16397);
and U18464 (N_18464,N_17887,N_16261);
or U18465 (N_18465,N_17003,N_17306);
or U18466 (N_18466,N_16871,N_16648);
xnor U18467 (N_18467,N_16033,N_17919);
or U18468 (N_18468,N_17109,N_16534);
or U18469 (N_18469,N_17424,N_17036);
or U18470 (N_18470,N_17012,N_17073);
and U18471 (N_18471,N_16215,N_17394);
nand U18472 (N_18472,N_17199,N_16062);
nand U18473 (N_18473,N_17027,N_16089);
nand U18474 (N_18474,N_17883,N_16182);
xnor U18475 (N_18475,N_17767,N_16146);
xor U18476 (N_18476,N_16999,N_16498);
nand U18477 (N_18477,N_16673,N_16305);
nand U18478 (N_18478,N_16742,N_16587);
or U18479 (N_18479,N_17393,N_16377);
or U18480 (N_18480,N_16050,N_17374);
and U18481 (N_18481,N_16617,N_17158);
nand U18482 (N_18482,N_17221,N_17500);
and U18483 (N_18483,N_16778,N_16643);
xor U18484 (N_18484,N_16759,N_16738);
or U18485 (N_18485,N_17461,N_17132);
nor U18486 (N_18486,N_16465,N_16877);
nor U18487 (N_18487,N_17442,N_16799);
xnor U18488 (N_18488,N_17656,N_16383);
and U18489 (N_18489,N_17886,N_17657);
nor U18490 (N_18490,N_16128,N_16025);
or U18491 (N_18491,N_16400,N_16311);
nand U18492 (N_18492,N_16575,N_17894);
or U18493 (N_18493,N_17597,N_17075);
nor U18494 (N_18494,N_16359,N_17616);
nand U18495 (N_18495,N_17818,N_16493);
xnor U18496 (N_18496,N_17996,N_17931);
nor U18497 (N_18497,N_17515,N_17687);
xor U18498 (N_18498,N_16771,N_17370);
or U18499 (N_18499,N_17699,N_16404);
or U18500 (N_18500,N_17179,N_16189);
xnor U18501 (N_18501,N_16562,N_16809);
or U18502 (N_18502,N_17600,N_17323);
or U18503 (N_18503,N_16813,N_17173);
xnor U18504 (N_18504,N_17000,N_17044);
nand U18505 (N_18505,N_16883,N_16432);
and U18506 (N_18506,N_16974,N_16277);
nor U18507 (N_18507,N_17752,N_17947);
or U18508 (N_18508,N_17680,N_16692);
nor U18509 (N_18509,N_17579,N_17859);
or U18510 (N_18510,N_16885,N_16797);
and U18511 (N_18511,N_16584,N_16469);
and U18512 (N_18512,N_16124,N_17150);
xnor U18513 (N_18513,N_17522,N_16755);
xor U18514 (N_18514,N_16893,N_16854);
and U18515 (N_18515,N_17976,N_17605);
and U18516 (N_18516,N_17586,N_17750);
nand U18517 (N_18517,N_17018,N_16422);
nor U18518 (N_18518,N_16361,N_16760);
nand U18519 (N_18519,N_16260,N_16074);
xnor U18520 (N_18520,N_17422,N_17239);
nor U18521 (N_18521,N_17609,N_17256);
nand U18522 (N_18522,N_16513,N_16250);
or U18523 (N_18523,N_17327,N_16911);
or U18524 (N_18524,N_17995,N_16831);
nor U18525 (N_18525,N_17249,N_17001);
nand U18526 (N_18526,N_17248,N_17439);
nand U18527 (N_18527,N_17955,N_17690);
nand U18528 (N_18528,N_17869,N_16254);
nor U18529 (N_18529,N_16270,N_17552);
or U18530 (N_18530,N_17371,N_17717);
nor U18531 (N_18531,N_17938,N_16040);
and U18532 (N_18532,N_16604,N_17039);
and U18533 (N_18533,N_17546,N_16542);
nor U18534 (N_18534,N_16631,N_17076);
or U18535 (N_18535,N_16317,N_17478);
nand U18536 (N_18536,N_17700,N_16341);
and U18537 (N_18537,N_16204,N_16152);
or U18538 (N_18538,N_16283,N_16343);
or U18539 (N_18539,N_16570,N_16143);
or U18540 (N_18540,N_17950,N_17771);
or U18541 (N_18541,N_17596,N_17568);
nand U18542 (N_18542,N_16398,N_17128);
or U18543 (N_18543,N_17398,N_17322);
and U18544 (N_18544,N_16393,N_16345);
nor U18545 (N_18545,N_17914,N_16660);
xor U18546 (N_18546,N_16894,N_16634);
xnor U18547 (N_18547,N_16036,N_17139);
and U18548 (N_18548,N_17337,N_17611);
xnor U18549 (N_18549,N_16136,N_16572);
nor U18550 (N_18550,N_16789,N_16399);
nor U18551 (N_18551,N_16612,N_16188);
or U18552 (N_18552,N_17713,N_17795);
or U18553 (N_18553,N_17766,N_16329);
nor U18554 (N_18554,N_16372,N_16607);
xor U18555 (N_18555,N_16666,N_16818);
xor U18556 (N_18556,N_16756,N_16408);
xor U18557 (N_18557,N_17009,N_17561);
and U18558 (N_18558,N_17411,N_16563);
xnor U18559 (N_18559,N_17275,N_16827);
or U18560 (N_18560,N_17250,N_16551);
nor U18561 (N_18561,N_16087,N_16971);
nor U18562 (N_18562,N_17740,N_16682);
nor U18563 (N_18563,N_17830,N_16667);
xnor U18564 (N_18564,N_17671,N_16839);
and U18565 (N_18565,N_17431,N_16445);
xor U18566 (N_18566,N_17388,N_16014);
xor U18567 (N_18567,N_17652,N_16179);
nand U18568 (N_18568,N_17763,N_17591);
nand U18569 (N_18569,N_16780,N_16144);
nand U18570 (N_18570,N_16191,N_17466);
xnor U18571 (N_18571,N_17772,N_16787);
or U18572 (N_18572,N_16727,N_16872);
nand U18573 (N_18573,N_16861,N_16964);
and U18574 (N_18574,N_16815,N_16969);
nor U18575 (N_18575,N_17043,N_17537);
xnor U18576 (N_18576,N_16100,N_17055);
xor U18577 (N_18577,N_16280,N_16937);
xor U18578 (N_18578,N_16276,N_16471);
and U18579 (N_18579,N_17497,N_16224);
and U18580 (N_18580,N_16451,N_17566);
nor U18581 (N_18581,N_16114,N_16683);
nand U18582 (N_18582,N_16810,N_17710);
or U18583 (N_18583,N_16661,N_17583);
xor U18584 (N_18584,N_17945,N_16968);
and U18585 (N_18585,N_17020,N_16483);
and U18586 (N_18586,N_17786,N_16129);
or U18587 (N_18587,N_17289,N_17175);
nor U18588 (N_18588,N_16295,N_17891);
or U18589 (N_18589,N_16676,N_16105);
nand U18590 (N_18590,N_17486,N_16769);
and U18591 (N_18591,N_17705,N_16700);
and U18592 (N_18592,N_16989,N_16049);
nor U18593 (N_18593,N_17998,N_16238);
nor U18594 (N_18594,N_17321,N_16611);
nor U18595 (N_18595,N_17300,N_16181);
xor U18596 (N_18596,N_17701,N_16987);
or U18597 (N_18597,N_16244,N_16641);
and U18598 (N_18598,N_16716,N_16253);
nand U18599 (N_18599,N_16338,N_16135);
nand U18600 (N_18600,N_16032,N_16490);
or U18601 (N_18601,N_17728,N_16456);
or U18602 (N_18602,N_17544,N_17099);
xor U18603 (N_18603,N_17726,N_17131);
or U18604 (N_18604,N_17555,N_17618);
nand U18605 (N_18605,N_16453,N_16624);
nor U18606 (N_18606,N_17146,N_17693);
or U18607 (N_18607,N_16614,N_17721);
xnor U18608 (N_18608,N_16892,N_16046);
xnor U18609 (N_18609,N_17450,N_16619);
xnor U18610 (N_18610,N_16170,N_17098);
nor U18611 (N_18611,N_17378,N_16368);
nand U18612 (N_18612,N_17399,N_17051);
nand U18613 (N_18613,N_16983,N_17287);
nand U18614 (N_18614,N_16268,N_16297);
nand U18615 (N_18615,N_16494,N_17140);
nand U18616 (N_18616,N_16228,N_17491);
nor U18617 (N_18617,N_16857,N_17202);
nor U18618 (N_18618,N_17377,N_16217);
xor U18619 (N_18619,N_17138,N_16446);
nand U18620 (N_18620,N_17071,N_16830);
nand U18621 (N_18621,N_16567,N_17293);
and U18622 (N_18622,N_16059,N_17836);
xnor U18623 (N_18623,N_17206,N_17781);
or U18624 (N_18624,N_17944,N_16416);
nor U18625 (N_18625,N_17480,N_16000);
or U18626 (N_18626,N_17628,N_16140);
nor U18627 (N_18627,N_17007,N_16821);
or U18628 (N_18628,N_16690,N_16120);
and U18629 (N_18629,N_16298,N_17401);
xnor U18630 (N_18630,N_16678,N_17973);
nor U18631 (N_18631,N_17603,N_16065);
xnor U18632 (N_18632,N_16623,N_17405);
nand U18633 (N_18633,N_17553,N_16153);
nand U18634 (N_18634,N_16782,N_16920);
and U18635 (N_18635,N_17841,N_16919);
or U18636 (N_18636,N_17651,N_17521);
or U18637 (N_18637,N_16406,N_16904);
and U18638 (N_18638,N_17312,N_17168);
and U18639 (N_18639,N_16726,N_16651);
xor U18640 (N_18640,N_17234,N_16023);
nor U18641 (N_18641,N_16748,N_16939);
and U18642 (N_18642,N_17904,N_17194);
and U18643 (N_18643,N_17330,N_16024);
nor U18644 (N_18644,N_16495,N_16723);
xnor U18645 (N_18645,N_17201,N_16326);
and U18646 (N_18646,N_17833,N_16323);
and U18647 (N_18647,N_16255,N_16069);
xnor U18648 (N_18648,N_17639,N_16160);
and U18649 (N_18649,N_16351,N_17053);
xnor U18650 (N_18650,N_17758,N_16931);
xnor U18651 (N_18651,N_17103,N_16379);
nand U18652 (N_18652,N_17430,N_17116);
or U18653 (N_18653,N_17787,N_17288);
nand U18654 (N_18654,N_17389,N_16216);
or U18655 (N_18655,N_16496,N_17691);
nand U18656 (N_18656,N_16366,N_16669);
nor U18657 (N_18657,N_16209,N_16290);
or U18658 (N_18658,N_16613,N_16549);
and U18659 (N_18659,N_17236,N_16450);
nand U18660 (N_18660,N_16304,N_16942);
nand U18661 (N_18661,N_17620,N_17529);
xnor U18662 (N_18662,N_16600,N_17107);
xnor U18663 (N_18663,N_17270,N_17069);
nor U18664 (N_18664,N_17205,N_16925);
nor U18665 (N_18665,N_17059,N_17837);
xnor U18666 (N_18666,N_16486,N_16702);
nor U18667 (N_18667,N_16309,N_17136);
xnor U18668 (N_18668,N_17190,N_16950);
nor U18669 (N_18669,N_17979,N_17353);
and U18670 (N_18670,N_17877,N_17855);
nand U18671 (N_18671,N_16510,N_17217);
xor U18672 (N_18672,N_17088,N_16077);
xnor U18673 (N_18673,N_17468,N_17733);
xnor U18674 (N_18674,N_17068,N_16791);
xnor U18675 (N_18675,N_17689,N_16860);
nor U18676 (N_18676,N_17097,N_16719);
xnor U18677 (N_18677,N_16714,N_16829);
and U18678 (N_18678,N_16758,N_16364);
xnor U18679 (N_18679,N_17196,N_16588);
xnor U18680 (N_18680,N_17218,N_17811);
xnor U18681 (N_18681,N_16879,N_16585);
or U18682 (N_18682,N_17292,N_16781);
or U18683 (N_18683,N_16605,N_16536);
and U18684 (N_18684,N_17637,N_17980);
and U18685 (N_18685,N_16668,N_17271);
or U18686 (N_18686,N_17114,N_16484);
nand U18687 (N_18687,N_17975,N_17447);
nand U18688 (N_18688,N_17382,N_16929);
nand U18689 (N_18689,N_17101,N_16164);
nand U18690 (N_18690,N_16459,N_17587);
and U18691 (N_18691,N_17707,N_17602);
xnor U18692 (N_18692,N_16777,N_16289);
or U18693 (N_18693,N_16745,N_16336);
nand U18694 (N_18694,N_16428,N_16744);
xor U18695 (N_18695,N_17517,N_17794);
or U18696 (N_18696,N_16107,N_17678);
xor U18697 (N_18697,N_16479,N_17106);
nor U18698 (N_18698,N_17520,N_16085);
and U18699 (N_18699,N_16694,N_16761);
nor U18700 (N_18700,N_16045,N_17329);
or U18701 (N_18701,N_16021,N_17046);
nand U18702 (N_18702,N_16357,N_17302);
and U18703 (N_18703,N_17863,N_16947);
nor U18704 (N_18704,N_16264,N_17756);
and U18705 (N_18705,N_17204,N_16862);
or U18706 (N_18706,N_16005,N_17415);
nand U18707 (N_18707,N_17942,N_16841);
xnor U18708 (N_18708,N_16527,N_17638);
nor U18709 (N_18709,N_16518,N_17535);
nor U18710 (N_18710,N_17987,N_16858);
or U18711 (N_18711,N_16064,N_16150);
and U18712 (N_18712,N_16664,N_17550);
and U18713 (N_18713,N_17663,N_16235);
nand U18714 (N_18714,N_17359,N_16207);
nand U18715 (N_18715,N_17354,N_16425);
nand U18716 (N_18716,N_17080,N_17483);
and U18717 (N_18717,N_16350,N_17964);
nand U18718 (N_18718,N_17352,N_17897);
nand U18719 (N_18719,N_16299,N_17164);
or U18720 (N_18720,N_17220,N_17254);
nand U18721 (N_18721,N_17247,N_16665);
or U18722 (N_18722,N_16018,N_17259);
nand U18723 (N_18723,N_17210,N_16142);
nand U18724 (N_18724,N_17849,N_16995);
nand U18725 (N_18725,N_16403,N_17364);
and U18726 (N_18726,N_17326,N_17120);
nor U18727 (N_18727,N_16622,N_17498);
nor U18728 (N_18728,N_17536,N_17943);
nand U18729 (N_18729,N_16056,N_16784);
and U18730 (N_18730,N_16772,N_16625);
xnor U18731 (N_18731,N_17593,N_16846);
and U18732 (N_18732,N_16557,N_16804);
and U18733 (N_18733,N_16917,N_16728);
or U18734 (N_18734,N_16417,N_17749);
nor U18735 (N_18735,N_16697,N_16526);
nand U18736 (N_18736,N_17313,N_16104);
nand U18737 (N_18737,N_17778,N_17558);
nor U18738 (N_18738,N_17505,N_17895);
xor U18739 (N_18739,N_16279,N_16353);
and U18740 (N_18740,N_17901,N_17780);
and U18741 (N_18741,N_16930,N_17123);
nand U18742 (N_18742,N_17990,N_16882);
xnor U18743 (N_18743,N_16531,N_16082);
and U18744 (N_18744,N_17298,N_16035);
or U18745 (N_18745,N_16068,N_17092);
nor U18746 (N_18746,N_16972,N_16449);
and U18747 (N_18747,N_16487,N_17458);
or U18748 (N_18748,N_17838,N_16747);
or U18749 (N_18749,N_17257,N_17735);
nor U18750 (N_18750,N_17056,N_17541);
and U18751 (N_18751,N_17086,N_17783);
nor U18752 (N_18752,N_17635,N_17711);
or U18753 (N_18753,N_16376,N_16828);
nor U18754 (N_18754,N_17570,N_16195);
or U18755 (N_18755,N_16544,N_17606);
xnor U18756 (N_18756,N_16042,N_17773);
nor U18757 (N_18757,N_17649,N_17245);
xnor U18758 (N_18758,N_17299,N_16696);
or U18759 (N_18759,N_16463,N_17067);
and U18760 (N_18760,N_17746,N_17473);
or U18761 (N_18761,N_17112,N_16768);
xnor U18762 (N_18762,N_17472,N_17410);
xnor U18763 (N_18763,N_16347,N_17380);
nand U18764 (N_18764,N_16090,N_17133);
nand U18765 (N_18765,N_17017,N_16630);
nand U18766 (N_18766,N_17304,N_17244);
nand U18767 (N_18767,N_16067,N_17708);
and U18768 (N_18768,N_16161,N_16367);
nor U18769 (N_18769,N_16517,N_16395);
or U18770 (N_18770,N_16481,N_17356);
xor U18771 (N_18771,N_16936,N_17924);
xnor U18772 (N_18772,N_17320,N_16601);
nand U18773 (N_18773,N_16026,N_16278);
xnor U18774 (N_18774,N_17867,N_17704);
or U18775 (N_18775,N_16007,N_17858);
and U18776 (N_18776,N_17592,N_17459);
or U18777 (N_18777,N_17358,N_16241);
nor U18778 (N_18778,N_17178,N_17933);
and U18779 (N_18779,N_17962,N_16856);
nor U18780 (N_18780,N_16155,N_16991);
or U18781 (N_18781,N_16628,N_16515);
xor U18782 (N_18782,N_16410,N_16602);
or U18783 (N_18783,N_17636,N_17499);
and U18784 (N_18784,N_17324,N_17490);
nand U18785 (N_18785,N_17095,N_16157);
nand U18786 (N_18786,N_16865,N_16713);
nand U18787 (N_18787,N_17562,N_17390);
and U18788 (N_18788,N_16608,N_16933);
or U18789 (N_18789,N_16978,N_17077);
nand U18790 (N_18790,N_16325,N_17647);
or U18791 (N_18791,N_16211,N_16193);
or U18792 (N_18792,N_17667,N_17023);
nand U18793 (N_18793,N_16348,N_17745);
nand U18794 (N_18794,N_16296,N_17400);
and U18795 (N_18795,N_16060,N_17623);
and U18796 (N_18796,N_16016,N_16130);
xor U18797 (N_18797,N_17557,N_17784);
nor U18798 (N_18798,N_16413,N_17827);
nand U18799 (N_18799,N_17375,N_17014);
and U18800 (N_18800,N_16699,N_17476);
nand U18801 (N_18801,N_16378,N_16687);
nand U18802 (N_18802,N_16382,N_16156);
and U18803 (N_18803,N_17507,N_17030);
or U18804 (N_18804,N_17225,N_17762);
xnor U18805 (N_18805,N_16703,N_16200);
or U18806 (N_18806,N_17856,N_17276);
nor U18807 (N_18807,N_17625,N_16940);
nor U18808 (N_18808,N_16663,N_17937);
xnor U18809 (N_18809,N_17413,N_16897);
xnor U18810 (N_18810,N_17982,N_17291);
xor U18811 (N_18811,N_17479,N_16205);
nand U18812 (N_18812,N_17512,N_17186);
or U18813 (N_18813,N_16340,N_17896);
and U18814 (N_18814,N_17927,N_16659);
or U18815 (N_18815,N_16307,N_16177);
xor U18816 (N_18816,N_17084,N_17816);
or U18817 (N_18817,N_17574,N_17427);
nand U18818 (N_18818,N_17589,N_16580);
xor U18819 (N_18819,N_17253,N_17823);
and U18820 (N_18820,N_16637,N_16415);
or U18821 (N_18821,N_16078,N_16616);
or U18822 (N_18822,N_17160,N_17038);
nand U18823 (N_18823,N_16847,N_16922);
and U18824 (N_18824,N_17672,N_17551);
nor U18825 (N_18825,N_17929,N_16118);
xor U18826 (N_18826,N_16330,N_16203);
nor U18827 (N_18827,N_17743,N_17731);
or U18828 (N_18828,N_17451,N_16941);
nor U18829 (N_18829,N_17283,N_17643);
nand U18830 (N_18830,N_17722,N_16421);
and U18831 (N_18831,N_16949,N_17066);
nand U18832 (N_18832,N_17754,N_16054);
xnor U18833 (N_18833,N_17645,N_17222);
or U18834 (N_18834,N_16806,N_16489);
nor U18835 (N_18835,N_16776,N_17011);
nand U18836 (N_18836,N_17751,N_17343);
xor U18837 (N_18837,N_16822,N_17921);
nor U18838 (N_18838,N_17661,N_17255);
nor U18839 (N_18839,N_16556,N_16331);
xnor U18840 (N_18840,N_17791,N_16269);
xor U18841 (N_18841,N_16392,N_17033);
nand U18842 (N_18842,N_16888,N_17426);
xnor U18843 (N_18843,N_16230,N_17622);
xnor U18844 (N_18844,N_16259,N_17588);
and U18845 (N_18845,N_17509,N_17977);
nand U18846 (N_18846,N_17846,N_16735);
nor U18847 (N_18847,N_16851,N_16173);
and U18848 (N_18848,N_17444,N_16186);
or U18849 (N_18849,N_16916,N_17503);
nand U18850 (N_18850,N_17880,N_16855);
nor U18851 (N_18851,N_16477,N_16448);
and U18852 (N_18852,N_17057,N_17004);
xnor U18853 (N_18853,N_16440,N_16335);
nor U18854 (N_18854,N_17612,N_17100);
and U18855 (N_18855,N_16976,N_16511);
xnor U18856 (N_18856,N_16274,N_16512);
nand U18857 (N_18857,N_16095,N_16501);
or U18858 (N_18858,N_17463,N_17448);
nor U18859 (N_18859,N_17485,N_17892);
nand U18860 (N_18860,N_17348,N_17860);
and U18861 (N_18861,N_16117,N_17482);
xnor U18862 (N_18862,N_16444,N_17502);
nand U18863 (N_18863,N_16475,N_17316);
nor U18864 (N_18864,N_16598,N_16874);
xnor U18865 (N_18865,N_17697,N_17839);
nor U18866 (N_18866,N_16654,N_17386);
and U18867 (N_18867,N_17154,N_17002);
nor U18868 (N_18868,N_17866,N_17578);
nor U18869 (N_18869,N_16506,N_17548);
nor U18870 (N_18870,N_17677,N_16053);
nand U18871 (N_18871,N_17999,N_17193);
nand U18872 (N_18872,N_17349,N_17296);
or U18873 (N_18873,N_16384,N_17681);
and U18874 (N_18874,N_17402,N_16954);
nor U18875 (N_18875,N_16344,N_16185);
nand U18876 (N_18876,N_16712,N_16452);
xor U18877 (N_18877,N_16842,N_17881);
or U18878 (N_18878,N_17598,N_16103);
and U18879 (N_18879,N_16711,N_16739);
and U18880 (N_18880,N_16167,N_16817);
or U18881 (N_18881,N_17951,N_17453);
nand U18882 (N_18882,N_16707,N_16823);
xnor U18883 (N_18883,N_17332,N_17096);
xor U18884 (N_18884,N_17899,N_16038);
or U18885 (N_18885,N_16878,N_16908);
nand U18886 (N_18886,N_17108,N_16354);
or U18887 (N_18887,N_17720,N_16844);
and U18888 (N_18888,N_16840,N_16210);
or U18889 (N_18889,N_16910,N_16647);
or U18890 (N_18890,N_17417,N_17319);
nand U18891 (N_18891,N_17414,N_16753);
nand U18892 (N_18892,N_17994,N_16190);
nand U18893 (N_18893,N_17334,N_16147);
xnor U18894 (N_18894,N_17493,N_16722);
or U18895 (N_18895,N_17384,N_17853);
and U18896 (N_18896,N_17280,N_17556);
nand U18897 (N_18897,N_17104,N_16537);
and U18898 (N_18898,N_16148,N_17367);
nand U18899 (N_18899,N_17991,N_17428);
and U18900 (N_18900,N_16423,N_17954);
nand U18901 (N_18901,N_16111,N_16093);
xor U18902 (N_18902,N_17213,N_17581);
xor U18903 (N_18903,N_16072,N_16532);
and U18904 (N_18904,N_16565,N_16816);
nor U18905 (N_18905,N_16119,N_17513);
nand U18906 (N_18906,N_16695,N_17290);
or U18907 (N_18907,N_16783,N_16548);
nor U18908 (N_18908,N_16943,N_17527);
and U18909 (N_18909,N_17650,N_16218);
nand U18910 (N_18910,N_16708,N_16220);
nor U18911 (N_18911,N_16048,N_17585);
or U18912 (N_18912,N_17021,N_17953);
or U18913 (N_18913,N_16132,N_17368);
and U18914 (N_18914,N_17514,N_16717);
and U18915 (N_18915,N_17260,N_16149);
nor U18916 (N_18916,N_16221,N_16184);
and U18917 (N_18917,N_17081,N_16174);
nor U18918 (N_18918,N_17725,N_17775);
or U18919 (N_18919,N_16080,N_17797);
nor U18920 (N_18920,N_17172,N_17496);
and U18921 (N_18921,N_17653,N_17956);
xnor U18922 (N_18922,N_16945,N_17967);
nor U18923 (N_18923,N_17928,N_16434);
or U18924 (N_18924,N_17761,N_17843);
and U18925 (N_18925,N_16313,N_16706);
or U18926 (N_18926,N_17344,N_16725);
nand U18927 (N_18927,N_16752,N_16172);
nand U18928 (N_18928,N_16029,N_16561);
xnor U18929 (N_18929,N_17126,N_16875);
xnor U18930 (N_18930,N_16051,N_16951);
nand U18931 (N_18931,N_17757,N_16757);
nor U18932 (N_18932,N_17272,N_16684);
nand U18933 (N_18933,N_16645,N_17872);
or U18934 (N_18934,N_17915,N_16004);
xor U18935 (N_18935,N_17900,N_16071);
or U18936 (N_18936,N_17301,N_16870);
nand U18937 (N_18937,N_17363,N_16375);
or U18938 (N_18938,N_17122,N_16063);
and U18939 (N_18939,N_17648,N_16530);
nor U18940 (N_18940,N_17188,N_17538);
and U18941 (N_18941,N_16774,N_17988);
xnor U18942 (N_18942,N_16653,N_16037);
nand U18943 (N_18943,N_17149,N_17265);
nand U18944 (N_18944,N_16178,N_16199);
or U18945 (N_18945,N_17902,N_17142);
nand U18946 (N_18946,N_17655,N_16332);
nor U18947 (N_18947,N_16662,N_16896);
and U18948 (N_18948,N_16358,N_16355);
or U18949 (N_18949,N_16360,N_17185);
nor U18950 (N_18950,N_16740,N_17634);
and U18951 (N_18951,N_16988,N_16610);
and U18952 (N_18952,N_17785,N_16058);
nor U18953 (N_18953,N_17965,N_17774);
xnor U18954 (N_18954,N_17286,N_17366);
nor U18955 (N_18955,N_17930,N_17851);
nor U18956 (N_18956,N_17335,N_16636);
or U18957 (N_18957,N_16981,N_17572);
and U18958 (N_18958,N_16901,N_17184);
nand U18959 (N_18959,N_16520,N_16319);
or U18960 (N_18960,N_16946,N_17531);
xnor U18961 (N_18961,N_16979,N_16521);
and U18962 (N_18962,N_17613,N_16670);
xnor U18963 (N_18963,N_17151,N_16407);
nand U18964 (N_18964,N_17134,N_16430);
xor U18965 (N_18965,N_16076,N_17734);
xor U18966 (N_18966,N_17695,N_16488);
xor U18967 (N_18967,N_17331,N_17748);
nor U18968 (N_18968,N_16686,N_16889);
or U18969 (N_18969,N_16552,N_17279);
nand U18970 (N_18970,N_17659,N_16480);
and U18971 (N_18971,N_16680,N_16242);
nand U18972 (N_18972,N_16099,N_16749);
xor U18973 (N_18973,N_17045,N_17189);
nor U18974 (N_18974,N_17890,N_16272);
and U18975 (N_18975,N_16835,N_17013);
nor U18976 (N_18976,N_16504,N_17730);
nor U18977 (N_18977,N_16838,N_17061);
nor U18978 (N_18978,N_16464,N_17130);
nor U18979 (N_18979,N_17434,N_16589);
and U18980 (N_18980,N_16139,N_16266);
nand U18981 (N_18981,N_16443,N_17936);
or U18982 (N_18982,N_17235,N_17284);
or U18983 (N_18983,N_17085,N_16867);
nand U18984 (N_18984,N_17789,N_16962);
nor U18985 (N_18985,N_17082,N_17467);
nand U18986 (N_18986,N_16101,N_16505);
or U18987 (N_18987,N_16629,N_17948);
and U18988 (N_18988,N_17641,N_16956);
nor U18989 (N_18989,N_17416,N_17005);
or U18990 (N_18990,N_17729,N_17508);
xnor U18991 (N_18991,N_16041,N_17263);
or U18992 (N_18992,N_17465,N_16698);
nand U18993 (N_18993,N_17642,N_16881);
nor U18994 (N_18994,N_17406,N_16022);
nand U18995 (N_18995,N_16638,N_16626);
xnor U18996 (N_18996,N_17171,N_16792);
nor U18997 (N_18997,N_17325,N_17079);
xor U18998 (N_18998,N_17679,N_16390);
and U18999 (N_18999,N_16845,N_16106);
and U19000 (N_19000,N_16798,N_17452);
or U19001 (N_19001,N_16558,N_17128);
nor U19002 (N_19002,N_17907,N_16985);
and U19003 (N_19003,N_16657,N_17306);
nand U19004 (N_19004,N_16399,N_17713);
nor U19005 (N_19005,N_16824,N_16079);
or U19006 (N_19006,N_16083,N_16949);
nand U19007 (N_19007,N_17053,N_16222);
nand U19008 (N_19008,N_17065,N_16395);
nor U19009 (N_19009,N_17030,N_16385);
xnor U19010 (N_19010,N_17985,N_17333);
and U19011 (N_19011,N_16919,N_17528);
nor U19012 (N_19012,N_17304,N_17876);
nand U19013 (N_19013,N_16424,N_16377);
nand U19014 (N_19014,N_16827,N_16924);
and U19015 (N_19015,N_16221,N_16514);
nand U19016 (N_19016,N_16946,N_16651);
nor U19017 (N_19017,N_16598,N_17406);
or U19018 (N_19018,N_16357,N_17242);
xnor U19019 (N_19019,N_17146,N_16299);
or U19020 (N_19020,N_17341,N_16679);
nand U19021 (N_19021,N_17340,N_17189);
nand U19022 (N_19022,N_17463,N_17335);
nor U19023 (N_19023,N_17297,N_16485);
xnor U19024 (N_19024,N_16458,N_17850);
nor U19025 (N_19025,N_17547,N_16626);
or U19026 (N_19026,N_16757,N_16498);
or U19027 (N_19027,N_17275,N_17233);
nand U19028 (N_19028,N_16427,N_17175);
nand U19029 (N_19029,N_17110,N_16297);
and U19030 (N_19030,N_17045,N_16137);
nand U19031 (N_19031,N_16092,N_17997);
or U19032 (N_19032,N_16133,N_16508);
or U19033 (N_19033,N_16582,N_17762);
xor U19034 (N_19034,N_17912,N_16275);
xnor U19035 (N_19035,N_16396,N_16613);
xor U19036 (N_19036,N_17548,N_17651);
or U19037 (N_19037,N_17535,N_16803);
nor U19038 (N_19038,N_16595,N_17975);
and U19039 (N_19039,N_17512,N_16856);
nor U19040 (N_19040,N_16036,N_16585);
and U19041 (N_19041,N_17074,N_17981);
nand U19042 (N_19042,N_16225,N_16370);
nand U19043 (N_19043,N_16697,N_17427);
and U19044 (N_19044,N_16271,N_17994);
xnor U19045 (N_19045,N_16287,N_16240);
or U19046 (N_19046,N_17122,N_17061);
and U19047 (N_19047,N_16674,N_17134);
nand U19048 (N_19048,N_16360,N_17644);
xor U19049 (N_19049,N_16581,N_16463);
xor U19050 (N_19050,N_17697,N_17724);
and U19051 (N_19051,N_17936,N_17605);
nand U19052 (N_19052,N_16272,N_16878);
xor U19053 (N_19053,N_16477,N_16485);
and U19054 (N_19054,N_16877,N_17470);
nand U19055 (N_19055,N_17754,N_17042);
or U19056 (N_19056,N_17174,N_16730);
and U19057 (N_19057,N_16641,N_17104);
nor U19058 (N_19058,N_16836,N_16406);
and U19059 (N_19059,N_16647,N_17285);
nor U19060 (N_19060,N_16587,N_17023);
or U19061 (N_19061,N_16494,N_16433);
or U19062 (N_19062,N_17942,N_17364);
or U19063 (N_19063,N_17026,N_16626);
nor U19064 (N_19064,N_16804,N_16798);
and U19065 (N_19065,N_16609,N_17406);
nor U19066 (N_19066,N_17465,N_17020);
nand U19067 (N_19067,N_16759,N_17106);
or U19068 (N_19068,N_16626,N_16865);
or U19069 (N_19069,N_16438,N_17547);
nor U19070 (N_19070,N_16773,N_16188);
or U19071 (N_19071,N_16151,N_16378);
nand U19072 (N_19072,N_16331,N_17426);
and U19073 (N_19073,N_17600,N_16216);
nand U19074 (N_19074,N_17008,N_17806);
and U19075 (N_19075,N_16398,N_17543);
xnor U19076 (N_19076,N_17913,N_17446);
and U19077 (N_19077,N_17505,N_16179);
or U19078 (N_19078,N_17030,N_17387);
or U19079 (N_19079,N_16928,N_16819);
and U19080 (N_19080,N_17065,N_17928);
nor U19081 (N_19081,N_17468,N_17067);
or U19082 (N_19082,N_16614,N_17511);
nor U19083 (N_19083,N_16880,N_16253);
xnor U19084 (N_19084,N_16700,N_16045);
nand U19085 (N_19085,N_16309,N_16658);
nand U19086 (N_19086,N_17333,N_17055);
nand U19087 (N_19087,N_17446,N_16532);
and U19088 (N_19088,N_17431,N_16907);
xnor U19089 (N_19089,N_17602,N_17485);
or U19090 (N_19090,N_17136,N_17426);
and U19091 (N_19091,N_17109,N_17576);
xnor U19092 (N_19092,N_16578,N_17063);
nand U19093 (N_19093,N_16953,N_16759);
and U19094 (N_19094,N_17743,N_17865);
xor U19095 (N_19095,N_17440,N_17644);
or U19096 (N_19096,N_17692,N_16269);
nor U19097 (N_19097,N_16977,N_17523);
nand U19098 (N_19098,N_17057,N_17098);
nand U19099 (N_19099,N_17300,N_17045);
nand U19100 (N_19100,N_17679,N_17977);
or U19101 (N_19101,N_17884,N_17776);
nor U19102 (N_19102,N_17865,N_16042);
or U19103 (N_19103,N_17210,N_16800);
nor U19104 (N_19104,N_17654,N_17231);
and U19105 (N_19105,N_16251,N_17998);
or U19106 (N_19106,N_17949,N_16656);
or U19107 (N_19107,N_17147,N_16595);
nand U19108 (N_19108,N_17400,N_17289);
and U19109 (N_19109,N_17768,N_17817);
or U19110 (N_19110,N_16514,N_16189);
and U19111 (N_19111,N_16174,N_17055);
nand U19112 (N_19112,N_16836,N_16033);
nor U19113 (N_19113,N_17714,N_16666);
and U19114 (N_19114,N_17487,N_17199);
or U19115 (N_19115,N_17637,N_16920);
nand U19116 (N_19116,N_16872,N_17527);
and U19117 (N_19117,N_17674,N_16087);
xor U19118 (N_19118,N_17947,N_16494);
and U19119 (N_19119,N_16698,N_16518);
or U19120 (N_19120,N_17668,N_16010);
and U19121 (N_19121,N_16084,N_16457);
xnor U19122 (N_19122,N_16107,N_16371);
and U19123 (N_19123,N_16468,N_16615);
and U19124 (N_19124,N_17042,N_17660);
xnor U19125 (N_19125,N_17827,N_17605);
nor U19126 (N_19126,N_16882,N_17677);
or U19127 (N_19127,N_17758,N_17130);
or U19128 (N_19128,N_16329,N_16693);
xnor U19129 (N_19129,N_17683,N_17687);
xor U19130 (N_19130,N_17482,N_16476);
xor U19131 (N_19131,N_17190,N_16042);
nand U19132 (N_19132,N_16652,N_16079);
xor U19133 (N_19133,N_17726,N_17800);
or U19134 (N_19134,N_17916,N_17639);
or U19135 (N_19135,N_16496,N_17334);
or U19136 (N_19136,N_17804,N_16123);
xor U19137 (N_19137,N_16581,N_16158);
or U19138 (N_19138,N_16853,N_17560);
xnor U19139 (N_19139,N_16488,N_16873);
nor U19140 (N_19140,N_17034,N_17773);
or U19141 (N_19141,N_17861,N_16642);
or U19142 (N_19142,N_16398,N_17657);
xnor U19143 (N_19143,N_16984,N_17874);
and U19144 (N_19144,N_16389,N_16532);
and U19145 (N_19145,N_17341,N_17258);
xnor U19146 (N_19146,N_16235,N_17896);
and U19147 (N_19147,N_16323,N_16816);
nand U19148 (N_19148,N_16315,N_17168);
xnor U19149 (N_19149,N_17250,N_17679);
nand U19150 (N_19150,N_16506,N_16255);
xor U19151 (N_19151,N_17210,N_16492);
xnor U19152 (N_19152,N_17237,N_16841);
and U19153 (N_19153,N_17135,N_16514);
nor U19154 (N_19154,N_17692,N_16686);
and U19155 (N_19155,N_17743,N_16283);
nor U19156 (N_19156,N_16133,N_16955);
nor U19157 (N_19157,N_17972,N_17036);
nand U19158 (N_19158,N_16462,N_16985);
and U19159 (N_19159,N_17320,N_17220);
xnor U19160 (N_19160,N_16077,N_16837);
and U19161 (N_19161,N_17040,N_16403);
nand U19162 (N_19162,N_16214,N_16986);
xnor U19163 (N_19163,N_16981,N_16627);
nor U19164 (N_19164,N_17064,N_16127);
or U19165 (N_19165,N_17960,N_16471);
or U19166 (N_19166,N_16971,N_16310);
and U19167 (N_19167,N_16536,N_16564);
and U19168 (N_19168,N_17415,N_17584);
and U19169 (N_19169,N_16133,N_16859);
and U19170 (N_19170,N_16103,N_17050);
or U19171 (N_19171,N_17040,N_16800);
xnor U19172 (N_19172,N_17709,N_16966);
and U19173 (N_19173,N_16261,N_16052);
xor U19174 (N_19174,N_16222,N_16927);
or U19175 (N_19175,N_17299,N_17430);
nor U19176 (N_19176,N_17121,N_17338);
nor U19177 (N_19177,N_16725,N_17114);
nor U19178 (N_19178,N_17253,N_17299);
nor U19179 (N_19179,N_16580,N_16655);
nand U19180 (N_19180,N_16768,N_17756);
nor U19181 (N_19181,N_16036,N_17535);
xnor U19182 (N_19182,N_16056,N_17627);
xnor U19183 (N_19183,N_17876,N_17379);
nand U19184 (N_19184,N_16036,N_16535);
and U19185 (N_19185,N_16537,N_16095);
or U19186 (N_19186,N_17879,N_17491);
and U19187 (N_19187,N_16677,N_17377);
xor U19188 (N_19188,N_16696,N_16249);
and U19189 (N_19189,N_16750,N_17561);
xor U19190 (N_19190,N_17015,N_16507);
xor U19191 (N_19191,N_17754,N_16725);
and U19192 (N_19192,N_16929,N_17354);
nand U19193 (N_19193,N_17097,N_16679);
nand U19194 (N_19194,N_17495,N_16660);
xnor U19195 (N_19195,N_17769,N_16792);
and U19196 (N_19196,N_17650,N_17246);
nand U19197 (N_19197,N_17347,N_16790);
nor U19198 (N_19198,N_17671,N_17343);
nor U19199 (N_19199,N_16402,N_17926);
nor U19200 (N_19200,N_16102,N_17973);
or U19201 (N_19201,N_16402,N_17431);
nor U19202 (N_19202,N_17586,N_16758);
or U19203 (N_19203,N_16955,N_17314);
nor U19204 (N_19204,N_16133,N_16682);
or U19205 (N_19205,N_16636,N_16915);
and U19206 (N_19206,N_17391,N_16964);
or U19207 (N_19207,N_17843,N_17647);
nand U19208 (N_19208,N_16757,N_16077);
nand U19209 (N_19209,N_17420,N_16376);
nand U19210 (N_19210,N_16025,N_17337);
nand U19211 (N_19211,N_16376,N_16665);
nand U19212 (N_19212,N_17192,N_16366);
and U19213 (N_19213,N_17425,N_16879);
nor U19214 (N_19214,N_17792,N_17489);
nand U19215 (N_19215,N_16556,N_16431);
nand U19216 (N_19216,N_16548,N_16433);
nor U19217 (N_19217,N_16007,N_16091);
and U19218 (N_19218,N_17347,N_16025);
nand U19219 (N_19219,N_16806,N_16236);
xor U19220 (N_19220,N_16710,N_16020);
or U19221 (N_19221,N_17663,N_17622);
or U19222 (N_19222,N_16835,N_16094);
nand U19223 (N_19223,N_16197,N_17590);
or U19224 (N_19224,N_17189,N_17529);
or U19225 (N_19225,N_16677,N_17737);
nand U19226 (N_19226,N_16063,N_17704);
nor U19227 (N_19227,N_17064,N_16729);
nand U19228 (N_19228,N_16388,N_17116);
or U19229 (N_19229,N_16645,N_16359);
xor U19230 (N_19230,N_16180,N_16606);
nor U19231 (N_19231,N_16045,N_16190);
nor U19232 (N_19232,N_16601,N_17903);
or U19233 (N_19233,N_17230,N_17787);
nand U19234 (N_19234,N_17056,N_17435);
or U19235 (N_19235,N_17057,N_17516);
or U19236 (N_19236,N_17917,N_17449);
nor U19237 (N_19237,N_17659,N_16835);
nand U19238 (N_19238,N_17105,N_16747);
and U19239 (N_19239,N_16167,N_16242);
or U19240 (N_19240,N_17315,N_17115);
and U19241 (N_19241,N_17431,N_16596);
xnor U19242 (N_19242,N_16739,N_16667);
nor U19243 (N_19243,N_16618,N_17660);
nor U19244 (N_19244,N_16697,N_16950);
nand U19245 (N_19245,N_17115,N_17829);
nand U19246 (N_19246,N_16525,N_16530);
xnor U19247 (N_19247,N_17390,N_17563);
or U19248 (N_19248,N_17143,N_16531);
or U19249 (N_19249,N_16194,N_17987);
and U19250 (N_19250,N_17339,N_17383);
or U19251 (N_19251,N_16056,N_16751);
nor U19252 (N_19252,N_17462,N_17133);
xor U19253 (N_19253,N_17038,N_16259);
nor U19254 (N_19254,N_17198,N_17862);
nor U19255 (N_19255,N_17157,N_17183);
and U19256 (N_19256,N_16644,N_17878);
and U19257 (N_19257,N_16449,N_16680);
or U19258 (N_19258,N_16328,N_16652);
xor U19259 (N_19259,N_16016,N_17978);
and U19260 (N_19260,N_16002,N_16614);
nand U19261 (N_19261,N_16043,N_16215);
and U19262 (N_19262,N_17225,N_16220);
or U19263 (N_19263,N_16611,N_17261);
nand U19264 (N_19264,N_17654,N_17090);
nand U19265 (N_19265,N_16910,N_16184);
or U19266 (N_19266,N_16307,N_17983);
or U19267 (N_19267,N_16290,N_16761);
nor U19268 (N_19268,N_16419,N_17216);
nor U19269 (N_19269,N_17683,N_17435);
xnor U19270 (N_19270,N_16723,N_16167);
nor U19271 (N_19271,N_16681,N_17799);
nor U19272 (N_19272,N_16371,N_17695);
and U19273 (N_19273,N_17223,N_16814);
nand U19274 (N_19274,N_17624,N_16561);
xor U19275 (N_19275,N_16109,N_17261);
or U19276 (N_19276,N_17076,N_17744);
xnor U19277 (N_19277,N_16974,N_16244);
or U19278 (N_19278,N_17943,N_17804);
xor U19279 (N_19279,N_16529,N_16627);
or U19280 (N_19280,N_17885,N_16923);
and U19281 (N_19281,N_16437,N_16647);
xor U19282 (N_19282,N_16819,N_16390);
and U19283 (N_19283,N_17098,N_17937);
nor U19284 (N_19284,N_17378,N_16888);
and U19285 (N_19285,N_17823,N_17767);
or U19286 (N_19286,N_17545,N_16920);
and U19287 (N_19287,N_16145,N_17534);
xor U19288 (N_19288,N_16329,N_16926);
nor U19289 (N_19289,N_16273,N_17013);
nand U19290 (N_19290,N_17050,N_16434);
nand U19291 (N_19291,N_17303,N_17861);
nand U19292 (N_19292,N_16254,N_16339);
nor U19293 (N_19293,N_16217,N_17191);
xor U19294 (N_19294,N_16660,N_17791);
nand U19295 (N_19295,N_17610,N_17076);
or U19296 (N_19296,N_16262,N_17922);
nor U19297 (N_19297,N_17065,N_16486);
nand U19298 (N_19298,N_17297,N_17056);
nor U19299 (N_19299,N_16651,N_16702);
xnor U19300 (N_19300,N_17600,N_17068);
or U19301 (N_19301,N_17258,N_17029);
or U19302 (N_19302,N_17507,N_16524);
and U19303 (N_19303,N_17087,N_16309);
and U19304 (N_19304,N_17767,N_17524);
nor U19305 (N_19305,N_16538,N_17613);
nand U19306 (N_19306,N_17075,N_17169);
or U19307 (N_19307,N_17608,N_17404);
or U19308 (N_19308,N_17365,N_16486);
nor U19309 (N_19309,N_17790,N_16049);
and U19310 (N_19310,N_17274,N_17004);
nand U19311 (N_19311,N_16749,N_16133);
xor U19312 (N_19312,N_16846,N_17650);
nor U19313 (N_19313,N_16221,N_17767);
nor U19314 (N_19314,N_16260,N_17738);
xnor U19315 (N_19315,N_16668,N_16760);
xnor U19316 (N_19316,N_16143,N_16698);
or U19317 (N_19317,N_16641,N_16416);
or U19318 (N_19318,N_17712,N_16220);
nand U19319 (N_19319,N_16321,N_17956);
nand U19320 (N_19320,N_17230,N_16818);
or U19321 (N_19321,N_17648,N_16834);
xnor U19322 (N_19322,N_16343,N_17921);
nand U19323 (N_19323,N_17378,N_17643);
nor U19324 (N_19324,N_16432,N_17875);
and U19325 (N_19325,N_16731,N_17846);
xnor U19326 (N_19326,N_17340,N_17030);
and U19327 (N_19327,N_17181,N_17527);
nor U19328 (N_19328,N_17964,N_16584);
xor U19329 (N_19329,N_16086,N_16688);
or U19330 (N_19330,N_16105,N_17485);
nor U19331 (N_19331,N_17051,N_17579);
nand U19332 (N_19332,N_17352,N_17389);
nor U19333 (N_19333,N_16841,N_16485);
nor U19334 (N_19334,N_16423,N_16502);
nand U19335 (N_19335,N_16967,N_16473);
or U19336 (N_19336,N_17704,N_17343);
xor U19337 (N_19337,N_17476,N_16095);
or U19338 (N_19338,N_17865,N_16747);
or U19339 (N_19339,N_16231,N_16407);
nand U19340 (N_19340,N_16192,N_16473);
and U19341 (N_19341,N_16960,N_16256);
xor U19342 (N_19342,N_17545,N_17749);
or U19343 (N_19343,N_17055,N_16585);
xnor U19344 (N_19344,N_17945,N_16977);
xor U19345 (N_19345,N_16086,N_16976);
nor U19346 (N_19346,N_16083,N_16659);
xnor U19347 (N_19347,N_16433,N_17958);
xor U19348 (N_19348,N_17568,N_17687);
nand U19349 (N_19349,N_16820,N_16768);
or U19350 (N_19350,N_17779,N_16850);
xor U19351 (N_19351,N_17115,N_17952);
and U19352 (N_19352,N_17498,N_17639);
or U19353 (N_19353,N_16934,N_17764);
nor U19354 (N_19354,N_16746,N_17956);
nor U19355 (N_19355,N_17953,N_17174);
or U19356 (N_19356,N_17977,N_16563);
nor U19357 (N_19357,N_17474,N_17009);
or U19358 (N_19358,N_16248,N_17141);
and U19359 (N_19359,N_16362,N_17226);
and U19360 (N_19360,N_17363,N_17651);
nand U19361 (N_19361,N_16588,N_16082);
nor U19362 (N_19362,N_16872,N_17456);
nand U19363 (N_19363,N_16046,N_16287);
nand U19364 (N_19364,N_16574,N_16674);
nor U19365 (N_19365,N_17394,N_16841);
xnor U19366 (N_19366,N_17027,N_17757);
xnor U19367 (N_19367,N_17560,N_16680);
xnor U19368 (N_19368,N_16224,N_17564);
or U19369 (N_19369,N_17797,N_17298);
and U19370 (N_19370,N_16269,N_16845);
nor U19371 (N_19371,N_16990,N_17735);
xor U19372 (N_19372,N_16381,N_16319);
nor U19373 (N_19373,N_16144,N_17730);
xnor U19374 (N_19374,N_16734,N_16963);
and U19375 (N_19375,N_17677,N_16057);
nor U19376 (N_19376,N_17707,N_16304);
nand U19377 (N_19377,N_16914,N_17972);
or U19378 (N_19378,N_16849,N_16814);
or U19379 (N_19379,N_16136,N_16085);
or U19380 (N_19380,N_17022,N_16081);
nor U19381 (N_19381,N_17725,N_17395);
or U19382 (N_19382,N_17681,N_17699);
or U19383 (N_19383,N_17227,N_16734);
nand U19384 (N_19384,N_17873,N_16602);
or U19385 (N_19385,N_16693,N_17474);
and U19386 (N_19386,N_17583,N_16029);
nor U19387 (N_19387,N_17652,N_17842);
and U19388 (N_19388,N_17263,N_17768);
and U19389 (N_19389,N_17972,N_17535);
xnor U19390 (N_19390,N_17500,N_16810);
nand U19391 (N_19391,N_16513,N_17803);
nor U19392 (N_19392,N_16433,N_16078);
or U19393 (N_19393,N_17855,N_17186);
xnor U19394 (N_19394,N_16468,N_17947);
or U19395 (N_19395,N_16003,N_17645);
xor U19396 (N_19396,N_16216,N_17666);
nor U19397 (N_19397,N_16106,N_17306);
nor U19398 (N_19398,N_16987,N_17215);
xor U19399 (N_19399,N_16426,N_17246);
xnor U19400 (N_19400,N_17253,N_16707);
nor U19401 (N_19401,N_17067,N_16056);
nor U19402 (N_19402,N_17341,N_17242);
xor U19403 (N_19403,N_16578,N_17568);
nor U19404 (N_19404,N_16162,N_16360);
and U19405 (N_19405,N_17740,N_16303);
or U19406 (N_19406,N_16804,N_17353);
nor U19407 (N_19407,N_16906,N_16787);
nor U19408 (N_19408,N_16547,N_16887);
xor U19409 (N_19409,N_17585,N_16161);
and U19410 (N_19410,N_17985,N_17224);
nor U19411 (N_19411,N_17933,N_17450);
or U19412 (N_19412,N_16739,N_17608);
nor U19413 (N_19413,N_16086,N_17008);
or U19414 (N_19414,N_16140,N_16008);
and U19415 (N_19415,N_16165,N_16208);
nand U19416 (N_19416,N_16494,N_17928);
or U19417 (N_19417,N_17297,N_17216);
and U19418 (N_19418,N_17757,N_17273);
xor U19419 (N_19419,N_17794,N_17428);
or U19420 (N_19420,N_16500,N_17279);
nor U19421 (N_19421,N_16157,N_17309);
nand U19422 (N_19422,N_17033,N_17825);
or U19423 (N_19423,N_17589,N_16429);
xnor U19424 (N_19424,N_17107,N_17054);
or U19425 (N_19425,N_17040,N_16827);
or U19426 (N_19426,N_16276,N_17378);
nand U19427 (N_19427,N_17678,N_17259);
nand U19428 (N_19428,N_16905,N_16019);
and U19429 (N_19429,N_17052,N_16489);
or U19430 (N_19430,N_17614,N_16697);
xnor U19431 (N_19431,N_16680,N_16192);
and U19432 (N_19432,N_17161,N_17070);
nor U19433 (N_19433,N_17783,N_16204);
and U19434 (N_19434,N_17720,N_17407);
and U19435 (N_19435,N_17720,N_17353);
or U19436 (N_19436,N_17279,N_17080);
and U19437 (N_19437,N_17249,N_17021);
or U19438 (N_19438,N_16494,N_16833);
and U19439 (N_19439,N_16318,N_17917);
nand U19440 (N_19440,N_16477,N_16356);
nor U19441 (N_19441,N_17624,N_16676);
nor U19442 (N_19442,N_16608,N_17471);
nor U19443 (N_19443,N_17713,N_16932);
nor U19444 (N_19444,N_16993,N_16697);
xor U19445 (N_19445,N_17889,N_17959);
or U19446 (N_19446,N_16599,N_17277);
nor U19447 (N_19447,N_17808,N_17259);
nand U19448 (N_19448,N_16118,N_17856);
xor U19449 (N_19449,N_17819,N_17001);
nor U19450 (N_19450,N_16426,N_17603);
nand U19451 (N_19451,N_17707,N_17467);
nor U19452 (N_19452,N_17964,N_16762);
xnor U19453 (N_19453,N_16898,N_16705);
nor U19454 (N_19454,N_17038,N_16191);
nand U19455 (N_19455,N_17451,N_16096);
nand U19456 (N_19456,N_16697,N_17739);
xnor U19457 (N_19457,N_17886,N_16863);
or U19458 (N_19458,N_16907,N_16434);
nor U19459 (N_19459,N_16428,N_17510);
or U19460 (N_19460,N_16592,N_16745);
and U19461 (N_19461,N_17975,N_17309);
xnor U19462 (N_19462,N_17474,N_17943);
nor U19463 (N_19463,N_17753,N_17129);
or U19464 (N_19464,N_17367,N_17727);
and U19465 (N_19465,N_16147,N_16074);
nor U19466 (N_19466,N_17768,N_16438);
and U19467 (N_19467,N_16865,N_16122);
or U19468 (N_19468,N_16999,N_16990);
or U19469 (N_19469,N_17624,N_16666);
or U19470 (N_19470,N_17865,N_16061);
or U19471 (N_19471,N_17012,N_16318);
xnor U19472 (N_19472,N_16949,N_16888);
and U19473 (N_19473,N_17922,N_16743);
nand U19474 (N_19474,N_17651,N_17520);
nand U19475 (N_19475,N_16502,N_16032);
or U19476 (N_19476,N_17588,N_16625);
and U19477 (N_19477,N_17643,N_17199);
nand U19478 (N_19478,N_16084,N_16427);
or U19479 (N_19479,N_16736,N_17698);
xnor U19480 (N_19480,N_17596,N_16889);
nand U19481 (N_19481,N_17016,N_17292);
xnor U19482 (N_19482,N_16514,N_16789);
xnor U19483 (N_19483,N_16776,N_17735);
nor U19484 (N_19484,N_16889,N_16220);
nor U19485 (N_19485,N_17924,N_16156);
nor U19486 (N_19486,N_16008,N_16300);
nor U19487 (N_19487,N_16654,N_16594);
or U19488 (N_19488,N_17105,N_16702);
and U19489 (N_19489,N_16639,N_16341);
nor U19490 (N_19490,N_16303,N_16075);
or U19491 (N_19491,N_16487,N_17856);
nor U19492 (N_19492,N_16216,N_17702);
xnor U19493 (N_19493,N_16242,N_17252);
nand U19494 (N_19494,N_17174,N_17435);
xnor U19495 (N_19495,N_17518,N_17164);
nor U19496 (N_19496,N_17552,N_16832);
or U19497 (N_19497,N_16890,N_16791);
xnor U19498 (N_19498,N_17311,N_17422);
xnor U19499 (N_19499,N_17674,N_17209);
xor U19500 (N_19500,N_16505,N_16726);
nand U19501 (N_19501,N_17283,N_16356);
and U19502 (N_19502,N_16600,N_17205);
or U19503 (N_19503,N_16903,N_16399);
and U19504 (N_19504,N_16626,N_17536);
or U19505 (N_19505,N_16045,N_16690);
nand U19506 (N_19506,N_16086,N_17345);
nand U19507 (N_19507,N_17922,N_17794);
nand U19508 (N_19508,N_17669,N_17288);
and U19509 (N_19509,N_16909,N_16599);
and U19510 (N_19510,N_16529,N_16173);
nor U19511 (N_19511,N_17426,N_16195);
nor U19512 (N_19512,N_17904,N_17233);
nor U19513 (N_19513,N_17234,N_17327);
or U19514 (N_19514,N_17230,N_16632);
or U19515 (N_19515,N_17379,N_16155);
nor U19516 (N_19516,N_17080,N_16162);
and U19517 (N_19517,N_16380,N_17337);
xor U19518 (N_19518,N_17860,N_16227);
or U19519 (N_19519,N_17008,N_16851);
or U19520 (N_19520,N_17638,N_16175);
xnor U19521 (N_19521,N_17142,N_17774);
nand U19522 (N_19522,N_16233,N_17453);
xnor U19523 (N_19523,N_16673,N_16971);
nor U19524 (N_19524,N_16895,N_17192);
or U19525 (N_19525,N_16227,N_16914);
nor U19526 (N_19526,N_16479,N_16231);
and U19527 (N_19527,N_16489,N_16595);
nand U19528 (N_19528,N_16256,N_16302);
nor U19529 (N_19529,N_16684,N_17791);
xor U19530 (N_19530,N_17844,N_16732);
xnor U19531 (N_19531,N_17607,N_17722);
xor U19532 (N_19532,N_16905,N_17663);
nand U19533 (N_19533,N_17915,N_16799);
and U19534 (N_19534,N_17626,N_17872);
nand U19535 (N_19535,N_17130,N_16827);
nand U19536 (N_19536,N_16806,N_17321);
and U19537 (N_19537,N_17676,N_17804);
or U19538 (N_19538,N_17213,N_16075);
nor U19539 (N_19539,N_16764,N_17044);
nand U19540 (N_19540,N_17388,N_17900);
xnor U19541 (N_19541,N_17324,N_17303);
xor U19542 (N_19542,N_16570,N_16378);
and U19543 (N_19543,N_17903,N_16690);
and U19544 (N_19544,N_16996,N_17704);
xnor U19545 (N_19545,N_17175,N_16747);
nand U19546 (N_19546,N_17426,N_16385);
and U19547 (N_19547,N_16941,N_17156);
and U19548 (N_19548,N_16083,N_17783);
and U19549 (N_19549,N_17762,N_16337);
nand U19550 (N_19550,N_17679,N_16712);
or U19551 (N_19551,N_17883,N_17138);
nand U19552 (N_19552,N_17674,N_17504);
nand U19553 (N_19553,N_16472,N_16823);
xor U19554 (N_19554,N_16645,N_16789);
and U19555 (N_19555,N_17719,N_17604);
nand U19556 (N_19556,N_17816,N_16702);
nand U19557 (N_19557,N_17440,N_16803);
xor U19558 (N_19558,N_16843,N_17371);
nand U19559 (N_19559,N_17736,N_16152);
xor U19560 (N_19560,N_16494,N_17893);
and U19561 (N_19561,N_16535,N_17419);
nand U19562 (N_19562,N_16731,N_16816);
xor U19563 (N_19563,N_17446,N_16472);
or U19564 (N_19564,N_16587,N_16138);
or U19565 (N_19565,N_16254,N_16474);
nand U19566 (N_19566,N_17396,N_16054);
or U19567 (N_19567,N_16161,N_17940);
xnor U19568 (N_19568,N_16227,N_17612);
xnor U19569 (N_19569,N_17983,N_17733);
nor U19570 (N_19570,N_16689,N_16678);
nand U19571 (N_19571,N_17421,N_16903);
and U19572 (N_19572,N_17677,N_16190);
and U19573 (N_19573,N_16528,N_16288);
and U19574 (N_19574,N_16833,N_16013);
xnor U19575 (N_19575,N_16108,N_16750);
or U19576 (N_19576,N_16016,N_17058);
or U19577 (N_19577,N_17575,N_16709);
nand U19578 (N_19578,N_16391,N_16397);
and U19579 (N_19579,N_16976,N_17179);
or U19580 (N_19580,N_17386,N_17040);
and U19581 (N_19581,N_16634,N_17172);
xnor U19582 (N_19582,N_16997,N_17861);
xor U19583 (N_19583,N_16489,N_16658);
xnor U19584 (N_19584,N_16380,N_16819);
nand U19585 (N_19585,N_16762,N_17665);
xor U19586 (N_19586,N_17362,N_17335);
or U19587 (N_19587,N_17893,N_16469);
and U19588 (N_19588,N_16184,N_16335);
xnor U19589 (N_19589,N_17424,N_17929);
nor U19590 (N_19590,N_16718,N_16928);
or U19591 (N_19591,N_16122,N_17671);
nor U19592 (N_19592,N_16389,N_17194);
xor U19593 (N_19593,N_17628,N_16028);
xnor U19594 (N_19594,N_16580,N_17919);
or U19595 (N_19595,N_17388,N_16415);
and U19596 (N_19596,N_16219,N_16374);
nand U19597 (N_19597,N_17263,N_16623);
xor U19598 (N_19598,N_16612,N_16199);
xor U19599 (N_19599,N_16861,N_16049);
and U19600 (N_19600,N_16789,N_16796);
nand U19601 (N_19601,N_17227,N_17861);
or U19602 (N_19602,N_17676,N_17880);
and U19603 (N_19603,N_17954,N_16063);
or U19604 (N_19604,N_17976,N_17630);
nand U19605 (N_19605,N_17498,N_17318);
nand U19606 (N_19606,N_17113,N_17023);
nand U19607 (N_19607,N_17682,N_16669);
or U19608 (N_19608,N_17660,N_17990);
nand U19609 (N_19609,N_16236,N_17083);
and U19610 (N_19610,N_17925,N_17946);
nor U19611 (N_19611,N_17379,N_16393);
and U19612 (N_19612,N_16245,N_16361);
nor U19613 (N_19613,N_17667,N_17806);
xnor U19614 (N_19614,N_16568,N_17358);
nand U19615 (N_19615,N_16367,N_16805);
xnor U19616 (N_19616,N_17497,N_16452);
and U19617 (N_19617,N_16900,N_17806);
nor U19618 (N_19618,N_17384,N_16466);
nor U19619 (N_19619,N_17718,N_17508);
nor U19620 (N_19620,N_17177,N_16736);
nor U19621 (N_19621,N_16267,N_17044);
or U19622 (N_19622,N_17028,N_16584);
xor U19623 (N_19623,N_17449,N_16434);
xnor U19624 (N_19624,N_16704,N_17211);
nand U19625 (N_19625,N_17692,N_17615);
nor U19626 (N_19626,N_16049,N_17903);
xor U19627 (N_19627,N_17853,N_16503);
nand U19628 (N_19628,N_16358,N_17541);
nor U19629 (N_19629,N_17561,N_17287);
nor U19630 (N_19630,N_17315,N_16146);
xor U19631 (N_19631,N_17947,N_17588);
nor U19632 (N_19632,N_17637,N_16022);
or U19633 (N_19633,N_17901,N_17858);
nor U19634 (N_19634,N_16752,N_16463);
and U19635 (N_19635,N_17352,N_16617);
and U19636 (N_19636,N_17200,N_16897);
nor U19637 (N_19637,N_16567,N_17947);
nor U19638 (N_19638,N_16108,N_17758);
nor U19639 (N_19639,N_16587,N_16998);
xnor U19640 (N_19640,N_17294,N_17820);
nand U19641 (N_19641,N_17176,N_17230);
and U19642 (N_19642,N_16497,N_16434);
nor U19643 (N_19643,N_16724,N_16957);
nand U19644 (N_19644,N_17932,N_17515);
nand U19645 (N_19645,N_17064,N_16228);
xnor U19646 (N_19646,N_16621,N_16956);
or U19647 (N_19647,N_16248,N_17717);
or U19648 (N_19648,N_17779,N_16413);
nand U19649 (N_19649,N_17036,N_17427);
or U19650 (N_19650,N_17432,N_17812);
xnor U19651 (N_19651,N_16919,N_16355);
or U19652 (N_19652,N_16010,N_16729);
or U19653 (N_19653,N_16386,N_17436);
xor U19654 (N_19654,N_16779,N_17995);
xnor U19655 (N_19655,N_17522,N_17616);
xnor U19656 (N_19656,N_17011,N_16484);
nand U19657 (N_19657,N_16796,N_17066);
and U19658 (N_19658,N_17196,N_16616);
nor U19659 (N_19659,N_17725,N_16186);
xor U19660 (N_19660,N_17391,N_17269);
xnor U19661 (N_19661,N_16965,N_16533);
or U19662 (N_19662,N_17660,N_17306);
nor U19663 (N_19663,N_17651,N_16119);
xnor U19664 (N_19664,N_16109,N_16025);
nand U19665 (N_19665,N_16994,N_17852);
nor U19666 (N_19666,N_16465,N_16051);
and U19667 (N_19667,N_17454,N_17324);
or U19668 (N_19668,N_17768,N_17083);
xnor U19669 (N_19669,N_17569,N_17836);
xor U19670 (N_19670,N_17095,N_17179);
xnor U19671 (N_19671,N_17893,N_17888);
nand U19672 (N_19672,N_17311,N_16739);
nand U19673 (N_19673,N_17799,N_16135);
xnor U19674 (N_19674,N_17871,N_16863);
nor U19675 (N_19675,N_17073,N_17339);
nor U19676 (N_19676,N_17737,N_17293);
or U19677 (N_19677,N_16510,N_16727);
nor U19678 (N_19678,N_17714,N_16987);
or U19679 (N_19679,N_17279,N_16952);
nor U19680 (N_19680,N_17118,N_17951);
nor U19681 (N_19681,N_16597,N_17794);
nand U19682 (N_19682,N_17699,N_16538);
or U19683 (N_19683,N_16273,N_16329);
and U19684 (N_19684,N_17045,N_16968);
or U19685 (N_19685,N_16928,N_16092);
nor U19686 (N_19686,N_16893,N_16708);
or U19687 (N_19687,N_17407,N_16202);
nand U19688 (N_19688,N_17368,N_17662);
and U19689 (N_19689,N_16911,N_16743);
and U19690 (N_19690,N_17322,N_16043);
xnor U19691 (N_19691,N_17800,N_16954);
xor U19692 (N_19692,N_17220,N_16123);
or U19693 (N_19693,N_17900,N_17190);
and U19694 (N_19694,N_17385,N_16065);
or U19695 (N_19695,N_16990,N_17011);
nand U19696 (N_19696,N_16016,N_17853);
nand U19697 (N_19697,N_16787,N_17183);
xor U19698 (N_19698,N_17856,N_16437);
xor U19699 (N_19699,N_16129,N_16397);
xor U19700 (N_19700,N_17877,N_16492);
nor U19701 (N_19701,N_17894,N_16709);
or U19702 (N_19702,N_17149,N_17578);
nor U19703 (N_19703,N_16720,N_17537);
xnor U19704 (N_19704,N_17960,N_17364);
nand U19705 (N_19705,N_16362,N_17032);
xnor U19706 (N_19706,N_17767,N_17750);
or U19707 (N_19707,N_16902,N_17765);
and U19708 (N_19708,N_16383,N_16682);
nand U19709 (N_19709,N_16308,N_17631);
xor U19710 (N_19710,N_16646,N_17702);
xnor U19711 (N_19711,N_16358,N_17356);
and U19712 (N_19712,N_17339,N_17609);
and U19713 (N_19713,N_17237,N_17047);
nor U19714 (N_19714,N_16774,N_16755);
nand U19715 (N_19715,N_17529,N_17023);
nand U19716 (N_19716,N_16205,N_17794);
or U19717 (N_19717,N_17370,N_17989);
or U19718 (N_19718,N_16350,N_17498);
nor U19719 (N_19719,N_16002,N_17851);
nor U19720 (N_19720,N_17914,N_17473);
xnor U19721 (N_19721,N_17974,N_16794);
and U19722 (N_19722,N_16704,N_16978);
nor U19723 (N_19723,N_16021,N_17465);
and U19724 (N_19724,N_17503,N_16064);
nand U19725 (N_19725,N_17062,N_16805);
nor U19726 (N_19726,N_17311,N_16909);
or U19727 (N_19727,N_17887,N_16991);
and U19728 (N_19728,N_16289,N_17747);
nor U19729 (N_19729,N_16156,N_16107);
or U19730 (N_19730,N_17551,N_16202);
xnor U19731 (N_19731,N_17678,N_16002);
and U19732 (N_19732,N_17218,N_17156);
nor U19733 (N_19733,N_16376,N_17098);
or U19734 (N_19734,N_17340,N_17426);
xor U19735 (N_19735,N_16431,N_16125);
or U19736 (N_19736,N_16453,N_16396);
and U19737 (N_19737,N_17080,N_17223);
or U19738 (N_19738,N_17753,N_16808);
nor U19739 (N_19739,N_17220,N_17554);
and U19740 (N_19740,N_17513,N_17025);
or U19741 (N_19741,N_17725,N_16462);
or U19742 (N_19742,N_17779,N_16033);
and U19743 (N_19743,N_17707,N_17681);
and U19744 (N_19744,N_17128,N_16933);
or U19745 (N_19745,N_16007,N_17973);
nor U19746 (N_19746,N_17003,N_16446);
nand U19747 (N_19747,N_16861,N_17081);
and U19748 (N_19748,N_17029,N_17533);
xor U19749 (N_19749,N_16748,N_17576);
nand U19750 (N_19750,N_17200,N_16512);
nand U19751 (N_19751,N_16646,N_17809);
xnor U19752 (N_19752,N_16920,N_16698);
nand U19753 (N_19753,N_16971,N_16891);
or U19754 (N_19754,N_17492,N_17932);
xnor U19755 (N_19755,N_17599,N_16688);
nor U19756 (N_19756,N_16855,N_16280);
nor U19757 (N_19757,N_17830,N_17874);
and U19758 (N_19758,N_17126,N_16248);
nand U19759 (N_19759,N_17892,N_17987);
or U19760 (N_19760,N_16486,N_16065);
nand U19761 (N_19761,N_16382,N_17903);
xnor U19762 (N_19762,N_16949,N_16234);
nor U19763 (N_19763,N_16552,N_17014);
xnor U19764 (N_19764,N_16843,N_17054);
or U19765 (N_19765,N_17810,N_17403);
nor U19766 (N_19766,N_17235,N_17988);
nor U19767 (N_19767,N_16986,N_17691);
or U19768 (N_19768,N_16623,N_17663);
or U19769 (N_19769,N_16603,N_16133);
xor U19770 (N_19770,N_16199,N_16913);
nand U19771 (N_19771,N_16862,N_17745);
and U19772 (N_19772,N_16822,N_17187);
nor U19773 (N_19773,N_17551,N_16930);
xor U19774 (N_19774,N_17064,N_16160);
nor U19775 (N_19775,N_17605,N_16571);
nor U19776 (N_19776,N_17006,N_16794);
and U19777 (N_19777,N_17185,N_16237);
nand U19778 (N_19778,N_17154,N_17310);
nand U19779 (N_19779,N_16045,N_17489);
xor U19780 (N_19780,N_17203,N_17362);
nor U19781 (N_19781,N_16865,N_16006);
nand U19782 (N_19782,N_16506,N_16984);
xor U19783 (N_19783,N_16863,N_17203);
nand U19784 (N_19784,N_17500,N_16529);
nor U19785 (N_19785,N_16731,N_17159);
nor U19786 (N_19786,N_16628,N_17361);
nor U19787 (N_19787,N_16038,N_16519);
and U19788 (N_19788,N_17714,N_17880);
nand U19789 (N_19789,N_16202,N_16092);
or U19790 (N_19790,N_17076,N_16488);
xor U19791 (N_19791,N_17462,N_16459);
nor U19792 (N_19792,N_17585,N_16828);
nor U19793 (N_19793,N_17861,N_16830);
nand U19794 (N_19794,N_17035,N_17191);
nor U19795 (N_19795,N_16024,N_16399);
or U19796 (N_19796,N_17188,N_17760);
and U19797 (N_19797,N_17837,N_16746);
and U19798 (N_19798,N_17459,N_16873);
or U19799 (N_19799,N_16646,N_16757);
nor U19800 (N_19800,N_17635,N_17510);
nor U19801 (N_19801,N_16466,N_17364);
nand U19802 (N_19802,N_16986,N_17179);
and U19803 (N_19803,N_16785,N_16714);
and U19804 (N_19804,N_17870,N_16546);
and U19805 (N_19805,N_16907,N_16873);
nor U19806 (N_19806,N_17198,N_16895);
nor U19807 (N_19807,N_17299,N_17153);
xnor U19808 (N_19808,N_17240,N_16154);
nor U19809 (N_19809,N_17430,N_16105);
and U19810 (N_19810,N_16361,N_16413);
or U19811 (N_19811,N_16573,N_17395);
nor U19812 (N_19812,N_16039,N_17421);
nor U19813 (N_19813,N_16567,N_17277);
or U19814 (N_19814,N_17795,N_16023);
and U19815 (N_19815,N_17907,N_16955);
or U19816 (N_19816,N_17269,N_16768);
and U19817 (N_19817,N_16522,N_17535);
or U19818 (N_19818,N_16465,N_16425);
nor U19819 (N_19819,N_17705,N_17499);
nand U19820 (N_19820,N_16352,N_17300);
or U19821 (N_19821,N_17499,N_17949);
or U19822 (N_19822,N_16982,N_17934);
or U19823 (N_19823,N_17885,N_16813);
and U19824 (N_19824,N_16237,N_16303);
xor U19825 (N_19825,N_16002,N_16783);
nor U19826 (N_19826,N_17271,N_16679);
xor U19827 (N_19827,N_17128,N_17420);
and U19828 (N_19828,N_17230,N_16337);
and U19829 (N_19829,N_16768,N_16966);
nor U19830 (N_19830,N_16519,N_17450);
nand U19831 (N_19831,N_16291,N_17541);
nor U19832 (N_19832,N_16016,N_16356);
nand U19833 (N_19833,N_16093,N_17676);
and U19834 (N_19834,N_17009,N_17771);
nor U19835 (N_19835,N_16359,N_16774);
xor U19836 (N_19836,N_17497,N_16920);
nand U19837 (N_19837,N_17583,N_16364);
or U19838 (N_19838,N_16190,N_17171);
nor U19839 (N_19839,N_16984,N_16747);
and U19840 (N_19840,N_16716,N_16352);
nor U19841 (N_19841,N_16466,N_16046);
nor U19842 (N_19842,N_16418,N_16321);
nor U19843 (N_19843,N_16001,N_16041);
nor U19844 (N_19844,N_17558,N_17457);
nand U19845 (N_19845,N_17550,N_16616);
nand U19846 (N_19846,N_16383,N_17411);
and U19847 (N_19847,N_17914,N_17794);
xor U19848 (N_19848,N_16622,N_16569);
or U19849 (N_19849,N_16413,N_16173);
or U19850 (N_19850,N_17656,N_17951);
nor U19851 (N_19851,N_16008,N_16479);
nor U19852 (N_19852,N_17660,N_17744);
or U19853 (N_19853,N_16388,N_16293);
and U19854 (N_19854,N_17696,N_17312);
or U19855 (N_19855,N_16534,N_16054);
xnor U19856 (N_19856,N_16549,N_16985);
or U19857 (N_19857,N_16437,N_16179);
xor U19858 (N_19858,N_16117,N_16114);
or U19859 (N_19859,N_17634,N_16737);
nand U19860 (N_19860,N_17598,N_16417);
nor U19861 (N_19861,N_17367,N_16115);
or U19862 (N_19862,N_16137,N_17267);
or U19863 (N_19863,N_17220,N_17869);
and U19864 (N_19864,N_16430,N_16046);
and U19865 (N_19865,N_17006,N_16698);
nand U19866 (N_19866,N_16147,N_17644);
or U19867 (N_19867,N_16664,N_17298);
nor U19868 (N_19868,N_17575,N_17332);
or U19869 (N_19869,N_17717,N_16752);
and U19870 (N_19870,N_17016,N_16946);
and U19871 (N_19871,N_17595,N_16164);
xnor U19872 (N_19872,N_17428,N_17455);
xor U19873 (N_19873,N_16336,N_16213);
and U19874 (N_19874,N_17022,N_17090);
nor U19875 (N_19875,N_17629,N_16150);
nor U19876 (N_19876,N_17395,N_17412);
nor U19877 (N_19877,N_17229,N_16800);
nand U19878 (N_19878,N_16290,N_17307);
nor U19879 (N_19879,N_16210,N_16797);
nor U19880 (N_19880,N_16112,N_16191);
xnor U19881 (N_19881,N_17112,N_16050);
or U19882 (N_19882,N_16587,N_17220);
xnor U19883 (N_19883,N_17251,N_16836);
xnor U19884 (N_19884,N_16700,N_16945);
and U19885 (N_19885,N_16964,N_17370);
or U19886 (N_19886,N_17057,N_16188);
nand U19887 (N_19887,N_16176,N_16632);
or U19888 (N_19888,N_17403,N_16880);
and U19889 (N_19889,N_17228,N_16454);
xor U19890 (N_19890,N_17483,N_16185);
xor U19891 (N_19891,N_17176,N_17079);
nand U19892 (N_19892,N_16095,N_17043);
xnor U19893 (N_19893,N_16209,N_17564);
nor U19894 (N_19894,N_16210,N_17118);
nand U19895 (N_19895,N_16767,N_17976);
nand U19896 (N_19896,N_17467,N_16890);
nand U19897 (N_19897,N_17398,N_16628);
and U19898 (N_19898,N_16639,N_17891);
nor U19899 (N_19899,N_16555,N_17761);
nor U19900 (N_19900,N_17283,N_16031);
nand U19901 (N_19901,N_17504,N_17886);
nand U19902 (N_19902,N_17593,N_17812);
or U19903 (N_19903,N_16714,N_17944);
xor U19904 (N_19904,N_17870,N_17409);
xnor U19905 (N_19905,N_17232,N_17192);
nor U19906 (N_19906,N_17761,N_17821);
nand U19907 (N_19907,N_16023,N_17144);
nand U19908 (N_19908,N_16277,N_17057);
xnor U19909 (N_19909,N_16506,N_17903);
nor U19910 (N_19910,N_17259,N_16133);
and U19911 (N_19911,N_17922,N_16921);
nand U19912 (N_19912,N_16946,N_17320);
xor U19913 (N_19913,N_17555,N_16923);
and U19914 (N_19914,N_16654,N_16344);
and U19915 (N_19915,N_16873,N_16177);
xor U19916 (N_19916,N_17347,N_17930);
and U19917 (N_19917,N_16775,N_17521);
and U19918 (N_19918,N_16018,N_16859);
and U19919 (N_19919,N_17699,N_17515);
xor U19920 (N_19920,N_17722,N_16441);
xnor U19921 (N_19921,N_16308,N_17633);
or U19922 (N_19922,N_17263,N_16841);
or U19923 (N_19923,N_16410,N_17385);
and U19924 (N_19924,N_17103,N_17901);
or U19925 (N_19925,N_16936,N_17530);
or U19926 (N_19926,N_16201,N_16394);
or U19927 (N_19927,N_17607,N_16238);
or U19928 (N_19928,N_17022,N_16248);
nand U19929 (N_19929,N_17023,N_16187);
or U19930 (N_19930,N_17408,N_17028);
nand U19931 (N_19931,N_17287,N_16236);
or U19932 (N_19932,N_17939,N_16615);
nand U19933 (N_19933,N_16472,N_17473);
and U19934 (N_19934,N_16854,N_17574);
or U19935 (N_19935,N_17431,N_17476);
or U19936 (N_19936,N_16068,N_16324);
or U19937 (N_19937,N_16662,N_16730);
or U19938 (N_19938,N_17069,N_17135);
or U19939 (N_19939,N_16312,N_17994);
and U19940 (N_19940,N_17138,N_17232);
nor U19941 (N_19941,N_17257,N_17046);
xor U19942 (N_19942,N_16475,N_17213);
nor U19943 (N_19943,N_16583,N_17337);
nand U19944 (N_19944,N_17774,N_17677);
xnor U19945 (N_19945,N_16862,N_17668);
or U19946 (N_19946,N_17956,N_16714);
or U19947 (N_19947,N_16337,N_16264);
nor U19948 (N_19948,N_16415,N_16863);
nor U19949 (N_19949,N_16051,N_17521);
and U19950 (N_19950,N_17057,N_17045);
nor U19951 (N_19951,N_17940,N_16545);
and U19952 (N_19952,N_17269,N_17972);
xor U19953 (N_19953,N_17261,N_17875);
nor U19954 (N_19954,N_16475,N_17190);
and U19955 (N_19955,N_16455,N_17549);
nand U19956 (N_19956,N_17467,N_17223);
nor U19957 (N_19957,N_16901,N_16323);
nor U19958 (N_19958,N_16289,N_16862);
nand U19959 (N_19959,N_16934,N_17371);
xnor U19960 (N_19960,N_17096,N_17015);
nor U19961 (N_19961,N_16759,N_16112);
xor U19962 (N_19962,N_17341,N_17948);
or U19963 (N_19963,N_17848,N_16483);
nor U19964 (N_19964,N_16544,N_17309);
nor U19965 (N_19965,N_17722,N_16538);
and U19966 (N_19966,N_16118,N_17772);
xor U19967 (N_19967,N_16928,N_17217);
and U19968 (N_19968,N_17107,N_16195);
nor U19969 (N_19969,N_17323,N_16049);
xnor U19970 (N_19970,N_16384,N_16901);
xor U19971 (N_19971,N_17491,N_17946);
xnor U19972 (N_19972,N_16126,N_16253);
nor U19973 (N_19973,N_17452,N_17377);
nor U19974 (N_19974,N_16035,N_16788);
or U19975 (N_19975,N_16076,N_16480);
nor U19976 (N_19976,N_17076,N_17777);
nand U19977 (N_19977,N_16115,N_17479);
or U19978 (N_19978,N_17496,N_16204);
or U19979 (N_19979,N_16864,N_17932);
and U19980 (N_19980,N_17725,N_17430);
nand U19981 (N_19981,N_16916,N_16373);
or U19982 (N_19982,N_16767,N_16386);
xor U19983 (N_19983,N_16453,N_17314);
nor U19984 (N_19984,N_17576,N_16247);
and U19985 (N_19985,N_16938,N_17134);
nand U19986 (N_19986,N_17492,N_17162);
or U19987 (N_19987,N_16308,N_17336);
or U19988 (N_19988,N_17222,N_16194);
or U19989 (N_19989,N_16733,N_16403);
xnor U19990 (N_19990,N_16154,N_17132);
nand U19991 (N_19991,N_16383,N_16937);
or U19992 (N_19992,N_17140,N_17968);
nand U19993 (N_19993,N_17612,N_16796);
and U19994 (N_19994,N_16710,N_16377);
nand U19995 (N_19995,N_16967,N_16893);
nand U19996 (N_19996,N_16513,N_16220);
xor U19997 (N_19997,N_17316,N_17631);
xnor U19998 (N_19998,N_16835,N_16883);
or U19999 (N_19999,N_17664,N_17456);
or UO_0 (O_0,N_18512,N_19174);
xnor UO_1 (O_1,N_18518,N_18077);
xnor UO_2 (O_2,N_18069,N_18705);
or UO_3 (O_3,N_19592,N_18453);
or UO_4 (O_4,N_18676,N_18403);
xor UO_5 (O_5,N_18855,N_18333);
xor UO_6 (O_6,N_19333,N_19080);
or UO_7 (O_7,N_19771,N_18416);
and UO_8 (O_8,N_18735,N_18529);
or UO_9 (O_9,N_18953,N_19320);
nor UO_10 (O_10,N_19444,N_19210);
and UO_11 (O_11,N_18085,N_19015);
xor UO_12 (O_12,N_18547,N_18960);
xnor UO_13 (O_13,N_18107,N_19537);
xor UO_14 (O_14,N_18183,N_19449);
and UO_15 (O_15,N_19119,N_19969);
xor UO_16 (O_16,N_18126,N_18563);
and UO_17 (O_17,N_18831,N_18010);
nand UO_18 (O_18,N_18712,N_19675);
and UO_19 (O_19,N_18003,N_18995);
or UO_20 (O_20,N_18498,N_18906);
nor UO_21 (O_21,N_18974,N_19654);
nand UO_22 (O_22,N_18141,N_19062);
and UO_23 (O_23,N_19912,N_19175);
and UO_24 (O_24,N_19861,N_19408);
nor UO_25 (O_25,N_19138,N_19763);
nand UO_26 (O_26,N_18905,N_18310);
and UO_27 (O_27,N_19284,N_18420);
or UO_28 (O_28,N_19042,N_18427);
nor UO_29 (O_29,N_18804,N_18426);
nand UO_30 (O_30,N_19837,N_18463);
and UO_31 (O_31,N_18955,N_19577);
nand UO_32 (O_32,N_18577,N_18760);
xor UO_33 (O_33,N_19456,N_18368);
xnor UO_34 (O_34,N_19113,N_19635);
nand UO_35 (O_35,N_18461,N_19129);
or UO_36 (O_36,N_18283,N_18023);
or UO_37 (O_37,N_19224,N_18894);
nand UO_38 (O_38,N_19669,N_19937);
xnor UO_39 (O_39,N_18241,N_19968);
and UO_40 (O_40,N_18424,N_18312);
nand UO_41 (O_41,N_19241,N_19493);
and UO_42 (O_42,N_18820,N_18800);
or UO_43 (O_43,N_19511,N_18353);
nand UO_44 (O_44,N_18150,N_18391);
nand UO_45 (O_45,N_18487,N_18553);
and UO_46 (O_46,N_18966,N_19013);
xnor UO_47 (O_47,N_18765,N_18914);
or UO_48 (O_48,N_19617,N_19327);
and UO_49 (O_49,N_19069,N_19889);
nand UO_50 (O_50,N_19691,N_19016);
xnor UO_51 (O_51,N_19351,N_19405);
and UO_52 (O_52,N_18789,N_19848);
or UO_53 (O_53,N_18798,N_18674);
nand UO_54 (O_54,N_18051,N_18394);
and UO_55 (O_55,N_19613,N_18342);
or UO_56 (O_56,N_19289,N_19481);
nand UO_57 (O_57,N_18637,N_19440);
xnor UO_58 (O_58,N_19860,N_19501);
and UO_59 (O_59,N_18387,N_19980);
nand UO_60 (O_60,N_18411,N_19921);
nand UO_61 (O_61,N_18635,N_19244);
nor UO_62 (O_62,N_19803,N_19801);
and UO_63 (O_63,N_19077,N_19994);
or UO_64 (O_64,N_19250,N_18042);
xor UO_65 (O_65,N_18471,N_19634);
or UO_66 (O_66,N_18136,N_19468);
or UO_67 (O_67,N_19382,N_19088);
nand UO_68 (O_68,N_19349,N_18532);
nor UO_69 (O_69,N_18555,N_19979);
and UO_70 (O_70,N_19923,N_19472);
or UO_71 (O_71,N_18599,N_18025);
or UO_72 (O_72,N_18358,N_18790);
and UO_73 (O_73,N_19671,N_19575);
or UO_74 (O_74,N_18928,N_19084);
and UO_75 (O_75,N_18040,N_19659);
and UO_76 (O_76,N_18679,N_19693);
and UO_77 (O_77,N_18337,N_19786);
or UO_78 (O_78,N_19153,N_19064);
nor UO_79 (O_79,N_18846,N_19115);
nand UO_80 (O_80,N_18445,N_19461);
nor UO_81 (O_81,N_18719,N_18489);
nor UO_82 (O_82,N_19962,N_19909);
nor UO_83 (O_83,N_19829,N_18805);
and UO_84 (O_84,N_19546,N_18548);
or UO_85 (O_85,N_18525,N_18541);
nand UO_86 (O_86,N_19309,N_19341);
and UO_87 (O_87,N_18724,N_18224);
nor UO_88 (O_88,N_18610,N_19977);
nand UO_89 (O_89,N_19974,N_19616);
nand UO_90 (O_90,N_19729,N_18474);
nand UO_91 (O_91,N_19010,N_19933);
or UO_92 (O_92,N_19802,N_19806);
or UO_93 (O_93,N_18048,N_18441);
nand UO_94 (O_94,N_18177,N_18649);
and UO_95 (O_95,N_19218,N_19116);
and UO_96 (O_96,N_19462,N_19820);
nand UO_97 (O_97,N_19499,N_18259);
xnor UO_98 (O_98,N_19151,N_19096);
nor UO_99 (O_99,N_19211,N_19401);
nor UO_100 (O_100,N_19756,N_18089);
xor UO_101 (O_101,N_19283,N_19240);
nand UO_102 (O_102,N_19025,N_19543);
nand UO_103 (O_103,N_19039,N_19878);
xnor UO_104 (O_104,N_19652,N_19960);
and UO_105 (O_105,N_19989,N_19325);
or UO_106 (O_106,N_19280,N_19790);
or UO_107 (O_107,N_18339,N_19818);
nand UO_108 (O_108,N_18513,N_18491);
or UO_109 (O_109,N_18982,N_19152);
nand UO_110 (O_110,N_18728,N_18866);
nor UO_111 (O_111,N_18060,N_19559);
nand UO_112 (O_112,N_18037,N_19387);
nand UO_113 (O_113,N_19752,N_18059);
nand UO_114 (O_114,N_18315,N_18115);
and UO_115 (O_115,N_18552,N_19736);
nand UO_116 (O_116,N_19413,N_18422);
xnor UO_117 (O_117,N_18576,N_18625);
and UO_118 (O_118,N_19530,N_18002);
nand UO_119 (O_119,N_18933,N_18351);
or UO_120 (O_120,N_18757,N_19102);
nand UO_121 (O_121,N_18496,N_19161);
or UO_122 (O_122,N_18980,N_19256);
or UO_123 (O_123,N_19058,N_19198);
or UO_124 (O_124,N_18912,N_18488);
or UO_125 (O_125,N_19604,N_18981);
xor UO_126 (O_126,N_18361,N_18954);
xor UO_127 (O_127,N_19593,N_18773);
or UO_128 (O_128,N_19620,N_19164);
xor UO_129 (O_129,N_18021,N_18247);
nand UO_130 (O_130,N_18444,N_19585);
nor UO_131 (O_131,N_18694,N_19538);
and UO_132 (O_132,N_18633,N_19590);
and UO_133 (O_133,N_18066,N_18588);
nand UO_134 (O_134,N_19451,N_19354);
and UO_135 (O_135,N_18882,N_19840);
and UO_136 (O_136,N_18043,N_19380);
nor UO_137 (O_137,N_19730,N_19733);
nand UO_138 (O_138,N_18780,N_18997);
nand UO_139 (O_139,N_18516,N_18743);
xnor UO_140 (O_140,N_18460,N_18213);
or UO_141 (O_141,N_18963,N_18880);
or UO_142 (O_142,N_18546,N_19513);
and UO_143 (O_143,N_18330,N_18891);
xor UO_144 (O_144,N_19514,N_18328);
nor UO_145 (O_145,N_18139,N_19184);
or UO_146 (O_146,N_19334,N_19862);
nand UO_147 (O_147,N_18636,N_19685);
and UO_148 (O_148,N_19090,N_18989);
nand UO_149 (O_149,N_19448,N_18840);
xor UO_150 (O_150,N_18589,N_19337);
nor UO_151 (O_151,N_18772,N_18785);
and UO_152 (O_152,N_19353,N_18381);
nand UO_153 (O_153,N_18559,N_19477);
nand UO_154 (O_154,N_19655,N_19781);
nand UO_155 (O_155,N_18159,N_19540);
and UO_156 (O_156,N_18155,N_18892);
and UO_157 (O_157,N_18691,N_18638);
and UO_158 (O_158,N_18741,N_18562);
nand UO_159 (O_159,N_18039,N_19163);
and UO_160 (O_160,N_18688,N_19021);
nand UO_161 (O_161,N_19965,N_18389);
or UO_162 (O_162,N_18202,N_19237);
nand UO_163 (O_163,N_19485,N_19875);
or UO_164 (O_164,N_19971,N_18192);
nand UO_165 (O_165,N_18402,N_19883);
or UO_166 (O_166,N_18868,N_18369);
nor UO_167 (O_167,N_19052,N_19067);
and UO_168 (O_168,N_18669,N_18404);
xor UO_169 (O_169,N_19074,N_18697);
or UO_170 (O_170,N_18538,N_19529);
xor UO_171 (O_171,N_19302,N_19916);
and UO_172 (O_172,N_18132,N_19087);
nor UO_173 (O_173,N_18539,N_19442);
or UO_174 (O_174,N_19640,N_18475);
xor UO_175 (O_175,N_18707,N_18469);
or UO_176 (O_176,N_18639,N_18074);
xor UO_177 (O_177,N_19199,N_18657);
xnor UO_178 (O_178,N_18194,N_19745);
and UO_179 (O_179,N_19951,N_18750);
and UO_180 (O_180,N_18929,N_18448);
or UO_181 (O_181,N_18684,N_18350);
nand UO_182 (O_182,N_19101,N_18414);
nand UO_183 (O_183,N_18581,N_18032);
nand UO_184 (O_184,N_18985,N_18284);
xor UO_185 (O_185,N_18845,N_19043);
nand UO_186 (O_186,N_18614,N_19407);
or UO_187 (O_187,N_19926,N_19457);
and UO_188 (O_188,N_19759,N_19255);
nand UO_189 (O_189,N_18147,N_19890);
nor UO_190 (O_190,N_18013,N_18797);
nor UO_191 (O_191,N_19484,N_19411);
nor UO_192 (O_192,N_19683,N_18045);
nand UO_193 (O_193,N_18366,N_19145);
nor UO_194 (O_194,N_18044,N_19421);
nand UO_195 (O_195,N_18062,N_19928);
or UO_196 (O_196,N_19191,N_18245);
xnor UO_197 (O_197,N_19336,N_18112);
nor UO_198 (O_198,N_18129,N_18844);
nor UO_199 (O_199,N_19506,N_18731);
or UO_200 (O_200,N_19120,N_19812);
and UO_201 (O_201,N_19929,N_18768);
nor UO_202 (O_202,N_18909,N_18854);
nand UO_203 (O_203,N_19375,N_19497);
xnor UO_204 (O_204,N_18087,N_18314);
nor UO_205 (O_205,N_19697,N_19223);
xnor UO_206 (O_206,N_19667,N_18097);
nor UO_207 (O_207,N_19012,N_19473);
nor UO_208 (O_208,N_19033,N_19170);
and UO_209 (O_209,N_18720,N_19983);
nor UO_210 (O_210,N_18571,N_19699);
and UO_211 (O_211,N_18747,N_19855);
nand UO_212 (O_212,N_19570,N_19315);
xor UO_213 (O_213,N_18158,N_18695);
nor UO_214 (O_214,N_18961,N_18199);
xnor UO_215 (O_215,N_18447,N_18430);
or UO_216 (O_216,N_18945,N_19135);
and UO_217 (O_217,N_18681,N_19075);
nor UO_218 (O_218,N_18716,N_19376);
xnor UO_219 (O_219,N_18825,N_19880);
or UO_220 (O_220,N_19679,N_18675);
xor UO_221 (O_221,N_18534,N_18265);
xor UO_222 (O_222,N_18907,N_19272);
nor UO_223 (O_223,N_18286,N_18551);
nor UO_224 (O_224,N_19982,N_19207);
and UO_225 (O_225,N_19674,N_18208);
nand UO_226 (O_226,N_19509,N_19834);
nand UO_227 (O_227,N_18261,N_19318);
nor UO_228 (O_228,N_18612,N_18618);
xnor UO_229 (O_229,N_18602,N_19718);
and UO_230 (O_230,N_18627,N_18918);
or UO_231 (O_231,N_18340,N_19807);
xor UO_232 (O_232,N_19757,N_19108);
xnor UO_233 (O_233,N_19859,N_18347);
or UO_234 (O_234,N_18439,N_19594);
nor UO_235 (O_235,N_19953,N_18298);
or UO_236 (O_236,N_18093,N_19008);
nand UO_237 (O_237,N_18826,N_18803);
or UO_238 (O_238,N_18285,N_18784);
nor UO_239 (O_239,N_19647,N_19963);
and UO_240 (O_240,N_18108,N_18617);
nand UO_241 (O_241,N_18917,N_19900);
nand UO_242 (O_242,N_19055,N_19954);
nor UO_243 (O_243,N_18165,N_19628);
xor UO_244 (O_244,N_18047,N_19083);
nand UO_245 (O_245,N_19518,N_19799);
nor UO_246 (O_246,N_18357,N_18049);
xor UO_247 (O_247,N_19731,N_19773);
and UO_248 (O_248,N_19841,N_19888);
xnor UO_249 (O_249,N_19521,N_19638);
and UO_250 (O_250,N_18570,N_18230);
xnor UO_251 (O_251,N_19808,N_19858);
xnor UO_252 (O_252,N_19660,N_18135);
and UO_253 (O_253,N_19479,N_19644);
and UO_254 (O_254,N_19073,N_18378);
xnor UO_255 (O_255,N_18792,N_19257);
or UO_256 (O_256,N_19774,N_18901);
nor UO_257 (O_257,N_18730,N_19505);
nor UO_258 (O_258,N_19027,N_19832);
xor UO_259 (O_259,N_19386,N_18289);
nand UO_260 (O_260,N_18379,N_18655);
nand UO_261 (O_261,N_18667,N_19189);
or UO_262 (O_262,N_19825,N_18941);
and UO_263 (O_263,N_18904,N_18659);
xor UO_264 (O_264,N_19238,N_18020);
nor UO_265 (O_265,N_18834,N_18472);
nor UO_266 (O_266,N_19678,N_19712);
or UO_267 (O_267,N_19169,N_18418);
nand UO_268 (O_268,N_18396,N_19778);
nand UO_269 (O_269,N_18902,N_18609);
or UO_270 (O_270,N_19903,N_19416);
or UO_271 (O_271,N_18949,N_19168);
and UO_272 (O_272,N_19625,N_19677);
xor UO_273 (O_273,N_18335,N_19984);
or UO_274 (O_274,N_19761,N_19232);
nand UO_275 (O_275,N_19838,N_18924);
nand UO_276 (O_276,N_19026,N_19051);
nor UO_277 (O_277,N_19639,N_19753);
and UO_278 (O_278,N_19927,N_19132);
or UO_279 (O_279,N_18729,N_19014);
and UO_280 (O_280,N_19830,N_19144);
or UO_281 (O_281,N_19406,N_18462);
or UO_282 (O_282,N_19340,N_18943);
xnor UO_283 (O_283,N_19545,N_18279);
or UO_284 (O_284,N_18256,N_18262);
and UO_285 (O_285,N_19057,N_19609);
or UO_286 (O_286,N_18575,N_18001);
nor UO_287 (O_287,N_19623,N_19262);
nand UO_288 (O_288,N_19071,N_18535);
xor UO_289 (O_289,N_18207,N_18287);
nand UO_290 (O_290,N_18174,N_18346);
and UO_291 (O_291,N_18948,N_19006);
and UO_292 (O_292,N_18668,N_18476);
and UO_293 (O_293,N_19725,N_19035);
nand UO_294 (O_294,N_19095,N_19653);
nand UO_295 (O_295,N_19948,N_19385);
xor UO_296 (O_296,N_19536,N_18407);
xor UO_297 (O_297,N_19265,N_18653);
or UO_298 (O_298,N_18721,N_18102);
nand UO_299 (O_299,N_18325,N_18269);
nand UO_300 (O_300,N_18095,N_18443);
and UO_301 (O_301,N_18367,N_19453);
nand UO_302 (O_302,N_18606,N_19397);
or UO_303 (O_303,N_19970,N_18345);
nor UO_304 (O_304,N_19767,N_18631);
and UO_305 (O_305,N_18561,N_19564);
xnor UO_306 (O_306,N_19760,N_19831);
or UO_307 (O_307,N_18992,N_19815);
and UO_308 (O_308,N_19915,N_18364);
and UO_309 (O_309,N_19631,N_18583);
nand UO_310 (O_310,N_19949,N_18543);
or UO_311 (O_311,N_18166,N_18011);
nor UO_312 (O_312,N_19597,N_19522);
xnor UO_313 (O_313,N_19158,N_18297);
nor UO_314 (O_314,N_19470,N_19601);
and UO_315 (O_315,N_18117,N_19269);
and UO_316 (O_316,N_18200,N_19343);
and UO_317 (O_317,N_19118,N_18796);
nor UO_318 (O_318,N_18178,N_18973);
xnor UO_319 (O_319,N_18812,N_19414);
nor UO_320 (O_320,N_18065,N_18500);
and UO_321 (O_321,N_18110,N_19017);
xnor UO_322 (O_322,N_19368,N_18425);
nor UO_323 (O_323,N_18016,N_19899);
or UO_324 (O_324,N_18740,N_19217);
nand UO_325 (O_325,N_18791,N_18843);
xor UO_326 (O_326,N_18073,N_18709);
xnor UO_327 (O_327,N_19464,N_18294);
or UO_328 (O_328,N_19556,N_19898);
or UO_329 (O_329,N_18832,N_19048);
nand UO_330 (O_330,N_18922,N_19222);
and UO_331 (O_331,N_18647,N_18006);
and UO_332 (O_332,N_19018,N_19724);
xnor UO_333 (O_333,N_19776,N_18229);
or UO_334 (O_334,N_19076,N_19050);
nor UO_335 (O_335,N_18591,N_18994);
and UO_336 (O_336,N_18786,N_18068);
and UO_337 (O_337,N_18334,N_18070);
and UO_338 (O_338,N_19373,N_18595);
and UO_339 (O_339,N_19156,N_19141);
or UO_340 (O_340,N_18715,N_19539);
nand UO_341 (O_341,N_19663,N_19358);
xor UO_342 (O_342,N_19117,N_18408);
nand UO_343 (O_343,N_19869,N_19508);
nand UO_344 (O_344,N_19091,N_18193);
nor UO_345 (O_345,N_19892,N_19193);
xnor UO_346 (O_346,N_18075,N_18125);
and UO_347 (O_347,N_18895,N_18468);
or UO_348 (O_348,N_19236,N_18217);
nor UO_349 (O_349,N_18623,N_19350);
and UO_350 (O_350,N_18244,N_18558);
or UO_351 (O_351,N_19229,N_18851);
nor UO_352 (O_352,N_18937,N_18392);
and UO_353 (O_353,N_19179,N_19323);
xor UO_354 (O_354,N_19185,N_18099);
nor UO_355 (O_355,N_18007,N_19772);
nor UO_356 (O_356,N_18828,N_18977);
nand UO_357 (O_357,N_19939,N_18662);
xor UO_358 (O_358,N_18009,N_19395);
nor UO_359 (O_359,N_19550,N_18026);
and UO_360 (O_360,N_18585,N_19698);
and UO_361 (O_361,N_18362,N_19205);
nand UO_362 (O_362,N_19409,N_18815);
nand UO_363 (O_363,N_18142,N_19094);
or UO_364 (O_364,N_18482,N_19765);
nand UO_365 (O_365,N_18755,N_19582);
nand UO_366 (O_366,N_18782,N_18264);
or UO_367 (O_367,N_19661,N_19910);
nor UO_368 (O_368,N_19636,N_19455);
nor UO_369 (O_369,N_19866,N_18920);
nand UO_370 (O_370,N_18931,N_19996);
xor UO_371 (O_371,N_18490,N_19780);
nand UO_372 (O_372,N_18678,N_19920);
xnor UO_373 (O_373,N_18384,N_19764);
nand UO_374 (O_374,N_18604,N_19572);
nand UO_375 (O_375,N_18466,N_19007);
nor UO_376 (O_376,N_18390,N_19360);
xnor UO_377 (O_377,N_19885,N_18749);
nor UO_378 (O_378,N_18956,N_18858);
nand UO_379 (O_379,N_19622,N_19985);
nor UO_380 (O_380,N_19103,N_18131);
and UO_381 (O_381,N_18829,N_18118);
nor UO_382 (O_382,N_19489,N_18574);
and UO_383 (O_383,N_18457,N_19306);
and UO_384 (O_384,N_19195,N_18748);
nand UO_385 (O_385,N_19228,N_18673);
nand UO_386 (O_386,N_18323,N_19646);
and UO_387 (O_387,N_19278,N_19288);
xnor UO_388 (O_388,N_19469,N_19847);
xnor UO_389 (O_389,N_19054,N_19936);
xnor UO_390 (O_390,N_18300,N_19642);
nor UO_391 (O_391,N_19417,N_19722);
or UO_392 (O_392,N_19552,N_19931);
and UO_393 (O_393,N_18754,N_19872);
or UO_394 (O_394,N_19686,N_19578);
nor UO_395 (O_395,N_18078,N_18303);
nor UO_396 (O_396,N_18876,N_18302);
and UO_397 (O_397,N_19785,N_19254);
xor UO_398 (O_398,N_19944,N_19099);
xnor UO_399 (O_399,N_19290,N_18533);
nor UO_400 (O_400,N_18189,N_19460);
nand UO_401 (O_401,N_19133,N_18024);
or UO_402 (O_402,N_19532,N_18801);
xnor UO_403 (O_403,N_18738,N_19868);
nor UO_404 (O_404,N_18238,N_18566);
xnor UO_405 (O_405,N_18355,N_18227);
or UO_406 (O_406,N_18616,N_18816);
xnor UO_407 (O_407,N_19268,N_19684);
or UO_408 (O_408,N_18950,N_18451);
xnor UO_409 (O_409,N_19314,N_18203);
nor UO_410 (O_410,N_18521,N_19178);
xor UO_411 (O_411,N_18000,N_19605);
nand UO_412 (O_412,N_18827,N_18580);
nor UO_413 (O_413,N_18877,N_18838);
nor UO_414 (O_414,N_19271,N_18484);
and UO_415 (O_415,N_19396,N_18932);
nand UO_416 (O_416,N_19361,N_19783);
or UO_417 (O_417,N_19924,N_19146);
nand UO_418 (O_418,N_18437,N_19172);
or UO_419 (O_419,N_18167,N_19946);
nand UO_420 (O_420,N_18654,N_19827);
xnor UO_421 (O_421,N_19041,N_19310);
or UO_422 (O_422,N_18210,N_19742);
or UO_423 (O_423,N_18584,N_18359);
or UO_424 (O_424,N_19563,N_19273);
nor UO_425 (O_425,N_19364,N_18911);
and UO_426 (O_426,N_18859,N_19192);
or UO_427 (O_427,N_19614,N_19001);
and UO_428 (O_428,N_18806,N_19426);
nor UO_429 (O_429,N_19127,N_19904);
xnor UO_430 (O_430,N_18419,N_19162);
xnor UO_431 (O_431,N_19298,N_19626);
xnor UO_432 (O_432,N_18372,N_18101);
and UO_433 (O_433,N_18004,N_19412);
and UO_434 (O_434,N_19296,N_18034);
xnor UO_435 (O_435,N_18096,N_18642);
xor UO_436 (O_436,N_18913,N_18725);
xor UO_437 (O_437,N_18664,N_19744);
and UO_438 (O_438,N_18693,N_18976);
xor UO_439 (O_439,N_18161,N_18593);
nor UO_440 (O_440,N_18925,N_18940);
xor UO_441 (O_441,N_18714,N_19398);
and UO_442 (O_442,N_18908,N_18670);
and UO_443 (O_443,N_18442,N_18934);
xnor UO_444 (O_444,N_19177,N_18544);
xnor UO_445 (O_445,N_18751,N_18276);
xnor UO_446 (O_446,N_19142,N_18191);
xor UO_447 (O_447,N_18458,N_18242);
xnor UO_448 (O_448,N_18507,N_18890);
xor UO_449 (O_449,N_18706,N_19527);
nor UO_450 (O_450,N_19584,N_18148);
and UO_451 (O_451,N_18250,N_18056);
nand UO_452 (O_452,N_18017,N_18927);
and UO_453 (O_453,N_18064,N_18744);
or UO_454 (O_454,N_18910,N_18253);
and UO_455 (O_455,N_18182,N_18291);
xnor UO_456 (O_456,N_19610,N_18732);
xor UO_457 (O_457,N_18299,N_18615);
xor UO_458 (O_458,N_18872,N_19180);
nand UO_459 (O_459,N_18536,N_18619);
nor UO_460 (O_460,N_18881,N_18438);
nand UO_461 (O_461,N_18900,N_19216);
or UO_462 (O_462,N_19150,N_18082);
nand UO_463 (O_463,N_19049,N_19507);
nand UO_464 (O_464,N_18779,N_18713);
nand UO_465 (O_465,N_18321,N_19392);
nor UO_466 (O_466,N_18650,N_19894);
or UO_467 (O_467,N_18807,N_18899);
nor UO_468 (O_468,N_19943,N_19573);
nor UO_469 (O_469,N_19641,N_19966);
nor UO_470 (O_470,N_19867,N_18061);
nor UO_471 (O_471,N_18519,N_19651);
xnor UO_472 (O_472,N_18326,N_18076);
nor UO_473 (O_473,N_19110,N_19727);
and UO_474 (O_474,N_19155,N_18479);
or UO_475 (O_475,N_18968,N_18204);
xor UO_476 (O_476,N_19703,N_18903);
nand UO_477 (O_477,N_18373,N_18103);
or UO_478 (O_478,N_19670,N_18090);
nor UO_479 (O_479,N_18327,N_18993);
or UO_480 (O_480,N_19843,N_19399);
or UO_481 (O_481,N_19432,N_19495);
or UO_482 (O_482,N_18506,N_18671);
nor UO_483 (O_483,N_19813,N_19362);
xnor UO_484 (O_484,N_19735,N_18578);
nand UO_485 (O_485,N_18172,N_18251);
and UO_486 (O_486,N_18187,N_19705);
or UO_487 (O_487,N_18811,N_18446);
xor UO_488 (O_488,N_18677,N_19833);
xnor UO_489 (O_489,N_19680,N_19856);
or UO_490 (O_490,N_19816,N_19329);
nand UO_491 (O_491,N_18098,N_19251);
and UO_492 (O_492,N_18030,N_18957);
nand UO_493 (O_493,N_19988,N_19919);
xor UO_494 (O_494,N_18465,N_18401);
nand UO_495 (O_495,N_18763,N_19285);
xnor UO_496 (O_496,N_19307,N_18802);
xnor UO_497 (O_497,N_19070,N_19467);
nor UO_498 (O_498,N_19533,N_19139);
nor UO_499 (O_499,N_18510,N_19884);
nor UO_500 (O_500,N_18220,N_18277);
xor UO_501 (O_501,N_19487,N_18234);
or UO_502 (O_502,N_18184,N_18862);
nand UO_503 (O_503,N_18423,N_18435);
or UO_504 (O_504,N_19557,N_19347);
nand UO_505 (O_505,N_18432,N_19081);
nand UO_506 (O_506,N_19821,N_19260);
nand UO_507 (O_507,N_18308,N_19068);
and UO_508 (O_508,N_18702,N_19082);
or UO_509 (O_509,N_19687,N_19851);
and UO_510 (O_510,N_18711,N_19516);
or UO_511 (O_511,N_18648,N_19770);
and UO_512 (O_512,N_19344,N_19471);
nand UO_513 (O_513,N_19377,N_18133);
or UO_514 (O_514,N_18304,N_19022);
nor UO_515 (O_515,N_19876,N_18257);
xnor UO_516 (O_516,N_18431,N_18557);
xnor UO_517 (O_517,N_19788,N_19754);
nor UO_518 (O_518,N_19183,N_19864);
nor UO_519 (O_519,N_18031,N_19842);
and UO_520 (O_520,N_18319,N_19419);
nor UO_521 (O_521,N_18524,N_18704);
and UO_522 (O_522,N_18722,N_18930);
nor UO_523 (O_523,N_18100,N_18233);
or UO_524 (O_524,N_19871,N_18274);
and UO_525 (O_525,N_19149,N_18978);
xnor UO_526 (O_526,N_19279,N_18582);
or UO_527 (O_527,N_19849,N_19028);
and UO_528 (O_528,N_18168,N_18162);
or UO_529 (O_529,N_18734,N_18413);
and UO_530 (O_530,N_19276,N_18385);
nand UO_531 (O_531,N_18690,N_18409);
and UO_532 (O_532,N_18497,N_19907);
xnor UO_533 (O_533,N_18620,N_18477);
xnor UO_534 (O_534,N_18128,N_18745);
nand UO_535 (O_535,N_19766,N_18850);
nand UO_536 (O_536,N_19492,N_18356);
xnor UO_537 (O_537,N_19136,N_19295);
nor UO_538 (O_538,N_19330,N_18371);
xnor UO_539 (O_539,N_18188,N_19901);
xnor UO_540 (O_540,N_19220,N_19692);
nand UO_541 (O_541,N_18218,N_18260);
and UO_542 (O_542,N_19877,N_19428);
nand UO_543 (O_543,N_18091,N_19715);
or UO_544 (O_544,N_19402,N_19292);
nor UO_545 (O_545,N_19458,N_19576);
nand UO_546 (O_546,N_19707,N_19305);
nand UO_547 (O_547,N_19450,N_18969);
and UO_548 (O_548,N_18318,N_19247);
nand UO_549 (O_549,N_19886,N_18038);
or UO_550 (O_550,N_19418,N_19689);
nand UO_551 (O_551,N_19166,N_19079);
or UO_552 (O_552,N_18886,N_18592);
and UO_553 (O_553,N_19316,N_19676);
nand UO_554 (O_554,N_19891,N_18863);
xor UO_555 (O_555,N_19032,N_19130);
xnor UO_556 (O_556,N_18766,N_19239);
nor UO_557 (O_557,N_18146,N_19297);
and UO_558 (O_558,N_19040,N_19500);
or UO_559 (O_559,N_18144,N_19287);
xor UO_560 (O_560,N_18053,N_19245);
nand UO_561 (O_561,N_18316,N_19758);
nand UO_562 (O_562,N_19599,N_19433);
nand UO_563 (O_563,N_19887,N_19266);
nor UO_564 (O_564,N_18848,N_19587);
nand UO_565 (O_565,N_18185,N_19606);
nor UO_566 (O_566,N_18511,N_19030);
or UO_567 (O_567,N_19308,N_19176);
nand UO_568 (O_568,N_19553,N_19917);
nand UO_569 (O_569,N_19131,N_19726);
or UO_570 (O_570,N_18470,N_18991);
or UO_571 (O_571,N_19664,N_18331);
xor UO_572 (O_572,N_18084,N_18660);
xor UO_573 (O_573,N_19439,N_18726);
nor UO_574 (O_574,N_18236,N_18586);
or UO_575 (O_575,N_19106,N_18205);
nor UO_576 (O_576,N_18079,N_19061);
nor UO_577 (O_577,N_18374,N_18889);
xor UO_578 (O_578,N_18433,N_19600);
nand UO_579 (O_579,N_19303,N_18774);
or UO_580 (O_580,N_18398,N_18239);
nor UO_581 (O_581,N_18349,N_18603);
and UO_582 (O_582,N_18568,N_19905);
xor UO_583 (O_583,N_18137,N_19122);
nand UO_584 (O_584,N_19947,N_19902);
nand UO_585 (O_585,N_18494,N_19657);
and UO_586 (O_586,N_19125,N_18415);
nand UO_587 (O_587,N_19304,N_19374);
or UO_588 (O_588,N_19562,N_19596);
nor UO_589 (O_589,N_19732,N_19248);
nand UO_590 (O_590,N_19544,N_19748);
or UO_591 (O_591,N_18005,N_19213);
nand UO_592 (O_592,N_18864,N_18282);
nand UO_593 (O_593,N_19734,N_18029);
nor UO_594 (O_594,N_18092,N_18998);
and UO_595 (O_595,N_18887,N_18149);
nor UO_596 (O_596,N_19950,N_18810);
xnor UO_597 (O_597,N_19121,N_19925);
and UO_598 (O_598,N_19147,N_18898);
or UO_599 (O_599,N_19388,N_18176);
nor UO_600 (O_600,N_19381,N_18153);
nor UO_601 (O_601,N_19086,N_18124);
nand UO_602 (O_602,N_19908,N_18388);
or UO_603 (O_603,N_18296,N_18232);
nor UO_604 (O_604,N_19611,N_19561);
nor UO_605 (O_605,N_18821,N_19976);
xor UO_606 (O_606,N_19721,N_18505);
xor UO_607 (O_607,N_18621,N_18195);
nor UO_608 (O_608,N_18046,N_19242);
xnor UO_609 (O_609,N_18134,N_18869);
nand UO_610 (O_610,N_18186,N_19342);
xnor UO_611 (O_611,N_18223,N_18306);
nor UO_612 (O_612,N_18666,N_19365);
and UO_613 (O_613,N_18057,N_19319);
or UO_614 (O_614,N_19787,N_18537);
and UO_615 (O_615,N_18450,N_19743);
nand UO_616 (O_616,N_18211,N_18028);
nand UO_617 (O_617,N_18703,N_18014);
or UO_618 (O_618,N_19294,N_19569);
nand UO_619 (O_619,N_19526,N_19789);
and UO_620 (O_620,N_18041,N_19154);
nor UO_621 (O_621,N_18503,N_18309);
nor UO_622 (O_622,N_19160,N_18867);
nor UO_623 (O_623,N_19463,N_19009);
or UO_624 (O_624,N_18594,N_18215);
or UO_625 (O_625,N_18123,N_18884);
nor UO_626 (O_626,N_19109,N_18179);
and UO_627 (O_627,N_18746,N_18417);
xor UO_628 (O_628,N_19852,N_19410);
or UO_629 (O_629,N_19800,N_19615);
xor UO_630 (O_630,N_19612,N_19085);
nand UO_631 (O_631,N_18540,N_18377);
xor UO_632 (O_632,N_19126,N_19066);
and UO_633 (O_633,N_19246,N_19717);
or UO_634 (O_634,N_19338,N_18054);
nor UO_635 (O_635,N_19531,N_18783);
or UO_636 (O_636,N_19893,N_18837);
nor UO_637 (O_637,N_18473,N_18814);
nor UO_638 (O_638,N_19112,N_18781);
and UO_639 (O_639,N_18410,N_19986);
nand UO_640 (O_640,N_19097,N_19688);
nand UO_641 (O_641,N_18959,N_19918);
nor UO_642 (O_642,N_19425,N_19044);
and UO_643 (O_643,N_18778,N_19701);
and UO_644 (O_644,N_18502,N_19494);
and UO_645 (O_645,N_18921,N_18508);
nand UO_646 (O_646,N_19695,N_18375);
xor UO_647 (O_647,N_18870,N_18456);
nor UO_648 (O_648,N_19356,N_19326);
nand UO_649 (O_649,N_18235,N_18564);
nand UO_650 (O_650,N_19063,N_19710);
nor UO_651 (O_651,N_19844,N_19775);
and UO_652 (O_652,N_19209,N_19512);
and UO_653 (O_653,N_19437,N_18600);
xnor UO_654 (O_654,N_19542,N_18464);
and UO_655 (O_655,N_18293,N_19879);
or UO_656 (O_656,N_19870,N_18382);
nand UO_657 (O_657,N_18143,N_19208);
xnor UO_658 (O_658,N_19630,N_19846);
xor UO_659 (O_659,N_18775,N_18893);
nor UO_660 (O_660,N_18597,N_19554);
nand UO_661 (O_661,N_19881,N_19665);
and UO_662 (O_662,N_19942,N_18972);
nand UO_663 (O_663,N_19046,N_19424);
nand UO_664 (O_664,N_19957,N_19036);
nor UO_665 (O_665,N_19331,N_19591);
and UO_666 (O_666,N_19270,N_19662);
nor UO_667 (O_667,N_18452,N_19762);
nor UO_668 (O_668,N_19299,N_19059);
or UO_669 (O_669,N_19441,N_18926);
nand UO_670 (O_670,N_19574,N_19791);
nand UO_671 (O_671,N_19235,N_19558);
xnor UO_672 (O_672,N_18971,N_19682);
nor UO_673 (O_673,N_19496,N_19714);
xor UO_674 (O_674,N_19465,N_18140);
nor UO_675 (O_675,N_18916,N_18946);
or UO_676 (O_676,N_18958,N_19352);
and UO_677 (O_677,N_19723,N_19391);
xnor UO_678 (O_678,N_18467,N_19882);
and UO_679 (O_679,N_19706,N_19475);
nor UO_680 (O_680,N_18699,N_18106);
and UO_681 (O_681,N_19589,N_19005);
and UO_682 (O_682,N_18018,N_19201);
and UO_683 (O_683,N_18228,N_19755);
nor UO_684 (O_684,N_18067,N_18645);
nand UO_685 (O_685,N_18332,N_19850);
nor UO_686 (O_686,N_19874,N_19317);
or UO_687 (O_687,N_18114,N_18254);
and UO_688 (O_688,N_19403,N_19602);
nor UO_689 (O_689,N_18938,N_19696);
and UO_690 (O_690,N_18601,N_19114);
or UO_691 (O_691,N_19274,N_19447);
and UO_692 (O_692,N_18109,N_19930);
xnor UO_693 (O_693,N_19673,N_19690);
and UO_694 (O_694,N_19031,N_19111);
nor UO_695 (O_695,N_18305,N_19648);
and UO_696 (O_696,N_19819,N_18701);
xor UO_697 (O_697,N_18360,N_18113);
nand UO_698 (O_698,N_18395,N_19140);
or UO_699 (O_699,N_18632,N_19474);
and UO_700 (O_700,N_18658,N_19482);
nand UO_701 (O_701,N_19603,N_18397);
nor UO_702 (O_702,N_18560,N_19157);
and UO_703 (O_703,N_19219,N_18240);
or UO_704 (O_704,N_18549,N_19023);
nand UO_705 (O_705,N_19510,N_18380);
nand UO_706 (O_706,N_18652,N_19443);
nor UO_707 (O_707,N_18343,N_18769);
or UO_708 (O_708,N_19956,N_18485);
or UO_709 (O_709,N_18988,N_19632);
and UO_710 (O_710,N_18163,N_19607);
nor UO_711 (O_711,N_19072,N_18975);
or UO_712 (O_712,N_18967,N_19914);
or UO_713 (O_713,N_19863,N_19534);
or UO_714 (O_714,N_18290,N_19434);
xnor UO_715 (O_715,N_19000,N_18033);
xnor UO_716 (O_716,N_19459,N_18281);
nor UO_717 (O_717,N_18935,N_18292);
nor UO_718 (O_718,N_19427,N_19922);
nand UO_719 (O_719,N_19252,N_18965);
xor UO_720 (O_720,N_18983,N_19400);
nor UO_721 (O_721,N_19993,N_19990);
xor UO_722 (O_722,N_19466,N_18739);
nand UO_723 (O_723,N_18896,N_18352);
xnor UO_724 (O_724,N_19935,N_19212);
or UO_725 (O_725,N_18267,N_19973);
or UO_726 (O_726,N_18157,N_19967);
nor UO_727 (O_727,N_19371,N_18545);
and UO_728 (O_728,N_18634,N_18984);
and UO_729 (O_729,N_19491,N_19581);
nand UO_730 (O_730,N_19817,N_18962);
nand UO_731 (O_731,N_19987,N_18145);
xor UO_732 (O_732,N_19190,N_18710);
or UO_733 (O_733,N_18164,N_19227);
nor UO_734 (O_734,N_18399,N_18400);
and UO_735 (O_735,N_18823,N_18311);
xor UO_736 (O_736,N_18528,N_18622);
nand UO_737 (O_737,N_18999,N_18515);
xnor UO_738 (O_738,N_18613,N_18680);
nand UO_739 (O_739,N_19649,N_19586);
and UO_740 (O_740,N_18243,N_18509);
nand UO_741 (O_741,N_19034,N_18111);
or UO_742 (O_742,N_19811,N_19197);
or UO_743 (O_743,N_19093,N_18329);
or UO_744 (O_744,N_18556,N_18492);
nor UO_745 (O_745,N_18818,N_19446);
xnor UO_746 (O_746,N_18406,N_19911);
and UO_747 (O_747,N_18841,N_18590);
or UO_748 (O_748,N_18344,N_19941);
nand UO_749 (O_749,N_18569,N_18169);
or UO_750 (O_750,N_18883,N_18231);
xor UO_751 (O_751,N_18687,N_18421);
nand UO_752 (O_752,N_19167,N_18341);
xor UO_753 (O_753,N_19835,N_19281);
or UO_754 (O_754,N_19498,N_19629);
and UO_755 (O_755,N_19004,N_19779);
nor UO_756 (O_756,N_18822,N_19488);
nand UO_757 (O_757,N_18879,N_19560);
nand UO_758 (O_758,N_18198,N_18209);
or UO_759 (O_759,N_18526,N_19003);
nand UO_760 (O_760,N_18273,N_19658);
and UO_761 (O_761,N_19794,N_19430);
xnor UO_762 (O_762,N_18156,N_19105);
nor UO_763 (O_763,N_18759,N_18605);
xnor UO_764 (O_764,N_19060,N_19964);
and UO_765 (O_765,N_19483,N_19384);
and UO_766 (O_766,N_19423,N_19565);
nand UO_767 (O_767,N_18121,N_19713);
or UO_768 (O_768,N_18776,N_19978);
and UO_769 (O_769,N_19568,N_19363);
nor UO_770 (O_770,N_18428,N_18270);
and UO_771 (O_771,N_18520,N_19857);
nand UO_772 (O_772,N_19598,N_18565);
xor UO_773 (O_773,N_18434,N_18871);
nand UO_774 (O_774,N_19165,N_18682);
nand UO_775 (O_775,N_19656,N_19519);
or UO_776 (O_776,N_18105,N_18348);
xnor UO_777 (O_777,N_18849,N_18830);
nand UO_778 (O_778,N_18365,N_19549);
and UO_779 (O_779,N_19826,N_19624);
xnor UO_780 (O_780,N_18449,N_19092);
nand UO_781 (O_781,N_19959,N_19480);
or UO_782 (O_782,N_19627,N_18338);
xnor UO_783 (O_783,N_18248,N_19301);
nor UO_784 (O_784,N_18012,N_18767);
nor UO_785 (O_785,N_19045,N_19369);
nand UO_786 (O_786,N_19263,N_19020);
nor UO_787 (O_787,N_18733,N_19311);
or UO_788 (O_788,N_19809,N_19504);
or UO_789 (O_789,N_18249,N_19137);
and UO_790 (O_790,N_18154,N_18762);
xnor UO_791 (O_791,N_18493,N_18320);
nor UO_792 (O_792,N_19258,N_19261);
xnor UO_793 (O_793,N_19694,N_19940);
xnor UO_794 (O_794,N_19422,N_19551);
or UO_795 (O_795,N_19814,N_19253);
nor UO_796 (O_796,N_18035,N_18201);
nand UO_797 (O_797,N_19913,N_19171);
nand UO_798 (O_798,N_19541,N_19445);
nand UO_799 (O_799,N_18393,N_18708);
and UO_800 (O_800,N_18915,N_19431);
nor UO_801 (O_801,N_19637,N_18237);
xor UO_802 (O_802,N_18454,N_19708);
nor UO_803 (O_803,N_19335,N_19024);
nor UO_804 (O_804,N_18171,N_19143);
nor UO_805 (O_805,N_18255,N_19517);
nand UO_806 (O_806,N_19332,N_18138);
xor UO_807 (O_807,N_18386,N_19571);
or UO_808 (O_808,N_19277,N_18088);
and UO_809 (O_809,N_18683,N_19895);
nand UO_810 (O_810,N_19828,N_19196);
nor UO_811 (O_811,N_18180,N_19520);
and UO_812 (O_812,N_19200,N_19259);
xor UO_813 (O_813,N_18429,N_18523);
or UO_814 (O_814,N_18736,N_19503);
xor UO_815 (O_815,N_18737,N_18809);
nand UO_816 (O_816,N_19339,N_19019);
and UO_817 (O_817,N_19991,N_19454);
nor UO_818 (O_818,N_19749,N_18698);
and UO_819 (O_819,N_19452,N_18919);
nand UO_820 (O_820,N_19792,N_18692);
nand UO_821 (O_821,N_19123,N_19955);
xnor UO_822 (O_822,N_19194,N_19672);
nand UO_823 (O_823,N_19173,N_18216);
xnor UO_824 (O_824,N_18656,N_18572);
and UO_825 (O_825,N_19769,N_19740);
xnor UO_826 (O_826,N_18027,N_18696);
and UO_827 (O_827,N_18483,N_19750);
xor UO_828 (O_828,N_19906,N_19393);
xor UO_829 (O_829,N_19580,N_19975);
nor UO_830 (O_830,N_19107,N_19502);
nand UO_831 (O_831,N_18104,N_18630);
xnor UO_832 (O_832,N_19567,N_18885);
xnor UO_833 (O_833,N_18643,N_19961);
xnor UO_834 (O_834,N_19313,N_19702);
or UO_835 (O_835,N_18225,N_19476);
nand UO_836 (O_836,N_18629,N_19588);
and UO_837 (O_837,N_18794,N_19321);
or UO_838 (O_838,N_19823,N_18579);
or UO_839 (O_839,N_18130,N_18122);
and UO_840 (O_840,N_18181,N_19186);
nand UO_841 (O_841,N_18022,N_18086);
or UO_842 (O_842,N_19608,N_18777);
or UO_843 (O_843,N_18936,N_18644);
xnor UO_844 (O_844,N_18756,N_18608);
or UO_845 (O_845,N_18275,N_18875);
nand UO_846 (O_846,N_18628,N_18354);
and UO_847 (O_847,N_18651,N_18874);
and UO_848 (O_848,N_19037,N_18127);
xor UO_849 (O_849,N_18554,N_19390);
xor UO_850 (O_850,N_18499,N_18478);
xor UO_851 (O_851,N_19804,N_19728);
nand UO_852 (O_852,N_19621,N_19394);
xor UO_853 (O_853,N_18083,N_19267);
or UO_854 (O_854,N_19243,N_18246);
nand UO_855 (O_855,N_19998,N_19065);
nor UO_856 (O_856,N_19666,N_18624);
or UO_857 (O_857,N_19746,N_18626);
nor UO_858 (O_858,N_18272,N_18944);
or UO_859 (O_859,N_19873,N_18376);
or UO_860 (O_860,N_18839,N_19226);
and UO_861 (O_861,N_19348,N_18799);
nor UO_862 (O_862,N_19370,N_18833);
nand UO_863 (O_863,N_19992,N_18152);
nor UO_864 (O_864,N_19089,N_18835);
or UO_865 (O_865,N_19793,N_18094);
xor UO_866 (O_866,N_19202,N_19372);
and UO_867 (O_867,N_19078,N_19378);
nor UO_868 (O_868,N_18252,N_18436);
or UO_869 (O_869,N_19897,N_18019);
xnor UO_870 (O_870,N_18795,N_19029);
or UO_871 (O_871,N_18856,N_18596);
xor UO_872 (O_872,N_18793,N_18970);
or UO_873 (O_873,N_19490,N_18322);
and UO_874 (O_874,N_19528,N_19282);
and UO_875 (O_875,N_19182,N_18072);
nand UO_876 (O_876,N_18263,N_19478);
nand UO_877 (O_877,N_18718,N_18990);
nand UO_878 (O_878,N_18542,N_19719);
and UO_879 (O_879,N_18530,N_18847);
xor UO_880 (O_880,N_19650,N_18480);
and UO_881 (O_881,N_19738,N_19429);
nor UO_882 (O_882,N_18080,N_18383);
and UO_883 (O_883,N_18514,N_19293);
nor UO_884 (O_884,N_18672,N_19328);
xnor UO_885 (O_885,N_18412,N_18050);
xnor UO_886 (O_886,N_18770,N_18550);
and UO_887 (O_887,N_19720,N_18036);
nand UO_888 (O_888,N_19322,N_19810);
and UO_889 (O_889,N_18226,N_18196);
nand UO_890 (O_890,N_19777,N_18861);
or UO_891 (O_891,N_19346,N_19523);
xnor UO_892 (O_892,N_18288,N_18641);
nor UO_893 (O_893,N_18222,N_19535);
nand UO_894 (O_894,N_18280,N_19134);
nor UO_895 (O_895,N_19436,N_19938);
xor UO_896 (O_896,N_18771,N_19681);
xor UO_897 (O_897,N_18787,N_19300);
nand UO_898 (O_898,N_19824,N_19234);
or UO_899 (O_899,N_19566,N_18459);
nand UO_900 (O_900,N_18819,N_19741);
or UO_901 (O_901,N_18689,N_18295);
nand UO_902 (O_902,N_18761,N_18808);
nor UO_903 (O_903,N_18116,N_18817);
and UO_904 (O_904,N_18405,N_18860);
xnor UO_905 (O_905,N_18370,N_19716);
nand UO_906 (O_906,N_18727,N_19822);
and UO_907 (O_907,N_19995,N_18611);
or UO_908 (O_908,N_19124,N_19548);
nand UO_909 (O_909,N_18278,N_19404);
nor UO_910 (O_910,N_18313,N_19355);
or UO_911 (O_911,N_18742,N_19420);
and UO_912 (O_912,N_19547,N_19181);
nor UO_913 (O_913,N_19958,N_19221);
or UO_914 (O_914,N_19896,N_18685);
nor UO_915 (O_915,N_18979,N_19230);
xor UO_916 (O_916,N_19366,N_18258);
and UO_917 (O_917,N_18015,N_19312);
and UO_918 (O_918,N_19805,N_18939);
or UO_919 (O_919,N_19711,N_18824);
nand UO_920 (O_920,N_19486,N_19214);
nand UO_921 (O_921,N_19100,N_19865);
xor UO_922 (O_922,N_19997,N_18587);
nor UO_923 (O_923,N_19188,N_19104);
nor UO_924 (O_924,N_19047,N_18455);
or UO_925 (O_925,N_18481,N_18788);
nor UO_926 (O_926,N_19383,N_19525);
nand UO_927 (O_927,N_19618,N_18753);
and UO_928 (O_928,N_18214,N_19187);
nor UO_929 (O_929,N_19972,N_18063);
nand UO_930 (O_930,N_18160,N_19053);
or UO_931 (O_931,N_19999,N_18888);
and UO_932 (O_932,N_18897,N_19203);
and UO_933 (O_933,N_19524,N_19357);
xor UO_934 (O_934,N_18119,N_18947);
or UO_935 (O_935,N_19619,N_19643);
nor UO_936 (O_936,N_19324,N_19739);
nor UO_937 (O_937,N_19359,N_18752);
nand UO_938 (O_938,N_19981,N_18175);
nor UO_939 (O_939,N_18501,N_18723);
nand UO_940 (O_940,N_19709,N_19438);
nand UO_941 (O_941,N_19782,N_19747);
and UO_942 (O_942,N_18071,N_18221);
or UO_943 (O_943,N_18271,N_19645);
nand UO_944 (O_944,N_18987,N_18504);
nor UO_945 (O_945,N_18661,N_18151);
nor UO_946 (O_946,N_19934,N_18646);
and UO_947 (O_947,N_18640,N_18857);
nand UO_948 (O_948,N_19345,N_18700);
xor UO_949 (O_949,N_18942,N_18717);
or UO_950 (O_950,N_19796,N_18607);
or UO_951 (O_951,N_19148,N_19002);
nor UO_952 (O_952,N_18212,N_19845);
nor UO_953 (O_953,N_19853,N_19264);
nand UO_954 (O_954,N_18813,N_19952);
and UO_955 (O_955,N_19204,N_19945);
xor UO_956 (O_956,N_19579,N_18052);
and UO_957 (O_957,N_18996,N_19751);
and UO_958 (O_958,N_18522,N_18842);
or UO_959 (O_959,N_18170,N_18317);
and UO_960 (O_960,N_19932,N_18336);
and UO_961 (O_961,N_18008,N_18923);
nand UO_962 (O_962,N_18120,N_19249);
nand UO_963 (O_963,N_18307,N_19098);
or UO_964 (O_964,N_18268,N_18852);
nand UO_965 (O_965,N_18486,N_18324);
nand UO_966 (O_966,N_18873,N_19275);
or UO_967 (O_967,N_19206,N_18764);
and UO_968 (O_968,N_19291,N_18190);
nor UO_969 (O_969,N_19389,N_19795);
and UO_970 (O_970,N_18986,N_18865);
xor UO_971 (O_971,N_19231,N_18440);
and UO_972 (O_972,N_19836,N_19415);
xor UO_973 (O_973,N_19367,N_19233);
and UO_974 (O_974,N_19854,N_19768);
nor UO_975 (O_975,N_18219,N_18964);
nor UO_976 (O_976,N_18567,N_18058);
nand UO_977 (O_977,N_18853,N_18573);
nor UO_978 (O_978,N_19056,N_19435);
nand UO_979 (O_979,N_19798,N_19583);
and UO_980 (O_980,N_18878,N_19797);
nand UO_981 (O_981,N_18081,N_19668);
xor UO_982 (O_982,N_19286,N_18951);
nor UO_983 (O_983,N_19215,N_18055);
xor UO_984 (O_984,N_19038,N_19700);
and UO_985 (O_985,N_18665,N_19128);
or UO_986 (O_986,N_19159,N_18197);
xnor UO_987 (O_987,N_18952,N_19704);
xnor UO_988 (O_988,N_18527,N_18531);
xnor UO_989 (O_989,N_18495,N_18266);
nand UO_990 (O_990,N_18173,N_19839);
xnor UO_991 (O_991,N_18663,N_19225);
xor UO_992 (O_992,N_19633,N_18598);
or UO_993 (O_993,N_18758,N_19555);
or UO_994 (O_994,N_18517,N_18206);
xnor UO_995 (O_995,N_19011,N_18301);
nor UO_996 (O_996,N_19595,N_19379);
or UO_997 (O_997,N_19737,N_18686);
and UO_998 (O_998,N_19515,N_18836);
nor UO_999 (O_999,N_19784,N_18363);
nand UO_1000 (O_1000,N_18567,N_19253);
or UO_1001 (O_1001,N_19109,N_18413);
and UO_1002 (O_1002,N_19020,N_19531);
or UO_1003 (O_1003,N_18764,N_18397);
nor UO_1004 (O_1004,N_18449,N_18134);
and UO_1005 (O_1005,N_19148,N_19932);
nand UO_1006 (O_1006,N_19321,N_18880);
or UO_1007 (O_1007,N_19110,N_19965);
nand UO_1008 (O_1008,N_18527,N_19029);
or UO_1009 (O_1009,N_18543,N_19924);
nor UO_1010 (O_1010,N_18627,N_18739);
nand UO_1011 (O_1011,N_19964,N_19980);
xor UO_1012 (O_1012,N_19366,N_18933);
nand UO_1013 (O_1013,N_18458,N_18604);
nand UO_1014 (O_1014,N_19102,N_18261);
or UO_1015 (O_1015,N_18095,N_19922);
and UO_1016 (O_1016,N_19066,N_19721);
and UO_1017 (O_1017,N_19599,N_19163);
or UO_1018 (O_1018,N_18290,N_18770);
or UO_1019 (O_1019,N_19094,N_18220);
or UO_1020 (O_1020,N_18501,N_18081);
or UO_1021 (O_1021,N_18549,N_19689);
nand UO_1022 (O_1022,N_18065,N_19165);
nor UO_1023 (O_1023,N_18348,N_18202);
nand UO_1024 (O_1024,N_18327,N_18270);
xor UO_1025 (O_1025,N_18347,N_19675);
nand UO_1026 (O_1026,N_18132,N_19098);
nand UO_1027 (O_1027,N_19059,N_19588);
nor UO_1028 (O_1028,N_18267,N_18901);
or UO_1029 (O_1029,N_19026,N_19053);
and UO_1030 (O_1030,N_18534,N_19019);
xor UO_1031 (O_1031,N_19290,N_18614);
nand UO_1032 (O_1032,N_18332,N_18093);
or UO_1033 (O_1033,N_18310,N_18975);
xor UO_1034 (O_1034,N_19480,N_19340);
and UO_1035 (O_1035,N_18221,N_19047);
nor UO_1036 (O_1036,N_19015,N_18816);
nand UO_1037 (O_1037,N_19220,N_18189);
nand UO_1038 (O_1038,N_19418,N_18928);
or UO_1039 (O_1039,N_19508,N_18283);
or UO_1040 (O_1040,N_19781,N_19772);
xnor UO_1041 (O_1041,N_19697,N_19922);
nor UO_1042 (O_1042,N_18855,N_19356);
nor UO_1043 (O_1043,N_19300,N_18860);
or UO_1044 (O_1044,N_18766,N_18505);
nor UO_1045 (O_1045,N_18487,N_18191);
xnor UO_1046 (O_1046,N_19598,N_18238);
xnor UO_1047 (O_1047,N_19307,N_18206);
nor UO_1048 (O_1048,N_19952,N_18828);
nor UO_1049 (O_1049,N_18031,N_18717);
xor UO_1050 (O_1050,N_18074,N_19748);
nor UO_1051 (O_1051,N_19599,N_19280);
nand UO_1052 (O_1052,N_18588,N_18079);
and UO_1053 (O_1053,N_18182,N_19787);
and UO_1054 (O_1054,N_19860,N_19897);
xnor UO_1055 (O_1055,N_18372,N_18274);
nand UO_1056 (O_1056,N_19131,N_19617);
nand UO_1057 (O_1057,N_19734,N_19409);
or UO_1058 (O_1058,N_19313,N_19417);
or UO_1059 (O_1059,N_18441,N_18348);
or UO_1060 (O_1060,N_18228,N_18276);
or UO_1061 (O_1061,N_19305,N_19410);
and UO_1062 (O_1062,N_19377,N_18311);
nand UO_1063 (O_1063,N_18386,N_19913);
nor UO_1064 (O_1064,N_19597,N_18921);
or UO_1065 (O_1065,N_19087,N_19095);
or UO_1066 (O_1066,N_19033,N_19699);
nand UO_1067 (O_1067,N_19762,N_18350);
nand UO_1068 (O_1068,N_18624,N_18792);
and UO_1069 (O_1069,N_19122,N_19368);
or UO_1070 (O_1070,N_19630,N_19568);
nor UO_1071 (O_1071,N_19048,N_19775);
nand UO_1072 (O_1072,N_19131,N_18454);
nor UO_1073 (O_1073,N_19279,N_18222);
xor UO_1074 (O_1074,N_19870,N_18001);
xor UO_1075 (O_1075,N_18040,N_19746);
and UO_1076 (O_1076,N_19803,N_18657);
nand UO_1077 (O_1077,N_18704,N_19211);
and UO_1078 (O_1078,N_19280,N_19548);
nor UO_1079 (O_1079,N_18587,N_18692);
nand UO_1080 (O_1080,N_18473,N_19621);
nand UO_1081 (O_1081,N_18839,N_18597);
nor UO_1082 (O_1082,N_19969,N_18552);
or UO_1083 (O_1083,N_19190,N_19770);
nand UO_1084 (O_1084,N_19509,N_18687);
xor UO_1085 (O_1085,N_18700,N_18589);
xnor UO_1086 (O_1086,N_18477,N_19793);
and UO_1087 (O_1087,N_18012,N_18166);
nor UO_1088 (O_1088,N_18541,N_18263);
nand UO_1089 (O_1089,N_18504,N_18300);
nor UO_1090 (O_1090,N_19494,N_18760);
and UO_1091 (O_1091,N_18977,N_18567);
or UO_1092 (O_1092,N_18797,N_18809);
xnor UO_1093 (O_1093,N_19264,N_19534);
and UO_1094 (O_1094,N_18913,N_18572);
nand UO_1095 (O_1095,N_19329,N_18057);
nand UO_1096 (O_1096,N_18262,N_19747);
xnor UO_1097 (O_1097,N_19755,N_18150);
or UO_1098 (O_1098,N_19687,N_18029);
nor UO_1099 (O_1099,N_18041,N_18627);
or UO_1100 (O_1100,N_19814,N_18349);
nor UO_1101 (O_1101,N_19544,N_19959);
nor UO_1102 (O_1102,N_19225,N_19493);
or UO_1103 (O_1103,N_18034,N_19397);
or UO_1104 (O_1104,N_19717,N_18105);
or UO_1105 (O_1105,N_19518,N_19841);
or UO_1106 (O_1106,N_18943,N_18987);
and UO_1107 (O_1107,N_19838,N_19898);
xor UO_1108 (O_1108,N_19881,N_19506);
nor UO_1109 (O_1109,N_19127,N_19510);
or UO_1110 (O_1110,N_19978,N_19063);
xnor UO_1111 (O_1111,N_18645,N_19772);
nor UO_1112 (O_1112,N_19475,N_18483);
xor UO_1113 (O_1113,N_18528,N_19288);
and UO_1114 (O_1114,N_18243,N_18417);
nand UO_1115 (O_1115,N_18494,N_19144);
xnor UO_1116 (O_1116,N_19463,N_18696);
or UO_1117 (O_1117,N_18657,N_18683);
or UO_1118 (O_1118,N_18307,N_18808);
or UO_1119 (O_1119,N_19266,N_18724);
nand UO_1120 (O_1120,N_18966,N_18422);
nor UO_1121 (O_1121,N_19608,N_18522);
nand UO_1122 (O_1122,N_19286,N_19237);
or UO_1123 (O_1123,N_19178,N_18677);
or UO_1124 (O_1124,N_18397,N_18688);
xnor UO_1125 (O_1125,N_19722,N_18072);
xor UO_1126 (O_1126,N_19046,N_18990);
nand UO_1127 (O_1127,N_18938,N_19307);
xor UO_1128 (O_1128,N_19894,N_19408);
nor UO_1129 (O_1129,N_19253,N_19866);
nand UO_1130 (O_1130,N_18440,N_19831);
or UO_1131 (O_1131,N_18817,N_19578);
and UO_1132 (O_1132,N_18894,N_19031);
and UO_1133 (O_1133,N_18014,N_18365);
xnor UO_1134 (O_1134,N_19073,N_19677);
nor UO_1135 (O_1135,N_19282,N_18111);
nor UO_1136 (O_1136,N_18063,N_18238);
or UO_1137 (O_1137,N_19885,N_18918);
nand UO_1138 (O_1138,N_19189,N_19411);
or UO_1139 (O_1139,N_19217,N_18258);
nor UO_1140 (O_1140,N_18754,N_19268);
nand UO_1141 (O_1141,N_19081,N_18905);
and UO_1142 (O_1142,N_18766,N_19615);
xor UO_1143 (O_1143,N_18478,N_19623);
nand UO_1144 (O_1144,N_19186,N_19911);
nor UO_1145 (O_1145,N_19787,N_19670);
nor UO_1146 (O_1146,N_19413,N_19161);
and UO_1147 (O_1147,N_19958,N_18338);
and UO_1148 (O_1148,N_18530,N_18745);
nor UO_1149 (O_1149,N_19025,N_19878);
nor UO_1150 (O_1150,N_19200,N_19371);
nor UO_1151 (O_1151,N_18763,N_18959);
nor UO_1152 (O_1152,N_18211,N_19441);
nor UO_1153 (O_1153,N_19962,N_18815);
nor UO_1154 (O_1154,N_19318,N_19578);
nand UO_1155 (O_1155,N_18456,N_18709);
and UO_1156 (O_1156,N_19639,N_19732);
nor UO_1157 (O_1157,N_18635,N_19625);
xor UO_1158 (O_1158,N_19590,N_19313);
nand UO_1159 (O_1159,N_19934,N_19049);
and UO_1160 (O_1160,N_19013,N_19627);
xnor UO_1161 (O_1161,N_18120,N_19663);
and UO_1162 (O_1162,N_18198,N_19719);
xnor UO_1163 (O_1163,N_18061,N_18273);
xor UO_1164 (O_1164,N_19280,N_18565);
and UO_1165 (O_1165,N_19151,N_18936);
nor UO_1166 (O_1166,N_18430,N_18236);
xnor UO_1167 (O_1167,N_18401,N_18189);
nor UO_1168 (O_1168,N_18113,N_18377);
nand UO_1169 (O_1169,N_19684,N_18072);
xnor UO_1170 (O_1170,N_18268,N_19995);
and UO_1171 (O_1171,N_18486,N_18460);
nor UO_1172 (O_1172,N_19615,N_19439);
and UO_1173 (O_1173,N_19097,N_19396);
xnor UO_1174 (O_1174,N_19059,N_18927);
nand UO_1175 (O_1175,N_19337,N_18938);
nand UO_1176 (O_1176,N_19348,N_18483);
nand UO_1177 (O_1177,N_19757,N_19739);
nor UO_1178 (O_1178,N_18819,N_19718);
nor UO_1179 (O_1179,N_19780,N_18425);
xnor UO_1180 (O_1180,N_18788,N_18993);
nand UO_1181 (O_1181,N_19812,N_18029);
and UO_1182 (O_1182,N_18680,N_19996);
or UO_1183 (O_1183,N_18867,N_19802);
and UO_1184 (O_1184,N_18707,N_18138);
or UO_1185 (O_1185,N_18176,N_18172);
nor UO_1186 (O_1186,N_19681,N_18592);
and UO_1187 (O_1187,N_19635,N_18296);
nand UO_1188 (O_1188,N_19202,N_18192);
nand UO_1189 (O_1189,N_19655,N_19496);
or UO_1190 (O_1190,N_18858,N_18823);
nand UO_1191 (O_1191,N_18742,N_19397);
xor UO_1192 (O_1192,N_18127,N_19445);
xnor UO_1193 (O_1193,N_19616,N_19276);
and UO_1194 (O_1194,N_19861,N_19644);
or UO_1195 (O_1195,N_19126,N_19546);
xnor UO_1196 (O_1196,N_18936,N_19862);
nor UO_1197 (O_1197,N_18783,N_18298);
or UO_1198 (O_1198,N_18052,N_19114);
xnor UO_1199 (O_1199,N_18072,N_19427);
and UO_1200 (O_1200,N_19963,N_19008);
xor UO_1201 (O_1201,N_19057,N_18820);
xnor UO_1202 (O_1202,N_19930,N_19517);
and UO_1203 (O_1203,N_18768,N_18930);
and UO_1204 (O_1204,N_18190,N_19676);
nand UO_1205 (O_1205,N_19777,N_19044);
nor UO_1206 (O_1206,N_19951,N_19601);
nor UO_1207 (O_1207,N_18941,N_18015);
or UO_1208 (O_1208,N_18606,N_19235);
and UO_1209 (O_1209,N_19620,N_19476);
or UO_1210 (O_1210,N_18083,N_18423);
and UO_1211 (O_1211,N_18916,N_18594);
xor UO_1212 (O_1212,N_18670,N_19758);
nand UO_1213 (O_1213,N_18517,N_18412);
nor UO_1214 (O_1214,N_19065,N_19619);
and UO_1215 (O_1215,N_18324,N_19746);
and UO_1216 (O_1216,N_18187,N_18125);
nor UO_1217 (O_1217,N_19276,N_19272);
and UO_1218 (O_1218,N_19038,N_19877);
nand UO_1219 (O_1219,N_18451,N_19939);
or UO_1220 (O_1220,N_18394,N_19379);
xor UO_1221 (O_1221,N_18737,N_19634);
nand UO_1222 (O_1222,N_18043,N_19180);
nor UO_1223 (O_1223,N_18092,N_18735);
nand UO_1224 (O_1224,N_18427,N_19033);
or UO_1225 (O_1225,N_19544,N_18599);
nor UO_1226 (O_1226,N_19851,N_19722);
xor UO_1227 (O_1227,N_19266,N_19391);
xor UO_1228 (O_1228,N_19959,N_18358);
and UO_1229 (O_1229,N_18279,N_19486);
xor UO_1230 (O_1230,N_18542,N_19716);
xnor UO_1231 (O_1231,N_19051,N_19477);
nor UO_1232 (O_1232,N_19179,N_18868);
nand UO_1233 (O_1233,N_19652,N_18071);
nor UO_1234 (O_1234,N_18719,N_18009);
nand UO_1235 (O_1235,N_19285,N_19471);
xnor UO_1236 (O_1236,N_19949,N_18450);
xnor UO_1237 (O_1237,N_18277,N_18732);
nor UO_1238 (O_1238,N_19981,N_19721);
nor UO_1239 (O_1239,N_18063,N_19621);
and UO_1240 (O_1240,N_19995,N_19161);
nand UO_1241 (O_1241,N_18449,N_18323);
nand UO_1242 (O_1242,N_19230,N_19539);
nand UO_1243 (O_1243,N_18185,N_19278);
and UO_1244 (O_1244,N_18493,N_18195);
xor UO_1245 (O_1245,N_19019,N_18990);
nor UO_1246 (O_1246,N_18585,N_19101);
or UO_1247 (O_1247,N_18165,N_19306);
or UO_1248 (O_1248,N_18180,N_18947);
or UO_1249 (O_1249,N_19640,N_19210);
and UO_1250 (O_1250,N_18531,N_18674);
xor UO_1251 (O_1251,N_18180,N_19499);
or UO_1252 (O_1252,N_19479,N_18420);
or UO_1253 (O_1253,N_18635,N_18150);
or UO_1254 (O_1254,N_19762,N_18858);
nor UO_1255 (O_1255,N_19877,N_19925);
and UO_1256 (O_1256,N_18260,N_19450);
nor UO_1257 (O_1257,N_18019,N_18490);
or UO_1258 (O_1258,N_18611,N_18234);
or UO_1259 (O_1259,N_19769,N_19764);
nor UO_1260 (O_1260,N_18363,N_19096);
nand UO_1261 (O_1261,N_19064,N_18301);
nor UO_1262 (O_1262,N_19890,N_18376);
xor UO_1263 (O_1263,N_19782,N_18594);
nand UO_1264 (O_1264,N_19457,N_19585);
xor UO_1265 (O_1265,N_19952,N_18356);
and UO_1266 (O_1266,N_18102,N_19777);
nor UO_1267 (O_1267,N_18963,N_19568);
nor UO_1268 (O_1268,N_18934,N_18214);
nor UO_1269 (O_1269,N_18875,N_18285);
nand UO_1270 (O_1270,N_18216,N_18506);
xnor UO_1271 (O_1271,N_18080,N_19391);
xnor UO_1272 (O_1272,N_19835,N_19575);
or UO_1273 (O_1273,N_19147,N_18777);
and UO_1274 (O_1274,N_19610,N_19792);
and UO_1275 (O_1275,N_19934,N_19573);
nand UO_1276 (O_1276,N_18581,N_19190);
or UO_1277 (O_1277,N_19282,N_19007);
nand UO_1278 (O_1278,N_19668,N_18287);
or UO_1279 (O_1279,N_19704,N_19322);
nand UO_1280 (O_1280,N_18193,N_18049);
nand UO_1281 (O_1281,N_19332,N_19331);
or UO_1282 (O_1282,N_19758,N_18935);
nor UO_1283 (O_1283,N_18532,N_19834);
or UO_1284 (O_1284,N_18231,N_19051);
or UO_1285 (O_1285,N_19847,N_18453);
xnor UO_1286 (O_1286,N_19048,N_19613);
or UO_1287 (O_1287,N_18921,N_18905);
nand UO_1288 (O_1288,N_19146,N_18801);
or UO_1289 (O_1289,N_18934,N_19297);
nor UO_1290 (O_1290,N_19894,N_18259);
xor UO_1291 (O_1291,N_19842,N_18018);
xnor UO_1292 (O_1292,N_19143,N_19507);
nor UO_1293 (O_1293,N_19887,N_18346);
nor UO_1294 (O_1294,N_18414,N_18081);
xnor UO_1295 (O_1295,N_19530,N_19855);
nand UO_1296 (O_1296,N_18091,N_19643);
nand UO_1297 (O_1297,N_19426,N_18821);
nor UO_1298 (O_1298,N_18817,N_19588);
and UO_1299 (O_1299,N_19718,N_19287);
and UO_1300 (O_1300,N_18220,N_18635);
xor UO_1301 (O_1301,N_18488,N_19579);
nand UO_1302 (O_1302,N_18070,N_18948);
and UO_1303 (O_1303,N_18504,N_18933);
and UO_1304 (O_1304,N_19774,N_19656);
nor UO_1305 (O_1305,N_19043,N_19074);
xor UO_1306 (O_1306,N_18258,N_18029);
nand UO_1307 (O_1307,N_18801,N_19820);
or UO_1308 (O_1308,N_19363,N_19252);
nand UO_1309 (O_1309,N_19964,N_19112);
nor UO_1310 (O_1310,N_19857,N_19955);
or UO_1311 (O_1311,N_18526,N_19732);
nand UO_1312 (O_1312,N_19916,N_18629);
and UO_1313 (O_1313,N_19953,N_18124);
nor UO_1314 (O_1314,N_18615,N_19302);
or UO_1315 (O_1315,N_19380,N_19401);
or UO_1316 (O_1316,N_18458,N_19121);
and UO_1317 (O_1317,N_19645,N_18331);
or UO_1318 (O_1318,N_19687,N_19774);
nand UO_1319 (O_1319,N_19989,N_18151);
xnor UO_1320 (O_1320,N_18682,N_18298);
nor UO_1321 (O_1321,N_18435,N_19667);
nand UO_1322 (O_1322,N_18464,N_19535);
xnor UO_1323 (O_1323,N_18889,N_18348);
and UO_1324 (O_1324,N_18400,N_19274);
nand UO_1325 (O_1325,N_19382,N_19825);
or UO_1326 (O_1326,N_19130,N_19645);
xor UO_1327 (O_1327,N_19087,N_18639);
nand UO_1328 (O_1328,N_18653,N_18477);
nor UO_1329 (O_1329,N_18011,N_19270);
and UO_1330 (O_1330,N_19442,N_18428);
nor UO_1331 (O_1331,N_19907,N_18447);
or UO_1332 (O_1332,N_18808,N_19812);
nor UO_1333 (O_1333,N_18729,N_19698);
and UO_1334 (O_1334,N_19537,N_19328);
and UO_1335 (O_1335,N_18903,N_19927);
xnor UO_1336 (O_1336,N_18048,N_19501);
nand UO_1337 (O_1337,N_19214,N_19201);
nor UO_1338 (O_1338,N_19575,N_18502);
nand UO_1339 (O_1339,N_18985,N_19243);
or UO_1340 (O_1340,N_18127,N_18375);
xor UO_1341 (O_1341,N_18130,N_18156);
xnor UO_1342 (O_1342,N_19988,N_19493);
nor UO_1343 (O_1343,N_18995,N_19129);
nand UO_1344 (O_1344,N_19260,N_19008);
xor UO_1345 (O_1345,N_19796,N_18345);
and UO_1346 (O_1346,N_19028,N_19102);
nor UO_1347 (O_1347,N_18838,N_19360);
xor UO_1348 (O_1348,N_18380,N_18854);
or UO_1349 (O_1349,N_19211,N_18153);
nor UO_1350 (O_1350,N_19173,N_18016);
xnor UO_1351 (O_1351,N_18414,N_18471);
nand UO_1352 (O_1352,N_19183,N_18961);
and UO_1353 (O_1353,N_19275,N_18568);
xnor UO_1354 (O_1354,N_19325,N_19156);
and UO_1355 (O_1355,N_19554,N_18398);
nor UO_1356 (O_1356,N_18642,N_18868);
and UO_1357 (O_1357,N_19569,N_19112);
nor UO_1358 (O_1358,N_19280,N_19976);
nor UO_1359 (O_1359,N_19422,N_18319);
and UO_1360 (O_1360,N_19047,N_18599);
nand UO_1361 (O_1361,N_19859,N_18015);
nand UO_1362 (O_1362,N_19294,N_18596);
and UO_1363 (O_1363,N_19248,N_18962);
nor UO_1364 (O_1364,N_18083,N_18323);
and UO_1365 (O_1365,N_19278,N_18992);
and UO_1366 (O_1366,N_19225,N_18713);
nor UO_1367 (O_1367,N_19350,N_19846);
nor UO_1368 (O_1368,N_19422,N_19227);
or UO_1369 (O_1369,N_18706,N_18707);
nand UO_1370 (O_1370,N_19771,N_19452);
nor UO_1371 (O_1371,N_18124,N_19090);
or UO_1372 (O_1372,N_19348,N_18720);
and UO_1373 (O_1373,N_18073,N_19051);
nand UO_1374 (O_1374,N_19059,N_19780);
nand UO_1375 (O_1375,N_18751,N_18539);
xor UO_1376 (O_1376,N_18002,N_19423);
or UO_1377 (O_1377,N_19406,N_19241);
nor UO_1378 (O_1378,N_18953,N_18258);
and UO_1379 (O_1379,N_19897,N_18782);
or UO_1380 (O_1380,N_18793,N_18053);
xnor UO_1381 (O_1381,N_18935,N_18258);
nand UO_1382 (O_1382,N_18937,N_18402);
or UO_1383 (O_1383,N_19247,N_18287);
and UO_1384 (O_1384,N_18180,N_19547);
nand UO_1385 (O_1385,N_19783,N_19636);
nand UO_1386 (O_1386,N_18371,N_19591);
and UO_1387 (O_1387,N_18809,N_18302);
nor UO_1388 (O_1388,N_18235,N_19443);
nor UO_1389 (O_1389,N_18730,N_19759);
xor UO_1390 (O_1390,N_18827,N_19566);
and UO_1391 (O_1391,N_19446,N_19925);
and UO_1392 (O_1392,N_19296,N_18714);
nand UO_1393 (O_1393,N_19426,N_18654);
nor UO_1394 (O_1394,N_18119,N_19398);
nand UO_1395 (O_1395,N_18013,N_19686);
xor UO_1396 (O_1396,N_19942,N_18009);
xnor UO_1397 (O_1397,N_18381,N_19399);
nor UO_1398 (O_1398,N_18062,N_18374);
nand UO_1399 (O_1399,N_19157,N_19388);
or UO_1400 (O_1400,N_18318,N_19974);
nor UO_1401 (O_1401,N_19232,N_19377);
nand UO_1402 (O_1402,N_19713,N_18641);
and UO_1403 (O_1403,N_18710,N_19690);
and UO_1404 (O_1404,N_19695,N_18537);
and UO_1405 (O_1405,N_19144,N_19281);
nand UO_1406 (O_1406,N_19426,N_18733);
or UO_1407 (O_1407,N_19030,N_19294);
or UO_1408 (O_1408,N_19546,N_18886);
and UO_1409 (O_1409,N_19542,N_18611);
and UO_1410 (O_1410,N_19959,N_19717);
and UO_1411 (O_1411,N_19989,N_19210);
or UO_1412 (O_1412,N_19500,N_18570);
or UO_1413 (O_1413,N_19071,N_18753);
and UO_1414 (O_1414,N_19144,N_19607);
nand UO_1415 (O_1415,N_19714,N_19204);
xor UO_1416 (O_1416,N_19500,N_19922);
and UO_1417 (O_1417,N_19961,N_19391);
xor UO_1418 (O_1418,N_18255,N_19867);
or UO_1419 (O_1419,N_19060,N_19267);
or UO_1420 (O_1420,N_19174,N_19956);
xnor UO_1421 (O_1421,N_19086,N_18112);
or UO_1422 (O_1422,N_18536,N_19745);
or UO_1423 (O_1423,N_19587,N_19360);
or UO_1424 (O_1424,N_18573,N_18677);
or UO_1425 (O_1425,N_18553,N_19000);
and UO_1426 (O_1426,N_18842,N_18694);
or UO_1427 (O_1427,N_18568,N_19586);
or UO_1428 (O_1428,N_18331,N_19600);
nand UO_1429 (O_1429,N_19000,N_19455);
xnor UO_1430 (O_1430,N_19790,N_19827);
nor UO_1431 (O_1431,N_19587,N_19613);
xor UO_1432 (O_1432,N_18869,N_19698);
or UO_1433 (O_1433,N_19234,N_18109);
nand UO_1434 (O_1434,N_18024,N_18702);
or UO_1435 (O_1435,N_19092,N_19977);
or UO_1436 (O_1436,N_18947,N_18496);
nor UO_1437 (O_1437,N_18229,N_19831);
nor UO_1438 (O_1438,N_19102,N_19242);
and UO_1439 (O_1439,N_18331,N_18973);
and UO_1440 (O_1440,N_18284,N_19180);
xor UO_1441 (O_1441,N_19002,N_19557);
xnor UO_1442 (O_1442,N_18375,N_18773);
and UO_1443 (O_1443,N_18466,N_18563);
or UO_1444 (O_1444,N_19764,N_19780);
and UO_1445 (O_1445,N_19444,N_19501);
nand UO_1446 (O_1446,N_19795,N_18912);
or UO_1447 (O_1447,N_18880,N_19863);
nor UO_1448 (O_1448,N_19012,N_19461);
nand UO_1449 (O_1449,N_18338,N_19067);
and UO_1450 (O_1450,N_19054,N_18666);
and UO_1451 (O_1451,N_18394,N_19265);
and UO_1452 (O_1452,N_18419,N_19141);
xnor UO_1453 (O_1453,N_18318,N_19774);
or UO_1454 (O_1454,N_18628,N_19245);
or UO_1455 (O_1455,N_19376,N_19926);
or UO_1456 (O_1456,N_18601,N_18348);
and UO_1457 (O_1457,N_19582,N_19507);
or UO_1458 (O_1458,N_19356,N_19198);
and UO_1459 (O_1459,N_19092,N_19437);
xnor UO_1460 (O_1460,N_19241,N_19779);
or UO_1461 (O_1461,N_18941,N_18700);
or UO_1462 (O_1462,N_19590,N_18197);
nand UO_1463 (O_1463,N_19878,N_18267);
and UO_1464 (O_1464,N_18187,N_19384);
and UO_1465 (O_1465,N_19453,N_18949);
and UO_1466 (O_1466,N_18377,N_18129);
and UO_1467 (O_1467,N_19641,N_18872);
or UO_1468 (O_1468,N_19343,N_18942);
xor UO_1469 (O_1469,N_18952,N_19388);
xnor UO_1470 (O_1470,N_18484,N_18575);
xnor UO_1471 (O_1471,N_18444,N_19722);
and UO_1472 (O_1472,N_18277,N_18923);
and UO_1473 (O_1473,N_18462,N_18162);
or UO_1474 (O_1474,N_19770,N_19397);
xor UO_1475 (O_1475,N_18946,N_19406);
nor UO_1476 (O_1476,N_19890,N_18827);
nand UO_1477 (O_1477,N_18472,N_18761);
or UO_1478 (O_1478,N_19534,N_18106);
and UO_1479 (O_1479,N_18258,N_19014);
nor UO_1480 (O_1480,N_19768,N_19008);
nand UO_1481 (O_1481,N_18766,N_19000);
and UO_1482 (O_1482,N_18576,N_18228);
or UO_1483 (O_1483,N_18315,N_19135);
nand UO_1484 (O_1484,N_19917,N_19996);
xnor UO_1485 (O_1485,N_19243,N_19887);
or UO_1486 (O_1486,N_19361,N_19382);
nand UO_1487 (O_1487,N_19394,N_18166);
xnor UO_1488 (O_1488,N_19458,N_19433);
xor UO_1489 (O_1489,N_18096,N_18909);
and UO_1490 (O_1490,N_18123,N_18381);
xnor UO_1491 (O_1491,N_18169,N_19631);
nor UO_1492 (O_1492,N_18306,N_19885);
and UO_1493 (O_1493,N_18224,N_18751);
nor UO_1494 (O_1494,N_18548,N_18561);
and UO_1495 (O_1495,N_19593,N_19127);
or UO_1496 (O_1496,N_19968,N_18091);
nand UO_1497 (O_1497,N_18782,N_19094);
and UO_1498 (O_1498,N_18912,N_18102);
and UO_1499 (O_1499,N_19281,N_19229);
xor UO_1500 (O_1500,N_19939,N_19940);
nand UO_1501 (O_1501,N_19855,N_19362);
xnor UO_1502 (O_1502,N_18221,N_19972);
and UO_1503 (O_1503,N_19921,N_18003);
nand UO_1504 (O_1504,N_18803,N_19282);
nor UO_1505 (O_1505,N_19353,N_18258);
or UO_1506 (O_1506,N_18116,N_19391);
or UO_1507 (O_1507,N_18507,N_19520);
xor UO_1508 (O_1508,N_19212,N_18868);
and UO_1509 (O_1509,N_18883,N_18523);
nand UO_1510 (O_1510,N_18355,N_19201);
xor UO_1511 (O_1511,N_18291,N_18695);
and UO_1512 (O_1512,N_18520,N_19742);
xnor UO_1513 (O_1513,N_19378,N_19200);
nand UO_1514 (O_1514,N_19143,N_19240);
nand UO_1515 (O_1515,N_18080,N_18475);
or UO_1516 (O_1516,N_19483,N_19724);
or UO_1517 (O_1517,N_19897,N_18209);
or UO_1518 (O_1518,N_19343,N_19832);
or UO_1519 (O_1519,N_19878,N_19368);
or UO_1520 (O_1520,N_19973,N_19143);
nand UO_1521 (O_1521,N_18640,N_19208);
nand UO_1522 (O_1522,N_19738,N_18755);
nand UO_1523 (O_1523,N_19649,N_18140);
xor UO_1524 (O_1524,N_18602,N_18852);
and UO_1525 (O_1525,N_19297,N_18476);
xnor UO_1526 (O_1526,N_19829,N_19759);
and UO_1527 (O_1527,N_18678,N_19982);
and UO_1528 (O_1528,N_19071,N_19942);
xnor UO_1529 (O_1529,N_18916,N_19817);
nand UO_1530 (O_1530,N_18695,N_18578);
or UO_1531 (O_1531,N_18886,N_18803);
or UO_1532 (O_1532,N_18159,N_19838);
or UO_1533 (O_1533,N_19203,N_19012);
nor UO_1534 (O_1534,N_19344,N_19149);
or UO_1535 (O_1535,N_19741,N_19120);
xnor UO_1536 (O_1536,N_18416,N_18947);
nor UO_1537 (O_1537,N_19938,N_18990);
nand UO_1538 (O_1538,N_19101,N_19751);
xnor UO_1539 (O_1539,N_19061,N_19655);
nand UO_1540 (O_1540,N_19767,N_19317);
or UO_1541 (O_1541,N_19149,N_19568);
xor UO_1542 (O_1542,N_19393,N_19416);
nor UO_1543 (O_1543,N_18188,N_19753);
nand UO_1544 (O_1544,N_18321,N_19373);
or UO_1545 (O_1545,N_19224,N_19786);
or UO_1546 (O_1546,N_18372,N_18562);
nor UO_1547 (O_1547,N_19037,N_18751);
and UO_1548 (O_1548,N_19832,N_19684);
xnor UO_1549 (O_1549,N_19825,N_18881);
nand UO_1550 (O_1550,N_19480,N_19676);
nand UO_1551 (O_1551,N_18493,N_19283);
and UO_1552 (O_1552,N_18205,N_18174);
nor UO_1553 (O_1553,N_19205,N_19446);
xor UO_1554 (O_1554,N_18060,N_18693);
xnor UO_1555 (O_1555,N_19639,N_18368);
xor UO_1556 (O_1556,N_19674,N_18632);
xor UO_1557 (O_1557,N_18622,N_19771);
nand UO_1558 (O_1558,N_19586,N_18058);
and UO_1559 (O_1559,N_18953,N_18225);
and UO_1560 (O_1560,N_18356,N_18198);
nor UO_1561 (O_1561,N_18573,N_19913);
and UO_1562 (O_1562,N_19354,N_18270);
nand UO_1563 (O_1563,N_19174,N_19856);
and UO_1564 (O_1564,N_18520,N_19277);
or UO_1565 (O_1565,N_19838,N_19739);
nor UO_1566 (O_1566,N_19784,N_19671);
xor UO_1567 (O_1567,N_18349,N_18389);
nor UO_1568 (O_1568,N_19713,N_18290);
or UO_1569 (O_1569,N_19958,N_18153);
nand UO_1570 (O_1570,N_18137,N_18189);
and UO_1571 (O_1571,N_19238,N_19763);
nand UO_1572 (O_1572,N_18029,N_19458);
xnor UO_1573 (O_1573,N_19651,N_18295);
or UO_1574 (O_1574,N_18741,N_18641);
nand UO_1575 (O_1575,N_18049,N_18609);
nor UO_1576 (O_1576,N_18985,N_19561);
nor UO_1577 (O_1577,N_19035,N_19472);
nand UO_1578 (O_1578,N_18423,N_18320);
nand UO_1579 (O_1579,N_18964,N_19642);
or UO_1580 (O_1580,N_19593,N_18737);
nand UO_1581 (O_1581,N_18125,N_18119);
nand UO_1582 (O_1582,N_18622,N_18723);
nor UO_1583 (O_1583,N_18327,N_19141);
or UO_1584 (O_1584,N_18716,N_18629);
xnor UO_1585 (O_1585,N_19452,N_18167);
and UO_1586 (O_1586,N_19723,N_19651);
nor UO_1587 (O_1587,N_19677,N_19359);
and UO_1588 (O_1588,N_18182,N_19736);
or UO_1589 (O_1589,N_18433,N_19646);
xnor UO_1590 (O_1590,N_18562,N_18681);
nand UO_1591 (O_1591,N_19942,N_18959);
or UO_1592 (O_1592,N_18706,N_18521);
nand UO_1593 (O_1593,N_19946,N_18658);
or UO_1594 (O_1594,N_19273,N_18793);
xor UO_1595 (O_1595,N_19944,N_19868);
nand UO_1596 (O_1596,N_18262,N_18933);
xnor UO_1597 (O_1597,N_19031,N_18527);
nand UO_1598 (O_1598,N_19577,N_18815);
or UO_1599 (O_1599,N_18321,N_18579);
nand UO_1600 (O_1600,N_19974,N_18772);
and UO_1601 (O_1601,N_18902,N_18106);
nand UO_1602 (O_1602,N_18928,N_19043);
xnor UO_1603 (O_1603,N_18158,N_19718);
or UO_1604 (O_1604,N_18142,N_18490);
nor UO_1605 (O_1605,N_19870,N_19837);
and UO_1606 (O_1606,N_18557,N_18539);
nand UO_1607 (O_1607,N_19843,N_18279);
nor UO_1608 (O_1608,N_19111,N_18863);
and UO_1609 (O_1609,N_19739,N_19880);
nand UO_1610 (O_1610,N_18563,N_18301);
nand UO_1611 (O_1611,N_18123,N_18091);
nor UO_1612 (O_1612,N_18681,N_19154);
nand UO_1613 (O_1613,N_18210,N_19936);
and UO_1614 (O_1614,N_19193,N_18500);
nor UO_1615 (O_1615,N_18777,N_18346);
and UO_1616 (O_1616,N_18388,N_18892);
or UO_1617 (O_1617,N_19469,N_18358);
nor UO_1618 (O_1618,N_19390,N_18937);
and UO_1619 (O_1619,N_18166,N_19688);
nand UO_1620 (O_1620,N_18498,N_18939);
or UO_1621 (O_1621,N_19524,N_18026);
nor UO_1622 (O_1622,N_18761,N_18506);
and UO_1623 (O_1623,N_19315,N_19195);
and UO_1624 (O_1624,N_19975,N_19787);
or UO_1625 (O_1625,N_19753,N_19389);
and UO_1626 (O_1626,N_18517,N_19769);
or UO_1627 (O_1627,N_18044,N_18938);
or UO_1628 (O_1628,N_18499,N_18167);
nor UO_1629 (O_1629,N_19386,N_19278);
nor UO_1630 (O_1630,N_18512,N_19285);
or UO_1631 (O_1631,N_18000,N_18551);
or UO_1632 (O_1632,N_18301,N_18787);
or UO_1633 (O_1633,N_19195,N_19496);
nor UO_1634 (O_1634,N_19228,N_19933);
nor UO_1635 (O_1635,N_18457,N_18303);
nand UO_1636 (O_1636,N_19864,N_19038);
nor UO_1637 (O_1637,N_19822,N_19044);
nand UO_1638 (O_1638,N_18191,N_19299);
or UO_1639 (O_1639,N_18582,N_19964);
and UO_1640 (O_1640,N_19510,N_19479);
nand UO_1641 (O_1641,N_19410,N_19110);
nor UO_1642 (O_1642,N_18073,N_18153);
nand UO_1643 (O_1643,N_19167,N_19423);
xor UO_1644 (O_1644,N_18762,N_18392);
xnor UO_1645 (O_1645,N_18431,N_19545);
or UO_1646 (O_1646,N_18321,N_18817);
nand UO_1647 (O_1647,N_19207,N_19378);
xnor UO_1648 (O_1648,N_18987,N_18146);
nor UO_1649 (O_1649,N_19504,N_19220);
nand UO_1650 (O_1650,N_18609,N_19914);
nor UO_1651 (O_1651,N_18669,N_19512);
or UO_1652 (O_1652,N_18937,N_18894);
nand UO_1653 (O_1653,N_19724,N_18761);
nor UO_1654 (O_1654,N_19485,N_18870);
nand UO_1655 (O_1655,N_19183,N_18765);
and UO_1656 (O_1656,N_18560,N_19211);
xor UO_1657 (O_1657,N_18757,N_18552);
xnor UO_1658 (O_1658,N_19379,N_18048);
nand UO_1659 (O_1659,N_19319,N_18235);
nand UO_1660 (O_1660,N_18090,N_19812);
xor UO_1661 (O_1661,N_19154,N_18688);
nand UO_1662 (O_1662,N_19136,N_18973);
nand UO_1663 (O_1663,N_19302,N_19931);
nand UO_1664 (O_1664,N_19386,N_18387);
xor UO_1665 (O_1665,N_18558,N_19082);
and UO_1666 (O_1666,N_18908,N_19206);
xnor UO_1667 (O_1667,N_19142,N_19467);
nor UO_1668 (O_1668,N_18568,N_19569);
xor UO_1669 (O_1669,N_18681,N_18081);
nor UO_1670 (O_1670,N_18407,N_19102);
nor UO_1671 (O_1671,N_18574,N_18436);
and UO_1672 (O_1672,N_18551,N_18947);
nor UO_1673 (O_1673,N_18277,N_19135);
and UO_1674 (O_1674,N_19575,N_19543);
and UO_1675 (O_1675,N_19584,N_18081);
nor UO_1676 (O_1676,N_18861,N_18574);
nand UO_1677 (O_1677,N_19451,N_19570);
and UO_1678 (O_1678,N_19319,N_18924);
nor UO_1679 (O_1679,N_18068,N_18829);
nand UO_1680 (O_1680,N_19909,N_19836);
nor UO_1681 (O_1681,N_19922,N_19912);
xnor UO_1682 (O_1682,N_19839,N_19677);
or UO_1683 (O_1683,N_18182,N_19447);
xor UO_1684 (O_1684,N_18310,N_18904);
nand UO_1685 (O_1685,N_18673,N_19802);
xor UO_1686 (O_1686,N_18180,N_19369);
xor UO_1687 (O_1687,N_19229,N_19330);
and UO_1688 (O_1688,N_19306,N_18628);
xor UO_1689 (O_1689,N_19484,N_18220);
xnor UO_1690 (O_1690,N_18915,N_18515);
or UO_1691 (O_1691,N_19214,N_18158);
nor UO_1692 (O_1692,N_18276,N_18584);
xnor UO_1693 (O_1693,N_18158,N_19317);
xnor UO_1694 (O_1694,N_19828,N_19844);
nand UO_1695 (O_1695,N_18867,N_19037);
and UO_1696 (O_1696,N_19084,N_19157);
or UO_1697 (O_1697,N_19576,N_18449);
or UO_1698 (O_1698,N_19673,N_19614);
and UO_1699 (O_1699,N_18269,N_19356);
xnor UO_1700 (O_1700,N_18993,N_19044);
and UO_1701 (O_1701,N_18806,N_18269);
nor UO_1702 (O_1702,N_19235,N_19434);
nand UO_1703 (O_1703,N_19147,N_18503);
or UO_1704 (O_1704,N_18212,N_19758);
nand UO_1705 (O_1705,N_19433,N_19308);
xnor UO_1706 (O_1706,N_19333,N_19501);
nand UO_1707 (O_1707,N_19944,N_18719);
nand UO_1708 (O_1708,N_19166,N_19988);
xnor UO_1709 (O_1709,N_18638,N_19739);
nor UO_1710 (O_1710,N_19571,N_19011);
nor UO_1711 (O_1711,N_18795,N_19374);
or UO_1712 (O_1712,N_19514,N_19528);
and UO_1713 (O_1713,N_18635,N_19380);
and UO_1714 (O_1714,N_18336,N_18193);
nor UO_1715 (O_1715,N_19559,N_18338);
nand UO_1716 (O_1716,N_19385,N_19367);
and UO_1717 (O_1717,N_19602,N_19007);
or UO_1718 (O_1718,N_19701,N_18586);
or UO_1719 (O_1719,N_19488,N_18192);
xnor UO_1720 (O_1720,N_18823,N_18511);
nand UO_1721 (O_1721,N_19101,N_18057);
or UO_1722 (O_1722,N_19817,N_18185);
or UO_1723 (O_1723,N_18213,N_18385);
xnor UO_1724 (O_1724,N_18016,N_18518);
or UO_1725 (O_1725,N_19619,N_19636);
or UO_1726 (O_1726,N_18932,N_19326);
and UO_1727 (O_1727,N_18901,N_19610);
and UO_1728 (O_1728,N_19145,N_19522);
xor UO_1729 (O_1729,N_19067,N_19992);
xnor UO_1730 (O_1730,N_18079,N_19339);
nor UO_1731 (O_1731,N_19175,N_19826);
or UO_1732 (O_1732,N_19278,N_19924);
nand UO_1733 (O_1733,N_19179,N_19271);
xor UO_1734 (O_1734,N_19760,N_19125);
or UO_1735 (O_1735,N_19872,N_18006);
nor UO_1736 (O_1736,N_18872,N_18317);
nor UO_1737 (O_1737,N_18004,N_19744);
or UO_1738 (O_1738,N_19032,N_18093);
and UO_1739 (O_1739,N_19010,N_19986);
nand UO_1740 (O_1740,N_18589,N_19303);
xnor UO_1741 (O_1741,N_18627,N_18828);
and UO_1742 (O_1742,N_19390,N_19580);
or UO_1743 (O_1743,N_19091,N_18424);
xor UO_1744 (O_1744,N_18488,N_19481);
and UO_1745 (O_1745,N_19742,N_18560);
or UO_1746 (O_1746,N_18636,N_19874);
or UO_1747 (O_1747,N_19566,N_18230);
nor UO_1748 (O_1748,N_19859,N_19954);
nand UO_1749 (O_1749,N_19144,N_18918);
nor UO_1750 (O_1750,N_19944,N_18116);
nand UO_1751 (O_1751,N_19618,N_18266);
and UO_1752 (O_1752,N_18993,N_18236);
xor UO_1753 (O_1753,N_18803,N_19360);
nand UO_1754 (O_1754,N_18497,N_18110);
xor UO_1755 (O_1755,N_19665,N_18924);
and UO_1756 (O_1756,N_19123,N_19037);
nor UO_1757 (O_1757,N_18317,N_18560);
nor UO_1758 (O_1758,N_19248,N_18539);
or UO_1759 (O_1759,N_18063,N_18983);
xnor UO_1760 (O_1760,N_19432,N_18681);
and UO_1761 (O_1761,N_19624,N_19906);
nor UO_1762 (O_1762,N_19347,N_19578);
nor UO_1763 (O_1763,N_18368,N_18985);
nand UO_1764 (O_1764,N_18042,N_19074);
and UO_1765 (O_1765,N_18118,N_18115);
or UO_1766 (O_1766,N_18023,N_19355);
or UO_1767 (O_1767,N_19773,N_19059);
or UO_1768 (O_1768,N_18430,N_18728);
nor UO_1769 (O_1769,N_18320,N_19553);
nand UO_1770 (O_1770,N_18713,N_19304);
and UO_1771 (O_1771,N_18313,N_18264);
or UO_1772 (O_1772,N_19567,N_19266);
nand UO_1773 (O_1773,N_19410,N_19002);
nor UO_1774 (O_1774,N_19398,N_19227);
and UO_1775 (O_1775,N_19121,N_18496);
nand UO_1776 (O_1776,N_19793,N_18351);
xnor UO_1777 (O_1777,N_19104,N_18932);
xor UO_1778 (O_1778,N_18112,N_18761);
and UO_1779 (O_1779,N_18690,N_19378);
or UO_1780 (O_1780,N_18681,N_18861);
and UO_1781 (O_1781,N_18368,N_18798);
or UO_1782 (O_1782,N_19476,N_18759);
or UO_1783 (O_1783,N_19694,N_19230);
nand UO_1784 (O_1784,N_19137,N_19802);
and UO_1785 (O_1785,N_18339,N_18217);
xnor UO_1786 (O_1786,N_18004,N_18288);
nor UO_1787 (O_1787,N_19655,N_19977);
xor UO_1788 (O_1788,N_18470,N_18945);
nand UO_1789 (O_1789,N_19229,N_19123);
xnor UO_1790 (O_1790,N_19511,N_18677);
xor UO_1791 (O_1791,N_18586,N_19967);
nand UO_1792 (O_1792,N_18491,N_19761);
and UO_1793 (O_1793,N_19967,N_18841);
nor UO_1794 (O_1794,N_18273,N_18202);
and UO_1795 (O_1795,N_19065,N_19343);
nor UO_1796 (O_1796,N_18746,N_18638);
nor UO_1797 (O_1797,N_19367,N_18235);
nand UO_1798 (O_1798,N_19867,N_18300);
and UO_1799 (O_1799,N_18810,N_18916);
or UO_1800 (O_1800,N_19904,N_19531);
xnor UO_1801 (O_1801,N_19817,N_18034);
nand UO_1802 (O_1802,N_19385,N_19687);
nand UO_1803 (O_1803,N_19762,N_19485);
and UO_1804 (O_1804,N_19608,N_18927);
nor UO_1805 (O_1805,N_18354,N_19270);
or UO_1806 (O_1806,N_19751,N_19858);
and UO_1807 (O_1807,N_19907,N_18359);
xor UO_1808 (O_1808,N_19288,N_18270);
nor UO_1809 (O_1809,N_19869,N_19741);
nor UO_1810 (O_1810,N_19943,N_19602);
nand UO_1811 (O_1811,N_19547,N_18492);
nor UO_1812 (O_1812,N_19405,N_19979);
nor UO_1813 (O_1813,N_18996,N_18096);
xnor UO_1814 (O_1814,N_18975,N_19117);
nor UO_1815 (O_1815,N_18627,N_19580);
or UO_1816 (O_1816,N_18892,N_19679);
or UO_1817 (O_1817,N_18280,N_18625);
nor UO_1818 (O_1818,N_18333,N_19938);
nand UO_1819 (O_1819,N_19528,N_19137);
nor UO_1820 (O_1820,N_19971,N_18538);
and UO_1821 (O_1821,N_19214,N_19641);
and UO_1822 (O_1822,N_19542,N_18451);
nor UO_1823 (O_1823,N_19972,N_19985);
or UO_1824 (O_1824,N_19053,N_18282);
nor UO_1825 (O_1825,N_19359,N_18153);
or UO_1826 (O_1826,N_19429,N_18215);
nand UO_1827 (O_1827,N_18966,N_19874);
and UO_1828 (O_1828,N_19848,N_19524);
nor UO_1829 (O_1829,N_19832,N_19159);
nor UO_1830 (O_1830,N_18098,N_19341);
or UO_1831 (O_1831,N_19503,N_18647);
nand UO_1832 (O_1832,N_19012,N_18272);
and UO_1833 (O_1833,N_18409,N_18464);
nand UO_1834 (O_1834,N_19668,N_18798);
xnor UO_1835 (O_1835,N_18458,N_18973);
nor UO_1836 (O_1836,N_18308,N_19564);
nand UO_1837 (O_1837,N_18724,N_19989);
nor UO_1838 (O_1838,N_19219,N_19167);
or UO_1839 (O_1839,N_19556,N_18167);
nor UO_1840 (O_1840,N_19099,N_18802);
or UO_1841 (O_1841,N_18507,N_18658);
nor UO_1842 (O_1842,N_19963,N_18199);
and UO_1843 (O_1843,N_19864,N_19731);
xor UO_1844 (O_1844,N_19152,N_19112);
or UO_1845 (O_1845,N_19640,N_19988);
and UO_1846 (O_1846,N_19327,N_18051);
xor UO_1847 (O_1847,N_19301,N_18351);
or UO_1848 (O_1848,N_19722,N_18715);
xor UO_1849 (O_1849,N_19194,N_18979);
and UO_1850 (O_1850,N_19423,N_18194);
or UO_1851 (O_1851,N_19868,N_18554);
or UO_1852 (O_1852,N_18980,N_18351);
nor UO_1853 (O_1853,N_18920,N_19406);
nand UO_1854 (O_1854,N_18153,N_19933);
or UO_1855 (O_1855,N_18419,N_19006);
and UO_1856 (O_1856,N_19459,N_18469);
nor UO_1857 (O_1857,N_19810,N_19892);
or UO_1858 (O_1858,N_18564,N_18477);
and UO_1859 (O_1859,N_18014,N_19296);
nand UO_1860 (O_1860,N_19408,N_18395);
or UO_1861 (O_1861,N_19445,N_18408);
or UO_1862 (O_1862,N_18960,N_18518);
and UO_1863 (O_1863,N_19081,N_19321);
or UO_1864 (O_1864,N_19688,N_19771);
and UO_1865 (O_1865,N_19767,N_18164);
and UO_1866 (O_1866,N_19288,N_18825);
nand UO_1867 (O_1867,N_19404,N_18885);
nand UO_1868 (O_1868,N_18017,N_18972);
or UO_1869 (O_1869,N_18837,N_18694);
and UO_1870 (O_1870,N_18406,N_18039);
and UO_1871 (O_1871,N_19556,N_19163);
and UO_1872 (O_1872,N_19051,N_18434);
or UO_1873 (O_1873,N_18904,N_18956);
nor UO_1874 (O_1874,N_19949,N_19051);
nor UO_1875 (O_1875,N_18316,N_19592);
nor UO_1876 (O_1876,N_18458,N_18768);
nand UO_1877 (O_1877,N_18676,N_19379);
nand UO_1878 (O_1878,N_19379,N_18128);
nor UO_1879 (O_1879,N_18620,N_18167);
and UO_1880 (O_1880,N_18035,N_19252);
or UO_1881 (O_1881,N_18346,N_18231);
and UO_1882 (O_1882,N_19072,N_19529);
nor UO_1883 (O_1883,N_19402,N_18075);
and UO_1884 (O_1884,N_18470,N_18200);
and UO_1885 (O_1885,N_18821,N_18622);
nor UO_1886 (O_1886,N_18134,N_18849);
or UO_1887 (O_1887,N_18560,N_18033);
xnor UO_1888 (O_1888,N_19565,N_18894);
and UO_1889 (O_1889,N_18070,N_19227);
xnor UO_1890 (O_1890,N_18509,N_19114);
nand UO_1891 (O_1891,N_18225,N_18600);
xnor UO_1892 (O_1892,N_18216,N_19060);
nor UO_1893 (O_1893,N_19396,N_19447);
xor UO_1894 (O_1894,N_19840,N_19907);
or UO_1895 (O_1895,N_18620,N_18945);
nand UO_1896 (O_1896,N_18415,N_18803);
nor UO_1897 (O_1897,N_19090,N_19097);
xnor UO_1898 (O_1898,N_18040,N_18626);
or UO_1899 (O_1899,N_18203,N_18876);
and UO_1900 (O_1900,N_19490,N_19376);
nand UO_1901 (O_1901,N_18627,N_19259);
nor UO_1902 (O_1902,N_18838,N_18193);
xor UO_1903 (O_1903,N_18243,N_18643);
nand UO_1904 (O_1904,N_18370,N_18417);
nand UO_1905 (O_1905,N_18927,N_18821);
xnor UO_1906 (O_1906,N_19384,N_19510);
nand UO_1907 (O_1907,N_19166,N_19175);
nand UO_1908 (O_1908,N_18192,N_18684);
or UO_1909 (O_1909,N_19846,N_19763);
nand UO_1910 (O_1910,N_19689,N_19313);
nand UO_1911 (O_1911,N_18422,N_19716);
nor UO_1912 (O_1912,N_19256,N_19566);
or UO_1913 (O_1913,N_19113,N_18726);
nand UO_1914 (O_1914,N_19897,N_18153);
and UO_1915 (O_1915,N_19087,N_18876);
nor UO_1916 (O_1916,N_18500,N_18026);
and UO_1917 (O_1917,N_19587,N_18092);
xnor UO_1918 (O_1918,N_19602,N_18091);
or UO_1919 (O_1919,N_19244,N_18120);
or UO_1920 (O_1920,N_18166,N_18181);
or UO_1921 (O_1921,N_18558,N_19832);
nand UO_1922 (O_1922,N_19943,N_18583);
nand UO_1923 (O_1923,N_18633,N_19906);
xnor UO_1924 (O_1924,N_19494,N_18910);
or UO_1925 (O_1925,N_19221,N_18659);
or UO_1926 (O_1926,N_19880,N_19738);
nor UO_1927 (O_1927,N_19545,N_18193);
xnor UO_1928 (O_1928,N_19303,N_19934);
xor UO_1929 (O_1929,N_18899,N_18045);
nor UO_1930 (O_1930,N_19036,N_19216);
nor UO_1931 (O_1931,N_18635,N_19063);
nand UO_1932 (O_1932,N_19851,N_19010);
nand UO_1933 (O_1933,N_18566,N_19758);
nor UO_1934 (O_1934,N_18910,N_19499);
nor UO_1935 (O_1935,N_18353,N_19532);
xor UO_1936 (O_1936,N_18292,N_19808);
or UO_1937 (O_1937,N_19516,N_18694);
nor UO_1938 (O_1938,N_18545,N_19834);
nand UO_1939 (O_1939,N_19705,N_19727);
xor UO_1940 (O_1940,N_19749,N_19441);
or UO_1941 (O_1941,N_18786,N_18498);
nand UO_1942 (O_1942,N_19342,N_19800);
nand UO_1943 (O_1943,N_19772,N_19549);
xnor UO_1944 (O_1944,N_19591,N_18159);
and UO_1945 (O_1945,N_19480,N_18891);
or UO_1946 (O_1946,N_19384,N_18624);
xnor UO_1947 (O_1947,N_19760,N_18451);
and UO_1948 (O_1948,N_19204,N_19116);
or UO_1949 (O_1949,N_19315,N_18841);
xor UO_1950 (O_1950,N_19119,N_18720);
or UO_1951 (O_1951,N_19778,N_19482);
and UO_1952 (O_1952,N_18156,N_18894);
nand UO_1953 (O_1953,N_19748,N_19531);
xor UO_1954 (O_1954,N_18587,N_19473);
or UO_1955 (O_1955,N_19030,N_19486);
and UO_1956 (O_1956,N_19260,N_18108);
xnor UO_1957 (O_1957,N_18152,N_18164);
nand UO_1958 (O_1958,N_18154,N_19446);
and UO_1959 (O_1959,N_18405,N_18903);
or UO_1960 (O_1960,N_19200,N_19413);
and UO_1961 (O_1961,N_18934,N_19942);
and UO_1962 (O_1962,N_18491,N_19795);
and UO_1963 (O_1963,N_18270,N_18085);
or UO_1964 (O_1964,N_19258,N_18606);
nand UO_1965 (O_1965,N_19952,N_19535);
nand UO_1966 (O_1966,N_18515,N_19414);
and UO_1967 (O_1967,N_19471,N_19035);
and UO_1968 (O_1968,N_18487,N_18038);
nor UO_1969 (O_1969,N_18586,N_19429);
and UO_1970 (O_1970,N_19342,N_18164);
and UO_1971 (O_1971,N_18973,N_19570);
or UO_1972 (O_1972,N_19121,N_19531);
or UO_1973 (O_1973,N_18943,N_19653);
nor UO_1974 (O_1974,N_19752,N_19929);
or UO_1975 (O_1975,N_18193,N_18045);
or UO_1976 (O_1976,N_18160,N_19201);
and UO_1977 (O_1977,N_18468,N_19738);
or UO_1978 (O_1978,N_19034,N_18110);
nand UO_1979 (O_1979,N_19944,N_18506);
xnor UO_1980 (O_1980,N_19011,N_19781);
xnor UO_1981 (O_1981,N_18778,N_19386);
xnor UO_1982 (O_1982,N_19487,N_19982);
nand UO_1983 (O_1983,N_18865,N_18971);
or UO_1984 (O_1984,N_19074,N_19841);
or UO_1985 (O_1985,N_18908,N_19846);
and UO_1986 (O_1986,N_19356,N_19335);
or UO_1987 (O_1987,N_18778,N_19416);
nor UO_1988 (O_1988,N_19106,N_19500);
nor UO_1989 (O_1989,N_18550,N_18269);
nor UO_1990 (O_1990,N_19821,N_18837);
xor UO_1991 (O_1991,N_19069,N_18089);
nor UO_1992 (O_1992,N_18249,N_18854);
xor UO_1993 (O_1993,N_19525,N_19072);
and UO_1994 (O_1994,N_18235,N_18375);
nand UO_1995 (O_1995,N_19308,N_18146);
nand UO_1996 (O_1996,N_19061,N_18052);
and UO_1997 (O_1997,N_19690,N_19975);
nand UO_1998 (O_1998,N_18802,N_19573);
and UO_1999 (O_1999,N_19099,N_19160);
or UO_2000 (O_2000,N_19215,N_18919);
nor UO_2001 (O_2001,N_19052,N_19575);
xor UO_2002 (O_2002,N_18071,N_19432);
nand UO_2003 (O_2003,N_19742,N_19737);
xnor UO_2004 (O_2004,N_18124,N_18029);
nor UO_2005 (O_2005,N_18448,N_19357);
and UO_2006 (O_2006,N_19676,N_18472);
and UO_2007 (O_2007,N_19908,N_18838);
or UO_2008 (O_2008,N_19298,N_19990);
nand UO_2009 (O_2009,N_18811,N_19649);
and UO_2010 (O_2010,N_19714,N_18335);
nor UO_2011 (O_2011,N_19571,N_18390);
xnor UO_2012 (O_2012,N_19587,N_18351);
nor UO_2013 (O_2013,N_18030,N_19755);
nor UO_2014 (O_2014,N_19276,N_18531);
xnor UO_2015 (O_2015,N_19748,N_19814);
nor UO_2016 (O_2016,N_18035,N_19094);
and UO_2017 (O_2017,N_18115,N_18777);
or UO_2018 (O_2018,N_19282,N_18533);
and UO_2019 (O_2019,N_18172,N_18301);
and UO_2020 (O_2020,N_19382,N_18462);
xnor UO_2021 (O_2021,N_18009,N_18499);
or UO_2022 (O_2022,N_19779,N_19684);
xnor UO_2023 (O_2023,N_19478,N_18887);
and UO_2024 (O_2024,N_19443,N_18957);
xnor UO_2025 (O_2025,N_18460,N_19201);
or UO_2026 (O_2026,N_18937,N_19161);
or UO_2027 (O_2027,N_18670,N_19011);
nand UO_2028 (O_2028,N_18125,N_18630);
nor UO_2029 (O_2029,N_19190,N_19292);
or UO_2030 (O_2030,N_19024,N_18180);
nand UO_2031 (O_2031,N_19556,N_19356);
and UO_2032 (O_2032,N_19566,N_19027);
or UO_2033 (O_2033,N_18654,N_19797);
xor UO_2034 (O_2034,N_19283,N_19816);
and UO_2035 (O_2035,N_18363,N_18986);
nand UO_2036 (O_2036,N_18204,N_19158);
and UO_2037 (O_2037,N_19504,N_18528);
nand UO_2038 (O_2038,N_18025,N_18658);
nand UO_2039 (O_2039,N_19464,N_19134);
nor UO_2040 (O_2040,N_19945,N_18123);
and UO_2041 (O_2041,N_18933,N_18948);
xor UO_2042 (O_2042,N_19816,N_19783);
nor UO_2043 (O_2043,N_18731,N_19981);
nand UO_2044 (O_2044,N_19845,N_19803);
or UO_2045 (O_2045,N_18792,N_19238);
and UO_2046 (O_2046,N_19391,N_18155);
nor UO_2047 (O_2047,N_18013,N_18076);
and UO_2048 (O_2048,N_19477,N_18810);
nor UO_2049 (O_2049,N_19812,N_18238);
xnor UO_2050 (O_2050,N_18708,N_18480);
or UO_2051 (O_2051,N_19120,N_18070);
nand UO_2052 (O_2052,N_19585,N_18066);
or UO_2053 (O_2053,N_18559,N_19862);
or UO_2054 (O_2054,N_19010,N_18785);
and UO_2055 (O_2055,N_19744,N_19768);
and UO_2056 (O_2056,N_19380,N_18415);
nand UO_2057 (O_2057,N_18872,N_19542);
or UO_2058 (O_2058,N_19546,N_18854);
and UO_2059 (O_2059,N_19577,N_19097);
or UO_2060 (O_2060,N_18583,N_18691);
nand UO_2061 (O_2061,N_19026,N_19913);
xor UO_2062 (O_2062,N_19031,N_18506);
xnor UO_2063 (O_2063,N_19276,N_19661);
or UO_2064 (O_2064,N_19976,N_19837);
and UO_2065 (O_2065,N_19932,N_19640);
nor UO_2066 (O_2066,N_18193,N_19628);
nor UO_2067 (O_2067,N_19482,N_18330);
nand UO_2068 (O_2068,N_19471,N_19458);
nand UO_2069 (O_2069,N_19533,N_19482);
xor UO_2070 (O_2070,N_18887,N_18055);
or UO_2071 (O_2071,N_18361,N_18672);
nand UO_2072 (O_2072,N_18575,N_19494);
and UO_2073 (O_2073,N_19875,N_18599);
or UO_2074 (O_2074,N_19815,N_19475);
and UO_2075 (O_2075,N_18102,N_18591);
or UO_2076 (O_2076,N_18395,N_19304);
or UO_2077 (O_2077,N_19226,N_19253);
nand UO_2078 (O_2078,N_19454,N_19591);
and UO_2079 (O_2079,N_18559,N_19154);
nor UO_2080 (O_2080,N_18923,N_18382);
or UO_2081 (O_2081,N_19541,N_18078);
xnor UO_2082 (O_2082,N_19931,N_19401);
and UO_2083 (O_2083,N_18271,N_19995);
or UO_2084 (O_2084,N_18365,N_19160);
or UO_2085 (O_2085,N_18088,N_18498);
xnor UO_2086 (O_2086,N_18628,N_18491);
nor UO_2087 (O_2087,N_19659,N_19069);
nor UO_2088 (O_2088,N_18224,N_19192);
nand UO_2089 (O_2089,N_19736,N_19893);
and UO_2090 (O_2090,N_18130,N_18652);
nand UO_2091 (O_2091,N_19259,N_18918);
nor UO_2092 (O_2092,N_18039,N_18741);
xor UO_2093 (O_2093,N_18508,N_18533);
or UO_2094 (O_2094,N_19430,N_18160);
nand UO_2095 (O_2095,N_19860,N_19398);
or UO_2096 (O_2096,N_18419,N_19654);
nand UO_2097 (O_2097,N_19326,N_19296);
nand UO_2098 (O_2098,N_18251,N_18661);
or UO_2099 (O_2099,N_18996,N_18510);
and UO_2100 (O_2100,N_19071,N_18284);
xnor UO_2101 (O_2101,N_19020,N_19375);
and UO_2102 (O_2102,N_19945,N_18138);
nor UO_2103 (O_2103,N_18218,N_18229);
nor UO_2104 (O_2104,N_19600,N_19232);
nand UO_2105 (O_2105,N_18661,N_19823);
nand UO_2106 (O_2106,N_19915,N_19818);
nor UO_2107 (O_2107,N_18532,N_18859);
and UO_2108 (O_2108,N_18526,N_19733);
or UO_2109 (O_2109,N_19454,N_19146);
xor UO_2110 (O_2110,N_19952,N_19206);
or UO_2111 (O_2111,N_18960,N_19145);
xnor UO_2112 (O_2112,N_18861,N_18423);
and UO_2113 (O_2113,N_18699,N_19846);
or UO_2114 (O_2114,N_18853,N_18905);
and UO_2115 (O_2115,N_18645,N_18883);
and UO_2116 (O_2116,N_18851,N_18996);
and UO_2117 (O_2117,N_19764,N_18825);
and UO_2118 (O_2118,N_19511,N_18433);
nor UO_2119 (O_2119,N_19438,N_19259);
nand UO_2120 (O_2120,N_18963,N_18683);
and UO_2121 (O_2121,N_19501,N_18226);
or UO_2122 (O_2122,N_19283,N_19971);
and UO_2123 (O_2123,N_18857,N_18874);
nand UO_2124 (O_2124,N_18098,N_18356);
xnor UO_2125 (O_2125,N_19260,N_18489);
xor UO_2126 (O_2126,N_19927,N_18587);
or UO_2127 (O_2127,N_19522,N_19354);
nor UO_2128 (O_2128,N_19563,N_18184);
xnor UO_2129 (O_2129,N_18478,N_18903);
xnor UO_2130 (O_2130,N_19650,N_19136);
and UO_2131 (O_2131,N_18363,N_18873);
and UO_2132 (O_2132,N_19578,N_18911);
nand UO_2133 (O_2133,N_19010,N_19507);
xnor UO_2134 (O_2134,N_19934,N_19058);
and UO_2135 (O_2135,N_18801,N_19331);
and UO_2136 (O_2136,N_19087,N_18577);
xnor UO_2137 (O_2137,N_19841,N_18308);
xnor UO_2138 (O_2138,N_18330,N_18903);
nand UO_2139 (O_2139,N_19778,N_18681);
or UO_2140 (O_2140,N_19808,N_19811);
and UO_2141 (O_2141,N_18844,N_18678);
nor UO_2142 (O_2142,N_18879,N_19802);
nor UO_2143 (O_2143,N_19258,N_18861);
nand UO_2144 (O_2144,N_19726,N_19041);
nand UO_2145 (O_2145,N_18406,N_19619);
or UO_2146 (O_2146,N_19181,N_18647);
nor UO_2147 (O_2147,N_18604,N_19761);
or UO_2148 (O_2148,N_18382,N_18765);
nand UO_2149 (O_2149,N_19006,N_19165);
or UO_2150 (O_2150,N_18815,N_18372);
nor UO_2151 (O_2151,N_18473,N_19144);
xnor UO_2152 (O_2152,N_18061,N_18874);
xnor UO_2153 (O_2153,N_19986,N_19530);
and UO_2154 (O_2154,N_18667,N_18257);
xor UO_2155 (O_2155,N_19597,N_19509);
nor UO_2156 (O_2156,N_18061,N_18279);
xnor UO_2157 (O_2157,N_18828,N_19328);
or UO_2158 (O_2158,N_18251,N_18981);
or UO_2159 (O_2159,N_18911,N_19515);
nand UO_2160 (O_2160,N_19689,N_18014);
nor UO_2161 (O_2161,N_19949,N_18479);
nand UO_2162 (O_2162,N_18811,N_18709);
nand UO_2163 (O_2163,N_19887,N_19688);
or UO_2164 (O_2164,N_19521,N_18176);
xnor UO_2165 (O_2165,N_18930,N_19126);
and UO_2166 (O_2166,N_19695,N_19456);
xor UO_2167 (O_2167,N_19894,N_19194);
nor UO_2168 (O_2168,N_18200,N_19675);
nand UO_2169 (O_2169,N_19451,N_18946);
or UO_2170 (O_2170,N_18190,N_19070);
nand UO_2171 (O_2171,N_18144,N_18326);
nor UO_2172 (O_2172,N_19236,N_19992);
or UO_2173 (O_2173,N_18983,N_18065);
xor UO_2174 (O_2174,N_18261,N_19122);
or UO_2175 (O_2175,N_18243,N_19906);
or UO_2176 (O_2176,N_19474,N_18070);
nor UO_2177 (O_2177,N_19072,N_19477);
nor UO_2178 (O_2178,N_18212,N_19384);
or UO_2179 (O_2179,N_18343,N_19140);
or UO_2180 (O_2180,N_18409,N_18152);
nand UO_2181 (O_2181,N_19321,N_18953);
nand UO_2182 (O_2182,N_19357,N_18660);
and UO_2183 (O_2183,N_19714,N_18273);
or UO_2184 (O_2184,N_19894,N_19089);
and UO_2185 (O_2185,N_18455,N_18681);
xnor UO_2186 (O_2186,N_19638,N_19218);
and UO_2187 (O_2187,N_19002,N_19846);
nand UO_2188 (O_2188,N_18516,N_19953);
or UO_2189 (O_2189,N_18130,N_19228);
or UO_2190 (O_2190,N_19869,N_18641);
nand UO_2191 (O_2191,N_19076,N_18289);
nand UO_2192 (O_2192,N_18245,N_19892);
nor UO_2193 (O_2193,N_19971,N_19402);
nor UO_2194 (O_2194,N_18963,N_19337);
and UO_2195 (O_2195,N_18299,N_18328);
or UO_2196 (O_2196,N_19227,N_19662);
and UO_2197 (O_2197,N_19015,N_19638);
nor UO_2198 (O_2198,N_18485,N_19034);
or UO_2199 (O_2199,N_18549,N_18804);
or UO_2200 (O_2200,N_18059,N_18925);
xor UO_2201 (O_2201,N_19982,N_19459);
nand UO_2202 (O_2202,N_18587,N_19996);
xor UO_2203 (O_2203,N_19702,N_18191);
nand UO_2204 (O_2204,N_19614,N_18909);
or UO_2205 (O_2205,N_18374,N_18812);
nor UO_2206 (O_2206,N_19549,N_19057);
and UO_2207 (O_2207,N_18270,N_19263);
nand UO_2208 (O_2208,N_19828,N_19385);
or UO_2209 (O_2209,N_18154,N_18747);
nand UO_2210 (O_2210,N_19869,N_18003);
xnor UO_2211 (O_2211,N_18958,N_18459);
and UO_2212 (O_2212,N_19212,N_19750);
nand UO_2213 (O_2213,N_19638,N_18698);
and UO_2214 (O_2214,N_19587,N_19800);
nand UO_2215 (O_2215,N_19805,N_18579);
xor UO_2216 (O_2216,N_18887,N_19765);
or UO_2217 (O_2217,N_19899,N_19556);
and UO_2218 (O_2218,N_19493,N_19954);
nand UO_2219 (O_2219,N_18472,N_19519);
or UO_2220 (O_2220,N_18862,N_18395);
and UO_2221 (O_2221,N_19269,N_19902);
nand UO_2222 (O_2222,N_18379,N_19437);
or UO_2223 (O_2223,N_18229,N_19901);
nor UO_2224 (O_2224,N_18481,N_18978);
xor UO_2225 (O_2225,N_18449,N_18136);
xor UO_2226 (O_2226,N_19553,N_19839);
nand UO_2227 (O_2227,N_18559,N_18521);
and UO_2228 (O_2228,N_19695,N_18798);
nand UO_2229 (O_2229,N_18345,N_18683);
and UO_2230 (O_2230,N_18133,N_18413);
or UO_2231 (O_2231,N_19036,N_18935);
or UO_2232 (O_2232,N_19148,N_18992);
and UO_2233 (O_2233,N_19940,N_18873);
xor UO_2234 (O_2234,N_18090,N_18177);
nand UO_2235 (O_2235,N_19965,N_19322);
xnor UO_2236 (O_2236,N_19242,N_18637);
nand UO_2237 (O_2237,N_19384,N_18350);
nand UO_2238 (O_2238,N_19746,N_18240);
and UO_2239 (O_2239,N_18234,N_19039);
and UO_2240 (O_2240,N_18894,N_18945);
nor UO_2241 (O_2241,N_18303,N_19240);
and UO_2242 (O_2242,N_19459,N_18429);
and UO_2243 (O_2243,N_18492,N_19047);
nand UO_2244 (O_2244,N_18328,N_19789);
nand UO_2245 (O_2245,N_19693,N_18655);
nand UO_2246 (O_2246,N_19317,N_19993);
or UO_2247 (O_2247,N_19820,N_18032);
nand UO_2248 (O_2248,N_19401,N_18134);
or UO_2249 (O_2249,N_18791,N_19256);
or UO_2250 (O_2250,N_19688,N_19432);
xor UO_2251 (O_2251,N_19678,N_18177);
or UO_2252 (O_2252,N_19621,N_18138);
or UO_2253 (O_2253,N_19259,N_18026);
and UO_2254 (O_2254,N_18650,N_19818);
nor UO_2255 (O_2255,N_18804,N_18181);
xor UO_2256 (O_2256,N_19183,N_18352);
or UO_2257 (O_2257,N_19415,N_18307);
xor UO_2258 (O_2258,N_19232,N_18879);
or UO_2259 (O_2259,N_19121,N_19254);
xor UO_2260 (O_2260,N_18427,N_18250);
nor UO_2261 (O_2261,N_19739,N_19764);
xor UO_2262 (O_2262,N_18304,N_18750);
or UO_2263 (O_2263,N_19242,N_19965);
and UO_2264 (O_2264,N_19382,N_18918);
nand UO_2265 (O_2265,N_18216,N_18181);
or UO_2266 (O_2266,N_18298,N_19938);
nor UO_2267 (O_2267,N_18490,N_18369);
xnor UO_2268 (O_2268,N_19431,N_18311);
nand UO_2269 (O_2269,N_18947,N_18910);
or UO_2270 (O_2270,N_19129,N_18154);
nor UO_2271 (O_2271,N_19644,N_19447);
and UO_2272 (O_2272,N_18421,N_18954);
nand UO_2273 (O_2273,N_18406,N_19520);
or UO_2274 (O_2274,N_19853,N_19924);
nor UO_2275 (O_2275,N_19984,N_18492);
and UO_2276 (O_2276,N_18049,N_19592);
or UO_2277 (O_2277,N_19265,N_19845);
nor UO_2278 (O_2278,N_18010,N_18948);
or UO_2279 (O_2279,N_19945,N_18507);
xor UO_2280 (O_2280,N_18216,N_19523);
nor UO_2281 (O_2281,N_18651,N_19574);
nand UO_2282 (O_2282,N_18262,N_18106);
and UO_2283 (O_2283,N_19797,N_18144);
and UO_2284 (O_2284,N_18586,N_18542);
or UO_2285 (O_2285,N_19599,N_19472);
or UO_2286 (O_2286,N_19255,N_19463);
nand UO_2287 (O_2287,N_18610,N_19822);
nor UO_2288 (O_2288,N_18808,N_19540);
and UO_2289 (O_2289,N_19898,N_18000);
nand UO_2290 (O_2290,N_19465,N_18495);
nand UO_2291 (O_2291,N_18199,N_19801);
xnor UO_2292 (O_2292,N_18456,N_18581);
and UO_2293 (O_2293,N_18491,N_19908);
and UO_2294 (O_2294,N_18410,N_18140);
nand UO_2295 (O_2295,N_19919,N_19477);
nand UO_2296 (O_2296,N_18274,N_18116);
nand UO_2297 (O_2297,N_18956,N_18240);
xnor UO_2298 (O_2298,N_19994,N_19558);
nand UO_2299 (O_2299,N_19035,N_19085);
nor UO_2300 (O_2300,N_18071,N_18913);
or UO_2301 (O_2301,N_18236,N_18779);
or UO_2302 (O_2302,N_19075,N_19541);
nor UO_2303 (O_2303,N_18560,N_19620);
or UO_2304 (O_2304,N_19347,N_19436);
or UO_2305 (O_2305,N_19096,N_19355);
nor UO_2306 (O_2306,N_19247,N_19342);
xor UO_2307 (O_2307,N_18115,N_19569);
or UO_2308 (O_2308,N_19840,N_18909);
xor UO_2309 (O_2309,N_18821,N_18882);
nand UO_2310 (O_2310,N_19697,N_19857);
or UO_2311 (O_2311,N_19488,N_18892);
nor UO_2312 (O_2312,N_18497,N_18767);
or UO_2313 (O_2313,N_18481,N_19767);
nor UO_2314 (O_2314,N_18337,N_19490);
nor UO_2315 (O_2315,N_19123,N_18653);
nand UO_2316 (O_2316,N_19760,N_19746);
nand UO_2317 (O_2317,N_19068,N_19376);
nand UO_2318 (O_2318,N_19991,N_19105);
xnor UO_2319 (O_2319,N_18910,N_19279);
and UO_2320 (O_2320,N_19026,N_18474);
nand UO_2321 (O_2321,N_18609,N_19272);
xnor UO_2322 (O_2322,N_19132,N_19676);
xnor UO_2323 (O_2323,N_18725,N_18258);
and UO_2324 (O_2324,N_18092,N_18272);
nor UO_2325 (O_2325,N_18354,N_18035);
nand UO_2326 (O_2326,N_18617,N_18994);
nand UO_2327 (O_2327,N_18574,N_18879);
and UO_2328 (O_2328,N_19464,N_18768);
or UO_2329 (O_2329,N_18771,N_19751);
xor UO_2330 (O_2330,N_19380,N_19854);
or UO_2331 (O_2331,N_19540,N_18527);
and UO_2332 (O_2332,N_18492,N_18103);
nor UO_2333 (O_2333,N_18616,N_18240);
nand UO_2334 (O_2334,N_19974,N_19603);
nand UO_2335 (O_2335,N_18962,N_18806);
or UO_2336 (O_2336,N_18114,N_19244);
nand UO_2337 (O_2337,N_19200,N_18142);
or UO_2338 (O_2338,N_19659,N_19063);
or UO_2339 (O_2339,N_19696,N_19891);
xor UO_2340 (O_2340,N_19088,N_19651);
or UO_2341 (O_2341,N_18996,N_18811);
xor UO_2342 (O_2342,N_18938,N_19178);
or UO_2343 (O_2343,N_19784,N_18909);
or UO_2344 (O_2344,N_19699,N_19702);
nand UO_2345 (O_2345,N_19483,N_19068);
nor UO_2346 (O_2346,N_19813,N_18323);
nor UO_2347 (O_2347,N_19211,N_18853);
or UO_2348 (O_2348,N_18906,N_19008);
and UO_2349 (O_2349,N_19352,N_18793);
nand UO_2350 (O_2350,N_19537,N_19438);
xor UO_2351 (O_2351,N_19319,N_19334);
nor UO_2352 (O_2352,N_19245,N_18903);
xnor UO_2353 (O_2353,N_18857,N_18708);
nand UO_2354 (O_2354,N_18230,N_19718);
and UO_2355 (O_2355,N_19531,N_19543);
nor UO_2356 (O_2356,N_19572,N_19918);
or UO_2357 (O_2357,N_18405,N_18441);
nor UO_2358 (O_2358,N_19247,N_19091);
nand UO_2359 (O_2359,N_19524,N_19496);
nand UO_2360 (O_2360,N_18291,N_19168);
or UO_2361 (O_2361,N_19420,N_19510);
or UO_2362 (O_2362,N_18093,N_18346);
and UO_2363 (O_2363,N_18447,N_18775);
xor UO_2364 (O_2364,N_18887,N_18474);
and UO_2365 (O_2365,N_18413,N_18567);
and UO_2366 (O_2366,N_19167,N_18354);
xnor UO_2367 (O_2367,N_18763,N_19878);
nand UO_2368 (O_2368,N_19684,N_19338);
xnor UO_2369 (O_2369,N_18813,N_19783);
nand UO_2370 (O_2370,N_18262,N_18228);
and UO_2371 (O_2371,N_18328,N_19906);
nand UO_2372 (O_2372,N_19952,N_18032);
and UO_2373 (O_2373,N_18274,N_18723);
nor UO_2374 (O_2374,N_19500,N_18364);
and UO_2375 (O_2375,N_18874,N_19757);
nand UO_2376 (O_2376,N_18371,N_18290);
nand UO_2377 (O_2377,N_18966,N_18908);
nor UO_2378 (O_2378,N_19283,N_19132);
nor UO_2379 (O_2379,N_19357,N_19211);
xnor UO_2380 (O_2380,N_19358,N_18789);
nand UO_2381 (O_2381,N_19019,N_19301);
nor UO_2382 (O_2382,N_18413,N_18148);
and UO_2383 (O_2383,N_19468,N_18068);
xor UO_2384 (O_2384,N_19957,N_18063);
xnor UO_2385 (O_2385,N_18486,N_18878);
or UO_2386 (O_2386,N_19298,N_19309);
and UO_2387 (O_2387,N_19083,N_19708);
or UO_2388 (O_2388,N_18836,N_19060);
nor UO_2389 (O_2389,N_18541,N_18834);
xor UO_2390 (O_2390,N_18417,N_18214);
or UO_2391 (O_2391,N_18653,N_19632);
nand UO_2392 (O_2392,N_18548,N_19964);
xnor UO_2393 (O_2393,N_19586,N_18645);
and UO_2394 (O_2394,N_19190,N_18480);
nor UO_2395 (O_2395,N_19111,N_19057);
or UO_2396 (O_2396,N_19587,N_18837);
and UO_2397 (O_2397,N_19816,N_18661);
nor UO_2398 (O_2398,N_18588,N_18518);
xor UO_2399 (O_2399,N_19645,N_18398);
xor UO_2400 (O_2400,N_18807,N_18641);
or UO_2401 (O_2401,N_18257,N_19192);
nor UO_2402 (O_2402,N_18755,N_18253);
nor UO_2403 (O_2403,N_19367,N_19474);
or UO_2404 (O_2404,N_18977,N_19176);
nand UO_2405 (O_2405,N_19602,N_18878);
xnor UO_2406 (O_2406,N_19434,N_18059);
or UO_2407 (O_2407,N_19819,N_19726);
and UO_2408 (O_2408,N_18922,N_19142);
nor UO_2409 (O_2409,N_19703,N_19696);
or UO_2410 (O_2410,N_18547,N_18683);
nand UO_2411 (O_2411,N_19250,N_18515);
xnor UO_2412 (O_2412,N_19208,N_18540);
nand UO_2413 (O_2413,N_18378,N_19575);
nand UO_2414 (O_2414,N_19271,N_18126);
nor UO_2415 (O_2415,N_18923,N_19807);
and UO_2416 (O_2416,N_19878,N_18318);
nor UO_2417 (O_2417,N_18718,N_18142);
nor UO_2418 (O_2418,N_18987,N_18759);
xnor UO_2419 (O_2419,N_19856,N_19271);
xnor UO_2420 (O_2420,N_18433,N_18223);
nand UO_2421 (O_2421,N_19509,N_19355);
and UO_2422 (O_2422,N_19307,N_19886);
nor UO_2423 (O_2423,N_19384,N_18261);
or UO_2424 (O_2424,N_19526,N_19069);
nand UO_2425 (O_2425,N_19009,N_19316);
xor UO_2426 (O_2426,N_19650,N_19317);
nand UO_2427 (O_2427,N_18379,N_18859);
nor UO_2428 (O_2428,N_19630,N_18260);
and UO_2429 (O_2429,N_19327,N_18827);
nand UO_2430 (O_2430,N_19875,N_18139);
nor UO_2431 (O_2431,N_18996,N_18617);
and UO_2432 (O_2432,N_18516,N_19146);
and UO_2433 (O_2433,N_18138,N_18170);
nor UO_2434 (O_2434,N_18003,N_18152);
nand UO_2435 (O_2435,N_18302,N_19988);
or UO_2436 (O_2436,N_18100,N_18046);
and UO_2437 (O_2437,N_18286,N_19061);
xnor UO_2438 (O_2438,N_19860,N_18039);
xor UO_2439 (O_2439,N_19431,N_18566);
nor UO_2440 (O_2440,N_19291,N_19932);
or UO_2441 (O_2441,N_18825,N_18096);
and UO_2442 (O_2442,N_19399,N_19220);
or UO_2443 (O_2443,N_18467,N_18651);
or UO_2444 (O_2444,N_19043,N_19675);
or UO_2445 (O_2445,N_18388,N_19679);
xor UO_2446 (O_2446,N_19805,N_18704);
nand UO_2447 (O_2447,N_19618,N_18249);
nand UO_2448 (O_2448,N_19386,N_18911);
and UO_2449 (O_2449,N_19937,N_19390);
and UO_2450 (O_2450,N_18137,N_18491);
nand UO_2451 (O_2451,N_18605,N_19868);
xnor UO_2452 (O_2452,N_19012,N_18665);
nor UO_2453 (O_2453,N_18323,N_18337);
or UO_2454 (O_2454,N_19367,N_18366);
or UO_2455 (O_2455,N_19732,N_18151);
or UO_2456 (O_2456,N_18581,N_18831);
and UO_2457 (O_2457,N_19080,N_18350);
nor UO_2458 (O_2458,N_19407,N_19532);
xnor UO_2459 (O_2459,N_18649,N_19621);
and UO_2460 (O_2460,N_18467,N_19212);
or UO_2461 (O_2461,N_18563,N_19584);
or UO_2462 (O_2462,N_19960,N_19562);
and UO_2463 (O_2463,N_18211,N_18143);
nor UO_2464 (O_2464,N_18362,N_18881);
or UO_2465 (O_2465,N_19510,N_19690);
nor UO_2466 (O_2466,N_19056,N_18665);
xor UO_2467 (O_2467,N_19889,N_18716);
or UO_2468 (O_2468,N_19858,N_19494);
nand UO_2469 (O_2469,N_18569,N_18906);
nor UO_2470 (O_2470,N_18195,N_18505);
xor UO_2471 (O_2471,N_18549,N_18722);
or UO_2472 (O_2472,N_18046,N_19858);
and UO_2473 (O_2473,N_18601,N_19119);
and UO_2474 (O_2474,N_19221,N_18593);
xnor UO_2475 (O_2475,N_18241,N_19159);
nand UO_2476 (O_2476,N_18208,N_19905);
and UO_2477 (O_2477,N_19366,N_18617);
nor UO_2478 (O_2478,N_19657,N_19572);
xnor UO_2479 (O_2479,N_19978,N_19933);
or UO_2480 (O_2480,N_18185,N_18085);
nor UO_2481 (O_2481,N_18661,N_18856);
nor UO_2482 (O_2482,N_19017,N_19861);
nor UO_2483 (O_2483,N_18406,N_18509);
xnor UO_2484 (O_2484,N_19547,N_19407);
and UO_2485 (O_2485,N_18101,N_19468);
or UO_2486 (O_2486,N_18920,N_18830);
and UO_2487 (O_2487,N_19861,N_18215);
or UO_2488 (O_2488,N_18907,N_18394);
and UO_2489 (O_2489,N_18810,N_19698);
xnor UO_2490 (O_2490,N_19428,N_18987);
xnor UO_2491 (O_2491,N_18849,N_19520);
xnor UO_2492 (O_2492,N_19349,N_19345);
nor UO_2493 (O_2493,N_18053,N_18845);
nand UO_2494 (O_2494,N_18275,N_19140);
and UO_2495 (O_2495,N_19724,N_19561);
nand UO_2496 (O_2496,N_19987,N_19994);
nor UO_2497 (O_2497,N_18510,N_19535);
nor UO_2498 (O_2498,N_19836,N_19474);
xnor UO_2499 (O_2499,N_18906,N_19628);
endmodule