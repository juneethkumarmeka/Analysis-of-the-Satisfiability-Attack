module basic_750_5000_1000_10_levels_1xor_9(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999;
or U0 (N_0,In_21,In_517);
or U1 (N_1,In_172,In_327);
nor U2 (N_2,In_705,In_649);
nand U3 (N_3,In_134,In_632);
nor U4 (N_4,In_611,In_371);
nor U5 (N_5,In_579,In_309);
nand U6 (N_6,In_616,In_137);
and U7 (N_7,In_56,In_426);
and U8 (N_8,In_532,In_477);
or U9 (N_9,In_476,In_293);
nand U10 (N_10,In_394,In_166);
nor U11 (N_11,In_332,In_279);
nand U12 (N_12,In_334,In_355);
nor U13 (N_13,In_229,In_40);
and U14 (N_14,In_523,In_231);
and U15 (N_15,In_31,In_527);
nor U16 (N_16,In_190,In_438);
nand U17 (N_17,In_429,In_609);
nand U18 (N_18,In_299,In_41);
and U19 (N_19,In_153,In_151);
and U20 (N_20,In_533,In_124);
nand U21 (N_21,In_487,In_553);
nand U22 (N_22,In_159,In_135);
nand U23 (N_23,In_602,In_681);
nor U24 (N_24,In_749,In_544);
nand U25 (N_25,In_294,In_490);
and U26 (N_26,In_635,In_526);
nor U27 (N_27,In_433,In_715);
nor U28 (N_28,In_703,In_312);
and U29 (N_29,In_746,In_621);
nor U30 (N_30,In_83,In_741);
nor U31 (N_31,In_434,In_292);
or U32 (N_32,In_23,In_317);
and U33 (N_33,In_641,In_217);
or U34 (N_34,In_674,In_634);
nand U35 (N_35,In_591,In_670);
or U36 (N_36,In_604,In_499);
and U37 (N_37,In_223,In_211);
nor U38 (N_38,In_492,In_330);
nand U39 (N_39,In_362,In_111);
nand U40 (N_40,In_745,In_64);
nor U41 (N_41,In_640,In_685);
or U42 (N_42,In_561,In_451);
nand U43 (N_43,In_558,In_38);
and U44 (N_44,In_704,In_677);
nor U45 (N_45,In_37,In_197);
nor U46 (N_46,In_315,In_306);
or U47 (N_47,In_186,In_267);
nand U48 (N_48,In_511,In_183);
nand U49 (N_49,In_208,In_418);
and U50 (N_50,In_264,In_243);
and U51 (N_51,In_732,In_97);
and U52 (N_52,In_198,In_385);
nor U53 (N_53,In_303,In_207);
nand U54 (N_54,In_78,In_592);
nand U55 (N_55,In_503,In_248);
or U56 (N_56,In_210,In_214);
nand U57 (N_57,In_324,In_227);
nor U58 (N_58,In_285,In_743);
or U59 (N_59,In_106,In_174);
and U60 (N_60,In_67,In_199);
nand U61 (N_61,In_577,In_466);
nor U62 (N_62,In_179,In_141);
nand U63 (N_63,In_564,In_431);
or U64 (N_64,In_373,In_475);
nand U65 (N_65,In_417,In_59);
and U66 (N_66,In_252,In_610);
nor U67 (N_67,In_486,In_667);
nor U68 (N_68,In_180,In_288);
and U69 (N_69,In_716,In_540);
nand U70 (N_70,In_238,In_201);
nor U71 (N_71,In_125,In_286);
nand U72 (N_72,In_349,In_10);
nand U73 (N_73,In_614,In_74);
and U74 (N_74,In_284,In_679);
nand U75 (N_75,In_557,In_206);
nand U76 (N_76,In_298,In_550);
nor U77 (N_77,In_96,In_444);
and U78 (N_78,In_268,In_407);
nand U79 (N_79,In_689,In_209);
and U80 (N_80,In_363,In_421);
nor U81 (N_81,In_571,In_430);
and U82 (N_82,In_615,In_542);
and U83 (N_83,In_569,In_622);
and U84 (N_84,In_529,In_545);
or U85 (N_85,In_383,In_501);
and U86 (N_86,In_627,In_608);
or U87 (N_87,In_521,In_226);
or U88 (N_88,In_247,In_404);
nor U89 (N_89,In_682,In_695);
and U90 (N_90,In_427,In_436);
and U91 (N_91,In_218,In_687);
nand U92 (N_92,In_414,In_702);
nand U93 (N_93,In_193,In_375);
or U94 (N_94,In_272,In_711);
or U95 (N_95,In_489,In_628);
and U96 (N_96,In_655,In_54);
nand U97 (N_97,In_20,In_601);
nand U98 (N_98,In_559,In_18);
nand U99 (N_99,In_405,In_391);
nand U100 (N_100,In_603,In_381);
or U101 (N_101,In_344,In_386);
nand U102 (N_102,In_388,In_566);
nand U103 (N_103,In_713,In_578);
nor U104 (N_104,In_519,In_524);
nand U105 (N_105,In_296,In_321);
nand U106 (N_106,In_255,In_43);
and U107 (N_107,In_496,In_335);
or U108 (N_108,In_63,In_563);
nand U109 (N_109,In_234,In_108);
or U110 (N_110,In_618,In_422);
nand U111 (N_111,In_650,In_484);
and U112 (N_112,In_28,In_465);
and U113 (N_113,In_26,In_360);
nand U114 (N_114,In_378,In_707);
nor U115 (N_115,In_379,In_395);
or U116 (N_116,In_352,In_177);
nand U117 (N_117,In_68,In_232);
nor U118 (N_118,In_338,In_12);
nand U119 (N_119,In_259,In_244);
nand U120 (N_120,In_122,In_437);
or U121 (N_121,In_361,In_187);
nand U122 (N_122,In_318,In_175);
nor U123 (N_123,In_301,In_380);
and U124 (N_124,In_195,In_7);
or U125 (N_125,In_428,In_680);
and U126 (N_126,In_441,In_205);
or U127 (N_127,In_498,In_246);
nor U128 (N_128,In_495,In_130);
nor U129 (N_129,In_42,In_514);
nand U130 (N_130,In_192,In_353);
nor U131 (N_131,In_95,In_277);
or U132 (N_132,In_710,In_712);
nand U133 (N_133,In_581,In_138);
and U134 (N_134,In_115,In_204);
and U135 (N_135,In_52,In_4);
and U136 (N_136,In_291,In_365);
nand U137 (N_137,In_188,In_552);
nand U138 (N_138,In_683,In_402);
nand U139 (N_139,In_637,In_302);
and U140 (N_140,In_88,In_189);
or U141 (N_141,In_176,In_154);
and U142 (N_142,In_9,In_148);
nand U143 (N_143,In_387,In_194);
and U144 (N_144,In_636,In_150);
nand U145 (N_145,In_358,In_722);
nor U146 (N_146,In_403,In_15);
or U147 (N_147,In_737,In_401);
nand U148 (N_148,In_350,In_399);
or U149 (N_149,In_225,In_598);
and U150 (N_150,In_432,In_528);
and U151 (N_151,In_121,In_516);
nor U152 (N_152,In_522,In_510);
xor U153 (N_153,In_657,In_734);
or U154 (N_154,In_376,In_480);
nor U155 (N_155,In_515,In_58);
nand U156 (N_156,In_14,In_398);
and U157 (N_157,In_76,In_708);
nor U158 (N_158,In_266,In_645);
nand U159 (N_159,In_457,In_102);
or U160 (N_160,In_587,In_230);
and U161 (N_161,In_724,In_273);
nand U162 (N_162,In_400,In_29);
or U163 (N_163,In_79,In_605);
nor U164 (N_164,In_123,In_164);
nor U165 (N_165,In_341,In_593);
or U166 (N_166,In_61,In_547);
nand U167 (N_167,In_625,In_90);
nor U168 (N_168,In_425,In_472);
nand U169 (N_169,In_468,In_747);
or U170 (N_170,In_212,In_48);
nor U171 (N_171,In_467,In_220);
nand U172 (N_172,In_448,In_580);
nor U173 (N_173,In_505,In_643);
xor U174 (N_174,In_196,In_551);
and U175 (N_175,In_348,In_261);
nor U176 (N_176,In_699,In_219);
xnor U177 (N_177,In_99,In_537);
or U178 (N_178,In_482,In_599);
or U179 (N_179,In_185,In_35);
or U180 (N_180,In_449,In_491);
nand U181 (N_181,In_478,In_369);
or U182 (N_182,In_184,In_459);
or U183 (N_183,In_697,In_98);
and U184 (N_184,In_339,In_668);
or U185 (N_185,In_411,In_72);
nor U186 (N_186,In_585,In_389);
and U187 (N_187,In_652,In_534);
or U188 (N_188,In_493,In_100);
or U189 (N_189,In_320,In_328);
nand U190 (N_190,In_659,In_626);
nand U191 (N_191,In_531,In_171);
nor U192 (N_192,In_583,In_576);
nor U193 (N_193,In_473,In_541);
nand U194 (N_194,In_744,In_89);
nor U195 (N_195,In_333,In_0);
and U196 (N_196,In_297,In_136);
nand U197 (N_197,In_377,In_45);
nand U198 (N_198,In_160,In_257);
nand U199 (N_199,In_463,In_629);
or U200 (N_200,In_686,In_104);
or U201 (N_201,In_666,In_367);
nor U202 (N_202,In_470,In_262);
or U203 (N_203,In_719,In_424);
and U204 (N_204,In_162,In_329);
nand U205 (N_205,In_535,In_105);
nand U206 (N_206,In_91,In_139);
nor U207 (N_207,In_93,In_308);
nor U208 (N_208,In_390,In_590);
and U209 (N_209,In_460,In_152);
nor U210 (N_210,In_423,In_718);
and U211 (N_211,In_239,In_256);
and U212 (N_212,In_60,In_118);
nor U213 (N_213,In_295,In_661);
nor U214 (N_214,In_27,In_656);
and U215 (N_215,In_420,In_584);
nor U216 (N_216,In_574,In_86);
nand U217 (N_217,In_631,In_222);
or U218 (N_218,In_570,In_723);
and U219 (N_219,In_2,In_364);
and U220 (N_220,In_664,In_447);
nor U221 (N_221,In_518,In_19);
and U222 (N_222,In_729,In_131);
nor U223 (N_223,In_606,In_6);
and U224 (N_224,In_692,In_156);
nor U225 (N_225,In_260,In_651);
nand U226 (N_226,In_241,In_413);
and U227 (N_227,In_654,In_454);
nor U228 (N_228,In_440,In_275);
and U229 (N_229,In_739,In_1);
nor U230 (N_230,In_412,In_82);
nand U231 (N_231,In_594,In_669);
nor U232 (N_232,In_158,In_55);
nand U233 (N_233,In_525,In_748);
or U234 (N_234,In_494,In_233);
nand U235 (N_235,In_730,In_619);
nor U236 (N_236,In_107,In_357);
nand U237 (N_237,In_254,In_546);
nand U238 (N_238,In_416,In_588);
nor U239 (N_239,In_727,In_165);
or U240 (N_240,In_245,In_513);
nor U241 (N_241,In_343,In_287);
nor U242 (N_242,In_445,In_543);
nand U243 (N_243,In_237,In_5);
and U244 (N_244,In_32,In_112);
nor U245 (N_245,In_36,In_178);
and U246 (N_246,In_149,In_374);
nand U247 (N_247,In_250,In_129);
or U248 (N_248,In_242,In_701);
nand U249 (N_249,In_85,In_520);
or U250 (N_250,In_568,In_575);
and U251 (N_251,In_471,In_224);
and U252 (N_252,In_392,In_117);
and U253 (N_253,In_648,In_589);
or U254 (N_254,In_120,In_340);
and U255 (N_255,In_110,In_693);
and U256 (N_256,In_132,In_314);
and U257 (N_257,In_446,In_549);
or U258 (N_258,In_356,In_662);
and U259 (N_259,In_142,In_8);
or U260 (N_260,In_479,In_500);
nand U261 (N_261,In_73,In_509);
and U262 (N_262,In_53,In_269);
or U263 (N_263,In_458,In_336);
and U264 (N_264,In_92,In_548);
nand U265 (N_265,In_720,In_69);
and U266 (N_266,In_539,In_271);
and U267 (N_267,In_216,In_65);
nor U268 (N_268,In_624,In_71);
nor U269 (N_269,In_507,In_3);
xnor U270 (N_270,In_530,In_596);
nor U271 (N_271,In_461,In_94);
nor U272 (N_272,In_304,In_161);
nor U273 (N_273,In_114,In_512);
or U274 (N_274,In_16,In_368);
or U275 (N_275,In_415,In_452);
or U276 (N_276,In_728,In_462);
nand U277 (N_277,In_396,In_87);
nor U278 (N_278,In_726,In_203);
or U279 (N_279,In_128,In_612);
or U280 (N_280,In_567,In_410);
and U281 (N_281,In_342,In_506);
and U282 (N_282,In_644,In_556);
nor U283 (N_283,In_191,In_310);
and U284 (N_284,In_11,In_289);
nor U285 (N_285,In_281,In_265);
nand U286 (N_286,In_44,In_167);
nand U287 (N_287,In_354,In_109);
or U288 (N_288,In_595,In_502);
nand U289 (N_289,In_740,In_103);
or U290 (N_290,In_168,In_282);
and U291 (N_291,In_62,In_181);
or U292 (N_292,In_311,In_642);
nand U293 (N_293,In_251,In_397);
or U294 (N_294,In_665,In_742);
or U295 (N_295,In_345,In_653);
nand U296 (N_296,In_57,In_173);
nand U297 (N_297,In_157,In_735);
nor U298 (N_298,In_323,In_435);
nand U299 (N_299,In_660,In_359);
nand U300 (N_300,In_393,In_536);
or U301 (N_301,In_200,In_170);
or U302 (N_302,In_565,In_84);
nor U303 (N_303,In_638,In_34);
nand U304 (N_304,In_366,In_313);
and U305 (N_305,In_49,In_326);
and U306 (N_306,In_613,In_671);
or U307 (N_307,In_351,In_658);
or U308 (N_308,In_169,In_455);
nand U309 (N_309,In_620,In_155);
or U310 (N_310,In_678,In_77);
nand U311 (N_311,In_623,In_75);
nand U312 (N_312,In_337,In_276);
nor U313 (N_313,In_607,In_675);
or U314 (N_314,In_442,In_554);
xor U315 (N_315,In_116,In_263);
or U316 (N_316,In_307,In_202);
nor U317 (N_317,In_147,In_586);
nand U318 (N_318,In_182,In_694);
nand U319 (N_319,In_384,In_300);
or U320 (N_320,In_143,In_346);
nand U321 (N_321,In_698,In_51);
nand U322 (N_322,In_163,In_280);
or U323 (N_323,In_101,In_582);
nor U324 (N_324,In_316,In_81);
or U325 (N_325,In_370,In_714);
or U326 (N_326,In_721,In_126);
nand U327 (N_327,In_319,In_688);
and U328 (N_328,In_419,In_630);
nor U329 (N_329,In_497,In_215);
or U330 (N_330,In_30,In_283);
and U331 (N_331,In_140,In_17);
nor U332 (N_332,In_700,In_560);
nand U333 (N_333,In_221,In_488);
xnor U334 (N_334,In_453,In_684);
nor U335 (N_335,In_690,In_573);
nand U336 (N_336,In_672,In_600);
nor U337 (N_337,In_240,In_443);
nand U338 (N_338,In_66,In_456);
or U339 (N_339,In_113,In_450);
and U340 (N_340,In_673,In_725);
or U341 (N_341,In_676,In_572);
or U342 (N_342,In_228,In_274);
nand U343 (N_343,In_278,In_709);
nand U344 (N_344,In_483,In_258);
nor U345 (N_345,In_22,In_538);
nor U346 (N_346,In_617,In_325);
xor U347 (N_347,In_46,In_13);
and U348 (N_348,In_39,In_47);
or U349 (N_349,In_691,In_409);
nor U350 (N_350,In_439,In_706);
nand U351 (N_351,In_504,In_80);
or U352 (N_352,In_597,In_305);
nor U353 (N_353,In_133,In_562);
or U354 (N_354,In_24,In_322);
and U355 (N_355,In_646,In_144);
nor U356 (N_356,In_408,In_696);
nor U357 (N_357,In_146,In_249);
nand U358 (N_358,In_663,In_736);
or U359 (N_359,In_270,In_733);
nor U360 (N_360,In_119,In_731);
or U361 (N_361,In_738,In_481);
and U362 (N_362,In_331,In_372);
nand U363 (N_363,In_469,In_70);
nand U364 (N_364,In_633,In_50);
and U365 (N_365,In_236,In_253);
or U366 (N_366,In_213,In_639);
nand U367 (N_367,In_290,In_717);
and U368 (N_368,In_508,In_33);
and U369 (N_369,In_474,In_485);
nor U370 (N_370,In_25,In_235);
nor U371 (N_371,In_406,In_647);
nor U372 (N_372,In_555,In_464);
nand U373 (N_373,In_145,In_382);
and U374 (N_374,In_127,In_347);
nand U375 (N_375,In_55,In_648);
or U376 (N_376,In_52,In_162);
and U377 (N_377,In_647,In_416);
or U378 (N_378,In_500,In_564);
and U379 (N_379,In_56,In_734);
nand U380 (N_380,In_419,In_192);
or U381 (N_381,In_280,In_203);
nand U382 (N_382,In_188,In_269);
nand U383 (N_383,In_326,In_409);
and U384 (N_384,In_312,In_202);
nand U385 (N_385,In_636,In_433);
nand U386 (N_386,In_161,In_412);
nand U387 (N_387,In_494,In_535);
nand U388 (N_388,In_193,In_692);
nand U389 (N_389,In_395,In_144);
and U390 (N_390,In_138,In_24);
nand U391 (N_391,In_320,In_171);
nor U392 (N_392,In_113,In_493);
nand U393 (N_393,In_356,In_253);
nand U394 (N_394,In_280,In_725);
nand U395 (N_395,In_230,In_130);
nor U396 (N_396,In_464,In_204);
nand U397 (N_397,In_556,In_45);
nor U398 (N_398,In_373,In_526);
nor U399 (N_399,In_24,In_274);
nor U400 (N_400,In_621,In_677);
nand U401 (N_401,In_712,In_320);
nor U402 (N_402,In_504,In_513);
nand U403 (N_403,In_693,In_467);
and U404 (N_404,In_10,In_655);
nor U405 (N_405,In_279,In_243);
and U406 (N_406,In_685,In_605);
nor U407 (N_407,In_518,In_20);
nor U408 (N_408,In_594,In_584);
or U409 (N_409,In_286,In_94);
or U410 (N_410,In_137,In_655);
nand U411 (N_411,In_6,In_122);
and U412 (N_412,In_504,In_213);
and U413 (N_413,In_596,In_250);
and U414 (N_414,In_686,In_705);
nand U415 (N_415,In_280,In_87);
nand U416 (N_416,In_568,In_105);
nor U417 (N_417,In_128,In_190);
nand U418 (N_418,In_333,In_88);
nor U419 (N_419,In_508,In_264);
or U420 (N_420,In_92,In_88);
or U421 (N_421,In_254,In_227);
nand U422 (N_422,In_546,In_313);
nor U423 (N_423,In_82,In_339);
or U424 (N_424,In_380,In_583);
nor U425 (N_425,In_545,In_611);
nor U426 (N_426,In_481,In_413);
nor U427 (N_427,In_571,In_627);
or U428 (N_428,In_506,In_715);
nor U429 (N_429,In_316,In_647);
nand U430 (N_430,In_629,In_464);
nor U431 (N_431,In_653,In_150);
and U432 (N_432,In_348,In_190);
nand U433 (N_433,In_461,In_394);
nor U434 (N_434,In_273,In_565);
nand U435 (N_435,In_254,In_121);
and U436 (N_436,In_412,In_738);
nor U437 (N_437,In_143,In_633);
or U438 (N_438,In_478,In_578);
and U439 (N_439,In_42,In_633);
and U440 (N_440,In_129,In_176);
nor U441 (N_441,In_476,In_510);
and U442 (N_442,In_468,In_531);
xor U443 (N_443,In_330,In_589);
or U444 (N_444,In_44,In_524);
or U445 (N_445,In_656,In_130);
or U446 (N_446,In_510,In_190);
or U447 (N_447,In_231,In_527);
nor U448 (N_448,In_526,In_631);
and U449 (N_449,In_80,In_406);
and U450 (N_450,In_610,In_108);
nor U451 (N_451,In_671,In_112);
nor U452 (N_452,In_604,In_528);
or U453 (N_453,In_380,In_581);
nor U454 (N_454,In_356,In_494);
nand U455 (N_455,In_65,In_439);
and U456 (N_456,In_236,In_508);
nand U457 (N_457,In_528,In_38);
nor U458 (N_458,In_281,In_10);
nand U459 (N_459,In_327,In_740);
nor U460 (N_460,In_243,In_5);
and U461 (N_461,In_606,In_439);
or U462 (N_462,In_351,In_742);
or U463 (N_463,In_206,In_126);
nand U464 (N_464,In_321,In_704);
nor U465 (N_465,In_503,In_530);
nor U466 (N_466,In_749,In_455);
nand U467 (N_467,In_161,In_616);
and U468 (N_468,In_295,In_387);
or U469 (N_469,In_303,In_696);
or U470 (N_470,In_284,In_556);
or U471 (N_471,In_512,In_437);
and U472 (N_472,In_478,In_493);
nor U473 (N_473,In_34,In_708);
and U474 (N_474,In_389,In_295);
or U475 (N_475,In_470,In_275);
nor U476 (N_476,In_417,In_357);
nor U477 (N_477,In_364,In_196);
or U478 (N_478,In_38,In_491);
and U479 (N_479,In_566,In_399);
nand U480 (N_480,In_713,In_221);
or U481 (N_481,In_103,In_509);
xnor U482 (N_482,In_282,In_675);
nand U483 (N_483,In_416,In_727);
nand U484 (N_484,In_101,In_23);
or U485 (N_485,In_10,In_251);
nand U486 (N_486,In_706,In_101);
nor U487 (N_487,In_701,In_184);
or U488 (N_488,In_568,In_287);
nor U489 (N_489,In_26,In_557);
or U490 (N_490,In_626,In_662);
or U491 (N_491,In_599,In_180);
and U492 (N_492,In_597,In_654);
or U493 (N_493,In_538,In_64);
nor U494 (N_494,In_706,In_65);
nor U495 (N_495,In_110,In_699);
nor U496 (N_496,In_737,In_744);
or U497 (N_497,In_478,In_393);
nor U498 (N_498,In_265,In_451);
and U499 (N_499,In_690,In_89);
or U500 (N_500,N_327,N_229);
or U501 (N_501,N_230,N_39);
and U502 (N_502,N_66,N_266);
nand U503 (N_503,N_270,N_453);
and U504 (N_504,N_171,N_153);
and U505 (N_505,N_143,N_430);
and U506 (N_506,N_427,N_370);
nor U507 (N_507,N_286,N_397);
or U508 (N_508,N_373,N_490);
nand U509 (N_509,N_142,N_364);
or U510 (N_510,N_409,N_496);
and U511 (N_511,N_354,N_303);
nand U512 (N_512,N_60,N_29);
or U513 (N_513,N_477,N_269);
nand U514 (N_514,N_402,N_157);
nand U515 (N_515,N_369,N_235);
nor U516 (N_516,N_140,N_62);
or U517 (N_517,N_37,N_411);
or U518 (N_518,N_146,N_495);
or U519 (N_519,N_461,N_422);
nand U520 (N_520,N_420,N_443);
nand U521 (N_521,N_459,N_35);
and U522 (N_522,N_456,N_86);
nor U523 (N_523,N_399,N_185);
nand U524 (N_524,N_0,N_281);
or U525 (N_525,N_425,N_323);
nor U526 (N_526,N_435,N_170);
or U527 (N_527,N_466,N_22);
and U528 (N_528,N_126,N_240);
nand U529 (N_529,N_321,N_268);
and U530 (N_530,N_325,N_221);
and U531 (N_531,N_247,N_335);
nor U532 (N_532,N_84,N_380);
and U533 (N_533,N_244,N_474);
or U534 (N_534,N_377,N_89);
nor U535 (N_535,N_21,N_43);
or U536 (N_536,N_297,N_294);
nand U537 (N_537,N_121,N_254);
and U538 (N_538,N_467,N_304);
and U539 (N_539,N_180,N_174);
nor U540 (N_540,N_317,N_245);
nand U541 (N_541,N_205,N_154);
nor U542 (N_542,N_457,N_438);
and U543 (N_543,N_276,N_289);
or U544 (N_544,N_250,N_55);
or U545 (N_545,N_478,N_15);
and U546 (N_546,N_24,N_190);
nand U547 (N_547,N_346,N_204);
nor U548 (N_548,N_342,N_107);
nand U549 (N_549,N_387,N_395);
or U550 (N_550,N_407,N_177);
or U551 (N_551,N_94,N_40);
or U552 (N_552,N_120,N_163);
nand U553 (N_553,N_67,N_368);
or U554 (N_554,N_429,N_374);
or U555 (N_555,N_446,N_178);
nand U556 (N_556,N_376,N_287);
nand U557 (N_557,N_152,N_57);
or U558 (N_558,N_439,N_217);
and U559 (N_559,N_108,N_95);
or U560 (N_560,N_432,N_49);
xor U561 (N_561,N_225,N_5);
and U562 (N_562,N_487,N_129);
or U563 (N_563,N_423,N_234);
or U564 (N_564,N_20,N_122);
or U565 (N_565,N_292,N_127);
nor U566 (N_566,N_18,N_262);
nor U567 (N_567,N_285,N_194);
and U568 (N_568,N_104,N_184);
or U569 (N_569,N_372,N_238);
and U570 (N_570,N_295,N_222);
or U571 (N_571,N_92,N_110);
nor U572 (N_572,N_460,N_41);
nand U573 (N_573,N_385,N_74);
or U574 (N_574,N_421,N_351);
and U575 (N_575,N_463,N_48);
nand U576 (N_576,N_176,N_389);
nor U577 (N_577,N_26,N_246);
nor U578 (N_578,N_75,N_156);
nand U579 (N_579,N_81,N_88);
and U580 (N_580,N_381,N_279);
and U581 (N_581,N_444,N_261);
nor U582 (N_582,N_408,N_480);
nor U583 (N_583,N_32,N_436);
nor U584 (N_584,N_348,N_314);
or U585 (N_585,N_58,N_263);
nand U586 (N_586,N_79,N_476);
and U587 (N_587,N_251,N_207);
nand U588 (N_588,N_412,N_10);
nand U589 (N_589,N_72,N_273);
nor U590 (N_590,N_458,N_186);
nand U591 (N_591,N_382,N_272);
nor U592 (N_592,N_50,N_305);
nand U593 (N_593,N_344,N_454);
and U594 (N_594,N_260,N_36);
or U595 (N_595,N_187,N_396);
and U596 (N_596,N_492,N_352);
and U597 (N_597,N_394,N_138);
nor U598 (N_598,N_291,N_306);
or U599 (N_599,N_119,N_313);
nand U600 (N_600,N_455,N_134);
nand U601 (N_601,N_253,N_302);
or U602 (N_602,N_416,N_181);
nand U603 (N_603,N_341,N_312);
nand U604 (N_604,N_133,N_497);
nor U605 (N_605,N_350,N_355);
or U606 (N_606,N_202,N_52);
nand U607 (N_607,N_53,N_216);
and U608 (N_608,N_17,N_197);
and U609 (N_609,N_7,N_219);
or U610 (N_610,N_363,N_71);
or U611 (N_611,N_330,N_417);
or U612 (N_612,N_293,N_123);
and U613 (N_613,N_148,N_223);
and U614 (N_614,N_145,N_203);
or U615 (N_615,N_308,N_8);
nand U616 (N_616,N_437,N_329);
or U617 (N_617,N_360,N_301);
nand U618 (N_618,N_19,N_257);
or U619 (N_619,N_210,N_331);
and U620 (N_620,N_78,N_173);
nand U621 (N_621,N_220,N_82);
or U622 (N_622,N_465,N_379);
nor U623 (N_623,N_431,N_320);
nor U624 (N_624,N_200,N_103);
nor U625 (N_625,N_80,N_311);
or U626 (N_626,N_182,N_16);
nand U627 (N_627,N_68,N_340);
and U628 (N_628,N_124,N_452);
or U629 (N_629,N_169,N_14);
nand U630 (N_630,N_224,N_117);
and U631 (N_631,N_278,N_198);
or U632 (N_632,N_319,N_144);
nand U633 (N_633,N_404,N_97);
nor U634 (N_634,N_132,N_214);
nor U635 (N_635,N_256,N_299);
and U636 (N_636,N_267,N_99);
and U637 (N_637,N_63,N_131);
nor U638 (N_638,N_403,N_59);
or U639 (N_639,N_118,N_491);
and U640 (N_640,N_392,N_34);
and U641 (N_641,N_398,N_499);
nor U642 (N_642,N_201,N_415);
nor U643 (N_643,N_424,N_468);
and U644 (N_644,N_471,N_162);
nand U645 (N_645,N_195,N_275);
or U646 (N_646,N_324,N_393);
or U647 (N_647,N_358,N_390);
or U648 (N_648,N_4,N_356);
nand U649 (N_649,N_464,N_111);
and U650 (N_650,N_484,N_433);
nor U651 (N_651,N_115,N_472);
and U652 (N_652,N_332,N_384);
nor U653 (N_653,N_333,N_338);
or U654 (N_654,N_61,N_159);
and U655 (N_655,N_69,N_30);
or U656 (N_656,N_296,N_349);
nor U657 (N_657,N_42,N_189);
or U658 (N_658,N_45,N_191);
or U659 (N_659,N_9,N_307);
nand U660 (N_660,N_440,N_70);
nand U661 (N_661,N_298,N_136);
nor U662 (N_662,N_212,N_54);
nor U663 (N_663,N_151,N_12);
nand U664 (N_664,N_371,N_318);
nand U665 (N_665,N_228,N_188);
and U666 (N_666,N_388,N_445);
nand U667 (N_667,N_375,N_38);
or U668 (N_668,N_258,N_322);
nor U669 (N_669,N_249,N_326);
nor U670 (N_670,N_357,N_280);
and U671 (N_671,N_284,N_316);
or U672 (N_672,N_167,N_353);
or U673 (N_673,N_237,N_386);
nor U674 (N_674,N_46,N_259);
nor U675 (N_675,N_206,N_6);
nor U676 (N_676,N_486,N_13);
or U677 (N_677,N_473,N_31);
xnor U678 (N_678,N_227,N_116);
or U679 (N_679,N_215,N_91);
or U680 (N_680,N_196,N_83);
or U681 (N_681,N_252,N_483);
nor U682 (N_682,N_141,N_105);
or U683 (N_683,N_343,N_498);
nand U684 (N_684,N_1,N_98);
and U685 (N_685,N_413,N_147);
or U686 (N_686,N_150,N_77);
nor U687 (N_687,N_248,N_428);
nor U688 (N_688,N_277,N_47);
or U689 (N_689,N_494,N_164);
nand U690 (N_690,N_130,N_64);
nand U691 (N_691,N_336,N_106);
or U692 (N_692,N_96,N_208);
nor U693 (N_693,N_475,N_192);
or U694 (N_694,N_426,N_366);
nand U695 (N_695,N_193,N_168);
nand U696 (N_696,N_113,N_367);
or U697 (N_697,N_489,N_135);
and U698 (N_698,N_434,N_93);
and U699 (N_699,N_288,N_482);
nor U700 (N_700,N_87,N_469);
and U701 (N_701,N_418,N_264);
or U702 (N_702,N_405,N_337);
nand U703 (N_703,N_419,N_165);
nand U704 (N_704,N_211,N_25);
and U705 (N_705,N_400,N_243);
nor U706 (N_706,N_213,N_315);
xor U707 (N_707,N_265,N_442);
nor U708 (N_708,N_450,N_447);
or U709 (N_709,N_449,N_462);
or U710 (N_710,N_493,N_283);
and U711 (N_711,N_334,N_158);
and U712 (N_712,N_282,N_175);
and U713 (N_713,N_183,N_361);
or U714 (N_714,N_76,N_239);
or U715 (N_715,N_448,N_125);
nor U716 (N_716,N_137,N_410);
nor U717 (N_717,N_155,N_2);
and U718 (N_718,N_51,N_28);
or U719 (N_719,N_485,N_44);
or U720 (N_720,N_347,N_112);
or U721 (N_721,N_27,N_255);
and U722 (N_722,N_236,N_242);
or U723 (N_723,N_241,N_378);
nand U724 (N_724,N_179,N_23);
nand U725 (N_725,N_139,N_232);
and U726 (N_726,N_101,N_90);
and U727 (N_727,N_365,N_383);
or U728 (N_728,N_309,N_33);
or U729 (N_729,N_109,N_209);
nor U730 (N_730,N_73,N_3);
nor U731 (N_731,N_345,N_233);
or U732 (N_732,N_339,N_56);
or U733 (N_733,N_406,N_470);
or U734 (N_734,N_310,N_11);
or U735 (N_735,N_114,N_290);
or U736 (N_736,N_199,N_274);
nand U737 (N_737,N_102,N_149);
or U738 (N_738,N_100,N_271);
or U739 (N_739,N_441,N_161);
nand U740 (N_740,N_414,N_391);
and U741 (N_741,N_218,N_128);
or U742 (N_742,N_328,N_85);
nand U743 (N_743,N_488,N_231);
nor U744 (N_744,N_160,N_359);
nand U745 (N_745,N_65,N_166);
and U746 (N_746,N_479,N_362);
nor U747 (N_747,N_172,N_300);
or U748 (N_748,N_226,N_451);
and U749 (N_749,N_481,N_401);
or U750 (N_750,N_153,N_22);
and U751 (N_751,N_163,N_370);
nor U752 (N_752,N_200,N_165);
or U753 (N_753,N_251,N_434);
or U754 (N_754,N_50,N_355);
or U755 (N_755,N_432,N_50);
nand U756 (N_756,N_345,N_4);
nand U757 (N_757,N_396,N_120);
nor U758 (N_758,N_182,N_358);
or U759 (N_759,N_303,N_120);
and U760 (N_760,N_70,N_459);
and U761 (N_761,N_92,N_400);
nand U762 (N_762,N_258,N_278);
and U763 (N_763,N_203,N_103);
or U764 (N_764,N_397,N_98);
nor U765 (N_765,N_80,N_413);
nor U766 (N_766,N_318,N_141);
and U767 (N_767,N_346,N_444);
nand U768 (N_768,N_222,N_378);
or U769 (N_769,N_109,N_73);
or U770 (N_770,N_341,N_304);
or U771 (N_771,N_411,N_178);
nor U772 (N_772,N_247,N_147);
or U773 (N_773,N_280,N_470);
or U774 (N_774,N_299,N_20);
nor U775 (N_775,N_274,N_104);
and U776 (N_776,N_416,N_439);
or U777 (N_777,N_404,N_484);
or U778 (N_778,N_431,N_84);
or U779 (N_779,N_335,N_278);
nand U780 (N_780,N_408,N_361);
and U781 (N_781,N_232,N_492);
and U782 (N_782,N_409,N_298);
or U783 (N_783,N_179,N_231);
nand U784 (N_784,N_113,N_379);
nand U785 (N_785,N_373,N_130);
or U786 (N_786,N_191,N_131);
nor U787 (N_787,N_455,N_387);
nand U788 (N_788,N_479,N_153);
nor U789 (N_789,N_199,N_337);
or U790 (N_790,N_432,N_244);
nand U791 (N_791,N_421,N_293);
nor U792 (N_792,N_72,N_426);
or U793 (N_793,N_1,N_278);
and U794 (N_794,N_264,N_424);
or U795 (N_795,N_244,N_24);
and U796 (N_796,N_323,N_381);
nand U797 (N_797,N_158,N_97);
or U798 (N_798,N_158,N_254);
and U799 (N_799,N_261,N_81);
nor U800 (N_800,N_8,N_296);
nand U801 (N_801,N_464,N_352);
nor U802 (N_802,N_404,N_377);
nor U803 (N_803,N_268,N_496);
or U804 (N_804,N_400,N_65);
and U805 (N_805,N_389,N_52);
or U806 (N_806,N_103,N_481);
or U807 (N_807,N_276,N_224);
nor U808 (N_808,N_82,N_486);
or U809 (N_809,N_128,N_160);
nand U810 (N_810,N_468,N_189);
and U811 (N_811,N_27,N_236);
and U812 (N_812,N_185,N_31);
nand U813 (N_813,N_384,N_41);
nor U814 (N_814,N_6,N_143);
or U815 (N_815,N_434,N_155);
nand U816 (N_816,N_246,N_130);
or U817 (N_817,N_298,N_104);
and U818 (N_818,N_445,N_461);
nor U819 (N_819,N_221,N_172);
or U820 (N_820,N_406,N_6);
and U821 (N_821,N_405,N_375);
and U822 (N_822,N_213,N_334);
or U823 (N_823,N_69,N_26);
and U824 (N_824,N_239,N_229);
and U825 (N_825,N_263,N_352);
or U826 (N_826,N_436,N_255);
nor U827 (N_827,N_208,N_484);
nor U828 (N_828,N_236,N_50);
and U829 (N_829,N_259,N_320);
or U830 (N_830,N_416,N_163);
or U831 (N_831,N_306,N_78);
nand U832 (N_832,N_368,N_440);
nand U833 (N_833,N_420,N_74);
or U834 (N_834,N_248,N_397);
or U835 (N_835,N_462,N_303);
nand U836 (N_836,N_385,N_332);
or U837 (N_837,N_217,N_409);
nand U838 (N_838,N_453,N_4);
or U839 (N_839,N_73,N_97);
and U840 (N_840,N_101,N_449);
nand U841 (N_841,N_158,N_0);
nor U842 (N_842,N_465,N_134);
or U843 (N_843,N_482,N_437);
or U844 (N_844,N_224,N_260);
and U845 (N_845,N_14,N_124);
or U846 (N_846,N_130,N_439);
nor U847 (N_847,N_268,N_150);
or U848 (N_848,N_391,N_411);
and U849 (N_849,N_82,N_490);
nor U850 (N_850,N_123,N_162);
or U851 (N_851,N_429,N_351);
and U852 (N_852,N_482,N_389);
or U853 (N_853,N_449,N_294);
nor U854 (N_854,N_328,N_292);
nand U855 (N_855,N_486,N_214);
nand U856 (N_856,N_424,N_38);
and U857 (N_857,N_312,N_213);
nand U858 (N_858,N_362,N_437);
nor U859 (N_859,N_455,N_259);
nand U860 (N_860,N_173,N_495);
and U861 (N_861,N_296,N_255);
nand U862 (N_862,N_202,N_362);
nand U863 (N_863,N_162,N_364);
or U864 (N_864,N_51,N_308);
nand U865 (N_865,N_212,N_303);
and U866 (N_866,N_411,N_57);
nand U867 (N_867,N_9,N_476);
and U868 (N_868,N_205,N_348);
nand U869 (N_869,N_435,N_138);
or U870 (N_870,N_370,N_231);
nor U871 (N_871,N_29,N_453);
nand U872 (N_872,N_108,N_253);
nor U873 (N_873,N_71,N_237);
nor U874 (N_874,N_298,N_322);
and U875 (N_875,N_495,N_301);
and U876 (N_876,N_86,N_423);
xnor U877 (N_877,N_311,N_304);
or U878 (N_878,N_126,N_101);
or U879 (N_879,N_326,N_297);
or U880 (N_880,N_327,N_358);
or U881 (N_881,N_338,N_16);
or U882 (N_882,N_265,N_299);
nand U883 (N_883,N_265,N_322);
or U884 (N_884,N_90,N_257);
nor U885 (N_885,N_364,N_202);
and U886 (N_886,N_483,N_27);
and U887 (N_887,N_244,N_389);
nand U888 (N_888,N_444,N_11);
nand U889 (N_889,N_406,N_389);
and U890 (N_890,N_162,N_174);
and U891 (N_891,N_358,N_482);
and U892 (N_892,N_491,N_495);
and U893 (N_893,N_175,N_344);
and U894 (N_894,N_130,N_11);
or U895 (N_895,N_145,N_198);
nor U896 (N_896,N_456,N_357);
nand U897 (N_897,N_331,N_324);
nor U898 (N_898,N_147,N_26);
nor U899 (N_899,N_456,N_260);
nor U900 (N_900,N_385,N_18);
or U901 (N_901,N_450,N_103);
nor U902 (N_902,N_274,N_463);
or U903 (N_903,N_424,N_127);
nand U904 (N_904,N_360,N_43);
nand U905 (N_905,N_319,N_312);
or U906 (N_906,N_212,N_258);
nor U907 (N_907,N_330,N_409);
and U908 (N_908,N_450,N_115);
nor U909 (N_909,N_303,N_344);
and U910 (N_910,N_485,N_129);
or U911 (N_911,N_257,N_447);
nor U912 (N_912,N_291,N_485);
and U913 (N_913,N_183,N_389);
nand U914 (N_914,N_205,N_407);
and U915 (N_915,N_438,N_13);
nand U916 (N_916,N_43,N_215);
and U917 (N_917,N_74,N_406);
and U918 (N_918,N_144,N_494);
nand U919 (N_919,N_262,N_92);
nand U920 (N_920,N_407,N_352);
nor U921 (N_921,N_459,N_383);
nand U922 (N_922,N_49,N_120);
nand U923 (N_923,N_495,N_180);
or U924 (N_924,N_395,N_230);
nor U925 (N_925,N_287,N_372);
and U926 (N_926,N_425,N_104);
nor U927 (N_927,N_70,N_17);
nor U928 (N_928,N_180,N_406);
and U929 (N_929,N_34,N_78);
nand U930 (N_930,N_114,N_264);
or U931 (N_931,N_336,N_196);
nand U932 (N_932,N_433,N_212);
and U933 (N_933,N_233,N_262);
and U934 (N_934,N_354,N_182);
nor U935 (N_935,N_213,N_407);
or U936 (N_936,N_361,N_5);
or U937 (N_937,N_316,N_312);
nor U938 (N_938,N_378,N_209);
or U939 (N_939,N_26,N_158);
nand U940 (N_940,N_367,N_464);
or U941 (N_941,N_68,N_223);
nand U942 (N_942,N_347,N_404);
or U943 (N_943,N_277,N_82);
and U944 (N_944,N_82,N_426);
nand U945 (N_945,N_433,N_300);
nor U946 (N_946,N_490,N_457);
nor U947 (N_947,N_307,N_359);
nand U948 (N_948,N_53,N_337);
or U949 (N_949,N_6,N_491);
nor U950 (N_950,N_404,N_240);
nand U951 (N_951,N_3,N_2);
and U952 (N_952,N_407,N_485);
nor U953 (N_953,N_138,N_101);
nor U954 (N_954,N_417,N_358);
nor U955 (N_955,N_399,N_465);
nand U956 (N_956,N_379,N_425);
nand U957 (N_957,N_446,N_125);
or U958 (N_958,N_401,N_10);
nor U959 (N_959,N_468,N_282);
nand U960 (N_960,N_104,N_424);
nand U961 (N_961,N_111,N_14);
nor U962 (N_962,N_67,N_16);
nand U963 (N_963,N_224,N_493);
and U964 (N_964,N_98,N_342);
nor U965 (N_965,N_432,N_366);
nand U966 (N_966,N_281,N_171);
nand U967 (N_967,N_117,N_280);
nand U968 (N_968,N_231,N_407);
nand U969 (N_969,N_188,N_263);
and U970 (N_970,N_78,N_104);
nand U971 (N_971,N_129,N_175);
nor U972 (N_972,N_340,N_417);
nand U973 (N_973,N_217,N_476);
nor U974 (N_974,N_467,N_287);
nor U975 (N_975,N_322,N_55);
or U976 (N_976,N_3,N_483);
nor U977 (N_977,N_437,N_151);
and U978 (N_978,N_249,N_461);
xor U979 (N_979,N_450,N_290);
and U980 (N_980,N_93,N_491);
nor U981 (N_981,N_204,N_69);
or U982 (N_982,N_474,N_495);
or U983 (N_983,N_38,N_339);
nor U984 (N_984,N_116,N_135);
nand U985 (N_985,N_160,N_191);
and U986 (N_986,N_268,N_97);
or U987 (N_987,N_63,N_372);
nor U988 (N_988,N_495,N_37);
nand U989 (N_989,N_233,N_53);
nor U990 (N_990,N_206,N_82);
nand U991 (N_991,N_68,N_171);
nor U992 (N_992,N_375,N_433);
and U993 (N_993,N_203,N_137);
or U994 (N_994,N_266,N_357);
or U995 (N_995,N_441,N_76);
and U996 (N_996,N_364,N_290);
or U997 (N_997,N_115,N_36);
nor U998 (N_998,N_225,N_242);
and U999 (N_999,N_120,N_355);
nor U1000 (N_1000,N_943,N_510);
or U1001 (N_1001,N_888,N_779);
or U1002 (N_1002,N_683,N_516);
or U1003 (N_1003,N_873,N_660);
and U1004 (N_1004,N_801,N_596);
nor U1005 (N_1005,N_629,N_965);
or U1006 (N_1006,N_747,N_946);
and U1007 (N_1007,N_983,N_894);
or U1008 (N_1008,N_817,N_927);
and U1009 (N_1009,N_881,N_846);
and U1010 (N_1010,N_824,N_852);
and U1011 (N_1011,N_640,N_522);
and U1012 (N_1012,N_891,N_521);
or U1013 (N_1013,N_854,N_614);
or U1014 (N_1014,N_830,N_744);
nor U1015 (N_1015,N_851,N_875);
or U1016 (N_1016,N_843,N_858);
or U1017 (N_1017,N_804,N_589);
or U1018 (N_1018,N_922,N_869);
or U1019 (N_1019,N_880,N_790);
nor U1020 (N_1020,N_636,N_821);
or U1021 (N_1021,N_716,N_714);
and U1022 (N_1022,N_606,N_872);
and U1023 (N_1023,N_917,N_930);
nand U1024 (N_1024,N_592,N_643);
nand U1025 (N_1025,N_656,N_600);
and U1026 (N_1026,N_708,N_595);
and U1027 (N_1027,N_591,N_644);
nor U1028 (N_1028,N_655,N_558);
nor U1029 (N_1029,N_561,N_538);
or U1030 (N_1030,N_912,N_584);
nand U1031 (N_1031,N_529,N_884);
nor U1032 (N_1032,N_559,N_502);
nand U1033 (N_1033,N_932,N_715);
or U1034 (N_1034,N_967,N_972);
and U1035 (N_1035,N_757,N_899);
nand U1036 (N_1036,N_878,N_676);
or U1037 (N_1037,N_862,N_731);
or U1038 (N_1038,N_908,N_637);
nand U1039 (N_1039,N_749,N_760);
nand U1040 (N_1040,N_641,N_580);
xor U1041 (N_1041,N_977,N_577);
nor U1042 (N_1042,N_975,N_619);
and U1043 (N_1043,N_933,N_630);
nand U1044 (N_1044,N_945,N_910);
and U1045 (N_1045,N_585,N_816);
or U1046 (N_1046,N_634,N_954);
and U1047 (N_1047,N_610,N_935);
nand U1048 (N_1048,N_885,N_971);
nor U1049 (N_1049,N_753,N_926);
and U1050 (N_1050,N_506,N_669);
xor U1051 (N_1051,N_989,N_914);
and U1052 (N_1052,N_859,N_962);
nand U1053 (N_1053,N_787,N_900);
nand U1054 (N_1054,N_680,N_772);
and U1055 (N_1055,N_730,N_662);
nand U1056 (N_1056,N_666,N_921);
nand U1057 (N_1057,N_621,N_523);
nor U1058 (N_1058,N_686,N_920);
and U1059 (N_1059,N_889,N_618);
or U1060 (N_1060,N_844,N_831);
and U1061 (N_1061,N_796,N_537);
and U1062 (N_1062,N_707,N_729);
nand U1063 (N_1063,N_952,N_527);
and U1064 (N_1064,N_979,N_574);
nor U1065 (N_1065,N_761,N_609);
nor U1066 (N_1066,N_705,N_564);
or U1067 (N_1067,N_916,N_622);
and U1068 (N_1068,N_611,N_674);
nor U1069 (N_1069,N_832,N_951);
and U1070 (N_1070,N_845,N_692);
nor U1071 (N_1071,N_995,N_807);
or U1072 (N_1072,N_996,N_847);
nand U1073 (N_1073,N_955,N_877);
and U1074 (N_1074,N_649,N_587);
or U1075 (N_1075,N_557,N_755);
nor U1076 (N_1076,N_672,N_631);
or U1077 (N_1077,N_868,N_737);
and U1078 (N_1078,N_515,N_632);
or U1079 (N_1079,N_986,N_890);
nor U1080 (N_1080,N_808,N_982);
and U1081 (N_1081,N_987,N_825);
and U1082 (N_1082,N_937,N_726);
nor U1083 (N_1083,N_850,N_950);
and U1084 (N_1084,N_528,N_598);
nor U1085 (N_1085,N_700,N_756);
or U1086 (N_1086,N_735,N_997);
nand U1087 (N_1087,N_980,N_803);
or U1088 (N_1088,N_572,N_604);
and U1089 (N_1089,N_752,N_998);
or U1090 (N_1090,N_918,N_849);
nor U1091 (N_1091,N_758,N_782);
or U1092 (N_1092,N_810,N_767);
nand U1093 (N_1093,N_841,N_969);
nor U1094 (N_1094,N_990,N_588);
and U1095 (N_1095,N_569,N_958);
or U1096 (N_1096,N_913,N_578);
nor U1097 (N_1097,N_551,N_993);
or U1098 (N_1098,N_879,N_525);
and U1099 (N_1099,N_765,N_524);
or U1100 (N_1100,N_679,N_860);
nor U1101 (N_1101,N_773,N_745);
nand U1102 (N_1102,N_593,N_904);
nor U1103 (N_1103,N_953,N_536);
and U1104 (N_1104,N_925,N_976);
nand U1105 (N_1105,N_549,N_541);
or U1106 (N_1106,N_780,N_981);
and U1107 (N_1107,N_652,N_770);
and U1108 (N_1108,N_697,N_764);
nor U1109 (N_1109,N_734,N_689);
or U1110 (N_1110,N_728,N_939);
or U1111 (N_1111,N_819,N_766);
nand U1112 (N_1112,N_533,N_783);
nor U1113 (N_1113,N_777,N_661);
and U1114 (N_1114,N_809,N_778);
nand U1115 (N_1115,N_546,N_806);
or U1116 (N_1116,N_658,N_897);
nand U1117 (N_1117,N_836,N_973);
and U1118 (N_1118,N_603,N_815);
or U1119 (N_1119,N_663,N_504);
nand U1120 (N_1120,N_601,N_519);
xor U1121 (N_1121,N_638,N_776);
and U1122 (N_1122,N_813,N_542);
and U1123 (N_1123,N_853,N_500);
and U1124 (N_1124,N_795,N_896);
or U1125 (N_1125,N_985,N_691);
and U1126 (N_1126,N_511,N_812);
xor U1127 (N_1127,N_840,N_893);
nor U1128 (N_1128,N_863,N_909);
or U1129 (N_1129,N_948,N_722);
and U1130 (N_1130,N_670,N_583);
or U1131 (N_1131,N_828,N_507);
or U1132 (N_1132,N_837,N_581);
nand U1133 (N_1133,N_648,N_931);
and U1134 (N_1134,N_704,N_724);
nand U1135 (N_1135,N_709,N_740);
nand U1136 (N_1136,N_822,N_750);
nor U1137 (N_1137,N_923,N_883);
nand U1138 (N_1138,N_867,N_882);
nor U1139 (N_1139,N_599,N_690);
nor U1140 (N_1140,N_798,N_657);
xor U1141 (N_1141,N_838,N_608);
nor U1142 (N_1142,N_991,N_586);
nand U1143 (N_1143,N_905,N_762);
or U1144 (N_1144,N_876,N_548);
nand U1145 (N_1145,N_626,N_685);
nor U1146 (N_1146,N_653,N_797);
and U1147 (N_1147,N_827,N_960);
nand U1148 (N_1148,N_906,N_539);
nand U1149 (N_1149,N_668,N_526);
nor U1150 (N_1150,N_713,N_763);
nor U1151 (N_1151,N_695,N_794);
and U1152 (N_1152,N_911,N_781);
nand U1153 (N_1153,N_675,N_769);
nor U1154 (N_1154,N_940,N_957);
or U1155 (N_1155,N_984,N_791);
or U1156 (N_1156,N_964,N_746);
nand U1157 (N_1157,N_861,N_503);
and U1158 (N_1158,N_673,N_968);
nand U1159 (N_1159,N_919,N_842);
or U1160 (N_1160,N_712,N_605);
nand U1161 (N_1161,N_624,N_650);
nor U1162 (N_1162,N_811,N_855);
or U1163 (N_1163,N_992,N_505);
or U1164 (N_1164,N_959,N_509);
nor U1165 (N_1165,N_871,N_751);
or U1166 (N_1166,N_562,N_696);
nor U1167 (N_1167,N_924,N_620);
nand U1168 (N_1168,N_571,N_739);
nand U1169 (N_1169,N_699,N_775);
nand U1170 (N_1170,N_759,N_800);
nor U1171 (N_1171,N_701,N_508);
and U1172 (N_1172,N_568,N_517);
or U1173 (N_1173,N_901,N_540);
or U1174 (N_1174,N_710,N_789);
and U1175 (N_1175,N_566,N_999);
and U1176 (N_1176,N_874,N_949);
nor U1177 (N_1177,N_887,N_677);
nor U1178 (N_1178,N_625,N_938);
and U1179 (N_1179,N_902,N_839);
nand U1180 (N_1180,N_547,N_639);
nor U1181 (N_1181,N_907,N_742);
nand U1182 (N_1182,N_667,N_554);
and U1183 (N_1183,N_563,N_870);
and U1184 (N_1184,N_978,N_545);
or U1185 (N_1185,N_741,N_687);
nand U1186 (N_1186,N_963,N_627);
nor U1187 (N_1187,N_693,N_535);
or U1188 (N_1188,N_834,N_820);
nor U1189 (N_1189,N_857,N_956);
nor U1190 (N_1190,N_895,N_865);
nor U1191 (N_1191,N_848,N_736);
or U1192 (N_1192,N_799,N_768);
or U1193 (N_1193,N_645,N_602);
nor U1194 (N_1194,N_552,N_616);
nor U1195 (N_1195,N_560,N_771);
or U1196 (N_1196,N_928,N_617);
or U1197 (N_1197,N_886,N_646);
nand U1198 (N_1198,N_553,N_966);
and U1199 (N_1199,N_970,N_514);
and U1200 (N_1200,N_681,N_994);
and U1201 (N_1201,N_573,N_936);
nand U1202 (N_1202,N_774,N_555);
nor U1203 (N_1203,N_788,N_698);
or U1204 (N_1204,N_654,N_635);
nor U1205 (N_1205,N_941,N_597);
nand U1206 (N_1206,N_607,N_544);
nor U1207 (N_1207,N_719,N_594);
or U1208 (N_1208,N_612,N_633);
nor U1209 (N_1209,N_684,N_929);
and U1210 (N_1210,N_590,N_721);
and U1211 (N_1211,N_664,N_579);
nor U1212 (N_1212,N_628,N_892);
nand U1213 (N_1213,N_534,N_501);
nor U1214 (N_1214,N_814,N_550);
nor U1215 (N_1215,N_833,N_651);
nor U1216 (N_1216,N_518,N_988);
or U1217 (N_1217,N_512,N_513);
or U1218 (N_1218,N_532,N_738);
nand U1219 (N_1219,N_934,N_733);
nor U1220 (N_1220,N_711,N_665);
and U1221 (N_1221,N_520,N_530);
and U1222 (N_1222,N_898,N_835);
or U1223 (N_1223,N_702,N_718);
and U1224 (N_1224,N_623,N_732);
nand U1225 (N_1225,N_717,N_556);
nor U1226 (N_1226,N_942,N_543);
or U1227 (N_1227,N_678,N_531);
and U1228 (N_1228,N_576,N_915);
or U1229 (N_1229,N_725,N_743);
or U1230 (N_1230,N_582,N_947);
nand U1231 (N_1231,N_647,N_720);
nand U1232 (N_1232,N_961,N_671);
or U1233 (N_1233,N_829,N_688);
nor U1234 (N_1234,N_565,N_748);
nor U1235 (N_1235,N_805,N_754);
nand U1236 (N_1236,N_727,N_864);
and U1237 (N_1237,N_567,N_786);
and U1238 (N_1238,N_694,N_866);
or U1239 (N_1239,N_784,N_903);
or U1240 (N_1240,N_642,N_802);
nand U1241 (N_1241,N_793,N_792);
or U1242 (N_1242,N_856,N_826);
nor U1243 (N_1243,N_682,N_659);
and U1244 (N_1244,N_706,N_944);
nor U1245 (N_1245,N_785,N_703);
or U1246 (N_1246,N_613,N_575);
or U1247 (N_1247,N_615,N_570);
nand U1248 (N_1248,N_818,N_823);
and U1249 (N_1249,N_723,N_974);
or U1250 (N_1250,N_544,N_988);
nand U1251 (N_1251,N_712,N_778);
nor U1252 (N_1252,N_568,N_669);
nand U1253 (N_1253,N_675,N_875);
nor U1254 (N_1254,N_860,N_613);
and U1255 (N_1255,N_761,N_557);
and U1256 (N_1256,N_720,N_670);
or U1257 (N_1257,N_622,N_595);
and U1258 (N_1258,N_985,N_800);
nor U1259 (N_1259,N_730,N_842);
nand U1260 (N_1260,N_558,N_588);
nor U1261 (N_1261,N_531,N_658);
or U1262 (N_1262,N_968,N_564);
nand U1263 (N_1263,N_967,N_568);
or U1264 (N_1264,N_560,N_645);
and U1265 (N_1265,N_807,N_748);
or U1266 (N_1266,N_720,N_944);
nand U1267 (N_1267,N_972,N_551);
and U1268 (N_1268,N_896,N_739);
or U1269 (N_1269,N_634,N_817);
nor U1270 (N_1270,N_579,N_694);
or U1271 (N_1271,N_515,N_558);
and U1272 (N_1272,N_544,N_659);
nor U1273 (N_1273,N_835,N_615);
nand U1274 (N_1274,N_770,N_880);
nor U1275 (N_1275,N_646,N_533);
and U1276 (N_1276,N_757,N_995);
nor U1277 (N_1277,N_539,N_627);
or U1278 (N_1278,N_970,N_994);
nor U1279 (N_1279,N_507,N_966);
or U1280 (N_1280,N_557,N_589);
nor U1281 (N_1281,N_771,N_888);
nand U1282 (N_1282,N_651,N_766);
or U1283 (N_1283,N_859,N_583);
nor U1284 (N_1284,N_960,N_838);
and U1285 (N_1285,N_671,N_672);
nor U1286 (N_1286,N_896,N_572);
nand U1287 (N_1287,N_719,N_577);
nor U1288 (N_1288,N_865,N_798);
nor U1289 (N_1289,N_527,N_972);
or U1290 (N_1290,N_876,N_897);
nor U1291 (N_1291,N_794,N_961);
or U1292 (N_1292,N_510,N_792);
or U1293 (N_1293,N_627,N_521);
xor U1294 (N_1294,N_820,N_665);
and U1295 (N_1295,N_998,N_982);
nor U1296 (N_1296,N_633,N_623);
and U1297 (N_1297,N_651,N_952);
and U1298 (N_1298,N_959,N_730);
nor U1299 (N_1299,N_548,N_924);
nand U1300 (N_1300,N_573,N_525);
or U1301 (N_1301,N_743,N_556);
nor U1302 (N_1302,N_676,N_914);
or U1303 (N_1303,N_966,N_897);
nor U1304 (N_1304,N_978,N_747);
and U1305 (N_1305,N_865,N_691);
and U1306 (N_1306,N_689,N_744);
nor U1307 (N_1307,N_770,N_943);
and U1308 (N_1308,N_650,N_675);
or U1309 (N_1309,N_678,N_975);
nand U1310 (N_1310,N_789,N_773);
nand U1311 (N_1311,N_822,N_948);
and U1312 (N_1312,N_504,N_931);
nor U1313 (N_1313,N_684,N_574);
and U1314 (N_1314,N_842,N_508);
nand U1315 (N_1315,N_649,N_620);
or U1316 (N_1316,N_880,N_834);
nor U1317 (N_1317,N_619,N_843);
nand U1318 (N_1318,N_535,N_702);
or U1319 (N_1319,N_669,N_583);
and U1320 (N_1320,N_697,N_974);
and U1321 (N_1321,N_950,N_519);
or U1322 (N_1322,N_767,N_835);
and U1323 (N_1323,N_772,N_611);
and U1324 (N_1324,N_932,N_535);
nor U1325 (N_1325,N_864,N_972);
and U1326 (N_1326,N_674,N_512);
and U1327 (N_1327,N_528,N_722);
nand U1328 (N_1328,N_838,N_708);
and U1329 (N_1329,N_750,N_926);
or U1330 (N_1330,N_964,N_620);
or U1331 (N_1331,N_622,N_989);
nand U1332 (N_1332,N_724,N_556);
or U1333 (N_1333,N_965,N_707);
nor U1334 (N_1334,N_961,N_942);
nor U1335 (N_1335,N_627,N_504);
and U1336 (N_1336,N_732,N_596);
nor U1337 (N_1337,N_972,N_926);
or U1338 (N_1338,N_785,N_605);
and U1339 (N_1339,N_535,N_572);
or U1340 (N_1340,N_622,N_542);
nand U1341 (N_1341,N_619,N_806);
or U1342 (N_1342,N_915,N_798);
nor U1343 (N_1343,N_793,N_637);
nand U1344 (N_1344,N_615,N_611);
nand U1345 (N_1345,N_705,N_519);
xor U1346 (N_1346,N_854,N_949);
nor U1347 (N_1347,N_504,N_848);
or U1348 (N_1348,N_573,N_940);
or U1349 (N_1349,N_999,N_623);
and U1350 (N_1350,N_656,N_920);
or U1351 (N_1351,N_802,N_658);
nor U1352 (N_1352,N_526,N_995);
or U1353 (N_1353,N_882,N_535);
nor U1354 (N_1354,N_817,N_896);
nor U1355 (N_1355,N_531,N_881);
or U1356 (N_1356,N_853,N_588);
or U1357 (N_1357,N_717,N_510);
or U1358 (N_1358,N_579,N_726);
nor U1359 (N_1359,N_759,N_505);
nand U1360 (N_1360,N_816,N_608);
or U1361 (N_1361,N_746,N_627);
and U1362 (N_1362,N_735,N_688);
or U1363 (N_1363,N_791,N_814);
or U1364 (N_1364,N_678,N_804);
nor U1365 (N_1365,N_524,N_539);
or U1366 (N_1366,N_558,N_594);
or U1367 (N_1367,N_855,N_677);
nor U1368 (N_1368,N_871,N_561);
xnor U1369 (N_1369,N_569,N_862);
or U1370 (N_1370,N_582,N_631);
or U1371 (N_1371,N_590,N_814);
or U1372 (N_1372,N_998,N_809);
nand U1373 (N_1373,N_887,N_512);
nand U1374 (N_1374,N_932,N_729);
nor U1375 (N_1375,N_586,N_781);
nand U1376 (N_1376,N_711,N_737);
nand U1377 (N_1377,N_532,N_720);
and U1378 (N_1378,N_605,N_833);
nor U1379 (N_1379,N_838,N_550);
nand U1380 (N_1380,N_844,N_999);
nor U1381 (N_1381,N_629,N_960);
and U1382 (N_1382,N_739,N_609);
nor U1383 (N_1383,N_569,N_731);
nand U1384 (N_1384,N_826,N_962);
or U1385 (N_1385,N_875,N_650);
nor U1386 (N_1386,N_732,N_542);
nor U1387 (N_1387,N_500,N_598);
and U1388 (N_1388,N_585,N_561);
nor U1389 (N_1389,N_533,N_515);
or U1390 (N_1390,N_667,N_922);
and U1391 (N_1391,N_543,N_813);
nor U1392 (N_1392,N_654,N_842);
nor U1393 (N_1393,N_750,N_796);
or U1394 (N_1394,N_858,N_521);
and U1395 (N_1395,N_550,N_960);
and U1396 (N_1396,N_507,N_723);
or U1397 (N_1397,N_674,N_578);
nand U1398 (N_1398,N_907,N_765);
and U1399 (N_1399,N_761,N_771);
nand U1400 (N_1400,N_775,N_717);
nand U1401 (N_1401,N_984,N_573);
or U1402 (N_1402,N_666,N_927);
and U1403 (N_1403,N_848,N_631);
and U1404 (N_1404,N_999,N_700);
and U1405 (N_1405,N_988,N_808);
nor U1406 (N_1406,N_847,N_936);
nor U1407 (N_1407,N_614,N_954);
nand U1408 (N_1408,N_721,N_904);
or U1409 (N_1409,N_893,N_873);
or U1410 (N_1410,N_609,N_504);
and U1411 (N_1411,N_858,N_886);
nand U1412 (N_1412,N_709,N_956);
nand U1413 (N_1413,N_683,N_630);
or U1414 (N_1414,N_517,N_700);
nand U1415 (N_1415,N_669,N_730);
nor U1416 (N_1416,N_971,N_572);
and U1417 (N_1417,N_785,N_536);
and U1418 (N_1418,N_578,N_734);
nor U1419 (N_1419,N_571,N_909);
nor U1420 (N_1420,N_605,N_738);
nand U1421 (N_1421,N_726,N_729);
nor U1422 (N_1422,N_864,N_749);
or U1423 (N_1423,N_657,N_588);
nand U1424 (N_1424,N_657,N_731);
or U1425 (N_1425,N_856,N_785);
nand U1426 (N_1426,N_604,N_703);
or U1427 (N_1427,N_773,N_999);
or U1428 (N_1428,N_821,N_824);
or U1429 (N_1429,N_634,N_814);
nand U1430 (N_1430,N_976,N_783);
and U1431 (N_1431,N_929,N_751);
and U1432 (N_1432,N_686,N_511);
or U1433 (N_1433,N_995,N_901);
and U1434 (N_1434,N_762,N_547);
nor U1435 (N_1435,N_806,N_632);
nor U1436 (N_1436,N_827,N_981);
or U1437 (N_1437,N_629,N_635);
nand U1438 (N_1438,N_779,N_904);
nor U1439 (N_1439,N_695,N_883);
and U1440 (N_1440,N_683,N_905);
and U1441 (N_1441,N_583,N_961);
nor U1442 (N_1442,N_963,N_602);
nor U1443 (N_1443,N_540,N_685);
and U1444 (N_1444,N_782,N_925);
and U1445 (N_1445,N_665,N_516);
nor U1446 (N_1446,N_748,N_998);
or U1447 (N_1447,N_554,N_743);
nand U1448 (N_1448,N_712,N_748);
nand U1449 (N_1449,N_946,N_569);
and U1450 (N_1450,N_822,N_883);
or U1451 (N_1451,N_998,N_723);
or U1452 (N_1452,N_740,N_638);
nand U1453 (N_1453,N_556,N_648);
nand U1454 (N_1454,N_989,N_980);
nand U1455 (N_1455,N_559,N_625);
and U1456 (N_1456,N_639,N_599);
or U1457 (N_1457,N_955,N_842);
or U1458 (N_1458,N_625,N_741);
and U1459 (N_1459,N_750,N_549);
or U1460 (N_1460,N_642,N_975);
and U1461 (N_1461,N_575,N_570);
and U1462 (N_1462,N_607,N_896);
nor U1463 (N_1463,N_931,N_750);
xor U1464 (N_1464,N_733,N_660);
nor U1465 (N_1465,N_852,N_689);
and U1466 (N_1466,N_583,N_534);
nand U1467 (N_1467,N_896,N_618);
and U1468 (N_1468,N_597,N_822);
or U1469 (N_1469,N_996,N_693);
and U1470 (N_1470,N_757,N_766);
nand U1471 (N_1471,N_943,N_892);
nand U1472 (N_1472,N_685,N_965);
nor U1473 (N_1473,N_685,N_971);
nand U1474 (N_1474,N_578,N_979);
or U1475 (N_1475,N_802,N_951);
or U1476 (N_1476,N_582,N_896);
or U1477 (N_1477,N_999,N_683);
and U1478 (N_1478,N_526,N_838);
or U1479 (N_1479,N_700,N_542);
nand U1480 (N_1480,N_659,N_988);
and U1481 (N_1481,N_726,N_823);
or U1482 (N_1482,N_607,N_715);
nand U1483 (N_1483,N_517,N_637);
nor U1484 (N_1484,N_584,N_940);
or U1485 (N_1485,N_902,N_621);
nor U1486 (N_1486,N_718,N_922);
nor U1487 (N_1487,N_523,N_855);
nand U1488 (N_1488,N_662,N_808);
nor U1489 (N_1489,N_865,N_622);
nand U1490 (N_1490,N_789,N_696);
nand U1491 (N_1491,N_815,N_724);
nor U1492 (N_1492,N_822,N_970);
nor U1493 (N_1493,N_622,N_659);
nand U1494 (N_1494,N_641,N_723);
nor U1495 (N_1495,N_906,N_860);
and U1496 (N_1496,N_532,N_875);
and U1497 (N_1497,N_788,N_588);
nor U1498 (N_1498,N_566,N_908);
nor U1499 (N_1499,N_758,N_739);
nor U1500 (N_1500,N_1348,N_1176);
or U1501 (N_1501,N_1185,N_1338);
and U1502 (N_1502,N_1288,N_1189);
and U1503 (N_1503,N_1123,N_1262);
nor U1504 (N_1504,N_1427,N_1492);
or U1505 (N_1505,N_1308,N_1089);
and U1506 (N_1506,N_1265,N_1070);
nor U1507 (N_1507,N_1449,N_1048);
nor U1508 (N_1508,N_1418,N_1243);
or U1509 (N_1509,N_1360,N_1320);
and U1510 (N_1510,N_1356,N_1045);
nand U1511 (N_1511,N_1291,N_1112);
or U1512 (N_1512,N_1098,N_1416);
and U1513 (N_1513,N_1464,N_1069);
and U1514 (N_1514,N_1402,N_1461);
nand U1515 (N_1515,N_1335,N_1211);
or U1516 (N_1516,N_1429,N_1354);
or U1517 (N_1517,N_1293,N_1026);
nand U1518 (N_1518,N_1314,N_1479);
or U1519 (N_1519,N_1008,N_1081);
or U1520 (N_1520,N_1454,N_1346);
or U1521 (N_1521,N_1025,N_1286);
nor U1522 (N_1522,N_1412,N_1234);
nor U1523 (N_1523,N_1287,N_1106);
and U1524 (N_1524,N_1030,N_1166);
and U1525 (N_1525,N_1364,N_1319);
nor U1526 (N_1526,N_1143,N_1303);
nand U1527 (N_1527,N_1079,N_1295);
or U1528 (N_1528,N_1192,N_1311);
nand U1529 (N_1529,N_1160,N_1157);
xnor U1530 (N_1530,N_1007,N_1087);
and U1531 (N_1531,N_1236,N_1318);
nand U1532 (N_1532,N_1339,N_1156);
and U1533 (N_1533,N_1063,N_1086);
and U1534 (N_1534,N_1221,N_1271);
and U1535 (N_1535,N_1175,N_1014);
nand U1536 (N_1536,N_1426,N_1344);
nor U1537 (N_1537,N_1013,N_1050);
and U1538 (N_1538,N_1135,N_1423);
nand U1539 (N_1539,N_1336,N_1369);
or U1540 (N_1540,N_1327,N_1386);
or U1541 (N_1541,N_1302,N_1396);
or U1542 (N_1542,N_1233,N_1217);
or U1543 (N_1543,N_1273,N_1486);
nor U1544 (N_1544,N_1202,N_1000);
and U1545 (N_1545,N_1433,N_1326);
nand U1546 (N_1546,N_1357,N_1181);
or U1547 (N_1547,N_1116,N_1379);
nor U1548 (N_1548,N_1082,N_1068);
and U1549 (N_1549,N_1408,N_1158);
nand U1550 (N_1550,N_1391,N_1052);
nand U1551 (N_1551,N_1366,N_1307);
nand U1552 (N_1552,N_1496,N_1254);
or U1553 (N_1553,N_1137,N_1072);
nor U1554 (N_1554,N_1446,N_1195);
nor U1555 (N_1555,N_1235,N_1264);
nand U1556 (N_1556,N_1184,N_1256);
or U1557 (N_1557,N_1019,N_1436);
or U1558 (N_1558,N_1219,N_1041);
nand U1559 (N_1559,N_1392,N_1470);
nor U1560 (N_1560,N_1096,N_1373);
or U1561 (N_1561,N_1476,N_1110);
nand U1562 (N_1562,N_1440,N_1055);
or U1563 (N_1563,N_1100,N_1215);
or U1564 (N_1564,N_1332,N_1377);
nor U1565 (N_1565,N_1150,N_1197);
nor U1566 (N_1566,N_1238,N_1297);
nand U1567 (N_1567,N_1294,N_1385);
and U1568 (N_1568,N_1465,N_1011);
nand U1569 (N_1569,N_1053,N_1397);
and U1570 (N_1570,N_1359,N_1206);
and U1571 (N_1571,N_1457,N_1249);
and U1572 (N_1572,N_1462,N_1452);
nor U1573 (N_1573,N_1413,N_1194);
or U1574 (N_1574,N_1138,N_1438);
nor U1575 (N_1575,N_1115,N_1174);
nand U1576 (N_1576,N_1161,N_1490);
nor U1577 (N_1577,N_1054,N_1310);
and U1578 (N_1578,N_1225,N_1404);
nor U1579 (N_1579,N_1400,N_1152);
or U1580 (N_1580,N_1378,N_1274);
nor U1581 (N_1581,N_1409,N_1071);
nor U1582 (N_1582,N_1283,N_1450);
or U1583 (N_1583,N_1093,N_1384);
or U1584 (N_1584,N_1399,N_1488);
or U1585 (N_1585,N_1127,N_1204);
or U1586 (N_1586,N_1066,N_1201);
or U1587 (N_1587,N_1276,N_1421);
nor U1588 (N_1588,N_1095,N_1227);
or U1589 (N_1589,N_1343,N_1441);
or U1590 (N_1590,N_1261,N_1005);
and U1591 (N_1591,N_1428,N_1101);
or U1592 (N_1592,N_1376,N_1442);
nor U1593 (N_1593,N_1059,N_1237);
nor U1594 (N_1594,N_1362,N_1431);
or U1595 (N_1595,N_1322,N_1222);
and U1596 (N_1596,N_1368,N_1499);
and U1597 (N_1597,N_1131,N_1419);
or U1598 (N_1598,N_1459,N_1275);
xnor U1599 (N_1599,N_1186,N_1078);
nor U1600 (N_1600,N_1043,N_1193);
or U1601 (N_1601,N_1444,N_1021);
nand U1602 (N_1602,N_1352,N_1482);
and U1603 (N_1603,N_1417,N_1477);
and U1604 (N_1604,N_1472,N_1231);
nor U1605 (N_1605,N_1341,N_1272);
nor U1606 (N_1606,N_1448,N_1263);
nand U1607 (N_1607,N_1375,N_1382);
nor U1608 (N_1608,N_1002,N_1179);
nand U1609 (N_1609,N_1109,N_1269);
and U1610 (N_1610,N_1229,N_1244);
or U1611 (N_1611,N_1010,N_1387);
nor U1612 (N_1612,N_1102,N_1478);
nor U1613 (N_1613,N_1120,N_1337);
nor U1614 (N_1614,N_1240,N_1094);
or U1615 (N_1615,N_1042,N_1453);
nand U1616 (N_1616,N_1355,N_1140);
nand U1617 (N_1617,N_1033,N_1199);
nand U1618 (N_1618,N_1411,N_1155);
nor U1619 (N_1619,N_1434,N_1209);
and U1620 (N_1620,N_1430,N_1139);
or U1621 (N_1621,N_1024,N_1208);
nor U1622 (N_1622,N_1258,N_1187);
and U1623 (N_1623,N_1334,N_1463);
and U1624 (N_1624,N_1108,N_1437);
nor U1625 (N_1625,N_1245,N_1046);
nand U1626 (N_1626,N_1333,N_1006);
nor U1627 (N_1627,N_1018,N_1267);
and U1628 (N_1628,N_1493,N_1124);
nor U1629 (N_1629,N_1169,N_1372);
nor U1630 (N_1630,N_1312,N_1277);
and U1631 (N_1631,N_1065,N_1388);
nand U1632 (N_1632,N_1001,N_1383);
nor U1633 (N_1633,N_1188,N_1145);
nor U1634 (N_1634,N_1458,N_1498);
nor U1635 (N_1635,N_1415,N_1038);
and U1636 (N_1636,N_1313,N_1381);
nand U1637 (N_1637,N_1132,N_1456);
nand U1638 (N_1638,N_1035,N_1250);
or U1639 (N_1639,N_1178,N_1130);
or U1640 (N_1640,N_1363,N_1474);
nand U1641 (N_1641,N_1228,N_1298);
and U1642 (N_1642,N_1136,N_1049);
nand U1643 (N_1643,N_1279,N_1214);
xor U1644 (N_1644,N_1317,N_1309);
nor U1645 (N_1645,N_1304,N_1015);
or U1646 (N_1646,N_1029,N_1420);
nor U1647 (N_1647,N_1495,N_1321);
or U1648 (N_1648,N_1036,N_1075);
and U1649 (N_1649,N_1347,N_1284);
or U1650 (N_1650,N_1191,N_1114);
and U1651 (N_1651,N_1028,N_1003);
nand U1652 (N_1652,N_1260,N_1061);
or U1653 (N_1653,N_1058,N_1424);
and U1654 (N_1654,N_1126,N_1009);
and U1655 (N_1655,N_1056,N_1022);
or U1656 (N_1656,N_1253,N_1374);
and U1657 (N_1657,N_1128,N_1047);
nor U1658 (N_1658,N_1281,N_1301);
nor U1659 (N_1659,N_1497,N_1296);
or U1660 (N_1660,N_1349,N_1380);
nor U1661 (N_1661,N_1350,N_1084);
and U1662 (N_1662,N_1146,N_1012);
or U1663 (N_1663,N_1305,N_1398);
nor U1664 (N_1664,N_1190,N_1073);
or U1665 (N_1665,N_1090,N_1289);
nand U1666 (N_1666,N_1371,N_1257);
nor U1667 (N_1667,N_1023,N_1425);
and U1668 (N_1668,N_1224,N_1345);
or U1669 (N_1669,N_1422,N_1351);
nor U1670 (N_1670,N_1151,N_1467);
or U1671 (N_1671,N_1092,N_1051);
nor U1672 (N_1672,N_1034,N_1203);
and U1673 (N_1673,N_1171,N_1113);
or U1674 (N_1674,N_1083,N_1057);
or U1675 (N_1675,N_1252,N_1141);
or U1676 (N_1676,N_1062,N_1445);
nor U1677 (N_1677,N_1270,N_1125);
nor U1678 (N_1678,N_1266,N_1370);
or U1679 (N_1679,N_1358,N_1020);
nor U1680 (N_1680,N_1148,N_1282);
or U1681 (N_1681,N_1091,N_1162);
and U1682 (N_1682,N_1122,N_1172);
or U1683 (N_1683,N_1394,N_1401);
nand U1684 (N_1684,N_1247,N_1133);
and U1685 (N_1685,N_1365,N_1154);
and U1686 (N_1686,N_1099,N_1395);
nand U1687 (N_1687,N_1468,N_1159);
or U1688 (N_1688,N_1105,N_1300);
nand U1689 (N_1689,N_1016,N_1487);
nor U1690 (N_1690,N_1315,N_1330);
or U1691 (N_1691,N_1103,N_1435);
nand U1692 (N_1692,N_1111,N_1325);
nor U1693 (N_1693,N_1183,N_1246);
or U1694 (N_1694,N_1447,N_1306);
or U1695 (N_1695,N_1403,N_1207);
nor U1696 (N_1696,N_1040,N_1278);
nor U1697 (N_1697,N_1085,N_1242);
nand U1698 (N_1698,N_1216,N_1205);
nor U1699 (N_1699,N_1248,N_1353);
and U1700 (N_1700,N_1167,N_1340);
nand U1701 (N_1701,N_1134,N_1230);
and U1702 (N_1702,N_1443,N_1491);
nand U1703 (N_1703,N_1119,N_1218);
nand U1704 (N_1704,N_1483,N_1406);
and U1705 (N_1705,N_1212,N_1439);
or U1706 (N_1706,N_1080,N_1292);
and U1707 (N_1707,N_1389,N_1129);
and U1708 (N_1708,N_1484,N_1121);
or U1709 (N_1709,N_1144,N_1432);
xor U1710 (N_1710,N_1039,N_1097);
nor U1711 (N_1711,N_1475,N_1323);
nand U1712 (N_1712,N_1361,N_1466);
and U1713 (N_1713,N_1268,N_1060);
nor U1714 (N_1714,N_1032,N_1280);
nand U1715 (N_1715,N_1481,N_1460);
or U1716 (N_1716,N_1494,N_1107);
and U1717 (N_1717,N_1471,N_1076);
or U1718 (N_1718,N_1210,N_1407);
or U1719 (N_1719,N_1414,N_1077);
and U1720 (N_1720,N_1393,N_1117);
and U1721 (N_1721,N_1285,N_1290);
or U1722 (N_1722,N_1299,N_1004);
nand U1723 (N_1723,N_1324,N_1196);
nor U1724 (N_1724,N_1064,N_1149);
and U1725 (N_1725,N_1480,N_1153);
or U1726 (N_1726,N_1037,N_1200);
or U1727 (N_1727,N_1232,N_1198);
nor U1728 (N_1728,N_1180,N_1251);
and U1729 (N_1729,N_1331,N_1031);
nor U1730 (N_1730,N_1226,N_1165);
nand U1731 (N_1731,N_1173,N_1451);
nand U1732 (N_1732,N_1182,N_1316);
nor U1733 (N_1733,N_1485,N_1405);
and U1734 (N_1734,N_1220,N_1469);
and U1735 (N_1735,N_1142,N_1410);
or U1736 (N_1736,N_1067,N_1342);
and U1737 (N_1737,N_1027,N_1164);
nand U1738 (N_1738,N_1489,N_1088);
nand U1739 (N_1739,N_1328,N_1241);
and U1740 (N_1740,N_1168,N_1163);
nand U1741 (N_1741,N_1259,N_1170);
nand U1742 (N_1742,N_1390,N_1177);
or U1743 (N_1743,N_1104,N_1367);
or U1744 (N_1744,N_1455,N_1239);
and U1745 (N_1745,N_1223,N_1118);
nand U1746 (N_1746,N_1329,N_1255);
nor U1747 (N_1747,N_1147,N_1473);
nor U1748 (N_1748,N_1017,N_1074);
or U1749 (N_1749,N_1213,N_1044);
nand U1750 (N_1750,N_1384,N_1161);
or U1751 (N_1751,N_1437,N_1197);
or U1752 (N_1752,N_1296,N_1238);
nor U1753 (N_1753,N_1490,N_1104);
and U1754 (N_1754,N_1440,N_1138);
nor U1755 (N_1755,N_1189,N_1383);
and U1756 (N_1756,N_1374,N_1434);
nor U1757 (N_1757,N_1181,N_1100);
nor U1758 (N_1758,N_1195,N_1112);
and U1759 (N_1759,N_1122,N_1029);
or U1760 (N_1760,N_1370,N_1366);
and U1761 (N_1761,N_1319,N_1217);
xnor U1762 (N_1762,N_1202,N_1391);
nor U1763 (N_1763,N_1146,N_1081);
and U1764 (N_1764,N_1202,N_1041);
or U1765 (N_1765,N_1012,N_1228);
or U1766 (N_1766,N_1229,N_1074);
nor U1767 (N_1767,N_1473,N_1389);
or U1768 (N_1768,N_1316,N_1377);
and U1769 (N_1769,N_1096,N_1061);
nor U1770 (N_1770,N_1426,N_1381);
nor U1771 (N_1771,N_1497,N_1155);
or U1772 (N_1772,N_1134,N_1163);
nor U1773 (N_1773,N_1195,N_1089);
nand U1774 (N_1774,N_1301,N_1380);
or U1775 (N_1775,N_1321,N_1042);
nand U1776 (N_1776,N_1424,N_1283);
and U1777 (N_1777,N_1037,N_1206);
or U1778 (N_1778,N_1494,N_1155);
or U1779 (N_1779,N_1206,N_1442);
or U1780 (N_1780,N_1410,N_1117);
or U1781 (N_1781,N_1123,N_1032);
nor U1782 (N_1782,N_1111,N_1231);
nor U1783 (N_1783,N_1181,N_1064);
nor U1784 (N_1784,N_1232,N_1432);
and U1785 (N_1785,N_1373,N_1424);
nand U1786 (N_1786,N_1040,N_1409);
or U1787 (N_1787,N_1355,N_1054);
nand U1788 (N_1788,N_1069,N_1253);
and U1789 (N_1789,N_1250,N_1255);
nand U1790 (N_1790,N_1159,N_1256);
xor U1791 (N_1791,N_1054,N_1244);
nand U1792 (N_1792,N_1432,N_1275);
nand U1793 (N_1793,N_1370,N_1088);
nand U1794 (N_1794,N_1209,N_1387);
nor U1795 (N_1795,N_1299,N_1063);
or U1796 (N_1796,N_1278,N_1158);
nor U1797 (N_1797,N_1493,N_1469);
or U1798 (N_1798,N_1283,N_1004);
or U1799 (N_1799,N_1016,N_1381);
and U1800 (N_1800,N_1157,N_1119);
nand U1801 (N_1801,N_1025,N_1347);
nand U1802 (N_1802,N_1047,N_1095);
or U1803 (N_1803,N_1086,N_1487);
and U1804 (N_1804,N_1035,N_1429);
or U1805 (N_1805,N_1035,N_1210);
or U1806 (N_1806,N_1242,N_1233);
and U1807 (N_1807,N_1138,N_1418);
nand U1808 (N_1808,N_1073,N_1379);
nand U1809 (N_1809,N_1429,N_1377);
or U1810 (N_1810,N_1384,N_1282);
nand U1811 (N_1811,N_1324,N_1243);
xor U1812 (N_1812,N_1370,N_1005);
nand U1813 (N_1813,N_1218,N_1391);
xor U1814 (N_1814,N_1072,N_1360);
nor U1815 (N_1815,N_1339,N_1011);
nand U1816 (N_1816,N_1396,N_1223);
nor U1817 (N_1817,N_1325,N_1261);
and U1818 (N_1818,N_1294,N_1416);
or U1819 (N_1819,N_1336,N_1261);
nor U1820 (N_1820,N_1214,N_1063);
and U1821 (N_1821,N_1104,N_1306);
nor U1822 (N_1822,N_1317,N_1438);
nand U1823 (N_1823,N_1365,N_1029);
nor U1824 (N_1824,N_1163,N_1034);
or U1825 (N_1825,N_1156,N_1082);
nor U1826 (N_1826,N_1394,N_1301);
nor U1827 (N_1827,N_1307,N_1310);
or U1828 (N_1828,N_1492,N_1454);
or U1829 (N_1829,N_1269,N_1183);
nor U1830 (N_1830,N_1012,N_1080);
nor U1831 (N_1831,N_1339,N_1258);
and U1832 (N_1832,N_1469,N_1104);
or U1833 (N_1833,N_1417,N_1086);
nand U1834 (N_1834,N_1485,N_1389);
nand U1835 (N_1835,N_1216,N_1224);
or U1836 (N_1836,N_1081,N_1489);
nand U1837 (N_1837,N_1045,N_1355);
or U1838 (N_1838,N_1038,N_1440);
and U1839 (N_1839,N_1463,N_1101);
nand U1840 (N_1840,N_1275,N_1479);
or U1841 (N_1841,N_1239,N_1083);
nor U1842 (N_1842,N_1210,N_1395);
nor U1843 (N_1843,N_1457,N_1118);
nand U1844 (N_1844,N_1461,N_1292);
nor U1845 (N_1845,N_1035,N_1041);
nor U1846 (N_1846,N_1011,N_1128);
or U1847 (N_1847,N_1071,N_1378);
nand U1848 (N_1848,N_1219,N_1404);
nand U1849 (N_1849,N_1135,N_1039);
or U1850 (N_1850,N_1302,N_1408);
or U1851 (N_1851,N_1465,N_1206);
or U1852 (N_1852,N_1443,N_1002);
and U1853 (N_1853,N_1031,N_1441);
nand U1854 (N_1854,N_1368,N_1488);
nor U1855 (N_1855,N_1415,N_1152);
nor U1856 (N_1856,N_1332,N_1404);
nand U1857 (N_1857,N_1369,N_1079);
or U1858 (N_1858,N_1222,N_1301);
nor U1859 (N_1859,N_1214,N_1481);
nor U1860 (N_1860,N_1167,N_1210);
nand U1861 (N_1861,N_1473,N_1292);
and U1862 (N_1862,N_1267,N_1397);
and U1863 (N_1863,N_1063,N_1405);
nand U1864 (N_1864,N_1183,N_1294);
and U1865 (N_1865,N_1088,N_1209);
nand U1866 (N_1866,N_1112,N_1340);
and U1867 (N_1867,N_1089,N_1033);
and U1868 (N_1868,N_1228,N_1326);
nand U1869 (N_1869,N_1139,N_1290);
nor U1870 (N_1870,N_1081,N_1253);
nor U1871 (N_1871,N_1451,N_1158);
and U1872 (N_1872,N_1206,N_1179);
nand U1873 (N_1873,N_1209,N_1159);
nor U1874 (N_1874,N_1301,N_1277);
and U1875 (N_1875,N_1257,N_1141);
or U1876 (N_1876,N_1496,N_1471);
nand U1877 (N_1877,N_1244,N_1023);
nand U1878 (N_1878,N_1388,N_1310);
and U1879 (N_1879,N_1180,N_1306);
nor U1880 (N_1880,N_1144,N_1196);
nor U1881 (N_1881,N_1479,N_1318);
nand U1882 (N_1882,N_1260,N_1009);
xnor U1883 (N_1883,N_1107,N_1303);
or U1884 (N_1884,N_1400,N_1097);
xnor U1885 (N_1885,N_1246,N_1064);
and U1886 (N_1886,N_1218,N_1491);
or U1887 (N_1887,N_1233,N_1276);
and U1888 (N_1888,N_1479,N_1102);
and U1889 (N_1889,N_1378,N_1404);
nand U1890 (N_1890,N_1408,N_1134);
nor U1891 (N_1891,N_1231,N_1299);
nor U1892 (N_1892,N_1050,N_1431);
and U1893 (N_1893,N_1233,N_1333);
or U1894 (N_1894,N_1114,N_1406);
or U1895 (N_1895,N_1136,N_1372);
and U1896 (N_1896,N_1272,N_1344);
nor U1897 (N_1897,N_1416,N_1342);
nor U1898 (N_1898,N_1253,N_1335);
or U1899 (N_1899,N_1380,N_1414);
nor U1900 (N_1900,N_1407,N_1306);
and U1901 (N_1901,N_1482,N_1305);
or U1902 (N_1902,N_1031,N_1094);
and U1903 (N_1903,N_1381,N_1178);
nand U1904 (N_1904,N_1358,N_1270);
and U1905 (N_1905,N_1402,N_1238);
and U1906 (N_1906,N_1454,N_1189);
nand U1907 (N_1907,N_1314,N_1060);
or U1908 (N_1908,N_1396,N_1393);
xnor U1909 (N_1909,N_1093,N_1223);
nand U1910 (N_1910,N_1034,N_1340);
xnor U1911 (N_1911,N_1158,N_1134);
xnor U1912 (N_1912,N_1009,N_1360);
nand U1913 (N_1913,N_1032,N_1333);
and U1914 (N_1914,N_1303,N_1059);
nand U1915 (N_1915,N_1321,N_1323);
nor U1916 (N_1916,N_1374,N_1333);
nor U1917 (N_1917,N_1294,N_1186);
nand U1918 (N_1918,N_1128,N_1116);
nor U1919 (N_1919,N_1268,N_1475);
xnor U1920 (N_1920,N_1247,N_1146);
or U1921 (N_1921,N_1192,N_1051);
and U1922 (N_1922,N_1212,N_1393);
nand U1923 (N_1923,N_1180,N_1445);
and U1924 (N_1924,N_1232,N_1194);
nand U1925 (N_1925,N_1183,N_1136);
or U1926 (N_1926,N_1378,N_1147);
nand U1927 (N_1927,N_1027,N_1403);
nor U1928 (N_1928,N_1153,N_1015);
and U1929 (N_1929,N_1015,N_1433);
nor U1930 (N_1930,N_1150,N_1207);
or U1931 (N_1931,N_1470,N_1424);
or U1932 (N_1932,N_1208,N_1416);
or U1933 (N_1933,N_1339,N_1199);
and U1934 (N_1934,N_1221,N_1009);
and U1935 (N_1935,N_1320,N_1109);
or U1936 (N_1936,N_1493,N_1294);
nor U1937 (N_1937,N_1476,N_1138);
or U1938 (N_1938,N_1488,N_1150);
or U1939 (N_1939,N_1366,N_1153);
and U1940 (N_1940,N_1405,N_1103);
nor U1941 (N_1941,N_1214,N_1497);
and U1942 (N_1942,N_1239,N_1037);
and U1943 (N_1943,N_1476,N_1310);
and U1944 (N_1944,N_1456,N_1499);
or U1945 (N_1945,N_1037,N_1173);
nor U1946 (N_1946,N_1387,N_1073);
or U1947 (N_1947,N_1332,N_1492);
nand U1948 (N_1948,N_1042,N_1490);
and U1949 (N_1949,N_1151,N_1431);
nor U1950 (N_1950,N_1153,N_1297);
or U1951 (N_1951,N_1096,N_1461);
nor U1952 (N_1952,N_1371,N_1148);
or U1953 (N_1953,N_1069,N_1055);
or U1954 (N_1954,N_1366,N_1303);
nor U1955 (N_1955,N_1065,N_1414);
or U1956 (N_1956,N_1018,N_1039);
or U1957 (N_1957,N_1290,N_1375);
or U1958 (N_1958,N_1129,N_1209);
nand U1959 (N_1959,N_1044,N_1394);
nor U1960 (N_1960,N_1471,N_1090);
nand U1961 (N_1961,N_1109,N_1283);
nor U1962 (N_1962,N_1182,N_1050);
nand U1963 (N_1963,N_1135,N_1454);
nor U1964 (N_1964,N_1238,N_1491);
and U1965 (N_1965,N_1416,N_1433);
nand U1966 (N_1966,N_1191,N_1419);
and U1967 (N_1967,N_1271,N_1494);
nor U1968 (N_1968,N_1084,N_1308);
or U1969 (N_1969,N_1299,N_1403);
nor U1970 (N_1970,N_1048,N_1080);
and U1971 (N_1971,N_1375,N_1260);
or U1972 (N_1972,N_1358,N_1401);
and U1973 (N_1973,N_1377,N_1403);
and U1974 (N_1974,N_1248,N_1192);
nor U1975 (N_1975,N_1403,N_1368);
nor U1976 (N_1976,N_1257,N_1248);
and U1977 (N_1977,N_1437,N_1192);
nand U1978 (N_1978,N_1025,N_1050);
nand U1979 (N_1979,N_1094,N_1184);
and U1980 (N_1980,N_1191,N_1495);
and U1981 (N_1981,N_1141,N_1100);
or U1982 (N_1982,N_1047,N_1262);
and U1983 (N_1983,N_1055,N_1000);
nand U1984 (N_1984,N_1105,N_1299);
nand U1985 (N_1985,N_1470,N_1098);
or U1986 (N_1986,N_1234,N_1321);
nand U1987 (N_1987,N_1230,N_1439);
or U1988 (N_1988,N_1285,N_1423);
or U1989 (N_1989,N_1189,N_1011);
nor U1990 (N_1990,N_1139,N_1193);
or U1991 (N_1991,N_1129,N_1099);
and U1992 (N_1992,N_1176,N_1031);
nor U1993 (N_1993,N_1247,N_1044);
or U1994 (N_1994,N_1142,N_1437);
and U1995 (N_1995,N_1139,N_1303);
or U1996 (N_1996,N_1124,N_1262);
and U1997 (N_1997,N_1060,N_1203);
nor U1998 (N_1998,N_1142,N_1043);
nand U1999 (N_1999,N_1022,N_1151);
and U2000 (N_2000,N_1825,N_1913);
nor U2001 (N_2001,N_1650,N_1709);
nand U2002 (N_2002,N_1658,N_1888);
or U2003 (N_2003,N_1837,N_1646);
nand U2004 (N_2004,N_1692,N_1931);
or U2005 (N_2005,N_1636,N_1889);
nand U2006 (N_2006,N_1832,N_1640);
nand U2007 (N_2007,N_1839,N_1723);
or U2008 (N_2008,N_1786,N_1679);
and U2009 (N_2009,N_1727,N_1951);
nand U2010 (N_2010,N_1719,N_1745);
nor U2011 (N_2011,N_1608,N_1859);
nor U2012 (N_2012,N_1663,N_1974);
and U2013 (N_2013,N_1739,N_1941);
or U2014 (N_2014,N_1821,N_1885);
and U2015 (N_2015,N_1753,N_1903);
nor U2016 (N_2016,N_1670,N_1830);
nand U2017 (N_2017,N_1639,N_1828);
nor U2018 (N_2018,N_1550,N_1642);
and U2019 (N_2019,N_1935,N_1824);
or U2020 (N_2020,N_1558,N_1629);
nand U2021 (N_2021,N_1996,N_1770);
nor U2022 (N_2022,N_1609,N_1734);
or U2023 (N_2023,N_1812,N_1509);
and U2024 (N_2024,N_1796,N_1652);
nand U2025 (N_2025,N_1699,N_1746);
nand U2026 (N_2026,N_1947,N_1882);
nor U2027 (N_2027,N_1876,N_1660);
nor U2028 (N_2028,N_1841,N_1514);
and U2029 (N_2029,N_1905,N_1827);
and U2030 (N_2030,N_1715,N_1501);
and U2031 (N_2031,N_1602,N_1879);
and U2032 (N_2032,N_1689,N_1867);
nor U2033 (N_2033,N_1568,N_1543);
nand U2034 (N_2034,N_1814,N_1732);
nor U2035 (N_2035,N_1611,N_1928);
nor U2036 (N_2036,N_1983,N_1891);
nor U2037 (N_2037,N_1648,N_1920);
nand U2038 (N_2038,N_1529,N_1620);
nand U2039 (N_2039,N_1549,N_1556);
nand U2040 (N_2040,N_1690,N_1680);
and U2041 (N_2041,N_1532,N_1701);
and U2042 (N_2042,N_1728,N_1762);
and U2043 (N_2043,N_1647,N_1655);
and U2044 (N_2044,N_1518,N_1772);
nand U2045 (N_2045,N_1681,N_1741);
and U2046 (N_2046,N_1822,N_1809);
or U2047 (N_2047,N_1700,N_1989);
or U2048 (N_2048,N_1523,N_1619);
and U2049 (N_2049,N_1998,N_1717);
nand U2050 (N_2050,N_1845,N_1502);
nand U2051 (N_2051,N_1542,N_1548);
or U2052 (N_2052,N_1969,N_1565);
nand U2053 (N_2053,N_1711,N_1731);
and U2054 (N_2054,N_1541,N_1554);
or U2055 (N_2055,N_1840,N_1693);
or U2056 (N_2056,N_1994,N_1942);
nor U2057 (N_2057,N_1966,N_1789);
nor U2058 (N_2058,N_1666,N_1536);
or U2059 (N_2059,N_1597,N_1850);
nor U2060 (N_2060,N_1952,N_1937);
or U2061 (N_2061,N_1616,N_1980);
nor U2062 (N_2062,N_1587,N_1531);
nand U2063 (N_2063,N_1826,N_1904);
and U2064 (N_2064,N_1643,N_1632);
and U2065 (N_2065,N_1665,N_1933);
or U2066 (N_2066,N_1671,N_1783);
or U2067 (N_2067,N_1683,N_1939);
nand U2068 (N_2068,N_1914,N_1831);
nor U2069 (N_2069,N_1898,N_1856);
or U2070 (N_2070,N_1583,N_1992);
nand U2071 (N_2071,N_1976,N_1984);
nor U2072 (N_2072,N_1964,N_1967);
and U2073 (N_2073,N_1718,N_1563);
and U2074 (N_2074,N_1712,N_1860);
nand U2075 (N_2075,N_1634,N_1869);
or U2076 (N_2076,N_1686,N_1641);
or U2077 (N_2077,N_1977,N_1887);
and U2078 (N_2078,N_1667,N_1582);
and U2079 (N_2079,N_1673,N_1930);
nor U2080 (N_2080,N_1798,N_1813);
nand U2081 (N_2081,N_1806,N_1697);
or U2082 (N_2082,N_1958,N_1743);
or U2083 (N_2083,N_1703,N_1768);
and U2084 (N_2084,N_1907,N_1704);
nor U2085 (N_2085,N_1979,N_1672);
or U2086 (N_2086,N_1927,N_1775);
or U2087 (N_2087,N_1978,N_1661);
and U2088 (N_2088,N_1545,N_1784);
or U2089 (N_2089,N_1591,N_1803);
and U2090 (N_2090,N_1787,N_1526);
and U2091 (N_2091,N_1932,N_1566);
nor U2092 (N_2092,N_1596,N_1589);
nor U2093 (N_2093,N_1940,N_1788);
and U2094 (N_2094,N_1972,N_1564);
nor U2095 (N_2095,N_1910,N_1833);
or U2096 (N_2096,N_1573,N_1706);
nand U2097 (N_2097,N_1559,N_1780);
and U2098 (N_2098,N_1630,N_1623);
nand U2099 (N_2099,N_1735,N_1504);
nand U2100 (N_2100,N_1748,N_1971);
and U2101 (N_2101,N_1644,N_1569);
or U2102 (N_2102,N_1881,N_1677);
nand U2103 (N_2103,N_1970,N_1778);
and U2104 (N_2104,N_1560,N_1777);
and U2105 (N_2105,N_1886,N_1987);
and U2106 (N_2106,N_1506,N_1656);
and U2107 (N_2107,N_1747,N_1848);
and U2108 (N_2108,N_1613,N_1875);
nand U2109 (N_2109,N_1749,N_1818);
or U2110 (N_2110,N_1600,N_1835);
and U2111 (N_2111,N_1870,N_1515);
and U2112 (N_2112,N_1968,N_1555);
and U2113 (N_2113,N_1657,N_1946);
nand U2114 (N_2114,N_1864,N_1815);
and U2115 (N_2115,N_1638,N_1936);
nand U2116 (N_2116,N_1764,N_1552);
and U2117 (N_2117,N_1763,N_1628);
nor U2118 (N_2118,N_1820,N_1577);
nand U2119 (N_2119,N_1584,N_1605);
nand U2120 (N_2120,N_1893,N_1988);
nand U2121 (N_2121,N_1802,N_1938);
nand U2122 (N_2122,N_1752,N_1981);
nand U2123 (N_2123,N_1954,N_1624);
nand U2124 (N_2124,N_1729,N_1525);
and U2125 (N_2125,N_1738,N_1924);
nor U2126 (N_2126,N_1571,N_1794);
nand U2127 (N_2127,N_1742,N_1829);
nand U2128 (N_2128,N_1847,N_1512);
and U2129 (N_2129,N_1858,N_1817);
and U2130 (N_2130,N_1800,N_1923);
or U2131 (N_2131,N_1694,N_1621);
and U2132 (N_2132,N_1503,N_1684);
and U2133 (N_2133,N_1575,N_1909);
nand U2134 (N_2134,N_1849,N_1855);
or U2135 (N_2135,N_1810,N_1906);
nor U2136 (N_2136,N_1900,N_1902);
nand U2137 (N_2137,N_1883,N_1949);
or U2138 (N_2138,N_1737,N_1908);
nor U2139 (N_2139,N_1615,N_1520);
or U2140 (N_2140,N_1676,N_1539);
nor U2141 (N_2141,N_1895,N_1961);
and U2142 (N_2142,N_1588,N_1510);
nand U2143 (N_2143,N_1999,N_1912);
nor U2144 (N_2144,N_1612,N_1767);
nand U2145 (N_2145,N_1948,N_1842);
nand U2146 (N_2146,N_1544,N_1843);
and U2147 (N_2147,N_1635,N_1865);
or U2148 (N_2148,N_1956,N_1547);
or U2149 (N_2149,N_1846,N_1607);
or U2150 (N_2150,N_1664,N_1576);
nor U2151 (N_2151,N_1540,N_1557);
nand U2152 (N_2152,N_1754,N_1595);
or U2153 (N_2153,N_1857,N_1807);
or U2154 (N_2154,N_1537,N_1505);
and U2155 (N_2155,N_1511,N_1945);
or U2156 (N_2156,N_1530,N_1795);
or U2157 (N_2157,N_1592,N_1553);
nor U2158 (N_2158,N_1926,N_1863);
xnor U2159 (N_2159,N_1844,N_1880);
nor U2160 (N_2160,N_1950,N_1603);
and U2161 (N_2161,N_1799,N_1579);
nand U2162 (N_2162,N_1790,N_1707);
or U2163 (N_2163,N_1668,N_1853);
and U2164 (N_2164,N_1797,N_1890);
or U2165 (N_2165,N_1685,N_1943);
nand U2166 (N_2166,N_1601,N_1751);
or U2167 (N_2167,N_1804,N_1760);
nor U2168 (N_2168,N_1819,N_1561);
or U2169 (N_2169,N_1873,N_1722);
nand U2170 (N_2170,N_1546,N_1758);
nand U2171 (N_2171,N_1617,N_1878);
nor U2172 (N_2172,N_1744,N_1522);
nand U2173 (N_2173,N_1538,N_1769);
nor U2174 (N_2174,N_1791,N_1622);
and U2175 (N_2175,N_1725,N_1733);
nor U2176 (N_2176,N_1586,N_1513);
nand U2177 (N_2177,N_1955,N_1776);
nor U2178 (N_2178,N_1517,N_1919);
nand U2179 (N_2179,N_1986,N_1585);
nor U2180 (N_2180,N_1765,N_1614);
or U2181 (N_2181,N_1963,N_1953);
or U2182 (N_2182,N_1695,N_1757);
nor U2183 (N_2183,N_1519,N_1633);
and U2184 (N_2184,N_1637,N_1578);
or U2185 (N_2185,N_1698,N_1781);
nand U2186 (N_2186,N_1674,N_1500);
nand U2187 (N_2187,N_1771,N_1570);
and U2188 (N_2188,N_1726,N_1721);
and U2189 (N_2189,N_1884,N_1929);
and U2190 (N_2190,N_1590,N_1714);
or U2191 (N_2191,N_1528,N_1997);
and U2192 (N_2192,N_1593,N_1610);
nor U2193 (N_2193,N_1572,N_1918);
or U2194 (N_2194,N_1625,N_1861);
or U2195 (N_2195,N_1805,N_1599);
nor U2196 (N_2196,N_1836,N_1598);
or U2197 (N_2197,N_1736,N_1892);
nand U2198 (N_2198,N_1604,N_1960);
nor U2199 (N_2199,N_1702,N_1862);
nor U2200 (N_2200,N_1651,N_1682);
nor U2201 (N_2201,N_1959,N_1713);
nand U2202 (N_2202,N_1527,N_1811);
nand U2203 (N_2203,N_1991,N_1533);
nand U2204 (N_2204,N_1962,N_1975);
and U2205 (N_2205,N_1785,N_1896);
nand U2206 (N_2206,N_1816,N_1911);
nand U2207 (N_2207,N_1627,N_1897);
and U2208 (N_2208,N_1934,N_1982);
nand U2209 (N_2209,N_1782,N_1838);
nor U2210 (N_2210,N_1730,N_1581);
nand U2211 (N_2211,N_1990,N_1877);
nand U2212 (N_2212,N_1894,N_1834);
and U2213 (N_2213,N_1773,N_1944);
or U2214 (N_2214,N_1965,N_1688);
or U2215 (N_2215,N_1779,N_1710);
and U2216 (N_2216,N_1606,N_1766);
and U2217 (N_2217,N_1874,N_1516);
or U2218 (N_2218,N_1669,N_1567);
nand U2219 (N_2219,N_1562,N_1759);
nor U2220 (N_2220,N_1678,N_1922);
nand U2221 (N_2221,N_1649,N_1662);
or U2222 (N_2222,N_1915,N_1675);
or U2223 (N_2223,N_1696,N_1808);
nor U2224 (N_2224,N_1521,N_1851);
and U2225 (N_2225,N_1507,N_1973);
nor U2226 (N_2226,N_1750,N_1985);
or U2227 (N_2227,N_1871,N_1724);
and U2228 (N_2228,N_1508,N_1631);
nand U2229 (N_2229,N_1854,N_1823);
nor U2230 (N_2230,N_1774,N_1755);
nor U2231 (N_2231,N_1653,N_1580);
nor U2232 (N_2232,N_1574,N_1921);
nand U2233 (N_2233,N_1995,N_1645);
or U2234 (N_2234,N_1792,N_1708);
nand U2235 (N_2235,N_1551,N_1740);
or U2236 (N_2236,N_1626,N_1687);
nor U2237 (N_2237,N_1901,N_1654);
nand U2238 (N_2238,N_1917,N_1793);
nor U2239 (N_2239,N_1761,N_1993);
and U2240 (N_2240,N_1756,N_1866);
nor U2241 (N_2241,N_1925,N_1594);
nand U2242 (N_2242,N_1852,N_1691);
nand U2243 (N_2243,N_1868,N_1618);
nand U2244 (N_2244,N_1720,N_1716);
or U2245 (N_2245,N_1916,N_1801);
nor U2246 (N_2246,N_1535,N_1534);
nor U2247 (N_2247,N_1659,N_1899);
nand U2248 (N_2248,N_1705,N_1524);
or U2249 (N_2249,N_1872,N_1957);
and U2250 (N_2250,N_1973,N_1540);
and U2251 (N_2251,N_1734,N_1562);
nand U2252 (N_2252,N_1644,N_1778);
nand U2253 (N_2253,N_1776,N_1889);
nor U2254 (N_2254,N_1847,N_1763);
nor U2255 (N_2255,N_1932,N_1849);
and U2256 (N_2256,N_1738,N_1765);
nand U2257 (N_2257,N_1672,N_1884);
nor U2258 (N_2258,N_1668,N_1671);
or U2259 (N_2259,N_1969,N_1789);
nand U2260 (N_2260,N_1602,N_1932);
and U2261 (N_2261,N_1981,N_1612);
and U2262 (N_2262,N_1721,N_1876);
or U2263 (N_2263,N_1599,N_1904);
nand U2264 (N_2264,N_1998,N_1849);
nand U2265 (N_2265,N_1747,N_1672);
nor U2266 (N_2266,N_1523,N_1947);
or U2267 (N_2267,N_1701,N_1750);
xor U2268 (N_2268,N_1600,N_1712);
and U2269 (N_2269,N_1900,N_1764);
nand U2270 (N_2270,N_1812,N_1558);
nand U2271 (N_2271,N_1792,N_1762);
nand U2272 (N_2272,N_1774,N_1882);
or U2273 (N_2273,N_1593,N_1830);
nor U2274 (N_2274,N_1757,N_1844);
nor U2275 (N_2275,N_1609,N_1967);
nand U2276 (N_2276,N_1995,N_1642);
nor U2277 (N_2277,N_1696,N_1637);
and U2278 (N_2278,N_1744,N_1984);
and U2279 (N_2279,N_1733,N_1547);
nand U2280 (N_2280,N_1823,N_1634);
or U2281 (N_2281,N_1584,N_1786);
nor U2282 (N_2282,N_1918,N_1711);
and U2283 (N_2283,N_1827,N_1635);
nand U2284 (N_2284,N_1580,N_1607);
or U2285 (N_2285,N_1824,N_1687);
or U2286 (N_2286,N_1843,N_1998);
and U2287 (N_2287,N_1519,N_1566);
nand U2288 (N_2288,N_1827,N_1927);
or U2289 (N_2289,N_1559,N_1917);
and U2290 (N_2290,N_1817,N_1618);
or U2291 (N_2291,N_1504,N_1594);
nor U2292 (N_2292,N_1896,N_1573);
nor U2293 (N_2293,N_1649,N_1544);
nor U2294 (N_2294,N_1955,N_1895);
and U2295 (N_2295,N_1977,N_1758);
or U2296 (N_2296,N_1977,N_1764);
nor U2297 (N_2297,N_1802,N_1952);
and U2298 (N_2298,N_1781,N_1686);
or U2299 (N_2299,N_1942,N_1816);
nand U2300 (N_2300,N_1941,N_1586);
or U2301 (N_2301,N_1648,N_1558);
and U2302 (N_2302,N_1547,N_1630);
or U2303 (N_2303,N_1823,N_1660);
nor U2304 (N_2304,N_1989,N_1786);
nand U2305 (N_2305,N_1848,N_1681);
and U2306 (N_2306,N_1729,N_1857);
and U2307 (N_2307,N_1613,N_1562);
and U2308 (N_2308,N_1816,N_1540);
or U2309 (N_2309,N_1530,N_1880);
nand U2310 (N_2310,N_1811,N_1871);
or U2311 (N_2311,N_1904,N_1749);
nor U2312 (N_2312,N_1854,N_1763);
or U2313 (N_2313,N_1871,N_1778);
nor U2314 (N_2314,N_1560,N_1513);
nand U2315 (N_2315,N_1709,N_1794);
or U2316 (N_2316,N_1812,N_1675);
and U2317 (N_2317,N_1511,N_1965);
and U2318 (N_2318,N_1704,N_1587);
nand U2319 (N_2319,N_1595,N_1581);
nor U2320 (N_2320,N_1770,N_1568);
nor U2321 (N_2321,N_1915,N_1521);
nand U2322 (N_2322,N_1572,N_1513);
or U2323 (N_2323,N_1902,N_1923);
and U2324 (N_2324,N_1629,N_1863);
nand U2325 (N_2325,N_1702,N_1691);
nand U2326 (N_2326,N_1844,N_1852);
nand U2327 (N_2327,N_1658,N_1986);
nor U2328 (N_2328,N_1920,N_1851);
nor U2329 (N_2329,N_1666,N_1700);
or U2330 (N_2330,N_1654,N_1520);
nor U2331 (N_2331,N_1643,N_1840);
or U2332 (N_2332,N_1678,N_1802);
nor U2333 (N_2333,N_1558,N_1538);
nand U2334 (N_2334,N_1628,N_1683);
or U2335 (N_2335,N_1912,N_1532);
nand U2336 (N_2336,N_1784,N_1594);
nand U2337 (N_2337,N_1670,N_1895);
and U2338 (N_2338,N_1705,N_1681);
nor U2339 (N_2339,N_1512,N_1715);
nor U2340 (N_2340,N_1997,N_1679);
nand U2341 (N_2341,N_1910,N_1804);
nand U2342 (N_2342,N_1911,N_1881);
nand U2343 (N_2343,N_1966,N_1660);
or U2344 (N_2344,N_1609,N_1705);
nand U2345 (N_2345,N_1541,N_1505);
nor U2346 (N_2346,N_1708,N_1642);
nand U2347 (N_2347,N_1806,N_1583);
and U2348 (N_2348,N_1885,N_1776);
nand U2349 (N_2349,N_1533,N_1806);
nand U2350 (N_2350,N_1603,N_1987);
or U2351 (N_2351,N_1898,N_1988);
and U2352 (N_2352,N_1760,N_1527);
nand U2353 (N_2353,N_1827,N_1986);
nor U2354 (N_2354,N_1740,N_1723);
and U2355 (N_2355,N_1862,N_1803);
or U2356 (N_2356,N_1727,N_1925);
or U2357 (N_2357,N_1913,N_1713);
nor U2358 (N_2358,N_1980,N_1631);
nor U2359 (N_2359,N_1554,N_1704);
and U2360 (N_2360,N_1766,N_1892);
or U2361 (N_2361,N_1525,N_1668);
or U2362 (N_2362,N_1548,N_1670);
nor U2363 (N_2363,N_1986,N_1591);
or U2364 (N_2364,N_1558,N_1909);
nand U2365 (N_2365,N_1855,N_1942);
nand U2366 (N_2366,N_1869,N_1516);
and U2367 (N_2367,N_1904,N_1945);
nor U2368 (N_2368,N_1671,N_1924);
or U2369 (N_2369,N_1926,N_1578);
and U2370 (N_2370,N_1891,N_1807);
or U2371 (N_2371,N_1918,N_1630);
and U2372 (N_2372,N_1768,N_1587);
and U2373 (N_2373,N_1968,N_1978);
or U2374 (N_2374,N_1931,N_1699);
or U2375 (N_2375,N_1599,N_1592);
or U2376 (N_2376,N_1845,N_1916);
and U2377 (N_2377,N_1532,N_1771);
and U2378 (N_2378,N_1728,N_1838);
or U2379 (N_2379,N_1860,N_1632);
or U2380 (N_2380,N_1908,N_1568);
and U2381 (N_2381,N_1715,N_1764);
nor U2382 (N_2382,N_1562,N_1629);
nand U2383 (N_2383,N_1935,N_1785);
or U2384 (N_2384,N_1990,N_1510);
or U2385 (N_2385,N_1648,N_1574);
or U2386 (N_2386,N_1660,N_1530);
or U2387 (N_2387,N_1554,N_1551);
and U2388 (N_2388,N_1902,N_1836);
or U2389 (N_2389,N_1691,N_1526);
nand U2390 (N_2390,N_1776,N_1796);
or U2391 (N_2391,N_1957,N_1868);
or U2392 (N_2392,N_1513,N_1650);
and U2393 (N_2393,N_1683,N_1688);
and U2394 (N_2394,N_1764,N_1869);
or U2395 (N_2395,N_1558,N_1617);
nor U2396 (N_2396,N_1938,N_1640);
nand U2397 (N_2397,N_1534,N_1638);
or U2398 (N_2398,N_1572,N_1567);
nand U2399 (N_2399,N_1925,N_1855);
and U2400 (N_2400,N_1633,N_1673);
or U2401 (N_2401,N_1909,N_1715);
and U2402 (N_2402,N_1759,N_1925);
or U2403 (N_2403,N_1970,N_1671);
or U2404 (N_2404,N_1932,N_1968);
nand U2405 (N_2405,N_1929,N_1579);
or U2406 (N_2406,N_1743,N_1563);
or U2407 (N_2407,N_1840,N_1612);
nor U2408 (N_2408,N_1632,N_1690);
nor U2409 (N_2409,N_1634,N_1974);
and U2410 (N_2410,N_1835,N_1966);
nand U2411 (N_2411,N_1586,N_1511);
and U2412 (N_2412,N_1912,N_1684);
or U2413 (N_2413,N_1702,N_1864);
and U2414 (N_2414,N_1869,N_1910);
and U2415 (N_2415,N_1724,N_1983);
or U2416 (N_2416,N_1943,N_1811);
xor U2417 (N_2417,N_1953,N_1780);
nand U2418 (N_2418,N_1633,N_1877);
nand U2419 (N_2419,N_1557,N_1812);
or U2420 (N_2420,N_1993,N_1808);
nand U2421 (N_2421,N_1634,N_1763);
nor U2422 (N_2422,N_1971,N_1962);
nor U2423 (N_2423,N_1914,N_1780);
nor U2424 (N_2424,N_1586,N_1722);
nand U2425 (N_2425,N_1901,N_1953);
nand U2426 (N_2426,N_1741,N_1573);
nor U2427 (N_2427,N_1513,N_1910);
nand U2428 (N_2428,N_1919,N_1680);
nand U2429 (N_2429,N_1958,N_1927);
and U2430 (N_2430,N_1993,N_1529);
nor U2431 (N_2431,N_1622,N_1829);
and U2432 (N_2432,N_1882,N_1606);
nand U2433 (N_2433,N_1892,N_1885);
and U2434 (N_2434,N_1562,N_1609);
nor U2435 (N_2435,N_1526,N_1946);
or U2436 (N_2436,N_1651,N_1612);
nor U2437 (N_2437,N_1965,N_1851);
and U2438 (N_2438,N_1802,N_1674);
nand U2439 (N_2439,N_1899,N_1962);
nand U2440 (N_2440,N_1741,N_1850);
and U2441 (N_2441,N_1656,N_1567);
or U2442 (N_2442,N_1999,N_1881);
nor U2443 (N_2443,N_1733,N_1842);
or U2444 (N_2444,N_1871,N_1705);
nor U2445 (N_2445,N_1714,N_1863);
xor U2446 (N_2446,N_1617,N_1606);
nand U2447 (N_2447,N_1929,N_1645);
nor U2448 (N_2448,N_1716,N_1783);
or U2449 (N_2449,N_1553,N_1607);
or U2450 (N_2450,N_1849,N_1623);
and U2451 (N_2451,N_1801,N_1643);
xnor U2452 (N_2452,N_1748,N_1569);
nand U2453 (N_2453,N_1967,N_1951);
nor U2454 (N_2454,N_1628,N_1633);
and U2455 (N_2455,N_1794,N_1966);
or U2456 (N_2456,N_1597,N_1717);
and U2457 (N_2457,N_1983,N_1611);
or U2458 (N_2458,N_1633,N_1935);
and U2459 (N_2459,N_1661,N_1519);
or U2460 (N_2460,N_1712,N_1899);
nand U2461 (N_2461,N_1866,N_1989);
nand U2462 (N_2462,N_1900,N_1924);
or U2463 (N_2463,N_1783,N_1986);
or U2464 (N_2464,N_1982,N_1571);
nand U2465 (N_2465,N_1831,N_1912);
nand U2466 (N_2466,N_1951,N_1684);
and U2467 (N_2467,N_1723,N_1840);
xor U2468 (N_2468,N_1813,N_1729);
xnor U2469 (N_2469,N_1890,N_1642);
and U2470 (N_2470,N_1963,N_1903);
nand U2471 (N_2471,N_1775,N_1872);
nand U2472 (N_2472,N_1883,N_1722);
or U2473 (N_2473,N_1512,N_1910);
nor U2474 (N_2474,N_1518,N_1980);
nand U2475 (N_2475,N_1637,N_1531);
or U2476 (N_2476,N_1646,N_1535);
nor U2477 (N_2477,N_1677,N_1782);
or U2478 (N_2478,N_1847,N_1507);
or U2479 (N_2479,N_1567,N_1944);
nor U2480 (N_2480,N_1799,N_1760);
nor U2481 (N_2481,N_1545,N_1815);
and U2482 (N_2482,N_1979,N_1703);
nand U2483 (N_2483,N_1919,N_1853);
nand U2484 (N_2484,N_1981,N_1599);
nor U2485 (N_2485,N_1721,N_1522);
and U2486 (N_2486,N_1551,N_1555);
nand U2487 (N_2487,N_1548,N_1843);
or U2488 (N_2488,N_1850,N_1779);
nand U2489 (N_2489,N_1760,N_1884);
nand U2490 (N_2490,N_1746,N_1840);
nor U2491 (N_2491,N_1720,N_1872);
or U2492 (N_2492,N_1506,N_1713);
nand U2493 (N_2493,N_1583,N_1808);
xnor U2494 (N_2494,N_1504,N_1701);
nand U2495 (N_2495,N_1999,N_1795);
nand U2496 (N_2496,N_1553,N_1753);
and U2497 (N_2497,N_1670,N_1842);
or U2498 (N_2498,N_1922,N_1773);
or U2499 (N_2499,N_1945,N_1846);
nand U2500 (N_2500,N_2179,N_2269);
and U2501 (N_2501,N_2390,N_2309);
nor U2502 (N_2502,N_2335,N_2461);
nand U2503 (N_2503,N_2305,N_2011);
or U2504 (N_2504,N_2300,N_2342);
nand U2505 (N_2505,N_2022,N_2105);
nor U2506 (N_2506,N_2338,N_2002);
nor U2507 (N_2507,N_2285,N_2456);
nor U2508 (N_2508,N_2268,N_2173);
and U2509 (N_2509,N_2228,N_2237);
or U2510 (N_2510,N_2183,N_2123);
and U2511 (N_2511,N_2312,N_2182);
nand U2512 (N_2512,N_2129,N_2274);
nor U2513 (N_2513,N_2201,N_2127);
nand U2514 (N_2514,N_2073,N_2012);
nor U2515 (N_2515,N_2157,N_2125);
and U2516 (N_2516,N_2346,N_2004);
and U2517 (N_2517,N_2333,N_2009);
and U2518 (N_2518,N_2055,N_2374);
nor U2519 (N_2519,N_2047,N_2408);
or U2520 (N_2520,N_2304,N_2024);
nor U2521 (N_2521,N_2033,N_2085);
nor U2522 (N_2522,N_2495,N_2441);
nand U2523 (N_2523,N_2243,N_2034);
and U2524 (N_2524,N_2056,N_2329);
and U2525 (N_2525,N_2153,N_2241);
and U2526 (N_2526,N_2496,N_2040);
or U2527 (N_2527,N_2164,N_2350);
and U2528 (N_2528,N_2299,N_2287);
nor U2529 (N_2529,N_2330,N_2370);
nor U2530 (N_2530,N_2439,N_2027);
nor U2531 (N_2531,N_2025,N_2006);
and U2532 (N_2532,N_2298,N_2000);
nor U2533 (N_2533,N_2210,N_2372);
nor U2534 (N_2534,N_2136,N_2071);
or U2535 (N_2535,N_2388,N_2355);
or U2536 (N_2536,N_2120,N_2239);
nand U2537 (N_2537,N_2231,N_2322);
nor U2538 (N_2538,N_2297,N_2483);
nor U2539 (N_2539,N_2475,N_2396);
xnor U2540 (N_2540,N_2045,N_2276);
xor U2541 (N_2541,N_2072,N_2489);
nand U2542 (N_2542,N_2499,N_2411);
or U2543 (N_2543,N_2178,N_2049);
and U2544 (N_2544,N_2263,N_2240);
nand U2545 (N_2545,N_2340,N_2395);
nand U2546 (N_2546,N_2194,N_2133);
and U2547 (N_2547,N_2115,N_2460);
and U2548 (N_2548,N_2198,N_2116);
nor U2549 (N_2549,N_2486,N_2223);
xnor U2550 (N_2550,N_2348,N_2387);
and U2551 (N_2551,N_2193,N_2169);
nor U2552 (N_2552,N_2061,N_2070);
nor U2553 (N_2553,N_2066,N_2467);
nand U2554 (N_2554,N_2255,N_2039);
and U2555 (N_2555,N_2165,N_2368);
or U2556 (N_2556,N_2093,N_2384);
nor U2557 (N_2557,N_2290,N_2319);
nor U2558 (N_2558,N_2067,N_2087);
and U2559 (N_2559,N_2209,N_2122);
and U2560 (N_2560,N_2422,N_2491);
nor U2561 (N_2561,N_2454,N_2477);
nor U2562 (N_2562,N_2075,N_2453);
and U2563 (N_2563,N_2236,N_2278);
or U2564 (N_2564,N_2135,N_2493);
or U2565 (N_2565,N_2341,N_2124);
nand U2566 (N_2566,N_2143,N_2036);
and U2567 (N_2567,N_2028,N_2168);
or U2568 (N_2568,N_2054,N_2212);
nor U2569 (N_2569,N_2280,N_2366);
nand U2570 (N_2570,N_2139,N_2147);
or U2571 (N_2571,N_2214,N_2320);
and U2572 (N_2572,N_2121,N_2302);
or U2573 (N_2573,N_2331,N_2277);
or U2574 (N_2574,N_2401,N_2177);
nand U2575 (N_2575,N_2259,N_2389);
and U2576 (N_2576,N_2421,N_2205);
nand U2577 (N_2577,N_2437,N_2138);
or U2578 (N_2578,N_2482,N_2215);
or U2579 (N_2579,N_2288,N_2472);
nand U2580 (N_2580,N_2469,N_2118);
nand U2581 (N_2581,N_2220,N_2050);
and U2582 (N_2582,N_2332,N_2434);
or U2583 (N_2583,N_2037,N_2038);
nor U2584 (N_2584,N_2371,N_2393);
and U2585 (N_2585,N_2398,N_2404);
nand U2586 (N_2586,N_2443,N_2052);
or U2587 (N_2587,N_2494,N_2289);
nor U2588 (N_2588,N_2058,N_2023);
and U2589 (N_2589,N_2099,N_2146);
or U2590 (N_2590,N_2046,N_2159);
nor U2591 (N_2591,N_2185,N_2447);
nor U2592 (N_2592,N_2271,N_2174);
or U2593 (N_2593,N_2232,N_2253);
nand U2594 (N_2594,N_2474,N_2292);
or U2595 (N_2595,N_2021,N_2065);
nor U2596 (N_2596,N_2427,N_2111);
nor U2597 (N_2597,N_2318,N_2378);
and U2598 (N_2598,N_2222,N_2266);
or U2599 (N_2599,N_2418,N_2150);
and U2600 (N_2600,N_2386,N_2369);
or U2601 (N_2601,N_2468,N_2286);
and U2602 (N_2602,N_2188,N_2078);
and U2603 (N_2603,N_2257,N_2128);
nor U2604 (N_2604,N_2323,N_2126);
and U2605 (N_2605,N_2248,N_2432);
nand U2606 (N_2606,N_2360,N_2195);
and U2607 (N_2607,N_2272,N_2016);
nand U2608 (N_2608,N_2132,N_2249);
nor U2609 (N_2609,N_2451,N_2315);
or U2610 (N_2610,N_2227,N_2156);
or U2611 (N_2611,N_2013,N_2385);
and U2612 (N_2612,N_2303,N_2353);
nand U2613 (N_2613,N_2470,N_2416);
and U2614 (N_2614,N_2196,N_2244);
nor U2615 (N_2615,N_2082,N_2362);
and U2616 (N_2616,N_2379,N_2308);
and U2617 (N_2617,N_2096,N_2083);
nor U2618 (N_2618,N_2351,N_2086);
or U2619 (N_2619,N_2254,N_2435);
nand U2620 (N_2620,N_2017,N_2191);
nor U2621 (N_2621,N_2192,N_2184);
or U2622 (N_2622,N_2283,N_2035);
and U2623 (N_2623,N_2317,N_2092);
nor U2624 (N_2624,N_2203,N_2463);
or U2625 (N_2625,N_2314,N_2079);
or U2626 (N_2626,N_2485,N_2026);
nand U2627 (N_2627,N_2490,N_2197);
or U2628 (N_2628,N_2258,N_2359);
or U2629 (N_2629,N_2161,N_2029);
nand U2630 (N_2630,N_2295,N_2336);
nand U2631 (N_2631,N_2020,N_2270);
nand U2632 (N_2632,N_2445,N_2252);
nor U2633 (N_2633,N_2113,N_2114);
or U2634 (N_2634,N_2217,N_2063);
or U2635 (N_2635,N_2446,N_2431);
nor U2636 (N_2636,N_2417,N_2264);
or U2637 (N_2637,N_2187,N_2402);
nand U2638 (N_2638,N_2391,N_2399);
and U2639 (N_2639,N_2084,N_2345);
or U2640 (N_2640,N_2471,N_2088);
and U2641 (N_2641,N_2175,N_2458);
or U2642 (N_2642,N_2337,N_2397);
xor U2643 (N_2643,N_2101,N_2204);
nand U2644 (N_2644,N_2448,N_2343);
nor U2645 (N_2645,N_2484,N_2301);
or U2646 (N_2646,N_2103,N_2488);
nor U2647 (N_2647,N_2015,N_2407);
nand U2648 (N_2648,N_2134,N_2356);
or U2649 (N_2649,N_2048,N_2074);
and U2650 (N_2650,N_2423,N_2339);
and U2651 (N_2651,N_2465,N_2457);
or U2652 (N_2652,N_2479,N_2365);
nand U2653 (N_2653,N_2076,N_2256);
nand U2654 (N_2654,N_2060,N_2375);
or U2655 (N_2655,N_2273,N_2310);
and U2656 (N_2656,N_2030,N_2415);
nand U2657 (N_2657,N_2167,N_2433);
and U2658 (N_2658,N_2367,N_2265);
nor U2659 (N_2659,N_2149,N_2154);
and U2660 (N_2660,N_2057,N_2327);
and U2661 (N_2661,N_2364,N_2207);
or U2662 (N_2662,N_2251,N_2442);
nand U2663 (N_2663,N_2090,N_2352);
nor U2664 (N_2664,N_2436,N_2452);
and U2665 (N_2665,N_2019,N_2152);
or U2666 (N_2666,N_2419,N_2449);
nor U2667 (N_2667,N_2238,N_2010);
and U2668 (N_2668,N_2383,N_2206);
and U2669 (N_2669,N_2100,N_2409);
nor U2670 (N_2670,N_2064,N_2466);
or U2671 (N_2671,N_2163,N_2296);
nand U2672 (N_2672,N_2328,N_2306);
nand U2673 (N_2673,N_2406,N_2069);
nand U2674 (N_2674,N_2291,N_2041);
and U2675 (N_2675,N_2293,N_2097);
or U2676 (N_2676,N_2426,N_2007);
nand U2677 (N_2677,N_2051,N_2032);
or U2678 (N_2678,N_2080,N_2081);
nor U2679 (N_2679,N_2361,N_2234);
nand U2680 (N_2680,N_2430,N_2382);
and U2681 (N_2681,N_2062,N_2162);
nand U2682 (N_2682,N_2279,N_2098);
nand U2683 (N_2683,N_2420,N_2429);
nor U2684 (N_2684,N_2166,N_2262);
or U2685 (N_2685,N_2104,N_2275);
and U2686 (N_2686,N_2381,N_2226);
or U2687 (N_2687,N_2110,N_2172);
nand U2688 (N_2688,N_2414,N_2089);
nand U2689 (N_2689,N_2245,N_2444);
and U2690 (N_2690,N_2144,N_2230);
nor U2691 (N_2691,N_2334,N_2148);
nand U2692 (N_2692,N_2455,N_2294);
or U2693 (N_2693,N_2005,N_2141);
nand U2694 (N_2694,N_2497,N_2311);
and U2695 (N_2695,N_2225,N_2003);
nand U2696 (N_2696,N_2044,N_2213);
nor U2697 (N_2697,N_2349,N_2284);
nand U2698 (N_2698,N_2109,N_2400);
and U2699 (N_2699,N_2031,N_2492);
or U2700 (N_2700,N_2459,N_2014);
nor U2701 (N_2701,N_2186,N_2487);
or U2702 (N_2702,N_2018,N_2068);
or U2703 (N_2703,N_2410,N_2440);
and U2704 (N_2704,N_2476,N_2373);
or U2705 (N_2705,N_2380,N_2094);
nand U2706 (N_2706,N_2464,N_2155);
nand U2707 (N_2707,N_2202,N_2095);
or U2708 (N_2708,N_2199,N_2181);
nor U2709 (N_2709,N_2216,N_2480);
nor U2710 (N_2710,N_2358,N_2438);
nand U2711 (N_2711,N_2171,N_2425);
nor U2712 (N_2712,N_2200,N_2324);
or U2713 (N_2713,N_2354,N_2108);
or U2714 (N_2714,N_2428,N_2102);
nand U2715 (N_2715,N_2077,N_2142);
and U2716 (N_2716,N_2158,N_2376);
nand U2717 (N_2717,N_2189,N_2347);
or U2718 (N_2718,N_2413,N_2107);
and U2719 (N_2719,N_2405,N_2307);
nor U2720 (N_2720,N_2137,N_2357);
and U2721 (N_2721,N_2053,N_2106);
or U2722 (N_2722,N_2218,N_2059);
and U2723 (N_2723,N_2042,N_2131);
or U2724 (N_2724,N_2246,N_2282);
nand U2725 (N_2725,N_2229,N_2260);
nand U2726 (N_2726,N_2151,N_2219);
or U2727 (N_2727,N_2412,N_2130);
nand U2728 (N_2728,N_2392,N_2462);
and U2729 (N_2729,N_2190,N_2394);
nand U2730 (N_2730,N_2281,N_2424);
nand U2731 (N_2731,N_2001,N_2235);
xor U2732 (N_2732,N_2180,N_2233);
nand U2733 (N_2733,N_2176,N_2224);
nand U2734 (N_2734,N_2498,N_2160);
nand U2735 (N_2735,N_2316,N_2211);
nor U2736 (N_2736,N_2119,N_2344);
nor U2737 (N_2737,N_2450,N_2321);
or U2738 (N_2738,N_2221,N_2112);
nand U2739 (N_2739,N_2261,N_2145);
nand U2740 (N_2740,N_2043,N_2326);
nand U2741 (N_2741,N_2091,N_2403);
nand U2742 (N_2742,N_2208,N_2117);
nand U2743 (N_2743,N_2140,N_2478);
or U2744 (N_2744,N_2377,N_2363);
xnor U2745 (N_2745,N_2250,N_2008);
and U2746 (N_2746,N_2267,N_2325);
or U2747 (N_2747,N_2481,N_2170);
nor U2748 (N_2748,N_2473,N_2313);
and U2749 (N_2749,N_2247,N_2242);
nor U2750 (N_2750,N_2491,N_2296);
nand U2751 (N_2751,N_2279,N_2476);
and U2752 (N_2752,N_2110,N_2101);
and U2753 (N_2753,N_2283,N_2016);
nor U2754 (N_2754,N_2254,N_2424);
nand U2755 (N_2755,N_2483,N_2400);
and U2756 (N_2756,N_2228,N_2264);
nor U2757 (N_2757,N_2067,N_2305);
or U2758 (N_2758,N_2009,N_2401);
and U2759 (N_2759,N_2390,N_2202);
nor U2760 (N_2760,N_2373,N_2396);
and U2761 (N_2761,N_2408,N_2323);
nor U2762 (N_2762,N_2100,N_2124);
or U2763 (N_2763,N_2275,N_2493);
and U2764 (N_2764,N_2338,N_2204);
and U2765 (N_2765,N_2022,N_2197);
and U2766 (N_2766,N_2046,N_2425);
and U2767 (N_2767,N_2154,N_2256);
and U2768 (N_2768,N_2408,N_2360);
and U2769 (N_2769,N_2122,N_2227);
and U2770 (N_2770,N_2295,N_2340);
nor U2771 (N_2771,N_2220,N_2214);
and U2772 (N_2772,N_2213,N_2269);
nor U2773 (N_2773,N_2453,N_2391);
and U2774 (N_2774,N_2005,N_2328);
nor U2775 (N_2775,N_2362,N_2024);
and U2776 (N_2776,N_2374,N_2322);
nor U2777 (N_2777,N_2445,N_2332);
nand U2778 (N_2778,N_2303,N_2024);
or U2779 (N_2779,N_2479,N_2035);
nor U2780 (N_2780,N_2274,N_2384);
nand U2781 (N_2781,N_2197,N_2465);
nor U2782 (N_2782,N_2091,N_2267);
or U2783 (N_2783,N_2128,N_2097);
or U2784 (N_2784,N_2156,N_2482);
and U2785 (N_2785,N_2267,N_2042);
and U2786 (N_2786,N_2150,N_2153);
nor U2787 (N_2787,N_2476,N_2189);
or U2788 (N_2788,N_2225,N_2149);
or U2789 (N_2789,N_2389,N_2383);
and U2790 (N_2790,N_2307,N_2002);
nor U2791 (N_2791,N_2297,N_2113);
nand U2792 (N_2792,N_2113,N_2488);
nor U2793 (N_2793,N_2317,N_2412);
or U2794 (N_2794,N_2084,N_2488);
or U2795 (N_2795,N_2401,N_2311);
nor U2796 (N_2796,N_2088,N_2224);
and U2797 (N_2797,N_2103,N_2204);
and U2798 (N_2798,N_2290,N_2204);
nor U2799 (N_2799,N_2489,N_2049);
and U2800 (N_2800,N_2117,N_2307);
or U2801 (N_2801,N_2063,N_2144);
and U2802 (N_2802,N_2140,N_2006);
nor U2803 (N_2803,N_2108,N_2209);
and U2804 (N_2804,N_2445,N_2267);
and U2805 (N_2805,N_2406,N_2437);
and U2806 (N_2806,N_2013,N_2194);
nor U2807 (N_2807,N_2283,N_2365);
nor U2808 (N_2808,N_2209,N_2372);
nor U2809 (N_2809,N_2367,N_2144);
and U2810 (N_2810,N_2292,N_2367);
or U2811 (N_2811,N_2045,N_2254);
xnor U2812 (N_2812,N_2098,N_2028);
nand U2813 (N_2813,N_2192,N_2268);
and U2814 (N_2814,N_2163,N_2255);
or U2815 (N_2815,N_2401,N_2161);
nand U2816 (N_2816,N_2118,N_2088);
or U2817 (N_2817,N_2266,N_2015);
nand U2818 (N_2818,N_2443,N_2115);
and U2819 (N_2819,N_2299,N_2090);
nand U2820 (N_2820,N_2168,N_2144);
nor U2821 (N_2821,N_2460,N_2170);
nand U2822 (N_2822,N_2392,N_2073);
and U2823 (N_2823,N_2326,N_2191);
nor U2824 (N_2824,N_2080,N_2013);
and U2825 (N_2825,N_2372,N_2268);
nand U2826 (N_2826,N_2463,N_2156);
or U2827 (N_2827,N_2387,N_2162);
nor U2828 (N_2828,N_2439,N_2064);
nor U2829 (N_2829,N_2055,N_2254);
and U2830 (N_2830,N_2224,N_2029);
nand U2831 (N_2831,N_2144,N_2251);
nor U2832 (N_2832,N_2332,N_2132);
and U2833 (N_2833,N_2316,N_2100);
and U2834 (N_2834,N_2357,N_2188);
nand U2835 (N_2835,N_2054,N_2267);
nand U2836 (N_2836,N_2164,N_2079);
nor U2837 (N_2837,N_2083,N_2095);
nor U2838 (N_2838,N_2045,N_2448);
or U2839 (N_2839,N_2118,N_2300);
or U2840 (N_2840,N_2055,N_2247);
nand U2841 (N_2841,N_2401,N_2469);
nor U2842 (N_2842,N_2005,N_2404);
nor U2843 (N_2843,N_2324,N_2488);
and U2844 (N_2844,N_2333,N_2344);
nor U2845 (N_2845,N_2014,N_2436);
nor U2846 (N_2846,N_2111,N_2084);
or U2847 (N_2847,N_2441,N_2473);
and U2848 (N_2848,N_2488,N_2214);
nor U2849 (N_2849,N_2336,N_2024);
nand U2850 (N_2850,N_2349,N_2446);
and U2851 (N_2851,N_2020,N_2273);
nand U2852 (N_2852,N_2476,N_2315);
and U2853 (N_2853,N_2439,N_2290);
or U2854 (N_2854,N_2127,N_2169);
and U2855 (N_2855,N_2189,N_2394);
or U2856 (N_2856,N_2106,N_2100);
nor U2857 (N_2857,N_2350,N_2360);
nor U2858 (N_2858,N_2267,N_2348);
nand U2859 (N_2859,N_2207,N_2490);
nor U2860 (N_2860,N_2130,N_2165);
or U2861 (N_2861,N_2384,N_2249);
nor U2862 (N_2862,N_2295,N_2177);
nand U2863 (N_2863,N_2158,N_2033);
nor U2864 (N_2864,N_2048,N_2421);
nor U2865 (N_2865,N_2433,N_2129);
and U2866 (N_2866,N_2219,N_2083);
nor U2867 (N_2867,N_2294,N_2013);
or U2868 (N_2868,N_2436,N_2435);
nand U2869 (N_2869,N_2315,N_2354);
or U2870 (N_2870,N_2076,N_2187);
nor U2871 (N_2871,N_2206,N_2214);
or U2872 (N_2872,N_2256,N_2214);
nor U2873 (N_2873,N_2186,N_2195);
nor U2874 (N_2874,N_2476,N_2168);
nor U2875 (N_2875,N_2462,N_2218);
nand U2876 (N_2876,N_2470,N_2152);
nand U2877 (N_2877,N_2251,N_2258);
nor U2878 (N_2878,N_2250,N_2126);
or U2879 (N_2879,N_2062,N_2430);
nand U2880 (N_2880,N_2459,N_2423);
nand U2881 (N_2881,N_2125,N_2153);
and U2882 (N_2882,N_2482,N_2431);
nor U2883 (N_2883,N_2490,N_2066);
or U2884 (N_2884,N_2253,N_2060);
and U2885 (N_2885,N_2437,N_2384);
or U2886 (N_2886,N_2478,N_2401);
nand U2887 (N_2887,N_2048,N_2209);
and U2888 (N_2888,N_2314,N_2310);
or U2889 (N_2889,N_2398,N_2105);
and U2890 (N_2890,N_2304,N_2379);
and U2891 (N_2891,N_2351,N_2180);
nand U2892 (N_2892,N_2098,N_2327);
and U2893 (N_2893,N_2421,N_2319);
and U2894 (N_2894,N_2027,N_2365);
nand U2895 (N_2895,N_2255,N_2149);
nor U2896 (N_2896,N_2339,N_2006);
or U2897 (N_2897,N_2197,N_2114);
nor U2898 (N_2898,N_2111,N_2091);
and U2899 (N_2899,N_2277,N_2203);
or U2900 (N_2900,N_2491,N_2184);
nor U2901 (N_2901,N_2091,N_2494);
and U2902 (N_2902,N_2060,N_2258);
or U2903 (N_2903,N_2485,N_2415);
xnor U2904 (N_2904,N_2237,N_2358);
or U2905 (N_2905,N_2066,N_2017);
or U2906 (N_2906,N_2278,N_2412);
nand U2907 (N_2907,N_2393,N_2305);
nor U2908 (N_2908,N_2103,N_2337);
nand U2909 (N_2909,N_2068,N_2107);
or U2910 (N_2910,N_2191,N_2323);
nand U2911 (N_2911,N_2129,N_2062);
nor U2912 (N_2912,N_2271,N_2255);
and U2913 (N_2913,N_2008,N_2289);
or U2914 (N_2914,N_2252,N_2441);
and U2915 (N_2915,N_2299,N_2274);
or U2916 (N_2916,N_2185,N_2122);
or U2917 (N_2917,N_2009,N_2448);
nor U2918 (N_2918,N_2368,N_2096);
nand U2919 (N_2919,N_2115,N_2378);
nor U2920 (N_2920,N_2060,N_2164);
or U2921 (N_2921,N_2170,N_2270);
nand U2922 (N_2922,N_2366,N_2049);
nand U2923 (N_2923,N_2125,N_2286);
nor U2924 (N_2924,N_2052,N_2490);
nor U2925 (N_2925,N_2373,N_2247);
nand U2926 (N_2926,N_2162,N_2285);
nor U2927 (N_2927,N_2068,N_2307);
nand U2928 (N_2928,N_2032,N_2368);
nand U2929 (N_2929,N_2022,N_2084);
nand U2930 (N_2930,N_2138,N_2398);
nand U2931 (N_2931,N_2264,N_2273);
nand U2932 (N_2932,N_2171,N_2481);
or U2933 (N_2933,N_2132,N_2215);
nor U2934 (N_2934,N_2463,N_2236);
nand U2935 (N_2935,N_2301,N_2363);
nand U2936 (N_2936,N_2127,N_2484);
nand U2937 (N_2937,N_2430,N_2441);
or U2938 (N_2938,N_2371,N_2201);
nor U2939 (N_2939,N_2127,N_2475);
nor U2940 (N_2940,N_2065,N_2486);
or U2941 (N_2941,N_2004,N_2023);
nand U2942 (N_2942,N_2128,N_2390);
and U2943 (N_2943,N_2174,N_2257);
nand U2944 (N_2944,N_2132,N_2075);
or U2945 (N_2945,N_2089,N_2172);
or U2946 (N_2946,N_2106,N_2125);
or U2947 (N_2947,N_2222,N_2396);
nor U2948 (N_2948,N_2313,N_2102);
or U2949 (N_2949,N_2277,N_2030);
nand U2950 (N_2950,N_2479,N_2394);
and U2951 (N_2951,N_2119,N_2353);
or U2952 (N_2952,N_2299,N_2352);
nor U2953 (N_2953,N_2396,N_2387);
nor U2954 (N_2954,N_2241,N_2377);
nor U2955 (N_2955,N_2329,N_2061);
and U2956 (N_2956,N_2257,N_2250);
and U2957 (N_2957,N_2137,N_2337);
nand U2958 (N_2958,N_2472,N_2074);
or U2959 (N_2959,N_2389,N_2479);
nor U2960 (N_2960,N_2265,N_2398);
nor U2961 (N_2961,N_2470,N_2255);
or U2962 (N_2962,N_2487,N_2456);
nor U2963 (N_2963,N_2348,N_2286);
nor U2964 (N_2964,N_2070,N_2439);
or U2965 (N_2965,N_2142,N_2355);
and U2966 (N_2966,N_2346,N_2045);
nor U2967 (N_2967,N_2457,N_2066);
or U2968 (N_2968,N_2024,N_2114);
and U2969 (N_2969,N_2207,N_2035);
nor U2970 (N_2970,N_2407,N_2061);
and U2971 (N_2971,N_2404,N_2450);
and U2972 (N_2972,N_2244,N_2085);
or U2973 (N_2973,N_2279,N_2227);
and U2974 (N_2974,N_2299,N_2321);
nand U2975 (N_2975,N_2084,N_2414);
xor U2976 (N_2976,N_2014,N_2122);
and U2977 (N_2977,N_2370,N_2193);
and U2978 (N_2978,N_2355,N_2100);
nor U2979 (N_2979,N_2377,N_2175);
nand U2980 (N_2980,N_2407,N_2296);
and U2981 (N_2981,N_2001,N_2175);
or U2982 (N_2982,N_2436,N_2486);
nand U2983 (N_2983,N_2252,N_2296);
and U2984 (N_2984,N_2463,N_2294);
or U2985 (N_2985,N_2423,N_2224);
nor U2986 (N_2986,N_2066,N_2093);
nor U2987 (N_2987,N_2375,N_2475);
nand U2988 (N_2988,N_2074,N_2041);
or U2989 (N_2989,N_2093,N_2006);
nor U2990 (N_2990,N_2401,N_2299);
or U2991 (N_2991,N_2254,N_2410);
or U2992 (N_2992,N_2254,N_2113);
xnor U2993 (N_2993,N_2460,N_2052);
nand U2994 (N_2994,N_2267,N_2097);
nor U2995 (N_2995,N_2342,N_2427);
nand U2996 (N_2996,N_2176,N_2361);
and U2997 (N_2997,N_2178,N_2311);
and U2998 (N_2998,N_2370,N_2220);
and U2999 (N_2999,N_2447,N_2255);
and U3000 (N_3000,N_2697,N_2821);
or U3001 (N_3001,N_2862,N_2897);
and U3002 (N_3002,N_2680,N_2551);
and U3003 (N_3003,N_2800,N_2503);
or U3004 (N_3004,N_2738,N_2568);
nor U3005 (N_3005,N_2716,N_2705);
nor U3006 (N_3006,N_2507,N_2781);
nand U3007 (N_3007,N_2855,N_2732);
nor U3008 (N_3008,N_2749,N_2943);
xnor U3009 (N_3009,N_2506,N_2779);
and U3010 (N_3010,N_2720,N_2901);
or U3011 (N_3011,N_2539,N_2528);
and U3012 (N_3012,N_2561,N_2964);
nand U3013 (N_3013,N_2547,N_2988);
nand U3014 (N_3014,N_2751,N_2755);
nor U3015 (N_3015,N_2757,N_2559);
nand U3016 (N_3016,N_2642,N_2954);
and U3017 (N_3017,N_2876,N_2823);
or U3018 (N_3018,N_2937,N_2887);
nand U3019 (N_3019,N_2583,N_2521);
nor U3020 (N_3020,N_2871,N_2625);
or U3021 (N_3021,N_2996,N_2917);
and U3022 (N_3022,N_2812,N_2604);
nor U3023 (N_3023,N_2577,N_2935);
and U3024 (N_3024,N_2828,N_2985);
nand U3025 (N_3025,N_2817,N_2692);
nand U3026 (N_3026,N_2574,N_2919);
nor U3027 (N_3027,N_2589,N_2508);
nand U3028 (N_3028,N_2960,N_2696);
or U3029 (N_3029,N_2957,N_2603);
and U3030 (N_3030,N_2984,N_2562);
and U3031 (N_3031,N_2729,N_2632);
nor U3032 (N_3032,N_2759,N_2747);
and U3033 (N_3033,N_2592,N_2861);
or U3034 (N_3034,N_2644,N_2804);
nand U3035 (N_3035,N_2573,N_2612);
nand U3036 (N_3036,N_2633,N_2989);
nand U3037 (N_3037,N_2753,N_2693);
nand U3038 (N_3038,N_2906,N_2504);
or U3039 (N_3039,N_2654,N_2582);
nor U3040 (N_3040,N_2646,N_2510);
nor U3041 (N_3041,N_2649,N_2616);
or U3042 (N_3042,N_2967,N_2997);
and U3043 (N_3043,N_2514,N_2842);
or U3044 (N_3044,N_2647,N_2601);
nand U3045 (N_3045,N_2548,N_2859);
nand U3046 (N_3046,N_2634,N_2814);
nor U3047 (N_3047,N_2735,N_2623);
nand U3048 (N_3048,N_2681,N_2927);
nand U3049 (N_3049,N_2678,N_2570);
nor U3050 (N_3050,N_2844,N_2666);
or U3051 (N_3051,N_2950,N_2768);
nor U3052 (N_3052,N_2933,N_2813);
and U3053 (N_3053,N_2934,N_2593);
and U3054 (N_3054,N_2661,N_2590);
nor U3055 (N_3055,N_2686,N_2707);
nand U3056 (N_3056,N_2882,N_2806);
or U3057 (N_3057,N_2762,N_2752);
or U3058 (N_3058,N_2908,N_2580);
nor U3059 (N_3059,N_2797,N_2888);
nand U3060 (N_3060,N_2667,N_2522);
and U3061 (N_3061,N_2785,N_2879);
nor U3062 (N_3062,N_2520,N_2530);
or U3063 (N_3063,N_2874,N_2981);
nand U3064 (N_3064,N_2941,N_2698);
or U3065 (N_3065,N_2763,N_2650);
nand U3066 (N_3066,N_2827,N_2926);
and U3067 (N_3067,N_2519,N_2717);
nor U3068 (N_3068,N_2911,N_2918);
xor U3069 (N_3069,N_2760,N_2578);
nand U3070 (N_3070,N_2587,N_2585);
nor U3071 (N_3071,N_2833,N_2898);
or U3072 (N_3072,N_2677,N_2944);
or U3073 (N_3073,N_2536,N_2659);
nand U3074 (N_3074,N_2959,N_2816);
or U3075 (N_3075,N_2932,N_2973);
nor U3076 (N_3076,N_2841,N_2711);
nor U3077 (N_3077,N_2907,N_2565);
and U3078 (N_3078,N_2775,N_2538);
xor U3079 (N_3079,N_2974,N_2928);
nor U3080 (N_3080,N_2792,N_2743);
nand U3081 (N_3081,N_2610,N_2533);
or U3082 (N_3082,N_2754,N_2982);
nand U3083 (N_3083,N_2839,N_2893);
nand U3084 (N_3084,N_2830,N_2790);
or U3085 (N_3085,N_2791,N_2535);
or U3086 (N_3086,N_2664,N_2892);
and U3087 (N_3087,N_2750,N_2772);
and U3088 (N_3088,N_2783,N_2673);
nor U3089 (N_3089,N_2836,N_2668);
and U3090 (N_3090,N_2727,N_2736);
nand U3091 (N_3091,N_2701,N_2730);
nand U3092 (N_3092,N_2709,N_2767);
nor U3093 (N_3093,N_2811,N_2948);
and U3094 (N_3094,N_2739,N_2682);
and U3095 (N_3095,N_2611,N_2877);
and U3096 (N_3096,N_2965,N_2929);
and U3097 (N_3097,N_2569,N_2558);
nor U3098 (N_3098,N_2872,N_2713);
or U3099 (N_3099,N_2626,N_2605);
and U3100 (N_3100,N_2665,N_2870);
nor U3101 (N_3101,N_2902,N_2986);
or U3102 (N_3102,N_2572,N_2949);
nand U3103 (N_3103,N_2869,N_2955);
or U3104 (N_3104,N_2660,N_2995);
or U3105 (N_3105,N_2845,N_2849);
or U3106 (N_3106,N_2607,N_2624);
nor U3107 (N_3107,N_2596,N_2599);
nand U3108 (N_3108,N_2600,N_2915);
or U3109 (N_3109,N_2773,N_2598);
and U3110 (N_3110,N_2904,N_2545);
and U3111 (N_3111,N_2653,N_2971);
and U3112 (N_3112,N_2723,N_2787);
nor U3113 (N_3113,N_2648,N_2631);
and U3114 (N_3114,N_2771,N_2684);
nand U3115 (N_3115,N_2541,N_2881);
or U3116 (N_3116,N_2591,N_2586);
or U3117 (N_3117,N_2880,N_2978);
nor U3118 (N_3118,N_2966,N_2801);
or U3119 (N_3119,N_2962,N_2746);
nor U3120 (N_3120,N_2993,N_2658);
or U3121 (N_3121,N_2655,N_2809);
nand U3122 (N_3122,N_2972,N_2714);
or U3123 (N_3123,N_2890,N_2706);
or U3124 (N_3124,N_2595,N_2776);
and U3125 (N_3125,N_2529,N_2617);
and U3126 (N_3126,N_2540,N_2704);
nor U3127 (N_3127,N_2818,N_2778);
or U3128 (N_3128,N_2774,N_2835);
and U3129 (N_3129,N_2525,N_2857);
and U3130 (N_3130,N_2737,N_2884);
and U3131 (N_3131,N_2721,N_2712);
or U3132 (N_3132,N_2761,N_2687);
or U3133 (N_3133,N_2537,N_2936);
and U3134 (N_3134,N_2685,N_2501);
and U3135 (N_3135,N_2724,N_2777);
nor U3136 (N_3136,N_2819,N_2575);
or U3137 (N_3137,N_2883,N_2858);
nand U3138 (N_3138,N_2756,N_2769);
nand U3139 (N_3139,N_2891,N_2793);
nor U3140 (N_3140,N_2983,N_2909);
or U3141 (N_3141,N_2715,N_2636);
nand U3142 (N_3142,N_2571,N_2651);
nand U3143 (N_3143,N_2848,N_2745);
and U3144 (N_3144,N_2670,N_2832);
and U3145 (N_3145,N_2780,N_2500);
and U3146 (N_3146,N_2675,N_2924);
or U3147 (N_3147,N_2826,N_2843);
nor U3148 (N_3148,N_2534,N_2786);
nor U3149 (N_3149,N_2979,N_2896);
or U3150 (N_3150,N_2822,N_2554);
and U3151 (N_3151,N_2663,N_2657);
nor U3152 (N_3152,N_2863,N_2576);
nand U3153 (N_3153,N_2690,N_2921);
and U3154 (N_3154,N_2951,N_2674);
nor U3155 (N_3155,N_2688,N_2563);
nand U3156 (N_3156,N_2608,N_2900);
or U3157 (N_3157,N_2992,N_2679);
or U3158 (N_3158,N_2628,N_2940);
nand U3159 (N_3159,N_2799,N_2878);
or U3160 (N_3160,N_2639,N_2526);
or U3161 (N_3161,N_2731,N_2810);
nand U3162 (N_3162,N_2524,N_2990);
nand U3163 (N_3163,N_2868,N_2546);
nor U3164 (N_3164,N_2567,N_2853);
nand U3165 (N_3165,N_2805,N_2629);
and U3166 (N_3166,N_2837,N_2764);
or U3167 (N_3167,N_2795,N_2511);
and U3168 (N_3168,N_2856,N_2922);
or U3169 (N_3169,N_2635,N_2829);
and U3170 (N_3170,N_2718,N_2584);
or U3171 (N_3171,N_2512,N_2505);
or U3172 (N_3172,N_2912,N_2834);
xnor U3173 (N_3173,N_2784,N_2854);
and U3174 (N_3174,N_2947,N_2980);
nand U3175 (N_3175,N_2825,N_2945);
nand U3176 (N_3176,N_2613,N_2553);
or U3177 (N_3177,N_2831,N_2676);
nand U3178 (N_3178,N_2758,N_2850);
or U3179 (N_3179,N_2549,N_2741);
nor U3180 (N_3180,N_2923,N_2588);
nand U3181 (N_3181,N_2998,N_2630);
or U3182 (N_3182,N_2637,N_2914);
and U3183 (N_3183,N_2700,N_2977);
xor U3184 (N_3184,N_2952,N_2838);
nand U3185 (N_3185,N_2953,N_2894);
or U3186 (N_3186,N_2770,N_2939);
nand U3187 (N_3187,N_2691,N_2802);
or U3188 (N_3188,N_2581,N_2815);
or U3189 (N_3189,N_2544,N_2734);
xnor U3190 (N_3190,N_2788,N_2566);
or U3191 (N_3191,N_2864,N_2671);
and U3192 (N_3192,N_2987,N_2557);
or U3193 (N_3193,N_2643,N_2641);
nor U3194 (N_3194,N_2638,N_2527);
or U3195 (N_3195,N_2963,N_2920);
nand U3196 (N_3196,N_2695,N_2803);
nand U3197 (N_3197,N_2689,N_2683);
nand U3198 (N_3198,N_2615,N_2913);
nand U3199 (N_3199,N_2961,N_2885);
nand U3200 (N_3200,N_2550,N_2846);
nand U3201 (N_3201,N_2930,N_2502);
and U3202 (N_3202,N_2725,N_2652);
nor U3203 (N_3203,N_2710,N_2820);
nor U3204 (N_3204,N_2609,N_2620);
and U3205 (N_3205,N_2602,N_2999);
nor U3206 (N_3206,N_2708,N_2532);
and U3207 (N_3207,N_2969,N_2728);
nand U3208 (N_3208,N_2621,N_2765);
and U3209 (N_3209,N_2824,N_2614);
nor U3210 (N_3210,N_2852,N_2873);
nor U3211 (N_3211,N_2956,N_2662);
or U3212 (N_3212,N_2694,N_2840);
and U3213 (N_3213,N_2606,N_2543);
or U3214 (N_3214,N_2627,N_2807);
nor U3215 (N_3215,N_2968,N_2640);
and U3216 (N_3216,N_2867,N_2847);
or U3217 (N_3217,N_2703,N_2931);
nand U3218 (N_3218,N_2560,N_2740);
nor U3219 (N_3219,N_2903,N_2656);
and U3220 (N_3220,N_2975,N_2513);
nand U3221 (N_3221,N_2579,N_2672);
or U3222 (N_3222,N_2991,N_2744);
or U3223 (N_3223,N_2886,N_2899);
and U3224 (N_3224,N_2925,N_2794);
nand U3225 (N_3225,N_2564,N_2622);
nor U3226 (N_3226,N_2875,N_2942);
nand U3227 (N_3227,N_2895,N_2748);
or U3228 (N_3228,N_2509,N_2618);
and U3229 (N_3229,N_2889,N_2958);
or U3230 (N_3230,N_2865,N_2523);
and U3231 (N_3231,N_2702,N_2976);
nand U3232 (N_3232,N_2542,N_2726);
nor U3233 (N_3233,N_2851,N_2515);
and U3234 (N_3234,N_2905,N_2866);
or U3235 (N_3235,N_2719,N_2645);
and U3236 (N_3236,N_2594,N_2597);
and U3237 (N_3237,N_2742,N_2798);
nand U3238 (N_3238,N_2910,N_2516);
nand U3239 (N_3239,N_2970,N_2733);
nand U3240 (N_3240,N_2555,N_2789);
and U3241 (N_3241,N_2531,N_2699);
nand U3242 (N_3242,N_2556,N_2552);
and U3243 (N_3243,N_2722,N_2517);
or U3244 (N_3244,N_2766,N_2518);
and U3245 (N_3245,N_2946,N_2619);
nor U3246 (N_3246,N_2860,N_2782);
or U3247 (N_3247,N_2796,N_2669);
nor U3248 (N_3248,N_2938,N_2916);
nor U3249 (N_3249,N_2994,N_2808);
and U3250 (N_3250,N_2529,N_2600);
xnor U3251 (N_3251,N_2760,N_2720);
or U3252 (N_3252,N_2783,N_2694);
nand U3253 (N_3253,N_2964,N_2779);
nor U3254 (N_3254,N_2613,N_2864);
nand U3255 (N_3255,N_2832,N_2708);
or U3256 (N_3256,N_2524,N_2719);
or U3257 (N_3257,N_2895,N_2728);
or U3258 (N_3258,N_2661,N_2994);
nand U3259 (N_3259,N_2691,N_2686);
nor U3260 (N_3260,N_2842,N_2638);
nor U3261 (N_3261,N_2668,N_2504);
nand U3262 (N_3262,N_2902,N_2557);
nor U3263 (N_3263,N_2712,N_2774);
or U3264 (N_3264,N_2670,N_2831);
or U3265 (N_3265,N_2781,N_2708);
or U3266 (N_3266,N_2616,N_2814);
nand U3267 (N_3267,N_2949,N_2766);
nor U3268 (N_3268,N_2841,N_2784);
nor U3269 (N_3269,N_2776,N_2828);
nand U3270 (N_3270,N_2730,N_2577);
nor U3271 (N_3271,N_2554,N_2540);
and U3272 (N_3272,N_2707,N_2554);
nand U3273 (N_3273,N_2709,N_2539);
nand U3274 (N_3274,N_2800,N_2526);
nor U3275 (N_3275,N_2888,N_2679);
and U3276 (N_3276,N_2524,N_2906);
or U3277 (N_3277,N_2974,N_2727);
or U3278 (N_3278,N_2809,N_2644);
nor U3279 (N_3279,N_2669,N_2881);
and U3280 (N_3280,N_2644,N_2737);
and U3281 (N_3281,N_2730,N_2510);
nor U3282 (N_3282,N_2712,N_2594);
nand U3283 (N_3283,N_2971,N_2696);
or U3284 (N_3284,N_2731,N_2619);
nor U3285 (N_3285,N_2604,N_2736);
nor U3286 (N_3286,N_2726,N_2973);
or U3287 (N_3287,N_2819,N_2714);
nand U3288 (N_3288,N_2563,N_2826);
nand U3289 (N_3289,N_2986,N_2725);
nor U3290 (N_3290,N_2936,N_2865);
nand U3291 (N_3291,N_2675,N_2746);
nand U3292 (N_3292,N_2565,N_2707);
nor U3293 (N_3293,N_2948,N_2965);
and U3294 (N_3294,N_2985,N_2768);
or U3295 (N_3295,N_2561,N_2583);
nand U3296 (N_3296,N_2784,N_2926);
nand U3297 (N_3297,N_2948,N_2785);
or U3298 (N_3298,N_2807,N_2669);
and U3299 (N_3299,N_2832,N_2776);
nor U3300 (N_3300,N_2982,N_2873);
or U3301 (N_3301,N_2757,N_2669);
nor U3302 (N_3302,N_2789,N_2625);
or U3303 (N_3303,N_2909,N_2984);
nand U3304 (N_3304,N_2948,N_2908);
nand U3305 (N_3305,N_2589,N_2715);
nor U3306 (N_3306,N_2658,N_2995);
and U3307 (N_3307,N_2569,N_2584);
and U3308 (N_3308,N_2819,N_2775);
and U3309 (N_3309,N_2775,N_2659);
and U3310 (N_3310,N_2709,N_2644);
and U3311 (N_3311,N_2690,N_2781);
and U3312 (N_3312,N_2566,N_2740);
nor U3313 (N_3313,N_2687,N_2815);
nand U3314 (N_3314,N_2908,N_2681);
nand U3315 (N_3315,N_2519,N_2508);
and U3316 (N_3316,N_2790,N_2746);
nand U3317 (N_3317,N_2892,N_2541);
and U3318 (N_3318,N_2730,N_2797);
nor U3319 (N_3319,N_2756,N_2947);
and U3320 (N_3320,N_2940,N_2786);
or U3321 (N_3321,N_2651,N_2580);
nand U3322 (N_3322,N_2723,N_2679);
or U3323 (N_3323,N_2864,N_2656);
nand U3324 (N_3324,N_2920,N_2849);
nor U3325 (N_3325,N_2861,N_2631);
and U3326 (N_3326,N_2823,N_2696);
nor U3327 (N_3327,N_2784,N_2613);
or U3328 (N_3328,N_2780,N_2854);
xor U3329 (N_3329,N_2747,N_2926);
and U3330 (N_3330,N_2694,N_2673);
or U3331 (N_3331,N_2887,N_2561);
or U3332 (N_3332,N_2762,N_2759);
nand U3333 (N_3333,N_2550,N_2903);
or U3334 (N_3334,N_2994,N_2634);
and U3335 (N_3335,N_2995,N_2712);
nand U3336 (N_3336,N_2899,N_2575);
and U3337 (N_3337,N_2780,N_2701);
nand U3338 (N_3338,N_2863,N_2548);
and U3339 (N_3339,N_2954,N_2969);
nor U3340 (N_3340,N_2509,N_2646);
nor U3341 (N_3341,N_2973,N_2873);
nand U3342 (N_3342,N_2995,N_2734);
or U3343 (N_3343,N_2538,N_2644);
nand U3344 (N_3344,N_2763,N_2620);
nand U3345 (N_3345,N_2956,N_2692);
nor U3346 (N_3346,N_2572,N_2701);
nand U3347 (N_3347,N_2518,N_2680);
and U3348 (N_3348,N_2513,N_2755);
and U3349 (N_3349,N_2882,N_2508);
nor U3350 (N_3350,N_2510,N_2597);
nand U3351 (N_3351,N_2580,N_2846);
or U3352 (N_3352,N_2513,N_2614);
nor U3353 (N_3353,N_2511,N_2986);
or U3354 (N_3354,N_2588,N_2762);
nand U3355 (N_3355,N_2507,N_2571);
and U3356 (N_3356,N_2651,N_2621);
and U3357 (N_3357,N_2616,N_2613);
nor U3358 (N_3358,N_2910,N_2909);
nor U3359 (N_3359,N_2792,N_2593);
or U3360 (N_3360,N_2709,N_2771);
or U3361 (N_3361,N_2877,N_2551);
and U3362 (N_3362,N_2728,N_2567);
and U3363 (N_3363,N_2904,N_2566);
and U3364 (N_3364,N_2615,N_2916);
and U3365 (N_3365,N_2735,N_2743);
or U3366 (N_3366,N_2866,N_2600);
nand U3367 (N_3367,N_2982,N_2592);
nand U3368 (N_3368,N_2661,N_2891);
and U3369 (N_3369,N_2873,N_2752);
and U3370 (N_3370,N_2589,N_2679);
or U3371 (N_3371,N_2749,N_2812);
or U3372 (N_3372,N_2643,N_2630);
or U3373 (N_3373,N_2999,N_2691);
nor U3374 (N_3374,N_2664,N_2513);
nand U3375 (N_3375,N_2631,N_2876);
nand U3376 (N_3376,N_2899,N_2806);
nand U3377 (N_3377,N_2883,N_2985);
or U3378 (N_3378,N_2760,N_2529);
or U3379 (N_3379,N_2790,N_2905);
nand U3380 (N_3380,N_2512,N_2741);
or U3381 (N_3381,N_2600,N_2873);
nand U3382 (N_3382,N_2942,N_2878);
or U3383 (N_3383,N_2547,N_2688);
or U3384 (N_3384,N_2841,N_2760);
or U3385 (N_3385,N_2536,N_2556);
nor U3386 (N_3386,N_2811,N_2853);
and U3387 (N_3387,N_2791,N_2534);
and U3388 (N_3388,N_2891,N_2503);
nand U3389 (N_3389,N_2544,N_2516);
or U3390 (N_3390,N_2551,N_2956);
and U3391 (N_3391,N_2772,N_2872);
and U3392 (N_3392,N_2770,N_2643);
nor U3393 (N_3393,N_2561,N_2659);
nor U3394 (N_3394,N_2750,N_2986);
nor U3395 (N_3395,N_2502,N_2766);
nor U3396 (N_3396,N_2540,N_2598);
nand U3397 (N_3397,N_2821,N_2722);
or U3398 (N_3398,N_2879,N_2609);
and U3399 (N_3399,N_2515,N_2773);
and U3400 (N_3400,N_2736,N_2504);
nand U3401 (N_3401,N_2839,N_2525);
nand U3402 (N_3402,N_2599,N_2738);
and U3403 (N_3403,N_2948,N_2900);
nand U3404 (N_3404,N_2576,N_2853);
nand U3405 (N_3405,N_2966,N_2644);
nor U3406 (N_3406,N_2830,N_2702);
nor U3407 (N_3407,N_2715,N_2603);
or U3408 (N_3408,N_2772,N_2963);
and U3409 (N_3409,N_2793,N_2698);
nor U3410 (N_3410,N_2935,N_2893);
xnor U3411 (N_3411,N_2554,N_2737);
or U3412 (N_3412,N_2895,N_2501);
nand U3413 (N_3413,N_2748,N_2687);
nand U3414 (N_3414,N_2770,N_2869);
and U3415 (N_3415,N_2853,N_2915);
and U3416 (N_3416,N_2709,N_2807);
nand U3417 (N_3417,N_2849,N_2800);
nand U3418 (N_3418,N_2685,N_2955);
nor U3419 (N_3419,N_2574,N_2757);
and U3420 (N_3420,N_2735,N_2674);
or U3421 (N_3421,N_2995,N_2965);
and U3422 (N_3422,N_2990,N_2896);
nor U3423 (N_3423,N_2815,N_2559);
or U3424 (N_3424,N_2719,N_2688);
and U3425 (N_3425,N_2610,N_2793);
and U3426 (N_3426,N_2515,N_2612);
nand U3427 (N_3427,N_2693,N_2864);
or U3428 (N_3428,N_2531,N_2760);
and U3429 (N_3429,N_2729,N_2610);
nor U3430 (N_3430,N_2583,N_2854);
or U3431 (N_3431,N_2750,N_2506);
nand U3432 (N_3432,N_2812,N_2926);
nor U3433 (N_3433,N_2916,N_2510);
nor U3434 (N_3434,N_2591,N_2946);
and U3435 (N_3435,N_2825,N_2741);
and U3436 (N_3436,N_2966,N_2584);
nand U3437 (N_3437,N_2924,N_2757);
and U3438 (N_3438,N_2777,N_2603);
or U3439 (N_3439,N_2666,N_2789);
nand U3440 (N_3440,N_2832,N_2558);
nor U3441 (N_3441,N_2687,N_2851);
and U3442 (N_3442,N_2507,N_2653);
and U3443 (N_3443,N_2789,N_2641);
nor U3444 (N_3444,N_2755,N_2594);
nor U3445 (N_3445,N_2514,N_2682);
nand U3446 (N_3446,N_2571,N_2728);
nor U3447 (N_3447,N_2743,N_2887);
and U3448 (N_3448,N_2781,N_2767);
xnor U3449 (N_3449,N_2987,N_2817);
and U3450 (N_3450,N_2793,N_2615);
nor U3451 (N_3451,N_2628,N_2542);
nand U3452 (N_3452,N_2582,N_2736);
nor U3453 (N_3453,N_2649,N_2838);
and U3454 (N_3454,N_2799,N_2960);
and U3455 (N_3455,N_2877,N_2732);
nand U3456 (N_3456,N_2563,N_2622);
nor U3457 (N_3457,N_2880,N_2694);
or U3458 (N_3458,N_2630,N_2963);
nor U3459 (N_3459,N_2891,N_2577);
and U3460 (N_3460,N_2548,N_2958);
nand U3461 (N_3461,N_2714,N_2547);
and U3462 (N_3462,N_2988,N_2630);
nand U3463 (N_3463,N_2716,N_2905);
and U3464 (N_3464,N_2683,N_2844);
nor U3465 (N_3465,N_2934,N_2502);
or U3466 (N_3466,N_2968,N_2542);
nand U3467 (N_3467,N_2936,N_2606);
and U3468 (N_3468,N_2758,N_2856);
or U3469 (N_3469,N_2808,N_2745);
nor U3470 (N_3470,N_2934,N_2804);
or U3471 (N_3471,N_2721,N_2807);
nor U3472 (N_3472,N_2537,N_2784);
nor U3473 (N_3473,N_2617,N_2805);
and U3474 (N_3474,N_2502,N_2896);
nand U3475 (N_3475,N_2557,N_2931);
and U3476 (N_3476,N_2966,N_2626);
and U3477 (N_3477,N_2520,N_2804);
nor U3478 (N_3478,N_2548,N_2547);
or U3479 (N_3479,N_2975,N_2841);
nor U3480 (N_3480,N_2546,N_2913);
nor U3481 (N_3481,N_2548,N_2522);
nand U3482 (N_3482,N_2774,N_2721);
and U3483 (N_3483,N_2944,N_2546);
and U3484 (N_3484,N_2948,N_2802);
or U3485 (N_3485,N_2874,N_2510);
nor U3486 (N_3486,N_2707,N_2763);
and U3487 (N_3487,N_2861,N_2532);
nand U3488 (N_3488,N_2854,N_2597);
or U3489 (N_3489,N_2712,N_2950);
and U3490 (N_3490,N_2670,N_2503);
and U3491 (N_3491,N_2552,N_2743);
and U3492 (N_3492,N_2860,N_2931);
nand U3493 (N_3493,N_2533,N_2963);
or U3494 (N_3494,N_2732,N_2931);
or U3495 (N_3495,N_2564,N_2796);
nand U3496 (N_3496,N_2862,N_2872);
and U3497 (N_3497,N_2545,N_2699);
nand U3498 (N_3498,N_2891,N_2511);
or U3499 (N_3499,N_2567,N_2731);
nor U3500 (N_3500,N_3232,N_3098);
nor U3501 (N_3501,N_3087,N_3344);
nand U3502 (N_3502,N_3131,N_3215);
and U3503 (N_3503,N_3420,N_3213);
nand U3504 (N_3504,N_3308,N_3440);
or U3505 (N_3505,N_3177,N_3080);
and U3506 (N_3506,N_3313,N_3153);
or U3507 (N_3507,N_3179,N_3126);
and U3508 (N_3508,N_3012,N_3424);
or U3509 (N_3509,N_3415,N_3419);
or U3510 (N_3510,N_3296,N_3475);
and U3511 (N_3511,N_3387,N_3411);
and U3512 (N_3512,N_3007,N_3101);
nor U3513 (N_3513,N_3228,N_3060);
and U3514 (N_3514,N_3452,N_3459);
nand U3515 (N_3515,N_3326,N_3188);
nor U3516 (N_3516,N_3493,N_3453);
and U3517 (N_3517,N_3107,N_3255);
nand U3518 (N_3518,N_3043,N_3373);
nand U3519 (N_3519,N_3046,N_3463);
nand U3520 (N_3520,N_3240,N_3067);
or U3521 (N_3521,N_3383,N_3031);
nand U3522 (N_3522,N_3049,N_3465);
nand U3523 (N_3523,N_3464,N_3477);
nand U3524 (N_3524,N_3246,N_3166);
or U3525 (N_3525,N_3321,N_3317);
or U3526 (N_3526,N_3156,N_3004);
nor U3527 (N_3527,N_3431,N_3462);
or U3528 (N_3528,N_3430,N_3360);
or U3529 (N_3529,N_3123,N_3348);
or U3530 (N_3530,N_3115,N_3081);
nor U3531 (N_3531,N_3097,N_3476);
and U3532 (N_3532,N_3402,N_3030);
nor U3533 (N_3533,N_3122,N_3342);
and U3534 (N_3534,N_3171,N_3155);
or U3535 (N_3535,N_3318,N_3418);
or U3536 (N_3536,N_3445,N_3434);
and U3537 (N_3537,N_3357,N_3479);
or U3538 (N_3538,N_3409,N_3303);
nor U3539 (N_3539,N_3039,N_3191);
nor U3540 (N_3540,N_3371,N_3273);
xor U3541 (N_3541,N_3154,N_3334);
nor U3542 (N_3542,N_3422,N_3110);
and U3543 (N_3543,N_3397,N_3490);
nor U3544 (N_3544,N_3149,N_3243);
and U3545 (N_3545,N_3234,N_3429);
nor U3546 (N_3546,N_3141,N_3088);
or U3547 (N_3547,N_3205,N_3203);
nand U3548 (N_3548,N_3437,N_3054);
or U3549 (N_3549,N_3251,N_3162);
nor U3550 (N_3550,N_3204,N_3066);
and U3551 (N_3551,N_3372,N_3070);
or U3552 (N_3552,N_3382,N_3005);
and U3553 (N_3553,N_3061,N_3354);
nor U3554 (N_3554,N_3036,N_3289);
nor U3555 (N_3555,N_3374,N_3423);
nand U3556 (N_3556,N_3394,N_3366);
nor U3557 (N_3557,N_3349,N_3237);
nand U3558 (N_3558,N_3355,N_3198);
or U3559 (N_3559,N_3019,N_3444);
nand U3560 (N_3560,N_3403,N_3167);
nor U3561 (N_3561,N_3169,N_3062);
nand U3562 (N_3562,N_3449,N_3158);
nor U3563 (N_3563,N_3033,N_3180);
or U3564 (N_3564,N_3274,N_3053);
and U3565 (N_3565,N_3024,N_3145);
nand U3566 (N_3566,N_3211,N_3146);
nor U3567 (N_3567,N_3231,N_3266);
or U3568 (N_3568,N_3186,N_3000);
and U3569 (N_3569,N_3302,N_3257);
nor U3570 (N_3570,N_3219,N_3077);
nor U3571 (N_3571,N_3172,N_3176);
nor U3572 (N_3572,N_3425,N_3079);
and U3573 (N_3573,N_3329,N_3460);
nand U3574 (N_3574,N_3144,N_3207);
nand U3575 (N_3575,N_3233,N_3224);
nand U3576 (N_3576,N_3104,N_3286);
or U3577 (N_3577,N_3168,N_3014);
nor U3578 (N_3578,N_3450,N_3405);
nand U3579 (N_3579,N_3142,N_3347);
nor U3580 (N_3580,N_3029,N_3263);
or U3581 (N_3581,N_3291,N_3482);
or U3582 (N_3582,N_3069,N_3100);
nor U3583 (N_3583,N_3353,N_3268);
nand U3584 (N_3584,N_3035,N_3305);
nand U3585 (N_3585,N_3106,N_3456);
nand U3586 (N_3586,N_3293,N_3252);
nor U3587 (N_3587,N_3116,N_3244);
nand U3588 (N_3588,N_3071,N_3178);
nor U3589 (N_3589,N_3442,N_3269);
and U3590 (N_3590,N_3316,N_3309);
or U3591 (N_3591,N_3471,N_3025);
xnor U3592 (N_3592,N_3367,N_3328);
nor U3593 (N_3593,N_3307,N_3271);
nand U3594 (N_3594,N_3287,N_3421);
or U3595 (N_3595,N_3325,N_3193);
and U3596 (N_3596,N_3103,N_3132);
nor U3597 (N_3597,N_3018,N_3384);
xor U3598 (N_3598,N_3454,N_3136);
and U3599 (N_3599,N_3413,N_3406);
and U3600 (N_3600,N_3378,N_3451);
nor U3601 (N_3601,N_3323,N_3338);
or U3602 (N_3602,N_3059,N_3466);
nand U3603 (N_3603,N_3276,N_3285);
or U3604 (N_3604,N_3135,N_3042);
nor U3605 (N_3605,N_3130,N_3022);
nand U3606 (N_3606,N_3094,N_3361);
or U3607 (N_3607,N_3073,N_3074);
nand U3608 (N_3608,N_3414,N_3364);
nand U3609 (N_3609,N_3143,N_3426);
nor U3610 (N_3610,N_3469,N_3212);
or U3611 (N_3611,N_3262,N_3008);
or U3612 (N_3612,N_3174,N_3381);
and U3613 (N_3613,N_3390,N_3259);
xnor U3614 (N_3614,N_3428,N_3256);
and U3615 (N_3615,N_3298,N_3474);
or U3616 (N_3616,N_3229,N_3391);
and U3617 (N_3617,N_3301,N_3404);
nand U3618 (N_3618,N_3056,N_3194);
or U3619 (N_3619,N_3461,N_3249);
or U3620 (N_3620,N_3222,N_3206);
nand U3621 (N_3621,N_3187,N_3435);
nand U3622 (N_3622,N_3486,N_3150);
or U3623 (N_3623,N_3218,N_3330);
nor U3624 (N_3624,N_3236,N_3032);
and U3625 (N_3625,N_3408,N_3284);
nor U3626 (N_3626,N_3282,N_3047);
or U3627 (N_3627,N_3072,N_3358);
or U3628 (N_3628,N_3300,N_3001);
nor U3629 (N_3629,N_3337,N_3091);
nand U3630 (N_3630,N_3368,N_3133);
nor U3631 (N_3631,N_3125,N_3346);
nor U3632 (N_3632,N_3470,N_3128);
or U3633 (N_3633,N_3161,N_3199);
nor U3634 (N_3634,N_3108,N_3105);
nor U3635 (N_3635,N_3084,N_3196);
nand U3636 (N_3636,N_3173,N_3340);
nor U3637 (N_3637,N_3028,N_3417);
nor U3638 (N_3638,N_3260,N_3495);
nand U3639 (N_3639,N_3458,N_3253);
and U3640 (N_3640,N_3138,N_3075);
and U3641 (N_3641,N_3245,N_3189);
or U3642 (N_3642,N_3157,N_3432);
or U3643 (N_3643,N_3235,N_3279);
nor U3644 (N_3644,N_3034,N_3443);
or U3645 (N_3645,N_3485,N_3350);
and U3646 (N_3646,N_3139,N_3151);
or U3647 (N_3647,N_3226,N_3214);
nor U3648 (N_3648,N_3264,N_3009);
nor U3649 (N_3649,N_3312,N_3006);
nand U3650 (N_3650,N_3011,N_3113);
nand U3651 (N_3651,N_3379,N_3090);
nor U3652 (N_3652,N_3190,N_3159);
nor U3653 (N_3653,N_3002,N_3208);
or U3654 (N_3654,N_3248,N_3119);
nor U3655 (N_3655,N_3481,N_3345);
nand U3656 (N_3656,N_3057,N_3064);
nand U3657 (N_3657,N_3015,N_3339);
or U3658 (N_3658,N_3221,N_3448);
nor U3659 (N_3659,N_3480,N_3356);
nor U3660 (N_3660,N_3265,N_3488);
or U3661 (N_3661,N_3102,N_3147);
or U3662 (N_3662,N_3068,N_3010);
nor U3663 (N_3663,N_3095,N_3467);
nand U3664 (N_3664,N_3395,N_3225);
nand U3665 (N_3665,N_3182,N_3398);
and U3666 (N_3666,N_3017,N_3164);
nor U3667 (N_3667,N_3333,N_3241);
nand U3668 (N_3668,N_3170,N_3376);
nand U3669 (N_3669,N_3306,N_3270);
nand U3670 (N_3670,N_3331,N_3399);
and U3671 (N_3671,N_3468,N_3148);
and U3672 (N_3672,N_3195,N_3044);
and U3673 (N_3673,N_3436,N_3254);
nand U3674 (N_3674,N_3280,N_3290);
nand U3675 (N_3675,N_3393,N_3239);
nand U3676 (N_3676,N_3386,N_3496);
nor U3677 (N_3677,N_3063,N_3335);
or U3678 (N_3678,N_3160,N_3117);
nor U3679 (N_3679,N_3341,N_3457);
nand U3680 (N_3680,N_3183,N_3048);
nor U3681 (N_3681,N_3499,N_3489);
and U3682 (N_3682,N_3278,N_3114);
nor U3683 (N_3683,N_3050,N_3086);
nor U3684 (N_3684,N_3013,N_3016);
and U3685 (N_3685,N_3314,N_3129);
and U3686 (N_3686,N_3497,N_3238);
nor U3687 (N_3687,N_3416,N_3375);
nor U3688 (N_3688,N_3400,N_3439);
or U3689 (N_3689,N_3491,N_3359);
nand U3690 (N_3690,N_3343,N_3118);
or U3691 (N_3691,N_3277,N_3027);
and U3692 (N_3692,N_3082,N_3227);
nor U3693 (N_3693,N_3315,N_3065);
nor U3694 (N_3694,N_3380,N_3076);
and U3695 (N_3695,N_3472,N_3021);
or U3696 (N_3696,N_3242,N_3362);
nor U3697 (N_3697,N_3003,N_3447);
or U3698 (N_3698,N_3370,N_3197);
nor U3699 (N_3699,N_3051,N_3336);
or U3700 (N_3700,N_3365,N_3281);
and U3701 (N_3701,N_3299,N_3089);
and U3702 (N_3702,N_3327,N_3217);
or U3703 (N_3703,N_3210,N_3184);
or U3704 (N_3704,N_3052,N_3163);
nand U3705 (N_3705,N_3137,N_3275);
and U3706 (N_3706,N_3446,N_3322);
nand U3707 (N_3707,N_3192,N_3473);
and U3708 (N_3708,N_3363,N_3045);
xnor U3709 (N_3709,N_3433,N_3220);
nand U3710 (N_3710,N_3258,N_3216);
or U3711 (N_3711,N_3484,N_3093);
nor U3712 (N_3712,N_3223,N_3038);
and U3713 (N_3713,N_3392,N_3085);
nand U3714 (N_3714,N_3037,N_3020);
or U3715 (N_3715,N_3202,N_3295);
and U3716 (N_3716,N_3388,N_3055);
and U3717 (N_3717,N_3247,N_3401);
nand U3718 (N_3718,N_3412,N_3492);
and U3719 (N_3719,N_3483,N_3283);
nor U3720 (N_3720,N_3478,N_3152);
nand U3721 (N_3721,N_3441,N_3272);
nor U3722 (N_3722,N_3185,N_3427);
and U3723 (N_3723,N_3209,N_3111);
nand U3724 (N_3724,N_3494,N_3438);
or U3725 (N_3725,N_3140,N_3134);
and U3726 (N_3726,N_3311,N_3083);
nand U3727 (N_3727,N_3099,N_3096);
and U3728 (N_3728,N_3267,N_3040);
nor U3729 (N_3729,N_3181,N_3026);
nand U3730 (N_3730,N_3250,N_3304);
and U3731 (N_3731,N_3078,N_3396);
or U3732 (N_3732,N_3023,N_3165);
nor U3733 (N_3733,N_3041,N_3324);
or U3734 (N_3734,N_3407,N_3121);
and U3735 (N_3735,N_3261,N_3369);
and U3736 (N_3736,N_3127,N_3230);
nor U3737 (N_3737,N_3351,N_3092);
or U3738 (N_3738,N_3332,N_3410);
nor U3739 (N_3739,N_3112,N_3294);
nor U3740 (N_3740,N_3200,N_3297);
nand U3741 (N_3741,N_3320,N_3292);
nand U3742 (N_3742,N_3455,N_3498);
nand U3743 (N_3743,N_3288,N_3377);
and U3744 (N_3744,N_3310,N_3385);
nor U3745 (N_3745,N_3319,N_3175);
nand U3746 (N_3746,N_3201,N_3120);
nand U3747 (N_3747,N_3109,N_3487);
nor U3748 (N_3748,N_3124,N_3389);
nor U3749 (N_3749,N_3058,N_3352);
and U3750 (N_3750,N_3412,N_3167);
nor U3751 (N_3751,N_3304,N_3177);
and U3752 (N_3752,N_3493,N_3469);
nor U3753 (N_3753,N_3176,N_3254);
and U3754 (N_3754,N_3231,N_3431);
nor U3755 (N_3755,N_3412,N_3441);
nor U3756 (N_3756,N_3427,N_3259);
or U3757 (N_3757,N_3381,N_3344);
or U3758 (N_3758,N_3354,N_3486);
and U3759 (N_3759,N_3010,N_3329);
nor U3760 (N_3760,N_3340,N_3077);
and U3761 (N_3761,N_3447,N_3442);
and U3762 (N_3762,N_3059,N_3002);
nor U3763 (N_3763,N_3190,N_3021);
or U3764 (N_3764,N_3394,N_3390);
or U3765 (N_3765,N_3339,N_3012);
and U3766 (N_3766,N_3121,N_3492);
and U3767 (N_3767,N_3318,N_3191);
xor U3768 (N_3768,N_3099,N_3294);
and U3769 (N_3769,N_3492,N_3060);
nor U3770 (N_3770,N_3321,N_3294);
nand U3771 (N_3771,N_3292,N_3431);
or U3772 (N_3772,N_3215,N_3012);
nand U3773 (N_3773,N_3436,N_3219);
nand U3774 (N_3774,N_3325,N_3056);
nand U3775 (N_3775,N_3018,N_3383);
and U3776 (N_3776,N_3484,N_3277);
nor U3777 (N_3777,N_3289,N_3056);
and U3778 (N_3778,N_3347,N_3053);
or U3779 (N_3779,N_3282,N_3126);
or U3780 (N_3780,N_3444,N_3146);
nand U3781 (N_3781,N_3470,N_3233);
and U3782 (N_3782,N_3033,N_3426);
nand U3783 (N_3783,N_3122,N_3023);
nand U3784 (N_3784,N_3162,N_3311);
nand U3785 (N_3785,N_3370,N_3200);
and U3786 (N_3786,N_3299,N_3329);
and U3787 (N_3787,N_3171,N_3249);
nand U3788 (N_3788,N_3397,N_3233);
or U3789 (N_3789,N_3230,N_3066);
nor U3790 (N_3790,N_3393,N_3328);
nor U3791 (N_3791,N_3494,N_3425);
and U3792 (N_3792,N_3413,N_3212);
nor U3793 (N_3793,N_3046,N_3406);
nor U3794 (N_3794,N_3346,N_3434);
nand U3795 (N_3795,N_3216,N_3397);
and U3796 (N_3796,N_3305,N_3456);
nor U3797 (N_3797,N_3088,N_3490);
or U3798 (N_3798,N_3441,N_3415);
xnor U3799 (N_3799,N_3170,N_3115);
nand U3800 (N_3800,N_3035,N_3242);
nand U3801 (N_3801,N_3158,N_3309);
nand U3802 (N_3802,N_3268,N_3139);
and U3803 (N_3803,N_3070,N_3014);
or U3804 (N_3804,N_3273,N_3078);
nand U3805 (N_3805,N_3115,N_3436);
nor U3806 (N_3806,N_3444,N_3044);
or U3807 (N_3807,N_3243,N_3124);
or U3808 (N_3808,N_3312,N_3345);
nor U3809 (N_3809,N_3427,N_3174);
nor U3810 (N_3810,N_3095,N_3269);
or U3811 (N_3811,N_3298,N_3429);
nor U3812 (N_3812,N_3096,N_3334);
or U3813 (N_3813,N_3485,N_3056);
and U3814 (N_3814,N_3064,N_3229);
nand U3815 (N_3815,N_3073,N_3222);
or U3816 (N_3816,N_3332,N_3377);
or U3817 (N_3817,N_3136,N_3278);
or U3818 (N_3818,N_3321,N_3359);
and U3819 (N_3819,N_3147,N_3008);
nand U3820 (N_3820,N_3091,N_3219);
or U3821 (N_3821,N_3200,N_3418);
and U3822 (N_3822,N_3460,N_3492);
nand U3823 (N_3823,N_3304,N_3470);
and U3824 (N_3824,N_3264,N_3439);
or U3825 (N_3825,N_3000,N_3130);
nand U3826 (N_3826,N_3118,N_3116);
nor U3827 (N_3827,N_3190,N_3379);
nor U3828 (N_3828,N_3414,N_3343);
and U3829 (N_3829,N_3357,N_3369);
nor U3830 (N_3830,N_3443,N_3342);
nor U3831 (N_3831,N_3036,N_3098);
nand U3832 (N_3832,N_3441,N_3245);
nor U3833 (N_3833,N_3071,N_3000);
nand U3834 (N_3834,N_3215,N_3458);
or U3835 (N_3835,N_3395,N_3076);
or U3836 (N_3836,N_3087,N_3115);
and U3837 (N_3837,N_3282,N_3453);
nor U3838 (N_3838,N_3457,N_3198);
nor U3839 (N_3839,N_3015,N_3186);
or U3840 (N_3840,N_3053,N_3182);
nor U3841 (N_3841,N_3229,N_3442);
nor U3842 (N_3842,N_3113,N_3170);
nand U3843 (N_3843,N_3252,N_3108);
xor U3844 (N_3844,N_3006,N_3109);
and U3845 (N_3845,N_3160,N_3312);
nor U3846 (N_3846,N_3368,N_3326);
and U3847 (N_3847,N_3195,N_3190);
or U3848 (N_3848,N_3071,N_3408);
and U3849 (N_3849,N_3140,N_3332);
and U3850 (N_3850,N_3125,N_3390);
and U3851 (N_3851,N_3198,N_3430);
or U3852 (N_3852,N_3373,N_3070);
nor U3853 (N_3853,N_3274,N_3055);
xor U3854 (N_3854,N_3230,N_3045);
and U3855 (N_3855,N_3357,N_3230);
and U3856 (N_3856,N_3213,N_3012);
nor U3857 (N_3857,N_3046,N_3426);
or U3858 (N_3858,N_3407,N_3199);
nand U3859 (N_3859,N_3447,N_3486);
nand U3860 (N_3860,N_3421,N_3234);
nor U3861 (N_3861,N_3040,N_3379);
and U3862 (N_3862,N_3092,N_3235);
nor U3863 (N_3863,N_3264,N_3416);
and U3864 (N_3864,N_3375,N_3028);
and U3865 (N_3865,N_3079,N_3227);
nor U3866 (N_3866,N_3227,N_3365);
and U3867 (N_3867,N_3043,N_3484);
nor U3868 (N_3868,N_3151,N_3327);
or U3869 (N_3869,N_3076,N_3259);
or U3870 (N_3870,N_3170,N_3274);
nand U3871 (N_3871,N_3053,N_3355);
nor U3872 (N_3872,N_3133,N_3285);
nor U3873 (N_3873,N_3409,N_3302);
nand U3874 (N_3874,N_3068,N_3027);
and U3875 (N_3875,N_3387,N_3095);
or U3876 (N_3876,N_3424,N_3079);
nand U3877 (N_3877,N_3193,N_3072);
or U3878 (N_3878,N_3215,N_3157);
or U3879 (N_3879,N_3198,N_3129);
and U3880 (N_3880,N_3261,N_3327);
and U3881 (N_3881,N_3033,N_3093);
or U3882 (N_3882,N_3363,N_3364);
and U3883 (N_3883,N_3019,N_3446);
nor U3884 (N_3884,N_3333,N_3096);
nor U3885 (N_3885,N_3279,N_3001);
and U3886 (N_3886,N_3012,N_3017);
nor U3887 (N_3887,N_3305,N_3118);
nor U3888 (N_3888,N_3328,N_3032);
nor U3889 (N_3889,N_3305,N_3377);
nand U3890 (N_3890,N_3385,N_3399);
and U3891 (N_3891,N_3095,N_3209);
nand U3892 (N_3892,N_3210,N_3467);
nand U3893 (N_3893,N_3127,N_3342);
nor U3894 (N_3894,N_3012,N_3071);
nor U3895 (N_3895,N_3165,N_3262);
nand U3896 (N_3896,N_3105,N_3211);
or U3897 (N_3897,N_3141,N_3161);
nand U3898 (N_3898,N_3168,N_3303);
nor U3899 (N_3899,N_3319,N_3259);
or U3900 (N_3900,N_3179,N_3292);
nor U3901 (N_3901,N_3430,N_3433);
or U3902 (N_3902,N_3456,N_3083);
or U3903 (N_3903,N_3139,N_3348);
nand U3904 (N_3904,N_3034,N_3487);
nor U3905 (N_3905,N_3147,N_3171);
or U3906 (N_3906,N_3389,N_3459);
and U3907 (N_3907,N_3421,N_3369);
and U3908 (N_3908,N_3446,N_3121);
and U3909 (N_3909,N_3085,N_3314);
nand U3910 (N_3910,N_3396,N_3011);
nand U3911 (N_3911,N_3290,N_3106);
nand U3912 (N_3912,N_3322,N_3281);
nand U3913 (N_3913,N_3255,N_3175);
or U3914 (N_3914,N_3119,N_3366);
nand U3915 (N_3915,N_3030,N_3005);
nand U3916 (N_3916,N_3495,N_3437);
nor U3917 (N_3917,N_3062,N_3449);
or U3918 (N_3918,N_3120,N_3192);
nor U3919 (N_3919,N_3344,N_3050);
or U3920 (N_3920,N_3012,N_3434);
and U3921 (N_3921,N_3083,N_3152);
nand U3922 (N_3922,N_3088,N_3498);
nand U3923 (N_3923,N_3363,N_3039);
nand U3924 (N_3924,N_3046,N_3483);
or U3925 (N_3925,N_3374,N_3368);
nor U3926 (N_3926,N_3031,N_3246);
or U3927 (N_3927,N_3366,N_3345);
nand U3928 (N_3928,N_3437,N_3163);
nor U3929 (N_3929,N_3385,N_3445);
nand U3930 (N_3930,N_3007,N_3384);
nor U3931 (N_3931,N_3039,N_3210);
nor U3932 (N_3932,N_3165,N_3286);
or U3933 (N_3933,N_3169,N_3095);
nand U3934 (N_3934,N_3257,N_3167);
and U3935 (N_3935,N_3123,N_3304);
or U3936 (N_3936,N_3273,N_3438);
nand U3937 (N_3937,N_3139,N_3454);
and U3938 (N_3938,N_3248,N_3358);
nor U3939 (N_3939,N_3021,N_3199);
and U3940 (N_3940,N_3473,N_3184);
nor U3941 (N_3941,N_3230,N_3210);
or U3942 (N_3942,N_3480,N_3069);
and U3943 (N_3943,N_3078,N_3055);
nor U3944 (N_3944,N_3032,N_3424);
nand U3945 (N_3945,N_3106,N_3244);
and U3946 (N_3946,N_3121,N_3481);
or U3947 (N_3947,N_3193,N_3256);
or U3948 (N_3948,N_3479,N_3245);
nor U3949 (N_3949,N_3130,N_3017);
nand U3950 (N_3950,N_3088,N_3022);
or U3951 (N_3951,N_3254,N_3035);
and U3952 (N_3952,N_3359,N_3202);
or U3953 (N_3953,N_3035,N_3421);
or U3954 (N_3954,N_3107,N_3446);
and U3955 (N_3955,N_3353,N_3297);
nor U3956 (N_3956,N_3350,N_3373);
and U3957 (N_3957,N_3104,N_3248);
or U3958 (N_3958,N_3166,N_3032);
and U3959 (N_3959,N_3277,N_3111);
or U3960 (N_3960,N_3212,N_3229);
or U3961 (N_3961,N_3032,N_3036);
nand U3962 (N_3962,N_3280,N_3070);
nand U3963 (N_3963,N_3480,N_3047);
and U3964 (N_3964,N_3109,N_3461);
or U3965 (N_3965,N_3057,N_3315);
or U3966 (N_3966,N_3139,N_3228);
or U3967 (N_3967,N_3196,N_3165);
nand U3968 (N_3968,N_3294,N_3477);
and U3969 (N_3969,N_3182,N_3386);
or U3970 (N_3970,N_3008,N_3220);
nor U3971 (N_3971,N_3400,N_3477);
and U3972 (N_3972,N_3469,N_3057);
nor U3973 (N_3973,N_3451,N_3141);
or U3974 (N_3974,N_3422,N_3155);
and U3975 (N_3975,N_3159,N_3222);
and U3976 (N_3976,N_3307,N_3483);
nand U3977 (N_3977,N_3001,N_3011);
nor U3978 (N_3978,N_3139,N_3430);
xor U3979 (N_3979,N_3400,N_3200);
nor U3980 (N_3980,N_3351,N_3341);
nand U3981 (N_3981,N_3288,N_3362);
nor U3982 (N_3982,N_3041,N_3345);
nand U3983 (N_3983,N_3243,N_3341);
or U3984 (N_3984,N_3216,N_3175);
nor U3985 (N_3985,N_3484,N_3366);
nand U3986 (N_3986,N_3177,N_3429);
and U3987 (N_3987,N_3276,N_3116);
or U3988 (N_3988,N_3026,N_3257);
and U3989 (N_3989,N_3197,N_3376);
nor U3990 (N_3990,N_3371,N_3083);
or U3991 (N_3991,N_3304,N_3074);
nand U3992 (N_3992,N_3124,N_3261);
nor U3993 (N_3993,N_3415,N_3062);
xor U3994 (N_3994,N_3230,N_3262);
and U3995 (N_3995,N_3130,N_3276);
nand U3996 (N_3996,N_3394,N_3078);
or U3997 (N_3997,N_3339,N_3095);
and U3998 (N_3998,N_3063,N_3486);
or U3999 (N_3999,N_3274,N_3305);
and U4000 (N_4000,N_3835,N_3995);
or U4001 (N_4001,N_3556,N_3551);
and U4002 (N_4002,N_3571,N_3758);
nand U4003 (N_4003,N_3520,N_3603);
or U4004 (N_4004,N_3627,N_3679);
and U4005 (N_4005,N_3595,N_3975);
nor U4006 (N_4006,N_3817,N_3553);
and U4007 (N_4007,N_3977,N_3508);
and U4008 (N_4008,N_3938,N_3747);
nand U4009 (N_4009,N_3545,N_3771);
or U4010 (N_4010,N_3648,N_3843);
and U4011 (N_4011,N_3557,N_3684);
or U4012 (N_4012,N_3926,N_3916);
or U4013 (N_4013,N_3583,N_3905);
nor U4014 (N_4014,N_3988,N_3879);
or U4015 (N_4015,N_3574,N_3895);
or U4016 (N_4016,N_3548,N_3955);
and U4017 (N_4017,N_3705,N_3527);
and U4018 (N_4018,N_3822,N_3830);
or U4019 (N_4019,N_3718,N_3581);
or U4020 (N_4020,N_3927,N_3788);
and U4021 (N_4021,N_3911,N_3946);
nor U4022 (N_4022,N_3956,N_3516);
nand U4023 (N_4023,N_3555,N_3722);
nand U4024 (N_4024,N_3763,N_3731);
nand U4025 (N_4025,N_3728,N_3529);
nand U4026 (N_4026,N_3781,N_3875);
and U4027 (N_4027,N_3866,N_3960);
and U4028 (N_4028,N_3588,N_3623);
nor U4029 (N_4029,N_3864,N_3576);
and U4030 (N_4030,N_3669,N_3855);
or U4031 (N_4031,N_3602,N_3900);
xnor U4032 (N_4032,N_3882,N_3532);
or U4033 (N_4033,N_3994,N_3767);
or U4034 (N_4034,N_3510,N_3608);
nor U4035 (N_4035,N_3974,N_3564);
nor U4036 (N_4036,N_3859,N_3600);
or U4037 (N_4037,N_3686,N_3785);
or U4038 (N_4038,N_3656,N_3642);
nand U4039 (N_4039,N_3552,N_3775);
nor U4040 (N_4040,N_3805,N_3562);
or U4041 (N_4041,N_3820,N_3888);
or U4042 (N_4042,N_3971,N_3650);
or U4043 (N_4043,N_3521,N_3784);
and U4044 (N_4044,N_3861,N_3518);
nor U4045 (N_4045,N_3856,N_3726);
and U4046 (N_4046,N_3837,N_3515);
nand U4047 (N_4047,N_3745,N_3725);
nor U4048 (N_4048,N_3565,N_3634);
nand U4049 (N_4049,N_3870,N_3885);
or U4050 (N_4050,N_3857,N_3958);
nor U4051 (N_4051,N_3964,N_3982);
or U4052 (N_4052,N_3867,N_3702);
nor U4053 (N_4053,N_3723,N_3724);
and U4054 (N_4054,N_3647,N_3945);
or U4055 (N_4055,N_3873,N_3792);
or U4056 (N_4056,N_3890,N_3904);
and U4057 (N_4057,N_3983,N_3672);
and U4058 (N_4058,N_3706,N_3751);
xor U4059 (N_4059,N_3733,N_3644);
and U4060 (N_4060,N_3554,N_3930);
and U4061 (N_4061,N_3736,N_3687);
nand U4062 (N_4062,N_3948,N_3746);
or U4063 (N_4063,N_3625,N_3940);
nand U4064 (N_4064,N_3766,N_3711);
nand U4065 (N_4065,N_3871,N_3538);
nand U4066 (N_4066,N_3793,N_3807);
nand U4067 (N_4067,N_3893,N_3735);
nand U4068 (N_4068,N_3840,N_3512);
nand U4069 (N_4069,N_3652,N_3847);
or U4070 (N_4070,N_3714,N_3522);
nand U4071 (N_4071,N_3743,N_3922);
or U4072 (N_4072,N_3637,N_3773);
nor U4073 (N_4073,N_3610,N_3523);
nor U4074 (N_4074,N_3984,N_3591);
or U4075 (N_4075,N_3883,N_3531);
and U4076 (N_4076,N_3823,N_3989);
nor U4077 (N_4077,N_3750,N_3813);
nor U4078 (N_4078,N_3617,N_3619);
nand U4079 (N_4079,N_3919,N_3566);
and U4080 (N_4080,N_3791,N_3730);
nand U4081 (N_4081,N_3663,N_3596);
and U4082 (N_4082,N_3671,N_3740);
nor U4083 (N_4083,N_3549,N_3782);
nand U4084 (N_4084,N_3721,N_3690);
nand U4085 (N_4085,N_3547,N_3661);
nand U4086 (N_4086,N_3601,N_3657);
nand U4087 (N_4087,N_3914,N_3836);
nor U4088 (N_4088,N_3673,N_3613);
nor U4089 (N_4089,N_3821,N_3993);
nor U4090 (N_4090,N_3704,N_3972);
or U4091 (N_4091,N_3812,N_3636);
or U4092 (N_4092,N_3951,N_3563);
or U4093 (N_4093,N_3825,N_3910);
nor U4094 (N_4094,N_3752,N_3999);
or U4095 (N_4095,N_3528,N_3645);
and U4096 (N_4096,N_3839,N_3921);
xnor U4097 (N_4097,N_3525,N_3710);
or U4098 (N_4098,N_3701,N_3933);
nor U4099 (N_4099,N_3901,N_3831);
nor U4100 (N_4100,N_3632,N_3963);
nor U4101 (N_4101,N_3973,N_3621);
xor U4102 (N_4102,N_3778,N_3950);
or U4103 (N_4103,N_3559,N_3981);
or U4104 (N_4104,N_3729,N_3590);
and U4105 (N_4105,N_3500,N_3903);
or U4106 (N_4106,N_3783,N_3920);
or U4107 (N_4107,N_3824,N_3978);
or U4108 (N_4108,N_3662,N_3717);
and U4109 (N_4109,N_3676,N_3809);
or U4110 (N_4110,N_3534,N_3509);
or U4111 (N_4111,N_3524,N_3540);
nor U4112 (N_4112,N_3877,N_3970);
nand U4113 (N_4113,N_3908,N_3818);
and U4114 (N_4114,N_3991,N_3694);
nor U4115 (N_4115,N_3570,N_3641);
xnor U4116 (N_4116,N_3878,N_3703);
nand U4117 (N_4117,N_3678,N_3691);
nor U4118 (N_4118,N_3614,N_3802);
or U4119 (N_4119,N_3707,N_3804);
and U4120 (N_4120,N_3742,N_3929);
nor U4121 (N_4121,N_3585,N_3827);
or U4122 (N_4122,N_3913,N_3841);
nor U4123 (N_4123,N_3819,N_3779);
nand U4124 (N_4124,N_3838,N_3580);
or U4125 (N_4125,N_3768,N_3851);
nor U4126 (N_4126,N_3698,N_3902);
nor U4127 (N_4127,N_3936,N_3667);
and U4128 (N_4128,N_3889,N_3789);
and U4129 (N_4129,N_3953,N_3598);
nor U4130 (N_4130,N_3616,N_3862);
or U4131 (N_4131,N_3561,N_3876);
or U4132 (N_4132,N_3689,N_3874);
and U4133 (N_4133,N_3957,N_3535);
or U4134 (N_4134,N_3530,N_3537);
or U4135 (N_4135,N_3573,N_3814);
or U4136 (N_4136,N_3918,N_3987);
and U4137 (N_4137,N_3578,N_3850);
and U4138 (N_4138,N_3898,N_3937);
and U4139 (N_4139,N_3624,N_3697);
and U4140 (N_4140,N_3786,N_3633);
nor U4141 (N_4141,N_3967,N_3593);
or U4142 (N_4142,N_3699,N_3604);
or U4143 (N_4143,N_3611,N_3849);
nand U4144 (N_4144,N_3666,N_3795);
and U4145 (N_4145,N_3780,N_3734);
nor U4146 (N_4146,N_3577,N_3536);
and U4147 (N_4147,N_3816,N_3806);
or U4148 (N_4148,N_3959,N_3749);
nand U4149 (N_4149,N_3759,N_3541);
and U4150 (N_4150,N_3845,N_3599);
and U4151 (N_4151,N_3715,N_3526);
nand U4152 (N_4152,N_3544,N_3865);
nand U4153 (N_4153,N_3727,N_3772);
nand U4154 (N_4154,N_3649,N_3976);
nand U4155 (N_4155,N_3719,N_3986);
nor U4156 (N_4156,N_3612,N_3700);
or U4157 (N_4157,N_3655,N_3801);
and U4158 (N_4158,N_3797,N_3777);
or U4159 (N_4159,N_3668,N_3880);
nor U4160 (N_4160,N_3560,N_3660);
nand U4161 (N_4161,N_3607,N_3584);
and U4162 (N_4162,N_3934,N_3646);
nand U4163 (N_4163,N_3844,N_3949);
nand U4164 (N_4164,N_3790,N_3635);
nor U4165 (N_4165,N_3692,N_3931);
nand U4166 (N_4166,N_3630,N_3980);
nand U4167 (N_4167,N_3770,N_3834);
nor U4168 (N_4168,N_3832,N_3799);
and U4169 (N_4169,N_3643,N_3869);
nand U4170 (N_4170,N_3764,N_3696);
and U4171 (N_4171,N_3962,N_3965);
nor U4172 (N_4172,N_3744,N_3558);
nor U4173 (N_4173,N_3606,N_3943);
or U4174 (N_4174,N_3757,N_3589);
nor U4175 (N_4175,N_3594,N_3969);
nand U4176 (N_4176,N_3952,N_3891);
or U4177 (N_4177,N_3979,N_3897);
nor U4178 (N_4178,N_3505,N_3543);
or U4179 (N_4179,N_3917,N_3848);
or U4180 (N_4180,N_3587,N_3815);
and U4181 (N_4181,N_3708,N_3659);
nor U4182 (N_4182,N_3892,N_3787);
nor U4183 (N_4183,N_3654,N_3996);
nand U4184 (N_4184,N_3681,N_3899);
and U4185 (N_4185,N_3896,N_3756);
or U4186 (N_4186,N_3502,N_3622);
nand U4187 (N_4187,N_3683,N_3693);
nor U4188 (N_4188,N_3658,N_3638);
nor U4189 (N_4189,N_3828,N_3761);
or U4190 (N_4190,N_3939,N_3688);
or U4191 (N_4191,N_3811,N_3829);
or U4192 (N_4192,N_3501,N_3852);
or U4193 (N_4193,N_3915,N_3738);
nand U4194 (N_4194,N_3968,N_3514);
nand U4195 (N_4195,N_3954,N_3695);
nor U4196 (N_4196,N_3924,N_3550);
or U4197 (N_4197,N_3629,N_3798);
nand U4198 (N_4198,N_3854,N_3932);
nand U4199 (N_4199,N_3928,N_3712);
nand U4200 (N_4200,N_3677,N_3941);
and U4201 (N_4201,N_3567,N_3572);
nand U4202 (N_4202,N_3796,N_3826);
nand U4203 (N_4203,N_3609,N_3620);
nand U4204 (N_4204,N_3539,N_3909);
nor U4205 (N_4205,N_3685,N_3626);
and U4206 (N_4206,N_3808,N_3716);
and U4207 (N_4207,N_3519,N_3513);
nor U4208 (N_4208,N_3713,N_3506);
or U4209 (N_4209,N_3769,N_3985);
nand U4210 (N_4210,N_3517,N_3762);
and U4211 (N_4211,N_3511,N_3753);
nor U4212 (N_4212,N_3615,N_3912);
nor U4213 (N_4213,N_3894,N_3853);
nand U4214 (N_4214,N_3794,N_3754);
nor U4215 (N_4215,N_3674,N_3906);
or U4216 (N_4216,N_3886,N_3992);
nand U4217 (N_4217,N_3868,N_3942);
nor U4218 (N_4218,N_3776,N_3582);
and U4219 (N_4219,N_3748,N_3833);
nor U4220 (N_4220,N_3680,N_3631);
nor U4221 (N_4221,N_3651,N_3507);
and U4222 (N_4222,N_3760,N_3884);
or U4223 (N_4223,N_3846,N_3503);
nor U4224 (N_4224,N_3504,N_3961);
nor U4225 (N_4225,N_3569,N_3739);
and U4226 (N_4226,N_3947,N_3575);
nand U4227 (N_4227,N_3966,N_3597);
or U4228 (N_4228,N_3737,N_3810);
and U4229 (N_4229,N_3670,N_3618);
or U4230 (N_4230,N_3665,N_3640);
nor U4231 (N_4231,N_3842,N_3732);
and U4232 (N_4232,N_3858,N_3800);
nand U4233 (N_4233,N_3586,N_3863);
or U4234 (N_4234,N_3881,N_3579);
nand U4235 (N_4235,N_3628,N_3925);
or U4236 (N_4236,N_3546,N_3682);
or U4237 (N_4237,N_3675,N_3923);
or U4238 (N_4238,N_3741,N_3533);
or U4239 (N_4239,N_3709,N_3664);
and U4240 (N_4240,N_3998,N_3997);
or U4241 (N_4241,N_3568,N_3872);
nor U4242 (N_4242,N_3653,N_3639);
or U4243 (N_4243,N_3605,N_3860);
nor U4244 (N_4244,N_3803,N_3592);
nor U4245 (N_4245,N_3944,N_3720);
or U4246 (N_4246,N_3990,N_3774);
xnor U4247 (N_4247,N_3755,N_3765);
or U4248 (N_4248,N_3542,N_3887);
nor U4249 (N_4249,N_3907,N_3935);
nor U4250 (N_4250,N_3673,N_3889);
nand U4251 (N_4251,N_3952,N_3583);
nand U4252 (N_4252,N_3810,N_3650);
nand U4253 (N_4253,N_3690,N_3551);
xnor U4254 (N_4254,N_3794,N_3711);
nand U4255 (N_4255,N_3581,N_3667);
and U4256 (N_4256,N_3688,N_3961);
or U4257 (N_4257,N_3530,N_3808);
nor U4258 (N_4258,N_3733,N_3983);
nor U4259 (N_4259,N_3726,N_3834);
nand U4260 (N_4260,N_3755,N_3648);
or U4261 (N_4261,N_3784,N_3794);
nor U4262 (N_4262,N_3653,N_3783);
xnor U4263 (N_4263,N_3772,N_3855);
or U4264 (N_4264,N_3980,N_3606);
and U4265 (N_4265,N_3714,N_3777);
nand U4266 (N_4266,N_3758,N_3563);
and U4267 (N_4267,N_3947,N_3691);
nor U4268 (N_4268,N_3993,N_3673);
or U4269 (N_4269,N_3686,N_3620);
nor U4270 (N_4270,N_3951,N_3510);
nor U4271 (N_4271,N_3614,N_3873);
and U4272 (N_4272,N_3922,N_3718);
nor U4273 (N_4273,N_3698,N_3792);
or U4274 (N_4274,N_3754,N_3576);
and U4275 (N_4275,N_3922,N_3684);
and U4276 (N_4276,N_3749,N_3912);
and U4277 (N_4277,N_3957,N_3959);
and U4278 (N_4278,N_3726,N_3737);
nand U4279 (N_4279,N_3609,N_3579);
or U4280 (N_4280,N_3795,N_3546);
or U4281 (N_4281,N_3700,N_3577);
nor U4282 (N_4282,N_3866,N_3877);
nor U4283 (N_4283,N_3856,N_3956);
nor U4284 (N_4284,N_3505,N_3896);
nor U4285 (N_4285,N_3530,N_3704);
nand U4286 (N_4286,N_3846,N_3762);
or U4287 (N_4287,N_3692,N_3646);
or U4288 (N_4288,N_3723,N_3510);
nor U4289 (N_4289,N_3959,N_3653);
nand U4290 (N_4290,N_3783,N_3925);
nand U4291 (N_4291,N_3748,N_3969);
or U4292 (N_4292,N_3848,N_3708);
nor U4293 (N_4293,N_3755,N_3818);
nor U4294 (N_4294,N_3611,N_3761);
nand U4295 (N_4295,N_3730,N_3591);
nand U4296 (N_4296,N_3828,N_3912);
and U4297 (N_4297,N_3674,N_3988);
or U4298 (N_4298,N_3736,N_3857);
nand U4299 (N_4299,N_3719,N_3924);
nand U4300 (N_4300,N_3547,N_3551);
and U4301 (N_4301,N_3581,N_3773);
or U4302 (N_4302,N_3871,N_3717);
nand U4303 (N_4303,N_3705,N_3964);
or U4304 (N_4304,N_3653,N_3641);
and U4305 (N_4305,N_3562,N_3855);
and U4306 (N_4306,N_3609,N_3582);
and U4307 (N_4307,N_3801,N_3803);
and U4308 (N_4308,N_3840,N_3594);
nor U4309 (N_4309,N_3744,N_3825);
xor U4310 (N_4310,N_3677,N_3533);
or U4311 (N_4311,N_3627,N_3843);
nand U4312 (N_4312,N_3704,N_3695);
nor U4313 (N_4313,N_3968,N_3726);
nand U4314 (N_4314,N_3658,N_3875);
nor U4315 (N_4315,N_3801,N_3513);
or U4316 (N_4316,N_3529,N_3917);
or U4317 (N_4317,N_3663,N_3634);
and U4318 (N_4318,N_3739,N_3501);
nor U4319 (N_4319,N_3964,N_3707);
and U4320 (N_4320,N_3649,N_3564);
nor U4321 (N_4321,N_3555,N_3590);
or U4322 (N_4322,N_3702,N_3861);
nor U4323 (N_4323,N_3580,N_3670);
or U4324 (N_4324,N_3783,N_3503);
or U4325 (N_4325,N_3650,N_3655);
or U4326 (N_4326,N_3991,N_3604);
nand U4327 (N_4327,N_3683,N_3794);
and U4328 (N_4328,N_3893,N_3921);
and U4329 (N_4329,N_3963,N_3696);
nor U4330 (N_4330,N_3958,N_3658);
or U4331 (N_4331,N_3843,N_3753);
nor U4332 (N_4332,N_3914,N_3641);
nand U4333 (N_4333,N_3564,N_3863);
or U4334 (N_4334,N_3706,N_3775);
and U4335 (N_4335,N_3639,N_3561);
nand U4336 (N_4336,N_3879,N_3551);
nor U4337 (N_4337,N_3712,N_3501);
nor U4338 (N_4338,N_3836,N_3624);
nor U4339 (N_4339,N_3712,N_3655);
and U4340 (N_4340,N_3655,N_3827);
and U4341 (N_4341,N_3884,N_3543);
nor U4342 (N_4342,N_3657,N_3832);
nand U4343 (N_4343,N_3916,N_3884);
or U4344 (N_4344,N_3592,N_3685);
nand U4345 (N_4345,N_3994,N_3815);
nand U4346 (N_4346,N_3588,N_3570);
or U4347 (N_4347,N_3740,N_3717);
nand U4348 (N_4348,N_3857,N_3780);
nand U4349 (N_4349,N_3825,N_3565);
nand U4350 (N_4350,N_3788,N_3819);
nor U4351 (N_4351,N_3569,N_3841);
nand U4352 (N_4352,N_3691,N_3577);
and U4353 (N_4353,N_3873,N_3933);
or U4354 (N_4354,N_3573,N_3603);
and U4355 (N_4355,N_3753,N_3778);
or U4356 (N_4356,N_3590,N_3843);
nand U4357 (N_4357,N_3662,N_3740);
nand U4358 (N_4358,N_3911,N_3783);
nand U4359 (N_4359,N_3883,N_3881);
nand U4360 (N_4360,N_3743,N_3993);
nor U4361 (N_4361,N_3725,N_3554);
and U4362 (N_4362,N_3881,N_3566);
nand U4363 (N_4363,N_3715,N_3702);
or U4364 (N_4364,N_3625,N_3595);
and U4365 (N_4365,N_3701,N_3581);
nand U4366 (N_4366,N_3873,N_3892);
and U4367 (N_4367,N_3934,N_3534);
nor U4368 (N_4368,N_3798,N_3646);
nand U4369 (N_4369,N_3615,N_3965);
or U4370 (N_4370,N_3887,N_3716);
and U4371 (N_4371,N_3636,N_3658);
nand U4372 (N_4372,N_3719,N_3763);
or U4373 (N_4373,N_3696,N_3721);
or U4374 (N_4374,N_3932,N_3830);
nand U4375 (N_4375,N_3778,N_3755);
or U4376 (N_4376,N_3584,N_3830);
or U4377 (N_4377,N_3659,N_3946);
and U4378 (N_4378,N_3776,N_3746);
nand U4379 (N_4379,N_3630,N_3657);
or U4380 (N_4380,N_3521,N_3752);
or U4381 (N_4381,N_3734,N_3789);
or U4382 (N_4382,N_3548,N_3901);
nand U4383 (N_4383,N_3529,N_3691);
or U4384 (N_4384,N_3565,N_3837);
nor U4385 (N_4385,N_3895,N_3776);
nor U4386 (N_4386,N_3567,N_3821);
or U4387 (N_4387,N_3679,N_3896);
or U4388 (N_4388,N_3521,N_3531);
nor U4389 (N_4389,N_3589,N_3771);
and U4390 (N_4390,N_3664,N_3541);
or U4391 (N_4391,N_3982,N_3684);
or U4392 (N_4392,N_3857,N_3542);
nor U4393 (N_4393,N_3698,N_3501);
nor U4394 (N_4394,N_3752,N_3737);
nor U4395 (N_4395,N_3546,N_3570);
or U4396 (N_4396,N_3831,N_3533);
and U4397 (N_4397,N_3838,N_3608);
nor U4398 (N_4398,N_3909,N_3530);
and U4399 (N_4399,N_3965,N_3913);
or U4400 (N_4400,N_3527,N_3891);
nand U4401 (N_4401,N_3988,N_3718);
and U4402 (N_4402,N_3839,N_3723);
nand U4403 (N_4403,N_3745,N_3917);
or U4404 (N_4404,N_3834,N_3941);
nand U4405 (N_4405,N_3942,N_3956);
and U4406 (N_4406,N_3645,N_3686);
or U4407 (N_4407,N_3523,N_3815);
and U4408 (N_4408,N_3930,N_3615);
or U4409 (N_4409,N_3846,N_3694);
and U4410 (N_4410,N_3720,N_3574);
nand U4411 (N_4411,N_3751,N_3853);
nor U4412 (N_4412,N_3731,N_3645);
nor U4413 (N_4413,N_3646,N_3576);
or U4414 (N_4414,N_3809,N_3929);
or U4415 (N_4415,N_3920,N_3548);
and U4416 (N_4416,N_3880,N_3720);
and U4417 (N_4417,N_3677,N_3936);
nor U4418 (N_4418,N_3993,N_3571);
nor U4419 (N_4419,N_3539,N_3753);
nor U4420 (N_4420,N_3885,N_3882);
nand U4421 (N_4421,N_3727,N_3853);
nor U4422 (N_4422,N_3905,N_3953);
and U4423 (N_4423,N_3864,N_3976);
or U4424 (N_4424,N_3995,N_3507);
nand U4425 (N_4425,N_3779,N_3964);
and U4426 (N_4426,N_3769,N_3538);
nor U4427 (N_4427,N_3961,N_3862);
or U4428 (N_4428,N_3626,N_3655);
xnor U4429 (N_4429,N_3537,N_3769);
nor U4430 (N_4430,N_3774,N_3786);
nor U4431 (N_4431,N_3501,N_3686);
or U4432 (N_4432,N_3886,N_3632);
or U4433 (N_4433,N_3791,N_3596);
and U4434 (N_4434,N_3504,N_3765);
or U4435 (N_4435,N_3547,N_3578);
nand U4436 (N_4436,N_3825,N_3660);
or U4437 (N_4437,N_3620,N_3737);
or U4438 (N_4438,N_3937,N_3729);
nor U4439 (N_4439,N_3698,N_3998);
nor U4440 (N_4440,N_3797,N_3819);
nand U4441 (N_4441,N_3788,N_3707);
and U4442 (N_4442,N_3509,N_3525);
or U4443 (N_4443,N_3994,N_3516);
nor U4444 (N_4444,N_3665,N_3557);
and U4445 (N_4445,N_3888,N_3525);
nor U4446 (N_4446,N_3559,N_3967);
and U4447 (N_4447,N_3938,N_3548);
or U4448 (N_4448,N_3582,N_3522);
or U4449 (N_4449,N_3750,N_3931);
nand U4450 (N_4450,N_3604,N_3688);
or U4451 (N_4451,N_3753,N_3836);
nand U4452 (N_4452,N_3585,N_3809);
and U4453 (N_4453,N_3607,N_3660);
nor U4454 (N_4454,N_3734,N_3791);
nand U4455 (N_4455,N_3874,N_3970);
and U4456 (N_4456,N_3748,N_3620);
nand U4457 (N_4457,N_3904,N_3732);
xor U4458 (N_4458,N_3622,N_3698);
nor U4459 (N_4459,N_3604,N_3795);
or U4460 (N_4460,N_3666,N_3712);
and U4461 (N_4461,N_3744,N_3989);
nor U4462 (N_4462,N_3851,N_3985);
and U4463 (N_4463,N_3708,N_3773);
or U4464 (N_4464,N_3580,N_3535);
nand U4465 (N_4465,N_3550,N_3709);
nor U4466 (N_4466,N_3913,N_3669);
and U4467 (N_4467,N_3628,N_3961);
nand U4468 (N_4468,N_3564,N_3995);
and U4469 (N_4469,N_3688,N_3937);
or U4470 (N_4470,N_3625,N_3598);
nand U4471 (N_4471,N_3945,N_3823);
or U4472 (N_4472,N_3833,N_3761);
nor U4473 (N_4473,N_3963,N_3508);
or U4474 (N_4474,N_3589,N_3801);
or U4475 (N_4475,N_3876,N_3989);
nor U4476 (N_4476,N_3659,N_3833);
nor U4477 (N_4477,N_3669,N_3691);
nor U4478 (N_4478,N_3909,N_3979);
nor U4479 (N_4479,N_3885,N_3817);
nand U4480 (N_4480,N_3853,N_3708);
nor U4481 (N_4481,N_3666,N_3585);
or U4482 (N_4482,N_3866,N_3722);
nor U4483 (N_4483,N_3846,N_3801);
or U4484 (N_4484,N_3722,N_3619);
nand U4485 (N_4485,N_3500,N_3604);
nand U4486 (N_4486,N_3843,N_3595);
nand U4487 (N_4487,N_3801,N_3509);
and U4488 (N_4488,N_3799,N_3877);
nand U4489 (N_4489,N_3745,N_3696);
nand U4490 (N_4490,N_3663,N_3883);
nand U4491 (N_4491,N_3526,N_3957);
and U4492 (N_4492,N_3551,N_3704);
nor U4493 (N_4493,N_3794,N_3500);
xor U4494 (N_4494,N_3920,N_3751);
nand U4495 (N_4495,N_3905,N_3840);
nor U4496 (N_4496,N_3728,N_3535);
nand U4497 (N_4497,N_3645,N_3625);
or U4498 (N_4498,N_3879,N_3546);
or U4499 (N_4499,N_3746,N_3749);
nand U4500 (N_4500,N_4428,N_4083);
nand U4501 (N_4501,N_4011,N_4365);
or U4502 (N_4502,N_4392,N_4035);
nand U4503 (N_4503,N_4148,N_4258);
nand U4504 (N_4504,N_4104,N_4355);
or U4505 (N_4505,N_4028,N_4447);
nand U4506 (N_4506,N_4055,N_4397);
and U4507 (N_4507,N_4107,N_4054);
and U4508 (N_4508,N_4477,N_4191);
and U4509 (N_4509,N_4364,N_4303);
nor U4510 (N_4510,N_4342,N_4015);
or U4511 (N_4511,N_4217,N_4131);
or U4512 (N_4512,N_4010,N_4346);
or U4513 (N_4513,N_4223,N_4067);
or U4514 (N_4514,N_4317,N_4375);
and U4515 (N_4515,N_4441,N_4044);
and U4516 (N_4516,N_4036,N_4125);
nand U4517 (N_4517,N_4225,N_4479);
and U4518 (N_4518,N_4394,N_4229);
nand U4519 (N_4519,N_4108,N_4013);
or U4520 (N_4520,N_4168,N_4467);
or U4521 (N_4521,N_4335,N_4000);
nor U4522 (N_4522,N_4182,N_4426);
nor U4523 (N_4523,N_4171,N_4421);
and U4524 (N_4524,N_4359,N_4481);
nor U4525 (N_4525,N_4149,N_4155);
nor U4526 (N_4526,N_4489,N_4360);
and U4527 (N_4527,N_4255,N_4179);
nor U4528 (N_4528,N_4174,N_4161);
or U4529 (N_4529,N_4178,N_4304);
nand U4530 (N_4530,N_4234,N_4320);
nor U4531 (N_4531,N_4358,N_4166);
and U4532 (N_4532,N_4429,N_4019);
or U4533 (N_4533,N_4387,N_4212);
xnor U4534 (N_4534,N_4159,N_4420);
and U4535 (N_4535,N_4193,N_4008);
or U4536 (N_4536,N_4145,N_4100);
and U4537 (N_4537,N_4361,N_4014);
nand U4538 (N_4538,N_4050,N_4404);
nand U4539 (N_4539,N_4490,N_4121);
or U4540 (N_4540,N_4456,N_4236);
or U4541 (N_4541,N_4460,N_4343);
or U4542 (N_4542,N_4114,N_4244);
nor U4543 (N_4543,N_4455,N_4332);
or U4544 (N_4544,N_4334,N_4286);
nor U4545 (N_4545,N_4115,N_4138);
nor U4546 (N_4546,N_4103,N_4160);
nor U4547 (N_4547,N_4336,N_4275);
nand U4548 (N_4548,N_4357,N_4246);
or U4549 (N_4549,N_4427,N_4068);
nor U4550 (N_4550,N_4450,N_4060);
nand U4551 (N_4551,N_4177,N_4063);
nand U4552 (N_4552,N_4051,N_4292);
and U4553 (N_4553,N_4081,N_4002);
nor U4554 (N_4554,N_4154,N_4491);
nand U4555 (N_4555,N_4459,N_4092);
nor U4556 (N_4556,N_4041,N_4312);
nand U4557 (N_4557,N_4118,N_4348);
nor U4558 (N_4558,N_4475,N_4205);
nor U4559 (N_4559,N_4274,N_4009);
or U4560 (N_4560,N_4362,N_4383);
or U4561 (N_4561,N_4465,N_4367);
and U4562 (N_4562,N_4314,N_4285);
and U4563 (N_4563,N_4442,N_4026);
nand U4564 (N_4564,N_4268,N_4064);
and U4565 (N_4565,N_4085,N_4293);
nand U4566 (N_4566,N_4452,N_4474);
nand U4567 (N_4567,N_4352,N_4127);
or U4568 (N_4568,N_4252,N_4142);
and U4569 (N_4569,N_4144,N_4038);
nor U4570 (N_4570,N_4073,N_4366);
and U4571 (N_4571,N_4102,N_4133);
or U4572 (N_4572,N_4445,N_4470);
and U4573 (N_4573,N_4084,N_4472);
or U4574 (N_4574,N_4416,N_4165);
nand U4575 (N_4575,N_4215,N_4313);
and U4576 (N_4576,N_4284,N_4095);
and U4577 (N_4577,N_4485,N_4399);
and U4578 (N_4578,N_4307,N_4087);
nor U4579 (N_4579,N_4153,N_4053);
nor U4580 (N_4580,N_4424,N_4403);
nor U4581 (N_4581,N_4120,N_4059);
nand U4582 (N_4582,N_4072,N_4024);
nor U4583 (N_4583,N_4037,N_4065);
and U4584 (N_4584,N_4356,N_4273);
or U4585 (N_4585,N_4116,N_4058);
and U4586 (N_4586,N_4278,N_4070);
nor U4587 (N_4587,N_4499,N_4400);
nor U4588 (N_4588,N_4388,N_4172);
or U4589 (N_4589,N_4486,N_4040);
or U4590 (N_4590,N_4451,N_4319);
nand U4591 (N_4591,N_4305,N_4079);
nor U4592 (N_4592,N_4266,N_4328);
nand U4593 (N_4593,N_4497,N_4419);
nor U4594 (N_4594,N_4439,N_4287);
nand U4595 (N_4595,N_4022,N_4281);
and U4596 (N_4596,N_4480,N_4230);
or U4597 (N_4597,N_4025,N_4156);
nand U4598 (N_4598,N_4458,N_4264);
and U4599 (N_4599,N_4323,N_4047);
nor U4600 (N_4600,N_4240,N_4373);
and U4601 (N_4601,N_4482,N_4422);
nand U4602 (N_4602,N_4123,N_4436);
nor U4603 (N_4603,N_4301,N_4327);
or U4604 (N_4604,N_4330,N_4146);
nor U4605 (N_4605,N_4325,N_4231);
and U4606 (N_4606,N_4297,N_4376);
nand U4607 (N_4607,N_4341,N_4391);
nor U4608 (N_4608,N_4170,N_4074);
or U4609 (N_4609,N_4350,N_4030);
and U4610 (N_4610,N_4412,N_4232);
nor U4611 (N_4611,N_4069,N_4031);
nand U4612 (N_4612,N_4483,N_4162);
or U4613 (N_4613,N_4315,N_4484);
or U4614 (N_4614,N_4487,N_4078);
nor U4615 (N_4615,N_4261,N_4141);
nand U4616 (N_4616,N_4071,N_4457);
and U4617 (N_4617,N_4222,N_4158);
nand U4618 (N_4618,N_4052,N_4094);
and U4619 (N_4619,N_4112,N_4128);
or U4620 (N_4620,N_4432,N_4076);
or U4621 (N_4621,N_4289,N_4017);
nand U4622 (N_4622,N_4126,N_4157);
and U4623 (N_4623,N_4408,N_4453);
nand U4624 (N_4624,N_4001,N_4196);
and U4625 (N_4625,N_4077,N_4163);
and U4626 (N_4626,N_4033,N_4414);
and U4627 (N_4627,N_4106,N_4117);
nand U4628 (N_4628,N_4433,N_4418);
nand U4629 (N_4629,N_4498,N_4093);
nand U4630 (N_4630,N_4318,N_4204);
and U4631 (N_4631,N_4132,N_4438);
or U4632 (N_4632,N_4294,N_4295);
nor U4633 (N_4633,N_4021,N_4454);
and U4634 (N_4634,N_4462,N_4034);
or U4635 (N_4635,N_4267,N_4492);
nor U4636 (N_4636,N_4221,N_4018);
or U4637 (N_4637,N_4351,N_4463);
nor U4638 (N_4638,N_4124,N_4396);
xor U4639 (N_4639,N_4371,N_4331);
nand U4640 (N_4640,N_4216,N_4277);
nor U4641 (N_4641,N_4242,N_4184);
and U4642 (N_4642,N_4005,N_4187);
and U4643 (N_4643,N_4353,N_4091);
and U4644 (N_4644,N_4004,N_4136);
nor U4645 (N_4645,N_4464,N_4238);
and U4646 (N_4646,N_4218,N_4340);
nand U4647 (N_4647,N_4099,N_4435);
nand U4648 (N_4648,N_4390,N_4046);
nand U4649 (N_4649,N_4039,N_4345);
nor U4650 (N_4650,N_4322,N_4338);
or U4651 (N_4651,N_4140,N_4368);
nand U4652 (N_4652,N_4235,N_4471);
or U4653 (N_4653,N_4259,N_4096);
or U4654 (N_4654,N_4233,N_4192);
and U4655 (N_4655,N_4382,N_4056);
or U4656 (N_4656,N_4282,N_4449);
or U4657 (N_4657,N_4310,N_4027);
or U4658 (N_4658,N_4023,N_4260);
and U4659 (N_4659,N_4150,N_4347);
or U4660 (N_4660,N_4185,N_4443);
xnor U4661 (N_4661,N_4029,N_4202);
or U4662 (N_4662,N_4151,N_4250);
or U4663 (N_4663,N_4300,N_4137);
or U4664 (N_4664,N_4398,N_4473);
or U4665 (N_4665,N_4245,N_4003);
nor U4666 (N_4666,N_4210,N_4113);
and U4667 (N_4667,N_4183,N_4379);
or U4668 (N_4668,N_4386,N_4385);
and U4669 (N_4669,N_4227,N_4478);
nand U4670 (N_4670,N_4251,N_4321);
nand U4671 (N_4671,N_4198,N_4135);
xor U4672 (N_4672,N_4049,N_4339);
nand U4673 (N_4673,N_4206,N_4105);
or U4674 (N_4674,N_4372,N_4254);
nand U4675 (N_4675,N_4493,N_4369);
and U4676 (N_4676,N_4007,N_4139);
nor U4677 (N_4677,N_4066,N_4377);
nor U4678 (N_4678,N_4173,N_4437);
nor U4679 (N_4679,N_4209,N_4283);
nand U4680 (N_4680,N_4256,N_4098);
and U4681 (N_4681,N_4263,N_4061);
and U4682 (N_4682,N_4265,N_4241);
nand U4683 (N_4683,N_4194,N_4190);
or U4684 (N_4684,N_4243,N_4344);
and U4685 (N_4685,N_4119,N_4374);
nand U4686 (N_4686,N_4111,N_4333);
and U4687 (N_4687,N_4337,N_4466);
nor U4688 (N_4688,N_4143,N_4197);
nor U4689 (N_4689,N_4262,N_4308);
nand U4690 (N_4690,N_4291,N_4211);
or U4691 (N_4691,N_4016,N_4164);
nor U4692 (N_4692,N_4446,N_4195);
nor U4693 (N_4693,N_4032,N_4224);
nand U4694 (N_4694,N_4354,N_4299);
or U4695 (N_4695,N_4257,N_4228);
nand U4696 (N_4696,N_4181,N_4279);
nand U4697 (N_4697,N_4272,N_4309);
or U4698 (N_4698,N_4496,N_4175);
and U4699 (N_4699,N_4363,N_4434);
nor U4700 (N_4700,N_4269,N_4169);
nand U4701 (N_4701,N_4208,N_4247);
nand U4702 (N_4702,N_4075,N_4249);
nand U4703 (N_4703,N_4296,N_4405);
nor U4704 (N_4704,N_4006,N_4042);
or U4705 (N_4705,N_4444,N_4089);
and U4706 (N_4706,N_4469,N_4237);
nand U4707 (N_4707,N_4280,N_4290);
and U4708 (N_4708,N_4349,N_4220);
or U4709 (N_4709,N_4213,N_4495);
and U4710 (N_4710,N_4461,N_4402);
nor U4711 (N_4711,N_4057,N_4413);
and U4712 (N_4712,N_4329,N_4270);
and U4713 (N_4713,N_4167,N_4048);
or U4714 (N_4714,N_4097,N_4045);
nor U4715 (N_4715,N_4415,N_4248);
or U4716 (N_4716,N_4122,N_4176);
nor U4717 (N_4717,N_4043,N_4430);
nor U4718 (N_4718,N_4088,N_4200);
nand U4719 (N_4719,N_4298,N_4326);
nand U4720 (N_4720,N_4381,N_4410);
and U4721 (N_4721,N_4306,N_4189);
nor U4722 (N_4722,N_4395,N_4080);
or U4723 (N_4723,N_4214,N_4110);
nand U4724 (N_4724,N_4423,N_4201);
nand U4725 (N_4725,N_4380,N_4276);
or U4726 (N_4726,N_4425,N_4109);
nor U4727 (N_4727,N_4203,N_4488);
or U4728 (N_4728,N_4086,N_4302);
or U4729 (N_4729,N_4134,N_4199);
nor U4730 (N_4730,N_4324,N_4082);
nand U4731 (N_4731,N_4219,N_4476);
nand U4732 (N_4732,N_4389,N_4411);
and U4733 (N_4733,N_4494,N_4448);
nor U4734 (N_4734,N_4180,N_4409);
nor U4735 (N_4735,N_4288,N_4147);
nor U4736 (N_4736,N_4188,N_4384);
and U4737 (N_4737,N_4401,N_4207);
nor U4738 (N_4738,N_4431,N_4012);
nor U4739 (N_4739,N_4406,N_4101);
nand U4740 (N_4740,N_4186,N_4062);
nand U4741 (N_4741,N_4152,N_4020);
nand U4742 (N_4742,N_4130,N_4253);
nand U4743 (N_4743,N_4239,N_4378);
nor U4744 (N_4744,N_4440,N_4407);
nand U4745 (N_4745,N_4393,N_4311);
and U4746 (N_4746,N_4226,N_4370);
nand U4747 (N_4747,N_4468,N_4129);
nor U4748 (N_4748,N_4417,N_4090);
nor U4749 (N_4749,N_4316,N_4271);
or U4750 (N_4750,N_4008,N_4493);
and U4751 (N_4751,N_4054,N_4213);
nand U4752 (N_4752,N_4265,N_4191);
nor U4753 (N_4753,N_4125,N_4074);
nor U4754 (N_4754,N_4328,N_4267);
nand U4755 (N_4755,N_4202,N_4265);
nand U4756 (N_4756,N_4373,N_4445);
or U4757 (N_4757,N_4497,N_4043);
and U4758 (N_4758,N_4353,N_4356);
and U4759 (N_4759,N_4485,N_4183);
nand U4760 (N_4760,N_4204,N_4178);
nor U4761 (N_4761,N_4156,N_4412);
nor U4762 (N_4762,N_4025,N_4389);
nor U4763 (N_4763,N_4062,N_4306);
nand U4764 (N_4764,N_4082,N_4240);
nand U4765 (N_4765,N_4172,N_4270);
and U4766 (N_4766,N_4126,N_4259);
and U4767 (N_4767,N_4494,N_4107);
nor U4768 (N_4768,N_4301,N_4424);
nand U4769 (N_4769,N_4151,N_4417);
nor U4770 (N_4770,N_4255,N_4319);
nor U4771 (N_4771,N_4119,N_4476);
nor U4772 (N_4772,N_4276,N_4130);
or U4773 (N_4773,N_4493,N_4378);
nand U4774 (N_4774,N_4333,N_4312);
nand U4775 (N_4775,N_4464,N_4414);
nor U4776 (N_4776,N_4174,N_4420);
and U4777 (N_4777,N_4025,N_4377);
nor U4778 (N_4778,N_4155,N_4080);
xor U4779 (N_4779,N_4135,N_4380);
nor U4780 (N_4780,N_4359,N_4476);
or U4781 (N_4781,N_4158,N_4126);
nor U4782 (N_4782,N_4177,N_4105);
and U4783 (N_4783,N_4299,N_4291);
or U4784 (N_4784,N_4411,N_4313);
or U4785 (N_4785,N_4354,N_4224);
and U4786 (N_4786,N_4421,N_4030);
or U4787 (N_4787,N_4495,N_4497);
or U4788 (N_4788,N_4167,N_4470);
nand U4789 (N_4789,N_4276,N_4040);
nor U4790 (N_4790,N_4024,N_4277);
and U4791 (N_4791,N_4165,N_4234);
nand U4792 (N_4792,N_4311,N_4255);
or U4793 (N_4793,N_4013,N_4028);
nor U4794 (N_4794,N_4427,N_4044);
nand U4795 (N_4795,N_4246,N_4156);
or U4796 (N_4796,N_4494,N_4119);
and U4797 (N_4797,N_4041,N_4386);
nand U4798 (N_4798,N_4433,N_4463);
or U4799 (N_4799,N_4084,N_4089);
nand U4800 (N_4800,N_4071,N_4181);
and U4801 (N_4801,N_4298,N_4169);
or U4802 (N_4802,N_4203,N_4374);
or U4803 (N_4803,N_4214,N_4203);
nor U4804 (N_4804,N_4145,N_4315);
and U4805 (N_4805,N_4461,N_4414);
nand U4806 (N_4806,N_4159,N_4161);
and U4807 (N_4807,N_4206,N_4199);
or U4808 (N_4808,N_4177,N_4044);
and U4809 (N_4809,N_4150,N_4372);
nor U4810 (N_4810,N_4358,N_4399);
and U4811 (N_4811,N_4247,N_4210);
nor U4812 (N_4812,N_4498,N_4344);
nand U4813 (N_4813,N_4048,N_4196);
or U4814 (N_4814,N_4338,N_4411);
and U4815 (N_4815,N_4109,N_4003);
nand U4816 (N_4816,N_4047,N_4128);
nand U4817 (N_4817,N_4193,N_4156);
and U4818 (N_4818,N_4495,N_4166);
nor U4819 (N_4819,N_4112,N_4347);
nand U4820 (N_4820,N_4211,N_4235);
nand U4821 (N_4821,N_4237,N_4363);
or U4822 (N_4822,N_4416,N_4111);
nand U4823 (N_4823,N_4448,N_4378);
nor U4824 (N_4824,N_4129,N_4154);
nor U4825 (N_4825,N_4079,N_4031);
and U4826 (N_4826,N_4419,N_4350);
or U4827 (N_4827,N_4219,N_4040);
and U4828 (N_4828,N_4399,N_4064);
and U4829 (N_4829,N_4251,N_4026);
nand U4830 (N_4830,N_4328,N_4323);
and U4831 (N_4831,N_4155,N_4373);
or U4832 (N_4832,N_4015,N_4475);
and U4833 (N_4833,N_4116,N_4161);
and U4834 (N_4834,N_4263,N_4476);
or U4835 (N_4835,N_4450,N_4454);
or U4836 (N_4836,N_4164,N_4130);
and U4837 (N_4837,N_4374,N_4404);
and U4838 (N_4838,N_4245,N_4275);
or U4839 (N_4839,N_4105,N_4134);
nor U4840 (N_4840,N_4339,N_4189);
nand U4841 (N_4841,N_4085,N_4448);
or U4842 (N_4842,N_4188,N_4342);
and U4843 (N_4843,N_4490,N_4152);
and U4844 (N_4844,N_4069,N_4432);
nand U4845 (N_4845,N_4109,N_4456);
and U4846 (N_4846,N_4482,N_4062);
nand U4847 (N_4847,N_4175,N_4051);
or U4848 (N_4848,N_4299,N_4199);
nor U4849 (N_4849,N_4405,N_4374);
or U4850 (N_4850,N_4339,N_4082);
nor U4851 (N_4851,N_4209,N_4377);
nand U4852 (N_4852,N_4067,N_4148);
nand U4853 (N_4853,N_4419,N_4461);
and U4854 (N_4854,N_4177,N_4214);
or U4855 (N_4855,N_4319,N_4218);
nand U4856 (N_4856,N_4271,N_4348);
nand U4857 (N_4857,N_4085,N_4056);
and U4858 (N_4858,N_4349,N_4195);
and U4859 (N_4859,N_4127,N_4048);
nor U4860 (N_4860,N_4025,N_4349);
and U4861 (N_4861,N_4460,N_4369);
nor U4862 (N_4862,N_4198,N_4043);
or U4863 (N_4863,N_4327,N_4112);
nand U4864 (N_4864,N_4342,N_4456);
nand U4865 (N_4865,N_4324,N_4453);
and U4866 (N_4866,N_4170,N_4423);
nor U4867 (N_4867,N_4388,N_4435);
nand U4868 (N_4868,N_4009,N_4117);
and U4869 (N_4869,N_4027,N_4391);
or U4870 (N_4870,N_4250,N_4031);
nor U4871 (N_4871,N_4487,N_4314);
nor U4872 (N_4872,N_4346,N_4038);
nor U4873 (N_4873,N_4170,N_4102);
nor U4874 (N_4874,N_4009,N_4139);
and U4875 (N_4875,N_4412,N_4246);
and U4876 (N_4876,N_4362,N_4308);
xnor U4877 (N_4877,N_4086,N_4105);
and U4878 (N_4878,N_4121,N_4478);
and U4879 (N_4879,N_4445,N_4071);
nand U4880 (N_4880,N_4048,N_4495);
nor U4881 (N_4881,N_4128,N_4183);
or U4882 (N_4882,N_4233,N_4139);
or U4883 (N_4883,N_4401,N_4376);
and U4884 (N_4884,N_4274,N_4479);
or U4885 (N_4885,N_4129,N_4120);
and U4886 (N_4886,N_4179,N_4144);
and U4887 (N_4887,N_4029,N_4002);
or U4888 (N_4888,N_4218,N_4249);
nor U4889 (N_4889,N_4100,N_4073);
nand U4890 (N_4890,N_4246,N_4101);
or U4891 (N_4891,N_4230,N_4145);
nor U4892 (N_4892,N_4214,N_4170);
nand U4893 (N_4893,N_4418,N_4259);
and U4894 (N_4894,N_4239,N_4111);
and U4895 (N_4895,N_4308,N_4121);
nor U4896 (N_4896,N_4430,N_4264);
or U4897 (N_4897,N_4160,N_4004);
and U4898 (N_4898,N_4413,N_4309);
nor U4899 (N_4899,N_4054,N_4417);
nor U4900 (N_4900,N_4272,N_4032);
or U4901 (N_4901,N_4084,N_4402);
nand U4902 (N_4902,N_4000,N_4444);
nand U4903 (N_4903,N_4320,N_4259);
nor U4904 (N_4904,N_4325,N_4334);
nand U4905 (N_4905,N_4017,N_4452);
nand U4906 (N_4906,N_4238,N_4075);
or U4907 (N_4907,N_4354,N_4452);
and U4908 (N_4908,N_4345,N_4156);
nor U4909 (N_4909,N_4290,N_4241);
nor U4910 (N_4910,N_4089,N_4409);
nor U4911 (N_4911,N_4480,N_4336);
or U4912 (N_4912,N_4255,N_4052);
or U4913 (N_4913,N_4438,N_4027);
or U4914 (N_4914,N_4259,N_4017);
nor U4915 (N_4915,N_4168,N_4066);
or U4916 (N_4916,N_4130,N_4225);
and U4917 (N_4917,N_4335,N_4217);
xnor U4918 (N_4918,N_4371,N_4035);
nor U4919 (N_4919,N_4441,N_4054);
nor U4920 (N_4920,N_4462,N_4096);
or U4921 (N_4921,N_4009,N_4302);
nand U4922 (N_4922,N_4412,N_4301);
xnor U4923 (N_4923,N_4419,N_4480);
and U4924 (N_4924,N_4221,N_4470);
and U4925 (N_4925,N_4345,N_4231);
and U4926 (N_4926,N_4168,N_4125);
nand U4927 (N_4927,N_4417,N_4150);
nor U4928 (N_4928,N_4331,N_4459);
nor U4929 (N_4929,N_4109,N_4081);
and U4930 (N_4930,N_4388,N_4338);
or U4931 (N_4931,N_4261,N_4052);
or U4932 (N_4932,N_4383,N_4228);
nand U4933 (N_4933,N_4127,N_4064);
and U4934 (N_4934,N_4308,N_4294);
or U4935 (N_4935,N_4434,N_4174);
or U4936 (N_4936,N_4322,N_4487);
nand U4937 (N_4937,N_4359,N_4226);
and U4938 (N_4938,N_4382,N_4155);
nor U4939 (N_4939,N_4385,N_4228);
or U4940 (N_4940,N_4291,N_4187);
nand U4941 (N_4941,N_4271,N_4180);
nand U4942 (N_4942,N_4498,N_4468);
nor U4943 (N_4943,N_4139,N_4462);
nand U4944 (N_4944,N_4218,N_4200);
nor U4945 (N_4945,N_4196,N_4159);
nor U4946 (N_4946,N_4256,N_4229);
or U4947 (N_4947,N_4254,N_4225);
nand U4948 (N_4948,N_4488,N_4338);
and U4949 (N_4949,N_4349,N_4131);
or U4950 (N_4950,N_4389,N_4229);
nand U4951 (N_4951,N_4246,N_4271);
and U4952 (N_4952,N_4112,N_4079);
nand U4953 (N_4953,N_4327,N_4136);
or U4954 (N_4954,N_4364,N_4401);
nor U4955 (N_4955,N_4193,N_4282);
or U4956 (N_4956,N_4266,N_4371);
or U4957 (N_4957,N_4229,N_4479);
or U4958 (N_4958,N_4027,N_4389);
nor U4959 (N_4959,N_4483,N_4185);
nand U4960 (N_4960,N_4160,N_4156);
xnor U4961 (N_4961,N_4128,N_4291);
and U4962 (N_4962,N_4299,N_4349);
and U4963 (N_4963,N_4086,N_4265);
or U4964 (N_4964,N_4376,N_4375);
nand U4965 (N_4965,N_4293,N_4363);
nor U4966 (N_4966,N_4001,N_4023);
nand U4967 (N_4967,N_4223,N_4258);
nand U4968 (N_4968,N_4122,N_4135);
and U4969 (N_4969,N_4345,N_4073);
or U4970 (N_4970,N_4499,N_4310);
and U4971 (N_4971,N_4336,N_4262);
nand U4972 (N_4972,N_4441,N_4304);
or U4973 (N_4973,N_4291,N_4222);
nor U4974 (N_4974,N_4282,N_4311);
or U4975 (N_4975,N_4418,N_4054);
nor U4976 (N_4976,N_4322,N_4194);
or U4977 (N_4977,N_4171,N_4493);
and U4978 (N_4978,N_4002,N_4241);
nand U4979 (N_4979,N_4170,N_4144);
nor U4980 (N_4980,N_4403,N_4087);
nor U4981 (N_4981,N_4321,N_4137);
and U4982 (N_4982,N_4349,N_4274);
and U4983 (N_4983,N_4403,N_4385);
and U4984 (N_4984,N_4391,N_4273);
or U4985 (N_4985,N_4026,N_4046);
and U4986 (N_4986,N_4250,N_4416);
xnor U4987 (N_4987,N_4018,N_4148);
nand U4988 (N_4988,N_4104,N_4311);
nand U4989 (N_4989,N_4387,N_4494);
nand U4990 (N_4990,N_4373,N_4053);
and U4991 (N_4991,N_4201,N_4017);
or U4992 (N_4992,N_4122,N_4439);
nand U4993 (N_4993,N_4265,N_4396);
nor U4994 (N_4994,N_4498,N_4111);
nand U4995 (N_4995,N_4255,N_4177);
or U4996 (N_4996,N_4003,N_4140);
nor U4997 (N_4997,N_4157,N_4213);
nor U4998 (N_4998,N_4007,N_4152);
nor U4999 (N_4999,N_4461,N_4210);
and UO_0 (O_0,N_4510,N_4837);
nand UO_1 (O_1,N_4756,N_4905);
nand UO_2 (O_2,N_4772,N_4954);
nand UO_3 (O_3,N_4561,N_4707);
and UO_4 (O_4,N_4949,N_4600);
or UO_5 (O_5,N_4721,N_4853);
nand UO_6 (O_6,N_4697,N_4701);
or UO_7 (O_7,N_4942,N_4613);
nand UO_8 (O_8,N_4585,N_4826);
nand UO_9 (O_9,N_4528,N_4946);
and UO_10 (O_10,N_4705,N_4931);
or UO_11 (O_11,N_4828,N_4529);
or UO_12 (O_12,N_4676,N_4717);
or UO_13 (O_13,N_4646,N_4879);
nor UO_14 (O_14,N_4806,N_4777);
or UO_15 (O_15,N_4752,N_4961);
nor UO_16 (O_16,N_4750,N_4790);
nand UO_17 (O_17,N_4770,N_4941);
and UO_18 (O_18,N_4531,N_4596);
nor UO_19 (O_19,N_4645,N_4923);
nor UO_20 (O_20,N_4698,N_4597);
or UO_21 (O_21,N_4798,N_4805);
and UO_22 (O_22,N_4735,N_4556);
and UO_23 (O_23,N_4587,N_4835);
nand UO_24 (O_24,N_4520,N_4714);
and UO_25 (O_25,N_4788,N_4847);
and UO_26 (O_26,N_4845,N_4882);
or UO_27 (O_27,N_4724,N_4868);
nand UO_28 (O_28,N_4661,N_4778);
or UO_29 (O_29,N_4896,N_4784);
nor UO_30 (O_30,N_4738,N_4821);
and UO_31 (O_31,N_4617,N_4981);
and UO_32 (O_32,N_4681,N_4878);
nand UO_33 (O_33,N_4508,N_4733);
nand UO_34 (O_34,N_4631,N_4774);
or UO_35 (O_35,N_4743,N_4918);
or UO_36 (O_36,N_4940,N_4582);
and UO_37 (O_37,N_4516,N_4865);
nand UO_38 (O_38,N_4749,N_4950);
and UO_39 (O_39,N_4550,N_4881);
nand UO_40 (O_40,N_4635,N_4848);
nand UO_41 (O_41,N_4824,N_4975);
nor UO_42 (O_42,N_4639,N_4511);
nand UO_43 (O_43,N_4892,N_4939);
and UO_44 (O_44,N_4518,N_4991);
or UO_45 (O_45,N_4519,N_4870);
nand UO_46 (O_46,N_4889,N_4786);
nor UO_47 (O_47,N_4998,N_4982);
and UO_48 (O_48,N_4906,N_4803);
nand UO_49 (O_49,N_4653,N_4539);
and UO_50 (O_50,N_4545,N_4685);
nor UO_51 (O_51,N_4968,N_4551);
nand UO_52 (O_52,N_4537,N_4827);
nor UO_53 (O_53,N_4789,N_4568);
nand UO_54 (O_54,N_4976,N_4920);
nor UO_55 (O_55,N_4504,N_4542);
nor UO_56 (O_56,N_4844,N_4863);
or UO_57 (O_57,N_4693,N_4605);
nor UO_58 (O_58,N_4572,N_4978);
and UO_59 (O_59,N_4754,N_4933);
nor UO_60 (O_60,N_4867,N_4802);
nand UO_61 (O_61,N_4783,N_4581);
and UO_62 (O_62,N_4830,N_4875);
nand UO_63 (O_63,N_4745,N_4758);
and UO_64 (O_64,N_4913,N_4618);
nor UO_65 (O_65,N_4718,N_4562);
or UO_66 (O_66,N_4921,N_4690);
and UO_67 (O_67,N_4570,N_4595);
nand UO_68 (O_68,N_4955,N_4934);
and UO_69 (O_69,N_4655,N_4814);
nand UO_70 (O_70,N_4994,N_4573);
and UO_71 (O_71,N_4993,N_4593);
nand UO_72 (O_72,N_4672,N_4914);
and UO_73 (O_73,N_4632,N_4773);
nor UO_74 (O_74,N_4692,N_4682);
nand UO_75 (O_75,N_4732,N_4804);
nand UO_76 (O_76,N_4709,N_4604);
nand UO_77 (O_77,N_4759,N_4967);
or UO_78 (O_78,N_4623,N_4677);
nand UO_79 (O_79,N_4696,N_4811);
or UO_80 (O_80,N_4795,N_4535);
nand UO_81 (O_81,N_4793,N_4796);
nand UO_82 (O_82,N_4671,N_4703);
nor UO_83 (O_83,N_4584,N_4995);
nor UO_84 (O_84,N_4959,N_4722);
nand UO_85 (O_85,N_4615,N_4546);
and UO_86 (O_86,N_4927,N_4842);
and UO_87 (O_87,N_4638,N_4549);
nand UO_88 (O_88,N_4829,N_4856);
or UO_89 (O_89,N_4876,N_4599);
xnor UO_90 (O_90,N_4836,N_4651);
nor UO_91 (O_91,N_4574,N_4740);
nand UO_92 (O_92,N_4607,N_4739);
and UO_93 (O_93,N_4898,N_4753);
or UO_94 (O_94,N_4997,N_4764);
or UO_95 (O_95,N_4598,N_4782);
and UO_96 (O_96,N_4747,N_4935);
or UO_97 (O_97,N_4833,N_4929);
and UO_98 (O_98,N_4684,N_4680);
and UO_99 (O_99,N_4660,N_4669);
or UO_100 (O_100,N_4970,N_4823);
nand UO_101 (O_101,N_4822,N_4964);
nor UO_102 (O_102,N_4943,N_4899);
nor UO_103 (O_103,N_4649,N_4616);
nor UO_104 (O_104,N_4885,N_4855);
nor UO_105 (O_105,N_4808,N_4736);
or UO_106 (O_106,N_4951,N_4800);
nand UO_107 (O_107,N_4577,N_4700);
or UO_108 (O_108,N_4502,N_4817);
and UO_109 (O_109,N_4711,N_4591);
and UO_110 (O_110,N_4769,N_4731);
and UO_111 (O_111,N_4971,N_4647);
nor UO_112 (O_112,N_4857,N_4579);
nand UO_113 (O_113,N_4636,N_4974);
nor UO_114 (O_114,N_4987,N_4633);
nor UO_115 (O_115,N_4544,N_4626);
nand UO_116 (O_116,N_4787,N_4999);
nand UO_117 (O_117,N_4849,N_4525);
nand UO_118 (O_118,N_4619,N_4917);
and UO_119 (O_119,N_4812,N_4872);
or UO_120 (O_120,N_4728,N_4864);
nor UO_121 (O_121,N_4586,N_4859);
and UO_122 (O_122,N_4761,N_4886);
nand UO_123 (O_123,N_4503,N_4694);
nand UO_124 (O_124,N_4891,N_4513);
or UO_125 (O_125,N_4780,N_4792);
nand UO_126 (O_126,N_4926,N_4507);
and UO_127 (O_127,N_4751,N_4742);
or UO_128 (O_128,N_4937,N_4530);
or UO_129 (O_129,N_4583,N_4763);
or UO_130 (O_130,N_4960,N_4894);
and UO_131 (O_131,N_4944,N_4624);
nor UO_132 (O_132,N_4990,N_4702);
nor UO_133 (O_133,N_4664,N_4558);
nor UO_134 (O_134,N_4904,N_4547);
nand UO_135 (O_135,N_4930,N_4858);
nand UO_136 (O_136,N_4601,N_4956);
nand UO_137 (O_137,N_4767,N_4526);
nor UO_138 (O_138,N_4992,N_4922);
and UO_139 (O_139,N_4972,N_4958);
or UO_140 (O_140,N_4688,N_4871);
nand UO_141 (O_141,N_4654,N_4797);
nor UO_142 (O_142,N_4720,N_4665);
nor UO_143 (O_143,N_4907,N_4678);
nor UO_144 (O_144,N_4683,N_4541);
nor UO_145 (O_145,N_4575,N_4565);
nor UO_146 (O_146,N_4602,N_4534);
nor UO_147 (O_147,N_4980,N_4928);
or UO_148 (O_148,N_4815,N_4533);
nand UO_149 (O_149,N_4536,N_4819);
nor UO_150 (O_150,N_4948,N_4887);
and UO_151 (O_151,N_4524,N_4839);
or UO_152 (O_152,N_4768,N_4622);
and UO_153 (O_153,N_4932,N_4608);
nor UO_154 (O_154,N_4912,N_4554);
or UO_155 (O_155,N_4877,N_4840);
nor UO_156 (O_156,N_4523,N_4625);
or UO_157 (O_157,N_4652,N_4675);
or UO_158 (O_158,N_4983,N_4755);
nand UO_159 (O_159,N_4820,N_4566);
or UO_160 (O_160,N_4816,N_4838);
nor UO_161 (O_161,N_4679,N_4637);
and UO_162 (O_162,N_4668,N_4686);
or UO_163 (O_163,N_4883,N_4947);
nor UO_164 (O_164,N_4910,N_4852);
nor UO_165 (O_165,N_4966,N_4590);
and UO_166 (O_166,N_4563,N_4843);
or UO_167 (O_167,N_4807,N_4667);
and UO_168 (O_168,N_4741,N_4716);
nor UO_169 (O_169,N_4785,N_4903);
nor UO_170 (O_170,N_4609,N_4710);
nor UO_171 (O_171,N_4952,N_4571);
xor UO_172 (O_172,N_4986,N_4874);
and UO_173 (O_173,N_4908,N_4517);
nor UO_174 (O_174,N_4532,N_4775);
and UO_175 (O_175,N_4614,N_4901);
nand UO_176 (O_176,N_4965,N_4687);
nor UO_177 (O_177,N_4580,N_4712);
nor UO_178 (O_178,N_4897,N_4522);
or UO_179 (O_179,N_4880,N_4620);
nand UO_180 (O_180,N_4500,N_4592);
nor UO_181 (O_181,N_4611,N_4977);
or UO_182 (O_182,N_4666,N_4854);
or UO_183 (O_183,N_4989,N_4984);
and UO_184 (O_184,N_4644,N_4726);
and UO_185 (O_185,N_4559,N_4776);
nor UO_186 (O_186,N_4569,N_4553);
and UO_187 (O_187,N_4866,N_4578);
nor UO_188 (O_188,N_4628,N_4893);
or UO_189 (O_189,N_4902,N_4634);
nor UO_190 (O_190,N_4670,N_4564);
and UO_191 (O_191,N_4725,N_4869);
and UO_192 (O_192,N_4936,N_4713);
and UO_193 (O_193,N_4794,N_4540);
nor UO_194 (O_194,N_4506,N_4945);
or UO_195 (O_195,N_4861,N_4734);
nand UO_196 (O_196,N_4727,N_4737);
nor UO_197 (O_197,N_4695,N_4860);
and UO_198 (O_198,N_4663,N_4691);
and UO_199 (O_199,N_4706,N_4729);
or UO_200 (O_200,N_4674,N_4801);
nand UO_201 (O_201,N_4909,N_4715);
nand UO_202 (O_202,N_4548,N_4643);
nor UO_203 (O_203,N_4630,N_4594);
and UO_204 (O_204,N_4650,N_4543);
nand UO_205 (O_205,N_4762,N_4527);
nand UO_206 (O_206,N_4621,N_4973);
nand UO_207 (O_207,N_4689,N_4746);
nand UO_208 (O_208,N_4825,N_4810);
nor UO_209 (O_209,N_4567,N_4719);
and UO_210 (O_210,N_4560,N_4779);
nand UO_211 (O_211,N_4841,N_4962);
or UO_212 (O_212,N_4509,N_4610);
xnor UO_213 (O_213,N_4834,N_4799);
nor UO_214 (O_214,N_4642,N_4873);
nor UO_215 (O_215,N_4552,N_4919);
and UO_216 (O_216,N_4514,N_4765);
or UO_217 (O_217,N_4915,N_4809);
nand UO_218 (O_218,N_4505,N_4699);
nand UO_219 (O_219,N_4832,N_4521);
or UO_220 (O_220,N_4888,N_4862);
or UO_221 (O_221,N_4771,N_4766);
or UO_222 (O_222,N_4629,N_4723);
nor UO_223 (O_223,N_4659,N_4657);
and UO_224 (O_224,N_4900,N_4953);
nand UO_225 (O_225,N_4791,N_4851);
or UO_226 (O_226,N_4818,N_4760);
and UO_227 (O_227,N_4979,N_4603);
or UO_228 (O_228,N_4831,N_4656);
and UO_229 (O_229,N_4938,N_4606);
and UO_230 (O_230,N_4969,N_4730);
and UO_231 (O_231,N_4708,N_4996);
nor UO_232 (O_232,N_4658,N_4895);
nand UO_233 (O_233,N_4925,N_4850);
and UO_234 (O_234,N_4640,N_4641);
nand UO_235 (O_235,N_4813,N_4648);
or UO_236 (O_236,N_4916,N_4627);
or UO_237 (O_237,N_4911,N_4512);
and UO_238 (O_238,N_4884,N_4963);
nand UO_239 (O_239,N_4988,N_4515);
nand UO_240 (O_240,N_4538,N_4576);
nand UO_241 (O_241,N_4924,N_4781);
nor UO_242 (O_242,N_4557,N_4501);
and UO_243 (O_243,N_4757,N_4588);
or UO_244 (O_244,N_4846,N_4555);
or UO_245 (O_245,N_4985,N_4662);
or UO_246 (O_246,N_4748,N_4890);
and UO_247 (O_247,N_4704,N_4744);
and UO_248 (O_248,N_4957,N_4612);
nor UO_249 (O_249,N_4673,N_4589);
and UO_250 (O_250,N_4743,N_4865);
nand UO_251 (O_251,N_4704,N_4742);
and UO_252 (O_252,N_4886,N_4599);
nor UO_253 (O_253,N_4551,N_4742);
nand UO_254 (O_254,N_4738,N_4776);
nor UO_255 (O_255,N_4692,N_4506);
and UO_256 (O_256,N_4777,N_4906);
and UO_257 (O_257,N_4873,N_4542);
and UO_258 (O_258,N_4610,N_4599);
or UO_259 (O_259,N_4567,N_4935);
and UO_260 (O_260,N_4663,N_4717);
nand UO_261 (O_261,N_4573,N_4702);
or UO_262 (O_262,N_4773,N_4887);
nand UO_263 (O_263,N_4529,N_4506);
and UO_264 (O_264,N_4845,N_4613);
or UO_265 (O_265,N_4892,N_4654);
nand UO_266 (O_266,N_4538,N_4635);
or UO_267 (O_267,N_4618,N_4662);
nand UO_268 (O_268,N_4776,N_4765);
and UO_269 (O_269,N_4975,N_4705);
nand UO_270 (O_270,N_4878,N_4620);
or UO_271 (O_271,N_4718,N_4825);
nor UO_272 (O_272,N_4543,N_4610);
nand UO_273 (O_273,N_4631,N_4523);
or UO_274 (O_274,N_4996,N_4674);
and UO_275 (O_275,N_4690,N_4966);
nand UO_276 (O_276,N_4929,N_4740);
nor UO_277 (O_277,N_4633,N_4557);
nand UO_278 (O_278,N_4566,N_4605);
nand UO_279 (O_279,N_4787,N_4845);
nand UO_280 (O_280,N_4905,N_4941);
or UO_281 (O_281,N_4819,N_4967);
or UO_282 (O_282,N_4895,N_4974);
nor UO_283 (O_283,N_4726,N_4949);
nand UO_284 (O_284,N_4884,N_4635);
or UO_285 (O_285,N_4542,N_4899);
or UO_286 (O_286,N_4666,N_4581);
nor UO_287 (O_287,N_4840,N_4943);
and UO_288 (O_288,N_4842,N_4777);
or UO_289 (O_289,N_4657,N_4665);
xnor UO_290 (O_290,N_4803,N_4532);
nand UO_291 (O_291,N_4932,N_4826);
or UO_292 (O_292,N_4735,N_4721);
or UO_293 (O_293,N_4580,N_4962);
nand UO_294 (O_294,N_4759,N_4632);
nand UO_295 (O_295,N_4544,N_4889);
or UO_296 (O_296,N_4716,N_4594);
or UO_297 (O_297,N_4828,N_4765);
and UO_298 (O_298,N_4586,N_4722);
or UO_299 (O_299,N_4596,N_4775);
nor UO_300 (O_300,N_4697,N_4549);
xnor UO_301 (O_301,N_4849,N_4621);
nand UO_302 (O_302,N_4865,N_4639);
or UO_303 (O_303,N_4696,N_4500);
nor UO_304 (O_304,N_4836,N_4942);
nand UO_305 (O_305,N_4630,N_4813);
nand UO_306 (O_306,N_4972,N_4751);
or UO_307 (O_307,N_4842,N_4679);
and UO_308 (O_308,N_4983,N_4924);
or UO_309 (O_309,N_4787,N_4559);
or UO_310 (O_310,N_4978,N_4930);
nand UO_311 (O_311,N_4843,N_4802);
or UO_312 (O_312,N_4803,N_4946);
or UO_313 (O_313,N_4809,N_4901);
and UO_314 (O_314,N_4812,N_4918);
nor UO_315 (O_315,N_4809,N_4732);
or UO_316 (O_316,N_4648,N_4725);
nor UO_317 (O_317,N_4962,N_4689);
nand UO_318 (O_318,N_4758,N_4951);
and UO_319 (O_319,N_4909,N_4904);
or UO_320 (O_320,N_4902,N_4726);
and UO_321 (O_321,N_4984,N_4943);
nand UO_322 (O_322,N_4913,N_4634);
or UO_323 (O_323,N_4983,N_4757);
and UO_324 (O_324,N_4776,N_4709);
xnor UO_325 (O_325,N_4755,N_4981);
or UO_326 (O_326,N_4505,N_4816);
or UO_327 (O_327,N_4872,N_4808);
nand UO_328 (O_328,N_4875,N_4869);
and UO_329 (O_329,N_4908,N_4777);
xnor UO_330 (O_330,N_4846,N_4907);
nor UO_331 (O_331,N_4681,N_4952);
and UO_332 (O_332,N_4531,N_4681);
or UO_333 (O_333,N_4678,N_4613);
and UO_334 (O_334,N_4684,N_4595);
nand UO_335 (O_335,N_4545,N_4713);
and UO_336 (O_336,N_4837,N_4853);
or UO_337 (O_337,N_4975,N_4543);
nand UO_338 (O_338,N_4764,N_4932);
nor UO_339 (O_339,N_4874,N_4529);
nand UO_340 (O_340,N_4775,N_4827);
and UO_341 (O_341,N_4640,N_4707);
nor UO_342 (O_342,N_4604,N_4724);
and UO_343 (O_343,N_4511,N_4781);
or UO_344 (O_344,N_4906,N_4734);
and UO_345 (O_345,N_4995,N_4645);
or UO_346 (O_346,N_4914,N_4704);
xnor UO_347 (O_347,N_4657,N_4909);
nor UO_348 (O_348,N_4513,N_4536);
and UO_349 (O_349,N_4677,N_4828);
or UO_350 (O_350,N_4806,N_4624);
nor UO_351 (O_351,N_4943,N_4564);
nand UO_352 (O_352,N_4781,N_4617);
nor UO_353 (O_353,N_4611,N_4863);
nand UO_354 (O_354,N_4963,N_4560);
and UO_355 (O_355,N_4983,N_4777);
nand UO_356 (O_356,N_4697,N_4562);
nand UO_357 (O_357,N_4862,N_4927);
nand UO_358 (O_358,N_4694,N_4616);
nor UO_359 (O_359,N_4737,N_4830);
nand UO_360 (O_360,N_4735,N_4662);
nand UO_361 (O_361,N_4825,N_4716);
nand UO_362 (O_362,N_4589,N_4566);
nand UO_363 (O_363,N_4553,N_4661);
or UO_364 (O_364,N_4916,N_4863);
nor UO_365 (O_365,N_4604,N_4967);
and UO_366 (O_366,N_4523,N_4524);
nand UO_367 (O_367,N_4876,N_4859);
nand UO_368 (O_368,N_4612,N_4944);
or UO_369 (O_369,N_4725,N_4828);
and UO_370 (O_370,N_4531,N_4989);
and UO_371 (O_371,N_4898,N_4819);
and UO_372 (O_372,N_4970,N_4615);
nand UO_373 (O_373,N_4773,N_4940);
and UO_374 (O_374,N_4618,N_4782);
or UO_375 (O_375,N_4574,N_4585);
nand UO_376 (O_376,N_4823,N_4991);
nand UO_377 (O_377,N_4854,N_4990);
and UO_378 (O_378,N_4894,N_4978);
and UO_379 (O_379,N_4565,N_4660);
nor UO_380 (O_380,N_4759,N_4879);
and UO_381 (O_381,N_4962,N_4517);
nor UO_382 (O_382,N_4810,N_4617);
nor UO_383 (O_383,N_4607,N_4513);
and UO_384 (O_384,N_4716,N_4788);
nand UO_385 (O_385,N_4679,N_4568);
nor UO_386 (O_386,N_4792,N_4735);
nor UO_387 (O_387,N_4564,N_4645);
and UO_388 (O_388,N_4700,N_4823);
and UO_389 (O_389,N_4881,N_4502);
or UO_390 (O_390,N_4637,N_4583);
and UO_391 (O_391,N_4623,N_4665);
nor UO_392 (O_392,N_4776,N_4835);
and UO_393 (O_393,N_4528,N_4785);
and UO_394 (O_394,N_4704,N_4762);
nor UO_395 (O_395,N_4843,N_4645);
nor UO_396 (O_396,N_4528,N_4795);
nor UO_397 (O_397,N_4736,N_4598);
xor UO_398 (O_398,N_4965,N_4654);
and UO_399 (O_399,N_4517,N_4558);
nor UO_400 (O_400,N_4897,N_4823);
nand UO_401 (O_401,N_4815,N_4943);
nand UO_402 (O_402,N_4836,N_4758);
nor UO_403 (O_403,N_4989,N_4567);
or UO_404 (O_404,N_4678,N_4667);
nor UO_405 (O_405,N_4897,N_4793);
and UO_406 (O_406,N_4506,N_4888);
or UO_407 (O_407,N_4795,N_4743);
or UO_408 (O_408,N_4848,N_4646);
or UO_409 (O_409,N_4965,N_4732);
nor UO_410 (O_410,N_4554,N_4627);
and UO_411 (O_411,N_4796,N_4562);
and UO_412 (O_412,N_4632,N_4531);
and UO_413 (O_413,N_4879,N_4660);
nor UO_414 (O_414,N_4980,N_4991);
nor UO_415 (O_415,N_4682,N_4770);
nand UO_416 (O_416,N_4985,N_4659);
and UO_417 (O_417,N_4978,N_4920);
and UO_418 (O_418,N_4663,N_4695);
nor UO_419 (O_419,N_4708,N_4947);
or UO_420 (O_420,N_4582,N_4800);
nand UO_421 (O_421,N_4616,N_4577);
nand UO_422 (O_422,N_4921,N_4696);
or UO_423 (O_423,N_4513,N_4935);
nor UO_424 (O_424,N_4914,N_4737);
or UO_425 (O_425,N_4605,N_4921);
nand UO_426 (O_426,N_4751,N_4766);
or UO_427 (O_427,N_4907,N_4988);
and UO_428 (O_428,N_4924,N_4551);
or UO_429 (O_429,N_4645,N_4935);
and UO_430 (O_430,N_4785,N_4711);
and UO_431 (O_431,N_4869,N_4908);
nor UO_432 (O_432,N_4811,N_4816);
and UO_433 (O_433,N_4585,N_4695);
nand UO_434 (O_434,N_4585,N_4615);
nor UO_435 (O_435,N_4941,N_4773);
nand UO_436 (O_436,N_4524,N_4712);
and UO_437 (O_437,N_4988,N_4826);
nand UO_438 (O_438,N_4774,N_4996);
nand UO_439 (O_439,N_4525,N_4768);
nor UO_440 (O_440,N_4909,N_4554);
nor UO_441 (O_441,N_4974,N_4611);
or UO_442 (O_442,N_4641,N_4974);
or UO_443 (O_443,N_4866,N_4558);
and UO_444 (O_444,N_4976,N_4817);
nand UO_445 (O_445,N_4545,N_4628);
nand UO_446 (O_446,N_4869,N_4646);
nand UO_447 (O_447,N_4751,N_4998);
or UO_448 (O_448,N_4586,N_4512);
nor UO_449 (O_449,N_4845,N_4725);
or UO_450 (O_450,N_4857,N_4921);
and UO_451 (O_451,N_4526,N_4567);
or UO_452 (O_452,N_4613,N_4745);
nor UO_453 (O_453,N_4646,N_4860);
and UO_454 (O_454,N_4742,N_4706);
nand UO_455 (O_455,N_4806,N_4869);
nand UO_456 (O_456,N_4962,N_4760);
nor UO_457 (O_457,N_4881,N_4818);
and UO_458 (O_458,N_4534,N_4829);
and UO_459 (O_459,N_4851,N_4578);
or UO_460 (O_460,N_4739,N_4510);
and UO_461 (O_461,N_4791,N_4937);
xnor UO_462 (O_462,N_4769,N_4869);
or UO_463 (O_463,N_4618,N_4874);
and UO_464 (O_464,N_4943,N_4623);
nand UO_465 (O_465,N_4984,N_4710);
or UO_466 (O_466,N_4602,N_4945);
nand UO_467 (O_467,N_4664,N_4739);
nand UO_468 (O_468,N_4748,N_4556);
and UO_469 (O_469,N_4862,N_4843);
and UO_470 (O_470,N_4957,N_4659);
nor UO_471 (O_471,N_4579,N_4745);
nand UO_472 (O_472,N_4523,N_4501);
and UO_473 (O_473,N_4688,N_4845);
nor UO_474 (O_474,N_4529,N_4890);
and UO_475 (O_475,N_4829,N_4656);
or UO_476 (O_476,N_4634,N_4933);
and UO_477 (O_477,N_4903,N_4829);
nand UO_478 (O_478,N_4719,N_4685);
nand UO_479 (O_479,N_4669,N_4680);
or UO_480 (O_480,N_4837,N_4805);
nand UO_481 (O_481,N_4678,N_4670);
and UO_482 (O_482,N_4804,N_4655);
and UO_483 (O_483,N_4852,N_4968);
and UO_484 (O_484,N_4819,N_4726);
or UO_485 (O_485,N_4888,N_4864);
nor UO_486 (O_486,N_4726,N_4719);
or UO_487 (O_487,N_4874,N_4599);
nor UO_488 (O_488,N_4560,N_4529);
or UO_489 (O_489,N_4930,N_4702);
xnor UO_490 (O_490,N_4522,N_4887);
nor UO_491 (O_491,N_4818,N_4563);
or UO_492 (O_492,N_4922,N_4769);
and UO_493 (O_493,N_4889,N_4927);
or UO_494 (O_494,N_4922,N_4975);
nand UO_495 (O_495,N_4961,N_4812);
and UO_496 (O_496,N_4534,N_4610);
and UO_497 (O_497,N_4898,N_4763);
nor UO_498 (O_498,N_4743,N_4809);
and UO_499 (O_499,N_4752,N_4872);
or UO_500 (O_500,N_4559,N_4838);
or UO_501 (O_501,N_4819,N_4854);
nor UO_502 (O_502,N_4987,N_4934);
and UO_503 (O_503,N_4691,N_4777);
or UO_504 (O_504,N_4645,N_4830);
and UO_505 (O_505,N_4734,N_4970);
or UO_506 (O_506,N_4635,N_4609);
or UO_507 (O_507,N_4786,N_4950);
nor UO_508 (O_508,N_4798,N_4747);
nand UO_509 (O_509,N_4575,N_4874);
and UO_510 (O_510,N_4505,N_4961);
or UO_511 (O_511,N_4877,N_4856);
nor UO_512 (O_512,N_4613,N_4689);
and UO_513 (O_513,N_4889,N_4622);
nor UO_514 (O_514,N_4694,N_4613);
or UO_515 (O_515,N_4521,N_4532);
nor UO_516 (O_516,N_4755,N_4706);
xnor UO_517 (O_517,N_4596,N_4626);
nor UO_518 (O_518,N_4614,N_4537);
or UO_519 (O_519,N_4679,N_4693);
nand UO_520 (O_520,N_4986,N_4971);
and UO_521 (O_521,N_4919,N_4618);
nand UO_522 (O_522,N_4513,N_4561);
nand UO_523 (O_523,N_4665,N_4694);
nor UO_524 (O_524,N_4696,N_4866);
nand UO_525 (O_525,N_4837,N_4854);
or UO_526 (O_526,N_4999,N_4560);
or UO_527 (O_527,N_4834,N_4581);
or UO_528 (O_528,N_4887,N_4633);
nand UO_529 (O_529,N_4901,N_4562);
nand UO_530 (O_530,N_4636,N_4575);
nor UO_531 (O_531,N_4697,N_4533);
or UO_532 (O_532,N_4870,N_4502);
nor UO_533 (O_533,N_4575,N_4816);
or UO_534 (O_534,N_4925,N_4653);
nor UO_535 (O_535,N_4660,N_4691);
nor UO_536 (O_536,N_4660,N_4538);
and UO_537 (O_537,N_4815,N_4924);
nor UO_538 (O_538,N_4928,N_4777);
or UO_539 (O_539,N_4884,N_4922);
nand UO_540 (O_540,N_4901,N_4945);
and UO_541 (O_541,N_4925,N_4629);
nor UO_542 (O_542,N_4914,N_4680);
or UO_543 (O_543,N_4708,N_4841);
nand UO_544 (O_544,N_4615,N_4567);
and UO_545 (O_545,N_4919,N_4891);
and UO_546 (O_546,N_4751,N_4565);
nand UO_547 (O_547,N_4918,N_4863);
nand UO_548 (O_548,N_4788,N_4561);
or UO_549 (O_549,N_4628,N_4734);
and UO_550 (O_550,N_4542,N_4612);
nand UO_551 (O_551,N_4571,N_4850);
and UO_552 (O_552,N_4666,N_4542);
and UO_553 (O_553,N_4536,N_4894);
nor UO_554 (O_554,N_4987,N_4781);
and UO_555 (O_555,N_4961,N_4766);
nor UO_556 (O_556,N_4990,N_4848);
nor UO_557 (O_557,N_4611,N_4876);
nor UO_558 (O_558,N_4636,N_4706);
nand UO_559 (O_559,N_4719,N_4563);
or UO_560 (O_560,N_4673,N_4505);
nand UO_561 (O_561,N_4778,N_4649);
nor UO_562 (O_562,N_4856,N_4755);
nor UO_563 (O_563,N_4929,N_4537);
or UO_564 (O_564,N_4799,N_4905);
nor UO_565 (O_565,N_4608,N_4917);
nor UO_566 (O_566,N_4835,N_4592);
and UO_567 (O_567,N_4523,N_4919);
nand UO_568 (O_568,N_4528,N_4752);
nand UO_569 (O_569,N_4659,N_4609);
or UO_570 (O_570,N_4714,N_4756);
nand UO_571 (O_571,N_4739,N_4612);
and UO_572 (O_572,N_4808,N_4777);
nand UO_573 (O_573,N_4616,N_4523);
or UO_574 (O_574,N_4934,N_4865);
nand UO_575 (O_575,N_4728,N_4588);
nor UO_576 (O_576,N_4717,N_4659);
and UO_577 (O_577,N_4881,N_4888);
nand UO_578 (O_578,N_4604,N_4926);
nor UO_579 (O_579,N_4755,N_4797);
or UO_580 (O_580,N_4939,N_4770);
or UO_581 (O_581,N_4535,N_4767);
nand UO_582 (O_582,N_4751,N_4634);
nand UO_583 (O_583,N_4530,N_4963);
and UO_584 (O_584,N_4713,N_4558);
and UO_585 (O_585,N_4710,N_4975);
nand UO_586 (O_586,N_4882,N_4957);
nand UO_587 (O_587,N_4751,N_4562);
or UO_588 (O_588,N_4958,N_4832);
and UO_589 (O_589,N_4526,N_4991);
and UO_590 (O_590,N_4508,N_4554);
or UO_591 (O_591,N_4920,N_4685);
nand UO_592 (O_592,N_4955,N_4938);
and UO_593 (O_593,N_4850,N_4554);
nand UO_594 (O_594,N_4752,N_4846);
and UO_595 (O_595,N_4643,N_4953);
or UO_596 (O_596,N_4877,N_4772);
nor UO_597 (O_597,N_4651,N_4794);
nand UO_598 (O_598,N_4619,N_4633);
and UO_599 (O_599,N_4696,N_4884);
or UO_600 (O_600,N_4525,N_4670);
nor UO_601 (O_601,N_4659,N_4961);
or UO_602 (O_602,N_4968,N_4936);
or UO_603 (O_603,N_4610,N_4955);
and UO_604 (O_604,N_4713,N_4908);
nand UO_605 (O_605,N_4996,N_4764);
and UO_606 (O_606,N_4963,N_4851);
nor UO_607 (O_607,N_4612,N_4583);
nor UO_608 (O_608,N_4697,N_4770);
or UO_609 (O_609,N_4757,N_4572);
or UO_610 (O_610,N_4979,N_4636);
nand UO_611 (O_611,N_4740,N_4763);
and UO_612 (O_612,N_4904,N_4561);
and UO_613 (O_613,N_4599,N_4870);
nand UO_614 (O_614,N_4904,N_4678);
or UO_615 (O_615,N_4549,N_4601);
or UO_616 (O_616,N_4835,N_4548);
nand UO_617 (O_617,N_4778,N_4930);
or UO_618 (O_618,N_4630,N_4640);
nand UO_619 (O_619,N_4658,N_4705);
and UO_620 (O_620,N_4990,N_4804);
or UO_621 (O_621,N_4619,N_4901);
nand UO_622 (O_622,N_4895,N_4851);
nor UO_623 (O_623,N_4718,N_4699);
nor UO_624 (O_624,N_4907,N_4956);
nand UO_625 (O_625,N_4717,N_4874);
nor UO_626 (O_626,N_4657,N_4737);
and UO_627 (O_627,N_4974,N_4577);
and UO_628 (O_628,N_4937,N_4817);
nand UO_629 (O_629,N_4738,N_4530);
nor UO_630 (O_630,N_4804,N_4960);
or UO_631 (O_631,N_4874,N_4588);
and UO_632 (O_632,N_4963,N_4787);
or UO_633 (O_633,N_4568,N_4769);
and UO_634 (O_634,N_4546,N_4552);
or UO_635 (O_635,N_4971,N_4749);
nand UO_636 (O_636,N_4997,N_4683);
nand UO_637 (O_637,N_4965,N_4879);
and UO_638 (O_638,N_4537,N_4747);
and UO_639 (O_639,N_4971,N_4531);
or UO_640 (O_640,N_4510,N_4835);
or UO_641 (O_641,N_4846,N_4724);
nand UO_642 (O_642,N_4859,N_4983);
nor UO_643 (O_643,N_4609,N_4702);
nor UO_644 (O_644,N_4815,N_4828);
or UO_645 (O_645,N_4771,N_4910);
nand UO_646 (O_646,N_4897,N_4886);
nor UO_647 (O_647,N_4960,N_4604);
nand UO_648 (O_648,N_4906,N_4792);
nor UO_649 (O_649,N_4721,N_4800);
nand UO_650 (O_650,N_4532,N_4537);
nor UO_651 (O_651,N_4862,N_4631);
nor UO_652 (O_652,N_4882,N_4965);
and UO_653 (O_653,N_4684,N_4809);
nand UO_654 (O_654,N_4871,N_4794);
or UO_655 (O_655,N_4958,N_4921);
and UO_656 (O_656,N_4728,N_4536);
and UO_657 (O_657,N_4864,N_4777);
and UO_658 (O_658,N_4958,N_4699);
or UO_659 (O_659,N_4609,N_4591);
nor UO_660 (O_660,N_4912,N_4783);
nand UO_661 (O_661,N_4712,N_4888);
and UO_662 (O_662,N_4627,N_4736);
nor UO_663 (O_663,N_4968,N_4948);
nor UO_664 (O_664,N_4521,N_4655);
and UO_665 (O_665,N_4644,N_4793);
or UO_666 (O_666,N_4576,N_4764);
nand UO_667 (O_667,N_4834,N_4940);
or UO_668 (O_668,N_4793,N_4948);
and UO_669 (O_669,N_4517,N_4666);
and UO_670 (O_670,N_4896,N_4732);
nand UO_671 (O_671,N_4995,N_4796);
nor UO_672 (O_672,N_4996,N_4532);
and UO_673 (O_673,N_4695,N_4953);
or UO_674 (O_674,N_4732,N_4920);
or UO_675 (O_675,N_4528,N_4669);
nand UO_676 (O_676,N_4594,N_4701);
or UO_677 (O_677,N_4943,N_4909);
nor UO_678 (O_678,N_4738,N_4522);
nand UO_679 (O_679,N_4699,N_4515);
nand UO_680 (O_680,N_4580,N_4842);
or UO_681 (O_681,N_4576,N_4731);
nand UO_682 (O_682,N_4740,N_4873);
and UO_683 (O_683,N_4809,N_4516);
and UO_684 (O_684,N_4761,N_4865);
and UO_685 (O_685,N_4964,N_4896);
and UO_686 (O_686,N_4595,N_4766);
and UO_687 (O_687,N_4754,N_4893);
or UO_688 (O_688,N_4694,N_4631);
or UO_689 (O_689,N_4839,N_4628);
nor UO_690 (O_690,N_4791,N_4636);
nand UO_691 (O_691,N_4528,N_4662);
or UO_692 (O_692,N_4988,N_4894);
nor UO_693 (O_693,N_4577,N_4969);
nand UO_694 (O_694,N_4579,N_4627);
and UO_695 (O_695,N_4716,N_4537);
nor UO_696 (O_696,N_4865,N_4924);
xnor UO_697 (O_697,N_4687,N_4913);
or UO_698 (O_698,N_4659,N_4903);
or UO_699 (O_699,N_4915,N_4647);
nand UO_700 (O_700,N_4825,N_4748);
and UO_701 (O_701,N_4658,N_4975);
or UO_702 (O_702,N_4739,N_4519);
or UO_703 (O_703,N_4956,N_4828);
and UO_704 (O_704,N_4996,N_4726);
and UO_705 (O_705,N_4510,N_4504);
and UO_706 (O_706,N_4701,N_4896);
nand UO_707 (O_707,N_4701,N_4504);
nor UO_708 (O_708,N_4591,N_4736);
nand UO_709 (O_709,N_4742,N_4750);
and UO_710 (O_710,N_4995,N_4625);
nor UO_711 (O_711,N_4606,N_4763);
and UO_712 (O_712,N_4877,N_4548);
xnor UO_713 (O_713,N_4751,N_4720);
nand UO_714 (O_714,N_4718,N_4591);
nand UO_715 (O_715,N_4846,N_4642);
nand UO_716 (O_716,N_4964,N_4781);
nand UO_717 (O_717,N_4597,N_4916);
and UO_718 (O_718,N_4500,N_4714);
nand UO_719 (O_719,N_4835,N_4746);
nand UO_720 (O_720,N_4929,N_4541);
or UO_721 (O_721,N_4712,N_4685);
and UO_722 (O_722,N_4581,N_4872);
and UO_723 (O_723,N_4929,N_4500);
and UO_724 (O_724,N_4615,N_4853);
and UO_725 (O_725,N_4677,N_4952);
and UO_726 (O_726,N_4651,N_4744);
nand UO_727 (O_727,N_4708,N_4620);
or UO_728 (O_728,N_4538,N_4781);
nor UO_729 (O_729,N_4814,N_4749);
nand UO_730 (O_730,N_4715,N_4663);
or UO_731 (O_731,N_4770,N_4506);
nand UO_732 (O_732,N_4771,N_4700);
nor UO_733 (O_733,N_4952,N_4533);
or UO_734 (O_734,N_4648,N_4502);
or UO_735 (O_735,N_4663,N_4552);
and UO_736 (O_736,N_4675,N_4794);
and UO_737 (O_737,N_4747,N_4712);
or UO_738 (O_738,N_4688,N_4722);
or UO_739 (O_739,N_4720,N_4766);
or UO_740 (O_740,N_4565,N_4628);
nor UO_741 (O_741,N_4549,N_4741);
and UO_742 (O_742,N_4691,N_4647);
nor UO_743 (O_743,N_4782,N_4588);
nor UO_744 (O_744,N_4689,N_4720);
and UO_745 (O_745,N_4583,N_4820);
nor UO_746 (O_746,N_4621,N_4946);
or UO_747 (O_747,N_4732,N_4579);
or UO_748 (O_748,N_4916,N_4677);
nor UO_749 (O_749,N_4733,N_4541);
or UO_750 (O_750,N_4929,N_4662);
and UO_751 (O_751,N_4511,N_4785);
nor UO_752 (O_752,N_4858,N_4688);
nor UO_753 (O_753,N_4672,N_4970);
xnor UO_754 (O_754,N_4609,N_4904);
or UO_755 (O_755,N_4672,N_4851);
nor UO_756 (O_756,N_4677,N_4736);
or UO_757 (O_757,N_4854,N_4936);
xnor UO_758 (O_758,N_4890,N_4736);
nor UO_759 (O_759,N_4725,N_4599);
or UO_760 (O_760,N_4728,N_4551);
nor UO_761 (O_761,N_4977,N_4923);
and UO_762 (O_762,N_4804,N_4615);
nand UO_763 (O_763,N_4595,N_4654);
nand UO_764 (O_764,N_4639,N_4642);
and UO_765 (O_765,N_4941,N_4665);
nor UO_766 (O_766,N_4908,N_4647);
nand UO_767 (O_767,N_4685,N_4792);
nand UO_768 (O_768,N_4759,N_4989);
nand UO_769 (O_769,N_4544,N_4741);
or UO_770 (O_770,N_4576,N_4732);
nor UO_771 (O_771,N_4936,N_4971);
nand UO_772 (O_772,N_4517,N_4846);
nand UO_773 (O_773,N_4932,N_4525);
and UO_774 (O_774,N_4715,N_4681);
or UO_775 (O_775,N_4852,N_4615);
nand UO_776 (O_776,N_4668,N_4988);
nand UO_777 (O_777,N_4863,N_4740);
or UO_778 (O_778,N_4537,N_4505);
and UO_779 (O_779,N_4852,N_4811);
nand UO_780 (O_780,N_4584,N_4550);
or UO_781 (O_781,N_4528,N_4902);
and UO_782 (O_782,N_4722,N_4990);
nand UO_783 (O_783,N_4561,N_4674);
or UO_784 (O_784,N_4577,N_4973);
nor UO_785 (O_785,N_4595,N_4990);
nor UO_786 (O_786,N_4534,N_4722);
and UO_787 (O_787,N_4623,N_4596);
nor UO_788 (O_788,N_4622,N_4938);
and UO_789 (O_789,N_4946,N_4721);
nand UO_790 (O_790,N_4708,N_4931);
nand UO_791 (O_791,N_4621,N_4531);
nor UO_792 (O_792,N_4577,N_4983);
and UO_793 (O_793,N_4916,N_4967);
or UO_794 (O_794,N_4790,N_4847);
or UO_795 (O_795,N_4740,N_4867);
nand UO_796 (O_796,N_4908,N_4743);
or UO_797 (O_797,N_4936,N_4922);
nor UO_798 (O_798,N_4909,N_4687);
and UO_799 (O_799,N_4795,N_4767);
or UO_800 (O_800,N_4553,N_4902);
or UO_801 (O_801,N_4513,N_4751);
nor UO_802 (O_802,N_4831,N_4920);
or UO_803 (O_803,N_4874,N_4820);
nor UO_804 (O_804,N_4893,N_4582);
nand UO_805 (O_805,N_4870,N_4740);
and UO_806 (O_806,N_4687,N_4835);
nand UO_807 (O_807,N_4958,N_4509);
nand UO_808 (O_808,N_4951,N_4943);
nor UO_809 (O_809,N_4828,N_4746);
or UO_810 (O_810,N_4852,N_4825);
nor UO_811 (O_811,N_4689,N_4897);
and UO_812 (O_812,N_4847,N_4823);
and UO_813 (O_813,N_4639,N_4581);
nor UO_814 (O_814,N_4964,N_4907);
nand UO_815 (O_815,N_4764,N_4724);
nand UO_816 (O_816,N_4811,N_4626);
nand UO_817 (O_817,N_4659,N_4776);
nand UO_818 (O_818,N_4606,N_4936);
nor UO_819 (O_819,N_4786,N_4513);
or UO_820 (O_820,N_4615,N_4682);
nor UO_821 (O_821,N_4574,N_4963);
nand UO_822 (O_822,N_4951,N_4984);
and UO_823 (O_823,N_4605,N_4882);
or UO_824 (O_824,N_4838,N_4810);
and UO_825 (O_825,N_4847,N_4879);
and UO_826 (O_826,N_4926,N_4803);
or UO_827 (O_827,N_4704,N_4829);
or UO_828 (O_828,N_4925,N_4677);
and UO_829 (O_829,N_4669,N_4966);
or UO_830 (O_830,N_4875,N_4969);
and UO_831 (O_831,N_4922,N_4757);
and UO_832 (O_832,N_4826,N_4820);
or UO_833 (O_833,N_4676,N_4799);
and UO_834 (O_834,N_4618,N_4972);
or UO_835 (O_835,N_4854,N_4559);
or UO_836 (O_836,N_4792,N_4837);
nand UO_837 (O_837,N_4782,N_4686);
or UO_838 (O_838,N_4759,N_4915);
nand UO_839 (O_839,N_4558,N_4698);
nor UO_840 (O_840,N_4602,N_4966);
nand UO_841 (O_841,N_4644,N_4775);
nand UO_842 (O_842,N_4860,N_4981);
or UO_843 (O_843,N_4929,N_4736);
nor UO_844 (O_844,N_4646,N_4639);
nor UO_845 (O_845,N_4904,N_4644);
nor UO_846 (O_846,N_4734,N_4545);
nand UO_847 (O_847,N_4549,N_4604);
or UO_848 (O_848,N_4617,N_4504);
nand UO_849 (O_849,N_4776,N_4673);
or UO_850 (O_850,N_4838,N_4736);
nor UO_851 (O_851,N_4741,N_4588);
or UO_852 (O_852,N_4697,N_4519);
and UO_853 (O_853,N_4678,N_4802);
nand UO_854 (O_854,N_4772,N_4810);
nand UO_855 (O_855,N_4901,N_4850);
nand UO_856 (O_856,N_4768,N_4644);
and UO_857 (O_857,N_4823,N_4961);
nor UO_858 (O_858,N_4689,N_4826);
nand UO_859 (O_859,N_4500,N_4720);
or UO_860 (O_860,N_4621,N_4782);
nand UO_861 (O_861,N_4925,N_4549);
nor UO_862 (O_862,N_4715,N_4811);
nor UO_863 (O_863,N_4669,N_4604);
or UO_864 (O_864,N_4888,N_4511);
nand UO_865 (O_865,N_4683,N_4641);
or UO_866 (O_866,N_4752,N_4706);
nor UO_867 (O_867,N_4818,N_4724);
nor UO_868 (O_868,N_4729,N_4606);
or UO_869 (O_869,N_4573,N_4968);
or UO_870 (O_870,N_4573,N_4570);
nor UO_871 (O_871,N_4593,N_4552);
nor UO_872 (O_872,N_4729,N_4692);
and UO_873 (O_873,N_4515,N_4747);
or UO_874 (O_874,N_4601,N_4587);
nand UO_875 (O_875,N_4861,N_4701);
nor UO_876 (O_876,N_4654,N_4735);
nor UO_877 (O_877,N_4960,N_4703);
nand UO_878 (O_878,N_4951,N_4589);
or UO_879 (O_879,N_4637,N_4516);
and UO_880 (O_880,N_4884,N_4984);
nor UO_881 (O_881,N_4875,N_4712);
nand UO_882 (O_882,N_4522,N_4585);
nand UO_883 (O_883,N_4639,N_4821);
nor UO_884 (O_884,N_4982,N_4587);
nand UO_885 (O_885,N_4881,N_4988);
and UO_886 (O_886,N_4803,N_4932);
nor UO_887 (O_887,N_4511,N_4859);
and UO_888 (O_888,N_4997,N_4703);
or UO_889 (O_889,N_4794,N_4672);
nor UO_890 (O_890,N_4876,N_4782);
nor UO_891 (O_891,N_4543,N_4797);
nand UO_892 (O_892,N_4630,N_4738);
nor UO_893 (O_893,N_4572,N_4739);
and UO_894 (O_894,N_4926,N_4712);
and UO_895 (O_895,N_4877,N_4755);
and UO_896 (O_896,N_4655,N_4701);
nor UO_897 (O_897,N_4988,N_4595);
or UO_898 (O_898,N_4630,N_4769);
nand UO_899 (O_899,N_4663,N_4694);
nand UO_900 (O_900,N_4716,N_4703);
nor UO_901 (O_901,N_4717,N_4920);
nor UO_902 (O_902,N_4932,N_4930);
nand UO_903 (O_903,N_4693,N_4768);
nand UO_904 (O_904,N_4591,N_4973);
nor UO_905 (O_905,N_4942,N_4877);
and UO_906 (O_906,N_4526,N_4834);
or UO_907 (O_907,N_4848,N_4877);
nand UO_908 (O_908,N_4595,N_4593);
and UO_909 (O_909,N_4503,N_4820);
and UO_910 (O_910,N_4728,N_4627);
nand UO_911 (O_911,N_4656,N_4858);
nor UO_912 (O_912,N_4708,N_4527);
nor UO_913 (O_913,N_4595,N_4634);
nand UO_914 (O_914,N_4534,N_4738);
or UO_915 (O_915,N_4870,N_4997);
nor UO_916 (O_916,N_4872,N_4687);
or UO_917 (O_917,N_4973,N_4549);
nand UO_918 (O_918,N_4668,N_4899);
nor UO_919 (O_919,N_4538,N_4662);
nor UO_920 (O_920,N_4883,N_4944);
and UO_921 (O_921,N_4890,N_4744);
nor UO_922 (O_922,N_4994,N_4653);
or UO_923 (O_923,N_4579,N_4913);
nor UO_924 (O_924,N_4962,N_4605);
and UO_925 (O_925,N_4642,N_4523);
or UO_926 (O_926,N_4684,N_4822);
or UO_927 (O_927,N_4698,N_4899);
or UO_928 (O_928,N_4667,N_4851);
nor UO_929 (O_929,N_4693,N_4556);
or UO_930 (O_930,N_4746,N_4694);
nor UO_931 (O_931,N_4739,N_4708);
nor UO_932 (O_932,N_4829,N_4726);
or UO_933 (O_933,N_4948,N_4808);
or UO_934 (O_934,N_4615,N_4565);
nand UO_935 (O_935,N_4655,N_4602);
and UO_936 (O_936,N_4534,N_4860);
and UO_937 (O_937,N_4813,N_4961);
or UO_938 (O_938,N_4769,N_4800);
nand UO_939 (O_939,N_4999,N_4588);
nor UO_940 (O_940,N_4653,N_4976);
or UO_941 (O_941,N_4910,N_4636);
or UO_942 (O_942,N_4546,N_4665);
nor UO_943 (O_943,N_4986,N_4966);
and UO_944 (O_944,N_4838,N_4768);
or UO_945 (O_945,N_4894,N_4967);
and UO_946 (O_946,N_4761,N_4685);
nor UO_947 (O_947,N_4549,N_4799);
nand UO_948 (O_948,N_4558,N_4687);
nor UO_949 (O_949,N_4596,N_4555);
or UO_950 (O_950,N_4849,N_4610);
and UO_951 (O_951,N_4937,N_4606);
or UO_952 (O_952,N_4746,N_4955);
nor UO_953 (O_953,N_4938,N_4939);
nor UO_954 (O_954,N_4716,N_4542);
or UO_955 (O_955,N_4980,N_4580);
or UO_956 (O_956,N_4930,N_4902);
and UO_957 (O_957,N_4781,N_4641);
nor UO_958 (O_958,N_4753,N_4656);
or UO_959 (O_959,N_4859,N_4844);
nand UO_960 (O_960,N_4656,N_4722);
nor UO_961 (O_961,N_4588,N_4962);
nand UO_962 (O_962,N_4715,N_4741);
xnor UO_963 (O_963,N_4860,N_4764);
or UO_964 (O_964,N_4717,N_4891);
and UO_965 (O_965,N_4637,N_4810);
nand UO_966 (O_966,N_4529,N_4953);
and UO_967 (O_967,N_4590,N_4659);
nand UO_968 (O_968,N_4831,N_4658);
or UO_969 (O_969,N_4986,N_4813);
nor UO_970 (O_970,N_4959,N_4861);
nand UO_971 (O_971,N_4978,N_4908);
or UO_972 (O_972,N_4556,N_4864);
or UO_973 (O_973,N_4546,N_4708);
nor UO_974 (O_974,N_4847,N_4987);
nand UO_975 (O_975,N_4871,N_4653);
or UO_976 (O_976,N_4533,N_4727);
nor UO_977 (O_977,N_4717,N_4836);
or UO_978 (O_978,N_4677,N_4912);
nor UO_979 (O_979,N_4801,N_4788);
nand UO_980 (O_980,N_4527,N_4600);
and UO_981 (O_981,N_4763,N_4610);
and UO_982 (O_982,N_4977,N_4532);
nor UO_983 (O_983,N_4946,N_4556);
nor UO_984 (O_984,N_4822,N_4742);
nor UO_985 (O_985,N_4729,N_4939);
nor UO_986 (O_986,N_4825,N_4806);
nor UO_987 (O_987,N_4686,N_4815);
nand UO_988 (O_988,N_4626,N_4535);
and UO_989 (O_989,N_4992,N_4715);
nor UO_990 (O_990,N_4714,N_4983);
and UO_991 (O_991,N_4720,N_4889);
or UO_992 (O_992,N_4659,N_4783);
nand UO_993 (O_993,N_4705,N_4616);
nor UO_994 (O_994,N_4732,N_4855);
nor UO_995 (O_995,N_4630,N_4788);
nor UO_996 (O_996,N_4878,N_4753);
and UO_997 (O_997,N_4718,N_4543);
nor UO_998 (O_998,N_4565,N_4827);
and UO_999 (O_999,N_4825,N_4904);
endmodule