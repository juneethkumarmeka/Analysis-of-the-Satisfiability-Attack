module basic_2000_20000_2500_25_levels_1xor_3(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999;
and U0 (N_0,In_1832,In_1781);
and U1 (N_1,In_76,In_211);
or U2 (N_2,In_1302,In_343);
nor U3 (N_3,In_300,In_762);
and U4 (N_4,In_1246,In_1917);
nor U5 (N_5,In_836,In_668);
nand U6 (N_6,In_523,In_1507);
nor U7 (N_7,In_129,In_355);
or U8 (N_8,In_12,In_698);
or U9 (N_9,In_414,In_958);
and U10 (N_10,In_530,In_89);
and U11 (N_11,In_2,In_205);
or U12 (N_12,In_715,In_815);
and U13 (N_13,In_1970,In_26);
nand U14 (N_14,In_311,In_1513);
or U15 (N_15,In_829,In_1236);
nand U16 (N_16,In_1481,In_734);
nor U17 (N_17,In_1399,In_1335);
and U18 (N_18,In_149,In_847);
nand U19 (N_19,In_1620,In_121);
nand U20 (N_20,In_957,In_1106);
nand U21 (N_21,In_156,In_552);
and U22 (N_22,In_1255,In_1313);
nor U23 (N_23,In_1024,In_585);
and U24 (N_24,In_475,In_1478);
or U25 (N_25,In_1558,In_1272);
nand U26 (N_26,In_747,In_545);
nand U27 (N_27,In_761,In_51);
and U28 (N_28,In_476,In_1654);
and U29 (N_29,In_1670,In_38);
nand U30 (N_30,In_727,In_204);
nand U31 (N_31,In_52,In_112);
or U32 (N_32,In_932,In_1695);
or U33 (N_33,In_1131,In_1805);
nand U34 (N_34,In_1322,In_1066);
and U35 (N_35,In_1646,In_831);
or U36 (N_36,In_213,In_411);
and U37 (N_37,In_1006,In_32);
nor U38 (N_38,In_1120,In_551);
nor U39 (N_39,In_1538,In_1264);
xor U40 (N_40,In_1325,In_499);
nor U41 (N_41,In_1133,In_1206);
or U42 (N_42,In_1569,In_1976);
or U43 (N_43,In_1678,In_1915);
nor U44 (N_44,In_303,In_309);
and U45 (N_45,In_192,In_925);
or U46 (N_46,In_1474,In_590);
or U47 (N_47,In_1005,In_1050);
or U48 (N_48,In_444,In_481);
and U49 (N_49,In_1825,In_262);
nand U50 (N_50,In_821,In_496);
nor U51 (N_51,In_1852,In_1922);
or U52 (N_52,In_1802,In_702);
nand U53 (N_53,In_1110,In_1531);
nor U54 (N_54,In_1925,In_1041);
nor U55 (N_55,In_1668,In_1998);
or U56 (N_56,In_943,In_75);
and U57 (N_57,In_998,In_507);
nand U58 (N_58,In_1116,In_1214);
and U59 (N_59,In_407,In_1383);
nor U60 (N_60,In_108,In_555);
or U61 (N_61,In_1426,In_1126);
and U62 (N_62,In_799,In_109);
nand U63 (N_63,In_498,In_738);
nand U64 (N_64,In_1659,In_660);
nor U65 (N_65,In_637,In_1866);
nand U66 (N_66,In_1934,In_1578);
nor U67 (N_67,In_61,In_1103);
or U68 (N_68,In_1550,In_1763);
nand U69 (N_69,In_621,In_512);
and U70 (N_70,In_1529,In_593);
or U71 (N_71,In_1964,In_1554);
nor U72 (N_72,In_1948,In_30);
or U73 (N_73,In_1703,In_1902);
or U74 (N_74,In_254,In_1197);
and U75 (N_75,In_1002,In_1095);
nand U76 (N_76,In_1499,In_751);
nor U77 (N_77,In_1109,In_986);
nand U78 (N_78,In_325,In_574);
and U79 (N_79,In_705,In_1848);
nor U80 (N_80,In_1527,In_1021);
and U81 (N_81,In_1138,In_1610);
nand U82 (N_82,In_361,In_1098);
nor U83 (N_83,In_996,In_1861);
nor U84 (N_84,In_1285,In_1308);
nand U85 (N_85,In_596,In_514);
and U86 (N_86,In_1331,In_1636);
nor U87 (N_87,In_1434,In_67);
or U88 (N_88,In_1039,In_603);
and U89 (N_89,In_914,In_510);
or U90 (N_90,In_859,In_1587);
nor U91 (N_91,In_468,In_676);
or U92 (N_92,In_169,In_1215);
or U93 (N_93,In_513,In_1705);
nand U94 (N_94,In_1018,In_1688);
and U95 (N_95,In_1762,In_1);
or U96 (N_96,In_106,In_173);
or U97 (N_97,In_1717,In_164);
and U98 (N_98,In_900,In_307);
nand U99 (N_99,In_1467,In_208);
or U100 (N_100,In_531,In_771);
nand U101 (N_101,In_1343,In_241);
nor U102 (N_102,In_1464,In_1580);
and U103 (N_103,In_1559,In_59);
nand U104 (N_104,In_1858,In_1985);
nor U105 (N_105,In_11,In_197);
nor U106 (N_106,In_1199,In_1704);
or U107 (N_107,In_728,In_1966);
nor U108 (N_108,In_759,In_455);
and U109 (N_109,In_260,In_147);
nand U110 (N_110,In_572,In_1774);
nand U111 (N_111,In_754,In_784);
or U112 (N_112,In_470,In_505);
or U113 (N_113,In_1873,In_1368);
nor U114 (N_114,In_820,In_1149);
nor U115 (N_115,In_394,In_1094);
and U116 (N_116,In_1952,In_934);
or U117 (N_117,In_1046,In_69);
or U118 (N_118,In_867,In_1223);
and U119 (N_119,In_1244,In_1818);
nand U120 (N_120,In_1552,In_1536);
or U121 (N_121,In_1471,In_678);
and U122 (N_122,In_1840,In_933);
or U123 (N_123,In_916,In_1652);
nand U124 (N_124,In_1674,In_1772);
nand U125 (N_125,In_1643,In_597);
and U126 (N_126,In_1437,In_1838);
nor U127 (N_127,In_691,In_722);
nor U128 (N_128,In_1993,In_1650);
and U129 (N_129,In_1594,In_923);
or U130 (N_130,In_1632,In_1248);
nand U131 (N_131,In_927,In_1905);
or U132 (N_132,In_1768,In_1773);
nand U133 (N_133,In_1614,In_285);
nor U134 (N_134,In_1961,In_1657);
nor U135 (N_135,In_351,In_1568);
nand U136 (N_136,In_618,In_221);
nor U137 (N_137,In_992,In_775);
or U138 (N_138,In_997,In_412);
or U139 (N_139,In_334,In_640);
and U140 (N_140,In_388,In_55);
nor U141 (N_141,In_263,In_1933);
nand U142 (N_142,In_35,In_1841);
nor U143 (N_143,In_605,In_1911);
nor U144 (N_144,In_1076,In_756);
nor U145 (N_145,In_1566,In_1789);
nand U146 (N_146,In_190,In_787);
or U147 (N_147,In_373,In_1876);
and U148 (N_148,In_1427,In_1582);
nor U149 (N_149,In_638,In_253);
nand U150 (N_150,In_716,In_97);
nand U151 (N_151,In_1565,In_993);
nand U152 (N_152,In_553,In_1546);
or U153 (N_153,In_864,In_1923);
nand U154 (N_154,In_124,In_1068);
and U155 (N_155,In_1386,In_1324);
nand U156 (N_156,In_1616,In_643);
or U157 (N_157,In_274,In_1301);
nor U158 (N_158,In_396,In_582);
nand U159 (N_159,In_318,In_1867);
nor U160 (N_160,In_162,In_717);
or U161 (N_161,In_764,In_130);
nor U162 (N_162,In_645,In_1300);
nand U163 (N_163,In_1227,In_1392);
or U164 (N_164,In_64,In_1907);
nor U165 (N_165,In_1353,In_460);
or U166 (N_166,In_1785,In_615);
nand U167 (N_167,In_85,In_1063);
and U168 (N_168,In_635,In_469);
and U169 (N_169,In_1350,In_1431);
and U170 (N_170,In_302,In_1412);
and U171 (N_171,In_65,In_338);
or U172 (N_172,In_1378,In_1183);
nand U173 (N_173,In_188,In_980);
and U174 (N_174,In_1526,In_1145);
and U175 (N_175,In_279,In_1401);
and U176 (N_176,In_1424,In_539);
or U177 (N_177,In_506,In_1433);
and U178 (N_178,In_180,In_199);
nor U179 (N_179,In_390,In_841);
or U180 (N_180,In_786,In_57);
nand U181 (N_181,In_966,In_973);
and U182 (N_182,In_508,In_752);
or U183 (N_183,In_1564,In_1776);
and U184 (N_184,In_662,In_904);
and U185 (N_185,In_406,In_1384);
and U186 (N_186,In_731,In_1168);
nand U187 (N_187,In_871,In_1791);
nor U188 (N_188,In_281,In_1254);
nor U189 (N_189,In_488,In_1816);
nand U190 (N_190,In_1760,In_589);
and U191 (N_191,In_389,In_1878);
or U192 (N_192,In_231,In_248);
nor U193 (N_193,In_432,In_382);
and U194 (N_194,In_686,In_275);
and U195 (N_195,In_1697,In_1675);
nor U196 (N_196,In_96,In_1330);
nor U197 (N_197,In_693,In_1294);
and U198 (N_198,In_570,In_1757);
nand U199 (N_199,In_1736,In_536);
or U200 (N_200,In_897,In_1243);
nand U201 (N_201,In_359,In_679);
nand U202 (N_202,In_667,In_1232);
nor U203 (N_203,In_940,In_6);
nor U204 (N_204,In_626,In_890);
or U205 (N_205,In_206,In_159);
nor U206 (N_206,In_988,In_1398);
nand U207 (N_207,In_1064,In_865);
nor U208 (N_208,In_1956,In_1344);
or U209 (N_209,In_1119,In_1411);
nor U210 (N_210,In_1879,In_360);
nand U211 (N_211,In_1169,In_910);
or U212 (N_212,In_104,In_1043);
nor U213 (N_213,In_824,In_1160);
or U214 (N_214,In_1758,In_1822);
or U215 (N_215,In_652,In_858);
nor U216 (N_216,In_987,In_749);
or U217 (N_217,In_167,In_181);
or U218 (N_218,In_1476,In_595);
nor U219 (N_219,In_1417,In_1851);
nor U220 (N_220,In_332,In_1159);
nor U221 (N_221,In_1814,In_519);
nand U222 (N_222,In_1171,In_1279);
nand U223 (N_223,In_802,In_410);
nor U224 (N_224,In_0,In_71);
or U225 (N_225,In_500,In_1714);
nor U226 (N_226,In_117,In_700);
nor U227 (N_227,In_979,In_1057);
nand U228 (N_228,In_244,In_1870);
nand U229 (N_229,In_1204,In_1836);
nor U230 (N_230,In_82,In_1102);
nand U231 (N_231,In_144,In_1919);
nor U232 (N_232,In_202,In_1699);
and U233 (N_233,In_1539,In_1249);
or U234 (N_234,In_1702,In_1056);
nor U235 (N_235,In_1731,In_1888);
or U236 (N_236,In_1777,In_758);
nor U237 (N_237,In_1549,In_225);
xnor U238 (N_238,In_1442,In_1400);
nor U239 (N_239,In_622,In_128);
nor U240 (N_240,In_1172,In_1872);
or U241 (N_241,In_1014,In_465);
nor U242 (N_242,In_15,In_368);
nand U243 (N_243,In_70,In_1282);
and U244 (N_244,In_520,In_354);
and U245 (N_245,In_466,In_1593);
or U246 (N_246,In_1782,In_1995);
nor U247 (N_247,In_1446,In_1196);
nand U248 (N_248,In_1557,In_636);
or U249 (N_249,In_264,In_1328);
nand U250 (N_250,In_322,In_1142);
and U251 (N_251,In_1257,In_1134);
and U252 (N_252,In_1741,In_1798);
or U253 (N_253,In_317,In_1058);
or U254 (N_254,In_218,In_1092);
nand U255 (N_255,In_863,In_477);
nor U256 (N_256,In_1892,In_1997);
or U257 (N_257,In_492,In_1860);
or U258 (N_258,In_895,In_464);
nand U259 (N_259,In_39,In_299);
nand U260 (N_260,In_4,In_1738);
and U261 (N_261,In_1337,In_245);
or U262 (N_262,In_1193,In_1069);
nor U263 (N_263,In_724,In_1684);
or U264 (N_264,In_1969,In_1755);
nand U265 (N_265,In_1287,In_1269);
and U266 (N_266,In_672,In_95);
or U267 (N_267,In_886,In_780);
nor U268 (N_268,In_653,In_1341);
nor U269 (N_269,In_803,In_21);
nor U270 (N_270,In_1960,In_398);
nor U271 (N_271,In_1391,In_341);
or U272 (N_272,In_1596,In_901);
or U273 (N_273,In_79,In_186);
nand U274 (N_274,In_814,In_546);
nor U275 (N_275,In_1543,In_1125);
nand U276 (N_276,In_86,In_1265);
or U277 (N_277,In_1886,In_1175);
nand U278 (N_278,In_563,In_400);
or U279 (N_279,In_1877,In_350);
nand U280 (N_280,In_669,In_798);
and U281 (N_281,In_684,In_982);
xnor U282 (N_282,In_326,In_1207);
nor U283 (N_283,In_1957,In_1490);
or U284 (N_284,In_1700,In_1649);
or U285 (N_285,In_1388,In_461);
and U286 (N_286,In_718,In_439);
nor U287 (N_287,In_1965,In_148);
or U288 (N_288,In_347,In_287);
xor U289 (N_289,In_330,In_687);
and U290 (N_290,In_493,In_557);
and U291 (N_291,In_538,In_66);
and U292 (N_292,In_1912,In_1304);
nand U293 (N_293,In_1259,In_591);
or U294 (N_294,In_1263,In_138);
or U295 (N_295,In_1454,In_27);
nand U296 (N_296,In_1184,In_319);
nand U297 (N_297,In_88,In_1036);
or U298 (N_298,In_402,In_223);
and U299 (N_299,In_1686,In_1622);
and U300 (N_300,In_1783,In_642);
nor U301 (N_301,In_1868,In_1205);
nand U302 (N_302,In_1091,In_879);
or U303 (N_303,In_1510,In_1979);
and U304 (N_304,In_954,In_975);
xor U305 (N_305,In_1638,In_1466);
nand U306 (N_306,In_189,In_1759);
and U307 (N_307,In_422,In_697);
or U308 (N_308,In_54,In_1753);
and U309 (N_309,In_1982,In_942);
and U310 (N_310,In_497,In_989);
and U311 (N_311,In_1174,In_1241);
nor U312 (N_312,In_294,In_651);
or U313 (N_313,In_978,In_1083);
or U314 (N_314,In_78,In_1975);
and U315 (N_315,In_160,In_1278);
xor U316 (N_316,In_735,In_1796);
nand U317 (N_317,In_946,In_823);
nand U318 (N_318,In_825,In_119);
nand U319 (N_319,In_887,In_1477);
nand U320 (N_320,In_650,In_579);
nor U321 (N_321,In_1831,In_230);
or U322 (N_322,In_1653,In_1605);
nor U323 (N_323,In_929,In_295);
or U324 (N_324,In_1967,In_706);
and U325 (N_325,In_102,In_1804);
nor U326 (N_326,In_1581,In_1994);
and U327 (N_327,In_111,In_1927);
nor U328 (N_328,In_1251,In_233);
and U329 (N_329,In_1093,In_280);
nand U330 (N_330,In_721,In_1493);
or U331 (N_331,In_1807,In_1533);
and U332 (N_332,In_586,In_196);
nand U333 (N_333,In_232,In_1747);
nor U334 (N_334,In_1573,In_84);
and U335 (N_335,In_1217,In_125);
nand U336 (N_336,In_1485,In_1245);
or U337 (N_337,In_701,In_1237);
nor U338 (N_338,In_386,In_1072);
nor U339 (N_339,In_1541,In_1617);
or U340 (N_340,In_905,In_746);
nor U341 (N_341,In_1007,In_1040);
nand U342 (N_342,In_380,In_1778);
nand U343 (N_343,In_1766,In_41);
nand U344 (N_344,In_571,In_1123);
nor U345 (N_345,In_908,In_1532);
nand U346 (N_346,In_215,In_1586);
nand U347 (N_347,In_559,In_708);
nor U348 (N_348,In_699,In_659);
nand U349 (N_349,In_610,In_625);
nor U350 (N_350,In_152,In_804);
or U351 (N_351,In_949,In_800);
nand U352 (N_352,In_576,In_725);
nand U353 (N_353,In_1191,In_770);
nand U354 (N_354,In_1899,In_1061);
and U355 (N_355,In_922,In_103);
nand U356 (N_356,In_1842,In_1710);
nor U357 (N_357,In_1153,In_1458);
nand U358 (N_358,In_1338,In_624);
or U359 (N_359,In_810,In_100);
or U360 (N_360,In_1909,In_310);
nand U361 (N_361,In_1274,In_760);
nand U362 (N_362,In_600,In_1971);
nor U363 (N_363,In_1658,In_1973);
or U364 (N_364,In_458,In_1959);
nor U365 (N_365,In_1111,In_1090);
nor U366 (N_366,In_1097,In_533);
nor U367 (N_367,In_425,In_1506);
nand U368 (N_368,In_118,In_959);
nor U369 (N_369,In_1887,In_379);
nand U370 (N_370,In_1370,In_1219);
and U371 (N_371,In_1001,In_413);
nor U372 (N_372,In_885,In_445);
and U373 (N_373,In_1509,In_837);
nor U374 (N_374,In_1187,In_293);
and U375 (N_375,In_665,In_1185);
nor U376 (N_376,In_1955,In_710);
and U377 (N_377,In_1320,In_1528);
nor U378 (N_378,In_503,In_1025);
and U379 (N_379,In_1084,In_335);
and U380 (N_380,In_736,In_1898);
or U381 (N_381,In_1329,In_1740);
or U382 (N_382,In_239,In_1000);
nand U383 (N_383,In_1640,In_1128);
or U384 (N_384,In_1026,In_1663);
or U385 (N_385,In_991,In_292);
and U386 (N_386,In_811,In_1662);
or U387 (N_387,In_792,In_312);
and U388 (N_388,In_1010,In_145);
nand U389 (N_389,In_1504,In_1972);
nand U390 (N_390,In_1500,In_540);
nand U391 (N_391,In_1497,In_794);
and U392 (N_392,In_839,In_1692);
and U393 (N_393,In_723,In_1498);
and U394 (N_394,In_730,In_28);
or U395 (N_395,In_812,In_1871);
nand U396 (N_396,In_1977,In_1053);
and U397 (N_397,In_1170,In_1044);
nor U398 (N_398,In_1415,In_1314);
nand U399 (N_399,In_1983,In_170);
nand U400 (N_400,In_1924,In_23);
nor U401 (N_401,In_242,In_598);
or U402 (N_402,In_1628,In_417);
or U403 (N_403,In_1754,In_1635);
or U404 (N_404,In_670,In_1694);
nand U405 (N_405,In_1718,In_1986);
nand U406 (N_406,In_489,In_1321);
and U407 (N_407,In_1920,In_741);
nor U408 (N_408,In_889,In_656);
nor U409 (N_409,In_838,In_483);
or U410 (N_410,In_113,In_945);
or U411 (N_411,In_1591,In_1136);
nand U412 (N_412,In_1429,In_1951);
nand U413 (N_413,In_1865,In_1806);
nor U414 (N_414,In_581,In_1020);
or U415 (N_415,In_1379,In_692);
or U416 (N_416,In_1828,In_1921);
nand U417 (N_417,In_1453,In_848);
nor U418 (N_418,In_139,In_153);
nor U419 (N_419,In_1987,In_1607);
nand U420 (N_420,In_1856,In_1612);
and U421 (N_421,In_448,In_1855);
and U422 (N_422,In_365,In_1362);
nand U423 (N_423,In_1690,In_602);
nor U424 (N_424,In_1537,In_748);
and U425 (N_425,In_1414,In_1089);
nand U426 (N_426,In_753,In_611);
and U427 (N_427,In_1055,In_1849);
nor U428 (N_428,In_774,In_1555);
or U429 (N_429,In_1834,In_486);
nor U430 (N_430,In_22,In_1530);
or U431 (N_431,In_1211,In_1101);
or U432 (N_432,In_866,In_346);
nor U433 (N_433,In_114,In_216);
nand U434 (N_434,In_1311,In_657);
nor U435 (N_435,In_339,In_480);
and U436 (N_436,In_234,In_387);
or U437 (N_437,In_1146,In_1216);
nand U438 (N_438,In_1845,In_1239);
and U439 (N_439,In_938,In_1812);
or U440 (N_440,In_1544,In_1928);
nand U441 (N_441,In_1830,In_1035);
or U442 (N_442,In_755,In_757);
and U443 (N_443,In_594,In_1266);
nand U444 (N_444,In_344,In_345);
and U445 (N_445,In_316,In_1460);
or U446 (N_446,In_1489,In_1656);
nor U447 (N_447,In_110,In_580);
nor U448 (N_448,In_1070,In_193);
nor U449 (N_449,In_1445,In_1711);
nor U450 (N_450,In_1182,In_367);
or U451 (N_451,In_1220,In_782);
nor U452 (N_452,In_712,In_1810);
nor U453 (N_453,In_378,In_43);
or U454 (N_454,In_482,In_861);
or U455 (N_455,In_1048,In_397);
and U456 (N_456,In_767,In_1488);
nor U457 (N_457,In_1230,In_37);
nand U458 (N_458,In_1441,In_151);
or U459 (N_459,In_709,In_282);
nand U460 (N_460,In_896,In_1028);
nand U461 (N_461,In_1150,In_9);
and U462 (N_462,In_970,In_851);
nor U463 (N_463,In_983,In_977);
nand U464 (N_464,In_833,In_101);
or U465 (N_465,In_1698,In_304);
and U466 (N_466,In_845,In_1289);
and U467 (N_467,In_971,In_1949);
or U468 (N_468,In_1273,In_19);
and U469 (N_469,In_247,In_1065);
and U470 (N_470,In_535,In_1903);
or U471 (N_471,In_74,In_1071);
or U472 (N_472,In_1880,In_524);
nor U473 (N_473,In_632,In_567);
nor U474 (N_474,In_501,In_1139);
or U475 (N_475,In_1882,In_577);
nand U476 (N_476,In_1307,In_1562);
or U477 (N_477,In_183,In_1642);
and U478 (N_478,In_1745,In_321);
and U479 (N_479,In_1615,In_772);
nand U480 (N_480,In_392,In_438);
and U481 (N_481,In_18,In_1863);
nor U482 (N_482,In_1075,In_1333);
nor U483 (N_483,In_601,In_1240);
nor U484 (N_484,In_329,In_1551);
and U485 (N_485,In_1835,In_385);
or U486 (N_486,In_227,In_337);
nor U487 (N_487,In_1715,In_1645);
or U488 (N_488,In_1945,In_875);
or U489 (N_489,In_251,In_1306);
nor U490 (N_490,In_1716,In_631);
and U491 (N_491,In_1895,In_537);
nor U492 (N_492,In_1918,In_1523);
nor U493 (N_493,In_614,In_306);
nand U494 (N_494,In_1455,In_578);
nand U495 (N_495,In_1815,In_917);
and U496 (N_496,In_1775,In_1900);
nor U497 (N_497,In_1937,In_426);
and U498 (N_498,In_1222,In_1770);
nor U499 (N_499,In_1022,In_48);
and U500 (N_500,In_473,In_876);
or U501 (N_501,In_1403,In_323);
and U502 (N_502,In_1801,In_1210);
nand U503 (N_503,In_1188,In_801);
or U504 (N_504,In_834,In_1229);
nand U505 (N_505,In_1719,In_1811);
or U506 (N_506,In_1761,In_1492);
or U507 (N_507,In_20,In_1570);
nor U508 (N_508,In_1127,In_462);
nand U509 (N_509,In_288,In_1790);
nand U510 (N_510,In_575,In_217);
and U511 (N_511,In_1588,In_381);
nor U512 (N_512,In_419,In_937);
nor U513 (N_513,In_171,In_1829);
nor U514 (N_514,In_1238,In_732);
nand U515 (N_515,In_1252,In_257);
nor U516 (N_516,In_1629,In_680);
or U517 (N_517,In_1108,In_1345);
nand U518 (N_518,In_92,In_607);
or U519 (N_519,In_1518,In_1047);
and U520 (N_520,In_1228,In_1276);
and U521 (N_521,In_168,In_1739);
nand U522 (N_522,In_1769,In_1496);
and U523 (N_523,In_1049,In_556);
or U524 (N_524,In_1505,In_1916);
nand U525 (N_525,In_542,In_1827);
and U526 (N_526,In_962,In_1857);
nor U527 (N_527,In_1361,In_1212);
or U528 (N_528,In_424,In_1077);
or U529 (N_529,In_1158,In_613);
nand U530 (N_530,In_509,In_1406);
nor U531 (N_531,In_924,In_1847);
nor U532 (N_532,In_1087,In_1202);
or U533 (N_533,In_1339,In_634);
or U534 (N_534,In_783,In_1723);
and U535 (N_535,In_349,In_1749);
or U536 (N_536,In_289,In_1482);
and U537 (N_537,In_370,In_1156);
nor U538 (N_538,In_1624,In_14);
nor U539 (N_539,In_1349,In_485);
nor U540 (N_540,In_1436,In_33);
nor U541 (N_541,In_1883,In_214);
or U542 (N_542,In_1501,In_1293);
or U543 (N_543,In_778,In_633);
nand U544 (N_544,In_1281,In_1443);
or U545 (N_545,In_1348,In_120);
nor U546 (N_546,In_713,In_1522);
and U547 (N_547,In_1332,In_25);
nand U548 (N_548,In_376,In_681);
and U549 (N_549,In_1376,In_967);
and U550 (N_550,In_891,In_878);
nand U551 (N_551,In_1450,In_1030);
nor U552 (N_552,In_1631,In_491);
nor U553 (N_553,In_1913,In_1511);
nor U554 (N_554,In_409,In_1954);
or U555 (N_555,In_131,In_1418);
nand U556 (N_556,In_1016,In_658);
nand U557 (N_557,In_797,In_1535);
or U558 (N_558,In_532,In_1648);
or U559 (N_559,In_1577,In_301);
or U560 (N_560,In_256,In_827);
nand U561 (N_561,In_29,In_862);
nor U562 (N_562,In_527,In_1813);
nor U563 (N_563,In_314,In_1465);
xnor U564 (N_564,In_1051,In_90);
and U565 (N_565,In_1371,In_1800);
nor U566 (N_566,In_56,In_628);
or U567 (N_567,In_547,In_136);
or U568 (N_568,In_951,In_1167);
or U569 (N_569,In_1784,In_1817);
nor U570 (N_570,In_313,In_198);
or U571 (N_571,In_920,In_1512);
and U572 (N_572,In_278,In_947);
nor U573 (N_573,In_1186,In_395);
and U574 (N_574,In_1319,In_819);
xor U575 (N_575,In_1448,In_1439);
and U576 (N_576,In_1494,In_817);
nand U577 (N_577,In_1560,In_939);
nor U578 (N_578,In_1606,In_1032);
nand U579 (N_579,In_146,In_969);
nand U580 (N_580,In_1080,In_1017);
nand U581 (N_581,In_83,In_793);
nand U582 (N_582,In_726,In_1837);
or U583 (N_583,In_142,In_1359);
or U584 (N_584,In_305,In_926);
or U585 (N_585,In_1405,In_1735);
nor U586 (N_586,In_1235,In_1859);
nand U587 (N_587,In_93,In_1958);
nor U588 (N_588,In_1377,In_1004);
and U589 (N_589,In_1669,In_298);
or U590 (N_590,In_165,In_1074);
and U591 (N_591,In_1152,In_1592);
nand U592 (N_592,In_122,In_284);
or U593 (N_593,In_163,In_62);
nor U594 (N_594,In_184,In_1824);
or U595 (N_595,In_868,In_1826);
or U596 (N_596,In_1929,In_172);
nand U597 (N_597,In_844,In_333);
xor U598 (N_598,In_573,In_990);
nand U599 (N_599,In_1910,In_290);
or U600 (N_600,In_1374,In_1440);
and U601 (N_601,In_1179,In_362);
nand U602 (N_602,In_1163,In_1585);
or U603 (N_603,In_1725,In_1630);
or U604 (N_604,In_919,In_846);
nand U605 (N_605,In_1764,In_1508);
nand U606 (N_606,In_240,In_974);
nand U607 (N_607,In_569,In_1981);
nand U608 (N_608,In_1935,In_955);
nor U609 (N_609,In_268,In_1721);
and U610 (N_610,In_222,In_1312);
nor U611 (N_611,In_1459,In_777);
nand U612 (N_612,In_880,In_1914);
or U613 (N_613,In_178,In_1942);
and U614 (N_614,In_1463,In_739);
and U615 (N_615,In_1233,In_1946);
nor U616 (N_616,In_1132,In_807);
nand U617 (N_617,In_1173,In_528);
nand U618 (N_618,In_789,In_654);
or U619 (N_619,In_1516,In_826);
or U620 (N_620,In_543,In_976);
or U621 (N_621,In_31,In_1121);
or U622 (N_622,In_1693,In_1943);
or U623 (N_623,In_1085,In_960);
nand U624 (N_624,In_17,In_1130);
nand U625 (N_625,In_1556,In_212);
or U626 (N_626,In_1462,In_8);
nor U627 (N_627,In_906,In_1161);
nor U628 (N_628,In_1939,In_550);
and U629 (N_629,In_1696,In_1468);
or U630 (N_630,In_1666,In_1479);
nand U631 (N_631,In_1088,In_1904);
nor U632 (N_632,In_707,In_415);
nor U633 (N_633,In_1795,In_179);
xnor U634 (N_634,In_1124,In_1893);
nor U635 (N_635,In_1520,In_10);
or U636 (N_636,In_1751,In_1253);
or U637 (N_637,In_1114,In_830);
or U638 (N_638,In_1779,In_915);
and U639 (N_639,In_822,In_272);
or U640 (N_640,In_1767,In_617);
xnor U641 (N_641,In_816,In_874);
or U642 (N_642,In_137,In_446);
nand U643 (N_643,In_911,In_1853);
or U644 (N_644,In_1165,In_1765);
nor U645 (N_645,In_737,In_207);
nor U646 (N_646,In_883,In_647);
nand U647 (N_647,In_42,In_1680);
nor U648 (N_648,In_1234,In_869);
nor U649 (N_649,In_1100,In_1380);
nor U650 (N_650,In_743,In_265);
nand U651 (N_651,In_641,In_592);
nand U652 (N_652,In_1664,In_177);
or U653 (N_653,In_348,In_719);
and U654 (N_654,In_913,In_1787);
or U655 (N_655,In_60,In_1305);
and U656 (N_656,In_58,In_1874);
nand U657 (N_657,In_200,In_1947);
or U658 (N_658,In_1316,In_1484);
or U659 (N_659,In_1938,In_1470);
or U660 (N_660,In_1176,In_529);
or U661 (N_661,In_1545,In_1797);
or U662 (N_662,In_490,In_195);
and U663 (N_663,In_1059,In_1148);
nor U664 (N_664,In_1155,In_1402);
and U665 (N_665,In_769,In_1571);
nand U666 (N_666,In_1722,In_843);
or U667 (N_667,In_935,In_429);
and U668 (N_668,In_1336,In_454);
nand U669 (N_669,In_881,In_805);
or U670 (N_670,In_261,In_1864);
or U671 (N_671,In_143,In_81);
or U672 (N_672,In_1786,In_1978);
nand U673 (N_673,In_965,In_1438);
nand U674 (N_674,In_3,In_1681);
or U675 (N_675,In_297,In_1037);
and U676 (N_676,In_194,In_1432);
nor U677 (N_677,In_1941,In_1444);
nand U678 (N_678,In_1992,In_1034);
and U679 (N_679,In_1280,In_1660);
and U680 (N_680,In_327,In_1154);
and U681 (N_681,In_161,In_1260);
nand U682 (N_682,In_384,In_1634);
and U683 (N_683,In_1326,In_1980);
or U684 (N_684,In_1671,In_1644);
and U685 (N_685,In_511,In_1944);
and U686 (N_686,In_541,In_1809);
and U687 (N_687,In_544,In_1486);
and U688 (N_688,In_36,In_729);
and U689 (N_689,In_1099,In_518);
or U690 (N_690,In_629,In_1015);
nand U691 (N_691,In_1846,In_809);
and U692 (N_692,In_369,In_1613);
and U693 (N_693,In_116,In_1286);
or U694 (N_694,In_1137,In_609);
nand U695 (N_695,In_1029,In_813);
nand U696 (N_696,In_134,In_1677);
nand U697 (N_697,In_1502,In_416);
nand U698 (N_698,In_1081,In_1340);
or U699 (N_699,In_588,In_1451);
nand U700 (N_700,In_1038,In_599);
xnor U701 (N_701,In_583,In_442);
nand U702 (N_702,In_342,In_1393);
and U703 (N_703,In_1355,In_1062);
nand U704 (N_704,In_157,In_1327);
nand U705 (N_705,In_564,In_1277);
and U706 (N_706,In_1365,In_852);
and U707 (N_707,In_1595,In_1991);
nand U708 (N_708,In_909,In_1572);
nand U709 (N_709,In_912,In_391);
and U710 (N_710,In_1862,In_34);
or U711 (N_711,In_1082,In_1673);
or U712 (N_712,In_1073,In_7);
nor U713 (N_713,In_854,In_1999);
nor U714 (N_714,In_1609,In_174);
and U715 (N_715,In_1743,In_358);
nor U716 (N_716,In_1428,In_1416);
or U717 (N_717,In_994,In_1707);
and U718 (N_718,In_1936,In_950);
nand U719 (N_719,In_521,In_478);
or U720 (N_720,In_286,In_1318);
nand U721 (N_721,In_745,In_456);
and U722 (N_722,In_1788,In_850);
or U723 (N_723,In_984,In_870);
or U724 (N_724,In_790,In_266);
and U725 (N_725,In_853,In_246);
or U726 (N_726,In_1687,In_773);
or U727 (N_727,In_1177,In_1891);
nor U728 (N_728,In_1144,In_267);
and U729 (N_729,In_1358,In_1584);
and U730 (N_730,In_115,In_930);
and U731 (N_731,In_1086,In_894);
and U732 (N_732,In_1421,In_1019);
nand U733 (N_733,In_1890,In_467);
nor U734 (N_734,In_175,In_907);
nor U735 (N_735,In_1599,In_1298);
and U736 (N_736,In_474,In_791);
and U737 (N_737,In_1023,In_1667);
or U738 (N_738,In_431,In_1651);
or U739 (N_739,In_893,In_363);
nor U740 (N_740,In_1356,In_1712);
and U741 (N_741,In_1147,In_1683);
nand U742 (N_742,In_1665,In_176);
nand U743 (N_743,In_1608,In_1346);
or U744 (N_744,In_1833,In_1799);
or U745 (N_745,In_1534,In_436);
nor U746 (N_746,In_856,In_123);
nor U747 (N_747,In_259,In_649);
nor U748 (N_748,In_1655,In_517);
nand U749 (N_749,In_1413,In_1884);
nand U750 (N_750,In_1096,In_1419);
nor U751 (N_751,In_1932,In_273);
nor U752 (N_752,In_502,In_393);
nor U753 (N_753,In_516,In_324);
nand U754 (N_754,In_1209,In_623);
or U755 (N_755,In_154,In_525);
or U756 (N_756,In_1792,In_1151);
nor U757 (N_757,In_133,In_451);
and U758 (N_758,In_1720,In_666);
and U759 (N_759,In_1691,In_1744);
nor U760 (N_760,In_1611,In_1729);
nor U761 (N_761,In_331,In_283);
nor U762 (N_762,In_806,In_1524);
nand U763 (N_763,In_1372,In_1122);
nand U764 (N_764,In_953,In_1394);
nor U765 (N_765,In_1198,In_1679);
xnor U766 (N_766,In_1875,In_377);
nor U767 (N_767,In_1843,In_276);
nor U768 (N_768,In_1583,In_855);
nand U769 (N_769,In_1381,In_682);
nor U770 (N_770,In_742,In_1271);
and U771 (N_771,In_420,In_548);
nand U772 (N_772,In_630,In_1449);
and U773 (N_773,In_5,In_1256);
and U774 (N_774,In_683,In_203);
or U775 (N_775,In_1342,In_1548);
or U776 (N_776,In_763,In_423);
and U777 (N_777,In_229,In_1748);
or U778 (N_778,In_1990,In_675);
or U779 (N_779,In_1115,In_892);
nor U780 (N_780,In_1619,In_1869);
and U781 (N_781,In_1730,In_1213);
and U782 (N_782,In_209,In_1601);
nor U783 (N_783,In_371,In_433);
and U784 (N_784,In_948,In_733);
or U785 (N_785,In_899,In_1033);
nor U786 (N_786,In_1224,In_1503);
nor U787 (N_787,In_674,In_1621);
and U788 (N_788,In_504,In_1250);
and U789 (N_789,In_399,In_720);
nor U790 (N_790,In_1563,In_1078);
or U791 (N_791,In_320,In_277);
nor U792 (N_792,In_1423,In_1894);
and U793 (N_793,In_98,In_872);
xor U794 (N_794,In_336,In_604);
and U795 (N_795,In_1360,In_201);
and U796 (N_796,In_646,In_1408);
or U797 (N_797,In_534,In_1475);
or U798 (N_798,In_44,In_24);
nor U799 (N_799,In_765,In_236);
nor U800 (N_800,In_842,N_400);
nor U801 (N_801,N_182,In_1011);
or U802 (N_802,N_242,N_627);
nand U803 (N_803,N_693,N_234);
nand U804 (N_804,N_56,N_426);
nor U805 (N_805,N_480,N_433);
nand U806 (N_806,In_1420,N_377);
and U807 (N_807,In_1288,In_1366);
nand U808 (N_808,N_456,N_449);
and U809 (N_809,N_227,In_1268);
or U810 (N_810,N_363,N_707);
nand U811 (N_811,N_745,N_429);
and U812 (N_812,N_76,In_902);
nor U813 (N_813,N_442,In_1157);
and U814 (N_814,N_639,N_121);
or U815 (N_815,In_91,N_628);
or U816 (N_816,N_616,In_1267);
and U817 (N_817,N_41,In_832);
or U818 (N_818,N_215,N_501);
or U819 (N_819,In_1931,N_83);
and U820 (N_820,N_686,N_372);
nor U821 (N_821,In_1375,N_589);
nand U822 (N_822,N_719,N_103);
or U823 (N_823,In_941,N_385);
or U824 (N_824,In_1218,N_559);
and U825 (N_825,N_416,In_1600);
or U826 (N_826,N_411,N_669);
nand U827 (N_827,N_713,In_1270);
or U828 (N_828,In_68,N_166);
and U829 (N_829,N_58,In_644);
and U830 (N_830,N_419,In_840);
or U831 (N_831,N_792,In_494);
or U832 (N_832,In_435,In_1553);
and U833 (N_833,N_785,In_150);
nor U834 (N_834,In_903,N_394);
nor U835 (N_835,N_648,In_447);
and U836 (N_836,In_126,N_356);
nor U837 (N_837,In_526,N_514);
nor U838 (N_838,In_1672,N_410);
nand U839 (N_839,N_632,In_1140);
nand U840 (N_840,In_158,N_663);
nand U841 (N_841,In_1027,N_647);
nor U842 (N_842,In_1752,N_551);
nand U843 (N_843,N_5,In_356);
nand U844 (N_844,In_995,N_232);
or U845 (N_845,N_233,N_230);
and U846 (N_846,N_642,In_1542);
nand U847 (N_847,N_269,In_1633);
or U848 (N_848,N_760,In_1701);
and U849 (N_849,In_372,N_577);
nand U850 (N_850,N_478,In_560);
nand U851 (N_851,In_1284,In_1395);
or U852 (N_852,N_343,N_683);
nand U853 (N_853,N_448,In_1819);
nand U854 (N_854,In_1452,N_615);
nand U855 (N_855,N_523,N_63);
nor U856 (N_856,In_612,N_398);
and U857 (N_857,In_963,In_357);
or U858 (N_858,N_279,N_2);
nand U859 (N_859,N_518,In_1129);
nand U860 (N_860,N_475,In_1821);
nand U861 (N_861,N_240,N_705);
and U862 (N_862,N_596,In_1625);
nor U863 (N_863,In_1299,N_178);
nor U864 (N_864,N_765,In_1623);
nand U865 (N_865,N_754,In_1283);
nand U866 (N_866,In_877,N_625);
nand U867 (N_867,In_779,N_689);
nand U868 (N_868,N_111,N_147);
and U869 (N_869,N_203,In_1309);
nand U870 (N_870,In_1750,N_365);
nand U871 (N_871,In_1823,N_72);
nand U872 (N_872,In_453,N_132);
nand U873 (N_873,In_704,N_584);
or U874 (N_874,In_1105,N_135);
nor U875 (N_875,N_560,N_297);
and U876 (N_876,N_374,N_31);
nor U877 (N_877,N_352,N_702);
or U878 (N_878,N_773,In_999);
xor U879 (N_879,N_23,In_1728);
nor U880 (N_880,N_751,In_249);
or U881 (N_881,N_198,In_956);
and U882 (N_882,N_487,In_1208);
and U883 (N_883,In_1181,N_220);
nand U884 (N_884,In_714,N_688);
xnor U885 (N_885,N_414,In_1351);
or U886 (N_886,In_1521,N_318);
nand U887 (N_887,N_600,N_154);
nand U888 (N_888,In_1647,N_299);
nand U889 (N_889,N_25,In_1135);
and U890 (N_890,N_316,N_355);
and U891 (N_891,In_49,In_1793);
nand U892 (N_892,N_503,N_432);
nand U893 (N_893,N_392,N_353);
nor U894 (N_894,In_219,N_703);
and U895 (N_895,N_753,In_243);
nor U896 (N_896,N_461,In_1295);
and U897 (N_897,In_1626,N_425);
or U898 (N_898,In_1113,N_155);
or U899 (N_899,N_793,N_573);
and U900 (N_900,In_1310,N_443);
nand U901 (N_901,N_264,In_258);
or U902 (N_902,N_77,In_471);
and U903 (N_903,N_27,N_435);
or U904 (N_904,In_690,N_60);
nor U905 (N_905,In_1194,N_75);
or U906 (N_906,In_228,N_641);
nor U907 (N_907,N_114,In_1003);
or U908 (N_908,In_255,In_1226);
nand U909 (N_909,In_1968,N_629);
nor U910 (N_910,N_38,N_303);
and U911 (N_911,N_160,In_487);
nand U912 (N_912,N_464,N_212);
and U913 (N_913,In_1771,N_52);
or U914 (N_914,In_1974,N_181);
nor U915 (N_915,N_491,N_507);
or U916 (N_916,In_437,N_43);
nor U917 (N_917,N_515,N_534);
or U918 (N_918,N_321,N_752);
and U919 (N_919,In_135,N_659);
nand U920 (N_920,N_750,N_192);
nor U921 (N_921,N_128,N_152);
and U922 (N_922,N_367,N_45);
or U923 (N_923,In_1404,N_228);
nand U924 (N_924,N_797,In_1315);
nor U925 (N_925,N_668,N_149);
nor U926 (N_926,N_309,N_253);
nor U927 (N_927,In_568,N_384);
nor U928 (N_928,In_1839,N_36);
or U929 (N_929,In_818,N_766);
nand U930 (N_930,N_106,N_117);
or U931 (N_931,In_1487,N_404);
nand U932 (N_932,In_1996,N_509);
nand U933 (N_933,N_272,N_273);
and U934 (N_934,In_616,N_500);
and U935 (N_935,In_515,In_1794);
nand U936 (N_936,In_140,In_1639);
and U937 (N_937,N_210,In_1618);
nand U938 (N_938,In_1410,N_180);
or U939 (N_939,N_772,In_220);
nand U940 (N_940,In_428,In_1430);
nor U941 (N_941,N_477,N_499);
nand U942 (N_942,In_1926,N_183);
and U943 (N_943,N_33,N_555);
or U944 (N_944,N_248,N_0);
and U945 (N_945,N_331,N_65);
or U946 (N_946,In_1303,N_50);
nand U947 (N_947,In_1906,N_73);
or U948 (N_948,N_603,In_1052);
or U949 (N_949,N_423,In_1013);
and U950 (N_950,In_964,In_383);
or U951 (N_951,N_214,N_34);
nor U952 (N_952,N_281,N_189);
nor U953 (N_953,In_1495,N_93);
nand U954 (N_954,N_175,In_472);
nor U955 (N_955,In_828,In_1676);
nor U956 (N_956,N_452,N_366);
or U957 (N_957,N_657,N_554);
or U958 (N_958,N_579,N_782);
or U959 (N_959,N_126,In_1603);
and U960 (N_960,In_781,N_7);
nor U961 (N_961,In_1323,N_631);
nor U962 (N_962,In_1225,N_148);
and U963 (N_963,N_723,N_85);
and U964 (N_964,N_422,In_364);
nor U965 (N_965,N_612,In_1352);
nand U966 (N_966,N_597,In_606);
or U967 (N_967,N_728,N_125);
and U968 (N_968,N_424,In_375);
nand U969 (N_969,In_1389,N_241);
or U970 (N_970,N_505,N_88);
or U971 (N_971,N_67,N_326);
and U972 (N_972,N_150,N_661);
nand U973 (N_973,N_474,N_9);
nor U974 (N_974,N_665,N_357);
nand U975 (N_975,N_613,In_296);
nor U976 (N_976,In_587,N_174);
and U977 (N_977,In_271,N_493);
nor U978 (N_978,In_1382,N_4);
or U979 (N_979,N_379,In_1390);
and U980 (N_980,N_463,N_346);
nand U981 (N_981,N_796,N_580);
and U982 (N_982,N_525,In_1515);
nor U983 (N_983,In_549,N_569);
nor U984 (N_984,N_345,In_1297);
nor U985 (N_985,N_789,N_566);
or U986 (N_986,In_1567,N_739);
nand U987 (N_987,N_136,N_710);
nand U988 (N_988,N_725,N_53);
and U989 (N_989,In_1896,In_1808);
nor U990 (N_990,N_497,N_610);
nor U991 (N_991,N_614,In_50);
or U992 (N_992,N_471,In_1435);
or U993 (N_993,N_335,N_138);
nand U994 (N_994,N_49,N_3);
and U995 (N_995,N_396,In_1820);
nand U996 (N_996,N_90,In_421);
nand U997 (N_997,In_94,N_70);
nor U998 (N_998,N_516,N_364);
or U999 (N_999,In_921,N_706);
nand U1000 (N_1000,N_284,In_695);
nand U1001 (N_1001,N_320,N_323);
nor U1002 (N_1002,In_457,In_1491);
nand U1003 (N_1003,N_687,In_566);
and U1004 (N_1004,N_635,N_609);
nor U1005 (N_1005,In_968,N_71);
nor U1006 (N_1006,N_791,In_1940);
nand U1007 (N_1007,N_245,N_222);
or U1008 (N_1008,N_113,In_191);
and U1009 (N_1009,N_735,N_64);
nand U1010 (N_1010,N_296,In_1540);
and U1011 (N_1011,N_328,In_694);
and U1012 (N_1012,N_496,N_225);
xnor U1013 (N_1013,In_1889,N_542);
nor U1014 (N_1014,N_768,N_709);
nor U1015 (N_1015,In_1367,In_441);
or U1016 (N_1016,In_1574,N_406);
and U1017 (N_1017,N_644,N_172);
and U1018 (N_1018,N_537,N_221);
and U1019 (N_1019,N_651,N_605);
nor U1020 (N_1020,N_213,N_165);
or U1021 (N_1021,In_1112,N_92);
nand U1022 (N_1022,N_684,N_412);
nor U1023 (N_1023,N_764,In_374);
nand U1024 (N_1024,N_418,N_124);
or U1025 (N_1025,In_16,In_1756);
nand U1026 (N_1026,In_1290,N_193);
or U1027 (N_1027,In_972,N_185);
and U1028 (N_1028,N_672,N_666);
and U1029 (N_1029,N_571,N_337);
or U1030 (N_1030,N_62,N_604);
and U1031 (N_1031,N_15,N_660);
and U1032 (N_1032,N_322,In_1425);
and U1033 (N_1033,N_680,N_633);
nand U1034 (N_1034,N_485,N_311);
and U1035 (N_1035,In_250,N_94);
or U1036 (N_1036,N_96,In_703);
and U1037 (N_1037,In_1575,N_658);
or U1038 (N_1038,In_1275,N_390);
or U1039 (N_1039,N_305,N_417);
and U1040 (N_1040,N_712,In_53);
and U1041 (N_1041,N_716,N_697);
nor U1042 (N_1042,N_54,N_506);
or U1043 (N_1043,In_127,N_585);
nand U1044 (N_1044,In_561,In_452);
and U1045 (N_1045,In_87,N_759);
or U1046 (N_1046,In_1042,In_182);
and U1047 (N_1047,N_558,N_774);
or U1048 (N_1048,N_591,N_109);
and U1049 (N_1049,N_531,In_238);
nor U1050 (N_1050,N_698,N_388);
and U1051 (N_1051,N_86,In_1901);
or U1052 (N_1052,N_209,In_1597);
and U1053 (N_1053,N_158,In_1472);
nor U1054 (N_1054,N_347,In_366);
or U1055 (N_1055,In_450,N_79);
or U1056 (N_1056,N_599,In_40);
nand U1057 (N_1057,N_142,In_1422);
or U1058 (N_1058,N_157,N_671);
nor U1059 (N_1059,In_80,N_622);
nand U1060 (N_1060,N_511,N_287);
and U1061 (N_1061,N_324,In_648);
or U1062 (N_1062,N_675,N_139);
nand U1063 (N_1063,In_664,N_14);
nand U1064 (N_1064,N_80,N_116);
or U1065 (N_1065,N_790,N_386);
or U1066 (N_1066,N_229,In_224);
nand U1067 (N_1067,In_1885,N_696);
or U1068 (N_1068,N_420,N_586);
nand U1069 (N_1069,In_785,N_315);
xnor U1070 (N_1070,In_928,N_389);
and U1071 (N_1071,N_202,N_69);
nor U1072 (N_1072,N_482,N_301);
or U1073 (N_1073,In_1682,N_489);
nand U1074 (N_1074,In_1396,N_244);
nand U1075 (N_1075,In_1713,N_459);
and U1076 (N_1076,In_1334,In_931);
nand U1077 (N_1077,In_1984,In_1689);
and U1078 (N_1078,In_1930,In_1480);
nand U1079 (N_1079,N_761,In_1009);
and U1080 (N_1080,N_513,N_163);
nand U1081 (N_1081,N_434,N_21);
nor U1082 (N_1082,In_768,N_749);
nand U1083 (N_1083,N_673,N_349);
and U1084 (N_1084,N_486,In_1296);
nor U1085 (N_1085,N_624,N_206);
nor U1086 (N_1086,N_360,N_397);
xor U1087 (N_1087,N_617,N_446);
nand U1088 (N_1088,In_1201,In_1708);
nand U1089 (N_1089,In_1060,N_99);
xnor U1090 (N_1090,N_718,N_217);
nor U1091 (N_1091,N_317,N_526);
and U1092 (N_1092,N_159,In_1514);
nor U1093 (N_1093,N_611,N_137);
nand U1094 (N_1094,N_767,In_1369);
nand U1095 (N_1095,N_522,N_29);
and U1096 (N_1096,N_46,N_8);
and U1097 (N_1097,In_857,N_451);
nand U1098 (N_1098,In_1407,N_237);
nand U1099 (N_1099,In_166,N_304);
nand U1100 (N_1100,In_884,In_1031);
nor U1101 (N_1101,N_747,In_1962);
and U1102 (N_1102,In_1473,In_1347);
nand U1103 (N_1103,N_179,N_556);
and U1104 (N_1104,N_19,N_572);
or U1105 (N_1105,N_574,In_1602);
nor U1106 (N_1106,N_415,N_219);
nand U1107 (N_1107,N_112,N_350);
nor U1108 (N_1108,N_484,N_286);
nand U1109 (N_1109,In_132,In_443);
nand U1110 (N_1110,N_757,N_643);
or U1111 (N_1111,In_408,N_543);
and U1112 (N_1112,N_325,N_775);
nor U1113 (N_1113,In_1724,N_607);
or U1114 (N_1114,In_404,N_494);
nor U1115 (N_1115,N_717,N_595);
xor U1116 (N_1116,N_495,N_457);
nor U1117 (N_1117,N_151,In_584);
nand U1118 (N_1118,N_441,In_63);
and U1119 (N_1119,N_24,In_440);
nand U1120 (N_1120,N_378,N_164);
and U1121 (N_1121,In_1221,N_582);
or U1122 (N_1122,N_568,N_87);
or U1123 (N_1123,N_359,N_679);
and U1124 (N_1124,N_521,In_73);
nand U1125 (N_1125,N_28,N_294);
or U1126 (N_1126,In_403,In_860);
or U1127 (N_1127,N_722,N_330);
and U1128 (N_1128,N_280,N_447);
and U1129 (N_1129,N_257,N_578);
nand U1130 (N_1130,In_1387,N_567);
nor U1131 (N_1131,In_740,N_621);
or U1132 (N_1132,N_479,N_541);
or U1133 (N_1133,N_454,N_236);
nor U1134 (N_1134,N_650,N_699);
nand U1135 (N_1135,N_786,In_961);
and U1136 (N_1136,N_78,N_517);
nor U1137 (N_1137,N_382,In_1733);
nor U1138 (N_1138,N_146,In_47);
nor U1139 (N_1139,N_141,N_342);
or U1140 (N_1140,N_780,In_1200);
nor U1141 (N_1141,N_387,In_1141);
or U1142 (N_1142,N_430,N_308);
nand U1143 (N_1143,In_427,N_667);
and U1144 (N_1144,N_289,In_673);
nor U1145 (N_1145,N_348,N_61);
and U1146 (N_1146,N_646,N_312);
or U1147 (N_1147,N_168,In_1203);
nor U1148 (N_1148,In_1604,N_730);
or U1149 (N_1149,N_226,In_1469);
nand U1150 (N_1150,In_1067,N_598);
nor U1151 (N_1151,In_340,N_467);
or U1152 (N_1152,In_1242,In_849);
and U1153 (N_1153,N_314,In_918);
or U1154 (N_1154,N_207,N_602);
or U1155 (N_1155,N_381,N_205);
nor U1156 (N_1156,In_418,N_338);
or U1157 (N_1157,In_1706,N_30);
nand U1158 (N_1158,N_562,In_185);
and U1159 (N_1159,In_1166,N_736);
and U1160 (N_1160,In_226,In_688);
or U1161 (N_1161,N_153,N_275);
nand U1162 (N_1162,In_430,In_1180);
or U1163 (N_1163,N_191,N_781);
nand U1164 (N_1164,In_788,N_721);
or U1165 (N_1165,N_188,N_436);
nor U1166 (N_1166,N_536,In_269);
and U1167 (N_1167,N_57,N_84);
and U1168 (N_1168,In_1953,N_177);
nor U1169 (N_1169,N_469,In_944);
and U1170 (N_1170,N_670,N_134);
and U1171 (N_1171,In_1881,N_654);
and U1172 (N_1172,N_700,N_504);
nand U1173 (N_1173,N_40,In_1079);
nor U1174 (N_1174,N_340,N_535);
nand U1175 (N_1175,N_89,N_795);
nor U1176 (N_1176,In_1258,In_1373);
nor U1177 (N_1177,In_796,In_1627);
nor U1178 (N_1178,N_545,In_107);
or U1179 (N_1179,N_630,In_873);
nand U1180 (N_1180,In_187,N_714);
nand U1181 (N_1181,In_141,N_450);
nand U1182 (N_1182,N_251,N_254);
nor U1183 (N_1183,In_105,N_738);
nand U1184 (N_1184,N_618,N_742);
nand U1185 (N_1185,N_208,N_199);
nand U1186 (N_1186,N_100,N_677);
or U1187 (N_1187,In_1598,In_401);
and U1188 (N_1188,N_211,N_727);
nor U1189 (N_1189,N_373,N_375);
nand U1190 (N_1190,In_479,N_231);
or U1191 (N_1191,N_488,N_37);
nor U1192 (N_1192,N_519,N_55);
nor U1193 (N_1193,N_262,In_235);
and U1194 (N_1194,In_522,N_553);
and U1195 (N_1195,N_319,N_402);
nor U1196 (N_1196,In_1164,In_1357);
and U1197 (N_1197,N_341,N_502);
nand U1198 (N_1198,N_458,N_581);
and U1199 (N_1199,N_235,N_238);
and U1200 (N_1200,N_468,N_549);
and U1201 (N_1201,In_1178,N_770);
or U1202 (N_1202,N_409,N_313);
nor U1203 (N_1203,In_1685,In_1519);
nand U1204 (N_1204,N_144,N_729);
nand U1205 (N_1205,In_808,N_476);
nand U1206 (N_1206,In_459,In_1045);
nand U1207 (N_1207,N_20,N_408);
and U1208 (N_1208,N_249,N_288);
or U1209 (N_1209,N_35,N_763);
or U1210 (N_1210,In_405,In_1989);
and U1211 (N_1211,N_776,N_133);
and U1212 (N_1212,In_985,N_498);
nor U1213 (N_1213,In_1726,N_17);
nor U1214 (N_1214,In_1247,N_354);
and U1215 (N_1215,In_1192,N_265);
nor U1216 (N_1216,N_285,N_561);
and U1217 (N_1217,N_362,N_255);
and U1218 (N_1218,N_638,N_704);
nand U1219 (N_1219,N_266,N_779);
and U1220 (N_1220,N_274,N_590);
nor U1221 (N_1221,In_1363,N_395);
nand U1222 (N_1222,N_748,In_888);
nand U1223 (N_1223,N_652,In_1118);
nor U1224 (N_1224,In_1661,N_97);
and U1225 (N_1225,N_293,N_246);
and U1226 (N_1226,N_583,N_102);
nand U1227 (N_1227,N_784,N_681);
or U1228 (N_1228,N_161,N_186);
nor U1229 (N_1229,N_104,In_155);
nor U1230 (N_1230,In_565,N_156);
nor U1231 (N_1231,N_200,N_427);
or U1232 (N_1232,N_606,N_115);
and U1233 (N_1233,N_122,N_737);
nand U1234 (N_1234,N_428,N_762);
and U1235 (N_1235,N_740,In_1709);
nand U1236 (N_1236,N_548,In_1561);
nor U1237 (N_1237,N_358,N_576);
nor U1238 (N_1238,N_176,In_1727);
xnor U1239 (N_1239,N_334,In_639);
nor U1240 (N_1240,N_758,N_532);
or U1241 (N_1241,N_587,N_247);
and U1242 (N_1242,N_119,N_798);
or U1243 (N_1243,N_259,In_46);
nor U1244 (N_1244,In_627,In_1104);
nand U1245 (N_1245,In_1897,N_720);
nor U1246 (N_1246,N_570,N_118);
and U1247 (N_1247,N_290,N_508);
or U1248 (N_1248,N_101,N_656);
nand U1249 (N_1249,In_1195,N_626);
nor U1250 (N_1250,N_544,N_530);
and U1251 (N_1251,N_339,In_795);
and U1252 (N_1252,N_283,N_620);
nor U1253 (N_1253,In_1576,In_1737);
or U1254 (N_1254,N_510,In_750);
and U1255 (N_1255,N_74,N_190);
nand U1256 (N_1256,N_66,N_540);
nand U1257 (N_1257,In_1054,In_1483);
or U1258 (N_1258,N_300,In_1190);
or U1259 (N_1259,In_1008,N_302);
or U1260 (N_1260,N_171,N_130);
or U1261 (N_1261,N_268,In_661);
nor U1262 (N_1262,In_1461,N_42);
nand U1263 (N_1263,In_1844,N_11);
nor U1264 (N_1264,N_685,In_1742);
and U1265 (N_1265,In_463,N_250);
or U1266 (N_1266,In_936,N_593);
and U1267 (N_1267,In_671,N_1);
nand U1268 (N_1268,N_440,N_676);
nor U1269 (N_1269,N_143,N_258);
or U1270 (N_1270,N_108,N_370);
xor U1271 (N_1271,N_39,In_1579);
and U1272 (N_1272,N_295,N_204);
or U1273 (N_1273,N_407,In_237);
nor U1274 (N_1274,In_1162,N_129);
and U1275 (N_1275,N_623,N_369);
or U1276 (N_1276,In_99,N_755);
or U1277 (N_1277,N_557,In_1261);
nand U1278 (N_1278,N_298,In_353);
nand U1279 (N_1279,N_473,N_453);
and U1280 (N_1280,N_674,N_276);
nand U1281 (N_1281,In_776,N_462);
nand U1282 (N_1282,In_1385,N_327);
nor U1283 (N_1283,N_383,N_197);
or U1284 (N_1284,N_405,In_835);
and U1285 (N_1285,In_1107,In_1189);
and U1286 (N_1286,N_131,N_371);
nand U1287 (N_1287,N_524,N_184);
and U1288 (N_1288,In_1547,In_1637);
nand U1289 (N_1289,N_120,In_77);
and U1290 (N_1290,N_634,N_282);
nor U1291 (N_1291,N_399,N_533);
and U1292 (N_1292,N_731,N_445);
or U1293 (N_1293,N_48,N_734);
and U1294 (N_1294,In_1456,In_45);
or U1295 (N_1295,In_1589,N_145);
or U1296 (N_1296,N_472,N_10);
nand U1297 (N_1297,In_689,N_361);
and U1298 (N_1298,In_562,N_439);
and U1299 (N_1299,N_655,N_6);
nor U1300 (N_1300,N_563,N_547);
nor U1301 (N_1301,N_744,N_592);
or U1302 (N_1302,N_59,N_756);
and U1303 (N_1303,N_12,In_270);
or U1304 (N_1304,In_1641,N_292);
or U1305 (N_1305,N_82,N_195);
nor U1306 (N_1306,N_194,N_601);
nand U1307 (N_1307,In_1734,In_328);
and U1308 (N_1308,In_1354,In_655);
nand U1309 (N_1309,N_787,N_243);
or U1310 (N_1310,N_575,In_495);
nand U1311 (N_1311,In_484,N_81);
nor U1312 (N_1312,In_1525,In_308);
nor U1313 (N_1313,N_277,N_788);
or U1314 (N_1314,N_636,In_1732);
nand U1315 (N_1315,N_127,In_210);
nand U1316 (N_1316,N_527,N_216);
or U1317 (N_1317,N_169,N_403);
and U1318 (N_1318,N_701,N_538);
or U1319 (N_1319,N_380,N_187);
or U1320 (N_1320,N_391,N_649);
and U1321 (N_1321,In_1780,N_490);
nor U1322 (N_1322,In_1364,N_260);
nand U1323 (N_1323,N_98,N_546);
and U1324 (N_1324,N_694,In_677);
and U1325 (N_1325,In_981,In_1012);
nor U1326 (N_1326,N_162,N_695);
nor U1327 (N_1327,In_620,N_329);
nor U1328 (N_1328,In_1950,N_691);
nor U1329 (N_1329,In_1409,In_554);
nor U1330 (N_1330,N_771,N_170);
nand U1331 (N_1331,N_743,N_267);
nor U1332 (N_1332,In_744,In_1803);
nor U1333 (N_1333,In_663,N_732);
and U1334 (N_1334,N_270,N_173);
and U1335 (N_1335,In_13,N_51);
or U1336 (N_1336,N_550,N_271);
and U1337 (N_1337,N_528,N_307);
nand U1338 (N_1338,N_107,In_898);
or U1339 (N_1339,N_336,N_783);
and U1340 (N_1340,In_291,N_466);
nand U1341 (N_1341,N_47,N_645);
or U1342 (N_1342,N_95,N_692);
nor U1343 (N_1343,N_741,N_44);
or U1344 (N_1344,N_291,N_637);
or U1345 (N_1345,N_91,N_22);
nand U1346 (N_1346,N_746,N_252);
nand U1347 (N_1347,N_196,N_110);
nand U1348 (N_1348,In_352,N_263);
and U1349 (N_1349,N_438,In_685);
and U1350 (N_1350,N_778,In_1292);
or U1351 (N_1351,N_708,N_393);
or U1352 (N_1352,In_1291,In_952);
nand U1353 (N_1353,In_1397,N_18);
nor U1354 (N_1354,In_1854,N_455);
nor U1355 (N_1355,N_711,In_315);
or U1356 (N_1356,N_769,N_565);
or U1357 (N_1357,In_1850,N_678);
or U1358 (N_1358,N_218,N_224);
nor U1359 (N_1359,In_711,N_653);
and U1360 (N_1360,In_1590,In_1262);
nor U1361 (N_1361,In_608,N_351);
nor U1362 (N_1362,N_588,N_794);
nor U1363 (N_1363,N_32,N_256);
xnor U1364 (N_1364,N_470,N_690);
or U1365 (N_1365,N_777,N_401);
nor U1366 (N_1366,In_619,In_1457);
and U1367 (N_1367,N_552,N_421);
or U1368 (N_1368,In_1143,N_465);
nand U1369 (N_1369,N_140,In_1988);
and U1370 (N_1370,N_68,N_512);
or U1371 (N_1371,N_460,N_492);
nand U1372 (N_1372,In_449,In_72);
and U1373 (N_1373,N_13,N_368);
xor U1374 (N_1374,N_239,N_594);
and U1375 (N_1375,In_766,N_664);
or U1376 (N_1376,In_1746,N_123);
nand U1377 (N_1377,N_306,N_799);
nand U1378 (N_1378,In_1117,N_437);
and U1379 (N_1379,N_724,N_444);
nor U1380 (N_1380,N_167,N_333);
or U1381 (N_1381,N_619,N_529);
nor U1382 (N_1382,N_520,In_1447);
nor U1383 (N_1383,In_558,N_481);
nor U1384 (N_1384,N_105,N_483);
nand U1385 (N_1385,In_1317,N_223);
and U1386 (N_1386,N_310,N_715);
nand U1387 (N_1387,N_344,N_201);
or U1388 (N_1388,In_696,N_662);
nor U1389 (N_1389,In_1908,N_413);
nand U1390 (N_1390,N_431,N_726);
nor U1391 (N_1391,N_682,In_1231);
nand U1392 (N_1392,In_1963,In_252);
nor U1393 (N_1393,N_16,In_434);
and U1394 (N_1394,N_26,N_278);
nand U1395 (N_1395,N_376,N_539);
or U1396 (N_1396,N_733,In_882);
nand U1397 (N_1397,N_608,N_261);
xor U1398 (N_1398,N_640,N_332);
nand U1399 (N_1399,N_564,In_1517);
or U1400 (N_1400,N_663,In_1457);
or U1401 (N_1401,In_981,In_449);
and U1402 (N_1402,N_134,N_761);
or U1403 (N_1403,In_1221,In_1190);
nand U1404 (N_1404,N_367,N_55);
or U1405 (N_1405,N_382,N_287);
nor U1406 (N_1406,N_497,N_447);
nand U1407 (N_1407,In_1226,N_410);
nand U1408 (N_1408,N_795,N_233);
and U1409 (N_1409,N_274,In_1525);
xnor U1410 (N_1410,N_570,N_360);
nand U1411 (N_1411,In_1931,N_431);
or U1412 (N_1412,N_59,N_577);
or U1413 (N_1413,In_1553,In_1950);
nand U1414 (N_1414,In_1410,In_226);
or U1415 (N_1415,N_254,In_1352);
and U1416 (N_1416,N_596,In_1487);
nand U1417 (N_1417,N_135,N_687);
nand U1418 (N_1418,N_641,N_228);
nand U1419 (N_1419,N_733,N_362);
nand U1420 (N_1420,In_1317,In_1166);
nand U1421 (N_1421,N_98,In_921);
nand U1422 (N_1422,N_639,N_120);
nor U1423 (N_1423,N_83,N_105);
xor U1424 (N_1424,N_243,N_253);
or U1425 (N_1425,N_305,N_661);
or U1426 (N_1426,N_25,N_692);
or U1427 (N_1427,N_243,In_1647);
or U1428 (N_1428,In_1724,N_786);
and U1429 (N_1429,In_936,In_1495);
and U1430 (N_1430,N_545,In_375);
and U1431 (N_1431,N_588,N_700);
nand U1432 (N_1432,In_1178,N_347);
and U1433 (N_1433,N_61,In_1567);
nand U1434 (N_1434,N_434,N_774);
and U1435 (N_1435,N_639,N_511);
nor U1436 (N_1436,N_678,N_450);
and U1437 (N_1437,N_325,N_540);
or U1438 (N_1438,N_431,In_1031);
nand U1439 (N_1439,In_1641,N_694);
or U1440 (N_1440,N_531,N_660);
nand U1441 (N_1441,In_1989,In_796);
xor U1442 (N_1442,In_135,In_941);
and U1443 (N_1443,N_404,N_778);
and U1444 (N_1444,In_418,In_985);
or U1445 (N_1445,In_558,N_309);
and U1446 (N_1446,N_556,N_318);
nor U1447 (N_1447,N_551,N_523);
and U1448 (N_1448,N_184,N_347);
nor U1449 (N_1449,N_443,In_1897);
nand U1450 (N_1450,N_601,N_471);
and U1451 (N_1451,N_414,N_164);
nor U1452 (N_1452,In_1310,N_694);
xor U1453 (N_1453,N_710,In_1052);
and U1454 (N_1454,N_286,N_725);
nor U1455 (N_1455,N_151,N_372);
nand U1456 (N_1456,In_1885,N_447);
and U1457 (N_1457,N_482,In_952);
nor U1458 (N_1458,In_694,N_681);
nand U1459 (N_1459,N_229,N_3);
nand U1460 (N_1460,In_105,N_12);
nand U1461 (N_1461,N_561,N_379);
nand U1462 (N_1462,N_571,In_1962);
nand U1463 (N_1463,N_101,N_293);
nor U1464 (N_1464,N_253,In_1140);
or U1465 (N_1465,N_701,N_372);
or U1466 (N_1466,N_697,In_1060);
nor U1467 (N_1467,N_695,N_632);
nor U1468 (N_1468,N_407,In_1283);
nand U1469 (N_1469,N_689,N_351);
nor U1470 (N_1470,N_676,N_661);
nor U1471 (N_1471,N_516,N_300);
nor U1472 (N_1472,N_765,N_438);
and U1473 (N_1473,In_677,In_1756);
nor U1474 (N_1474,In_1310,N_72);
and U1475 (N_1475,N_192,N_706);
nand U1476 (N_1476,In_77,In_238);
and U1477 (N_1477,N_470,N_594);
nor U1478 (N_1478,In_94,N_18);
nand U1479 (N_1479,In_1600,N_186);
and U1480 (N_1480,N_587,N_545);
nor U1481 (N_1481,In_49,N_615);
and U1482 (N_1482,N_122,N_523);
nor U1483 (N_1483,N_750,N_541);
nand U1484 (N_1484,N_252,N_325);
nand U1485 (N_1485,N_344,N_249);
or U1486 (N_1486,In_1547,N_149);
and U1487 (N_1487,In_936,N_97);
nor U1488 (N_1488,In_443,N_249);
and U1489 (N_1489,N_724,N_315);
nand U1490 (N_1490,N_686,N_537);
or U1491 (N_1491,In_1480,In_269);
and U1492 (N_1492,N_688,In_1261);
nand U1493 (N_1493,N_727,N_247);
nand U1494 (N_1494,N_334,N_479);
nor U1495 (N_1495,N_705,N_130);
nor U1496 (N_1496,N_396,N_465);
and U1497 (N_1497,N_768,N_393);
or U1498 (N_1498,N_522,In_328);
and U1499 (N_1499,In_46,In_68);
nand U1500 (N_1500,In_1685,N_526);
nand U1501 (N_1501,In_877,In_1472);
and U1502 (N_1502,N_742,N_279);
or U1503 (N_1503,N_547,N_734);
nand U1504 (N_1504,N_66,N_554);
or U1505 (N_1505,In_441,N_462);
and U1506 (N_1506,N_602,N_84);
and U1507 (N_1507,In_1247,N_18);
or U1508 (N_1508,N_531,In_1367);
or U1509 (N_1509,N_641,N_415);
or U1510 (N_1510,In_94,N_334);
or U1511 (N_1511,N_31,N_334);
and U1512 (N_1512,N_674,N_744);
nand U1513 (N_1513,In_1590,In_421);
nor U1514 (N_1514,N_481,N_329);
or U1515 (N_1515,In_566,In_1409);
nor U1516 (N_1516,In_1283,N_296);
or U1517 (N_1517,In_1896,N_490);
nand U1518 (N_1518,N_324,N_366);
nor U1519 (N_1519,N_24,N_378);
and U1520 (N_1520,N_169,N_534);
and U1521 (N_1521,In_664,In_968);
nor U1522 (N_1522,N_371,N_293);
and U1523 (N_1523,N_311,In_1641);
and U1524 (N_1524,In_1974,In_1926);
nand U1525 (N_1525,N_682,N_86);
nor U1526 (N_1526,N_599,N_501);
or U1527 (N_1527,In_673,N_273);
nor U1528 (N_1528,In_639,N_149);
and U1529 (N_1529,N_217,In_1897);
nor U1530 (N_1530,N_573,N_530);
or U1531 (N_1531,In_1195,N_518);
or U1532 (N_1532,N_325,In_1746);
nand U1533 (N_1533,N_10,In_1931);
nand U1534 (N_1534,In_1708,N_741);
nor U1535 (N_1535,N_665,In_898);
nand U1536 (N_1536,N_379,N_308);
or U1537 (N_1537,N_751,N_301);
nand U1538 (N_1538,N_31,N_562);
nor U1539 (N_1539,N_283,In_127);
and U1540 (N_1540,N_136,N_221);
or U1541 (N_1541,N_204,N_309);
nand U1542 (N_1542,N_585,N_288);
or U1543 (N_1543,N_292,In_627);
or U1544 (N_1544,In_1930,In_1009);
or U1545 (N_1545,N_416,N_682);
and U1546 (N_1546,N_631,In_1839);
nor U1547 (N_1547,In_1901,N_575);
or U1548 (N_1548,N_599,N_244);
nor U1549 (N_1549,N_297,N_581);
or U1550 (N_1550,In_1706,N_492);
nor U1551 (N_1551,N_365,N_580);
and U1552 (N_1552,In_68,N_715);
nor U1553 (N_1553,N_644,N_715);
or U1554 (N_1554,N_439,N_267);
nor U1555 (N_1555,In_1288,N_298);
nor U1556 (N_1556,In_1009,N_705);
or U1557 (N_1557,N_446,N_767);
and U1558 (N_1558,In_1012,N_396);
nand U1559 (N_1559,N_327,N_569);
nor U1560 (N_1560,N_752,N_356);
or U1561 (N_1561,N_746,In_1984);
nor U1562 (N_1562,N_253,N_277);
and U1563 (N_1563,N_682,In_383);
or U1564 (N_1564,In_1625,In_1157);
or U1565 (N_1565,N_265,In_1542);
or U1566 (N_1566,N_370,N_346);
nand U1567 (N_1567,N_542,In_1430);
and U1568 (N_1568,N_392,In_270);
nand U1569 (N_1569,In_487,N_657);
xor U1570 (N_1570,In_1409,N_294);
or U1571 (N_1571,N_102,N_10);
and U1572 (N_1572,In_1288,In_484);
nor U1573 (N_1573,N_213,In_956);
or U1574 (N_1574,In_1885,N_120);
nand U1575 (N_1575,N_36,N_271);
nand U1576 (N_1576,N_655,N_632);
nor U1577 (N_1577,N_535,In_828);
and U1578 (N_1578,N_505,N_118);
nand U1579 (N_1579,In_72,N_6);
nor U1580 (N_1580,N_360,N_157);
or U1581 (N_1581,In_995,N_751);
nand U1582 (N_1582,In_1008,N_10);
nor U1583 (N_1583,N_482,N_783);
nor U1584 (N_1584,In_1996,N_404);
nand U1585 (N_1585,N_265,N_732);
nand U1586 (N_1586,N_258,N_233);
nand U1587 (N_1587,In_1514,N_183);
and U1588 (N_1588,N_417,In_53);
and U1589 (N_1589,In_689,N_593);
nor U1590 (N_1590,In_941,In_459);
nor U1591 (N_1591,In_1389,N_735);
nor U1592 (N_1592,In_849,N_683);
nand U1593 (N_1593,N_428,N_123);
and U1594 (N_1594,N_175,N_294);
nand U1595 (N_1595,N_310,N_374);
and U1596 (N_1596,N_590,N_114);
and U1597 (N_1597,N_248,In_1517);
or U1598 (N_1598,N_593,N_501);
or U1599 (N_1599,In_1950,N_255);
and U1600 (N_1600,N_1228,N_1390);
or U1601 (N_1601,N_1511,N_1208);
nand U1602 (N_1602,N_1412,N_1165);
nand U1603 (N_1603,N_1264,N_1513);
nand U1604 (N_1604,N_904,N_956);
and U1605 (N_1605,N_1089,N_822);
or U1606 (N_1606,N_1189,N_1419);
nor U1607 (N_1607,N_1414,N_1094);
and U1608 (N_1608,N_1118,N_1032);
and U1609 (N_1609,N_1170,N_1048);
and U1610 (N_1610,N_1049,N_1432);
or U1611 (N_1611,N_1338,N_1096);
nor U1612 (N_1612,N_1534,N_1254);
nand U1613 (N_1613,N_917,N_1398);
or U1614 (N_1614,N_1238,N_1200);
nor U1615 (N_1615,N_1594,N_1525);
nor U1616 (N_1616,N_1372,N_1197);
nor U1617 (N_1617,N_1084,N_1476);
or U1618 (N_1618,N_898,N_807);
nor U1619 (N_1619,N_1471,N_1082);
nand U1620 (N_1620,N_1058,N_1069);
and U1621 (N_1621,N_1485,N_1126);
or U1622 (N_1622,N_1002,N_1070);
or U1623 (N_1623,N_1098,N_903);
nand U1624 (N_1624,N_840,N_1212);
xnor U1625 (N_1625,N_1143,N_968);
nand U1626 (N_1626,N_970,N_1052);
or U1627 (N_1627,N_1510,N_1233);
nor U1628 (N_1628,N_1310,N_1240);
nor U1629 (N_1629,N_1251,N_1059);
and U1630 (N_1630,N_805,N_1072);
nand U1631 (N_1631,N_1330,N_856);
nand U1632 (N_1632,N_1507,N_1029);
and U1633 (N_1633,N_1191,N_947);
or U1634 (N_1634,N_1113,N_1137);
nor U1635 (N_1635,N_1092,N_1304);
and U1636 (N_1636,N_936,N_1409);
and U1637 (N_1637,N_1363,N_1364);
xor U1638 (N_1638,N_819,N_1421);
and U1639 (N_1639,N_1076,N_967);
or U1640 (N_1640,N_1258,N_809);
and U1641 (N_1641,N_1306,N_900);
nor U1642 (N_1642,N_1248,N_1066);
or U1643 (N_1643,N_1382,N_1087);
or U1644 (N_1644,N_1033,N_901);
nand U1645 (N_1645,N_1289,N_1370);
and U1646 (N_1646,N_801,N_1568);
and U1647 (N_1647,N_1539,N_995);
nand U1648 (N_1648,N_1475,N_1544);
nand U1649 (N_1649,N_1524,N_1566);
or U1650 (N_1650,N_1314,N_1149);
or U1651 (N_1651,N_1351,N_1599);
nor U1652 (N_1652,N_1331,N_1298);
and U1653 (N_1653,N_1522,N_1071);
and U1654 (N_1654,N_919,N_1576);
nand U1655 (N_1655,N_1546,N_1027);
or U1656 (N_1656,N_1337,N_1038);
and U1657 (N_1657,N_1487,N_1423);
nor U1658 (N_1658,N_1211,N_977);
nand U1659 (N_1659,N_1270,N_1287);
or U1660 (N_1660,N_1293,N_1178);
nor U1661 (N_1661,N_1464,N_1416);
nand U1662 (N_1662,N_1352,N_1272);
nor U1663 (N_1663,N_1177,N_1396);
nand U1664 (N_1664,N_993,N_1426);
nor U1665 (N_1665,N_1110,N_1360);
or U1666 (N_1666,N_1425,N_1107);
nand U1667 (N_1667,N_1242,N_1493);
and U1668 (N_1668,N_1533,N_1588);
nor U1669 (N_1669,N_1129,N_1342);
or U1670 (N_1670,N_1144,N_1388);
or U1671 (N_1671,N_1296,N_1561);
or U1672 (N_1672,N_905,N_1168);
or U1673 (N_1673,N_1543,N_844);
and U1674 (N_1674,N_1462,N_1291);
or U1675 (N_1675,N_1325,N_1132);
nand U1676 (N_1676,N_1210,N_1173);
nand U1677 (N_1677,N_1035,N_923);
or U1678 (N_1678,N_938,N_1369);
and U1679 (N_1679,N_1009,N_1060);
nand U1680 (N_1680,N_1551,N_969);
or U1681 (N_1681,N_957,N_1246);
nand U1682 (N_1682,N_1295,N_1452);
nor U1683 (N_1683,N_1275,N_1316);
or U1684 (N_1684,N_1044,N_1181);
nand U1685 (N_1685,N_1108,N_1245);
and U1686 (N_1686,N_1010,N_1499);
nand U1687 (N_1687,N_1365,N_1121);
or U1688 (N_1688,N_951,N_1252);
and U1689 (N_1689,N_1570,N_1237);
nand U1690 (N_1690,N_1063,N_889);
nor U1691 (N_1691,N_1083,N_1263);
nand U1692 (N_1692,N_1103,N_850);
or U1693 (N_1693,N_1013,N_1117);
and U1694 (N_1694,N_821,N_1313);
nand U1695 (N_1695,N_954,N_1508);
nor U1696 (N_1696,N_1196,N_961);
nand U1697 (N_1697,N_1285,N_1180);
nand U1698 (N_1698,N_1589,N_1241);
nand U1699 (N_1699,N_833,N_914);
nand U1700 (N_1700,N_866,N_959);
or U1701 (N_1701,N_983,N_1091);
and U1702 (N_1702,N_1549,N_930);
nand U1703 (N_1703,N_1185,N_1582);
nor U1704 (N_1704,N_1006,N_820);
or U1705 (N_1705,N_1505,N_1175);
nand U1706 (N_1706,N_1250,N_1504);
nand U1707 (N_1707,N_1068,N_860);
nor U1708 (N_1708,N_1016,N_1481);
nand U1709 (N_1709,N_857,N_1535);
nor U1710 (N_1710,N_1407,N_1111);
nand U1711 (N_1711,N_1024,N_1008);
nand U1712 (N_1712,N_808,N_1440);
and U1713 (N_1713,N_1519,N_1547);
or U1714 (N_1714,N_1274,N_1453);
and U1715 (N_1715,N_949,N_1301);
or U1716 (N_1716,N_1431,N_989);
nand U1717 (N_1717,N_1430,N_1494);
or U1718 (N_1718,N_926,N_952);
and U1719 (N_1719,N_848,N_1427);
nor U1720 (N_1720,N_884,N_1190);
nand U1721 (N_1721,N_1176,N_1573);
and U1722 (N_1722,N_1000,N_1007);
nor U1723 (N_1723,N_1577,N_1429);
xor U1724 (N_1724,N_1389,N_1053);
nor U1725 (N_1725,N_843,N_1232);
or U1726 (N_1726,N_1575,N_1183);
and U1727 (N_1727,N_1478,N_1518);
or U1728 (N_1728,N_921,N_1514);
nor U1729 (N_1729,N_1347,N_1062);
and U1730 (N_1730,N_1156,N_803);
and U1731 (N_1731,N_1267,N_1202);
and U1732 (N_1732,N_1090,N_1552);
and U1733 (N_1733,N_1184,N_1413);
nand U1734 (N_1734,N_896,N_873);
nand U1735 (N_1735,N_1135,N_1222);
nand U1736 (N_1736,N_1154,N_1278);
or U1737 (N_1737,N_916,N_1186);
nand U1738 (N_1738,N_1217,N_1131);
or U1739 (N_1739,N_1377,N_1437);
or U1740 (N_1740,N_1284,N_1290);
nor U1741 (N_1741,N_1124,N_1147);
or U1742 (N_1742,N_1537,N_1381);
nor U1743 (N_1743,N_1417,N_1410);
or U1744 (N_1744,N_1580,N_988);
nor U1745 (N_1745,N_915,N_1468);
nand U1746 (N_1746,N_1520,N_1495);
nor U1747 (N_1747,N_1327,N_892);
nand U1748 (N_1748,N_1502,N_1030);
and U1749 (N_1749,N_1442,N_1253);
nand U1750 (N_1750,N_1554,N_1459);
or U1751 (N_1751,N_1473,N_980);
or U1752 (N_1752,N_1555,N_1122);
and U1753 (N_1753,N_881,N_1393);
nand U1754 (N_1754,N_875,N_1503);
and U1755 (N_1755,N_817,N_1260);
nor U1756 (N_1756,N_1448,N_1578);
nor U1757 (N_1757,N_1061,N_940);
nand U1758 (N_1758,N_1492,N_1422);
nor U1759 (N_1759,N_1465,N_1333);
and U1760 (N_1760,N_1309,N_1336);
nand U1761 (N_1761,N_981,N_1065);
nand U1762 (N_1762,N_877,N_1012);
nand U1763 (N_1763,N_1257,N_1457);
nand U1764 (N_1764,N_1023,N_1564);
and U1765 (N_1765,N_1559,N_1404);
nand U1766 (N_1766,N_1483,N_1350);
nand U1767 (N_1767,N_906,N_1400);
and U1768 (N_1768,N_1307,N_1596);
and U1769 (N_1769,N_1073,N_1281);
xor U1770 (N_1770,N_1540,N_945);
nor U1771 (N_1771,N_838,N_907);
nand U1772 (N_1772,N_1401,N_1215);
and U1773 (N_1773,N_1420,N_1488);
nor U1774 (N_1774,N_1585,N_1560);
nor U1775 (N_1775,N_958,N_1584);
and U1776 (N_1776,N_1315,N_1406);
or U1777 (N_1777,N_1075,N_1277);
nor U1778 (N_1778,N_1467,N_876);
nor U1779 (N_1779,N_909,N_1358);
or U1780 (N_1780,N_1501,N_1374);
or U1781 (N_1781,N_872,N_879);
nand U1782 (N_1782,N_972,N_1288);
nand U1783 (N_1783,N_1162,N_1171);
or U1784 (N_1784,N_1286,N_1256);
nand U1785 (N_1785,N_964,N_1034);
or U1786 (N_1786,N_1179,N_1067);
nand U1787 (N_1787,N_913,N_944);
nor U1788 (N_1788,N_1055,N_870);
and U1789 (N_1789,N_1120,N_1234);
nor U1790 (N_1790,N_1490,N_1138);
nand U1791 (N_1791,N_882,N_1188);
nor U1792 (N_1792,N_1155,N_1036);
nand U1793 (N_1793,N_1335,N_894);
and U1794 (N_1794,N_1074,N_1346);
nand U1795 (N_1795,N_1099,N_1198);
and U1796 (N_1796,N_1158,N_994);
and U1797 (N_1797,N_946,N_1500);
nor U1798 (N_1798,N_1341,N_1102);
or U1799 (N_1799,N_868,N_1593);
and U1800 (N_1800,N_1086,N_1153);
nor U1801 (N_1801,N_1395,N_854);
nor U1802 (N_1802,N_1526,N_1164);
nor U1803 (N_1803,N_971,N_1088);
or U1804 (N_1804,N_1187,N_1109);
or U1805 (N_1805,N_990,N_1343);
nor U1806 (N_1806,N_1141,N_1380);
or U1807 (N_1807,N_1025,N_1322);
and U1808 (N_1808,N_1265,N_1486);
xor U1809 (N_1809,N_1408,N_948);
nand U1810 (N_1810,N_1302,N_1031);
and U1811 (N_1811,N_1095,N_1050);
nor U1812 (N_1812,N_810,N_934);
nand U1813 (N_1813,N_1216,N_1591);
or U1814 (N_1814,N_1116,N_1105);
nor U1815 (N_1815,N_1283,N_1041);
nand U1816 (N_1816,N_929,N_1039);
nor U1817 (N_1817,N_832,N_924);
or U1818 (N_1818,N_1446,N_1362);
nor U1819 (N_1819,N_886,N_1026);
nand U1820 (N_1820,N_1563,N_862);
or U1821 (N_1821,N_1045,N_891);
nor U1822 (N_1822,N_847,N_1498);
and U1823 (N_1823,N_1064,N_859);
nor U1824 (N_1824,N_1454,N_1332);
nor U1825 (N_1825,N_812,N_1182);
or U1826 (N_1826,N_842,N_1199);
or U1827 (N_1827,N_1451,N_1455);
nand U1828 (N_1828,N_890,N_1139);
nor U1829 (N_1829,N_823,N_1128);
and U1830 (N_1830,N_826,N_1345);
or U1831 (N_1831,N_939,N_1586);
or U1832 (N_1832,N_1461,N_1279);
and U1833 (N_1833,N_1472,N_1203);
or U1834 (N_1834,N_1097,N_1349);
or U1835 (N_1835,N_897,N_852);
nand U1836 (N_1836,N_815,N_1312);
or U1837 (N_1837,N_871,N_1040);
or U1838 (N_1838,N_1324,N_1292);
and U1839 (N_1839,N_1001,N_1474);
and U1840 (N_1840,N_1460,N_1541);
and U1841 (N_1841,N_1375,N_943);
or U1842 (N_1842,N_992,N_1348);
and U1843 (N_1843,N_1411,N_1367);
or U1844 (N_1844,N_1236,N_813);
nand U1845 (N_1845,N_839,N_950);
nand U1846 (N_1846,N_1479,N_1043);
and U1847 (N_1847,N_966,N_1046);
or U1848 (N_1848,N_1249,N_1469);
nand U1849 (N_1849,N_1506,N_1100);
and U1850 (N_1850,N_841,N_806);
and U1851 (N_1851,N_973,N_1078);
nand U1852 (N_1852,N_1444,N_830);
nand U1853 (N_1853,N_1392,N_1015);
and U1854 (N_1854,N_1042,N_1019);
or U1855 (N_1855,N_1515,N_1572);
nand U1856 (N_1856,N_1399,N_1266);
nor U1857 (N_1857,N_835,N_984);
and U1858 (N_1858,N_1394,N_1590);
and U1859 (N_1859,N_1536,N_895);
nor U1860 (N_1860,N_1428,N_1230);
and U1861 (N_1861,N_963,N_1353);
or U1862 (N_1862,N_1418,N_925);
nand U1863 (N_1863,N_1509,N_1466);
nor U1864 (N_1864,N_1136,N_1359);
and U1865 (N_1865,N_1201,N_1329);
nor U1866 (N_1866,N_1447,N_1209);
nand U1867 (N_1867,N_1553,N_902);
and U1868 (N_1868,N_1161,N_1166);
nor U1869 (N_1869,N_927,N_975);
nand U1870 (N_1870,N_997,N_1357);
nor U1871 (N_1871,N_853,N_1273);
xor U1872 (N_1872,N_1127,N_1403);
nor U1873 (N_1873,N_928,N_1402);
nor U1874 (N_1874,N_1268,N_1597);
or U1875 (N_1875,N_1017,N_1424);
and U1876 (N_1876,N_1021,N_1458);
nand U1877 (N_1877,N_1300,N_834);
and U1878 (N_1878,N_1262,N_1221);
nand U1879 (N_1879,N_955,N_1523);
and U1880 (N_1880,N_1150,N_1435);
nor U1881 (N_1881,N_1206,N_1548);
nor U1882 (N_1882,N_1558,N_1383);
nand U1883 (N_1883,N_1169,N_1583);
nor U1884 (N_1884,N_1361,N_811);
nor U1885 (N_1885,N_1114,N_1319);
nand U1886 (N_1886,N_1157,N_1320);
nor U1887 (N_1887,N_1449,N_1512);
and U1888 (N_1888,N_1480,N_1517);
or U1889 (N_1889,N_1521,N_867);
and U1890 (N_1890,N_1484,N_1530);
or U1891 (N_1891,N_1456,N_1595);
nor U1892 (N_1892,N_1080,N_1311);
or U1893 (N_1893,N_1318,N_1556);
and U1894 (N_1894,N_1334,N_1101);
and U1895 (N_1895,N_829,N_1112);
and U1896 (N_1896,N_855,N_953);
nand U1897 (N_1897,N_1477,N_1214);
nand U1898 (N_1898,N_1218,N_1294);
or U1899 (N_1899,N_1328,N_858);
nand U1900 (N_1900,N_1125,N_1243);
nand U1901 (N_1901,N_1276,N_931);
nand U1902 (N_1902,N_1305,N_814);
nand U1903 (N_1903,N_1356,N_935);
nor U1904 (N_1904,N_1443,N_887);
or U1905 (N_1905,N_1308,N_1571);
nand U1906 (N_1906,N_1378,N_899);
nor U1907 (N_1907,N_863,N_837);
or U1908 (N_1908,N_1271,N_1592);
nor U1909 (N_1909,N_1227,N_1445);
nor U1910 (N_1910,N_1531,N_985);
and U1911 (N_1911,N_1354,N_1204);
nor U1912 (N_1912,N_1282,N_1567);
and U1913 (N_1913,N_1133,N_1077);
or U1914 (N_1914,N_1532,N_1441);
nor U1915 (N_1915,N_1193,N_910);
and U1916 (N_1916,N_1145,N_1172);
and U1917 (N_1917,N_846,N_1142);
or U1918 (N_1918,N_1219,N_880);
or U1919 (N_1919,N_1545,N_869);
and U1920 (N_1920,N_816,N_1387);
and U1921 (N_1921,N_1255,N_893);
nand U1922 (N_1922,N_1056,N_1439);
nor U1923 (N_1923,N_1205,N_996);
nor U1924 (N_1924,N_827,N_1079);
nand U1925 (N_1925,N_883,N_999);
nor U1926 (N_1926,N_1497,N_942);
and U1927 (N_1927,N_849,N_1436);
and U1928 (N_1928,N_1384,N_1003);
nand U1929 (N_1929,N_888,N_831);
and U1930 (N_1930,N_1491,N_1081);
or U1931 (N_1931,N_802,N_1280);
or U1932 (N_1932,N_874,N_1174);
and U1933 (N_1933,N_1119,N_1220);
nand U1934 (N_1934,N_804,N_1368);
nand U1935 (N_1935,N_1482,N_1579);
nand U1936 (N_1936,N_1226,N_1229);
nand U1937 (N_1937,N_908,N_987);
nor U1938 (N_1938,N_1397,N_818);
or U1939 (N_1939,N_1123,N_1011);
nor U1940 (N_1940,N_937,N_1542);
nand U1941 (N_1941,N_1018,N_1047);
nand U1942 (N_1942,N_962,N_1528);
nor U1943 (N_1943,N_864,N_1085);
and U1944 (N_1944,N_1529,N_1148);
nand U1945 (N_1945,N_1167,N_1463);
nor U1946 (N_1946,N_933,N_1005);
nand U1947 (N_1947,N_800,N_1489);
and U1948 (N_1948,N_1391,N_974);
and U1949 (N_1949,N_1450,N_1057);
nor U1950 (N_1950,N_1516,N_828);
or U1951 (N_1951,N_1130,N_1574);
nor U1952 (N_1952,N_1366,N_1223);
nor U1953 (N_1953,N_865,N_885);
and U1954 (N_1954,N_1159,N_878);
and U1955 (N_1955,N_1244,N_1231);
and U1956 (N_1956,N_824,N_1259);
nor U1957 (N_1957,N_979,N_1317);
nor U1958 (N_1958,N_1207,N_851);
or U1959 (N_1959,N_1598,N_1192);
and U1960 (N_1960,N_1355,N_1470);
nand U1961 (N_1961,N_1303,N_1022);
or U1962 (N_1962,N_1297,N_1323);
nand U1963 (N_1963,N_1247,N_922);
nand U1964 (N_1964,N_1093,N_1340);
and U1965 (N_1965,N_1213,N_1051);
and U1966 (N_1966,N_1134,N_986);
or U1967 (N_1967,N_1321,N_1496);
or U1968 (N_1968,N_1379,N_911);
nand U1969 (N_1969,N_1569,N_1140);
or U1970 (N_1970,N_1261,N_1037);
and U1971 (N_1971,N_1344,N_1020);
nor U1972 (N_1972,N_1195,N_825);
or U1973 (N_1973,N_991,N_1004);
and U1974 (N_1974,N_941,N_1550);
and U1975 (N_1975,N_845,N_1562);
or U1976 (N_1976,N_1269,N_1386);
or U1977 (N_1977,N_1433,N_918);
or U1978 (N_1978,N_1565,N_1225);
nor U1979 (N_1979,N_1104,N_1299);
nor U1980 (N_1980,N_1028,N_920);
nor U1981 (N_1981,N_1376,N_1194);
nor U1982 (N_1982,N_912,N_1557);
and U1983 (N_1983,N_1239,N_1371);
nor U1984 (N_1984,N_1160,N_1152);
nand U1985 (N_1985,N_978,N_1415);
and U1986 (N_1986,N_1146,N_1438);
xnor U1987 (N_1987,N_1163,N_1106);
nor U1988 (N_1988,N_1014,N_1339);
or U1989 (N_1989,N_1385,N_1235);
and U1990 (N_1990,N_1405,N_998);
and U1991 (N_1991,N_1527,N_965);
or U1992 (N_1992,N_1538,N_1151);
nand U1993 (N_1993,N_1326,N_1587);
or U1994 (N_1994,N_1373,N_1115);
nor U1995 (N_1995,N_1434,N_1054);
or U1996 (N_1996,N_836,N_861);
nor U1997 (N_1997,N_1581,N_960);
xnor U1998 (N_1998,N_982,N_1224);
and U1999 (N_1999,N_932,N_976);
nor U2000 (N_2000,N_1341,N_1349);
nor U2001 (N_2001,N_1339,N_960);
and U2002 (N_2002,N_1376,N_1340);
and U2003 (N_2003,N_1597,N_1013);
nor U2004 (N_2004,N_906,N_1577);
and U2005 (N_2005,N_948,N_1596);
and U2006 (N_2006,N_938,N_806);
or U2007 (N_2007,N_1369,N_1518);
or U2008 (N_2008,N_1237,N_1319);
nor U2009 (N_2009,N_1014,N_879);
or U2010 (N_2010,N_909,N_1247);
nor U2011 (N_2011,N_841,N_1110);
and U2012 (N_2012,N_1515,N_914);
and U2013 (N_2013,N_930,N_831);
nand U2014 (N_2014,N_1138,N_1301);
and U2015 (N_2015,N_1573,N_800);
nor U2016 (N_2016,N_1020,N_883);
and U2017 (N_2017,N_1332,N_1266);
and U2018 (N_2018,N_1164,N_1284);
nor U2019 (N_2019,N_933,N_926);
nand U2020 (N_2020,N_831,N_1051);
nor U2021 (N_2021,N_862,N_1297);
nand U2022 (N_2022,N_965,N_874);
nand U2023 (N_2023,N_1038,N_1046);
and U2024 (N_2024,N_1553,N_1258);
or U2025 (N_2025,N_1538,N_1031);
or U2026 (N_2026,N_1420,N_1380);
nand U2027 (N_2027,N_871,N_1049);
nor U2028 (N_2028,N_1513,N_1445);
nand U2029 (N_2029,N_1072,N_1501);
or U2030 (N_2030,N_1586,N_973);
nand U2031 (N_2031,N_1239,N_1463);
or U2032 (N_2032,N_1318,N_1250);
nand U2033 (N_2033,N_1003,N_965);
or U2034 (N_2034,N_1330,N_1345);
or U2035 (N_2035,N_1332,N_1256);
or U2036 (N_2036,N_1066,N_1093);
nor U2037 (N_2037,N_1125,N_1217);
nor U2038 (N_2038,N_1446,N_1110);
nor U2039 (N_2039,N_949,N_1183);
nand U2040 (N_2040,N_811,N_974);
and U2041 (N_2041,N_897,N_1279);
nand U2042 (N_2042,N_1575,N_920);
nand U2043 (N_2043,N_1174,N_942);
nor U2044 (N_2044,N_1063,N_1203);
nor U2045 (N_2045,N_1309,N_1261);
or U2046 (N_2046,N_1184,N_1502);
or U2047 (N_2047,N_898,N_1453);
and U2048 (N_2048,N_1271,N_1083);
or U2049 (N_2049,N_1325,N_853);
nand U2050 (N_2050,N_1435,N_843);
nand U2051 (N_2051,N_880,N_1598);
and U2052 (N_2052,N_1216,N_1258);
nor U2053 (N_2053,N_1468,N_965);
and U2054 (N_2054,N_1225,N_833);
and U2055 (N_2055,N_1129,N_1142);
nand U2056 (N_2056,N_1185,N_1274);
nor U2057 (N_2057,N_1122,N_1271);
or U2058 (N_2058,N_1338,N_824);
and U2059 (N_2059,N_1439,N_974);
nor U2060 (N_2060,N_1362,N_1223);
nand U2061 (N_2061,N_1177,N_874);
and U2062 (N_2062,N_1552,N_1469);
and U2063 (N_2063,N_802,N_1022);
nand U2064 (N_2064,N_1491,N_1557);
and U2065 (N_2065,N_1097,N_959);
nand U2066 (N_2066,N_1100,N_940);
nand U2067 (N_2067,N_1232,N_1003);
nor U2068 (N_2068,N_1095,N_948);
or U2069 (N_2069,N_1440,N_931);
or U2070 (N_2070,N_1292,N_1191);
and U2071 (N_2071,N_1171,N_1026);
or U2072 (N_2072,N_1423,N_1214);
and U2073 (N_2073,N_941,N_896);
or U2074 (N_2074,N_1082,N_1465);
nand U2075 (N_2075,N_1070,N_1434);
nand U2076 (N_2076,N_823,N_1007);
or U2077 (N_2077,N_1497,N_935);
nand U2078 (N_2078,N_1494,N_1102);
and U2079 (N_2079,N_876,N_1177);
and U2080 (N_2080,N_1341,N_1039);
nand U2081 (N_2081,N_840,N_1533);
nor U2082 (N_2082,N_1409,N_1480);
or U2083 (N_2083,N_1050,N_1186);
or U2084 (N_2084,N_1058,N_1442);
nor U2085 (N_2085,N_1399,N_895);
or U2086 (N_2086,N_1175,N_1498);
or U2087 (N_2087,N_1591,N_1385);
nand U2088 (N_2088,N_898,N_1282);
and U2089 (N_2089,N_908,N_1506);
and U2090 (N_2090,N_1494,N_1588);
nand U2091 (N_2091,N_1004,N_1115);
and U2092 (N_2092,N_1193,N_1309);
nand U2093 (N_2093,N_953,N_1115);
and U2094 (N_2094,N_1202,N_952);
and U2095 (N_2095,N_1589,N_1471);
nor U2096 (N_2096,N_1114,N_1589);
nor U2097 (N_2097,N_808,N_802);
nor U2098 (N_2098,N_1317,N_1478);
and U2099 (N_2099,N_1150,N_1345);
and U2100 (N_2100,N_1172,N_1093);
nor U2101 (N_2101,N_996,N_1186);
nand U2102 (N_2102,N_1444,N_1008);
or U2103 (N_2103,N_824,N_1529);
and U2104 (N_2104,N_958,N_837);
or U2105 (N_2105,N_1467,N_1508);
nand U2106 (N_2106,N_1364,N_1577);
or U2107 (N_2107,N_931,N_1016);
nand U2108 (N_2108,N_1333,N_953);
nor U2109 (N_2109,N_1461,N_1374);
or U2110 (N_2110,N_1325,N_1154);
or U2111 (N_2111,N_1497,N_1041);
nand U2112 (N_2112,N_1407,N_1464);
xor U2113 (N_2113,N_1435,N_1199);
nand U2114 (N_2114,N_1564,N_1598);
nand U2115 (N_2115,N_836,N_893);
nor U2116 (N_2116,N_806,N_1126);
nor U2117 (N_2117,N_812,N_1225);
or U2118 (N_2118,N_1454,N_944);
nor U2119 (N_2119,N_970,N_1127);
or U2120 (N_2120,N_1306,N_1032);
and U2121 (N_2121,N_911,N_1437);
nand U2122 (N_2122,N_1457,N_1509);
or U2123 (N_2123,N_1229,N_1516);
and U2124 (N_2124,N_1028,N_826);
nand U2125 (N_2125,N_1419,N_875);
or U2126 (N_2126,N_1293,N_992);
nand U2127 (N_2127,N_1214,N_1109);
or U2128 (N_2128,N_1425,N_1039);
nor U2129 (N_2129,N_1233,N_895);
nor U2130 (N_2130,N_1227,N_940);
nor U2131 (N_2131,N_1014,N_998);
and U2132 (N_2132,N_1154,N_1078);
nor U2133 (N_2133,N_1330,N_1103);
nand U2134 (N_2134,N_1365,N_1332);
and U2135 (N_2135,N_1344,N_943);
nor U2136 (N_2136,N_1463,N_985);
nand U2137 (N_2137,N_1526,N_1583);
and U2138 (N_2138,N_1303,N_912);
or U2139 (N_2139,N_967,N_1118);
nand U2140 (N_2140,N_1432,N_1308);
nand U2141 (N_2141,N_1409,N_1218);
nand U2142 (N_2142,N_1013,N_1030);
and U2143 (N_2143,N_1556,N_1340);
nand U2144 (N_2144,N_1544,N_823);
nand U2145 (N_2145,N_1072,N_1561);
and U2146 (N_2146,N_1256,N_1352);
nor U2147 (N_2147,N_1442,N_817);
or U2148 (N_2148,N_1039,N_1185);
nand U2149 (N_2149,N_856,N_1225);
nor U2150 (N_2150,N_1339,N_852);
and U2151 (N_2151,N_1136,N_1355);
nor U2152 (N_2152,N_919,N_1345);
and U2153 (N_2153,N_1074,N_923);
nand U2154 (N_2154,N_1433,N_1304);
nor U2155 (N_2155,N_1587,N_945);
nor U2156 (N_2156,N_1454,N_970);
and U2157 (N_2157,N_1398,N_1103);
nor U2158 (N_2158,N_1011,N_1049);
and U2159 (N_2159,N_881,N_1076);
nand U2160 (N_2160,N_1478,N_1410);
nand U2161 (N_2161,N_1078,N_846);
nor U2162 (N_2162,N_1282,N_1029);
and U2163 (N_2163,N_1121,N_1596);
or U2164 (N_2164,N_1198,N_1548);
and U2165 (N_2165,N_1472,N_1372);
nand U2166 (N_2166,N_975,N_1113);
or U2167 (N_2167,N_1144,N_914);
and U2168 (N_2168,N_1398,N_1122);
nor U2169 (N_2169,N_1427,N_1116);
and U2170 (N_2170,N_1173,N_1179);
nand U2171 (N_2171,N_1371,N_943);
nor U2172 (N_2172,N_902,N_1409);
and U2173 (N_2173,N_1446,N_1225);
and U2174 (N_2174,N_1143,N_844);
and U2175 (N_2175,N_1471,N_1462);
nor U2176 (N_2176,N_1533,N_1307);
nor U2177 (N_2177,N_802,N_1117);
nor U2178 (N_2178,N_1184,N_984);
nand U2179 (N_2179,N_1310,N_1231);
and U2180 (N_2180,N_1279,N_1282);
nor U2181 (N_2181,N_1475,N_1084);
or U2182 (N_2182,N_965,N_1293);
nand U2183 (N_2183,N_1148,N_1117);
nand U2184 (N_2184,N_1261,N_997);
and U2185 (N_2185,N_1174,N_926);
nand U2186 (N_2186,N_1470,N_930);
nand U2187 (N_2187,N_1180,N_1291);
or U2188 (N_2188,N_1267,N_967);
and U2189 (N_2189,N_1581,N_1004);
nand U2190 (N_2190,N_1399,N_1126);
nor U2191 (N_2191,N_1387,N_1414);
and U2192 (N_2192,N_1484,N_937);
or U2193 (N_2193,N_1091,N_907);
xor U2194 (N_2194,N_817,N_1106);
nor U2195 (N_2195,N_1235,N_1397);
nor U2196 (N_2196,N_1270,N_1319);
or U2197 (N_2197,N_1489,N_1110);
and U2198 (N_2198,N_1395,N_1244);
nor U2199 (N_2199,N_1376,N_1533);
nor U2200 (N_2200,N_1171,N_1548);
nand U2201 (N_2201,N_818,N_1158);
and U2202 (N_2202,N_1521,N_1198);
and U2203 (N_2203,N_914,N_1399);
nor U2204 (N_2204,N_1283,N_1415);
nor U2205 (N_2205,N_1055,N_1058);
or U2206 (N_2206,N_1585,N_1065);
and U2207 (N_2207,N_1276,N_1414);
nor U2208 (N_2208,N_843,N_1471);
or U2209 (N_2209,N_1382,N_1404);
nor U2210 (N_2210,N_1040,N_1135);
nor U2211 (N_2211,N_844,N_978);
and U2212 (N_2212,N_954,N_892);
nand U2213 (N_2213,N_824,N_1266);
or U2214 (N_2214,N_1038,N_1305);
nand U2215 (N_2215,N_1481,N_1068);
nor U2216 (N_2216,N_925,N_1034);
or U2217 (N_2217,N_991,N_1484);
nand U2218 (N_2218,N_1525,N_807);
nand U2219 (N_2219,N_938,N_1337);
nor U2220 (N_2220,N_1144,N_1564);
nand U2221 (N_2221,N_803,N_1225);
or U2222 (N_2222,N_1286,N_1557);
nand U2223 (N_2223,N_1185,N_1463);
and U2224 (N_2224,N_862,N_1195);
and U2225 (N_2225,N_1580,N_1257);
and U2226 (N_2226,N_1115,N_1299);
nor U2227 (N_2227,N_1092,N_977);
nor U2228 (N_2228,N_1225,N_1357);
and U2229 (N_2229,N_1424,N_915);
or U2230 (N_2230,N_1491,N_871);
nand U2231 (N_2231,N_857,N_1573);
nand U2232 (N_2232,N_1500,N_841);
nand U2233 (N_2233,N_1227,N_900);
nand U2234 (N_2234,N_1005,N_1260);
or U2235 (N_2235,N_902,N_1589);
nand U2236 (N_2236,N_1476,N_1374);
and U2237 (N_2237,N_1508,N_1325);
or U2238 (N_2238,N_823,N_1078);
or U2239 (N_2239,N_1199,N_1440);
and U2240 (N_2240,N_1073,N_1426);
and U2241 (N_2241,N_828,N_1427);
and U2242 (N_2242,N_1572,N_1302);
nor U2243 (N_2243,N_1128,N_1152);
or U2244 (N_2244,N_1387,N_1404);
and U2245 (N_2245,N_1088,N_1066);
and U2246 (N_2246,N_1252,N_1478);
nand U2247 (N_2247,N_867,N_1376);
nand U2248 (N_2248,N_827,N_1307);
nor U2249 (N_2249,N_1241,N_1530);
nand U2250 (N_2250,N_1130,N_967);
or U2251 (N_2251,N_1482,N_1140);
xnor U2252 (N_2252,N_959,N_1490);
nor U2253 (N_2253,N_1543,N_1045);
or U2254 (N_2254,N_1344,N_1397);
and U2255 (N_2255,N_1347,N_1243);
and U2256 (N_2256,N_1345,N_1112);
or U2257 (N_2257,N_1152,N_1452);
nor U2258 (N_2258,N_1453,N_1135);
nand U2259 (N_2259,N_1328,N_901);
nand U2260 (N_2260,N_1593,N_1353);
or U2261 (N_2261,N_1018,N_1578);
nand U2262 (N_2262,N_1065,N_871);
or U2263 (N_2263,N_829,N_988);
nor U2264 (N_2264,N_1563,N_1138);
nand U2265 (N_2265,N_1431,N_956);
nand U2266 (N_2266,N_1091,N_825);
nor U2267 (N_2267,N_1193,N_1383);
and U2268 (N_2268,N_1423,N_1365);
nor U2269 (N_2269,N_819,N_1023);
or U2270 (N_2270,N_1447,N_1070);
nand U2271 (N_2271,N_809,N_1042);
nand U2272 (N_2272,N_1333,N_1446);
or U2273 (N_2273,N_1190,N_922);
nor U2274 (N_2274,N_1117,N_1428);
nor U2275 (N_2275,N_1447,N_886);
nor U2276 (N_2276,N_918,N_1183);
or U2277 (N_2277,N_880,N_1080);
and U2278 (N_2278,N_1158,N_1511);
and U2279 (N_2279,N_1161,N_1110);
and U2280 (N_2280,N_1278,N_944);
nand U2281 (N_2281,N_1113,N_1270);
or U2282 (N_2282,N_1292,N_1178);
nand U2283 (N_2283,N_1554,N_1538);
nand U2284 (N_2284,N_1163,N_1040);
nand U2285 (N_2285,N_1552,N_1031);
nand U2286 (N_2286,N_1100,N_1451);
nand U2287 (N_2287,N_854,N_1318);
nand U2288 (N_2288,N_1435,N_1393);
nor U2289 (N_2289,N_1164,N_1262);
or U2290 (N_2290,N_1488,N_1407);
nand U2291 (N_2291,N_872,N_1039);
or U2292 (N_2292,N_1307,N_828);
or U2293 (N_2293,N_1046,N_1298);
and U2294 (N_2294,N_828,N_831);
nor U2295 (N_2295,N_1333,N_1599);
or U2296 (N_2296,N_1444,N_908);
or U2297 (N_2297,N_1074,N_1399);
and U2298 (N_2298,N_1214,N_858);
nand U2299 (N_2299,N_1197,N_1559);
or U2300 (N_2300,N_869,N_1383);
and U2301 (N_2301,N_1539,N_1437);
nand U2302 (N_2302,N_1107,N_1503);
nand U2303 (N_2303,N_1049,N_1174);
nand U2304 (N_2304,N_862,N_953);
and U2305 (N_2305,N_1507,N_1411);
or U2306 (N_2306,N_1379,N_1054);
and U2307 (N_2307,N_1441,N_963);
and U2308 (N_2308,N_1592,N_1047);
nand U2309 (N_2309,N_1324,N_1369);
or U2310 (N_2310,N_852,N_942);
and U2311 (N_2311,N_1316,N_991);
nand U2312 (N_2312,N_1532,N_836);
nor U2313 (N_2313,N_1568,N_1527);
or U2314 (N_2314,N_922,N_1320);
or U2315 (N_2315,N_931,N_1358);
nor U2316 (N_2316,N_892,N_1173);
or U2317 (N_2317,N_989,N_1382);
and U2318 (N_2318,N_827,N_1434);
and U2319 (N_2319,N_889,N_1235);
or U2320 (N_2320,N_1559,N_894);
nand U2321 (N_2321,N_1348,N_881);
and U2322 (N_2322,N_879,N_915);
and U2323 (N_2323,N_1369,N_1184);
and U2324 (N_2324,N_1182,N_1092);
or U2325 (N_2325,N_1171,N_1309);
nor U2326 (N_2326,N_934,N_1590);
and U2327 (N_2327,N_1439,N_1103);
and U2328 (N_2328,N_1479,N_1114);
and U2329 (N_2329,N_1098,N_881);
or U2330 (N_2330,N_1003,N_1548);
and U2331 (N_2331,N_1241,N_1536);
or U2332 (N_2332,N_884,N_1251);
and U2333 (N_2333,N_1558,N_1143);
and U2334 (N_2334,N_1360,N_1404);
and U2335 (N_2335,N_1346,N_1044);
nand U2336 (N_2336,N_1219,N_1318);
nor U2337 (N_2337,N_1139,N_1470);
and U2338 (N_2338,N_1153,N_1104);
or U2339 (N_2339,N_1167,N_1004);
xor U2340 (N_2340,N_966,N_1072);
and U2341 (N_2341,N_1554,N_1031);
and U2342 (N_2342,N_1088,N_1073);
and U2343 (N_2343,N_960,N_970);
or U2344 (N_2344,N_1598,N_899);
nor U2345 (N_2345,N_1575,N_839);
and U2346 (N_2346,N_993,N_1167);
and U2347 (N_2347,N_1510,N_1146);
xor U2348 (N_2348,N_1043,N_1514);
nor U2349 (N_2349,N_1320,N_919);
nand U2350 (N_2350,N_1291,N_1326);
nor U2351 (N_2351,N_1454,N_903);
and U2352 (N_2352,N_801,N_1339);
or U2353 (N_2353,N_1195,N_1225);
nor U2354 (N_2354,N_1001,N_1479);
and U2355 (N_2355,N_1307,N_837);
nor U2356 (N_2356,N_1567,N_1339);
and U2357 (N_2357,N_1545,N_1076);
or U2358 (N_2358,N_1275,N_915);
nor U2359 (N_2359,N_1477,N_910);
or U2360 (N_2360,N_1492,N_1335);
and U2361 (N_2361,N_1351,N_1125);
or U2362 (N_2362,N_1220,N_1081);
nor U2363 (N_2363,N_1358,N_880);
and U2364 (N_2364,N_1508,N_818);
nand U2365 (N_2365,N_1423,N_1368);
nand U2366 (N_2366,N_1368,N_1036);
or U2367 (N_2367,N_996,N_979);
nand U2368 (N_2368,N_1240,N_1096);
nand U2369 (N_2369,N_956,N_1563);
nand U2370 (N_2370,N_1576,N_1339);
or U2371 (N_2371,N_1314,N_1564);
nor U2372 (N_2372,N_1404,N_1122);
or U2373 (N_2373,N_1122,N_1287);
nor U2374 (N_2374,N_1371,N_1449);
and U2375 (N_2375,N_878,N_1190);
nand U2376 (N_2376,N_959,N_935);
nand U2377 (N_2377,N_913,N_1152);
nor U2378 (N_2378,N_1014,N_1485);
nand U2379 (N_2379,N_1293,N_889);
and U2380 (N_2380,N_1161,N_1286);
or U2381 (N_2381,N_886,N_1098);
nor U2382 (N_2382,N_1503,N_1179);
or U2383 (N_2383,N_1457,N_1193);
nor U2384 (N_2384,N_1479,N_1556);
nand U2385 (N_2385,N_1427,N_1192);
nand U2386 (N_2386,N_1452,N_1034);
nor U2387 (N_2387,N_946,N_1204);
and U2388 (N_2388,N_1370,N_1137);
and U2389 (N_2389,N_1242,N_1331);
nand U2390 (N_2390,N_1424,N_1535);
or U2391 (N_2391,N_1082,N_1175);
nand U2392 (N_2392,N_848,N_964);
and U2393 (N_2393,N_929,N_1018);
xnor U2394 (N_2394,N_1434,N_843);
or U2395 (N_2395,N_1098,N_1492);
or U2396 (N_2396,N_1528,N_1008);
and U2397 (N_2397,N_1513,N_959);
and U2398 (N_2398,N_1414,N_976);
and U2399 (N_2399,N_1350,N_1000);
nand U2400 (N_2400,N_2159,N_1824);
nor U2401 (N_2401,N_1676,N_2395);
nand U2402 (N_2402,N_1718,N_2290);
or U2403 (N_2403,N_1703,N_2312);
nor U2404 (N_2404,N_1789,N_1760);
or U2405 (N_2405,N_1684,N_2227);
nand U2406 (N_2406,N_1813,N_2381);
nor U2407 (N_2407,N_2267,N_1691);
and U2408 (N_2408,N_1957,N_1756);
nand U2409 (N_2409,N_2299,N_1977);
and U2410 (N_2410,N_2178,N_2135);
nor U2411 (N_2411,N_2286,N_2317);
or U2412 (N_2412,N_2048,N_1913);
or U2413 (N_2413,N_2077,N_1801);
and U2414 (N_2414,N_2343,N_1783);
nand U2415 (N_2415,N_2165,N_1617);
or U2416 (N_2416,N_2132,N_1959);
nand U2417 (N_2417,N_2065,N_1941);
nand U2418 (N_2418,N_2131,N_1704);
and U2419 (N_2419,N_1900,N_2150);
and U2420 (N_2420,N_2331,N_1793);
or U2421 (N_2421,N_2216,N_2330);
and U2422 (N_2422,N_2107,N_1880);
nor U2423 (N_2423,N_2021,N_1980);
nand U2424 (N_2424,N_2321,N_2119);
nand U2425 (N_2425,N_2251,N_1920);
or U2426 (N_2426,N_2003,N_2042);
nand U2427 (N_2427,N_1808,N_2380);
or U2428 (N_2428,N_1889,N_2170);
or U2429 (N_2429,N_2039,N_2089);
nand U2430 (N_2430,N_2137,N_2248);
and U2431 (N_2431,N_1794,N_2105);
nand U2432 (N_2432,N_1636,N_2151);
or U2433 (N_2433,N_2311,N_2175);
or U2434 (N_2434,N_1811,N_2180);
and U2435 (N_2435,N_2262,N_1631);
and U2436 (N_2436,N_2392,N_2364);
or U2437 (N_2437,N_1884,N_1975);
or U2438 (N_2438,N_1670,N_2253);
or U2439 (N_2439,N_2288,N_2366);
or U2440 (N_2440,N_2399,N_2111);
and U2441 (N_2441,N_1846,N_2293);
nor U2442 (N_2442,N_2204,N_1613);
nand U2443 (N_2443,N_2088,N_2052);
nor U2444 (N_2444,N_2080,N_2349);
nor U2445 (N_2445,N_2144,N_2063);
nand U2446 (N_2446,N_2238,N_2026);
nor U2447 (N_2447,N_2007,N_2022);
and U2448 (N_2448,N_2079,N_1997);
or U2449 (N_2449,N_1985,N_2398);
nor U2450 (N_2450,N_2016,N_2091);
and U2451 (N_2451,N_2250,N_2241);
and U2452 (N_2452,N_1868,N_1697);
nor U2453 (N_2453,N_2085,N_1864);
nor U2454 (N_2454,N_1615,N_1807);
and U2455 (N_2455,N_2076,N_1767);
nor U2456 (N_2456,N_2045,N_1969);
and U2457 (N_2457,N_2242,N_2305);
and U2458 (N_2458,N_1648,N_1638);
nor U2459 (N_2459,N_1902,N_1744);
and U2460 (N_2460,N_2001,N_1961);
nand U2461 (N_2461,N_2138,N_1683);
nand U2462 (N_2462,N_1943,N_2228);
nor U2463 (N_2463,N_1640,N_2154);
nand U2464 (N_2464,N_1641,N_2211);
and U2465 (N_2465,N_1962,N_2314);
nor U2466 (N_2466,N_1799,N_2086);
nand U2467 (N_2467,N_2073,N_1982);
and U2468 (N_2468,N_1994,N_2361);
nor U2469 (N_2469,N_2391,N_1669);
and U2470 (N_2470,N_2056,N_1633);
nor U2471 (N_2471,N_2316,N_1782);
or U2472 (N_2472,N_2213,N_2136);
nor U2473 (N_2473,N_2081,N_1779);
nand U2474 (N_2474,N_2327,N_1918);
and U2475 (N_2475,N_1628,N_1649);
or U2476 (N_2476,N_2249,N_1922);
and U2477 (N_2477,N_2143,N_1983);
xnor U2478 (N_2478,N_2110,N_1841);
or U2479 (N_2479,N_2212,N_2353);
and U2480 (N_2480,N_2122,N_2058);
or U2481 (N_2481,N_1623,N_2329);
and U2482 (N_2482,N_1692,N_2221);
nor U2483 (N_2483,N_1914,N_1787);
nand U2484 (N_2484,N_2372,N_2225);
and U2485 (N_2485,N_1986,N_2145);
or U2486 (N_2486,N_1600,N_1901);
or U2487 (N_2487,N_2351,N_2087);
or U2488 (N_2488,N_1788,N_1805);
nor U2489 (N_2489,N_1780,N_2005);
and U2490 (N_2490,N_1947,N_2215);
nor U2491 (N_2491,N_1791,N_1812);
nand U2492 (N_2492,N_1618,N_1777);
nand U2493 (N_2493,N_1928,N_1828);
and U2494 (N_2494,N_1652,N_1890);
or U2495 (N_2495,N_2129,N_1845);
nand U2496 (N_2496,N_2027,N_2345);
nand U2497 (N_2497,N_2390,N_2199);
xnor U2498 (N_2498,N_2033,N_2394);
and U2499 (N_2499,N_2342,N_1700);
nor U2500 (N_2500,N_1899,N_1898);
nand U2501 (N_2501,N_2050,N_1849);
nor U2502 (N_2502,N_1651,N_1912);
nor U2503 (N_2503,N_2103,N_1608);
nand U2504 (N_2504,N_2373,N_1964);
nor U2505 (N_2505,N_2169,N_1878);
nand U2506 (N_2506,N_2340,N_1911);
and U2507 (N_2507,N_1929,N_2009);
and U2508 (N_2508,N_1860,N_2246);
or U2509 (N_2509,N_1809,N_1842);
nand U2510 (N_2510,N_2220,N_2263);
nor U2511 (N_2511,N_2356,N_2237);
and U2512 (N_2512,N_2096,N_1866);
nand U2513 (N_2513,N_2294,N_1992);
or U2514 (N_2514,N_1891,N_2335);
and U2515 (N_2515,N_2023,N_1850);
and U2516 (N_2516,N_1705,N_2320);
or U2517 (N_2517,N_1619,N_2285);
nor U2518 (N_2518,N_1896,N_1650);
nor U2519 (N_2519,N_1908,N_2352);
and U2520 (N_2520,N_2280,N_1690);
or U2521 (N_2521,N_2222,N_1952);
nor U2522 (N_2522,N_1978,N_2120);
and U2523 (N_2523,N_1723,N_1987);
or U2524 (N_2524,N_2245,N_2210);
nor U2525 (N_2525,N_2208,N_1689);
nand U2526 (N_2526,N_1655,N_2383);
or U2527 (N_2527,N_2125,N_2011);
xnor U2528 (N_2528,N_2232,N_2376);
nor U2529 (N_2529,N_2185,N_1803);
nand U2530 (N_2530,N_1792,N_2386);
or U2531 (N_2531,N_1888,N_2350);
nor U2532 (N_2532,N_2236,N_1932);
nand U2533 (N_2533,N_1865,N_2206);
nand U2534 (N_2534,N_1719,N_1639);
or U2535 (N_2535,N_1642,N_1610);
or U2536 (N_2536,N_1784,N_1972);
nor U2537 (N_2537,N_2082,N_2355);
nand U2538 (N_2538,N_2004,N_2139);
nand U2539 (N_2539,N_2078,N_2176);
and U2540 (N_2540,N_2283,N_1736);
or U2541 (N_2541,N_1867,N_1979);
nor U2542 (N_2542,N_2269,N_2322);
xnor U2543 (N_2543,N_2074,N_1698);
nor U2544 (N_2544,N_1764,N_1806);
xor U2545 (N_2545,N_2147,N_1693);
nand U2546 (N_2546,N_2190,N_2191);
nand U2547 (N_2547,N_1763,N_2113);
and U2548 (N_2548,N_2189,N_1624);
nor U2549 (N_2549,N_1708,N_2346);
nand U2550 (N_2550,N_1678,N_2046);
nor U2551 (N_2551,N_2123,N_2300);
and U2552 (N_2552,N_1823,N_1872);
nand U2553 (N_2553,N_1630,N_1858);
and U2554 (N_2554,N_2053,N_1673);
nand U2555 (N_2555,N_2298,N_1916);
nor U2556 (N_2556,N_2226,N_1906);
nor U2557 (N_2557,N_1717,N_2229);
and U2558 (N_2558,N_1797,N_2302);
nor U2559 (N_2559,N_2396,N_1739);
and U2560 (N_2560,N_2083,N_2171);
and U2561 (N_2561,N_1817,N_2292);
nor U2562 (N_2562,N_2179,N_2274);
nand U2563 (N_2563,N_2070,N_1645);
nor U2564 (N_2564,N_2233,N_1758);
or U2565 (N_2565,N_2344,N_2028);
nor U2566 (N_2566,N_2348,N_2124);
nand U2567 (N_2567,N_2297,N_1728);
or U2568 (N_2568,N_1815,N_1602);
and U2569 (N_2569,N_1629,N_1861);
nor U2570 (N_2570,N_2393,N_1729);
nor U2571 (N_2571,N_2117,N_2020);
nor U2572 (N_2572,N_2062,N_2198);
and U2573 (N_2573,N_1917,N_2130);
or U2574 (N_2574,N_1948,N_2024);
or U2575 (N_2575,N_2173,N_1702);
nor U2576 (N_2576,N_2370,N_2244);
nand U2577 (N_2577,N_2201,N_1800);
nand U2578 (N_2578,N_1894,N_2047);
and U2579 (N_2579,N_1835,N_1679);
or U2580 (N_2580,N_1897,N_1990);
or U2581 (N_2581,N_2034,N_1869);
nor U2582 (N_2582,N_1790,N_2193);
nor U2583 (N_2583,N_1935,N_1715);
nor U2584 (N_2584,N_1772,N_1930);
nand U2585 (N_2585,N_1857,N_2307);
and U2586 (N_2586,N_1965,N_2224);
and U2587 (N_2587,N_2128,N_1838);
nand U2588 (N_2588,N_2397,N_1656);
nand U2589 (N_2589,N_2060,N_2303);
and U2590 (N_2590,N_2036,N_1741);
nor U2591 (N_2591,N_1895,N_2032);
nand U2592 (N_2592,N_2319,N_1749);
and U2593 (N_2593,N_1768,N_1770);
and U2594 (N_2594,N_1802,N_1796);
nand U2595 (N_2595,N_1747,N_2101);
nand U2596 (N_2596,N_1765,N_2369);
or U2597 (N_2597,N_1635,N_2153);
or U2598 (N_2598,N_1646,N_2059);
nand U2599 (N_2599,N_1950,N_1968);
nand U2600 (N_2600,N_1944,N_1604);
or U2601 (N_2601,N_1714,N_2258);
nor U2602 (N_2602,N_1611,N_1634);
nand U2603 (N_2603,N_1625,N_1688);
nor U2604 (N_2604,N_2134,N_1847);
or U2605 (N_2605,N_2168,N_1722);
or U2606 (N_2606,N_1925,N_2234);
nor U2607 (N_2607,N_2090,N_1664);
or U2608 (N_2608,N_1993,N_1721);
nor U2609 (N_2609,N_1949,N_1832);
or U2610 (N_2610,N_1874,N_2072);
or U2611 (N_2611,N_2095,N_1755);
and U2612 (N_2612,N_1605,N_1766);
nor U2613 (N_2613,N_1776,N_1798);
or U2614 (N_2614,N_1680,N_2013);
nand U2615 (N_2615,N_2140,N_1999);
nor U2616 (N_2616,N_2325,N_1709);
or U2617 (N_2617,N_2161,N_2014);
and U2618 (N_2618,N_2239,N_2157);
nand U2619 (N_2619,N_2341,N_2309);
nor U2620 (N_2620,N_2219,N_2162);
and U2621 (N_2621,N_2360,N_1762);
or U2622 (N_2622,N_2000,N_2037);
or U2623 (N_2623,N_1870,N_2377);
nand U2624 (N_2624,N_2146,N_1998);
or U2625 (N_2625,N_2200,N_2166);
nand U2626 (N_2626,N_2266,N_2205);
nand U2627 (N_2627,N_1915,N_1954);
or U2628 (N_2628,N_2315,N_2357);
nor U2629 (N_2629,N_2338,N_1989);
nor U2630 (N_2630,N_2359,N_1887);
nor U2631 (N_2631,N_2092,N_1699);
nor U2632 (N_2632,N_1674,N_1785);
nor U2633 (N_2633,N_1853,N_2094);
or U2634 (N_2634,N_2289,N_2277);
nand U2635 (N_2635,N_2108,N_2031);
nand U2636 (N_2636,N_2182,N_2044);
or U2637 (N_2637,N_1687,N_1851);
and U2638 (N_2638,N_2209,N_1738);
nor U2639 (N_2639,N_1707,N_2389);
or U2640 (N_2640,N_2141,N_1654);
and U2641 (N_2641,N_1834,N_1840);
or U2642 (N_2642,N_1743,N_2093);
nand U2643 (N_2643,N_2337,N_1816);
nor U2644 (N_2644,N_2055,N_1833);
nand U2645 (N_2645,N_2030,N_2121);
or U2646 (N_2646,N_2214,N_2257);
and U2647 (N_2647,N_1672,N_2382);
nand U2648 (N_2648,N_2084,N_2041);
or U2649 (N_2649,N_1778,N_1923);
or U2650 (N_2650,N_2002,N_2167);
and U2651 (N_2651,N_1621,N_2387);
or U2652 (N_2652,N_1885,N_1825);
nand U2653 (N_2653,N_1875,N_2049);
nor U2654 (N_2654,N_2223,N_2230);
nor U2655 (N_2655,N_2152,N_1660);
or U2656 (N_2656,N_2336,N_1671);
and U2657 (N_2657,N_1677,N_1725);
nand U2658 (N_2658,N_2069,N_2282);
nor U2659 (N_2659,N_2254,N_2273);
nor U2660 (N_2660,N_2155,N_2304);
and U2661 (N_2661,N_2243,N_1942);
nor U2662 (N_2662,N_1752,N_1614);
or U2663 (N_2663,N_2247,N_2367);
and U2664 (N_2664,N_2164,N_1706);
and U2665 (N_2665,N_1657,N_1606);
nor U2666 (N_2666,N_2010,N_1730);
or U2667 (N_2667,N_2183,N_2324);
or U2668 (N_2668,N_2231,N_2339);
nor U2669 (N_2669,N_1938,N_1748);
nor U2670 (N_2670,N_2099,N_2363);
or U2671 (N_2671,N_2043,N_1726);
nor U2672 (N_2672,N_1818,N_2116);
nor U2673 (N_2673,N_1881,N_1996);
nand U2674 (N_2674,N_1607,N_2365);
nor U2675 (N_2675,N_2054,N_2265);
nor U2676 (N_2676,N_1667,N_1742);
nand U2677 (N_2677,N_2012,N_1960);
nor U2678 (N_2678,N_2109,N_1883);
nor U2679 (N_2679,N_2035,N_2197);
or U2680 (N_2680,N_1821,N_2284);
or U2681 (N_2681,N_2252,N_1662);
nand U2682 (N_2682,N_2374,N_1740);
nor U2683 (N_2683,N_2371,N_1661);
and U2684 (N_2684,N_1750,N_1926);
and U2685 (N_2685,N_1893,N_1933);
and U2686 (N_2686,N_1771,N_2102);
or U2687 (N_2687,N_1871,N_1774);
or U2688 (N_2688,N_2067,N_1627);
nand U2689 (N_2689,N_1694,N_2313);
and U2690 (N_2690,N_1967,N_1754);
nor U2691 (N_2691,N_1863,N_2115);
or U2692 (N_2692,N_2015,N_1711);
nor U2693 (N_2693,N_2160,N_2066);
nor U2694 (N_2694,N_1886,N_1668);
or U2695 (N_2695,N_1644,N_2075);
and U2696 (N_2696,N_1647,N_1695);
nor U2697 (N_2697,N_1620,N_2068);
nor U2698 (N_2698,N_2328,N_1844);
and U2699 (N_2699,N_1734,N_2281);
nand U2700 (N_2700,N_1712,N_2126);
nor U2701 (N_2701,N_2172,N_1781);
nand U2702 (N_2702,N_2271,N_2163);
nand U2703 (N_2703,N_2196,N_1746);
or U2704 (N_2704,N_2295,N_2156);
nor U2705 (N_2705,N_2235,N_1603);
nor U2706 (N_2706,N_1988,N_1795);
or U2707 (N_2707,N_2195,N_2019);
and U2708 (N_2708,N_1675,N_1940);
or U2709 (N_2709,N_2306,N_2008);
and U2710 (N_2710,N_1852,N_1724);
nand U2711 (N_2711,N_2057,N_2217);
nand U2712 (N_2712,N_1963,N_1843);
xor U2713 (N_2713,N_2385,N_2184);
nor U2714 (N_2714,N_1659,N_1984);
nor U2715 (N_2715,N_1953,N_1757);
nor U2716 (N_2716,N_1637,N_2187);
and U2717 (N_2717,N_1761,N_1981);
nand U2718 (N_2718,N_1830,N_2061);
and U2719 (N_2719,N_2332,N_2181);
nand U2720 (N_2720,N_1601,N_1859);
or U2721 (N_2721,N_1970,N_2203);
nand U2722 (N_2722,N_2275,N_1810);
nand U2723 (N_2723,N_2362,N_1622);
and U2724 (N_2724,N_1753,N_2097);
and U2725 (N_2725,N_2270,N_1946);
nor U2726 (N_2726,N_2278,N_1819);
or U2727 (N_2727,N_1955,N_1745);
or U2728 (N_2728,N_1716,N_1616);
and U2729 (N_2729,N_1848,N_1653);
nor U2730 (N_2730,N_2255,N_2127);
nand U2731 (N_2731,N_1831,N_2276);
or U2732 (N_2732,N_1909,N_1919);
nand U2733 (N_2733,N_1626,N_1910);
or U2734 (N_2734,N_2192,N_1685);
nor U2735 (N_2735,N_2104,N_2207);
nor U2736 (N_2736,N_2142,N_2308);
and U2737 (N_2737,N_2378,N_1973);
nor U2738 (N_2738,N_1826,N_1934);
or U2739 (N_2739,N_1971,N_2118);
and U2740 (N_2740,N_1696,N_1663);
or U2741 (N_2741,N_1732,N_1995);
nor U2742 (N_2742,N_1686,N_1873);
nand U2743 (N_2743,N_1666,N_1609);
nand U2744 (N_2744,N_1876,N_2018);
or U2745 (N_2745,N_2071,N_1879);
and U2746 (N_2746,N_2158,N_1827);
or U2747 (N_2747,N_2017,N_1877);
and U2748 (N_2748,N_1839,N_2174);
nor U2749 (N_2749,N_1976,N_2334);
or U2750 (N_2750,N_2029,N_1904);
or U2751 (N_2751,N_2006,N_1937);
or U2752 (N_2752,N_2296,N_1775);
and U2753 (N_2753,N_1804,N_2025);
nor U2754 (N_2754,N_2261,N_1855);
or U2755 (N_2755,N_1936,N_1921);
or U2756 (N_2756,N_2106,N_2098);
nor U2757 (N_2757,N_1958,N_2379);
and U2758 (N_2758,N_2038,N_1814);
and U2759 (N_2759,N_2149,N_2051);
or U2760 (N_2760,N_1837,N_1836);
nor U2761 (N_2761,N_2040,N_1727);
and U2762 (N_2762,N_1720,N_2375);
or U2763 (N_2763,N_2114,N_2354);
or U2764 (N_2764,N_1862,N_1951);
or U2765 (N_2765,N_1905,N_1733);
nand U2766 (N_2766,N_1713,N_2188);
nand U2767 (N_2767,N_2358,N_1786);
nor U2768 (N_2768,N_2301,N_1903);
and U2769 (N_2769,N_1854,N_2368);
nand U2770 (N_2770,N_1701,N_1682);
nand U2771 (N_2771,N_1974,N_1822);
nand U2772 (N_2772,N_2100,N_2202);
and U2773 (N_2773,N_2133,N_2218);
or U2774 (N_2774,N_1710,N_1665);
nand U2775 (N_2775,N_2388,N_1931);
nand U2776 (N_2776,N_1829,N_1632);
and U2777 (N_2777,N_1658,N_2064);
nor U2778 (N_2778,N_1907,N_2268);
or U2779 (N_2779,N_2260,N_1927);
nor U2780 (N_2780,N_2264,N_1945);
or U2781 (N_2781,N_1751,N_1939);
or U2782 (N_2782,N_2326,N_1773);
or U2783 (N_2783,N_1735,N_2272);
nand U2784 (N_2784,N_2384,N_1759);
or U2785 (N_2785,N_2259,N_2347);
nor U2786 (N_2786,N_1737,N_2177);
and U2787 (N_2787,N_1924,N_2186);
nand U2788 (N_2788,N_1991,N_1731);
or U2789 (N_2789,N_2194,N_1856);
or U2790 (N_2790,N_1820,N_1643);
or U2791 (N_2791,N_2318,N_1892);
and U2792 (N_2792,N_1966,N_2240);
nor U2793 (N_2793,N_1612,N_2148);
nor U2794 (N_2794,N_1769,N_2323);
nand U2795 (N_2795,N_1681,N_1956);
nand U2796 (N_2796,N_2256,N_2287);
nor U2797 (N_2797,N_2279,N_2291);
and U2798 (N_2798,N_2310,N_2112);
or U2799 (N_2799,N_1882,N_2333);
nand U2800 (N_2800,N_2229,N_2383);
nand U2801 (N_2801,N_2285,N_2117);
and U2802 (N_2802,N_2025,N_2293);
nor U2803 (N_2803,N_1945,N_2341);
nor U2804 (N_2804,N_1886,N_1673);
and U2805 (N_2805,N_2365,N_2212);
or U2806 (N_2806,N_2365,N_2034);
nor U2807 (N_2807,N_1981,N_2389);
nor U2808 (N_2808,N_2208,N_1821);
nand U2809 (N_2809,N_2186,N_2288);
or U2810 (N_2810,N_2078,N_1785);
and U2811 (N_2811,N_1844,N_1679);
and U2812 (N_2812,N_1755,N_2042);
nor U2813 (N_2813,N_2195,N_1823);
nand U2814 (N_2814,N_1985,N_2160);
nor U2815 (N_2815,N_2034,N_1660);
nand U2816 (N_2816,N_1647,N_1925);
nand U2817 (N_2817,N_2392,N_2282);
and U2818 (N_2818,N_1787,N_1715);
or U2819 (N_2819,N_2375,N_1921);
and U2820 (N_2820,N_1836,N_1805);
nand U2821 (N_2821,N_1912,N_2141);
and U2822 (N_2822,N_1974,N_2340);
or U2823 (N_2823,N_1669,N_2182);
nand U2824 (N_2824,N_1693,N_2349);
nor U2825 (N_2825,N_1640,N_1842);
nand U2826 (N_2826,N_1852,N_1889);
nand U2827 (N_2827,N_1928,N_1714);
nor U2828 (N_2828,N_1636,N_1972);
nor U2829 (N_2829,N_1871,N_1714);
and U2830 (N_2830,N_2051,N_1749);
or U2831 (N_2831,N_2120,N_2122);
nand U2832 (N_2832,N_1776,N_1679);
nand U2833 (N_2833,N_2159,N_1872);
nor U2834 (N_2834,N_1846,N_2122);
and U2835 (N_2835,N_2254,N_1826);
or U2836 (N_2836,N_2267,N_2316);
nand U2837 (N_2837,N_1968,N_1906);
nor U2838 (N_2838,N_2304,N_2369);
nand U2839 (N_2839,N_2150,N_2104);
nor U2840 (N_2840,N_1977,N_1721);
or U2841 (N_2841,N_1807,N_2122);
and U2842 (N_2842,N_1822,N_1838);
nor U2843 (N_2843,N_2098,N_1680);
nor U2844 (N_2844,N_1817,N_1740);
nor U2845 (N_2845,N_1779,N_2059);
nor U2846 (N_2846,N_1795,N_1705);
or U2847 (N_2847,N_1866,N_2181);
nor U2848 (N_2848,N_2394,N_2189);
and U2849 (N_2849,N_2363,N_2176);
nand U2850 (N_2850,N_1941,N_1991);
and U2851 (N_2851,N_1997,N_1703);
or U2852 (N_2852,N_1797,N_1917);
nor U2853 (N_2853,N_2387,N_2070);
and U2854 (N_2854,N_2051,N_2001);
nand U2855 (N_2855,N_1692,N_2007);
nor U2856 (N_2856,N_1728,N_2033);
and U2857 (N_2857,N_2241,N_2239);
nand U2858 (N_2858,N_1612,N_2314);
and U2859 (N_2859,N_2365,N_2388);
and U2860 (N_2860,N_2195,N_1951);
or U2861 (N_2861,N_2016,N_1681);
or U2862 (N_2862,N_1702,N_1935);
and U2863 (N_2863,N_1987,N_2023);
nand U2864 (N_2864,N_2097,N_2273);
nand U2865 (N_2865,N_2176,N_1645);
or U2866 (N_2866,N_1741,N_2330);
and U2867 (N_2867,N_1976,N_2260);
nor U2868 (N_2868,N_1688,N_1730);
and U2869 (N_2869,N_1664,N_2244);
nor U2870 (N_2870,N_1713,N_2020);
or U2871 (N_2871,N_2374,N_1962);
or U2872 (N_2872,N_2019,N_1772);
xor U2873 (N_2873,N_2227,N_2037);
and U2874 (N_2874,N_2039,N_2307);
or U2875 (N_2875,N_1746,N_1859);
or U2876 (N_2876,N_1671,N_1736);
and U2877 (N_2877,N_1686,N_1979);
nand U2878 (N_2878,N_1988,N_1828);
or U2879 (N_2879,N_2202,N_2155);
or U2880 (N_2880,N_2358,N_2200);
and U2881 (N_2881,N_2036,N_2166);
or U2882 (N_2882,N_1845,N_2361);
nor U2883 (N_2883,N_1873,N_1954);
nand U2884 (N_2884,N_1717,N_1810);
nand U2885 (N_2885,N_1808,N_2059);
or U2886 (N_2886,N_2181,N_2182);
nand U2887 (N_2887,N_2398,N_1711);
nand U2888 (N_2888,N_2268,N_1948);
nor U2889 (N_2889,N_2091,N_1854);
nand U2890 (N_2890,N_1911,N_1635);
nor U2891 (N_2891,N_2134,N_1829);
nor U2892 (N_2892,N_1857,N_2209);
and U2893 (N_2893,N_2153,N_1756);
or U2894 (N_2894,N_1891,N_1677);
and U2895 (N_2895,N_2171,N_2298);
nor U2896 (N_2896,N_2179,N_1894);
nor U2897 (N_2897,N_2095,N_1849);
nand U2898 (N_2898,N_2327,N_2258);
or U2899 (N_2899,N_2155,N_2073);
nand U2900 (N_2900,N_1997,N_1922);
nor U2901 (N_2901,N_1742,N_1942);
nor U2902 (N_2902,N_1997,N_2342);
or U2903 (N_2903,N_1935,N_1956);
and U2904 (N_2904,N_2095,N_1669);
and U2905 (N_2905,N_1835,N_1792);
nand U2906 (N_2906,N_1798,N_1730);
nor U2907 (N_2907,N_1710,N_2219);
or U2908 (N_2908,N_1868,N_2351);
nand U2909 (N_2909,N_2394,N_1690);
and U2910 (N_2910,N_2274,N_1858);
or U2911 (N_2911,N_1739,N_2203);
or U2912 (N_2912,N_1730,N_2068);
nor U2913 (N_2913,N_1771,N_2269);
and U2914 (N_2914,N_2213,N_1930);
nor U2915 (N_2915,N_2115,N_2126);
nor U2916 (N_2916,N_2104,N_2061);
and U2917 (N_2917,N_2086,N_1954);
or U2918 (N_2918,N_1756,N_1870);
nor U2919 (N_2919,N_2359,N_2332);
nand U2920 (N_2920,N_1963,N_2331);
or U2921 (N_2921,N_2306,N_1835);
or U2922 (N_2922,N_1724,N_2065);
nor U2923 (N_2923,N_1915,N_1678);
nor U2924 (N_2924,N_1928,N_2150);
or U2925 (N_2925,N_1971,N_2222);
nand U2926 (N_2926,N_1674,N_1830);
and U2927 (N_2927,N_1800,N_1683);
or U2928 (N_2928,N_1713,N_1725);
or U2929 (N_2929,N_2013,N_2193);
nor U2930 (N_2930,N_1601,N_1799);
nor U2931 (N_2931,N_1947,N_1921);
or U2932 (N_2932,N_2387,N_1841);
nand U2933 (N_2933,N_2340,N_1811);
or U2934 (N_2934,N_2064,N_2143);
nor U2935 (N_2935,N_1841,N_2171);
or U2936 (N_2936,N_2110,N_1693);
nand U2937 (N_2937,N_2200,N_1876);
and U2938 (N_2938,N_2259,N_1766);
or U2939 (N_2939,N_1952,N_2291);
nor U2940 (N_2940,N_2115,N_2304);
and U2941 (N_2941,N_1653,N_1604);
nand U2942 (N_2942,N_1614,N_1937);
nand U2943 (N_2943,N_2243,N_2039);
nand U2944 (N_2944,N_2069,N_2051);
nor U2945 (N_2945,N_1634,N_1883);
and U2946 (N_2946,N_2195,N_2264);
nand U2947 (N_2947,N_1715,N_2381);
and U2948 (N_2948,N_1912,N_1754);
or U2949 (N_2949,N_1798,N_2330);
nand U2950 (N_2950,N_2209,N_1733);
and U2951 (N_2951,N_1653,N_1817);
and U2952 (N_2952,N_2250,N_1838);
and U2953 (N_2953,N_2281,N_1811);
nor U2954 (N_2954,N_2172,N_1871);
or U2955 (N_2955,N_2135,N_1654);
or U2956 (N_2956,N_2280,N_2349);
or U2957 (N_2957,N_2240,N_1770);
nor U2958 (N_2958,N_1837,N_2216);
or U2959 (N_2959,N_2205,N_2053);
nor U2960 (N_2960,N_1909,N_1731);
and U2961 (N_2961,N_1829,N_1950);
nor U2962 (N_2962,N_1616,N_1732);
nor U2963 (N_2963,N_2175,N_2389);
and U2964 (N_2964,N_1775,N_1870);
nor U2965 (N_2965,N_1678,N_1673);
or U2966 (N_2966,N_1954,N_2303);
nor U2967 (N_2967,N_2301,N_2372);
or U2968 (N_2968,N_2083,N_1727);
and U2969 (N_2969,N_2296,N_2170);
nor U2970 (N_2970,N_2378,N_2254);
and U2971 (N_2971,N_2393,N_1943);
nand U2972 (N_2972,N_2214,N_2057);
nand U2973 (N_2973,N_2179,N_1937);
nor U2974 (N_2974,N_2053,N_1839);
xor U2975 (N_2975,N_2224,N_1644);
and U2976 (N_2976,N_1614,N_1772);
nor U2977 (N_2977,N_2326,N_2076);
and U2978 (N_2978,N_2212,N_2327);
xor U2979 (N_2979,N_1861,N_1675);
nor U2980 (N_2980,N_2301,N_1968);
and U2981 (N_2981,N_1669,N_1698);
nand U2982 (N_2982,N_2295,N_2074);
nand U2983 (N_2983,N_1966,N_1894);
nor U2984 (N_2984,N_2197,N_1698);
nor U2985 (N_2985,N_2028,N_1986);
nor U2986 (N_2986,N_2204,N_1821);
nand U2987 (N_2987,N_2095,N_1940);
nand U2988 (N_2988,N_1677,N_2261);
nor U2989 (N_2989,N_1953,N_1897);
nand U2990 (N_2990,N_2354,N_1982);
nand U2991 (N_2991,N_2099,N_2009);
nor U2992 (N_2992,N_1650,N_1850);
nor U2993 (N_2993,N_1644,N_1768);
xnor U2994 (N_2994,N_1900,N_2154);
or U2995 (N_2995,N_1819,N_2335);
nor U2996 (N_2996,N_1706,N_2240);
nand U2997 (N_2997,N_2025,N_2295);
nand U2998 (N_2998,N_2088,N_2191);
or U2999 (N_2999,N_1762,N_1976);
nand U3000 (N_3000,N_1606,N_1933);
nor U3001 (N_3001,N_2075,N_1641);
nor U3002 (N_3002,N_1632,N_1952);
nor U3003 (N_3003,N_1678,N_1738);
nor U3004 (N_3004,N_1708,N_1923);
nand U3005 (N_3005,N_2093,N_1975);
or U3006 (N_3006,N_1632,N_1661);
and U3007 (N_3007,N_1940,N_1727);
nand U3008 (N_3008,N_2084,N_2300);
or U3009 (N_3009,N_2272,N_1901);
nand U3010 (N_3010,N_1847,N_1684);
or U3011 (N_3011,N_1728,N_2260);
or U3012 (N_3012,N_1745,N_1729);
nor U3013 (N_3013,N_2249,N_1735);
nand U3014 (N_3014,N_1919,N_2101);
and U3015 (N_3015,N_1933,N_1854);
nor U3016 (N_3016,N_2361,N_1777);
nand U3017 (N_3017,N_2379,N_2230);
nor U3018 (N_3018,N_2347,N_1666);
nor U3019 (N_3019,N_1907,N_2107);
nor U3020 (N_3020,N_2248,N_2338);
and U3021 (N_3021,N_1897,N_2248);
nor U3022 (N_3022,N_2225,N_1945);
nor U3023 (N_3023,N_2097,N_2290);
or U3024 (N_3024,N_2139,N_1758);
nor U3025 (N_3025,N_1661,N_2187);
nor U3026 (N_3026,N_2349,N_1851);
or U3027 (N_3027,N_1897,N_2092);
and U3028 (N_3028,N_1792,N_2056);
nor U3029 (N_3029,N_1627,N_2398);
nand U3030 (N_3030,N_2059,N_1939);
xnor U3031 (N_3031,N_2351,N_1718);
nor U3032 (N_3032,N_2378,N_2136);
nand U3033 (N_3033,N_1727,N_1846);
nor U3034 (N_3034,N_1993,N_1632);
nor U3035 (N_3035,N_1883,N_1749);
or U3036 (N_3036,N_2241,N_2291);
nor U3037 (N_3037,N_2146,N_1968);
and U3038 (N_3038,N_2355,N_2069);
xor U3039 (N_3039,N_2220,N_1987);
or U3040 (N_3040,N_1885,N_1797);
nand U3041 (N_3041,N_2073,N_1907);
nor U3042 (N_3042,N_2317,N_1745);
nand U3043 (N_3043,N_2001,N_1815);
or U3044 (N_3044,N_1679,N_1837);
nor U3045 (N_3045,N_2212,N_1785);
or U3046 (N_3046,N_1751,N_2078);
nor U3047 (N_3047,N_1842,N_2233);
or U3048 (N_3048,N_2282,N_1658);
and U3049 (N_3049,N_1627,N_1734);
or U3050 (N_3050,N_1703,N_1816);
or U3051 (N_3051,N_2035,N_2389);
and U3052 (N_3052,N_1760,N_1671);
and U3053 (N_3053,N_2202,N_2063);
nor U3054 (N_3054,N_1802,N_1604);
nor U3055 (N_3055,N_2317,N_1688);
or U3056 (N_3056,N_1898,N_2363);
and U3057 (N_3057,N_2027,N_1924);
nor U3058 (N_3058,N_2029,N_1843);
or U3059 (N_3059,N_1884,N_1894);
xor U3060 (N_3060,N_1976,N_2088);
nand U3061 (N_3061,N_1763,N_1603);
or U3062 (N_3062,N_2193,N_1645);
nand U3063 (N_3063,N_1829,N_1641);
and U3064 (N_3064,N_1687,N_1924);
nor U3065 (N_3065,N_1886,N_2162);
nand U3066 (N_3066,N_1871,N_1925);
or U3067 (N_3067,N_2278,N_2355);
or U3068 (N_3068,N_2107,N_2349);
nor U3069 (N_3069,N_1766,N_1990);
or U3070 (N_3070,N_1943,N_2046);
nor U3071 (N_3071,N_2158,N_2377);
and U3072 (N_3072,N_1839,N_1879);
nand U3073 (N_3073,N_1639,N_2129);
or U3074 (N_3074,N_2354,N_1617);
xor U3075 (N_3075,N_1856,N_1757);
nor U3076 (N_3076,N_1732,N_2221);
nand U3077 (N_3077,N_1621,N_1995);
nand U3078 (N_3078,N_1642,N_1866);
and U3079 (N_3079,N_1700,N_1689);
or U3080 (N_3080,N_2179,N_1748);
and U3081 (N_3081,N_2085,N_1718);
nand U3082 (N_3082,N_2353,N_2074);
or U3083 (N_3083,N_1834,N_2127);
nor U3084 (N_3084,N_1893,N_2074);
and U3085 (N_3085,N_2058,N_1706);
nor U3086 (N_3086,N_2069,N_2382);
nand U3087 (N_3087,N_1952,N_1763);
and U3088 (N_3088,N_1751,N_2028);
and U3089 (N_3089,N_2239,N_1790);
nand U3090 (N_3090,N_1955,N_2331);
nand U3091 (N_3091,N_2167,N_2020);
and U3092 (N_3092,N_1929,N_1977);
and U3093 (N_3093,N_2057,N_1628);
nand U3094 (N_3094,N_2199,N_2010);
and U3095 (N_3095,N_1953,N_1877);
nor U3096 (N_3096,N_2256,N_1675);
or U3097 (N_3097,N_2303,N_1755);
and U3098 (N_3098,N_1932,N_1639);
or U3099 (N_3099,N_2246,N_1664);
and U3100 (N_3100,N_1898,N_1696);
and U3101 (N_3101,N_2207,N_2260);
nor U3102 (N_3102,N_2175,N_2253);
nor U3103 (N_3103,N_1637,N_2217);
nand U3104 (N_3104,N_2132,N_1926);
or U3105 (N_3105,N_1808,N_1775);
nor U3106 (N_3106,N_1665,N_2286);
or U3107 (N_3107,N_2039,N_1924);
or U3108 (N_3108,N_2249,N_1847);
or U3109 (N_3109,N_1670,N_2146);
nand U3110 (N_3110,N_1657,N_2048);
and U3111 (N_3111,N_2112,N_2012);
and U3112 (N_3112,N_1690,N_1803);
nand U3113 (N_3113,N_2065,N_2219);
nor U3114 (N_3114,N_2238,N_2199);
or U3115 (N_3115,N_2243,N_1706);
or U3116 (N_3116,N_2302,N_1907);
nor U3117 (N_3117,N_2337,N_2079);
nor U3118 (N_3118,N_2087,N_2194);
nor U3119 (N_3119,N_2361,N_2183);
nor U3120 (N_3120,N_1796,N_1678);
xor U3121 (N_3121,N_1946,N_2387);
or U3122 (N_3122,N_2080,N_2093);
or U3123 (N_3123,N_2270,N_1709);
nor U3124 (N_3124,N_1943,N_2019);
and U3125 (N_3125,N_2398,N_1944);
nor U3126 (N_3126,N_1722,N_1818);
nor U3127 (N_3127,N_1883,N_1879);
xor U3128 (N_3128,N_2222,N_1918);
nor U3129 (N_3129,N_1673,N_1634);
and U3130 (N_3130,N_1651,N_2088);
nand U3131 (N_3131,N_2135,N_2165);
nor U3132 (N_3132,N_2278,N_2307);
nor U3133 (N_3133,N_1912,N_2394);
or U3134 (N_3134,N_2278,N_2045);
or U3135 (N_3135,N_2374,N_2234);
nor U3136 (N_3136,N_1683,N_1902);
or U3137 (N_3137,N_2270,N_2250);
nand U3138 (N_3138,N_2391,N_1972);
nor U3139 (N_3139,N_1722,N_2025);
nor U3140 (N_3140,N_1936,N_1855);
and U3141 (N_3141,N_1831,N_1894);
or U3142 (N_3142,N_1975,N_1668);
nand U3143 (N_3143,N_2045,N_1906);
nand U3144 (N_3144,N_1719,N_1676);
nand U3145 (N_3145,N_1647,N_1911);
nand U3146 (N_3146,N_2073,N_2126);
and U3147 (N_3147,N_2171,N_2039);
or U3148 (N_3148,N_2395,N_2295);
and U3149 (N_3149,N_2238,N_1866);
nor U3150 (N_3150,N_2159,N_1882);
xnor U3151 (N_3151,N_2308,N_1730);
nor U3152 (N_3152,N_1786,N_2227);
and U3153 (N_3153,N_1701,N_2287);
or U3154 (N_3154,N_1755,N_2211);
or U3155 (N_3155,N_1701,N_2022);
nand U3156 (N_3156,N_2196,N_1907);
or U3157 (N_3157,N_2024,N_1978);
and U3158 (N_3158,N_1623,N_2081);
nor U3159 (N_3159,N_2373,N_1651);
nand U3160 (N_3160,N_1673,N_2262);
and U3161 (N_3161,N_2050,N_2053);
nor U3162 (N_3162,N_1799,N_2272);
nor U3163 (N_3163,N_1931,N_2048);
or U3164 (N_3164,N_2307,N_2042);
or U3165 (N_3165,N_1667,N_2044);
or U3166 (N_3166,N_2081,N_2039);
and U3167 (N_3167,N_2393,N_1970);
and U3168 (N_3168,N_2305,N_2227);
nand U3169 (N_3169,N_2219,N_1871);
or U3170 (N_3170,N_2178,N_1710);
and U3171 (N_3171,N_2387,N_2399);
nor U3172 (N_3172,N_1606,N_1766);
nand U3173 (N_3173,N_2225,N_2294);
or U3174 (N_3174,N_2324,N_2094);
or U3175 (N_3175,N_1920,N_2269);
and U3176 (N_3176,N_2130,N_2117);
nand U3177 (N_3177,N_2397,N_2006);
nor U3178 (N_3178,N_1762,N_1602);
nand U3179 (N_3179,N_1993,N_1889);
and U3180 (N_3180,N_2384,N_1641);
or U3181 (N_3181,N_2100,N_2122);
or U3182 (N_3182,N_2092,N_1786);
and U3183 (N_3183,N_2379,N_1999);
or U3184 (N_3184,N_1961,N_2171);
and U3185 (N_3185,N_1949,N_2169);
and U3186 (N_3186,N_1886,N_1608);
nand U3187 (N_3187,N_1663,N_1916);
or U3188 (N_3188,N_1853,N_2089);
nor U3189 (N_3189,N_2336,N_1867);
nand U3190 (N_3190,N_2028,N_2257);
nand U3191 (N_3191,N_2070,N_1947);
and U3192 (N_3192,N_2018,N_2384);
xnor U3193 (N_3193,N_1816,N_1667);
and U3194 (N_3194,N_1771,N_2206);
xnor U3195 (N_3195,N_1604,N_2300);
or U3196 (N_3196,N_2266,N_2286);
and U3197 (N_3197,N_2325,N_1840);
or U3198 (N_3198,N_1848,N_2363);
or U3199 (N_3199,N_2284,N_1745);
nor U3200 (N_3200,N_2886,N_2738);
or U3201 (N_3201,N_2732,N_2621);
and U3202 (N_3202,N_3117,N_2848);
and U3203 (N_3203,N_2747,N_2505);
nor U3204 (N_3204,N_3168,N_2903);
or U3205 (N_3205,N_2553,N_2824);
nand U3206 (N_3206,N_2658,N_3094);
nor U3207 (N_3207,N_2464,N_3030);
or U3208 (N_3208,N_2499,N_2922);
and U3209 (N_3209,N_2831,N_2742);
nor U3210 (N_3210,N_2841,N_2737);
nand U3211 (N_3211,N_2457,N_3010);
and U3212 (N_3212,N_2497,N_2483);
or U3213 (N_3213,N_3006,N_2911);
or U3214 (N_3214,N_2984,N_3143);
nand U3215 (N_3215,N_2432,N_3134);
nand U3216 (N_3216,N_2489,N_2863);
nor U3217 (N_3217,N_3160,N_2468);
nand U3218 (N_3218,N_2525,N_3183);
or U3219 (N_3219,N_2630,N_2754);
xnor U3220 (N_3220,N_2818,N_3068);
or U3221 (N_3221,N_2555,N_2588);
nand U3222 (N_3222,N_3036,N_3179);
nor U3223 (N_3223,N_3028,N_2511);
nand U3224 (N_3224,N_2615,N_3079);
or U3225 (N_3225,N_3163,N_3098);
nor U3226 (N_3226,N_2982,N_2961);
nor U3227 (N_3227,N_2673,N_2939);
nand U3228 (N_3228,N_3164,N_2513);
nor U3229 (N_3229,N_2437,N_2977);
or U3230 (N_3230,N_2444,N_2484);
nand U3231 (N_3231,N_3108,N_3085);
nor U3232 (N_3232,N_2461,N_2563);
nand U3233 (N_3233,N_2800,N_2427);
or U3234 (N_3234,N_2685,N_2634);
and U3235 (N_3235,N_2814,N_3007);
nand U3236 (N_3236,N_2642,N_3195);
or U3237 (N_3237,N_2589,N_3138);
or U3238 (N_3238,N_2493,N_2907);
nor U3239 (N_3239,N_2893,N_2807);
and U3240 (N_3240,N_2959,N_2908);
nand U3241 (N_3241,N_2935,N_3105);
nand U3242 (N_3242,N_3084,N_2676);
and U3243 (N_3243,N_3073,N_2775);
nand U3244 (N_3244,N_2606,N_3186);
or U3245 (N_3245,N_2920,N_2500);
and U3246 (N_3246,N_2998,N_2750);
nor U3247 (N_3247,N_2622,N_3058);
nor U3248 (N_3248,N_3170,N_3121);
nand U3249 (N_3249,N_2610,N_3037);
nor U3250 (N_3250,N_2633,N_2593);
and U3251 (N_3251,N_2986,N_3092);
and U3252 (N_3252,N_2845,N_2929);
or U3253 (N_3253,N_2751,N_2960);
or U3254 (N_3254,N_2828,N_2717);
nor U3255 (N_3255,N_2956,N_3193);
and U3256 (N_3256,N_2520,N_2646);
nand U3257 (N_3257,N_2569,N_2561);
or U3258 (N_3258,N_2704,N_2504);
nor U3259 (N_3259,N_2546,N_2657);
or U3260 (N_3260,N_3124,N_2957);
nand U3261 (N_3261,N_2867,N_3054);
or U3262 (N_3262,N_2411,N_3038);
xnor U3263 (N_3263,N_2554,N_3070);
nor U3264 (N_3264,N_3076,N_3145);
nand U3265 (N_3265,N_2441,N_2989);
or U3266 (N_3266,N_2875,N_2502);
or U3267 (N_3267,N_2883,N_3180);
nor U3268 (N_3268,N_2729,N_2844);
and U3269 (N_3269,N_2476,N_2482);
nand U3270 (N_3270,N_2522,N_2906);
nand U3271 (N_3271,N_2644,N_2995);
nand U3272 (N_3272,N_3057,N_2643);
and U3273 (N_3273,N_2470,N_2709);
or U3274 (N_3274,N_3154,N_2774);
or U3275 (N_3275,N_2506,N_2971);
nand U3276 (N_3276,N_3078,N_2746);
xnor U3277 (N_3277,N_2947,N_2650);
nor U3278 (N_3278,N_3133,N_2528);
nand U3279 (N_3279,N_2452,N_2614);
xor U3280 (N_3280,N_2869,N_3115);
nand U3281 (N_3281,N_3018,N_2762);
nor U3282 (N_3282,N_2462,N_2779);
nand U3283 (N_3283,N_2933,N_3005);
or U3284 (N_3284,N_2877,N_2696);
and U3285 (N_3285,N_2888,N_2976);
nand U3286 (N_3286,N_2429,N_2575);
and U3287 (N_3287,N_3106,N_2790);
nor U3288 (N_3288,N_2519,N_3026);
nand U3289 (N_3289,N_2594,N_2735);
nand U3290 (N_3290,N_2759,N_2764);
nand U3291 (N_3291,N_2940,N_2878);
or U3292 (N_3292,N_2892,N_2983);
nor U3293 (N_3293,N_3104,N_2787);
nand U3294 (N_3294,N_3009,N_2937);
and U3295 (N_3295,N_3102,N_2412);
nor U3296 (N_3296,N_2866,N_3136);
and U3297 (N_3297,N_2918,N_2994);
and U3298 (N_3298,N_2993,N_2916);
or U3299 (N_3299,N_2455,N_3065);
nor U3300 (N_3300,N_2778,N_2475);
and U3301 (N_3301,N_2765,N_2486);
and U3302 (N_3302,N_2661,N_2856);
and U3303 (N_3303,N_2469,N_2474);
nand U3304 (N_3304,N_3110,N_2549);
nor U3305 (N_3305,N_2805,N_3047);
nor U3306 (N_3306,N_2636,N_2722);
or U3307 (N_3307,N_2900,N_2923);
or U3308 (N_3308,N_3161,N_2773);
nand U3309 (N_3309,N_2819,N_2958);
nor U3310 (N_3310,N_2910,N_3112);
and U3311 (N_3311,N_2527,N_3033);
nor U3312 (N_3312,N_2966,N_2731);
nor U3313 (N_3313,N_2946,N_2855);
and U3314 (N_3314,N_2660,N_2419);
or U3315 (N_3315,N_2820,N_2739);
and U3316 (N_3316,N_2537,N_2840);
nand U3317 (N_3317,N_3192,N_2625);
nor U3318 (N_3318,N_2585,N_2400);
nor U3319 (N_3319,N_2967,N_2620);
nand U3320 (N_3320,N_2424,N_2656);
or U3321 (N_3321,N_3199,N_2882);
or U3322 (N_3322,N_2689,N_3130);
or U3323 (N_3323,N_2487,N_3017);
nand U3324 (N_3324,N_2955,N_2899);
nand U3325 (N_3325,N_2712,N_2627);
xor U3326 (N_3326,N_2683,N_2703);
and U3327 (N_3327,N_2843,N_2822);
or U3328 (N_3328,N_2928,N_3191);
or U3329 (N_3329,N_3126,N_2975);
nand U3330 (N_3330,N_2826,N_2686);
nor U3331 (N_3331,N_2458,N_3155);
nor U3332 (N_3332,N_2401,N_2943);
and U3333 (N_3333,N_2490,N_3188);
and U3334 (N_3334,N_2577,N_2491);
nand U3335 (N_3335,N_2770,N_2952);
nand U3336 (N_3336,N_2838,N_2426);
nand U3337 (N_3337,N_2420,N_2927);
and U3338 (N_3338,N_2782,N_3116);
and U3339 (N_3339,N_3091,N_2980);
or U3340 (N_3340,N_2654,N_3120);
nor U3341 (N_3341,N_2926,N_2969);
or U3342 (N_3342,N_2439,N_2786);
and U3343 (N_3343,N_2416,N_2748);
and U3344 (N_3344,N_2783,N_2868);
and U3345 (N_3345,N_2410,N_3069);
nand U3346 (N_3346,N_2972,N_2635);
nand U3347 (N_3347,N_2485,N_2815);
and U3348 (N_3348,N_2640,N_2618);
and U3349 (N_3349,N_2433,N_2453);
or U3350 (N_3350,N_2430,N_3067);
and U3351 (N_3351,N_3063,N_2626);
nor U3352 (N_3352,N_2551,N_2478);
nor U3353 (N_3353,N_2789,N_3041);
nor U3354 (N_3354,N_2571,N_2645);
and U3355 (N_3355,N_3197,N_2719);
nand U3356 (N_3356,N_2873,N_2827);
and U3357 (N_3357,N_2586,N_2930);
nand U3358 (N_3358,N_2707,N_2812);
and U3359 (N_3359,N_2481,N_2521);
and U3360 (N_3360,N_2752,N_3083);
nand U3361 (N_3361,N_2604,N_3146);
nand U3362 (N_3362,N_2798,N_3128);
or U3363 (N_3363,N_2792,N_2564);
and U3364 (N_3364,N_2725,N_2694);
nand U3365 (N_3365,N_3049,N_2898);
nor U3366 (N_3366,N_3086,N_3175);
and U3367 (N_3367,N_2817,N_3074);
nor U3368 (N_3368,N_2498,N_2587);
xnor U3369 (N_3369,N_2407,N_2896);
nand U3370 (N_3370,N_2858,N_2945);
and U3371 (N_3371,N_2727,N_2545);
or U3372 (N_3372,N_3035,N_2700);
nor U3373 (N_3373,N_2755,N_2954);
nor U3374 (N_3374,N_2756,N_3149);
or U3375 (N_3375,N_2950,N_2757);
and U3376 (N_3376,N_2876,N_2842);
or U3377 (N_3377,N_2602,N_2723);
or U3378 (N_3378,N_2990,N_2881);
or U3379 (N_3379,N_2591,N_2699);
and U3380 (N_3380,N_2810,N_2825);
or U3381 (N_3381,N_3165,N_2417);
and U3382 (N_3382,N_2510,N_3118);
and U3383 (N_3383,N_3046,N_2578);
and U3384 (N_3384,N_2421,N_2936);
and U3385 (N_3385,N_2523,N_2821);
nor U3386 (N_3386,N_2864,N_2816);
nor U3387 (N_3387,N_2582,N_3023);
or U3388 (N_3388,N_2418,N_3196);
nor U3389 (N_3389,N_3189,N_3013);
nor U3390 (N_3390,N_2772,N_2999);
nand U3391 (N_3391,N_2833,N_2413);
or U3392 (N_3392,N_2605,N_3034);
nand U3393 (N_3393,N_3184,N_2665);
and U3394 (N_3394,N_2434,N_2508);
nand U3395 (N_3395,N_2785,N_2509);
or U3396 (N_3396,N_2663,N_2583);
and U3397 (N_3397,N_2566,N_2889);
and U3398 (N_3398,N_3150,N_3148);
and U3399 (N_3399,N_2613,N_2579);
nand U3400 (N_3400,N_2953,N_3159);
or U3401 (N_3401,N_2733,N_2865);
or U3402 (N_3402,N_2791,N_2557);
or U3403 (N_3403,N_2607,N_3080);
nor U3404 (N_3404,N_2891,N_2542);
nand U3405 (N_3405,N_2574,N_2897);
or U3406 (N_3406,N_2720,N_2580);
nor U3407 (N_3407,N_2516,N_2668);
nand U3408 (N_3408,N_2612,N_2973);
or U3409 (N_3409,N_2802,N_2496);
nand U3410 (N_3410,N_2598,N_2674);
or U3411 (N_3411,N_2619,N_2596);
and U3412 (N_3412,N_2771,N_2526);
nand U3413 (N_3413,N_2690,N_2862);
or U3414 (N_3414,N_2649,N_3119);
and U3415 (N_3415,N_3114,N_2595);
or U3416 (N_3416,N_2492,N_2501);
nor U3417 (N_3417,N_2985,N_2761);
and U3418 (N_3418,N_2988,N_3055);
and U3419 (N_3419,N_3187,N_3052);
or U3420 (N_3420,N_2403,N_2987);
nor U3421 (N_3421,N_3088,N_2978);
or U3422 (N_3422,N_3002,N_3066);
or U3423 (N_3423,N_2544,N_3181);
xor U3424 (N_3424,N_2541,N_2617);
or U3425 (N_3425,N_2652,N_3031);
or U3426 (N_3426,N_3096,N_2647);
nor U3427 (N_3427,N_2423,N_2533);
or U3428 (N_3428,N_2438,N_3100);
nor U3429 (N_3429,N_2550,N_2447);
or U3430 (N_3430,N_2885,N_2599);
or U3431 (N_3431,N_3172,N_2964);
and U3432 (N_3432,N_3051,N_2415);
or U3433 (N_3433,N_3095,N_3107);
nand U3434 (N_3434,N_3093,N_2488);
nor U3435 (N_3435,N_2965,N_2446);
nand U3436 (N_3436,N_2749,N_2616);
or U3437 (N_3437,N_2758,N_3061);
and U3438 (N_3438,N_2473,N_2666);
or U3439 (N_3439,N_2846,N_3198);
and U3440 (N_3440,N_2466,N_2835);
nor U3441 (N_3441,N_3027,N_2874);
or U3442 (N_3442,N_3153,N_2472);
nand U3443 (N_3443,N_2721,N_2479);
or U3444 (N_3444,N_2861,N_2670);
and U3445 (N_3445,N_2776,N_2829);
and U3446 (N_3446,N_2912,N_3000);
nor U3447 (N_3447,N_2548,N_2451);
or U3448 (N_3448,N_2693,N_2655);
and U3449 (N_3449,N_2839,N_2901);
or U3450 (N_3450,N_2780,N_2968);
or U3451 (N_3451,N_2781,N_3015);
nor U3452 (N_3452,N_2795,N_2706);
xor U3453 (N_3453,N_2408,N_2796);
or U3454 (N_3454,N_3053,N_2543);
and U3455 (N_3455,N_3012,N_2924);
nor U3456 (N_3456,N_2671,N_2871);
or U3457 (N_3457,N_2456,N_3129);
nor U3458 (N_3458,N_2440,N_3132);
and U3459 (N_3459,N_2974,N_2979);
or U3460 (N_3460,N_2465,N_3060);
or U3461 (N_3461,N_2409,N_3185);
or U3462 (N_3462,N_3082,N_2743);
nor U3463 (N_3463,N_3166,N_2480);
nand U3464 (N_3464,N_2879,N_2672);
or U3465 (N_3465,N_3139,N_2951);
or U3466 (N_3466,N_2887,N_2857);
nor U3467 (N_3467,N_2823,N_2431);
and U3468 (N_3468,N_2809,N_2450);
nor U3469 (N_3469,N_2405,N_2422);
and U3470 (N_3470,N_2837,N_2777);
nand U3471 (N_3471,N_2449,N_2714);
or U3472 (N_3472,N_3142,N_2734);
nand U3473 (N_3473,N_2463,N_2745);
and U3474 (N_3474,N_2531,N_2797);
and U3475 (N_3475,N_3123,N_3004);
nand U3476 (N_3476,N_3162,N_2547);
and U3477 (N_3477,N_2859,N_2851);
nor U3478 (N_3478,N_2904,N_3090);
nand U3479 (N_3479,N_3025,N_3024);
and U3480 (N_3480,N_3048,N_2556);
xnor U3481 (N_3481,N_2870,N_3056);
or U3482 (N_3482,N_2705,N_2894);
or U3483 (N_3483,N_2890,N_3178);
nand U3484 (N_3484,N_3151,N_2530);
nand U3485 (N_3485,N_2684,N_2808);
nand U3486 (N_3486,N_2942,N_2648);
and U3487 (N_3487,N_3087,N_2702);
nand U3488 (N_3488,N_3043,N_2836);
nand U3489 (N_3489,N_2559,N_2536);
or U3490 (N_3490,N_2552,N_2507);
nand U3491 (N_3491,N_3174,N_2949);
or U3492 (N_3492,N_2597,N_2425);
or U3493 (N_3493,N_2406,N_2806);
or U3494 (N_3494,N_3089,N_2801);
nand U3495 (N_3495,N_2641,N_3194);
nand U3496 (N_3496,N_3050,N_2629);
nor U3497 (N_3497,N_3157,N_2692);
and U3498 (N_3498,N_2662,N_2695);
and U3499 (N_3499,N_3099,N_2584);
nor U3500 (N_3500,N_2850,N_2915);
nand U3501 (N_3501,N_2688,N_2623);
nand U3502 (N_3502,N_2515,N_2766);
nor U3503 (N_3503,N_3062,N_2460);
or U3504 (N_3504,N_3039,N_2996);
and U3505 (N_3505,N_2728,N_2414);
or U3506 (N_3506,N_2639,N_2560);
or U3507 (N_3507,N_2849,N_3077);
nand U3508 (N_3508,N_2697,N_2736);
and U3509 (N_3509,N_3011,N_2428);
and U3510 (N_3510,N_3003,N_2562);
and U3511 (N_3511,N_3140,N_2651);
nor U3512 (N_3512,N_2494,N_2963);
nor U3513 (N_3513,N_3171,N_2445);
nand U3514 (N_3514,N_2667,N_2794);
and U3515 (N_3515,N_2852,N_2948);
nor U3516 (N_3516,N_2512,N_3173);
and U3517 (N_3517,N_2603,N_2803);
nor U3518 (N_3518,N_2740,N_2535);
nor U3519 (N_3519,N_2799,N_2628);
or U3520 (N_3520,N_2471,N_2675);
or U3521 (N_3521,N_2934,N_2788);
nor U3522 (N_3522,N_3019,N_3176);
and U3523 (N_3523,N_3147,N_2679);
nand U3524 (N_3524,N_2880,N_2919);
nor U3525 (N_3525,N_2708,N_2724);
and U3526 (N_3526,N_2730,N_2611);
xnor U3527 (N_3527,N_3001,N_2970);
or U3528 (N_3528,N_2710,N_3075);
or U3529 (N_3529,N_2534,N_3081);
and U3530 (N_3530,N_2711,N_2435);
and U3531 (N_3531,N_3131,N_2454);
or U3532 (N_3532,N_2830,N_2631);
nand U3533 (N_3533,N_2701,N_2726);
and U3534 (N_3534,N_2677,N_2570);
xor U3535 (N_3535,N_3167,N_2941);
and U3536 (N_3536,N_2608,N_2698);
nor U3537 (N_3537,N_2592,N_2436);
and U3538 (N_3538,N_3152,N_3016);
nand U3539 (N_3539,N_2914,N_2590);
and U3540 (N_3540,N_2517,N_3040);
nor U3541 (N_3541,N_3109,N_2529);
and U3542 (N_3542,N_2687,N_2902);
or U3543 (N_3543,N_2576,N_3182);
or U3544 (N_3544,N_3064,N_2518);
nand U3545 (N_3545,N_3122,N_3156);
and U3546 (N_3546,N_3111,N_2637);
nor U3547 (N_3547,N_2909,N_2669);
nor U3548 (N_3548,N_3137,N_2741);
nor U3549 (N_3549,N_3097,N_3044);
nand U3550 (N_3550,N_2997,N_2691);
nor U3551 (N_3551,N_2448,N_2600);
or U3552 (N_3552,N_2467,N_3029);
or U3553 (N_3553,N_2632,N_2784);
nor U3554 (N_3554,N_2834,N_2459);
or U3555 (N_3555,N_3072,N_2753);
or U3556 (N_3556,N_2847,N_3071);
or U3557 (N_3557,N_2503,N_2678);
or U3558 (N_3558,N_2913,N_2477);
nor U3559 (N_3559,N_2832,N_2514);
or U3560 (N_3560,N_2539,N_2917);
nand U3561 (N_3561,N_2682,N_2715);
nand U3562 (N_3562,N_3141,N_2853);
and U3563 (N_3563,N_2568,N_2905);
or U3564 (N_3564,N_3177,N_2638);
and U3565 (N_3565,N_2558,N_2581);
nor U3566 (N_3566,N_3144,N_2767);
and U3567 (N_3567,N_3125,N_3022);
nor U3568 (N_3568,N_2962,N_3059);
or U3569 (N_3569,N_2872,N_2925);
nor U3570 (N_3570,N_2854,N_2404);
and U3571 (N_3571,N_2402,N_2981);
or U3572 (N_3572,N_2495,N_2932);
nor U3573 (N_3573,N_3045,N_2992);
and U3574 (N_3574,N_3190,N_3158);
and U3575 (N_3575,N_2938,N_3103);
nand U3576 (N_3576,N_3127,N_2931);
or U3577 (N_3577,N_2921,N_2760);
and U3578 (N_3578,N_2664,N_2680);
or U3579 (N_3579,N_2769,N_3032);
nor U3580 (N_3580,N_2768,N_3021);
nand U3581 (N_3581,N_2532,N_3008);
nor U3582 (N_3582,N_2860,N_3014);
or U3583 (N_3583,N_2718,N_2538);
and U3584 (N_3584,N_2713,N_2884);
nand U3585 (N_3585,N_2895,N_3169);
nor U3586 (N_3586,N_2716,N_2609);
nor U3587 (N_3587,N_2811,N_2572);
nand U3588 (N_3588,N_2804,N_2744);
and U3589 (N_3589,N_2565,N_2601);
or U3590 (N_3590,N_3135,N_2681);
nand U3591 (N_3591,N_3042,N_2763);
or U3592 (N_3592,N_2524,N_3020);
or U3593 (N_3593,N_2653,N_2443);
and U3594 (N_3594,N_2813,N_2793);
nand U3595 (N_3595,N_2944,N_2659);
xor U3596 (N_3596,N_2567,N_2624);
nor U3597 (N_3597,N_2442,N_2573);
nand U3598 (N_3598,N_2540,N_3113);
nor U3599 (N_3599,N_3101,N_2991);
xnor U3600 (N_3600,N_3148,N_3044);
or U3601 (N_3601,N_3177,N_2688);
nor U3602 (N_3602,N_2863,N_3063);
or U3603 (N_3603,N_2682,N_2872);
xnor U3604 (N_3604,N_2856,N_2547);
or U3605 (N_3605,N_2593,N_2637);
nor U3606 (N_3606,N_2907,N_2770);
or U3607 (N_3607,N_2716,N_2655);
and U3608 (N_3608,N_2447,N_2764);
or U3609 (N_3609,N_2642,N_2508);
and U3610 (N_3610,N_3081,N_2545);
nand U3611 (N_3611,N_2840,N_3107);
or U3612 (N_3612,N_3193,N_2936);
nor U3613 (N_3613,N_3017,N_2781);
or U3614 (N_3614,N_2560,N_2528);
and U3615 (N_3615,N_2997,N_2798);
nor U3616 (N_3616,N_2842,N_2709);
nor U3617 (N_3617,N_2874,N_2787);
nor U3618 (N_3618,N_3112,N_2438);
xnor U3619 (N_3619,N_2726,N_2548);
nand U3620 (N_3620,N_2645,N_2436);
nand U3621 (N_3621,N_2761,N_2675);
nor U3622 (N_3622,N_3011,N_3128);
and U3623 (N_3623,N_2957,N_2484);
nand U3624 (N_3624,N_2857,N_2754);
and U3625 (N_3625,N_2607,N_2926);
and U3626 (N_3626,N_2796,N_2563);
nand U3627 (N_3627,N_2802,N_2531);
nand U3628 (N_3628,N_3128,N_2849);
nand U3629 (N_3629,N_2958,N_2427);
and U3630 (N_3630,N_3076,N_2819);
and U3631 (N_3631,N_2489,N_3184);
or U3632 (N_3632,N_3103,N_3045);
and U3633 (N_3633,N_2595,N_2905);
and U3634 (N_3634,N_2476,N_2547);
xor U3635 (N_3635,N_2851,N_3009);
nor U3636 (N_3636,N_2974,N_2711);
nor U3637 (N_3637,N_2931,N_3085);
nand U3638 (N_3638,N_2476,N_3167);
nand U3639 (N_3639,N_3066,N_3156);
nor U3640 (N_3640,N_2757,N_2980);
nand U3641 (N_3641,N_2999,N_2786);
and U3642 (N_3642,N_2531,N_2772);
nor U3643 (N_3643,N_3171,N_2708);
nand U3644 (N_3644,N_2421,N_2873);
nand U3645 (N_3645,N_3151,N_2439);
or U3646 (N_3646,N_3131,N_3190);
or U3647 (N_3647,N_3172,N_2464);
nand U3648 (N_3648,N_2758,N_3070);
and U3649 (N_3649,N_2538,N_3045);
and U3650 (N_3650,N_3122,N_2965);
nand U3651 (N_3651,N_2519,N_2803);
and U3652 (N_3652,N_2598,N_3172);
or U3653 (N_3653,N_2948,N_2807);
and U3654 (N_3654,N_2983,N_2609);
nor U3655 (N_3655,N_2531,N_2866);
nand U3656 (N_3656,N_3137,N_3024);
nand U3657 (N_3657,N_2622,N_2401);
nor U3658 (N_3658,N_3062,N_3104);
nand U3659 (N_3659,N_2763,N_3137);
or U3660 (N_3660,N_3016,N_2843);
and U3661 (N_3661,N_2888,N_2804);
and U3662 (N_3662,N_3059,N_2547);
or U3663 (N_3663,N_2907,N_2977);
nand U3664 (N_3664,N_3019,N_2628);
or U3665 (N_3665,N_2867,N_2961);
or U3666 (N_3666,N_2440,N_2634);
or U3667 (N_3667,N_3085,N_3019);
nor U3668 (N_3668,N_2689,N_2515);
and U3669 (N_3669,N_2711,N_2698);
nand U3670 (N_3670,N_2839,N_2767);
and U3671 (N_3671,N_3123,N_2603);
and U3672 (N_3672,N_3180,N_3160);
nor U3673 (N_3673,N_2833,N_2789);
or U3674 (N_3674,N_2614,N_2707);
nand U3675 (N_3675,N_2495,N_2404);
nand U3676 (N_3676,N_3137,N_3188);
nand U3677 (N_3677,N_3138,N_2608);
nor U3678 (N_3678,N_2419,N_2717);
and U3679 (N_3679,N_2703,N_2663);
and U3680 (N_3680,N_2464,N_2709);
nand U3681 (N_3681,N_2867,N_2800);
nor U3682 (N_3682,N_2871,N_3188);
and U3683 (N_3683,N_3139,N_2730);
or U3684 (N_3684,N_2985,N_2979);
nand U3685 (N_3685,N_3143,N_2611);
or U3686 (N_3686,N_2747,N_3072);
or U3687 (N_3687,N_2529,N_2655);
nor U3688 (N_3688,N_3157,N_2724);
nand U3689 (N_3689,N_3130,N_3150);
or U3690 (N_3690,N_2466,N_2483);
nand U3691 (N_3691,N_3183,N_3158);
or U3692 (N_3692,N_3188,N_2830);
or U3693 (N_3693,N_2741,N_2945);
and U3694 (N_3694,N_2968,N_2664);
nor U3695 (N_3695,N_2583,N_2535);
nor U3696 (N_3696,N_2997,N_2746);
nand U3697 (N_3697,N_3069,N_2498);
and U3698 (N_3698,N_2981,N_2976);
nor U3699 (N_3699,N_3052,N_2475);
or U3700 (N_3700,N_2663,N_2524);
or U3701 (N_3701,N_2666,N_2941);
nand U3702 (N_3702,N_2897,N_2596);
nor U3703 (N_3703,N_2503,N_2848);
nand U3704 (N_3704,N_2527,N_2806);
or U3705 (N_3705,N_3013,N_2430);
nand U3706 (N_3706,N_2762,N_2453);
nand U3707 (N_3707,N_2534,N_2894);
nand U3708 (N_3708,N_3142,N_2527);
nand U3709 (N_3709,N_2673,N_2987);
nand U3710 (N_3710,N_2986,N_2858);
nand U3711 (N_3711,N_2523,N_2831);
nor U3712 (N_3712,N_2753,N_3098);
nor U3713 (N_3713,N_2653,N_2673);
and U3714 (N_3714,N_2507,N_3089);
and U3715 (N_3715,N_2950,N_3004);
nor U3716 (N_3716,N_3019,N_2838);
nor U3717 (N_3717,N_2580,N_2697);
and U3718 (N_3718,N_2853,N_2581);
or U3719 (N_3719,N_2730,N_2795);
nand U3720 (N_3720,N_3158,N_2629);
xnor U3721 (N_3721,N_3074,N_2777);
or U3722 (N_3722,N_2884,N_3181);
nor U3723 (N_3723,N_2482,N_2960);
nand U3724 (N_3724,N_2457,N_3079);
and U3725 (N_3725,N_2748,N_2975);
and U3726 (N_3726,N_2707,N_2494);
nand U3727 (N_3727,N_2946,N_2967);
or U3728 (N_3728,N_2561,N_2898);
and U3729 (N_3729,N_3074,N_2736);
or U3730 (N_3730,N_2406,N_2581);
or U3731 (N_3731,N_2851,N_2564);
and U3732 (N_3732,N_2456,N_2978);
or U3733 (N_3733,N_2570,N_3011);
and U3734 (N_3734,N_3129,N_2606);
xnor U3735 (N_3735,N_2793,N_2967);
and U3736 (N_3736,N_2939,N_3010);
nor U3737 (N_3737,N_2637,N_2920);
or U3738 (N_3738,N_3002,N_2622);
and U3739 (N_3739,N_2447,N_2629);
nand U3740 (N_3740,N_2565,N_2422);
and U3741 (N_3741,N_2778,N_2997);
nor U3742 (N_3742,N_3191,N_2868);
and U3743 (N_3743,N_3104,N_2734);
nor U3744 (N_3744,N_2746,N_3111);
or U3745 (N_3745,N_3053,N_2568);
nand U3746 (N_3746,N_2450,N_2949);
nor U3747 (N_3747,N_3142,N_3016);
xor U3748 (N_3748,N_2575,N_2678);
and U3749 (N_3749,N_2687,N_3115);
or U3750 (N_3750,N_3161,N_2923);
nor U3751 (N_3751,N_2881,N_3060);
nor U3752 (N_3752,N_3197,N_2947);
nor U3753 (N_3753,N_2928,N_2871);
and U3754 (N_3754,N_3129,N_3038);
or U3755 (N_3755,N_2818,N_2647);
and U3756 (N_3756,N_2863,N_3119);
and U3757 (N_3757,N_3032,N_2835);
nor U3758 (N_3758,N_2552,N_2700);
nor U3759 (N_3759,N_3131,N_2567);
and U3760 (N_3760,N_2953,N_2578);
and U3761 (N_3761,N_2832,N_2699);
nand U3762 (N_3762,N_2517,N_2912);
xnor U3763 (N_3763,N_3159,N_2789);
nor U3764 (N_3764,N_3108,N_2881);
nand U3765 (N_3765,N_2511,N_2512);
or U3766 (N_3766,N_2880,N_3024);
or U3767 (N_3767,N_3103,N_2563);
nand U3768 (N_3768,N_2537,N_3036);
and U3769 (N_3769,N_3107,N_3084);
nor U3770 (N_3770,N_2989,N_2575);
and U3771 (N_3771,N_2413,N_2928);
nand U3772 (N_3772,N_2682,N_3062);
nand U3773 (N_3773,N_2593,N_3182);
nand U3774 (N_3774,N_3174,N_3124);
and U3775 (N_3775,N_3077,N_2923);
or U3776 (N_3776,N_2477,N_2708);
nand U3777 (N_3777,N_2562,N_2911);
xnor U3778 (N_3778,N_3190,N_2571);
and U3779 (N_3779,N_2878,N_3133);
nor U3780 (N_3780,N_2441,N_3058);
nor U3781 (N_3781,N_2945,N_2747);
nand U3782 (N_3782,N_2653,N_2910);
or U3783 (N_3783,N_2817,N_2525);
nor U3784 (N_3784,N_2970,N_2765);
and U3785 (N_3785,N_3116,N_2914);
nor U3786 (N_3786,N_2538,N_2638);
and U3787 (N_3787,N_3160,N_2950);
nand U3788 (N_3788,N_2535,N_3156);
nor U3789 (N_3789,N_2632,N_2616);
nand U3790 (N_3790,N_3189,N_2431);
nand U3791 (N_3791,N_2645,N_3018);
nand U3792 (N_3792,N_2817,N_2777);
nand U3793 (N_3793,N_2890,N_2746);
or U3794 (N_3794,N_2809,N_2980);
nor U3795 (N_3795,N_2713,N_2831);
nand U3796 (N_3796,N_3020,N_2420);
or U3797 (N_3797,N_2916,N_2602);
or U3798 (N_3798,N_2686,N_2688);
nor U3799 (N_3799,N_2657,N_2560);
or U3800 (N_3800,N_2413,N_2743);
nand U3801 (N_3801,N_2428,N_2487);
and U3802 (N_3802,N_2613,N_2448);
nor U3803 (N_3803,N_2465,N_2934);
and U3804 (N_3804,N_2570,N_2736);
and U3805 (N_3805,N_3008,N_3187);
nand U3806 (N_3806,N_2996,N_2890);
nor U3807 (N_3807,N_2834,N_2623);
nand U3808 (N_3808,N_3144,N_3101);
or U3809 (N_3809,N_2785,N_3115);
and U3810 (N_3810,N_3183,N_2906);
nor U3811 (N_3811,N_2761,N_2832);
and U3812 (N_3812,N_3163,N_3010);
nor U3813 (N_3813,N_2986,N_2637);
nor U3814 (N_3814,N_2993,N_2712);
or U3815 (N_3815,N_2880,N_2971);
and U3816 (N_3816,N_3168,N_2691);
and U3817 (N_3817,N_3160,N_3021);
or U3818 (N_3818,N_2448,N_2913);
and U3819 (N_3819,N_2967,N_3044);
or U3820 (N_3820,N_2565,N_2734);
and U3821 (N_3821,N_2534,N_2517);
nor U3822 (N_3822,N_3069,N_2665);
and U3823 (N_3823,N_2924,N_3176);
or U3824 (N_3824,N_2647,N_2850);
and U3825 (N_3825,N_2954,N_3059);
nor U3826 (N_3826,N_3189,N_2762);
nand U3827 (N_3827,N_2666,N_3085);
or U3828 (N_3828,N_2934,N_2972);
and U3829 (N_3829,N_2460,N_2595);
nor U3830 (N_3830,N_2456,N_2704);
nor U3831 (N_3831,N_2882,N_3080);
and U3832 (N_3832,N_2440,N_2956);
nand U3833 (N_3833,N_2655,N_2919);
nand U3834 (N_3834,N_2681,N_2787);
nor U3835 (N_3835,N_2856,N_2733);
or U3836 (N_3836,N_2669,N_2812);
nand U3837 (N_3837,N_2910,N_2816);
and U3838 (N_3838,N_3061,N_2621);
nor U3839 (N_3839,N_2832,N_3091);
nor U3840 (N_3840,N_3015,N_2675);
nand U3841 (N_3841,N_2594,N_3024);
nand U3842 (N_3842,N_3175,N_3145);
or U3843 (N_3843,N_2403,N_2768);
nand U3844 (N_3844,N_3056,N_2435);
or U3845 (N_3845,N_3095,N_2528);
nand U3846 (N_3846,N_3135,N_3123);
or U3847 (N_3847,N_2442,N_2864);
or U3848 (N_3848,N_2741,N_2460);
or U3849 (N_3849,N_2584,N_2876);
nand U3850 (N_3850,N_2598,N_2751);
and U3851 (N_3851,N_3089,N_3103);
and U3852 (N_3852,N_2418,N_2924);
nor U3853 (N_3853,N_2577,N_2493);
or U3854 (N_3854,N_3177,N_2840);
nand U3855 (N_3855,N_2999,N_2434);
nand U3856 (N_3856,N_3052,N_2933);
nand U3857 (N_3857,N_2464,N_3153);
and U3858 (N_3858,N_2724,N_2639);
nor U3859 (N_3859,N_3135,N_3193);
nor U3860 (N_3860,N_2764,N_2682);
nor U3861 (N_3861,N_3023,N_2619);
nand U3862 (N_3862,N_2554,N_2814);
and U3863 (N_3863,N_2912,N_2540);
nor U3864 (N_3864,N_3090,N_2517);
or U3865 (N_3865,N_3007,N_2741);
xor U3866 (N_3866,N_2718,N_3113);
nor U3867 (N_3867,N_2734,N_2682);
nand U3868 (N_3868,N_2743,N_2925);
nor U3869 (N_3869,N_2519,N_2860);
and U3870 (N_3870,N_2466,N_3126);
or U3871 (N_3871,N_2447,N_2529);
nand U3872 (N_3872,N_3131,N_2904);
and U3873 (N_3873,N_2884,N_2646);
nor U3874 (N_3874,N_2535,N_2468);
nand U3875 (N_3875,N_2657,N_2975);
and U3876 (N_3876,N_3186,N_2919);
nand U3877 (N_3877,N_2890,N_3038);
and U3878 (N_3878,N_2871,N_2457);
nor U3879 (N_3879,N_2728,N_2765);
nand U3880 (N_3880,N_2647,N_3029);
or U3881 (N_3881,N_2521,N_2830);
or U3882 (N_3882,N_3063,N_2807);
nand U3883 (N_3883,N_3003,N_3102);
or U3884 (N_3884,N_2929,N_2607);
or U3885 (N_3885,N_2836,N_2850);
or U3886 (N_3886,N_2930,N_2552);
and U3887 (N_3887,N_2436,N_3072);
nor U3888 (N_3888,N_3115,N_3091);
or U3889 (N_3889,N_2955,N_2516);
and U3890 (N_3890,N_2409,N_2840);
and U3891 (N_3891,N_2922,N_2852);
nor U3892 (N_3892,N_3007,N_2468);
or U3893 (N_3893,N_2555,N_2568);
nand U3894 (N_3894,N_2714,N_2420);
or U3895 (N_3895,N_3098,N_3139);
nor U3896 (N_3896,N_2906,N_2632);
nand U3897 (N_3897,N_3125,N_2713);
and U3898 (N_3898,N_2482,N_3105);
nand U3899 (N_3899,N_2737,N_2976);
or U3900 (N_3900,N_2961,N_2695);
and U3901 (N_3901,N_2534,N_3110);
and U3902 (N_3902,N_3026,N_2514);
nand U3903 (N_3903,N_3153,N_2750);
nand U3904 (N_3904,N_2948,N_2594);
xor U3905 (N_3905,N_3062,N_2860);
and U3906 (N_3906,N_3091,N_2590);
nor U3907 (N_3907,N_3141,N_2859);
and U3908 (N_3908,N_3120,N_3148);
or U3909 (N_3909,N_3094,N_3070);
and U3910 (N_3910,N_2416,N_3184);
nor U3911 (N_3911,N_2823,N_2733);
or U3912 (N_3912,N_2901,N_2553);
and U3913 (N_3913,N_3094,N_2774);
or U3914 (N_3914,N_2891,N_2541);
nand U3915 (N_3915,N_2615,N_3193);
and U3916 (N_3916,N_2615,N_2630);
nor U3917 (N_3917,N_2435,N_2740);
and U3918 (N_3918,N_2888,N_3032);
or U3919 (N_3919,N_2679,N_2867);
nor U3920 (N_3920,N_2574,N_3169);
and U3921 (N_3921,N_2683,N_3054);
nor U3922 (N_3922,N_2928,N_2842);
nand U3923 (N_3923,N_2543,N_2957);
or U3924 (N_3924,N_2595,N_2579);
nand U3925 (N_3925,N_2430,N_2523);
nor U3926 (N_3926,N_3153,N_3109);
and U3927 (N_3927,N_2479,N_2766);
or U3928 (N_3928,N_2419,N_2598);
nor U3929 (N_3929,N_2520,N_2855);
nand U3930 (N_3930,N_2673,N_2950);
nand U3931 (N_3931,N_2968,N_2933);
nor U3932 (N_3932,N_2895,N_2893);
or U3933 (N_3933,N_2771,N_2769);
and U3934 (N_3934,N_2707,N_3013);
and U3935 (N_3935,N_2650,N_3195);
nand U3936 (N_3936,N_2958,N_2913);
and U3937 (N_3937,N_2659,N_2560);
nor U3938 (N_3938,N_2789,N_2578);
or U3939 (N_3939,N_2822,N_2434);
and U3940 (N_3940,N_3103,N_3163);
or U3941 (N_3941,N_2867,N_3132);
or U3942 (N_3942,N_3199,N_3004);
or U3943 (N_3943,N_2539,N_2718);
xnor U3944 (N_3944,N_3180,N_2621);
nor U3945 (N_3945,N_3098,N_3159);
and U3946 (N_3946,N_2840,N_2816);
or U3947 (N_3947,N_2643,N_3079);
and U3948 (N_3948,N_3125,N_3066);
xor U3949 (N_3949,N_3086,N_2460);
nand U3950 (N_3950,N_2831,N_2837);
and U3951 (N_3951,N_2810,N_2952);
nor U3952 (N_3952,N_2477,N_2603);
nand U3953 (N_3953,N_3177,N_2880);
nor U3954 (N_3954,N_3081,N_2485);
nor U3955 (N_3955,N_2826,N_2777);
nand U3956 (N_3956,N_2631,N_2408);
or U3957 (N_3957,N_2503,N_2658);
or U3958 (N_3958,N_2780,N_2924);
nand U3959 (N_3959,N_3186,N_2471);
nor U3960 (N_3960,N_2401,N_2415);
nor U3961 (N_3961,N_2494,N_2737);
nor U3962 (N_3962,N_3169,N_2470);
xor U3963 (N_3963,N_2408,N_3148);
and U3964 (N_3964,N_2785,N_2424);
nand U3965 (N_3965,N_3066,N_2430);
nor U3966 (N_3966,N_2460,N_2747);
and U3967 (N_3967,N_3170,N_2907);
and U3968 (N_3968,N_2907,N_2516);
or U3969 (N_3969,N_2500,N_2740);
or U3970 (N_3970,N_3038,N_2630);
nor U3971 (N_3971,N_2594,N_2931);
and U3972 (N_3972,N_2700,N_2648);
nor U3973 (N_3973,N_3067,N_3040);
or U3974 (N_3974,N_2626,N_2798);
nor U3975 (N_3975,N_2486,N_2974);
or U3976 (N_3976,N_2980,N_2424);
and U3977 (N_3977,N_2645,N_2504);
and U3978 (N_3978,N_2854,N_2511);
or U3979 (N_3979,N_3135,N_3198);
and U3980 (N_3980,N_2753,N_3140);
nand U3981 (N_3981,N_2544,N_2821);
and U3982 (N_3982,N_2768,N_2624);
or U3983 (N_3983,N_2698,N_3166);
or U3984 (N_3984,N_2526,N_2713);
or U3985 (N_3985,N_2558,N_2570);
nand U3986 (N_3986,N_2828,N_2911);
and U3987 (N_3987,N_2470,N_2683);
and U3988 (N_3988,N_2657,N_2581);
nor U3989 (N_3989,N_2412,N_2460);
or U3990 (N_3990,N_2741,N_2586);
or U3991 (N_3991,N_2973,N_2724);
nand U3992 (N_3992,N_2467,N_2871);
nand U3993 (N_3993,N_3160,N_2921);
nor U3994 (N_3994,N_3035,N_2580);
nor U3995 (N_3995,N_2713,N_2903);
and U3996 (N_3996,N_3188,N_2806);
nand U3997 (N_3997,N_3051,N_2647);
nand U3998 (N_3998,N_2942,N_2564);
and U3999 (N_3999,N_3142,N_2956);
nand U4000 (N_4000,N_3345,N_3683);
and U4001 (N_4001,N_3652,N_3281);
nor U4002 (N_4002,N_3508,N_3850);
or U4003 (N_4003,N_3504,N_3638);
or U4004 (N_4004,N_3763,N_3323);
nor U4005 (N_4005,N_3496,N_3677);
nand U4006 (N_4006,N_3516,N_3482);
nand U4007 (N_4007,N_3915,N_3995);
nor U4008 (N_4008,N_3484,N_3996);
and U4009 (N_4009,N_3497,N_3834);
nor U4010 (N_4010,N_3548,N_3353);
nand U4011 (N_4011,N_3424,N_3234);
and U4012 (N_4012,N_3208,N_3705);
nand U4013 (N_4013,N_3700,N_3619);
and U4014 (N_4014,N_3520,N_3667);
nand U4015 (N_4015,N_3313,N_3576);
nand U4016 (N_4016,N_3750,N_3434);
nor U4017 (N_4017,N_3493,N_3852);
nand U4018 (N_4018,N_3775,N_3556);
and U4019 (N_4019,N_3807,N_3615);
nand U4020 (N_4020,N_3620,N_3416);
nand U4021 (N_4021,N_3495,N_3490);
nor U4022 (N_4022,N_3384,N_3499);
nor U4023 (N_4023,N_3542,N_3918);
or U4024 (N_4024,N_3610,N_3747);
or U4025 (N_4025,N_3588,N_3832);
or U4026 (N_4026,N_3465,N_3488);
nand U4027 (N_4027,N_3579,N_3571);
nor U4028 (N_4028,N_3304,N_3535);
or U4029 (N_4029,N_3803,N_3238);
nand U4030 (N_4030,N_3794,N_3317);
nor U4031 (N_4031,N_3798,N_3987);
or U4032 (N_4032,N_3716,N_3528);
or U4033 (N_4033,N_3557,N_3373);
nor U4034 (N_4034,N_3280,N_3975);
or U4035 (N_4035,N_3336,N_3882);
nand U4036 (N_4036,N_3779,N_3252);
or U4037 (N_4037,N_3917,N_3367);
or U4038 (N_4038,N_3724,N_3818);
or U4039 (N_4039,N_3318,N_3637);
and U4040 (N_4040,N_3876,N_3358);
or U4041 (N_4041,N_3693,N_3210);
nor U4042 (N_4042,N_3746,N_3892);
nand U4043 (N_4043,N_3645,N_3942);
nor U4044 (N_4044,N_3671,N_3228);
nand U4045 (N_4045,N_3951,N_3214);
or U4046 (N_4046,N_3733,N_3697);
nor U4047 (N_4047,N_3333,N_3563);
or U4048 (N_4048,N_3607,N_3532);
nand U4049 (N_4049,N_3346,N_3360);
nor U4050 (N_4050,N_3522,N_3795);
or U4051 (N_4051,N_3659,N_3331);
and U4052 (N_4052,N_3782,N_3821);
and U4053 (N_4053,N_3586,N_3498);
nor U4054 (N_4054,N_3564,N_3463);
and U4055 (N_4055,N_3405,N_3853);
or U4056 (N_4056,N_3663,N_3829);
or U4057 (N_4057,N_3666,N_3748);
nand U4058 (N_4058,N_3558,N_3344);
nand U4059 (N_4059,N_3787,N_3608);
xnor U4060 (N_4060,N_3978,N_3617);
nand U4061 (N_4061,N_3738,N_3453);
or U4062 (N_4062,N_3765,N_3276);
nor U4063 (N_4063,N_3526,N_3397);
and U4064 (N_4064,N_3656,N_3560);
or U4065 (N_4065,N_3991,N_3236);
or U4066 (N_4066,N_3785,N_3898);
nand U4067 (N_4067,N_3849,N_3545);
or U4068 (N_4068,N_3664,N_3739);
nor U4069 (N_4069,N_3525,N_3591);
nand U4070 (N_4070,N_3613,N_3896);
or U4071 (N_4071,N_3639,N_3540);
nor U4072 (N_4072,N_3814,N_3992);
nand U4073 (N_4073,N_3534,N_3854);
nor U4074 (N_4074,N_3875,N_3438);
nor U4075 (N_4075,N_3552,N_3362);
and U4076 (N_4076,N_3772,N_3809);
nand U4077 (N_4077,N_3768,N_3261);
nor U4078 (N_4078,N_3893,N_3343);
nor U4079 (N_4079,N_3606,N_3900);
or U4080 (N_4080,N_3451,N_3941);
or U4081 (N_4081,N_3783,N_3519);
or U4082 (N_4082,N_3710,N_3206);
or U4083 (N_4083,N_3272,N_3887);
nand U4084 (N_4084,N_3650,N_3403);
nor U4085 (N_4085,N_3521,N_3931);
nand U4086 (N_4086,N_3396,N_3725);
and U4087 (N_4087,N_3865,N_3695);
nor U4088 (N_4088,N_3267,N_3417);
or U4089 (N_4089,N_3582,N_3474);
nand U4090 (N_4090,N_3209,N_3847);
or U4091 (N_4091,N_3948,N_3611);
or U4092 (N_4092,N_3956,N_3481);
nand U4093 (N_4093,N_3366,N_3347);
or U4094 (N_4094,N_3904,N_3365);
nand U4095 (N_4095,N_3432,N_3329);
xor U4096 (N_4096,N_3780,N_3550);
nor U4097 (N_4097,N_3623,N_3997);
or U4098 (N_4098,N_3225,N_3324);
nand U4099 (N_4099,N_3791,N_3943);
or U4100 (N_4100,N_3503,N_3801);
or U4101 (N_4101,N_3910,N_3229);
and U4102 (N_4102,N_3311,N_3784);
and U4103 (N_4103,N_3622,N_3927);
and U4104 (N_4104,N_3250,N_3665);
nand U4105 (N_4105,N_3593,N_3433);
xnor U4106 (N_4106,N_3502,N_3653);
and U4107 (N_4107,N_3407,N_3744);
or U4108 (N_4108,N_3934,N_3492);
nand U4109 (N_4109,N_3570,N_3300);
nand U4110 (N_4110,N_3937,N_3573);
nor U4111 (N_4111,N_3448,N_3858);
nor U4112 (N_4112,N_3844,N_3673);
and U4113 (N_4113,N_3627,N_3647);
or U4114 (N_4114,N_3726,N_3719);
nand U4115 (N_4115,N_3328,N_3295);
or U4116 (N_4116,N_3761,N_3421);
or U4117 (N_4117,N_3246,N_3363);
or U4118 (N_4118,N_3518,N_3636);
nor U4119 (N_4119,N_3444,N_3305);
or U4120 (N_4120,N_3441,N_3709);
and U4121 (N_4121,N_3413,N_3699);
nand U4122 (N_4122,N_3599,N_3804);
nor U4123 (N_4123,N_3303,N_3544);
nand U4124 (N_4124,N_3901,N_3201);
xnor U4125 (N_4125,N_3480,N_3885);
nor U4126 (N_4126,N_3958,N_3897);
nand U4127 (N_4127,N_3269,N_3342);
and U4128 (N_4128,N_3376,N_3501);
or U4129 (N_4129,N_3530,N_3781);
or U4130 (N_4130,N_3813,N_3741);
or U4131 (N_4131,N_3730,N_3307);
nor U4132 (N_4132,N_3301,N_3868);
nor U4133 (N_4133,N_3754,N_3967);
nand U4134 (N_4134,N_3551,N_3979);
nor U4135 (N_4135,N_3972,N_3831);
nand U4136 (N_4136,N_3988,N_3728);
or U4137 (N_4137,N_3239,N_3878);
or U4138 (N_4138,N_3398,N_3477);
or U4139 (N_4139,N_3812,N_3965);
nand U4140 (N_4140,N_3760,N_3378);
nor U4141 (N_4141,N_3604,N_3450);
nand U4142 (N_4142,N_3793,N_3790);
nand U4143 (N_4143,N_3447,N_3660);
or U4144 (N_4144,N_3263,N_3762);
nor U4145 (N_4145,N_3436,N_3428);
and U4146 (N_4146,N_3568,N_3734);
and U4147 (N_4147,N_3288,N_3251);
nand U4148 (N_4148,N_3479,N_3316);
nor U4149 (N_4149,N_3751,N_3980);
nor U4150 (N_4150,N_3543,N_3335);
and U4151 (N_4151,N_3283,N_3952);
nand U4152 (N_4152,N_3833,N_3701);
or U4153 (N_4153,N_3856,N_3869);
nand U4154 (N_4154,N_3439,N_3240);
nand U4155 (N_4155,N_3386,N_3233);
nor U4156 (N_4156,N_3581,N_3265);
nand U4157 (N_4157,N_3810,N_3609);
or U4158 (N_4158,N_3629,N_3392);
and U4159 (N_4159,N_3412,N_3402);
and U4160 (N_4160,N_3302,N_3224);
or U4161 (N_4161,N_3248,N_3533);
nor U4162 (N_4162,N_3583,N_3244);
or U4163 (N_4163,N_3736,N_3703);
and U4164 (N_4164,N_3939,N_3322);
and U4165 (N_4165,N_3862,N_3334);
nand U4166 (N_4166,N_3387,N_3855);
or U4167 (N_4167,N_3954,N_3422);
and U4168 (N_4168,N_3848,N_3879);
and U4169 (N_4169,N_3889,N_3601);
nor U4170 (N_4170,N_3685,N_3907);
nand U4171 (N_4171,N_3430,N_3391);
and U4172 (N_4172,N_3668,N_3555);
nand U4173 (N_4173,N_3680,N_3921);
nor U4174 (N_4174,N_3237,N_3640);
or U4175 (N_4175,N_3735,N_3830);
and U4176 (N_4176,N_3310,N_3870);
or U4177 (N_4177,N_3674,N_3319);
or U4178 (N_4178,N_3511,N_3899);
nand U4179 (N_4179,N_3565,N_3827);
and U4180 (N_4180,N_3936,N_3688);
or U4181 (N_4181,N_3908,N_3971);
nor U4182 (N_4182,N_3976,N_3257);
or U4183 (N_4183,N_3932,N_3625);
nand U4184 (N_4184,N_3999,N_3815);
or U4185 (N_4185,N_3415,N_3286);
xor U4186 (N_4186,N_3510,N_3994);
nand U4187 (N_4187,N_3602,N_3580);
nor U4188 (N_4188,N_3443,N_3561);
or U4189 (N_4189,N_3213,N_3471);
nor U4190 (N_4190,N_3903,N_3399);
nor U4191 (N_4191,N_3454,N_3473);
or U4192 (N_4192,N_3634,N_3420);
nor U4193 (N_4193,N_3644,N_3370);
nor U4194 (N_4194,N_3461,N_3431);
nand U4195 (N_4195,N_3249,N_3678);
xor U4196 (N_4196,N_3618,N_3478);
nand U4197 (N_4197,N_3633,N_3773);
nand U4198 (N_4198,N_3788,N_3863);
or U4199 (N_4199,N_3905,N_3590);
or U4200 (N_4200,N_3986,N_3717);
and U4201 (N_4201,N_3486,N_3946);
nand U4202 (N_4202,N_3388,N_3745);
and U4203 (N_4203,N_3374,N_3554);
or U4204 (N_4204,N_3714,N_3840);
and U4205 (N_4205,N_3817,N_3449);
and U4206 (N_4206,N_3916,N_3825);
and U4207 (N_4207,N_3694,N_3361);
and U4208 (N_4208,N_3594,N_3977);
and U4209 (N_4209,N_3395,N_3711);
or U4210 (N_4210,N_3727,N_3872);
nor U4211 (N_4211,N_3457,N_3642);
nor U4212 (N_4212,N_3381,N_3340);
or U4213 (N_4213,N_3955,N_3802);
and U4214 (N_4214,N_3820,N_3427);
nor U4215 (N_4215,N_3553,N_3274);
nor U4216 (N_4216,N_3506,N_3296);
nor U4217 (N_4217,N_3839,N_3982);
and U4218 (N_4218,N_3458,N_3846);
nand U4219 (N_4219,N_3983,N_3891);
and U4220 (N_4220,N_3669,N_3949);
nand U4221 (N_4221,N_3969,N_3860);
or U4222 (N_4222,N_3299,N_3874);
nand U4223 (N_4223,N_3749,N_3587);
or U4224 (N_4224,N_3349,N_3658);
nand U4225 (N_4225,N_3414,N_3468);
or U4226 (N_4226,N_3217,N_3922);
and U4227 (N_4227,N_3824,N_3718);
xnor U4228 (N_4228,N_3298,N_3256);
and U4229 (N_4229,N_3293,N_3743);
nor U4230 (N_4230,N_3966,N_3359);
nor U4231 (N_4231,N_3989,N_3616);
and U4232 (N_4232,N_3585,N_3805);
nand U4233 (N_4233,N_3828,N_3321);
or U4234 (N_4234,N_3327,N_3306);
or U4235 (N_4235,N_3445,N_3753);
or U4236 (N_4236,N_3512,N_3375);
nand U4237 (N_4237,N_3687,N_3740);
or U4238 (N_4238,N_3819,N_3757);
nand U4239 (N_4239,N_3411,N_3984);
nand U4240 (N_4240,N_3758,N_3963);
nand U4241 (N_4241,N_3686,N_3935);
or U4242 (N_4242,N_3584,N_3940);
and U4243 (N_4243,N_3938,N_3998);
nor U4244 (N_4244,N_3404,N_3462);
nor U4245 (N_4245,N_3626,N_3212);
and U4246 (N_4246,N_3559,N_3843);
and U4247 (N_4247,N_3309,N_3221);
nor U4248 (N_4248,N_3547,N_3778);
and U4249 (N_4249,N_3595,N_3628);
and U4250 (N_4250,N_3429,N_3837);
and U4251 (N_4251,N_3270,N_3655);
and U4252 (N_4252,N_3575,N_3348);
nor U4253 (N_4253,N_3401,N_3389);
nand U4254 (N_4254,N_3871,N_3993);
nand U4255 (N_4255,N_3377,N_3207);
nand U4256 (N_4256,N_3646,N_3215);
nor U4257 (N_4257,N_3483,N_3676);
or U4258 (N_4258,N_3661,N_3235);
nand U4259 (N_4259,N_3467,N_3247);
and U4260 (N_4260,N_3792,N_3877);
xor U4261 (N_4261,N_3258,N_3596);
and U4262 (N_4262,N_3764,N_3895);
nor U4263 (N_4263,N_3278,N_3435);
or U4264 (N_4264,N_3851,N_3767);
or U4265 (N_4265,N_3418,N_3308);
nand U4266 (N_4266,N_3867,N_3704);
nor U4267 (N_4267,N_3243,N_3385);
nor U4268 (N_4268,N_3888,N_3797);
nand U4269 (N_4269,N_3312,N_3505);
nand U4270 (N_4270,N_3369,N_3964);
nand U4271 (N_4271,N_3919,N_3379);
nor U4272 (N_4272,N_3672,N_3913);
nand U4273 (N_4273,N_3538,N_3929);
or U4274 (N_4274,N_3230,N_3702);
or U4275 (N_4275,N_3489,N_3253);
or U4276 (N_4276,N_3605,N_3408);
xnor U4277 (N_4277,N_3771,N_3220);
nand U4278 (N_4278,N_3475,N_3894);
nor U4279 (N_4279,N_3950,N_3957);
nand U4280 (N_4280,N_3287,N_3691);
or U4281 (N_4281,N_3393,N_3372);
nand U4282 (N_4282,N_3406,N_3974);
nand U4283 (N_4283,N_3341,N_3670);
nor U4284 (N_4284,N_3279,N_3657);
nand U4285 (N_4285,N_3861,N_3339);
and U4286 (N_4286,N_3513,N_3866);
and U4287 (N_4287,N_3826,N_3721);
xnor U4288 (N_4288,N_3924,N_3314);
nor U4289 (N_4289,N_3800,N_3284);
and U4290 (N_4290,N_3291,N_3789);
nand U4291 (N_4291,N_3715,N_3507);
and U4292 (N_4292,N_3752,N_3546);
and U4293 (N_4293,N_3643,N_3260);
and U4294 (N_4294,N_3944,N_3320);
nor U4295 (N_4295,N_3271,N_3460);
nor U4296 (N_4296,N_3442,N_3631);
or U4297 (N_4297,N_3524,N_3600);
and U4298 (N_4298,N_3566,N_3696);
nor U4299 (N_4299,N_3682,N_3732);
nand U4300 (N_4300,N_3419,N_3902);
and U4301 (N_4301,N_3597,N_3297);
nor U4302 (N_4302,N_3290,N_3592);
and U4303 (N_4303,N_3226,N_3689);
and U4304 (N_4304,N_3662,N_3472);
or U4305 (N_4305,N_3383,N_3731);
nor U4306 (N_4306,N_3205,N_3452);
nor U4307 (N_4307,N_3737,N_3242);
nor U4308 (N_4308,N_3254,N_3338);
nand U4309 (N_4309,N_3612,N_3681);
and U4310 (N_4310,N_3960,N_3961);
or U4311 (N_4311,N_3883,N_3536);
or U4312 (N_4312,N_3835,N_3985);
and U4313 (N_4313,N_3509,N_3933);
xor U4314 (N_4314,N_3273,N_3811);
nand U4315 (N_4315,N_3218,N_3569);
and U4316 (N_4316,N_3410,N_3864);
and U4317 (N_4317,N_3541,N_3884);
or U4318 (N_4318,N_3945,N_3337);
nand U4319 (N_4319,N_3523,N_3285);
nand U4320 (N_4320,N_3836,N_3262);
nand U4321 (N_4321,N_3776,N_3466);
or U4322 (N_4322,N_3470,N_3911);
and U4323 (N_4323,N_3351,N_3822);
and U4324 (N_4324,N_3517,N_3264);
nor U4325 (N_4325,N_3589,N_3423);
nand U4326 (N_4326,N_3906,N_3742);
and U4327 (N_4327,N_3712,N_3537);
or U4328 (N_4328,N_3690,N_3970);
nand U4329 (N_4329,N_3614,N_3574);
or U4330 (N_4330,N_3920,N_3890);
or U4331 (N_4331,N_3294,N_3603);
nor U4332 (N_4332,N_3953,N_3227);
or U4333 (N_4333,N_3368,N_3756);
nand U4334 (N_4334,N_3531,N_3514);
or U4335 (N_4335,N_3223,N_3654);
nor U4336 (N_4336,N_3487,N_3766);
and U4337 (N_4337,N_3491,N_3873);
or U4338 (N_4338,N_3881,N_3382);
and U4339 (N_4339,N_3857,N_3909);
nor U4340 (N_4340,N_3292,N_3332);
or U4341 (N_4341,N_3231,N_3759);
or U4342 (N_4342,N_3354,N_3713);
or U4343 (N_4343,N_3371,N_3706);
or U4344 (N_4344,N_3926,N_3315);
or U4345 (N_4345,N_3440,N_3476);
and U4346 (N_4346,N_3648,N_3649);
nand U4347 (N_4347,N_3838,N_3529);
nand U4348 (N_4348,N_3621,N_3216);
and U4349 (N_4349,N_3204,N_3277);
and U4350 (N_4350,N_3232,N_3698);
and U4351 (N_4351,N_3259,N_3330);
nand U4352 (N_4352,N_3222,N_3203);
nand U4353 (N_4353,N_3679,N_3708);
nor U4354 (N_4354,N_3456,N_3282);
or U4355 (N_4355,N_3409,N_3266);
nor U4356 (N_4356,N_3842,N_3464);
nor U4357 (N_4357,N_3325,N_3245);
or U4358 (N_4358,N_3437,N_3572);
or U4359 (N_4359,N_3426,N_3289);
or U4360 (N_4360,N_3380,N_3947);
nand U4361 (N_4361,N_3796,N_3968);
nor U4362 (N_4362,N_3485,N_3981);
nand U4363 (N_4363,N_3930,N_3500);
nor U4364 (N_4364,N_3255,N_3959);
nor U4365 (N_4365,N_3707,N_3425);
nand U4366 (N_4366,N_3400,N_3356);
or U4367 (N_4367,N_3630,N_3914);
nor U4368 (N_4368,N_3729,N_3675);
nand U4369 (N_4369,N_3816,N_3202);
nor U4370 (N_4370,N_3973,N_3275);
and U4371 (N_4371,N_3200,N_3808);
and U4372 (N_4372,N_3469,N_3515);
nand U4373 (N_4373,N_3268,N_3549);
nand U4374 (N_4374,N_3880,N_3455);
or U4375 (N_4375,N_3446,N_3355);
or U4376 (N_4376,N_3962,N_3527);
and U4377 (N_4377,N_3769,N_3755);
nand U4378 (N_4378,N_3723,N_3886);
or U4379 (N_4379,N_3578,N_3598);
or U4380 (N_4380,N_3390,N_3241);
nand U4381 (N_4381,N_3912,N_3494);
and U4382 (N_4382,N_3352,N_3990);
and U4383 (N_4383,N_3770,N_3624);
nor U4384 (N_4384,N_3651,N_3357);
and U4385 (N_4385,N_3845,N_3567);
or U4386 (N_4386,N_3641,N_3923);
or U4387 (N_4387,N_3777,N_3219);
nor U4388 (N_4388,N_3925,N_3722);
or U4389 (N_4389,N_3684,N_3562);
nand U4390 (N_4390,N_3350,N_3211);
nand U4391 (N_4391,N_3806,N_3326);
or U4392 (N_4392,N_3632,N_3577);
nand U4393 (N_4393,N_3786,N_3720);
nor U4394 (N_4394,N_3859,N_3364);
nor U4395 (N_4395,N_3692,N_3823);
nand U4396 (N_4396,N_3841,N_3394);
and U4397 (N_4397,N_3774,N_3928);
and U4398 (N_4398,N_3799,N_3539);
nand U4399 (N_4399,N_3635,N_3459);
nand U4400 (N_4400,N_3205,N_3464);
and U4401 (N_4401,N_3969,N_3401);
and U4402 (N_4402,N_3227,N_3217);
or U4403 (N_4403,N_3389,N_3391);
and U4404 (N_4404,N_3541,N_3967);
and U4405 (N_4405,N_3855,N_3703);
nand U4406 (N_4406,N_3729,N_3660);
and U4407 (N_4407,N_3626,N_3686);
and U4408 (N_4408,N_3490,N_3645);
or U4409 (N_4409,N_3605,N_3798);
or U4410 (N_4410,N_3271,N_3819);
nor U4411 (N_4411,N_3711,N_3444);
nand U4412 (N_4412,N_3342,N_3605);
nor U4413 (N_4413,N_3459,N_3260);
nor U4414 (N_4414,N_3200,N_3933);
nor U4415 (N_4415,N_3404,N_3518);
nand U4416 (N_4416,N_3728,N_3456);
nor U4417 (N_4417,N_3699,N_3859);
and U4418 (N_4418,N_3596,N_3959);
nand U4419 (N_4419,N_3604,N_3620);
and U4420 (N_4420,N_3928,N_3818);
nand U4421 (N_4421,N_3521,N_3724);
and U4422 (N_4422,N_3565,N_3752);
or U4423 (N_4423,N_3282,N_3399);
nand U4424 (N_4424,N_3829,N_3619);
nand U4425 (N_4425,N_3587,N_3993);
nor U4426 (N_4426,N_3738,N_3626);
or U4427 (N_4427,N_3306,N_3948);
or U4428 (N_4428,N_3203,N_3988);
nor U4429 (N_4429,N_3475,N_3962);
nand U4430 (N_4430,N_3562,N_3289);
and U4431 (N_4431,N_3334,N_3235);
or U4432 (N_4432,N_3276,N_3783);
nand U4433 (N_4433,N_3388,N_3827);
and U4434 (N_4434,N_3371,N_3509);
nand U4435 (N_4435,N_3420,N_3767);
nand U4436 (N_4436,N_3220,N_3467);
nor U4437 (N_4437,N_3982,N_3284);
nand U4438 (N_4438,N_3901,N_3496);
and U4439 (N_4439,N_3716,N_3654);
or U4440 (N_4440,N_3954,N_3467);
and U4441 (N_4441,N_3487,N_3461);
or U4442 (N_4442,N_3508,N_3532);
nor U4443 (N_4443,N_3909,N_3658);
or U4444 (N_4444,N_3618,N_3294);
and U4445 (N_4445,N_3883,N_3778);
and U4446 (N_4446,N_3764,N_3981);
nor U4447 (N_4447,N_3494,N_3733);
nor U4448 (N_4448,N_3973,N_3563);
nand U4449 (N_4449,N_3616,N_3735);
and U4450 (N_4450,N_3344,N_3219);
and U4451 (N_4451,N_3938,N_3250);
nor U4452 (N_4452,N_3668,N_3844);
nand U4453 (N_4453,N_3643,N_3419);
nand U4454 (N_4454,N_3243,N_3827);
nor U4455 (N_4455,N_3709,N_3869);
and U4456 (N_4456,N_3755,N_3388);
xor U4457 (N_4457,N_3349,N_3226);
and U4458 (N_4458,N_3766,N_3953);
nor U4459 (N_4459,N_3247,N_3547);
and U4460 (N_4460,N_3707,N_3362);
and U4461 (N_4461,N_3389,N_3989);
or U4462 (N_4462,N_3250,N_3791);
or U4463 (N_4463,N_3881,N_3706);
nand U4464 (N_4464,N_3412,N_3644);
or U4465 (N_4465,N_3572,N_3950);
or U4466 (N_4466,N_3825,N_3268);
and U4467 (N_4467,N_3929,N_3636);
or U4468 (N_4468,N_3283,N_3744);
and U4469 (N_4469,N_3708,N_3845);
nor U4470 (N_4470,N_3284,N_3688);
and U4471 (N_4471,N_3315,N_3796);
nor U4472 (N_4472,N_3687,N_3404);
or U4473 (N_4473,N_3219,N_3932);
and U4474 (N_4474,N_3564,N_3743);
and U4475 (N_4475,N_3669,N_3307);
nor U4476 (N_4476,N_3978,N_3499);
and U4477 (N_4477,N_3421,N_3625);
or U4478 (N_4478,N_3828,N_3657);
or U4479 (N_4479,N_3692,N_3460);
or U4480 (N_4480,N_3482,N_3992);
nand U4481 (N_4481,N_3609,N_3499);
nor U4482 (N_4482,N_3982,N_3761);
nor U4483 (N_4483,N_3526,N_3912);
or U4484 (N_4484,N_3819,N_3324);
nor U4485 (N_4485,N_3727,N_3730);
or U4486 (N_4486,N_3997,N_3418);
or U4487 (N_4487,N_3762,N_3550);
nor U4488 (N_4488,N_3264,N_3613);
nor U4489 (N_4489,N_3665,N_3860);
nor U4490 (N_4490,N_3769,N_3287);
nor U4491 (N_4491,N_3408,N_3908);
nand U4492 (N_4492,N_3870,N_3935);
nor U4493 (N_4493,N_3604,N_3664);
nand U4494 (N_4494,N_3506,N_3743);
or U4495 (N_4495,N_3206,N_3450);
nand U4496 (N_4496,N_3875,N_3988);
nor U4497 (N_4497,N_3294,N_3963);
or U4498 (N_4498,N_3692,N_3671);
or U4499 (N_4499,N_3859,N_3988);
nor U4500 (N_4500,N_3832,N_3677);
and U4501 (N_4501,N_3708,N_3894);
nand U4502 (N_4502,N_3984,N_3648);
nor U4503 (N_4503,N_3433,N_3338);
or U4504 (N_4504,N_3689,N_3289);
and U4505 (N_4505,N_3448,N_3462);
nand U4506 (N_4506,N_3914,N_3255);
and U4507 (N_4507,N_3298,N_3465);
or U4508 (N_4508,N_3912,N_3424);
nor U4509 (N_4509,N_3862,N_3803);
or U4510 (N_4510,N_3258,N_3300);
or U4511 (N_4511,N_3614,N_3916);
nand U4512 (N_4512,N_3545,N_3332);
nand U4513 (N_4513,N_3650,N_3647);
or U4514 (N_4514,N_3385,N_3374);
nor U4515 (N_4515,N_3588,N_3874);
nor U4516 (N_4516,N_3458,N_3485);
nor U4517 (N_4517,N_3476,N_3252);
and U4518 (N_4518,N_3819,N_3838);
nand U4519 (N_4519,N_3937,N_3273);
nand U4520 (N_4520,N_3357,N_3731);
nand U4521 (N_4521,N_3921,N_3633);
and U4522 (N_4522,N_3286,N_3789);
or U4523 (N_4523,N_3550,N_3721);
or U4524 (N_4524,N_3491,N_3986);
or U4525 (N_4525,N_3617,N_3241);
or U4526 (N_4526,N_3607,N_3507);
nor U4527 (N_4527,N_3296,N_3744);
nor U4528 (N_4528,N_3672,N_3612);
and U4529 (N_4529,N_3721,N_3438);
and U4530 (N_4530,N_3759,N_3335);
or U4531 (N_4531,N_3525,N_3585);
nor U4532 (N_4532,N_3614,N_3839);
nor U4533 (N_4533,N_3269,N_3714);
nand U4534 (N_4534,N_3621,N_3523);
and U4535 (N_4535,N_3962,N_3599);
and U4536 (N_4536,N_3473,N_3954);
or U4537 (N_4537,N_3477,N_3785);
or U4538 (N_4538,N_3766,N_3704);
and U4539 (N_4539,N_3365,N_3349);
nor U4540 (N_4540,N_3778,N_3876);
or U4541 (N_4541,N_3957,N_3698);
nand U4542 (N_4542,N_3876,N_3939);
or U4543 (N_4543,N_3238,N_3243);
nor U4544 (N_4544,N_3925,N_3915);
or U4545 (N_4545,N_3726,N_3217);
nor U4546 (N_4546,N_3563,N_3515);
or U4547 (N_4547,N_3552,N_3290);
and U4548 (N_4548,N_3545,N_3527);
or U4549 (N_4549,N_3724,N_3511);
nor U4550 (N_4550,N_3627,N_3529);
nand U4551 (N_4551,N_3973,N_3733);
nand U4552 (N_4552,N_3533,N_3999);
nor U4553 (N_4553,N_3629,N_3721);
and U4554 (N_4554,N_3926,N_3269);
and U4555 (N_4555,N_3976,N_3540);
and U4556 (N_4556,N_3930,N_3577);
nor U4557 (N_4557,N_3458,N_3370);
or U4558 (N_4558,N_3524,N_3400);
nor U4559 (N_4559,N_3811,N_3667);
or U4560 (N_4560,N_3447,N_3499);
nand U4561 (N_4561,N_3214,N_3950);
nor U4562 (N_4562,N_3414,N_3717);
xnor U4563 (N_4563,N_3970,N_3955);
nor U4564 (N_4564,N_3765,N_3536);
nor U4565 (N_4565,N_3526,N_3236);
nor U4566 (N_4566,N_3253,N_3863);
nand U4567 (N_4567,N_3936,N_3594);
nand U4568 (N_4568,N_3251,N_3274);
nor U4569 (N_4569,N_3629,N_3547);
nand U4570 (N_4570,N_3505,N_3437);
nand U4571 (N_4571,N_3233,N_3984);
and U4572 (N_4572,N_3718,N_3693);
and U4573 (N_4573,N_3330,N_3982);
or U4574 (N_4574,N_3773,N_3313);
or U4575 (N_4575,N_3853,N_3605);
and U4576 (N_4576,N_3754,N_3938);
and U4577 (N_4577,N_3317,N_3224);
nor U4578 (N_4578,N_3472,N_3369);
and U4579 (N_4579,N_3249,N_3807);
and U4580 (N_4580,N_3243,N_3217);
xor U4581 (N_4581,N_3554,N_3407);
or U4582 (N_4582,N_3769,N_3922);
nor U4583 (N_4583,N_3706,N_3488);
or U4584 (N_4584,N_3293,N_3338);
xnor U4585 (N_4585,N_3608,N_3802);
nand U4586 (N_4586,N_3486,N_3352);
nor U4587 (N_4587,N_3761,N_3231);
and U4588 (N_4588,N_3834,N_3839);
nor U4589 (N_4589,N_3531,N_3341);
or U4590 (N_4590,N_3390,N_3306);
nor U4591 (N_4591,N_3631,N_3610);
nor U4592 (N_4592,N_3629,N_3407);
nand U4593 (N_4593,N_3701,N_3263);
or U4594 (N_4594,N_3245,N_3993);
or U4595 (N_4595,N_3969,N_3361);
or U4596 (N_4596,N_3206,N_3243);
nand U4597 (N_4597,N_3368,N_3991);
nand U4598 (N_4598,N_3661,N_3812);
nor U4599 (N_4599,N_3595,N_3600);
or U4600 (N_4600,N_3931,N_3693);
nand U4601 (N_4601,N_3219,N_3444);
nor U4602 (N_4602,N_3987,N_3782);
nor U4603 (N_4603,N_3291,N_3963);
or U4604 (N_4604,N_3485,N_3384);
and U4605 (N_4605,N_3486,N_3667);
and U4606 (N_4606,N_3414,N_3722);
nor U4607 (N_4607,N_3453,N_3204);
nand U4608 (N_4608,N_3757,N_3616);
or U4609 (N_4609,N_3248,N_3673);
or U4610 (N_4610,N_3699,N_3931);
or U4611 (N_4611,N_3701,N_3809);
and U4612 (N_4612,N_3490,N_3484);
and U4613 (N_4613,N_3545,N_3914);
or U4614 (N_4614,N_3867,N_3502);
nor U4615 (N_4615,N_3961,N_3508);
nand U4616 (N_4616,N_3515,N_3283);
and U4617 (N_4617,N_3839,N_3997);
nand U4618 (N_4618,N_3806,N_3840);
nand U4619 (N_4619,N_3795,N_3807);
or U4620 (N_4620,N_3407,N_3775);
or U4621 (N_4621,N_3985,N_3779);
nor U4622 (N_4622,N_3316,N_3418);
nor U4623 (N_4623,N_3873,N_3804);
and U4624 (N_4624,N_3421,N_3587);
and U4625 (N_4625,N_3325,N_3311);
nand U4626 (N_4626,N_3764,N_3457);
nor U4627 (N_4627,N_3423,N_3366);
nor U4628 (N_4628,N_3991,N_3589);
nand U4629 (N_4629,N_3990,N_3374);
nand U4630 (N_4630,N_3310,N_3972);
or U4631 (N_4631,N_3347,N_3565);
nand U4632 (N_4632,N_3375,N_3242);
or U4633 (N_4633,N_3482,N_3578);
nor U4634 (N_4634,N_3530,N_3255);
nor U4635 (N_4635,N_3827,N_3769);
nand U4636 (N_4636,N_3285,N_3521);
or U4637 (N_4637,N_3725,N_3662);
nor U4638 (N_4638,N_3660,N_3352);
nand U4639 (N_4639,N_3993,N_3779);
nor U4640 (N_4640,N_3433,N_3986);
and U4641 (N_4641,N_3736,N_3773);
nor U4642 (N_4642,N_3718,N_3363);
nand U4643 (N_4643,N_3575,N_3746);
nor U4644 (N_4644,N_3371,N_3745);
or U4645 (N_4645,N_3806,N_3324);
and U4646 (N_4646,N_3577,N_3776);
nand U4647 (N_4647,N_3350,N_3526);
and U4648 (N_4648,N_3383,N_3281);
or U4649 (N_4649,N_3275,N_3450);
and U4650 (N_4650,N_3903,N_3898);
and U4651 (N_4651,N_3338,N_3699);
nor U4652 (N_4652,N_3753,N_3730);
and U4653 (N_4653,N_3487,N_3565);
nor U4654 (N_4654,N_3530,N_3970);
and U4655 (N_4655,N_3328,N_3462);
nand U4656 (N_4656,N_3292,N_3337);
and U4657 (N_4657,N_3307,N_3892);
and U4658 (N_4658,N_3413,N_3486);
nor U4659 (N_4659,N_3921,N_3435);
and U4660 (N_4660,N_3601,N_3656);
and U4661 (N_4661,N_3465,N_3529);
and U4662 (N_4662,N_3216,N_3304);
nor U4663 (N_4663,N_3993,N_3999);
nor U4664 (N_4664,N_3497,N_3513);
nand U4665 (N_4665,N_3631,N_3411);
or U4666 (N_4666,N_3938,N_3538);
nor U4667 (N_4667,N_3615,N_3662);
nor U4668 (N_4668,N_3746,N_3419);
or U4669 (N_4669,N_3555,N_3553);
nor U4670 (N_4670,N_3937,N_3666);
or U4671 (N_4671,N_3340,N_3970);
nand U4672 (N_4672,N_3235,N_3391);
nand U4673 (N_4673,N_3575,N_3555);
and U4674 (N_4674,N_3984,N_3551);
nor U4675 (N_4675,N_3907,N_3808);
nand U4676 (N_4676,N_3203,N_3372);
and U4677 (N_4677,N_3907,N_3690);
nand U4678 (N_4678,N_3421,N_3407);
and U4679 (N_4679,N_3562,N_3242);
nand U4680 (N_4680,N_3568,N_3559);
nand U4681 (N_4681,N_3900,N_3570);
or U4682 (N_4682,N_3206,N_3609);
or U4683 (N_4683,N_3680,N_3562);
nor U4684 (N_4684,N_3854,N_3316);
nor U4685 (N_4685,N_3803,N_3544);
and U4686 (N_4686,N_3742,N_3994);
nor U4687 (N_4687,N_3523,N_3306);
nor U4688 (N_4688,N_3677,N_3852);
or U4689 (N_4689,N_3919,N_3786);
or U4690 (N_4690,N_3780,N_3398);
and U4691 (N_4691,N_3201,N_3930);
and U4692 (N_4692,N_3986,N_3793);
and U4693 (N_4693,N_3989,N_3402);
or U4694 (N_4694,N_3583,N_3921);
nor U4695 (N_4695,N_3823,N_3603);
and U4696 (N_4696,N_3828,N_3890);
xnor U4697 (N_4697,N_3913,N_3651);
nand U4698 (N_4698,N_3923,N_3215);
and U4699 (N_4699,N_3729,N_3739);
nor U4700 (N_4700,N_3338,N_3380);
nor U4701 (N_4701,N_3882,N_3808);
or U4702 (N_4702,N_3583,N_3554);
nor U4703 (N_4703,N_3366,N_3322);
nor U4704 (N_4704,N_3946,N_3536);
and U4705 (N_4705,N_3387,N_3368);
and U4706 (N_4706,N_3762,N_3326);
or U4707 (N_4707,N_3894,N_3511);
nand U4708 (N_4708,N_3809,N_3784);
nand U4709 (N_4709,N_3329,N_3489);
nand U4710 (N_4710,N_3811,N_3965);
and U4711 (N_4711,N_3694,N_3594);
nor U4712 (N_4712,N_3707,N_3429);
and U4713 (N_4713,N_3515,N_3935);
or U4714 (N_4714,N_3934,N_3769);
and U4715 (N_4715,N_3346,N_3271);
nor U4716 (N_4716,N_3499,N_3319);
and U4717 (N_4717,N_3959,N_3806);
nand U4718 (N_4718,N_3694,N_3218);
xnor U4719 (N_4719,N_3600,N_3690);
or U4720 (N_4720,N_3331,N_3886);
or U4721 (N_4721,N_3618,N_3470);
and U4722 (N_4722,N_3808,N_3979);
nand U4723 (N_4723,N_3402,N_3915);
or U4724 (N_4724,N_3826,N_3264);
or U4725 (N_4725,N_3749,N_3762);
nor U4726 (N_4726,N_3221,N_3773);
nor U4727 (N_4727,N_3206,N_3397);
and U4728 (N_4728,N_3748,N_3284);
nor U4729 (N_4729,N_3527,N_3832);
nand U4730 (N_4730,N_3736,N_3456);
or U4731 (N_4731,N_3243,N_3883);
and U4732 (N_4732,N_3325,N_3444);
nand U4733 (N_4733,N_3549,N_3248);
or U4734 (N_4734,N_3278,N_3555);
and U4735 (N_4735,N_3268,N_3217);
and U4736 (N_4736,N_3716,N_3405);
nor U4737 (N_4737,N_3310,N_3349);
or U4738 (N_4738,N_3622,N_3439);
nor U4739 (N_4739,N_3635,N_3204);
nand U4740 (N_4740,N_3333,N_3546);
nor U4741 (N_4741,N_3985,N_3468);
or U4742 (N_4742,N_3773,N_3650);
and U4743 (N_4743,N_3785,N_3532);
nor U4744 (N_4744,N_3611,N_3850);
nand U4745 (N_4745,N_3598,N_3839);
nand U4746 (N_4746,N_3902,N_3209);
or U4747 (N_4747,N_3842,N_3238);
and U4748 (N_4748,N_3606,N_3667);
nor U4749 (N_4749,N_3235,N_3823);
and U4750 (N_4750,N_3959,N_3243);
nor U4751 (N_4751,N_3881,N_3994);
or U4752 (N_4752,N_3867,N_3233);
nand U4753 (N_4753,N_3961,N_3745);
and U4754 (N_4754,N_3365,N_3647);
or U4755 (N_4755,N_3883,N_3783);
and U4756 (N_4756,N_3295,N_3876);
nand U4757 (N_4757,N_3359,N_3397);
nand U4758 (N_4758,N_3551,N_3636);
or U4759 (N_4759,N_3876,N_3410);
nand U4760 (N_4760,N_3621,N_3288);
or U4761 (N_4761,N_3258,N_3595);
nand U4762 (N_4762,N_3776,N_3490);
nand U4763 (N_4763,N_3239,N_3773);
or U4764 (N_4764,N_3746,N_3930);
and U4765 (N_4765,N_3964,N_3982);
or U4766 (N_4766,N_3848,N_3454);
nand U4767 (N_4767,N_3549,N_3650);
nor U4768 (N_4768,N_3864,N_3902);
and U4769 (N_4769,N_3847,N_3536);
nor U4770 (N_4770,N_3256,N_3741);
or U4771 (N_4771,N_3993,N_3677);
and U4772 (N_4772,N_3292,N_3247);
and U4773 (N_4773,N_3721,N_3347);
nor U4774 (N_4774,N_3979,N_3950);
nand U4775 (N_4775,N_3903,N_3609);
or U4776 (N_4776,N_3753,N_3956);
and U4777 (N_4777,N_3732,N_3421);
and U4778 (N_4778,N_3403,N_3335);
or U4779 (N_4779,N_3208,N_3224);
and U4780 (N_4780,N_3246,N_3422);
or U4781 (N_4781,N_3505,N_3834);
nand U4782 (N_4782,N_3435,N_3897);
nor U4783 (N_4783,N_3961,N_3360);
and U4784 (N_4784,N_3252,N_3770);
nand U4785 (N_4785,N_3644,N_3858);
or U4786 (N_4786,N_3215,N_3243);
or U4787 (N_4787,N_3990,N_3383);
nor U4788 (N_4788,N_3329,N_3247);
and U4789 (N_4789,N_3524,N_3240);
and U4790 (N_4790,N_3615,N_3967);
nor U4791 (N_4791,N_3912,N_3255);
or U4792 (N_4792,N_3946,N_3256);
or U4793 (N_4793,N_3985,N_3950);
nor U4794 (N_4794,N_3401,N_3514);
nand U4795 (N_4795,N_3586,N_3265);
nand U4796 (N_4796,N_3795,N_3838);
or U4797 (N_4797,N_3318,N_3852);
and U4798 (N_4798,N_3549,N_3700);
and U4799 (N_4799,N_3868,N_3830);
nor U4800 (N_4800,N_4770,N_4659);
or U4801 (N_4801,N_4641,N_4116);
and U4802 (N_4802,N_4099,N_4692);
or U4803 (N_4803,N_4695,N_4069);
nand U4804 (N_4804,N_4506,N_4230);
or U4805 (N_4805,N_4460,N_4163);
and U4806 (N_4806,N_4318,N_4756);
nor U4807 (N_4807,N_4119,N_4246);
or U4808 (N_4808,N_4202,N_4053);
nand U4809 (N_4809,N_4214,N_4113);
or U4810 (N_4810,N_4580,N_4187);
nor U4811 (N_4811,N_4540,N_4665);
nor U4812 (N_4812,N_4670,N_4628);
nand U4813 (N_4813,N_4104,N_4279);
or U4814 (N_4814,N_4209,N_4363);
nand U4815 (N_4815,N_4072,N_4698);
or U4816 (N_4816,N_4043,N_4168);
or U4817 (N_4817,N_4229,N_4590);
nand U4818 (N_4818,N_4410,N_4624);
nor U4819 (N_4819,N_4489,N_4056);
or U4820 (N_4820,N_4132,N_4255);
and U4821 (N_4821,N_4338,N_4123);
nand U4822 (N_4822,N_4402,N_4058);
nand U4823 (N_4823,N_4419,N_4503);
nand U4824 (N_4824,N_4257,N_4742);
and U4825 (N_4825,N_4423,N_4059);
or U4826 (N_4826,N_4693,N_4632);
or U4827 (N_4827,N_4436,N_4252);
nand U4828 (N_4828,N_4074,N_4592);
nor U4829 (N_4829,N_4373,N_4730);
or U4830 (N_4830,N_4519,N_4125);
nor U4831 (N_4831,N_4623,N_4518);
and U4832 (N_4832,N_4155,N_4388);
nor U4833 (N_4833,N_4383,N_4536);
nand U4834 (N_4834,N_4677,N_4650);
or U4835 (N_4835,N_4028,N_4378);
nor U4836 (N_4836,N_4182,N_4067);
nor U4837 (N_4837,N_4443,N_4703);
and U4838 (N_4838,N_4535,N_4548);
or U4839 (N_4839,N_4395,N_4728);
and U4840 (N_4840,N_4306,N_4139);
or U4841 (N_4841,N_4578,N_4581);
nand U4842 (N_4842,N_4292,N_4424);
nor U4843 (N_4843,N_4169,N_4459);
and U4844 (N_4844,N_4017,N_4153);
nor U4845 (N_4845,N_4406,N_4227);
or U4846 (N_4846,N_4405,N_4490);
or U4847 (N_4847,N_4060,N_4534);
and U4848 (N_4848,N_4587,N_4267);
and U4849 (N_4849,N_4064,N_4207);
nand U4850 (N_4850,N_4295,N_4159);
or U4851 (N_4851,N_4513,N_4583);
nand U4852 (N_4852,N_4030,N_4105);
or U4853 (N_4853,N_4316,N_4717);
nor U4854 (N_4854,N_4615,N_4366);
and U4855 (N_4855,N_4706,N_4746);
nor U4856 (N_4856,N_4263,N_4184);
or U4857 (N_4857,N_4517,N_4510);
and U4858 (N_4858,N_4667,N_4653);
nor U4859 (N_4859,N_4085,N_4057);
nand U4860 (N_4860,N_4342,N_4287);
and U4861 (N_4861,N_4718,N_4694);
and U4862 (N_4862,N_4784,N_4013);
or U4863 (N_4863,N_4157,N_4183);
nor U4864 (N_4864,N_4725,N_4062);
nor U4865 (N_4865,N_4430,N_4304);
nor U4866 (N_4866,N_4759,N_4411);
nand U4867 (N_4867,N_4264,N_4451);
nor U4868 (N_4868,N_4780,N_4764);
and U4869 (N_4869,N_4269,N_4744);
or U4870 (N_4870,N_4646,N_4337);
nor U4871 (N_4871,N_4731,N_4418);
nor U4872 (N_4872,N_4468,N_4170);
or U4873 (N_4873,N_4450,N_4538);
and U4874 (N_4874,N_4754,N_4775);
nand U4875 (N_4875,N_4788,N_4003);
and U4876 (N_4876,N_4470,N_4205);
and U4877 (N_4877,N_4322,N_4432);
or U4878 (N_4878,N_4595,N_4111);
or U4879 (N_4879,N_4721,N_4068);
or U4880 (N_4880,N_4765,N_4236);
or U4881 (N_4881,N_4140,N_4012);
or U4882 (N_4882,N_4189,N_4714);
nand U4883 (N_4883,N_4179,N_4626);
or U4884 (N_4884,N_4124,N_4296);
nor U4885 (N_4885,N_4127,N_4479);
nor U4886 (N_4886,N_4211,N_4158);
and U4887 (N_4887,N_4114,N_4772);
and U4888 (N_4888,N_4096,N_4095);
nor U4889 (N_4889,N_4572,N_4630);
nand U4890 (N_4890,N_4621,N_4782);
and U4891 (N_4891,N_4607,N_4370);
and U4892 (N_4892,N_4781,N_4672);
and U4893 (N_4893,N_4385,N_4799);
nand U4894 (N_4894,N_4444,N_4729);
nand U4895 (N_4895,N_4549,N_4250);
nand U4896 (N_4896,N_4537,N_4259);
nor U4897 (N_4897,N_4226,N_4633);
and U4898 (N_4898,N_4018,N_4006);
nand U4899 (N_4899,N_4225,N_4708);
and U4900 (N_4900,N_4285,N_4458);
nand U4901 (N_4901,N_4228,N_4223);
nand U4902 (N_4902,N_4610,N_4608);
nor U4903 (N_4903,N_4545,N_4086);
nor U4904 (N_4904,N_4574,N_4025);
and U4905 (N_4905,N_4502,N_4663);
or U4906 (N_4906,N_4673,N_4685);
or U4907 (N_4907,N_4351,N_4231);
or U4908 (N_4908,N_4551,N_4190);
nor U4909 (N_4909,N_4492,N_4319);
or U4910 (N_4910,N_4379,N_4128);
nor U4911 (N_4911,N_4658,N_4483);
nor U4912 (N_4912,N_4606,N_4559);
nor U4913 (N_4913,N_4245,N_4041);
nor U4914 (N_4914,N_4117,N_4154);
nor U4915 (N_4915,N_4529,N_4611);
nor U4916 (N_4916,N_4773,N_4253);
nor U4917 (N_4917,N_4200,N_4616);
nand U4918 (N_4918,N_4499,N_4464);
or U4919 (N_4919,N_4431,N_4216);
nor U4920 (N_4920,N_4629,N_4674);
or U4921 (N_4921,N_4270,N_4651);
or U4922 (N_4922,N_4346,N_4527);
nor U4923 (N_4923,N_4533,N_4272);
nand U4924 (N_4924,N_4361,N_4177);
or U4925 (N_4925,N_4682,N_4711);
or U4926 (N_4926,N_4634,N_4577);
or U4927 (N_4927,N_4348,N_4009);
and U4928 (N_4928,N_4080,N_4311);
nand U4929 (N_4929,N_4582,N_4409);
and U4930 (N_4930,N_4643,N_4303);
nor U4931 (N_4931,N_4120,N_4709);
nand U4932 (N_4932,N_4389,N_4493);
and U4933 (N_4933,N_4349,N_4232);
nand U4934 (N_4934,N_4106,N_4798);
and U4935 (N_4935,N_4397,N_4484);
nor U4936 (N_4936,N_4305,N_4426);
nor U4937 (N_4937,N_4477,N_4102);
and U4938 (N_4938,N_4568,N_4707);
or U4939 (N_4939,N_4103,N_4690);
and U4940 (N_4940,N_4049,N_4218);
and U4941 (N_4941,N_4181,N_4520);
nor U4942 (N_4942,N_4261,N_4330);
nand U4943 (N_4943,N_4761,N_4283);
and U4944 (N_4944,N_4427,N_4525);
or U4945 (N_4945,N_4314,N_4199);
nand U4946 (N_4946,N_4666,N_4593);
and U4947 (N_4947,N_4065,N_4332);
xor U4948 (N_4948,N_4648,N_4413);
nand U4949 (N_4949,N_4191,N_4194);
and U4950 (N_4950,N_4357,N_4515);
or U4951 (N_4951,N_4093,N_4462);
and U4952 (N_4952,N_4089,N_4282);
and U4953 (N_4953,N_4408,N_4763);
nand U4954 (N_4954,N_4212,N_4591);
nand U4955 (N_4955,N_4523,N_4473);
and U4956 (N_4956,N_4662,N_4531);
or U4957 (N_4957,N_4455,N_4073);
or U4958 (N_4958,N_4317,N_4147);
and U4959 (N_4959,N_4329,N_4552);
nand U4960 (N_4960,N_4078,N_4481);
or U4961 (N_4961,N_4735,N_4596);
and U4962 (N_4962,N_4055,N_4689);
nor U4963 (N_4963,N_4241,N_4291);
nor U4964 (N_4964,N_4237,N_4751);
nand U4965 (N_4965,N_4040,N_4452);
and U4966 (N_4966,N_4433,N_4343);
nand U4967 (N_4967,N_4206,N_4456);
nor U4968 (N_4968,N_4441,N_4010);
and U4969 (N_4969,N_4213,N_4027);
nor U4970 (N_4970,N_4647,N_4723);
and U4971 (N_4971,N_4779,N_4571);
and U4972 (N_4972,N_4563,N_4129);
and U4973 (N_4973,N_4740,N_4268);
nand U4974 (N_4974,N_4288,N_4133);
or U4975 (N_4975,N_4752,N_4193);
nor U4976 (N_4976,N_4716,N_4614);
and U4977 (N_4977,N_4710,N_4768);
and U4978 (N_4978,N_4079,N_4428);
nand U4979 (N_4979,N_4618,N_4495);
and U4980 (N_4980,N_4371,N_4249);
nand U4981 (N_4981,N_4469,N_4727);
nand U4982 (N_4982,N_4284,N_4032);
and U4983 (N_4983,N_4739,N_4134);
or U4984 (N_4984,N_4774,N_4434);
nand U4985 (N_4985,N_4586,N_4247);
nor U4986 (N_4986,N_4446,N_4457);
nand U4987 (N_4987,N_4425,N_4180);
and U4988 (N_4988,N_4248,N_4145);
and U4989 (N_4989,N_4704,N_4350);
and U4990 (N_4990,N_4115,N_4174);
and U4991 (N_4991,N_4325,N_4654);
and U4992 (N_4992,N_4299,N_4612);
nand U4993 (N_4993,N_4466,N_4414);
nor U4994 (N_4994,N_4576,N_4126);
nand U4995 (N_4995,N_4321,N_4748);
and U4996 (N_4996,N_4637,N_4656);
nor U4997 (N_4997,N_4442,N_4192);
or U4998 (N_4998,N_4491,N_4471);
or U4999 (N_4999,N_4084,N_4448);
or U5000 (N_5000,N_4273,N_4386);
nor U5001 (N_5001,N_4594,N_4556);
nand U5002 (N_5002,N_4570,N_4235);
or U5003 (N_5003,N_4108,N_4308);
nand U5004 (N_5004,N_4365,N_4565);
and U5005 (N_5005,N_4684,N_4394);
nor U5006 (N_5006,N_4737,N_4603);
nor U5007 (N_5007,N_4324,N_4627);
nand U5008 (N_5008,N_4101,N_4256);
nor U5009 (N_5009,N_4328,N_4546);
or U5010 (N_5010,N_4793,N_4429);
and U5011 (N_5011,N_4239,N_4175);
nor U5012 (N_5012,N_4691,N_4029);
nor U5013 (N_5013,N_4390,N_4008);
or U5014 (N_5014,N_4242,N_4403);
nand U5015 (N_5015,N_4355,N_4575);
and U5016 (N_5016,N_4541,N_4617);
and U5017 (N_5017,N_4340,N_4033);
or U5018 (N_5018,N_4286,N_4715);
nor U5019 (N_5019,N_4776,N_4507);
nand U5020 (N_5020,N_4185,N_4486);
nand U5021 (N_5021,N_4146,N_4688);
nand U5022 (N_5022,N_4360,N_4075);
nor U5023 (N_5023,N_4001,N_4050);
and U5024 (N_5024,N_4655,N_4795);
nand U5025 (N_5025,N_4494,N_4220);
and U5026 (N_5026,N_4094,N_4726);
or U5027 (N_5027,N_4121,N_4031);
and U5028 (N_5028,N_4664,N_4475);
and U5029 (N_5029,N_4312,N_4165);
nand U5030 (N_5030,N_4732,N_4234);
nand U5031 (N_5031,N_4152,N_4671);
nor U5032 (N_5032,N_4258,N_4609);
or U5033 (N_5033,N_4465,N_4112);
nor U5034 (N_5034,N_4301,N_4500);
and U5035 (N_5035,N_4136,N_4024);
and U5036 (N_5036,N_4445,N_4061);
nand U5037 (N_5037,N_4530,N_4021);
or U5038 (N_5038,N_4547,N_4543);
or U5039 (N_5039,N_4555,N_4757);
nand U5040 (N_5040,N_4561,N_4352);
nand U5041 (N_5041,N_4160,N_4110);
or U5042 (N_5042,N_4020,N_4642);
or U5043 (N_5043,N_4487,N_4047);
nand U5044 (N_5044,N_4790,N_4036);
nor U5045 (N_5045,N_4196,N_4198);
or U5046 (N_5046,N_4797,N_4144);
or U5047 (N_5047,N_4401,N_4300);
and U5048 (N_5048,N_4749,N_4156);
nor U5049 (N_5049,N_4638,N_4573);
nand U5050 (N_5050,N_4562,N_4313);
nor U5051 (N_5051,N_4417,N_4222);
nor U5052 (N_5052,N_4393,N_4090);
nand U5053 (N_5053,N_4254,N_4794);
or U5054 (N_5054,N_4310,N_4092);
or U5055 (N_5055,N_4142,N_4336);
xor U5056 (N_5056,N_4496,N_4720);
nand U5057 (N_5057,N_4400,N_4070);
or U5058 (N_5058,N_4597,N_4497);
nand U5059 (N_5059,N_4512,N_4161);
and U5060 (N_5060,N_4364,N_4369);
nor U5061 (N_5061,N_4046,N_4038);
or U5062 (N_5062,N_4713,N_4767);
or U5063 (N_5063,N_4712,N_4696);
nor U5064 (N_5064,N_4353,N_4544);
nor U5065 (N_5065,N_4356,N_4368);
or U5066 (N_5066,N_4521,N_4109);
and U5067 (N_5067,N_4374,N_4063);
or U5068 (N_5068,N_4553,N_4498);
nand U5069 (N_5069,N_4381,N_4240);
or U5070 (N_5070,N_4440,N_4091);
and U5071 (N_5071,N_4195,N_4143);
nand U5072 (N_5072,N_4474,N_4557);
and U5073 (N_5073,N_4290,N_4702);
nor U5074 (N_5074,N_4275,N_4081);
nand U5075 (N_5075,N_4392,N_4331);
and U5076 (N_5076,N_4044,N_4644);
nand U5077 (N_5077,N_4326,N_4422);
nor U5078 (N_5078,N_4605,N_4293);
and U5079 (N_5079,N_4449,N_4148);
and U5080 (N_5080,N_4039,N_4420);
or U5081 (N_5081,N_4380,N_4783);
or U5082 (N_5082,N_4107,N_4197);
nand U5083 (N_5083,N_4755,N_4243);
or U5084 (N_5084,N_4435,N_4511);
xnor U5085 (N_5085,N_4640,N_4204);
nor U5086 (N_5086,N_4088,N_4260);
nor U5087 (N_5087,N_4224,N_4649);
or U5088 (N_5088,N_4657,N_4604);
nand U5089 (N_5089,N_4130,N_4620);
nor U5090 (N_5090,N_4785,N_4554);
or U5091 (N_5091,N_4387,N_4645);
nand U5092 (N_5092,N_4508,N_4384);
or U5093 (N_5093,N_4558,N_4528);
and U5094 (N_5094,N_4743,N_4164);
xnor U5095 (N_5095,N_4289,N_4741);
nor U5096 (N_5096,N_4705,N_4678);
nand U5097 (N_5097,N_4722,N_4376);
nand U5098 (N_5098,N_4482,N_4699);
nor U5099 (N_5099,N_4051,N_4005);
nand U5100 (N_5100,N_4524,N_4208);
and U5101 (N_5101,N_4004,N_4244);
or U5102 (N_5102,N_4738,N_4485);
nand U5103 (N_5103,N_4201,N_4472);
or U5104 (N_5104,N_4323,N_4334);
nand U5105 (N_5105,N_4463,N_4042);
nor U5106 (N_5106,N_4514,N_4437);
nand U5107 (N_5107,N_4302,N_4362);
nand U5108 (N_5108,N_4598,N_4377);
nor U5109 (N_5109,N_4736,N_4421);
or U5110 (N_5110,N_4309,N_4686);
nand U5111 (N_5111,N_4467,N_4600);
nand U5112 (N_5112,N_4335,N_4167);
nand U5113 (N_5113,N_4675,N_4266);
nand U5114 (N_5114,N_4100,N_4122);
nand U5115 (N_5115,N_4271,N_4588);
and U5116 (N_5116,N_4026,N_4747);
and U5117 (N_5117,N_4636,N_4054);
nand U5118 (N_5118,N_4344,N_4215);
and U5119 (N_5119,N_4137,N_4461);
nor U5120 (N_5120,N_4320,N_4048);
and U5121 (N_5121,N_4791,N_4777);
or U5122 (N_5122,N_4173,N_4097);
nor U5123 (N_5123,N_4135,N_4679);
or U5124 (N_5124,N_4345,N_4382);
nor U5125 (N_5125,N_4622,N_4087);
and U5126 (N_5126,N_4083,N_4786);
and U5127 (N_5127,N_4203,N_4045);
and U5128 (N_5128,N_4480,N_4034);
nor U5129 (N_5129,N_4687,N_4542);
or U5130 (N_5130,N_4066,N_4023);
and U5131 (N_5131,N_4082,N_4758);
nor U5132 (N_5132,N_4141,N_4416);
and U5133 (N_5133,N_4149,N_4327);
and U5134 (N_5134,N_4014,N_4560);
nor U5135 (N_5135,N_4526,N_4447);
or U5136 (N_5136,N_4007,N_4399);
nor U5137 (N_5137,N_4019,N_4238);
and U5138 (N_5138,N_4000,N_4697);
nor U5139 (N_5139,N_4276,N_4118);
and U5140 (N_5140,N_4298,N_4412);
and U5141 (N_5141,N_4398,N_4166);
or U5142 (N_5142,N_4262,N_4661);
nor U5143 (N_5143,N_4076,N_4439);
or U5144 (N_5144,N_4488,N_4652);
and U5145 (N_5145,N_4639,N_4476);
nor U5146 (N_5146,N_4233,N_4186);
nor U5147 (N_5147,N_4683,N_4769);
nor U5148 (N_5148,N_4307,N_4796);
xnor U5149 (N_5149,N_4567,N_4219);
nor U5150 (N_5150,N_4766,N_4002);
and U5151 (N_5151,N_4011,N_4660);
nor U5152 (N_5152,N_4354,N_4367);
nor U5153 (N_5153,N_4505,N_4171);
and U5154 (N_5154,N_4052,N_4071);
nand U5155 (N_5155,N_4619,N_4037);
and U5156 (N_5156,N_4733,N_4265);
and U5157 (N_5157,N_4522,N_4719);
or U5158 (N_5158,N_4391,N_4359);
nor U5159 (N_5159,N_4599,N_4294);
nand U5160 (N_5160,N_4584,N_4022);
or U5161 (N_5161,N_4625,N_4151);
nand U5162 (N_5162,N_4589,N_4753);
and U5163 (N_5163,N_4404,N_4792);
nand U5164 (N_5164,N_4635,N_4566);
or U5165 (N_5165,N_4701,N_4789);
nor U5166 (N_5166,N_4750,N_4501);
and U5167 (N_5167,N_4762,N_4339);
and U5168 (N_5168,N_4358,N_4669);
and U5169 (N_5169,N_4724,N_4016);
nor U5170 (N_5170,N_4564,N_4407);
and U5171 (N_5171,N_4172,N_4138);
or U5172 (N_5172,N_4631,N_4680);
or U5173 (N_5173,N_4585,N_4532);
and U5174 (N_5174,N_4415,N_4098);
or U5175 (N_5175,N_4150,N_4787);
nand U5176 (N_5176,N_4015,N_4771);
and U5177 (N_5177,N_4613,N_4509);
or U5178 (N_5178,N_4077,N_4278);
and U5179 (N_5179,N_4539,N_4178);
nand U5180 (N_5180,N_4333,N_4176);
or U5181 (N_5181,N_4396,N_4516);
and U5182 (N_5182,N_4188,N_4372);
nand U5183 (N_5183,N_4760,N_4281);
nand U5184 (N_5184,N_4478,N_4778);
and U5185 (N_5185,N_4341,N_4277);
or U5186 (N_5186,N_4131,N_4602);
and U5187 (N_5187,N_4700,N_4297);
or U5188 (N_5188,N_4601,N_4221);
nand U5189 (N_5189,N_4274,N_4668);
nor U5190 (N_5190,N_4438,N_4504);
nor U5191 (N_5191,N_4315,N_4210);
nor U5192 (N_5192,N_4681,N_4676);
or U5193 (N_5193,N_4280,N_4217);
nand U5194 (N_5194,N_4569,N_4454);
nand U5195 (N_5195,N_4745,N_4453);
nand U5196 (N_5196,N_4162,N_4251);
nand U5197 (N_5197,N_4035,N_4734);
or U5198 (N_5198,N_4347,N_4579);
nand U5199 (N_5199,N_4550,N_4375);
or U5200 (N_5200,N_4652,N_4169);
or U5201 (N_5201,N_4615,N_4072);
nor U5202 (N_5202,N_4315,N_4374);
and U5203 (N_5203,N_4550,N_4576);
and U5204 (N_5204,N_4345,N_4225);
nor U5205 (N_5205,N_4251,N_4363);
and U5206 (N_5206,N_4632,N_4130);
nand U5207 (N_5207,N_4298,N_4006);
or U5208 (N_5208,N_4035,N_4728);
nor U5209 (N_5209,N_4289,N_4120);
and U5210 (N_5210,N_4592,N_4336);
nor U5211 (N_5211,N_4672,N_4542);
or U5212 (N_5212,N_4316,N_4262);
or U5213 (N_5213,N_4300,N_4192);
nand U5214 (N_5214,N_4424,N_4487);
nand U5215 (N_5215,N_4179,N_4513);
nor U5216 (N_5216,N_4043,N_4428);
or U5217 (N_5217,N_4198,N_4798);
nand U5218 (N_5218,N_4289,N_4660);
and U5219 (N_5219,N_4087,N_4147);
nor U5220 (N_5220,N_4177,N_4157);
and U5221 (N_5221,N_4504,N_4561);
and U5222 (N_5222,N_4520,N_4482);
and U5223 (N_5223,N_4335,N_4268);
or U5224 (N_5224,N_4405,N_4727);
nor U5225 (N_5225,N_4321,N_4054);
or U5226 (N_5226,N_4151,N_4165);
nor U5227 (N_5227,N_4596,N_4388);
nor U5228 (N_5228,N_4518,N_4116);
nor U5229 (N_5229,N_4599,N_4594);
and U5230 (N_5230,N_4160,N_4291);
nand U5231 (N_5231,N_4510,N_4371);
or U5232 (N_5232,N_4635,N_4294);
nand U5233 (N_5233,N_4227,N_4786);
nor U5234 (N_5234,N_4028,N_4433);
nand U5235 (N_5235,N_4000,N_4230);
or U5236 (N_5236,N_4571,N_4780);
nor U5237 (N_5237,N_4486,N_4219);
and U5238 (N_5238,N_4214,N_4409);
and U5239 (N_5239,N_4699,N_4251);
or U5240 (N_5240,N_4459,N_4790);
nor U5241 (N_5241,N_4611,N_4441);
and U5242 (N_5242,N_4292,N_4251);
or U5243 (N_5243,N_4678,N_4332);
nand U5244 (N_5244,N_4475,N_4746);
nand U5245 (N_5245,N_4386,N_4425);
nand U5246 (N_5246,N_4480,N_4180);
nand U5247 (N_5247,N_4219,N_4516);
or U5248 (N_5248,N_4067,N_4068);
nand U5249 (N_5249,N_4149,N_4509);
nor U5250 (N_5250,N_4462,N_4709);
nand U5251 (N_5251,N_4181,N_4089);
nor U5252 (N_5252,N_4722,N_4363);
or U5253 (N_5253,N_4260,N_4002);
or U5254 (N_5254,N_4240,N_4176);
nand U5255 (N_5255,N_4426,N_4418);
and U5256 (N_5256,N_4766,N_4613);
or U5257 (N_5257,N_4220,N_4621);
nor U5258 (N_5258,N_4269,N_4488);
nand U5259 (N_5259,N_4747,N_4634);
or U5260 (N_5260,N_4105,N_4493);
nand U5261 (N_5261,N_4284,N_4392);
or U5262 (N_5262,N_4138,N_4625);
nand U5263 (N_5263,N_4488,N_4614);
or U5264 (N_5264,N_4439,N_4445);
and U5265 (N_5265,N_4330,N_4214);
nor U5266 (N_5266,N_4391,N_4234);
nand U5267 (N_5267,N_4728,N_4005);
or U5268 (N_5268,N_4321,N_4204);
nand U5269 (N_5269,N_4264,N_4307);
nor U5270 (N_5270,N_4274,N_4359);
and U5271 (N_5271,N_4474,N_4552);
or U5272 (N_5272,N_4171,N_4720);
or U5273 (N_5273,N_4376,N_4686);
nor U5274 (N_5274,N_4698,N_4204);
nand U5275 (N_5275,N_4661,N_4211);
or U5276 (N_5276,N_4664,N_4016);
and U5277 (N_5277,N_4764,N_4125);
nor U5278 (N_5278,N_4384,N_4246);
nor U5279 (N_5279,N_4669,N_4489);
nor U5280 (N_5280,N_4635,N_4414);
or U5281 (N_5281,N_4774,N_4161);
nor U5282 (N_5282,N_4244,N_4448);
or U5283 (N_5283,N_4070,N_4124);
nor U5284 (N_5284,N_4563,N_4708);
or U5285 (N_5285,N_4610,N_4576);
nor U5286 (N_5286,N_4599,N_4120);
nor U5287 (N_5287,N_4673,N_4410);
nor U5288 (N_5288,N_4361,N_4343);
or U5289 (N_5289,N_4020,N_4695);
nor U5290 (N_5290,N_4052,N_4100);
nand U5291 (N_5291,N_4514,N_4041);
or U5292 (N_5292,N_4037,N_4408);
or U5293 (N_5293,N_4116,N_4513);
or U5294 (N_5294,N_4668,N_4533);
nand U5295 (N_5295,N_4132,N_4314);
nand U5296 (N_5296,N_4787,N_4296);
nand U5297 (N_5297,N_4124,N_4502);
or U5298 (N_5298,N_4158,N_4541);
and U5299 (N_5299,N_4609,N_4618);
and U5300 (N_5300,N_4728,N_4781);
and U5301 (N_5301,N_4350,N_4130);
nor U5302 (N_5302,N_4176,N_4768);
nand U5303 (N_5303,N_4455,N_4032);
nor U5304 (N_5304,N_4612,N_4249);
and U5305 (N_5305,N_4488,N_4580);
nand U5306 (N_5306,N_4612,N_4331);
or U5307 (N_5307,N_4048,N_4377);
and U5308 (N_5308,N_4016,N_4060);
nor U5309 (N_5309,N_4764,N_4458);
and U5310 (N_5310,N_4715,N_4071);
and U5311 (N_5311,N_4736,N_4246);
or U5312 (N_5312,N_4370,N_4755);
or U5313 (N_5313,N_4498,N_4705);
nand U5314 (N_5314,N_4798,N_4078);
nor U5315 (N_5315,N_4307,N_4122);
nand U5316 (N_5316,N_4371,N_4050);
nand U5317 (N_5317,N_4344,N_4725);
nor U5318 (N_5318,N_4440,N_4443);
nor U5319 (N_5319,N_4290,N_4399);
and U5320 (N_5320,N_4582,N_4284);
nand U5321 (N_5321,N_4181,N_4541);
or U5322 (N_5322,N_4589,N_4411);
and U5323 (N_5323,N_4699,N_4372);
nand U5324 (N_5324,N_4674,N_4695);
and U5325 (N_5325,N_4198,N_4714);
nor U5326 (N_5326,N_4350,N_4077);
or U5327 (N_5327,N_4398,N_4107);
or U5328 (N_5328,N_4029,N_4033);
nor U5329 (N_5329,N_4201,N_4454);
nand U5330 (N_5330,N_4575,N_4398);
nor U5331 (N_5331,N_4094,N_4518);
nor U5332 (N_5332,N_4554,N_4056);
and U5333 (N_5333,N_4277,N_4382);
nor U5334 (N_5334,N_4692,N_4276);
nor U5335 (N_5335,N_4301,N_4078);
nor U5336 (N_5336,N_4297,N_4465);
and U5337 (N_5337,N_4722,N_4657);
nor U5338 (N_5338,N_4641,N_4612);
xnor U5339 (N_5339,N_4681,N_4528);
xnor U5340 (N_5340,N_4075,N_4381);
nor U5341 (N_5341,N_4227,N_4458);
and U5342 (N_5342,N_4164,N_4326);
and U5343 (N_5343,N_4463,N_4556);
or U5344 (N_5344,N_4356,N_4564);
nand U5345 (N_5345,N_4088,N_4674);
nor U5346 (N_5346,N_4634,N_4669);
nor U5347 (N_5347,N_4512,N_4216);
and U5348 (N_5348,N_4418,N_4061);
nor U5349 (N_5349,N_4704,N_4434);
or U5350 (N_5350,N_4671,N_4578);
nor U5351 (N_5351,N_4606,N_4738);
nor U5352 (N_5352,N_4333,N_4227);
nand U5353 (N_5353,N_4711,N_4248);
and U5354 (N_5354,N_4305,N_4034);
or U5355 (N_5355,N_4152,N_4753);
nand U5356 (N_5356,N_4798,N_4455);
and U5357 (N_5357,N_4006,N_4437);
and U5358 (N_5358,N_4126,N_4686);
nand U5359 (N_5359,N_4573,N_4391);
or U5360 (N_5360,N_4129,N_4102);
or U5361 (N_5361,N_4501,N_4735);
nor U5362 (N_5362,N_4142,N_4507);
and U5363 (N_5363,N_4682,N_4223);
nand U5364 (N_5364,N_4649,N_4698);
nor U5365 (N_5365,N_4361,N_4359);
nor U5366 (N_5366,N_4516,N_4427);
and U5367 (N_5367,N_4370,N_4731);
and U5368 (N_5368,N_4543,N_4458);
nor U5369 (N_5369,N_4038,N_4681);
and U5370 (N_5370,N_4046,N_4285);
nand U5371 (N_5371,N_4478,N_4506);
or U5372 (N_5372,N_4652,N_4003);
or U5373 (N_5373,N_4575,N_4572);
and U5374 (N_5374,N_4009,N_4394);
or U5375 (N_5375,N_4003,N_4707);
or U5376 (N_5376,N_4557,N_4358);
or U5377 (N_5377,N_4200,N_4724);
and U5378 (N_5378,N_4674,N_4189);
nor U5379 (N_5379,N_4192,N_4089);
and U5380 (N_5380,N_4322,N_4198);
nor U5381 (N_5381,N_4741,N_4140);
nand U5382 (N_5382,N_4320,N_4164);
nand U5383 (N_5383,N_4602,N_4358);
or U5384 (N_5384,N_4404,N_4686);
nor U5385 (N_5385,N_4137,N_4614);
nand U5386 (N_5386,N_4374,N_4307);
or U5387 (N_5387,N_4305,N_4250);
nand U5388 (N_5388,N_4664,N_4617);
and U5389 (N_5389,N_4773,N_4524);
or U5390 (N_5390,N_4049,N_4263);
or U5391 (N_5391,N_4051,N_4101);
or U5392 (N_5392,N_4037,N_4217);
or U5393 (N_5393,N_4300,N_4396);
or U5394 (N_5394,N_4334,N_4066);
and U5395 (N_5395,N_4220,N_4107);
nand U5396 (N_5396,N_4069,N_4306);
nand U5397 (N_5397,N_4245,N_4583);
nor U5398 (N_5398,N_4688,N_4192);
and U5399 (N_5399,N_4198,N_4486);
nand U5400 (N_5400,N_4034,N_4540);
and U5401 (N_5401,N_4695,N_4447);
nand U5402 (N_5402,N_4719,N_4772);
nor U5403 (N_5403,N_4441,N_4630);
nor U5404 (N_5404,N_4572,N_4121);
nor U5405 (N_5405,N_4085,N_4180);
nand U5406 (N_5406,N_4680,N_4685);
nand U5407 (N_5407,N_4307,N_4306);
and U5408 (N_5408,N_4584,N_4173);
nand U5409 (N_5409,N_4066,N_4350);
nand U5410 (N_5410,N_4595,N_4564);
nand U5411 (N_5411,N_4035,N_4776);
or U5412 (N_5412,N_4110,N_4277);
or U5413 (N_5413,N_4555,N_4453);
and U5414 (N_5414,N_4006,N_4469);
and U5415 (N_5415,N_4633,N_4220);
or U5416 (N_5416,N_4708,N_4323);
and U5417 (N_5417,N_4294,N_4760);
and U5418 (N_5418,N_4041,N_4675);
xnor U5419 (N_5419,N_4199,N_4331);
nor U5420 (N_5420,N_4280,N_4641);
or U5421 (N_5421,N_4167,N_4434);
nand U5422 (N_5422,N_4488,N_4464);
nor U5423 (N_5423,N_4695,N_4281);
nand U5424 (N_5424,N_4182,N_4712);
nor U5425 (N_5425,N_4295,N_4527);
nor U5426 (N_5426,N_4544,N_4163);
and U5427 (N_5427,N_4388,N_4482);
or U5428 (N_5428,N_4167,N_4170);
and U5429 (N_5429,N_4226,N_4641);
or U5430 (N_5430,N_4380,N_4673);
or U5431 (N_5431,N_4710,N_4261);
or U5432 (N_5432,N_4067,N_4663);
nor U5433 (N_5433,N_4381,N_4057);
nand U5434 (N_5434,N_4115,N_4658);
nand U5435 (N_5435,N_4635,N_4633);
nor U5436 (N_5436,N_4280,N_4054);
nand U5437 (N_5437,N_4170,N_4152);
nand U5438 (N_5438,N_4032,N_4482);
and U5439 (N_5439,N_4409,N_4407);
nor U5440 (N_5440,N_4770,N_4625);
or U5441 (N_5441,N_4334,N_4294);
or U5442 (N_5442,N_4396,N_4460);
nor U5443 (N_5443,N_4078,N_4750);
nand U5444 (N_5444,N_4037,N_4088);
or U5445 (N_5445,N_4259,N_4760);
and U5446 (N_5446,N_4044,N_4026);
or U5447 (N_5447,N_4117,N_4383);
or U5448 (N_5448,N_4619,N_4149);
nand U5449 (N_5449,N_4330,N_4129);
xor U5450 (N_5450,N_4039,N_4061);
or U5451 (N_5451,N_4209,N_4548);
nor U5452 (N_5452,N_4683,N_4357);
nor U5453 (N_5453,N_4714,N_4234);
and U5454 (N_5454,N_4443,N_4735);
nor U5455 (N_5455,N_4457,N_4769);
nand U5456 (N_5456,N_4583,N_4058);
xnor U5457 (N_5457,N_4667,N_4341);
nand U5458 (N_5458,N_4454,N_4668);
and U5459 (N_5459,N_4237,N_4526);
or U5460 (N_5460,N_4036,N_4617);
nor U5461 (N_5461,N_4739,N_4439);
or U5462 (N_5462,N_4394,N_4133);
nor U5463 (N_5463,N_4275,N_4381);
and U5464 (N_5464,N_4699,N_4477);
or U5465 (N_5465,N_4578,N_4751);
nand U5466 (N_5466,N_4088,N_4415);
or U5467 (N_5467,N_4042,N_4010);
or U5468 (N_5468,N_4196,N_4776);
or U5469 (N_5469,N_4132,N_4155);
or U5470 (N_5470,N_4156,N_4302);
nand U5471 (N_5471,N_4435,N_4219);
and U5472 (N_5472,N_4672,N_4068);
or U5473 (N_5473,N_4626,N_4753);
or U5474 (N_5474,N_4735,N_4163);
nor U5475 (N_5475,N_4239,N_4165);
nand U5476 (N_5476,N_4347,N_4092);
and U5477 (N_5477,N_4339,N_4260);
or U5478 (N_5478,N_4368,N_4218);
or U5479 (N_5479,N_4178,N_4565);
nand U5480 (N_5480,N_4240,N_4166);
nor U5481 (N_5481,N_4769,N_4681);
nor U5482 (N_5482,N_4003,N_4436);
nand U5483 (N_5483,N_4257,N_4261);
nand U5484 (N_5484,N_4489,N_4091);
and U5485 (N_5485,N_4262,N_4675);
and U5486 (N_5486,N_4122,N_4213);
nor U5487 (N_5487,N_4474,N_4151);
and U5488 (N_5488,N_4676,N_4075);
or U5489 (N_5489,N_4153,N_4737);
nor U5490 (N_5490,N_4563,N_4787);
nor U5491 (N_5491,N_4117,N_4700);
or U5492 (N_5492,N_4716,N_4779);
or U5493 (N_5493,N_4145,N_4796);
and U5494 (N_5494,N_4154,N_4251);
or U5495 (N_5495,N_4288,N_4338);
nor U5496 (N_5496,N_4385,N_4485);
and U5497 (N_5497,N_4746,N_4695);
or U5498 (N_5498,N_4085,N_4775);
nand U5499 (N_5499,N_4048,N_4656);
or U5500 (N_5500,N_4123,N_4538);
nor U5501 (N_5501,N_4135,N_4383);
or U5502 (N_5502,N_4442,N_4740);
or U5503 (N_5503,N_4015,N_4783);
xor U5504 (N_5504,N_4443,N_4408);
and U5505 (N_5505,N_4167,N_4252);
nor U5506 (N_5506,N_4116,N_4303);
nand U5507 (N_5507,N_4201,N_4262);
nand U5508 (N_5508,N_4337,N_4232);
nand U5509 (N_5509,N_4619,N_4722);
or U5510 (N_5510,N_4290,N_4334);
nand U5511 (N_5511,N_4025,N_4534);
and U5512 (N_5512,N_4436,N_4548);
and U5513 (N_5513,N_4539,N_4742);
and U5514 (N_5514,N_4437,N_4049);
nor U5515 (N_5515,N_4030,N_4755);
and U5516 (N_5516,N_4492,N_4504);
and U5517 (N_5517,N_4552,N_4212);
and U5518 (N_5518,N_4040,N_4449);
and U5519 (N_5519,N_4742,N_4283);
or U5520 (N_5520,N_4109,N_4230);
and U5521 (N_5521,N_4100,N_4467);
nand U5522 (N_5522,N_4321,N_4265);
and U5523 (N_5523,N_4278,N_4131);
nand U5524 (N_5524,N_4490,N_4397);
nor U5525 (N_5525,N_4350,N_4628);
nor U5526 (N_5526,N_4717,N_4325);
nand U5527 (N_5527,N_4514,N_4153);
and U5528 (N_5528,N_4394,N_4309);
or U5529 (N_5529,N_4781,N_4486);
and U5530 (N_5530,N_4790,N_4376);
and U5531 (N_5531,N_4646,N_4015);
or U5532 (N_5532,N_4536,N_4175);
or U5533 (N_5533,N_4651,N_4733);
and U5534 (N_5534,N_4110,N_4626);
or U5535 (N_5535,N_4769,N_4514);
and U5536 (N_5536,N_4469,N_4020);
and U5537 (N_5537,N_4676,N_4188);
nor U5538 (N_5538,N_4349,N_4175);
and U5539 (N_5539,N_4653,N_4027);
nand U5540 (N_5540,N_4267,N_4092);
nand U5541 (N_5541,N_4196,N_4187);
or U5542 (N_5542,N_4215,N_4479);
nand U5543 (N_5543,N_4338,N_4221);
or U5544 (N_5544,N_4602,N_4119);
and U5545 (N_5545,N_4732,N_4775);
or U5546 (N_5546,N_4357,N_4016);
or U5547 (N_5547,N_4517,N_4246);
or U5548 (N_5548,N_4041,N_4415);
or U5549 (N_5549,N_4762,N_4503);
and U5550 (N_5550,N_4474,N_4119);
nor U5551 (N_5551,N_4665,N_4409);
and U5552 (N_5552,N_4380,N_4711);
or U5553 (N_5553,N_4318,N_4675);
nor U5554 (N_5554,N_4069,N_4438);
nand U5555 (N_5555,N_4386,N_4668);
and U5556 (N_5556,N_4062,N_4091);
nand U5557 (N_5557,N_4521,N_4261);
nand U5558 (N_5558,N_4298,N_4242);
or U5559 (N_5559,N_4449,N_4687);
nand U5560 (N_5560,N_4007,N_4530);
or U5561 (N_5561,N_4301,N_4110);
and U5562 (N_5562,N_4070,N_4213);
and U5563 (N_5563,N_4339,N_4124);
or U5564 (N_5564,N_4633,N_4395);
and U5565 (N_5565,N_4083,N_4576);
nor U5566 (N_5566,N_4630,N_4360);
nor U5567 (N_5567,N_4276,N_4649);
nor U5568 (N_5568,N_4086,N_4731);
and U5569 (N_5569,N_4474,N_4273);
and U5570 (N_5570,N_4626,N_4734);
or U5571 (N_5571,N_4127,N_4733);
nand U5572 (N_5572,N_4762,N_4704);
or U5573 (N_5573,N_4057,N_4627);
and U5574 (N_5574,N_4697,N_4274);
nand U5575 (N_5575,N_4665,N_4293);
nor U5576 (N_5576,N_4226,N_4097);
nand U5577 (N_5577,N_4783,N_4688);
xor U5578 (N_5578,N_4633,N_4071);
or U5579 (N_5579,N_4651,N_4242);
nand U5580 (N_5580,N_4508,N_4136);
nor U5581 (N_5581,N_4055,N_4187);
and U5582 (N_5582,N_4287,N_4586);
or U5583 (N_5583,N_4723,N_4633);
or U5584 (N_5584,N_4135,N_4130);
nand U5585 (N_5585,N_4160,N_4238);
nand U5586 (N_5586,N_4184,N_4740);
nand U5587 (N_5587,N_4523,N_4505);
and U5588 (N_5588,N_4094,N_4024);
or U5589 (N_5589,N_4574,N_4232);
or U5590 (N_5590,N_4362,N_4014);
or U5591 (N_5591,N_4198,N_4190);
nor U5592 (N_5592,N_4611,N_4541);
nand U5593 (N_5593,N_4651,N_4664);
nor U5594 (N_5594,N_4304,N_4341);
nand U5595 (N_5595,N_4311,N_4098);
or U5596 (N_5596,N_4084,N_4504);
nand U5597 (N_5597,N_4038,N_4590);
nand U5598 (N_5598,N_4032,N_4579);
or U5599 (N_5599,N_4151,N_4212);
nand U5600 (N_5600,N_4954,N_5057);
nor U5601 (N_5601,N_5165,N_5573);
nor U5602 (N_5602,N_5234,N_5504);
or U5603 (N_5603,N_5264,N_4835);
nor U5604 (N_5604,N_4976,N_4843);
nor U5605 (N_5605,N_5408,N_4983);
or U5606 (N_5606,N_5021,N_5169);
or U5607 (N_5607,N_4864,N_5113);
nand U5608 (N_5608,N_4827,N_5235);
nor U5609 (N_5609,N_5214,N_5503);
or U5610 (N_5610,N_5424,N_5252);
or U5611 (N_5611,N_5281,N_4850);
and U5612 (N_5612,N_5293,N_5501);
nor U5613 (N_5613,N_5413,N_5362);
and U5614 (N_5614,N_4854,N_5225);
or U5615 (N_5615,N_5376,N_4979);
or U5616 (N_5616,N_5120,N_5472);
nand U5617 (N_5617,N_5114,N_5555);
nand U5618 (N_5618,N_4956,N_5195);
and U5619 (N_5619,N_5525,N_4831);
and U5620 (N_5620,N_5529,N_4806);
or U5621 (N_5621,N_5290,N_5218);
nor U5622 (N_5622,N_5550,N_5422);
nand U5623 (N_5623,N_4987,N_5453);
nor U5624 (N_5624,N_4945,N_5368);
and U5625 (N_5625,N_5521,N_5464);
and U5626 (N_5626,N_5569,N_4840);
and U5627 (N_5627,N_5013,N_5539);
or U5628 (N_5628,N_5260,N_5327);
nand U5629 (N_5629,N_5510,N_5534);
and U5630 (N_5630,N_5032,N_5219);
nor U5631 (N_5631,N_5551,N_5258);
xnor U5632 (N_5632,N_4959,N_4994);
or U5633 (N_5633,N_5434,N_5243);
nor U5634 (N_5634,N_4950,N_4800);
xor U5635 (N_5635,N_4975,N_5331);
nor U5636 (N_5636,N_5035,N_5137);
and U5637 (N_5637,N_5296,N_5076);
nand U5638 (N_5638,N_5066,N_5152);
and U5639 (N_5639,N_4995,N_5528);
nor U5640 (N_5640,N_5392,N_4890);
and U5641 (N_5641,N_5109,N_5536);
nor U5642 (N_5642,N_5179,N_5340);
nor U5643 (N_5643,N_5242,N_4955);
and U5644 (N_5644,N_4962,N_4913);
or U5645 (N_5645,N_5479,N_4927);
nand U5646 (N_5646,N_5344,N_4918);
nor U5647 (N_5647,N_5565,N_5090);
or U5648 (N_5648,N_5053,N_5207);
nor U5649 (N_5649,N_5126,N_5583);
and U5650 (N_5650,N_5108,N_5423);
or U5651 (N_5651,N_5305,N_5028);
nand U5652 (N_5652,N_4924,N_5564);
and U5653 (N_5653,N_5485,N_5083);
nor U5654 (N_5654,N_5025,N_5072);
nor U5655 (N_5655,N_5325,N_5261);
nor U5656 (N_5656,N_5415,N_4919);
nor U5657 (N_5657,N_5540,N_5561);
nand U5658 (N_5658,N_4804,N_5236);
or U5659 (N_5659,N_5224,N_5213);
nand U5660 (N_5660,N_5597,N_5102);
and U5661 (N_5661,N_5315,N_5123);
nor U5662 (N_5662,N_5342,N_4882);
nand U5663 (N_5663,N_4920,N_4822);
and U5664 (N_5664,N_5526,N_4928);
nand U5665 (N_5665,N_4915,N_4977);
nor U5666 (N_5666,N_4951,N_5239);
and U5667 (N_5667,N_5462,N_5011);
nor U5668 (N_5668,N_5227,N_5567);
nand U5669 (N_5669,N_5447,N_4925);
and U5670 (N_5670,N_5221,N_5100);
nand U5671 (N_5671,N_5240,N_5187);
and U5672 (N_5672,N_4938,N_4974);
and U5673 (N_5673,N_5105,N_5267);
and U5674 (N_5674,N_5420,N_5382);
nand U5675 (N_5675,N_5578,N_5506);
and U5676 (N_5676,N_4997,N_5532);
or U5677 (N_5677,N_5067,N_4949);
or U5678 (N_5678,N_5377,N_5553);
and U5679 (N_5679,N_5388,N_4874);
or U5680 (N_5680,N_5118,N_5353);
nand U5681 (N_5681,N_4818,N_5458);
and U5682 (N_5682,N_4978,N_4813);
nand U5683 (N_5683,N_5358,N_5301);
nand U5684 (N_5684,N_5265,N_5037);
nand U5685 (N_5685,N_5444,N_4873);
and U5686 (N_5686,N_5049,N_4923);
or U5687 (N_5687,N_4847,N_5404);
nor U5688 (N_5688,N_5463,N_5093);
and U5689 (N_5689,N_4887,N_5369);
and U5690 (N_5690,N_5217,N_5593);
or U5691 (N_5691,N_5473,N_5257);
nor U5692 (N_5692,N_5098,N_5289);
nor U5693 (N_5693,N_5212,N_5470);
nand U5694 (N_5694,N_4893,N_5156);
and U5695 (N_5695,N_5520,N_5186);
nor U5696 (N_5696,N_5365,N_5394);
nand U5697 (N_5697,N_5230,N_4870);
nor U5698 (N_5698,N_5367,N_4931);
and U5699 (N_5699,N_5441,N_5096);
nand U5700 (N_5700,N_4972,N_4914);
nor U5701 (N_5701,N_4941,N_5074);
nand U5702 (N_5702,N_5581,N_4940);
and U5703 (N_5703,N_5129,N_4869);
or U5704 (N_5704,N_5385,N_4985);
nand U5705 (N_5705,N_5507,N_5428);
nand U5706 (N_5706,N_4871,N_5188);
and U5707 (N_5707,N_5192,N_4932);
or U5708 (N_5708,N_5176,N_5405);
and U5709 (N_5709,N_5497,N_5430);
or U5710 (N_5710,N_5223,N_5416);
nor U5711 (N_5711,N_4820,N_5446);
nand U5712 (N_5712,N_5081,N_5039);
nor U5713 (N_5713,N_4982,N_5101);
nor U5714 (N_5714,N_5598,N_5075);
and U5715 (N_5715,N_5406,N_5518);
nand U5716 (N_5716,N_4990,N_5249);
and U5717 (N_5717,N_4910,N_5489);
nand U5718 (N_5718,N_5030,N_5560);
nand U5719 (N_5719,N_5373,N_4848);
or U5720 (N_5720,N_5208,N_5517);
nor U5721 (N_5721,N_5095,N_5233);
or U5722 (N_5722,N_5487,N_5266);
nand U5723 (N_5723,N_4898,N_5397);
and U5724 (N_5724,N_5492,N_5481);
and U5725 (N_5725,N_5566,N_5092);
nand U5726 (N_5726,N_5542,N_5078);
nand U5727 (N_5727,N_5513,N_5454);
nand U5728 (N_5728,N_5117,N_5171);
or U5729 (N_5729,N_4885,N_5448);
and U5730 (N_5730,N_5229,N_4842);
nor U5731 (N_5731,N_5070,N_5425);
or U5732 (N_5732,N_5094,N_5545);
and U5733 (N_5733,N_5194,N_5193);
nand U5734 (N_5734,N_5041,N_5461);
or U5735 (N_5735,N_5563,N_4971);
nand U5736 (N_5736,N_5482,N_5357);
or U5737 (N_5737,N_4826,N_5595);
or U5738 (N_5738,N_5309,N_5389);
or U5739 (N_5739,N_5549,N_4845);
nand U5740 (N_5740,N_5157,N_5530);
nand U5741 (N_5741,N_5390,N_4830);
nor U5742 (N_5742,N_5572,N_4879);
nor U5743 (N_5743,N_5255,N_5148);
nor U5744 (N_5744,N_5299,N_5414);
nand U5745 (N_5745,N_5269,N_4872);
and U5746 (N_5746,N_5062,N_5048);
or U5747 (N_5747,N_4996,N_5263);
or U5748 (N_5748,N_5082,N_5106);
nor U5749 (N_5749,N_5379,N_5181);
or U5750 (N_5750,N_5211,N_5477);
nor U5751 (N_5751,N_5274,N_5310);
nor U5752 (N_5752,N_5499,N_5135);
xor U5753 (N_5753,N_5185,N_5403);
nand U5754 (N_5754,N_5571,N_5437);
or U5755 (N_5755,N_5173,N_5537);
xor U5756 (N_5756,N_4894,N_5402);
nand U5757 (N_5757,N_4935,N_4895);
or U5758 (N_5758,N_5189,N_5144);
and U5759 (N_5759,N_5014,N_5204);
nor U5760 (N_5760,N_4947,N_5084);
nand U5761 (N_5761,N_5199,N_5089);
nand U5762 (N_5762,N_5107,N_5352);
and U5763 (N_5763,N_5064,N_5139);
nor U5764 (N_5764,N_4829,N_5330);
and U5765 (N_5765,N_5311,N_5427);
nor U5766 (N_5766,N_4837,N_5543);
and U5767 (N_5767,N_5411,N_5387);
nand U5768 (N_5768,N_4909,N_5099);
and U5769 (N_5769,N_5245,N_5592);
nand U5770 (N_5770,N_4967,N_5280);
and U5771 (N_5771,N_4917,N_5505);
nor U5772 (N_5772,N_5004,N_5418);
and U5773 (N_5773,N_5329,N_4846);
or U5774 (N_5774,N_5457,N_5574);
nor U5775 (N_5775,N_5326,N_5548);
nor U5776 (N_5776,N_5132,N_5237);
nand U5777 (N_5777,N_5085,N_4816);
or U5778 (N_5778,N_5486,N_5121);
nand U5779 (N_5779,N_5097,N_5409);
and U5780 (N_5780,N_5306,N_4828);
nor U5781 (N_5781,N_5196,N_5334);
nor U5782 (N_5782,N_5375,N_5345);
nand U5783 (N_5783,N_5439,N_5210);
nor U5784 (N_5784,N_5559,N_5412);
or U5785 (N_5785,N_5313,N_5466);
nand U5786 (N_5786,N_5359,N_5314);
nand U5787 (N_5787,N_5450,N_5577);
nand U5788 (N_5788,N_4908,N_4888);
or U5789 (N_5789,N_4948,N_4933);
nand U5790 (N_5790,N_4992,N_5174);
or U5791 (N_5791,N_5594,N_5511);
nand U5792 (N_5792,N_5295,N_4892);
nand U5793 (N_5793,N_5146,N_5287);
or U5794 (N_5794,N_5465,N_5585);
nor U5795 (N_5795,N_5378,N_5546);
nand U5796 (N_5796,N_5271,N_5339);
nor U5797 (N_5797,N_5086,N_4906);
and U5798 (N_5798,N_4939,N_5206);
and U5799 (N_5799,N_5459,N_4881);
and U5800 (N_5800,N_5442,N_5562);
or U5801 (N_5801,N_5319,N_5300);
nor U5802 (N_5802,N_5502,N_5535);
or U5803 (N_5803,N_5080,N_5127);
and U5804 (N_5804,N_4876,N_4960);
or U5805 (N_5805,N_4946,N_4862);
or U5806 (N_5806,N_4905,N_5209);
nor U5807 (N_5807,N_5145,N_4942);
nand U5808 (N_5808,N_5159,N_5163);
or U5809 (N_5809,N_4926,N_5393);
nor U5810 (N_5810,N_5480,N_5079);
nor U5811 (N_5811,N_5200,N_5527);
nand U5812 (N_5812,N_5318,N_5508);
nor U5813 (N_5813,N_5308,N_5356);
or U5814 (N_5814,N_5116,N_5069);
nand U5815 (N_5815,N_5302,N_5468);
nand U5816 (N_5816,N_5045,N_5033);
or U5817 (N_5817,N_4814,N_5366);
nor U5818 (N_5818,N_4981,N_5488);
nand U5819 (N_5819,N_5575,N_5130);
nor U5820 (N_5820,N_4904,N_4877);
nor U5821 (N_5821,N_5040,N_5364);
nand U5822 (N_5822,N_5162,N_5347);
and U5823 (N_5823,N_4808,N_5350);
nor U5824 (N_5824,N_5558,N_5346);
and U5825 (N_5825,N_4802,N_5104);
nor U5826 (N_5826,N_4878,N_5003);
or U5827 (N_5827,N_5321,N_5278);
or U5828 (N_5828,N_4821,N_5476);
and U5829 (N_5829,N_5250,N_4824);
nor U5830 (N_5830,N_5410,N_5401);
and U5831 (N_5831,N_5044,N_5332);
nand U5832 (N_5832,N_5544,N_5320);
and U5833 (N_5833,N_5228,N_5125);
and U5834 (N_5834,N_5022,N_5361);
and U5835 (N_5835,N_5134,N_4834);
or U5836 (N_5836,N_4853,N_5582);
nand U5837 (N_5837,N_5531,N_5110);
nand U5838 (N_5838,N_5399,N_5478);
nand U5839 (N_5839,N_5024,N_5043);
nor U5840 (N_5840,N_5167,N_5141);
nor U5841 (N_5841,N_5026,N_4969);
or U5842 (N_5842,N_4986,N_4807);
nand U5843 (N_5843,N_5036,N_5498);
and U5844 (N_5844,N_5262,N_5142);
xor U5845 (N_5845,N_4851,N_5231);
or U5846 (N_5846,N_5433,N_4810);
nand U5847 (N_5847,N_5533,N_5452);
nor U5848 (N_5848,N_5500,N_5493);
or U5849 (N_5849,N_4856,N_5432);
nand U5850 (N_5850,N_5371,N_5061);
nand U5851 (N_5851,N_4823,N_4998);
nor U5852 (N_5852,N_5407,N_4833);
and U5853 (N_5853,N_5060,N_5580);
nand U5854 (N_5854,N_5522,N_5557);
and U5855 (N_5855,N_4957,N_4859);
nand U5856 (N_5856,N_5133,N_5323);
nor U5857 (N_5857,N_4943,N_5475);
or U5858 (N_5858,N_5283,N_5455);
and U5859 (N_5859,N_4964,N_4965);
nand U5860 (N_5860,N_5435,N_5354);
nor U5861 (N_5861,N_5286,N_5016);
nand U5862 (N_5862,N_5587,N_4973);
nand U5863 (N_5863,N_5491,N_5259);
nor U5864 (N_5864,N_5222,N_5324);
or U5865 (N_5865,N_4858,N_5031);
nor U5866 (N_5866,N_5547,N_5417);
nor U5867 (N_5867,N_5068,N_5570);
nor U5868 (N_5868,N_4841,N_5147);
or U5869 (N_5869,N_4832,N_5523);
or U5870 (N_5870,N_5005,N_5182);
or U5871 (N_5871,N_5322,N_5248);
or U5872 (N_5872,N_5282,N_5449);
nand U5873 (N_5873,N_5277,N_4863);
or U5874 (N_5874,N_4901,N_5483);
or U5875 (N_5875,N_5002,N_5077);
or U5876 (N_5876,N_5328,N_5576);
nand U5877 (N_5877,N_4891,N_5164);
nand U5878 (N_5878,N_5556,N_5112);
nand U5879 (N_5879,N_5538,N_5268);
nor U5880 (N_5880,N_5512,N_5056);
nor U5881 (N_5881,N_5177,N_5333);
xnor U5882 (N_5882,N_5238,N_5552);
and U5883 (N_5883,N_5124,N_5276);
nor U5884 (N_5884,N_5019,N_5579);
and U5885 (N_5885,N_5275,N_5136);
or U5886 (N_5886,N_5190,N_5029);
nand U5887 (N_5887,N_5297,N_5015);
nor U5888 (N_5888,N_5111,N_4817);
xnor U5889 (N_5889,N_5215,N_4903);
or U5890 (N_5890,N_5241,N_5119);
nand U5891 (N_5891,N_5451,N_4825);
and U5892 (N_5892,N_5027,N_5599);
and U5893 (N_5893,N_5380,N_5471);
and U5894 (N_5894,N_5284,N_4897);
nand U5895 (N_5895,N_4968,N_5584);
nand U5896 (N_5896,N_5372,N_4989);
nand U5897 (N_5897,N_5063,N_5303);
and U5898 (N_5898,N_5051,N_4902);
nor U5899 (N_5899,N_5055,N_5596);
or U5900 (N_5900,N_5370,N_5205);
and U5901 (N_5901,N_5059,N_4855);
or U5902 (N_5902,N_5256,N_5184);
xnor U5903 (N_5903,N_5253,N_5158);
nor U5904 (N_5904,N_4849,N_4911);
nor U5905 (N_5905,N_5247,N_5515);
or U5906 (N_5906,N_5589,N_4819);
nand U5907 (N_5907,N_5140,N_5054);
or U5908 (N_5908,N_4999,N_5456);
or U5909 (N_5909,N_5178,N_5431);
and U5910 (N_5910,N_5443,N_4934);
nand U5911 (N_5911,N_4868,N_5467);
nor U5912 (N_5912,N_5091,N_5153);
nor U5913 (N_5913,N_5460,N_4875);
nor U5914 (N_5914,N_5202,N_4936);
and U5915 (N_5915,N_5317,N_5201);
nor U5916 (N_5916,N_5509,N_5272);
or U5917 (N_5917,N_4812,N_5285);
nor U5918 (N_5918,N_4839,N_4860);
or U5919 (N_5919,N_5586,N_5519);
nand U5920 (N_5920,N_5143,N_4889);
nand U5921 (N_5921,N_4912,N_4899);
nor U5922 (N_5922,N_5590,N_5343);
and U5923 (N_5923,N_5484,N_5440);
and U5924 (N_5924,N_5047,N_5383);
and U5925 (N_5925,N_4861,N_4866);
nand U5926 (N_5926,N_4937,N_5175);
and U5927 (N_5927,N_5254,N_5294);
and U5928 (N_5928,N_5338,N_4966);
nor U5929 (N_5929,N_5588,N_5020);
xnor U5930 (N_5930,N_5349,N_4884);
nand U5931 (N_5931,N_4961,N_5216);
or U5932 (N_5932,N_5150,N_5042);
or U5933 (N_5933,N_5203,N_4993);
nand U5934 (N_5934,N_5273,N_5400);
and U5935 (N_5935,N_4991,N_5128);
nor U5936 (N_5936,N_5138,N_5469);
nor U5937 (N_5937,N_5474,N_5052);
nand U5938 (N_5938,N_5046,N_4836);
nor U5939 (N_5939,N_4809,N_5154);
nor U5940 (N_5940,N_5220,N_5183);
nor U5941 (N_5941,N_4970,N_4980);
and U5942 (N_5942,N_4865,N_5087);
nand U5943 (N_5943,N_5151,N_5017);
or U5944 (N_5944,N_5298,N_5426);
or U5945 (N_5945,N_5251,N_5244);
and U5946 (N_5946,N_4900,N_5554);
and U5947 (N_5947,N_5155,N_4811);
nand U5948 (N_5948,N_5270,N_5149);
nor U5949 (N_5949,N_5291,N_4944);
and U5950 (N_5950,N_4922,N_4886);
nand U5951 (N_5951,N_5312,N_5168);
or U5952 (N_5952,N_5341,N_5058);
and U5953 (N_5953,N_4805,N_5514);
and U5954 (N_5954,N_5073,N_5384);
or U5955 (N_5955,N_5386,N_5122);
nor U5956 (N_5956,N_5419,N_5348);
nor U5957 (N_5957,N_4963,N_5337);
nand U5958 (N_5958,N_5006,N_5292);
nand U5959 (N_5959,N_5191,N_5018);
nand U5960 (N_5960,N_5496,N_5131);
and U5961 (N_5961,N_4916,N_4930);
nand U5962 (N_5962,N_5351,N_4958);
nor U5963 (N_5963,N_5232,N_5065);
nand U5964 (N_5964,N_5429,N_5335);
or U5965 (N_5965,N_5494,N_5395);
nor U5966 (N_5966,N_5197,N_5246);
nand U5967 (N_5967,N_5304,N_5023);
and U5968 (N_5968,N_5038,N_5288);
nand U5969 (N_5969,N_5172,N_5445);
nand U5970 (N_5970,N_5421,N_5363);
or U5971 (N_5971,N_5307,N_5007);
nor U5972 (N_5972,N_5071,N_5170);
nor U5973 (N_5973,N_5226,N_5568);
nand U5974 (N_5974,N_4815,N_4896);
and U5975 (N_5975,N_5115,N_4907);
nand U5976 (N_5976,N_5516,N_4857);
or U5977 (N_5977,N_5398,N_4952);
and U5978 (N_5978,N_5591,N_4838);
nand U5979 (N_5979,N_4852,N_5008);
nand U5980 (N_5980,N_5166,N_4801);
or U5981 (N_5981,N_5490,N_5541);
nor U5982 (N_5982,N_4803,N_5381);
nand U5983 (N_5983,N_5198,N_5438);
nor U5984 (N_5984,N_5279,N_5009);
or U5985 (N_5985,N_4844,N_5160);
nand U5986 (N_5986,N_5050,N_5524);
nand U5987 (N_5987,N_5000,N_5336);
and U5988 (N_5988,N_4988,N_4867);
nand U5989 (N_5989,N_4984,N_5374);
nor U5990 (N_5990,N_4953,N_5001);
and U5991 (N_5991,N_5103,N_5010);
nor U5992 (N_5992,N_5034,N_5355);
nor U5993 (N_5993,N_5180,N_5391);
or U5994 (N_5994,N_5088,N_5436);
or U5995 (N_5995,N_4929,N_5495);
or U5996 (N_5996,N_4883,N_5161);
nor U5997 (N_5997,N_5316,N_4921);
nor U5998 (N_5998,N_5012,N_5360);
or U5999 (N_5999,N_4880,N_5396);
or U6000 (N_6000,N_5585,N_4992);
nand U6001 (N_6001,N_5077,N_5260);
nand U6002 (N_6002,N_5227,N_5423);
or U6003 (N_6003,N_4932,N_4985);
and U6004 (N_6004,N_5377,N_4933);
or U6005 (N_6005,N_5219,N_5453);
and U6006 (N_6006,N_5541,N_5533);
xnor U6007 (N_6007,N_5172,N_4852);
nand U6008 (N_6008,N_5296,N_5589);
and U6009 (N_6009,N_5319,N_5168);
or U6010 (N_6010,N_5587,N_5041);
and U6011 (N_6011,N_5403,N_5215);
or U6012 (N_6012,N_5524,N_5430);
nor U6013 (N_6013,N_5505,N_5395);
or U6014 (N_6014,N_5266,N_5037);
nor U6015 (N_6015,N_4925,N_5098);
nand U6016 (N_6016,N_4826,N_5312);
nor U6017 (N_6017,N_5093,N_4884);
or U6018 (N_6018,N_4832,N_5213);
or U6019 (N_6019,N_5546,N_5346);
nor U6020 (N_6020,N_5354,N_4826);
and U6021 (N_6021,N_5161,N_5105);
nand U6022 (N_6022,N_5527,N_5402);
nor U6023 (N_6023,N_4854,N_5253);
nand U6024 (N_6024,N_5050,N_5261);
nand U6025 (N_6025,N_5148,N_5191);
nor U6026 (N_6026,N_4958,N_5558);
nand U6027 (N_6027,N_5278,N_5528);
xor U6028 (N_6028,N_5234,N_5283);
nor U6029 (N_6029,N_5215,N_5018);
or U6030 (N_6030,N_5477,N_4822);
nor U6031 (N_6031,N_4931,N_5227);
and U6032 (N_6032,N_5486,N_5333);
and U6033 (N_6033,N_5097,N_5306);
nand U6034 (N_6034,N_4953,N_5094);
nand U6035 (N_6035,N_4961,N_5102);
or U6036 (N_6036,N_5311,N_4953);
nand U6037 (N_6037,N_5181,N_4921);
nand U6038 (N_6038,N_4906,N_5089);
nor U6039 (N_6039,N_5528,N_5140);
or U6040 (N_6040,N_5258,N_5152);
nor U6041 (N_6041,N_5550,N_5483);
nand U6042 (N_6042,N_5387,N_4937);
nor U6043 (N_6043,N_5335,N_4812);
nand U6044 (N_6044,N_5260,N_5203);
or U6045 (N_6045,N_5194,N_5370);
nand U6046 (N_6046,N_4809,N_5138);
and U6047 (N_6047,N_5144,N_5224);
nor U6048 (N_6048,N_4800,N_5119);
or U6049 (N_6049,N_5487,N_5185);
and U6050 (N_6050,N_5097,N_5322);
nor U6051 (N_6051,N_5450,N_5026);
and U6052 (N_6052,N_5325,N_5429);
nand U6053 (N_6053,N_4810,N_4910);
nand U6054 (N_6054,N_5440,N_4998);
nand U6055 (N_6055,N_5125,N_4920);
and U6056 (N_6056,N_5169,N_5320);
nor U6057 (N_6057,N_5289,N_5415);
nor U6058 (N_6058,N_4990,N_5300);
nand U6059 (N_6059,N_5330,N_5597);
nor U6060 (N_6060,N_5584,N_4978);
or U6061 (N_6061,N_5417,N_4959);
and U6062 (N_6062,N_4947,N_5030);
or U6063 (N_6063,N_4801,N_5308);
nor U6064 (N_6064,N_5386,N_4915);
nor U6065 (N_6065,N_5598,N_5177);
nor U6066 (N_6066,N_5201,N_5292);
nand U6067 (N_6067,N_5245,N_4830);
or U6068 (N_6068,N_5487,N_4995);
or U6069 (N_6069,N_5291,N_5149);
and U6070 (N_6070,N_4906,N_5266);
and U6071 (N_6071,N_4880,N_5459);
nand U6072 (N_6072,N_5246,N_5153);
and U6073 (N_6073,N_5474,N_5566);
and U6074 (N_6074,N_5516,N_5073);
or U6075 (N_6075,N_5364,N_4910);
and U6076 (N_6076,N_5258,N_5015);
and U6077 (N_6077,N_5233,N_5491);
and U6078 (N_6078,N_5374,N_5599);
and U6079 (N_6079,N_4812,N_5310);
nand U6080 (N_6080,N_4858,N_4869);
and U6081 (N_6081,N_5105,N_5187);
and U6082 (N_6082,N_5579,N_4859);
and U6083 (N_6083,N_5013,N_5110);
or U6084 (N_6084,N_4945,N_5052);
nor U6085 (N_6085,N_4816,N_5249);
nand U6086 (N_6086,N_5213,N_5587);
nor U6087 (N_6087,N_5259,N_5514);
nor U6088 (N_6088,N_5018,N_4983);
nor U6089 (N_6089,N_5593,N_5491);
nor U6090 (N_6090,N_5314,N_4919);
nor U6091 (N_6091,N_5060,N_5157);
or U6092 (N_6092,N_5046,N_5004);
or U6093 (N_6093,N_4964,N_5451);
or U6094 (N_6094,N_5134,N_5166);
nand U6095 (N_6095,N_5017,N_5452);
or U6096 (N_6096,N_5205,N_4906);
or U6097 (N_6097,N_5004,N_5434);
and U6098 (N_6098,N_5165,N_5157);
nor U6099 (N_6099,N_5227,N_5018);
nand U6100 (N_6100,N_5152,N_5196);
nand U6101 (N_6101,N_5168,N_5438);
and U6102 (N_6102,N_5211,N_5283);
and U6103 (N_6103,N_5079,N_5560);
or U6104 (N_6104,N_4819,N_4813);
nand U6105 (N_6105,N_5058,N_5564);
or U6106 (N_6106,N_5225,N_4890);
nand U6107 (N_6107,N_5521,N_5500);
nor U6108 (N_6108,N_5230,N_5112);
nand U6109 (N_6109,N_4879,N_4801);
and U6110 (N_6110,N_5076,N_5586);
nand U6111 (N_6111,N_5095,N_5520);
nand U6112 (N_6112,N_5095,N_4984);
nor U6113 (N_6113,N_5009,N_4907);
nand U6114 (N_6114,N_5107,N_5222);
xor U6115 (N_6115,N_5451,N_4833);
nand U6116 (N_6116,N_5389,N_5368);
and U6117 (N_6117,N_5067,N_5197);
and U6118 (N_6118,N_5156,N_5051);
and U6119 (N_6119,N_5232,N_4884);
nor U6120 (N_6120,N_4822,N_5098);
nand U6121 (N_6121,N_4948,N_5492);
or U6122 (N_6122,N_5592,N_5052);
nor U6123 (N_6123,N_5390,N_5037);
and U6124 (N_6124,N_5183,N_4995);
nand U6125 (N_6125,N_5063,N_5260);
and U6126 (N_6126,N_5153,N_5282);
and U6127 (N_6127,N_5362,N_5203);
nor U6128 (N_6128,N_4944,N_4965);
nand U6129 (N_6129,N_5385,N_5487);
and U6130 (N_6130,N_5403,N_5024);
or U6131 (N_6131,N_5559,N_5423);
nand U6132 (N_6132,N_5023,N_4801);
xnor U6133 (N_6133,N_4813,N_5270);
nor U6134 (N_6134,N_5373,N_5437);
and U6135 (N_6135,N_5311,N_5419);
nor U6136 (N_6136,N_5135,N_5589);
and U6137 (N_6137,N_5512,N_5030);
nand U6138 (N_6138,N_4899,N_5072);
nor U6139 (N_6139,N_5139,N_5023);
nand U6140 (N_6140,N_5224,N_5370);
or U6141 (N_6141,N_4812,N_5579);
nand U6142 (N_6142,N_5006,N_5041);
and U6143 (N_6143,N_5408,N_5151);
and U6144 (N_6144,N_4933,N_5222);
or U6145 (N_6145,N_4963,N_5183);
and U6146 (N_6146,N_5534,N_4950);
nand U6147 (N_6147,N_4803,N_5163);
nor U6148 (N_6148,N_5308,N_5099);
nand U6149 (N_6149,N_5374,N_5226);
or U6150 (N_6150,N_4951,N_4819);
nand U6151 (N_6151,N_4906,N_5384);
nand U6152 (N_6152,N_4816,N_5482);
nor U6153 (N_6153,N_5563,N_5346);
or U6154 (N_6154,N_5113,N_5206);
nor U6155 (N_6155,N_5542,N_5141);
or U6156 (N_6156,N_4832,N_5333);
nand U6157 (N_6157,N_5147,N_5586);
and U6158 (N_6158,N_5271,N_5081);
nand U6159 (N_6159,N_5531,N_5544);
nand U6160 (N_6160,N_5239,N_5031);
and U6161 (N_6161,N_4888,N_5030);
and U6162 (N_6162,N_4915,N_5133);
or U6163 (N_6163,N_5554,N_4814);
or U6164 (N_6164,N_4938,N_5507);
nor U6165 (N_6165,N_4936,N_5404);
or U6166 (N_6166,N_5508,N_4924);
nand U6167 (N_6167,N_4860,N_5580);
nor U6168 (N_6168,N_4875,N_5304);
nand U6169 (N_6169,N_5418,N_5033);
nand U6170 (N_6170,N_5550,N_4970);
nor U6171 (N_6171,N_5461,N_4895);
nand U6172 (N_6172,N_5138,N_4829);
nor U6173 (N_6173,N_4955,N_5009);
or U6174 (N_6174,N_4872,N_5223);
nand U6175 (N_6175,N_5177,N_4990);
and U6176 (N_6176,N_5545,N_5090);
nor U6177 (N_6177,N_5004,N_5436);
and U6178 (N_6178,N_5461,N_5206);
nand U6179 (N_6179,N_4950,N_5075);
nor U6180 (N_6180,N_4992,N_5283);
or U6181 (N_6181,N_4962,N_4938);
and U6182 (N_6182,N_5562,N_5065);
nor U6183 (N_6183,N_5213,N_5300);
and U6184 (N_6184,N_5270,N_5135);
nand U6185 (N_6185,N_5515,N_5106);
and U6186 (N_6186,N_5542,N_5271);
or U6187 (N_6187,N_5277,N_5091);
or U6188 (N_6188,N_5337,N_5236);
and U6189 (N_6189,N_5119,N_5106);
nand U6190 (N_6190,N_5416,N_5090);
and U6191 (N_6191,N_4850,N_4828);
nand U6192 (N_6192,N_5213,N_5478);
and U6193 (N_6193,N_5283,N_4980);
nand U6194 (N_6194,N_5225,N_4929);
nor U6195 (N_6195,N_5117,N_4925);
nor U6196 (N_6196,N_5116,N_5186);
nor U6197 (N_6197,N_5137,N_4841);
nor U6198 (N_6198,N_5165,N_4948);
nand U6199 (N_6199,N_5056,N_5072);
nor U6200 (N_6200,N_5406,N_4842);
nor U6201 (N_6201,N_4846,N_4998);
or U6202 (N_6202,N_5548,N_4825);
and U6203 (N_6203,N_4995,N_5517);
nand U6204 (N_6204,N_5547,N_5020);
nor U6205 (N_6205,N_5015,N_4906);
nor U6206 (N_6206,N_4891,N_5133);
nand U6207 (N_6207,N_5366,N_4806);
nor U6208 (N_6208,N_4955,N_5269);
nor U6209 (N_6209,N_5126,N_5510);
or U6210 (N_6210,N_5483,N_5517);
nor U6211 (N_6211,N_5240,N_5561);
or U6212 (N_6212,N_5583,N_4995);
nand U6213 (N_6213,N_5220,N_5336);
nor U6214 (N_6214,N_5402,N_5121);
or U6215 (N_6215,N_5355,N_5041);
or U6216 (N_6216,N_5448,N_5575);
or U6217 (N_6217,N_5244,N_5570);
or U6218 (N_6218,N_5476,N_5084);
and U6219 (N_6219,N_5231,N_5216);
and U6220 (N_6220,N_5516,N_5338);
nand U6221 (N_6221,N_5028,N_5485);
nand U6222 (N_6222,N_5233,N_5184);
nand U6223 (N_6223,N_5211,N_5537);
or U6224 (N_6224,N_4852,N_5034);
nand U6225 (N_6225,N_5088,N_5396);
and U6226 (N_6226,N_5039,N_5315);
nand U6227 (N_6227,N_4839,N_5238);
nand U6228 (N_6228,N_4915,N_5309);
nor U6229 (N_6229,N_5433,N_5140);
nor U6230 (N_6230,N_5448,N_5431);
nand U6231 (N_6231,N_4914,N_4865);
nand U6232 (N_6232,N_4866,N_5394);
and U6233 (N_6233,N_5085,N_4854);
nand U6234 (N_6234,N_5599,N_4982);
or U6235 (N_6235,N_5507,N_5328);
and U6236 (N_6236,N_5284,N_5041);
nand U6237 (N_6237,N_4903,N_5101);
nor U6238 (N_6238,N_4807,N_5264);
nor U6239 (N_6239,N_4896,N_5091);
nand U6240 (N_6240,N_5574,N_5110);
and U6241 (N_6241,N_4958,N_5424);
nor U6242 (N_6242,N_4833,N_4964);
and U6243 (N_6243,N_5551,N_5572);
or U6244 (N_6244,N_5328,N_4971);
and U6245 (N_6245,N_4987,N_5340);
and U6246 (N_6246,N_5316,N_5161);
and U6247 (N_6247,N_5239,N_5367);
nor U6248 (N_6248,N_5560,N_4990);
nor U6249 (N_6249,N_5310,N_5260);
and U6250 (N_6250,N_5597,N_5183);
and U6251 (N_6251,N_5454,N_4973);
or U6252 (N_6252,N_5125,N_5326);
nand U6253 (N_6253,N_4955,N_4840);
or U6254 (N_6254,N_5118,N_5492);
nand U6255 (N_6255,N_5451,N_5186);
and U6256 (N_6256,N_5290,N_5217);
nand U6257 (N_6257,N_4843,N_4985);
or U6258 (N_6258,N_5440,N_5572);
nor U6259 (N_6259,N_5193,N_5396);
nor U6260 (N_6260,N_5130,N_5241);
or U6261 (N_6261,N_4892,N_5362);
or U6262 (N_6262,N_5541,N_4868);
nand U6263 (N_6263,N_5141,N_5247);
nand U6264 (N_6264,N_4898,N_4992);
nand U6265 (N_6265,N_4857,N_5166);
or U6266 (N_6266,N_5249,N_4911);
nor U6267 (N_6267,N_5242,N_5051);
and U6268 (N_6268,N_4987,N_5118);
nor U6269 (N_6269,N_5595,N_5442);
or U6270 (N_6270,N_4902,N_5437);
nor U6271 (N_6271,N_4911,N_5572);
and U6272 (N_6272,N_4881,N_4913);
nor U6273 (N_6273,N_5089,N_5006);
or U6274 (N_6274,N_5576,N_5534);
nand U6275 (N_6275,N_5333,N_5167);
nor U6276 (N_6276,N_4881,N_5534);
or U6277 (N_6277,N_5223,N_5251);
nor U6278 (N_6278,N_4842,N_4900);
and U6279 (N_6279,N_5297,N_5205);
or U6280 (N_6280,N_5128,N_4954);
nand U6281 (N_6281,N_5217,N_5442);
or U6282 (N_6282,N_5116,N_5088);
nand U6283 (N_6283,N_4821,N_5491);
and U6284 (N_6284,N_5057,N_5494);
and U6285 (N_6285,N_4915,N_5176);
nor U6286 (N_6286,N_5471,N_5003);
nor U6287 (N_6287,N_4870,N_5057);
nor U6288 (N_6288,N_5210,N_5276);
and U6289 (N_6289,N_4921,N_4846);
or U6290 (N_6290,N_5065,N_4947);
or U6291 (N_6291,N_5492,N_5305);
nand U6292 (N_6292,N_5080,N_5280);
and U6293 (N_6293,N_5088,N_4931);
or U6294 (N_6294,N_5334,N_5058);
nand U6295 (N_6295,N_5107,N_4852);
or U6296 (N_6296,N_5036,N_5495);
nor U6297 (N_6297,N_5062,N_5324);
or U6298 (N_6298,N_5347,N_5110);
nor U6299 (N_6299,N_5461,N_5180);
nand U6300 (N_6300,N_5426,N_5129);
nor U6301 (N_6301,N_5214,N_5056);
or U6302 (N_6302,N_5272,N_4859);
and U6303 (N_6303,N_5242,N_4981);
nand U6304 (N_6304,N_5026,N_5411);
nand U6305 (N_6305,N_5477,N_5153);
and U6306 (N_6306,N_5028,N_5374);
nand U6307 (N_6307,N_5353,N_5057);
and U6308 (N_6308,N_4893,N_5175);
nand U6309 (N_6309,N_5101,N_5374);
xnor U6310 (N_6310,N_5183,N_4845);
or U6311 (N_6311,N_4909,N_5242);
or U6312 (N_6312,N_4832,N_5011);
nand U6313 (N_6313,N_5258,N_4825);
nand U6314 (N_6314,N_4920,N_5437);
nor U6315 (N_6315,N_4852,N_5264);
nand U6316 (N_6316,N_5367,N_5103);
or U6317 (N_6317,N_5465,N_5206);
and U6318 (N_6318,N_5393,N_5181);
nand U6319 (N_6319,N_5211,N_5042);
nand U6320 (N_6320,N_5397,N_4917);
nand U6321 (N_6321,N_5205,N_4913);
or U6322 (N_6322,N_5064,N_5117);
nand U6323 (N_6323,N_5102,N_5329);
nand U6324 (N_6324,N_4848,N_5237);
nand U6325 (N_6325,N_5381,N_5167);
or U6326 (N_6326,N_5035,N_5160);
nand U6327 (N_6327,N_5475,N_4863);
nand U6328 (N_6328,N_5521,N_5391);
nor U6329 (N_6329,N_5311,N_5048);
nor U6330 (N_6330,N_4833,N_5450);
or U6331 (N_6331,N_5149,N_5264);
nor U6332 (N_6332,N_5171,N_5519);
or U6333 (N_6333,N_5519,N_5420);
or U6334 (N_6334,N_5257,N_5383);
or U6335 (N_6335,N_5431,N_5544);
nand U6336 (N_6336,N_5581,N_4893);
nor U6337 (N_6337,N_4919,N_5573);
and U6338 (N_6338,N_5187,N_5250);
nand U6339 (N_6339,N_5478,N_5004);
nand U6340 (N_6340,N_4955,N_5444);
nand U6341 (N_6341,N_5118,N_4832);
nor U6342 (N_6342,N_5273,N_5010);
nand U6343 (N_6343,N_5186,N_4830);
nor U6344 (N_6344,N_5057,N_5562);
nor U6345 (N_6345,N_4957,N_5089);
or U6346 (N_6346,N_5239,N_5323);
nand U6347 (N_6347,N_5259,N_5591);
xnor U6348 (N_6348,N_5348,N_5175);
nor U6349 (N_6349,N_5549,N_5365);
nor U6350 (N_6350,N_5314,N_5464);
nor U6351 (N_6351,N_5241,N_5269);
and U6352 (N_6352,N_4943,N_5103);
or U6353 (N_6353,N_5458,N_4839);
or U6354 (N_6354,N_5585,N_5561);
nand U6355 (N_6355,N_5333,N_5476);
nor U6356 (N_6356,N_5390,N_5335);
nand U6357 (N_6357,N_5542,N_5514);
and U6358 (N_6358,N_4973,N_5076);
or U6359 (N_6359,N_5428,N_5499);
or U6360 (N_6360,N_5546,N_5068);
and U6361 (N_6361,N_5352,N_5227);
and U6362 (N_6362,N_5147,N_4817);
nand U6363 (N_6363,N_4851,N_5381);
and U6364 (N_6364,N_5518,N_4951);
and U6365 (N_6365,N_5530,N_5514);
or U6366 (N_6366,N_4992,N_5187);
nor U6367 (N_6367,N_5343,N_5113);
and U6368 (N_6368,N_4853,N_5251);
and U6369 (N_6369,N_5040,N_4964);
and U6370 (N_6370,N_5316,N_5262);
or U6371 (N_6371,N_5040,N_5035);
nand U6372 (N_6372,N_5352,N_5255);
or U6373 (N_6373,N_5019,N_4906);
or U6374 (N_6374,N_5132,N_5516);
or U6375 (N_6375,N_4961,N_5378);
or U6376 (N_6376,N_5276,N_5460);
and U6377 (N_6377,N_4970,N_4857);
nand U6378 (N_6378,N_5574,N_4984);
and U6379 (N_6379,N_5044,N_5209);
or U6380 (N_6380,N_5460,N_4941);
nor U6381 (N_6381,N_4898,N_5319);
and U6382 (N_6382,N_4886,N_4816);
nor U6383 (N_6383,N_5048,N_5444);
and U6384 (N_6384,N_4940,N_4853);
or U6385 (N_6385,N_5118,N_4844);
or U6386 (N_6386,N_5135,N_5091);
and U6387 (N_6387,N_4834,N_4984);
nand U6388 (N_6388,N_5145,N_5460);
xor U6389 (N_6389,N_5186,N_5512);
or U6390 (N_6390,N_5414,N_4914);
nor U6391 (N_6391,N_4897,N_5522);
nor U6392 (N_6392,N_5553,N_4935);
nand U6393 (N_6393,N_4843,N_5219);
or U6394 (N_6394,N_5576,N_5343);
nor U6395 (N_6395,N_5054,N_5507);
nor U6396 (N_6396,N_5183,N_5124);
nand U6397 (N_6397,N_5366,N_4878);
nor U6398 (N_6398,N_5051,N_4813);
nor U6399 (N_6399,N_4910,N_4834);
or U6400 (N_6400,N_5646,N_5934);
or U6401 (N_6401,N_5874,N_5641);
nand U6402 (N_6402,N_5681,N_6167);
nor U6403 (N_6403,N_5910,N_5808);
or U6404 (N_6404,N_6103,N_6014);
and U6405 (N_6405,N_5915,N_5952);
or U6406 (N_6406,N_6079,N_5731);
nor U6407 (N_6407,N_6262,N_5979);
nor U6408 (N_6408,N_6343,N_5601);
nor U6409 (N_6409,N_5827,N_6199);
xnor U6410 (N_6410,N_5961,N_6152);
nor U6411 (N_6411,N_6148,N_6141);
or U6412 (N_6412,N_5656,N_5793);
nor U6413 (N_6413,N_5799,N_6390);
nor U6414 (N_6414,N_6030,N_6312);
nor U6415 (N_6415,N_6234,N_6365);
nor U6416 (N_6416,N_6047,N_5689);
or U6417 (N_6417,N_5992,N_5653);
or U6418 (N_6418,N_6303,N_5691);
nand U6419 (N_6419,N_5813,N_5842);
nor U6420 (N_6420,N_6389,N_5861);
or U6421 (N_6421,N_6092,N_6118);
nand U6422 (N_6422,N_5945,N_5715);
or U6423 (N_6423,N_5790,N_6138);
nor U6424 (N_6424,N_5780,N_5875);
or U6425 (N_6425,N_6319,N_5685);
nor U6426 (N_6426,N_5865,N_6113);
nor U6427 (N_6427,N_5752,N_6003);
nor U6428 (N_6428,N_6130,N_5809);
nand U6429 (N_6429,N_6158,N_5758);
or U6430 (N_6430,N_5697,N_6393);
nand U6431 (N_6431,N_6194,N_5880);
nand U6432 (N_6432,N_6102,N_5779);
and U6433 (N_6433,N_5608,N_6143);
and U6434 (N_6434,N_6311,N_5928);
nor U6435 (N_6435,N_5706,N_5632);
or U6436 (N_6436,N_5777,N_6112);
nand U6437 (N_6437,N_6168,N_5603);
nor U6438 (N_6438,N_5918,N_5848);
and U6439 (N_6439,N_6381,N_5907);
and U6440 (N_6440,N_5782,N_5607);
or U6441 (N_6441,N_5645,N_5901);
and U6442 (N_6442,N_6058,N_6046);
nor U6443 (N_6443,N_6302,N_6172);
nor U6444 (N_6444,N_6107,N_6159);
nor U6445 (N_6445,N_5951,N_5680);
nand U6446 (N_6446,N_6098,N_6214);
nand U6447 (N_6447,N_5696,N_5887);
nor U6448 (N_6448,N_6219,N_5924);
or U6449 (N_6449,N_6322,N_6139);
nor U6450 (N_6450,N_6074,N_6069);
or U6451 (N_6451,N_6129,N_5710);
nor U6452 (N_6452,N_6292,N_5817);
nor U6453 (N_6453,N_5713,N_6095);
or U6454 (N_6454,N_6227,N_6018);
nor U6455 (N_6455,N_6323,N_5755);
and U6456 (N_6456,N_6002,N_5998);
or U6457 (N_6457,N_5933,N_5738);
nand U6458 (N_6458,N_5778,N_5684);
nor U6459 (N_6459,N_5911,N_5611);
and U6460 (N_6460,N_6105,N_5830);
or U6461 (N_6461,N_5668,N_6368);
or U6462 (N_6462,N_6283,N_5703);
nand U6463 (N_6463,N_6220,N_6256);
nor U6464 (N_6464,N_5843,N_6305);
nor U6465 (N_6465,N_6359,N_5702);
nor U6466 (N_6466,N_5683,N_6073);
nand U6467 (N_6467,N_5869,N_5804);
and U6468 (N_6468,N_6300,N_5826);
nor U6469 (N_6469,N_6109,N_5797);
and U6470 (N_6470,N_6171,N_6071);
or U6471 (N_6471,N_6308,N_5635);
and U6472 (N_6472,N_6057,N_5655);
and U6473 (N_6473,N_6086,N_6282);
and U6474 (N_6474,N_6090,N_6328);
or U6475 (N_6475,N_6280,N_5638);
nand U6476 (N_6476,N_5935,N_6068);
or U6477 (N_6477,N_5651,N_6181);
nand U6478 (N_6478,N_5980,N_5665);
and U6479 (N_6479,N_6096,N_6396);
nand U6480 (N_6480,N_5629,N_6244);
and U6481 (N_6481,N_5970,N_5949);
nor U6482 (N_6482,N_5682,N_6080);
or U6483 (N_6483,N_5663,N_5993);
nor U6484 (N_6484,N_6075,N_5825);
nand U6485 (N_6485,N_6378,N_6287);
nand U6486 (N_6486,N_6379,N_5771);
nor U6487 (N_6487,N_5737,N_5605);
nor U6488 (N_6488,N_6193,N_5895);
nor U6489 (N_6489,N_5909,N_6123);
nand U6490 (N_6490,N_5727,N_6110);
nand U6491 (N_6491,N_6173,N_5751);
and U6492 (N_6492,N_6091,N_5805);
nor U6493 (N_6493,N_5630,N_5876);
and U6494 (N_6494,N_5904,N_6094);
xor U6495 (N_6495,N_5765,N_5705);
nor U6496 (N_6496,N_5905,N_5798);
and U6497 (N_6497,N_6276,N_5840);
or U6498 (N_6498,N_5678,N_6072);
or U6499 (N_6499,N_5821,N_5967);
nand U6500 (N_6500,N_5926,N_6019);
nor U6501 (N_6501,N_6081,N_6257);
nor U6502 (N_6502,N_6325,N_6082);
or U6503 (N_6503,N_6087,N_5983);
nand U6504 (N_6504,N_5745,N_5836);
and U6505 (N_6505,N_6229,N_6358);
nor U6506 (N_6506,N_6165,N_6254);
or U6507 (N_6507,N_6156,N_6197);
nor U6508 (N_6508,N_6232,N_6395);
and U6509 (N_6509,N_6179,N_6119);
or U6510 (N_6510,N_5740,N_6314);
and U6511 (N_6511,N_5671,N_6392);
nand U6512 (N_6512,N_5768,N_5723);
nand U6513 (N_6513,N_5832,N_5772);
or U6514 (N_6514,N_6348,N_5812);
nand U6515 (N_6515,N_5900,N_6364);
nand U6516 (N_6516,N_6127,N_5718);
nor U6517 (N_6517,N_5894,N_5927);
and U6518 (N_6518,N_5649,N_6182);
xnor U6519 (N_6519,N_6385,N_6012);
nor U6520 (N_6520,N_5857,N_5898);
nand U6521 (N_6521,N_6230,N_5652);
nand U6522 (N_6522,N_5921,N_6178);
nor U6523 (N_6523,N_5664,N_5971);
and U6524 (N_6524,N_5747,N_5859);
nor U6525 (N_6525,N_5714,N_6166);
or U6526 (N_6526,N_5717,N_6192);
nor U6527 (N_6527,N_6088,N_6242);
nor U6528 (N_6528,N_6144,N_6128);
and U6529 (N_6529,N_6341,N_5882);
nor U6530 (N_6530,N_5853,N_6035);
nand U6531 (N_6531,N_6013,N_5988);
and U6532 (N_6532,N_6340,N_6032);
nor U6533 (N_6533,N_5606,N_5627);
nor U6534 (N_6534,N_5667,N_6051);
nor U6535 (N_6535,N_6376,N_6268);
and U6536 (N_6536,N_6063,N_6010);
nor U6537 (N_6537,N_6021,N_6020);
nor U6538 (N_6538,N_6238,N_5726);
and U6539 (N_6539,N_5672,N_5863);
or U6540 (N_6540,N_6334,N_6045);
nor U6541 (N_6541,N_6140,N_5829);
nor U6542 (N_6542,N_5987,N_5837);
nand U6543 (N_6543,N_5756,N_6085);
or U6544 (N_6544,N_6089,N_5938);
nand U6545 (N_6545,N_6034,N_5619);
nand U6546 (N_6546,N_5846,N_6059);
and U6547 (N_6547,N_6083,N_6246);
nand U6548 (N_6548,N_6356,N_5614);
nor U6549 (N_6549,N_5610,N_5801);
nand U6550 (N_6550,N_6186,N_5620);
and U6551 (N_6551,N_6187,N_5989);
or U6552 (N_6552,N_5815,N_5658);
nand U6553 (N_6553,N_6295,N_6125);
and U6554 (N_6554,N_5975,N_6296);
or U6555 (N_6555,N_6028,N_6147);
and U6556 (N_6556,N_5650,N_5800);
or U6557 (N_6557,N_5981,N_5890);
nand U6558 (N_6558,N_5735,N_5974);
and U6559 (N_6559,N_6155,N_5913);
and U6560 (N_6560,N_5639,N_5704);
or U6561 (N_6561,N_6272,N_6136);
and U6562 (N_6562,N_6064,N_6346);
nand U6563 (N_6563,N_6249,N_5749);
nor U6564 (N_6564,N_6053,N_6241);
and U6565 (N_6565,N_6329,N_5953);
or U6566 (N_6566,N_6289,N_6367);
or U6567 (N_6567,N_5733,N_5708);
and U6568 (N_6568,N_6317,N_5858);
nor U6569 (N_6569,N_6204,N_5783);
or U6570 (N_6570,N_6237,N_6160);
nand U6571 (N_6571,N_5719,N_5695);
and U6572 (N_6572,N_5786,N_6039);
nand U6573 (N_6573,N_5637,N_6264);
nand U6574 (N_6574,N_6366,N_5600);
or U6575 (N_6575,N_6200,N_5643);
nand U6576 (N_6576,N_5899,N_5613);
nor U6577 (N_6577,N_5986,N_6399);
or U6578 (N_6578,N_6279,N_6335);
nor U6579 (N_6579,N_6363,N_6371);
nand U6580 (N_6580,N_5795,N_6351);
or U6581 (N_6581,N_5767,N_5792);
and U6582 (N_6582,N_5742,N_5660);
and U6583 (N_6583,N_6217,N_6216);
and U6584 (N_6584,N_5892,N_6233);
nand U6585 (N_6585,N_6189,N_6121);
nand U6586 (N_6586,N_6061,N_5764);
nand U6587 (N_6587,N_5636,N_6060);
nand U6588 (N_6588,N_5769,N_5688);
or U6589 (N_6589,N_6387,N_5947);
or U6590 (N_6590,N_5960,N_5622);
nor U6591 (N_6591,N_5676,N_6225);
nor U6592 (N_6592,N_5822,N_6122);
or U6593 (N_6593,N_5902,N_5766);
nor U6594 (N_6594,N_6261,N_6037);
nand U6595 (N_6595,N_5621,N_5838);
and U6596 (N_6596,N_5939,N_5834);
nand U6597 (N_6597,N_6142,N_5647);
or U6598 (N_6598,N_5709,N_6209);
nand U6599 (N_6599,N_5673,N_5806);
nor U6600 (N_6600,N_5716,N_6153);
and U6601 (N_6601,N_5872,N_6150);
or U6602 (N_6602,N_6116,N_5849);
or U6603 (N_6603,N_6115,N_6223);
nand U6604 (N_6604,N_6391,N_5634);
nand U6605 (N_6605,N_5877,N_6077);
or U6606 (N_6606,N_5624,N_5725);
nor U6607 (N_6607,N_5976,N_5852);
or U6608 (N_6608,N_6043,N_5868);
or U6609 (N_6609,N_6008,N_6011);
nor U6610 (N_6610,N_5850,N_6065);
and U6611 (N_6611,N_5881,N_6006);
nand U6612 (N_6612,N_6333,N_6036);
nand U6613 (N_6613,N_6126,N_6176);
nand U6614 (N_6614,N_5956,N_5674);
nand U6615 (N_6615,N_6318,N_6342);
and U6616 (N_6616,N_6327,N_6285);
nand U6617 (N_6617,N_6245,N_5879);
nand U6618 (N_6618,N_5612,N_6164);
nand U6619 (N_6619,N_5724,N_6101);
nor U6620 (N_6620,N_5864,N_6022);
nor U6621 (N_6621,N_6211,N_5785);
nand U6622 (N_6622,N_6286,N_6208);
nor U6623 (N_6623,N_5626,N_5739);
or U6624 (N_6624,N_6345,N_5761);
nand U6625 (N_6625,N_5677,N_5811);
and U6626 (N_6626,N_5885,N_5760);
or U6627 (N_6627,N_6100,N_6271);
nand U6628 (N_6628,N_6330,N_6062);
nand U6629 (N_6629,N_5966,N_6222);
nand U6630 (N_6630,N_6236,N_6267);
and U6631 (N_6631,N_5720,N_5996);
nor U6632 (N_6632,N_5730,N_6084);
and U6633 (N_6633,N_6038,N_6290);
or U6634 (N_6634,N_6203,N_6324);
nand U6635 (N_6635,N_6108,N_5687);
and U6636 (N_6636,N_5914,N_6076);
and U6637 (N_6637,N_6394,N_5721);
or U6638 (N_6638,N_6029,N_6066);
or U6639 (N_6639,N_5734,N_6078);
nor U6640 (N_6640,N_5625,N_5823);
nand U6641 (N_6641,N_6093,N_5916);
nand U6642 (N_6642,N_5922,N_5753);
nand U6643 (N_6643,N_6120,N_5897);
and U6644 (N_6644,N_5839,N_5920);
and U6645 (N_6645,N_5991,N_5912);
and U6646 (N_6646,N_5936,N_6210);
nand U6647 (N_6647,N_6055,N_5616);
nand U6648 (N_6648,N_5642,N_6117);
nand U6649 (N_6649,N_5741,N_6339);
and U6650 (N_6650,N_6054,N_5754);
and U6651 (N_6651,N_5893,N_6134);
or U6652 (N_6652,N_5906,N_5762);
or U6653 (N_6653,N_6265,N_6005);
nor U6654 (N_6654,N_6332,N_5886);
and U6655 (N_6655,N_5690,N_5648);
or U6656 (N_6656,N_6111,N_5814);
nand U6657 (N_6657,N_5867,N_5824);
and U6658 (N_6658,N_6248,N_6042);
nand U6659 (N_6659,N_6023,N_6201);
and U6660 (N_6660,N_6048,N_5854);
nor U6661 (N_6661,N_5803,N_5955);
nor U6662 (N_6662,N_6354,N_5973);
and U6663 (N_6663,N_6007,N_5962);
nor U6664 (N_6664,N_5787,N_6070);
or U6665 (N_6665,N_5700,N_6106);
nand U6666 (N_6666,N_6025,N_6009);
or U6667 (N_6667,N_5776,N_5618);
nand U6668 (N_6668,N_6269,N_6024);
nor U6669 (N_6669,N_5657,N_5957);
nor U6670 (N_6670,N_5954,N_6154);
nor U6671 (N_6671,N_6380,N_6137);
and U6672 (N_6672,N_6360,N_6162);
nand U6673 (N_6673,N_6228,N_6031);
or U6674 (N_6674,N_6337,N_6250);
nor U6675 (N_6675,N_5888,N_6163);
nor U6676 (N_6676,N_5969,N_5644);
nand U6677 (N_6677,N_6049,N_6321);
or U6678 (N_6678,N_5847,N_6369);
nand U6679 (N_6679,N_6350,N_6353);
or U6680 (N_6680,N_6313,N_5944);
nor U6681 (N_6681,N_6374,N_6251);
nor U6682 (N_6682,N_5965,N_6259);
and U6683 (N_6683,N_5978,N_5711);
nand U6684 (N_6684,N_6050,N_6326);
nor U6685 (N_6685,N_5609,N_6177);
nor U6686 (N_6686,N_6310,N_6375);
and U6687 (N_6687,N_6170,N_6016);
nand U6688 (N_6688,N_5679,N_5628);
and U6689 (N_6689,N_5763,N_6263);
and U6690 (N_6690,N_5732,N_5977);
nand U6691 (N_6691,N_6382,N_6239);
or U6692 (N_6692,N_5744,N_6301);
or U6693 (N_6693,N_5844,N_6355);
and U6694 (N_6694,N_6352,N_6299);
or U6695 (N_6695,N_5666,N_5810);
nor U6696 (N_6696,N_6386,N_6243);
or U6697 (N_6697,N_6370,N_6114);
nor U6698 (N_6698,N_6252,N_5759);
nor U6699 (N_6699,N_6331,N_6133);
or U6700 (N_6700,N_6213,N_5770);
and U6701 (N_6701,N_6149,N_6198);
nor U6702 (N_6702,N_5884,N_6255);
nor U6703 (N_6703,N_5950,N_5931);
nor U6704 (N_6704,N_5984,N_6388);
or U6705 (N_6705,N_5932,N_6309);
nand U6706 (N_6706,N_5923,N_5985);
nor U6707 (N_6707,N_5669,N_5845);
or U6708 (N_6708,N_5990,N_6253);
or U6709 (N_6709,N_5750,N_5878);
or U6710 (N_6710,N_5903,N_5889);
and U6711 (N_6711,N_6067,N_5860);
nor U6712 (N_6712,N_6384,N_6215);
nor U6713 (N_6713,N_6026,N_6044);
nand U6714 (N_6714,N_5729,N_6104);
nor U6715 (N_6715,N_5694,N_6212);
and U6716 (N_6716,N_5699,N_6131);
nor U6717 (N_6717,N_6015,N_6235);
or U6718 (N_6718,N_6027,N_6247);
and U6719 (N_6719,N_5775,N_5623);
or U6720 (N_6720,N_5948,N_5942);
nand U6721 (N_6721,N_5796,N_5940);
or U6722 (N_6722,N_6336,N_6266);
nor U6723 (N_6723,N_5871,N_5617);
nor U6724 (N_6724,N_5722,N_5789);
or U6725 (N_6725,N_6196,N_5982);
nor U6726 (N_6726,N_5925,N_5662);
nand U6727 (N_6727,N_5819,N_5693);
or U6728 (N_6728,N_6297,N_6001);
nand U6729 (N_6729,N_6260,N_5781);
nor U6730 (N_6730,N_6383,N_6017);
nand U6731 (N_6731,N_5728,N_6306);
and U6732 (N_6732,N_5972,N_5841);
or U6733 (N_6733,N_6146,N_6185);
and U6734 (N_6734,N_5917,N_5896);
nand U6735 (N_6735,N_6207,N_6097);
or U6736 (N_6736,N_6056,N_6298);
nand U6737 (N_6737,N_5633,N_6398);
nor U6738 (N_6738,N_5686,N_6307);
nor U6739 (N_6739,N_5794,N_5615);
nand U6740 (N_6740,N_6052,N_5748);
or U6741 (N_6741,N_6099,N_5968);
nor U6742 (N_6742,N_5640,N_6191);
or U6743 (N_6743,N_6205,N_6347);
nand U6744 (N_6744,N_5802,N_5773);
and U6745 (N_6745,N_5602,N_5958);
nor U6746 (N_6746,N_6161,N_5698);
nand U6747 (N_6747,N_6258,N_5943);
and U6748 (N_6748,N_5692,N_6124);
or U6749 (N_6749,N_5631,N_5675);
or U6750 (N_6750,N_5604,N_6357);
nor U6751 (N_6751,N_5995,N_6278);
or U6752 (N_6752,N_5856,N_5964);
nand U6753 (N_6753,N_5908,N_6277);
and U6754 (N_6754,N_6188,N_5712);
nor U6755 (N_6755,N_6174,N_5784);
or U6756 (N_6756,N_5659,N_6169);
nor U6757 (N_6757,N_6270,N_5937);
nand U6758 (N_6758,N_5736,N_6132);
and U6759 (N_6759,N_5670,N_5870);
or U6760 (N_6760,N_6349,N_6397);
nand U6761 (N_6761,N_5855,N_6221);
or U6762 (N_6762,N_5994,N_6362);
nand U6763 (N_6763,N_5788,N_5707);
nor U6764 (N_6764,N_6315,N_5654);
nand U6765 (N_6765,N_6281,N_5891);
nor U6766 (N_6766,N_6304,N_6000);
or U6767 (N_6767,N_6183,N_6004);
nand U6768 (N_6768,N_5820,N_6145);
nand U6769 (N_6769,N_6294,N_5746);
or U6770 (N_6770,N_6202,N_6338);
and U6771 (N_6771,N_5929,N_5791);
and U6772 (N_6772,N_6041,N_6288);
nor U6773 (N_6773,N_5851,N_6218);
nor U6774 (N_6774,N_6240,N_6373);
nand U6775 (N_6775,N_5946,N_5873);
nor U6776 (N_6776,N_5831,N_5930);
and U6777 (N_6777,N_6231,N_5883);
and U6778 (N_6778,N_6284,N_5807);
and U6779 (N_6779,N_6372,N_5866);
xnor U6780 (N_6780,N_6274,N_6184);
and U6781 (N_6781,N_6344,N_5774);
and U6782 (N_6782,N_5743,N_6361);
or U6783 (N_6783,N_5757,N_6316);
and U6784 (N_6784,N_6320,N_5833);
nor U6785 (N_6785,N_6377,N_5835);
or U6786 (N_6786,N_5828,N_5701);
and U6787 (N_6787,N_5997,N_6040);
and U6788 (N_6788,N_6151,N_5661);
nor U6789 (N_6789,N_6175,N_6190);
or U6790 (N_6790,N_6157,N_6273);
nor U6791 (N_6791,N_6135,N_6275);
nor U6792 (N_6792,N_5818,N_6224);
nor U6793 (N_6793,N_6291,N_6195);
or U6794 (N_6794,N_5816,N_5862);
or U6795 (N_6795,N_5999,N_6206);
nor U6796 (N_6796,N_5919,N_5963);
or U6797 (N_6797,N_5959,N_6226);
nor U6798 (N_6798,N_6180,N_6033);
or U6799 (N_6799,N_6293,N_5941);
or U6800 (N_6800,N_6187,N_5902);
xnor U6801 (N_6801,N_5742,N_6186);
or U6802 (N_6802,N_6230,N_5806);
nor U6803 (N_6803,N_5619,N_5940);
or U6804 (N_6804,N_5715,N_5714);
or U6805 (N_6805,N_6192,N_6271);
and U6806 (N_6806,N_5907,N_5630);
or U6807 (N_6807,N_5956,N_6199);
nand U6808 (N_6808,N_5690,N_6134);
nand U6809 (N_6809,N_5613,N_6109);
or U6810 (N_6810,N_5873,N_6323);
or U6811 (N_6811,N_6306,N_6277);
nand U6812 (N_6812,N_6220,N_5924);
nand U6813 (N_6813,N_6324,N_5957);
nor U6814 (N_6814,N_6027,N_5688);
or U6815 (N_6815,N_5952,N_6272);
and U6816 (N_6816,N_6327,N_6180);
nand U6817 (N_6817,N_5972,N_5703);
nand U6818 (N_6818,N_6075,N_6353);
nand U6819 (N_6819,N_5600,N_5941);
or U6820 (N_6820,N_6270,N_5917);
and U6821 (N_6821,N_6005,N_6124);
or U6822 (N_6822,N_6070,N_6136);
nor U6823 (N_6823,N_6172,N_5749);
or U6824 (N_6824,N_5781,N_5666);
or U6825 (N_6825,N_5776,N_5775);
or U6826 (N_6826,N_5976,N_6050);
and U6827 (N_6827,N_5974,N_5787);
nor U6828 (N_6828,N_6342,N_5863);
nor U6829 (N_6829,N_5749,N_5793);
nand U6830 (N_6830,N_5973,N_5897);
and U6831 (N_6831,N_5734,N_5999);
nand U6832 (N_6832,N_5805,N_5726);
nor U6833 (N_6833,N_5747,N_6349);
nor U6834 (N_6834,N_5667,N_6049);
and U6835 (N_6835,N_5747,N_5898);
nand U6836 (N_6836,N_5792,N_5657);
or U6837 (N_6837,N_6007,N_5722);
or U6838 (N_6838,N_5892,N_6186);
nor U6839 (N_6839,N_5976,N_6377);
nor U6840 (N_6840,N_6282,N_6376);
and U6841 (N_6841,N_5812,N_5793);
or U6842 (N_6842,N_6023,N_6043);
or U6843 (N_6843,N_5989,N_5893);
and U6844 (N_6844,N_5991,N_5973);
or U6845 (N_6845,N_5743,N_6314);
and U6846 (N_6846,N_6102,N_6288);
nand U6847 (N_6847,N_6124,N_5640);
and U6848 (N_6848,N_5757,N_5832);
or U6849 (N_6849,N_5897,N_6080);
nand U6850 (N_6850,N_5795,N_6238);
nand U6851 (N_6851,N_6360,N_5695);
or U6852 (N_6852,N_6264,N_5941);
and U6853 (N_6853,N_5618,N_6135);
and U6854 (N_6854,N_5656,N_5731);
nand U6855 (N_6855,N_5830,N_5963);
and U6856 (N_6856,N_5681,N_6121);
or U6857 (N_6857,N_5934,N_5988);
and U6858 (N_6858,N_5733,N_6106);
or U6859 (N_6859,N_5882,N_5602);
or U6860 (N_6860,N_5722,N_6086);
and U6861 (N_6861,N_5904,N_5966);
nand U6862 (N_6862,N_5711,N_5768);
or U6863 (N_6863,N_5922,N_6007);
nand U6864 (N_6864,N_6273,N_5903);
nor U6865 (N_6865,N_6320,N_5603);
and U6866 (N_6866,N_6349,N_5609);
nand U6867 (N_6867,N_6330,N_6355);
and U6868 (N_6868,N_5748,N_6071);
or U6869 (N_6869,N_6002,N_5795);
nand U6870 (N_6870,N_5901,N_6120);
nor U6871 (N_6871,N_6191,N_6141);
and U6872 (N_6872,N_6084,N_5611);
nand U6873 (N_6873,N_6072,N_6160);
nor U6874 (N_6874,N_5773,N_6267);
nor U6875 (N_6875,N_6232,N_5679);
nor U6876 (N_6876,N_6290,N_5662);
nor U6877 (N_6877,N_5890,N_5745);
nor U6878 (N_6878,N_5948,N_6348);
and U6879 (N_6879,N_5797,N_5687);
and U6880 (N_6880,N_5747,N_6254);
nor U6881 (N_6881,N_5900,N_5894);
nand U6882 (N_6882,N_5749,N_5708);
nor U6883 (N_6883,N_6292,N_6041);
or U6884 (N_6884,N_6032,N_6218);
and U6885 (N_6885,N_5842,N_6390);
nor U6886 (N_6886,N_6199,N_5613);
and U6887 (N_6887,N_5877,N_5604);
nor U6888 (N_6888,N_5814,N_6122);
or U6889 (N_6889,N_5963,N_5862);
or U6890 (N_6890,N_5958,N_5953);
or U6891 (N_6891,N_5878,N_6137);
and U6892 (N_6892,N_6358,N_6257);
or U6893 (N_6893,N_5842,N_5626);
and U6894 (N_6894,N_6009,N_6152);
nor U6895 (N_6895,N_6304,N_5994);
nor U6896 (N_6896,N_6333,N_5650);
nor U6897 (N_6897,N_5916,N_5605);
and U6898 (N_6898,N_6221,N_6174);
nor U6899 (N_6899,N_5695,N_5697);
and U6900 (N_6900,N_5726,N_5815);
nor U6901 (N_6901,N_5876,N_5702);
nand U6902 (N_6902,N_5609,N_5884);
nor U6903 (N_6903,N_6178,N_6268);
xor U6904 (N_6904,N_6160,N_5891);
or U6905 (N_6905,N_6033,N_6368);
or U6906 (N_6906,N_5988,N_6299);
nor U6907 (N_6907,N_6236,N_6022);
or U6908 (N_6908,N_5998,N_6241);
and U6909 (N_6909,N_5721,N_5897);
and U6910 (N_6910,N_5814,N_5629);
nand U6911 (N_6911,N_5807,N_5912);
and U6912 (N_6912,N_5915,N_6294);
or U6913 (N_6913,N_6278,N_6047);
and U6914 (N_6914,N_6316,N_5646);
nor U6915 (N_6915,N_5735,N_5896);
or U6916 (N_6916,N_5993,N_5911);
and U6917 (N_6917,N_5609,N_6052);
nand U6918 (N_6918,N_5641,N_6234);
or U6919 (N_6919,N_5853,N_6389);
or U6920 (N_6920,N_6276,N_6023);
or U6921 (N_6921,N_5714,N_6058);
nand U6922 (N_6922,N_6195,N_6036);
or U6923 (N_6923,N_5946,N_5602);
nor U6924 (N_6924,N_5820,N_6386);
and U6925 (N_6925,N_6364,N_5910);
and U6926 (N_6926,N_5836,N_6365);
or U6927 (N_6927,N_6386,N_5656);
or U6928 (N_6928,N_5899,N_5730);
nand U6929 (N_6929,N_5628,N_5909);
nor U6930 (N_6930,N_6160,N_6228);
nor U6931 (N_6931,N_5752,N_5831);
and U6932 (N_6932,N_6085,N_6286);
nor U6933 (N_6933,N_5880,N_6319);
nor U6934 (N_6934,N_6256,N_6252);
or U6935 (N_6935,N_5785,N_5741);
and U6936 (N_6936,N_5881,N_5979);
or U6937 (N_6937,N_5837,N_5963);
nor U6938 (N_6938,N_6222,N_5760);
and U6939 (N_6939,N_6248,N_5872);
nor U6940 (N_6940,N_5827,N_5793);
and U6941 (N_6941,N_5799,N_5755);
nand U6942 (N_6942,N_5752,N_6219);
or U6943 (N_6943,N_5874,N_5876);
and U6944 (N_6944,N_6029,N_5991);
nand U6945 (N_6945,N_6379,N_5997);
and U6946 (N_6946,N_6053,N_5647);
nand U6947 (N_6947,N_6040,N_5709);
and U6948 (N_6948,N_5828,N_5807);
and U6949 (N_6949,N_5903,N_6116);
nor U6950 (N_6950,N_5979,N_6078);
or U6951 (N_6951,N_6010,N_5600);
nand U6952 (N_6952,N_5984,N_6378);
or U6953 (N_6953,N_5695,N_5847);
and U6954 (N_6954,N_5608,N_5643);
or U6955 (N_6955,N_5736,N_5611);
nor U6956 (N_6956,N_5834,N_6101);
nand U6957 (N_6957,N_6392,N_6106);
and U6958 (N_6958,N_6248,N_6118);
nand U6959 (N_6959,N_6150,N_5686);
nand U6960 (N_6960,N_5690,N_5707);
and U6961 (N_6961,N_6098,N_6117);
or U6962 (N_6962,N_6020,N_6231);
or U6963 (N_6963,N_5983,N_5621);
or U6964 (N_6964,N_6126,N_6003);
nor U6965 (N_6965,N_6199,N_5801);
or U6966 (N_6966,N_6209,N_5997);
nand U6967 (N_6967,N_5669,N_5969);
and U6968 (N_6968,N_6153,N_6275);
nand U6969 (N_6969,N_6350,N_5867);
nor U6970 (N_6970,N_5784,N_6234);
and U6971 (N_6971,N_5728,N_5996);
nand U6972 (N_6972,N_5687,N_6245);
or U6973 (N_6973,N_5660,N_5639);
and U6974 (N_6974,N_5834,N_6061);
and U6975 (N_6975,N_6282,N_5877);
and U6976 (N_6976,N_6107,N_6186);
nor U6977 (N_6977,N_6144,N_5783);
nor U6978 (N_6978,N_6374,N_5661);
and U6979 (N_6979,N_6085,N_6244);
nor U6980 (N_6980,N_6395,N_5624);
nor U6981 (N_6981,N_6380,N_6314);
nand U6982 (N_6982,N_6160,N_5983);
or U6983 (N_6983,N_6162,N_6359);
or U6984 (N_6984,N_6161,N_6389);
and U6985 (N_6985,N_5847,N_6261);
nor U6986 (N_6986,N_5902,N_6369);
nand U6987 (N_6987,N_5703,N_6346);
or U6988 (N_6988,N_6170,N_6110);
and U6989 (N_6989,N_5848,N_5624);
nand U6990 (N_6990,N_6289,N_6137);
nor U6991 (N_6991,N_6133,N_5774);
xor U6992 (N_6992,N_6241,N_6394);
or U6993 (N_6993,N_6115,N_5827);
or U6994 (N_6994,N_5660,N_5695);
or U6995 (N_6995,N_6118,N_6391);
nor U6996 (N_6996,N_5705,N_5913);
nand U6997 (N_6997,N_5718,N_6300);
or U6998 (N_6998,N_6183,N_5998);
and U6999 (N_6999,N_6300,N_6064);
nor U7000 (N_7000,N_6331,N_6064);
or U7001 (N_7001,N_6024,N_5940);
nand U7002 (N_7002,N_6114,N_6056);
nor U7003 (N_7003,N_6362,N_5613);
nand U7004 (N_7004,N_5688,N_5818);
nor U7005 (N_7005,N_6367,N_6172);
nand U7006 (N_7006,N_5919,N_6370);
or U7007 (N_7007,N_5731,N_6158);
or U7008 (N_7008,N_6303,N_6034);
and U7009 (N_7009,N_6021,N_5813);
and U7010 (N_7010,N_6367,N_5681);
nand U7011 (N_7011,N_5999,N_6197);
nand U7012 (N_7012,N_5736,N_6388);
nor U7013 (N_7013,N_6124,N_5913);
or U7014 (N_7014,N_6331,N_5940);
and U7015 (N_7015,N_5844,N_6000);
or U7016 (N_7016,N_5885,N_6371);
nor U7017 (N_7017,N_5890,N_5750);
or U7018 (N_7018,N_5788,N_6371);
or U7019 (N_7019,N_5795,N_6396);
or U7020 (N_7020,N_5913,N_5877);
or U7021 (N_7021,N_5751,N_5836);
and U7022 (N_7022,N_6139,N_6275);
and U7023 (N_7023,N_6245,N_5650);
nand U7024 (N_7024,N_5805,N_5618);
nand U7025 (N_7025,N_6396,N_6127);
nand U7026 (N_7026,N_5709,N_6000);
or U7027 (N_7027,N_6124,N_6266);
nor U7028 (N_7028,N_6034,N_5621);
nor U7029 (N_7029,N_6281,N_5648);
and U7030 (N_7030,N_5950,N_5969);
or U7031 (N_7031,N_6380,N_6100);
nand U7032 (N_7032,N_6294,N_6240);
nand U7033 (N_7033,N_6121,N_5756);
nand U7034 (N_7034,N_5912,N_6362);
or U7035 (N_7035,N_5683,N_6160);
and U7036 (N_7036,N_5841,N_5617);
or U7037 (N_7037,N_5725,N_5976);
xnor U7038 (N_7038,N_6336,N_5857);
nor U7039 (N_7039,N_5728,N_5859);
nand U7040 (N_7040,N_6220,N_6015);
nand U7041 (N_7041,N_6067,N_5995);
and U7042 (N_7042,N_6164,N_5638);
nand U7043 (N_7043,N_5946,N_6315);
and U7044 (N_7044,N_5821,N_5891);
nand U7045 (N_7045,N_6229,N_5973);
and U7046 (N_7046,N_6070,N_6033);
or U7047 (N_7047,N_5804,N_6297);
and U7048 (N_7048,N_5830,N_5819);
nor U7049 (N_7049,N_5840,N_5922);
or U7050 (N_7050,N_5890,N_5930);
and U7051 (N_7051,N_6064,N_5800);
or U7052 (N_7052,N_6366,N_6381);
nor U7053 (N_7053,N_6159,N_6095);
or U7054 (N_7054,N_5783,N_5748);
nor U7055 (N_7055,N_5965,N_6320);
and U7056 (N_7056,N_6269,N_6382);
nor U7057 (N_7057,N_5876,N_6195);
or U7058 (N_7058,N_5649,N_5936);
nor U7059 (N_7059,N_6134,N_6200);
nand U7060 (N_7060,N_5918,N_5705);
or U7061 (N_7061,N_5772,N_6069);
or U7062 (N_7062,N_6124,N_5944);
or U7063 (N_7063,N_5925,N_6226);
and U7064 (N_7064,N_6078,N_6277);
nand U7065 (N_7065,N_6114,N_6238);
or U7066 (N_7066,N_6286,N_6331);
nand U7067 (N_7067,N_6237,N_5662);
or U7068 (N_7068,N_5737,N_5619);
or U7069 (N_7069,N_6363,N_6310);
nand U7070 (N_7070,N_5846,N_6237);
nor U7071 (N_7071,N_6299,N_5610);
nand U7072 (N_7072,N_6315,N_6327);
nor U7073 (N_7073,N_6359,N_6349);
or U7074 (N_7074,N_6178,N_6194);
or U7075 (N_7075,N_6020,N_6027);
and U7076 (N_7076,N_6040,N_6146);
and U7077 (N_7077,N_6046,N_6000);
nor U7078 (N_7078,N_5808,N_6301);
nand U7079 (N_7079,N_6328,N_6302);
or U7080 (N_7080,N_6174,N_5635);
and U7081 (N_7081,N_5914,N_6067);
or U7082 (N_7082,N_5854,N_6196);
or U7083 (N_7083,N_5791,N_6006);
or U7084 (N_7084,N_5857,N_6041);
or U7085 (N_7085,N_5743,N_6007);
nand U7086 (N_7086,N_5719,N_5642);
xnor U7087 (N_7087,N_5761,N_5759);
nand U7088 (N_7088,N_6097,N_5653);
nor U7089 (N_7089,N_5664,N_5717);
nor U7090 (N_7090,N_5680,N_5790);
or U7091 (N_7091,N_5727,N_5869);
and U7092 (N_7092,N_6063,N_5701);
or U7093 (N_7093,N_6186,N_6010);
nor U7094 (N_7094,N_6179,N_6291);
and U7095 (N_7095,N_5858,N_5751);
nor U7096 (N_7096,N_5922,N_6339);
or U7097 (N_7097,N_6190,N_5908);
xnor U7098 (N_7098,N_6098,N_5995);
nor U7099 (N_7099,N_5913,N_5675);
nor U7100 (N_7100,N_6127,N_5822);
nand U7101 (N_7101,N_5833,N_5847);
and U7102 (N_7102,N_6209,N_5791);
nand U7103 (N_7103,N_6286,N_5787);
nand U7104 (N_7104,N_5876,N_6335);
nand U7105 (N_7105,N_6156,N_6257);
or U7106 (N_7106,N_6243,N_5852);
nor U7107 (N_7107,N_6102,N_5882);
or U7108 (N_7108,N_5766,N_6192);
or U7109 (N_7109,N_6394,N_6148);
nand U7110 (N_7110,N_6039,N_6088);
and U7111 (N_7111,N_6289,N_5804);
or U7112 (N_7112,N_6172,N_5964);
nor U7113 (N_7113,N_6339,N_5803);
nor U7114 (N_7114,N_5916,N_6257);
and U7115 (N_7115,N_5770,N_5660);
and U7116 (N_7116,N_5673,N_5823);
or U7117 (N_7117,N_5809,N_6020);
or U7118 (N_7118,N_5668,N_6096);
or U7119 (N_7119,N_6359,N_5914);
nor U7120 (N_7120,N_5845,N_5948);
nor U7121 (N_7121,N_6286,N_5965);
nand U7122 (N_7122,N_6312,N_6193);
or U7123 (N_7123,N_6280,N_6114);
nor U7124 (N_7124,N_6214,N_6194);
nand U7125 (N_7125,N_6312,N_5922);
nand U7126 (N_7126,N_5742,N_5712);
nor U7127 (N_7127,N_6206,N_6251);
or U7128 (N_7128,N_5976,N_5784);
or U7129 (N_7129,N_5681,N_5764);
or U7130 (N_7130,N_6162,N_6252);
nor U7131 (N_7131,N_6036,N_6060);
or U7132 (N_7132,N_5601,N_6006);
nor U7133 (N_7133,N_6180,N_5986);
nand U7134 (N_7134,N_6093,N_5798);
and U7135 (N_7135,N_6188,N_5982);
nor U7136 (N_7136,N_6008,N_5865);
nand U7137 (N_7137,N_6258,N_6158);
nand U7138 (N_7138,N_6226,N_5645);
nor U7139 (N_7139,N_5796,N_5786);
and U7140 (N_7140,N_6284,N_6392);
or U7141 (N_7141,N_5937,N_5796);
nor U7142 (N_7142,N_5965,N_6208);
and U7143 (N_7143,N_6294,N_6337);
and U7144 (N_7144,N_5659,N_6025);
nand U7145 (N_7145,N_5741,N_6387);
and U7146 (N_7146,N_5898,N_6284);
and U7147 (N_7147,N_5938,N_6394);
or U7148 (N_7148,N_5789,N_6097);
and U7149 (N_7149,N_5938,N_6158);
or U7150 (N_7150,N_5653,N_6070);
or U7151 (N_7151,N_6254,N_5858);
nand U7152 (N_7152,N_6375,N_5789);
nor U7153 (N_7153,N_5886,N_6078);
nand U7154 (N_7154,N_6352,N_5989);
or U7155 (N_7155,N_5943,N_6285);
nor U7156 (N_7156,N_6166,N_5809);
nor U7157 (N_7157,N_5709,N_6207);
nand U7158 (N_7158,N_6103,N_6162);
xnor U7159 (N_7159,N_6205,N_6114);
nand U7160 (N_7160,N_5744,N_5787);
nand U7161 (N_7161,N_5697,N_6028);
or U7162 (N_7162,N_6184,N_6323);
nor U7163 (N_7163,N_5634,N_5866);
nor U7164 (N_7164,N_5952,N_6321);
and U7165 (N_7165,N_6024,N_5713);
nand U7166 (N_7166,N_6320,N_6006);
nor U7167 (N_7167,N_5872,N_5755);
nand U7168 (N_7168,N_6181,N_6001);
or U7169 (N_7169,N_5635,N_6043);
and U7170 (N_7170,N_5715,N_6359);
nor U7171 (N_7171,N_5759,N_5988);
nand U7172 (N_7172,N_6234,N_6140);
or U7173 (N_7173,N_6219,N_6311);
nor U7174 (N_7174,N_5848,N_5925);
or U7175 (N_7175,N_5700,N_5699);
nand U7176 (N_7176,N_6218,N_6222);
nand U7177 (N_7177,N_5849,N_5713);
and U7178 (N_7178,N_5822,N_6059);
and U7179 (N_7179,N_5741,N_5639);
nor U7180 (N_7180,N_6390,N_5863);
nor U7181 (N_7181,N_5612,N_5814);
or U7182 (N_7182,N_6154,N_5618);
nand U7183 (N_7183,N_5742,N_6332);
nor U7184 (N_7184,N_6358,N_6116);
and U7185 (N_7185,N_6276,N_5716);
or U7186 (N_7186,N_5975,N_6374);
nand U7187 (N_7187,N_6192,N_6325);
nand U7188 (N_7188,N_6263,N_6349);
nor U7189 (N_7189,N_6299,N_6096);
or U7190 (N_7190,N_6129,N_5659);
xor U7191 (N_7191,N_5990,N_6297);
nand U7192 (N_7192,N_5628,N_5837);
and U7193 (N_7193,N_6387,N_5933);
or U7194 (N_7194,N_5779,N_6046);
or U7195 (N_7195,N_5725,N_6063);
or U7196 (N_7196,N_6212,N_6102);
or U7197 (N_7197,N_6303,N_5666);
or U7198 (N_7198,N_5694,N_6363);
nand U7199 (N_7199,N_5776,N_6071);
or U7200 (N_7200,N_6884,N_7161);
nor U7201 (N_7201,N_6628,N_6509);
nand U7202 (N_7202,N_6402,N_6842);
nor U7203 (N_7203,N_6439,N_6919);
nor U7204 (N_7204,N_7179,N_6976);
and U7205 (N_7205,N_6987,N_7131);
nor U7206 (N_7206,N_6409,N_7187);
and U7207 (N_7207,N_6971,N_6486);
or U7208 (N_7208,N_7098,N_6800);
nor U7209 (N_7209,N_6672,N_6744);
and U7210 (N_7210,N_7065,N_6621);
or U7211 (N_7211,N_6730,N_6946);
or U7212 (N_7212,N_6640,N_6878);
and U7213 (N_7213,N_6969,N_7117);
or U7214 (N_7214,N_6892,N_6851);
and U7215 (N_7215,N_7151,N_6605);
nor U7216 (N_7216,N_7101,N_6548);
xor U7217 (N_7217,N_7041,N_6822);
or U7218 (N_7218,N_6570,N_6556);
and U7219 (N_7219,N_6807,N_6644);
nor U7220 (N_7220,N_7149,N_6827);
nand U7221 (N_7221,N_7140,N_6420);
or U7222 (N_7222,N_6533,N_6604);
and U7223 (N_7223,N_6664,N_6510);
and U7224 (N_7224,N_7192,N_7076);
nor U7225 (N_7225,N_6841,N_6748);
nor U7226 (N_7226,N_7113,N_7163);
nor U7227 (N_7227,N_6889,N_6867);
nor U7228 (N_7228,N_6525,N_7199);
or U7229 (N_7229,N_6810,N_6787);
and U7230 (N_7230,N_6790,N_6865);
nand U7231 (N_7231,N_6562,N_6922);
or U7232 (N_7232,N_6653,N_6530);
nand U7233 (N_7233,N_6584,N_6534);
nor U7234 (N_7234,N_6482,N_6665);
or U7235 (N_7235,N_6953,N_7027);
nor U7236 (N_7236,N_6606,N_6581);
and U7237 (N_7237,N_6782,N_7123);
or U7238 (N_7238,N_6972,N_6825);
nor U7239 (N_7239,N_6542,N_6569);
nand U7240 (N_7240,N_6465,N_7004);
nor U7241 (N_7241,N_7046,N_6583);
nand U7242 (N_7242,N_6757,N_6982);
or U7243 (N_7243,N_6863,N_7068);
nor U7244 (N_7244,N_6591,N_6968);
or U7245 (N_7245,N_6661,N_6687);
and U7246 (N_7246,N_7168,N_6876);
or U7247 (N_7247,N_6668,N_6907);
nor U7248 (N_7248,N_6610,N_6903);
or U7249 (N_7249,N_6905,N_6738);
nor U7250 (N_7250,N_6513,N_7082);
nor U7251 (N_7251,N_7026,N_6688);
nor U7252 (N_7252,N_7162,N_6769);
and U7253 (N_7253,N_6400,N_7066);
nand U7254 (N_7254,N_6835,N_6958);
and U7255 (N_7255,N_7059,N_7094);
and U7256 (N_7256,N_6566,N_7050);
and U7257 (N_7257,N_6543,N_6720);
nor U7258 (N_7258,N_6762,N_7037);
or U7259 (N_7259,N_7114,N_6796);
nand U7260 (N_7260,N_6597,N_6499);
nand U7261 (N_7261,N_6537,N_6472);
nand U7262 (N_7262,N_6888,N_6558);
nand U7263 (N_7263,N_6430,N_6930);
nand U7264 (N_7264,N_7054,N_7132);
and U7265 (N_7265,N_6444,N_6812);
xor U7266 (N_7266,N_6742,N_6941);
nor U7267 (N_7267,N_6467,N_7074);
and U7268 (N_7268,N_6455,N_6788);
nor U7269 (N_7269,N_7127,N_6928);
xor U7270 (N_7270,N_7100,N_6718);
or U7271 (N_7271,N_6483,N_6421);
nand U7272 (N_7272,N_6641,N_6850);
or U7273 (N_7273,N_7104,N_7012);
nand U7274 (N_7274,N_6838,N_6829);
nand U7275 (N_7275,N_6526,N_6823);
and U7276 (N_7276,N_6567,N_6476);
nor U7277 (N_7277,N_6475,N_6849);
or U7278 (N_7278,N_6574,N_6778);
or U7279 (N_7279,N_6652,N_6600);
and U7280 (N_7280,N_7099,N_7049);
nand U7281 (N_7281,N_7048,N_6480);
or U7282 (N_7282,N_7045,N_6760);
and U7283 (N_7283,N_6714,N_6559);
nand U7284 (N_7284,N_7080,N_6425);
nor U7285 (N_7285,N_6708,N_6925);
or U7286 (N_7286,N_7152,N_7014);
nor U7287 (N_7287,N_6855,N_6939);
nor U7288 (N_7288,N_6754,N_7015);
nor U7289 (N_7289,N_6772,N_6684);
xnor U7290 (N_7290,N_7178,N_6471);
or U7291 (N_7291,N_6921,N_6458);
and U7292 (N_7292,N_7024,N_6485);
or U7293 (N_7293,N_6655,N_6761);
nor U7294 (N_7294,N_6989,N_7181);
nor U7295 (N_7295,N_7064,N_6636);
nand U7296 (N_7296,N_6834,N_6697);
xor U7297 (N_7297,N_6759,N_6632);
nand U7298 (N_7298,N_7003,N_6786);
or U7299 (N_7299,N_7125,N_6879);
or U7300 (N_7300,N_6477,N_6685);
and U7301 (N_7301,N_6413,N_6898);
nor U7302 (N_7302,N_7088,N_7121);
nand U7303 (N_7303,N_6705,N_6695);
nand U7304 (N_7304,N_6724,N_6920);
nand U7305 (N_7305,N_6831,N_6774);
nand U7306 (N_7306,N_7111,N_7171);
nand U7307 (N_7307,N_7154,N_6869);
nand U7308 (N_7308,N_6582,N_7182);
nor U7309 (N_7309,N_7159,N_6650);
nor U7310 (N_7310,N_7010,N_6433);
nor U7311 (N_7311,N_6657,N_6478);
and U7312 (N_7312,N_7002,N_6518);
or U7313 (N_7313,N_7028,N_7142);
nand U7314 (N_7314,N_6495,N_6915);
or U7315 (N_7315,N_6852,N_6484);
nand U7316 (N_7316,N_6722,N_6965);
nand U7317 (N_7317,N_7057,N_6906);
nand U7318 (N_7318,N_6881,N_6417);
nand U7319 (N_7319,N_7139,N_6734);
and U7320 (N_7320,N_6438,N_6511);
nor U7321 (N_7321,N_7023,N_7183);
nand U7322 (N_7322,N_6904,N_6616);
nor U7323 (N_7323,N_7155,N_6932);
or U7324 (N_7324,N_6929,N_6816);
and U7325 (N_7325,N_6549,N_6431);
or U7326 (N_7326,N_7020,N_6527);
or U7327 (N_7327,N_6998,N_6442);
nor U7328 (N_7328,N_6437,N_6590);
nand U7329 (N_7329,N_7085,N_6840);
and U7330 (N_7330,N_6412,N_6427);
and U7331 (N_7331,N_6912,N_6805);
and U7332 (N_7332,N_6733,N_7033);
nor U7333 (N_7333,N_6967,N_7089);
and U7334 (N_7334,N_7193,N_7119);
nand U7335 (N_7335,N_7150,N_6575);
or U7336 (N_7336,N_6634,N_6815);
nor U7337 (N_7337,N_6633,N_6502);
nor U7338 (N_7338,N_7128,N_6675);
nor U7339 (N_7339,N_7141,N_7035);
nor U7340 (N_7340,N_6962,N_6726);
or U7341 (N_7341,N_6847,N_6736);
or U7342 (N_7342,N_6448,N_6910);
or U7343 (N_7343,N_6899,N_6457);
nand U7344 (N_7344,N_6789,N_6961);
and U7345 (N_7345,N_7073,N_6897);
or U7346 (N_7346,N_6691,N_6490);
and U7347 (N_7347,N_6622,N_6456);
and U7348 (N_7348,N_6523,N_6909);
and U7349 (N_7349,N_6602,N_6704);
or U7350 (N_7350,N_7115,N_6565);
nor U7351 (N_7351,N_7186,N_7170);
and U7352 (N_7352,N_7146,N_6945);
and U7353 (N_7353,N_6515,N_6864);
nand U7354 (N_7354,N_6401,N_7034);
and U7355 (N_7355,N_6450,N_6498);
nand U7356 (N_7356,N_6445,N_7079);
nor U7357 (N_7357,N_6978,N_7043);
nand U7358 (N_7358,N_7039,N_7031);
or U7359 (N_7359,N_7135,N_6696);
nor U7360 (N_7360,N_6463,N_7018);
or U7361 (N_7361,N_7105,N_6700);
nor U7362 (N_7362,N_6435,N_6415);
and U7363 (N_7363,N_6447,N_6753);
or U7364 (N_7364,N_7157,N_6817);
nor U7365 (N_7365,N_6955,N_7148);
nand U7366 (N_7366,N_6853,N_6469);
and U7367 (N_7367,N_6618,N_6625);
and U7368 (N_7368,N_6758,N_6940);
nor U7369 (N_7369,N_7052,N_7136);
and U7370 (N_7370,N_6950,N_6844);
nor U7371 (N_7371,N_7008,N_6792);
or U7372 (N_7372,N_6991,N_7165);
xnor U7373 (N_7373,N_6882,N_6671);
and U7374 (N_7374,N_6607,N_6639);
nor U7375 (N_7375,N_6706,N_6839);
nand U7376 (N_7376,N_7005,N_6927);
nand U7377 (N_7377,N_7077,N_7169);
or U7378 (N_7378,N_7083,N_6833);
nor U7379 (N_7379,N_6689,N_6578);
and U7380 (N_7380,N_6620,N_7091);
or U7381 (N_7381,N_6938,N_6493);
nor U7382 (N_7382,N_6573,N_6690);
or U7383 (N_7383,N_6837,N_6751);
nand U7384 (N_7384,N_6725,N_7180);
nand U7385 (N_7385,N_6803,N_6768);
and U7386 (N_7386,N_6426,N_6702);
nand U7387 (N_7387,N_6773,N_6494);
and U7388 (N_7388,N_6503,N_6710);
or U7389 (N_7389,N_6612,N_6561);
nor U7390 (N_7390,N_6871,N_7189);
nand U7391 (N_7391,N_6861,N_6693);
and U7392 (N_7392,N_7167,N_6843);
nand U7393 (N_7393,N_6902,N_6770);
nor U7394 (N_7394,N_7145,N_6500);
nand U7395 (N_7395,N_6995,N_6544);
nor U7396 (N_7396,N_6505,N_6872);
nand U7397 (N_7397,N_6667,N_6659);
nor U7398 (N_7398,N_6423,N_7070);
nand U7399 (N_7399,N_6595,N_6996);
or U7400 (N_7400,N_7197,N_6846);
and U7401 (N_7401,N_6877,N_6609);
nand U7402 (N_7402,N_7102,N_6755);
or U7403 (N_7403,N_6454,N_6646);
or U7404 (N_7404,N_6436,N_6731);
nand U7405 (N_7405,N_6579,N_6679);
and U7406 (N_7406,N_6703,N_6993);
nor U7407 (N_7407,N_6686,N_6799);
and U7408 (N_7408,N_6658,N_6429);
and U7409 (N_7409,N_6418,N_7061);
and U7410 (N_7410,N_7194,N_6784);
and U7411 (N_7411,N_6519,N_6896);
nor U7412 (N_7412,N_7006,N_6763);
nand U7413 (N_7413,N_6553,N_6983);
nor U7414 (N_7414,N_6577,N_6428);
and U7415 (N_7415,N_6830,N_6593);
and U7416 (N_7416,N_6911,N_6917);
nor U7417 (N_7417,N_6947,N_6529);
nand U7418 (N_7418,N_6986,N_6524);
and U7419 (N_7419,N_6951,N_7177);
and U7420 (N_7420,N_6520,N_6900);
nor U7421 (N_7421,N_6984,N_7086);
and U7422 (N_7422,N_6740,N_6645);
nand U7423 (N_7423,N_6883,N_6552);
or U7424 (N_7424,N_6776,N_7185);
and U7425 (N_7425,N_6443,N_7107);
xnor U7426 (N_7426,N_6453,N_6432);
nor U7427 (N_7427,N_6715,N_7124);
or U7428 (N_7428,N_6707,N_7011);
or U7429 (N_7429,N_6651,N_6875);
and U7430 (N_7430,N_6977,N_6594);
nand U7431 (N_7431,N_6473,N_6462);
nor U7432 (N_7432,N_6727,N_6414);
nand U7433 (N_7433,N_6956,N_6403);
and U7434 (N_7434,N_6747,N_6973);
nand U7435 (N_7435,N_7106,N_6459);
nor U7436 (N_7436,N_6756,N_6516);
nand U7437 (N_7437,N_6845,N_6979);
nor U7438 (N_7438,N_7087,N_7051);
nand U7439 (N_7439,N_7032,N_6464);
nand U7440 (N_7440,N_6508,N_7195);
nor U7441 (N_7441,N_6924,N_6893);
nor U7442 (N_7442,N_6775,N_6551);
nand U7443 (N_7443,N_6935,N_6746);
nand U7444 (N_7444,N_6674,N_6894);
nor U7445 (N_7445,N_6656,N_7056);
or U7446 (N_7446,N_6629,N_7129);
or U7447 (N_7447,N_6441,N_6613);
nand U7448 (N_7448,N_6623,N_6683);
nor U7449 (N_7449,N_7110,N_6908);
or U7450 (N_7450,N_6780,N_7009);
or U7451 (N_7451,N_6635,N_6966);
or U7452 (N_7452,N_6804,N_7016);
nand U7453 (N_7453,N_6603,N_7160);
nor U7454 (N_7454,N_6557,N_6913);
nor U7455 (N_7455,N_6619,N_6791);
nor U7456 (N_7456,N_6808,N_7060);
nand U7457 (N_7457,N_7137,N_6678);
and U7458 (N_7458,N_6531,N_6440);
xnor U7459 (N_7459,N_6507,N_6624);
and U7460 (N_7460,N_7071,N_6836);
or U7461 (N_7461,N_6764,N_6598);
nor U7462 (N_7462,N_6649,N_6794);
or U7463 (N_7463,N_7158,N_6474);
and U7464 (N_7464,N_6642,N_6970);
nor U7465 (N_7465,N_6701,N_6630);
or U7466 (N_7466,N_6434,N_6818);
nand U7467 (N_7467,N_6488,N_6676);
nor U7468 (N_7468,N_7075,N_6901);
nor U7469 (N_7469,N_7133,N_6820);
or U7470 (N_7470,N_7025,N_7038);
nor U7471 (N_7471,N_6564,N_7069);
nand U7472 (N_7472,N_7156,N_7184);
nor U7473 (N_7473,N_6824,N_6611);
nand U7474 (N_7474,N_6895,N_6862);
nand U7475 (N_7475,N_6848,N_7017);
nand U7476 (N_7476,N_6713,N_7053);
and U7477 (N_7477,N_6813,N_7030);
or U7478 (N_7478,N_6601,N_6615);
nand U7479 (N_7479,N_7095,N_7103);
nand U7480 (N_7480,N_6536,N_6638);
or U7481 (N_7481,N_6948,N_6735);
nor U7482 (N_7482,N_6496,N_6481);
nor U7483 (N_7483,N_6419,N_6944);
nand U7484 (N_7484,N_6497,N_6501);
and U7485 (N_7485,N_7112,N_7072);
nor U7486 (N_7486,N_6739,N_6980);
or U7487 (N_7487,N_6677,N_7174);
nor U7488 (N_7488,N_6614,N_6745);
or U7489 (N_7489,N_6451,N_6999);
or U7490 (N_7490,N_6767,N_6416);
or U7491 (N_7491,N_6729,N_6937);
nand U7492 (N_7492,N_6555,N_6662);
or U7493 (N_7493,N_6860,N_6694);
nor U7494 (N_7494,N_6589,N_7093);
and U7495 (N_7495,N_6468,N_6680);
and U7496 (N_7496,N_6424,N_7130);
nand U7497 (N_7497,N_7022,N_6406);
nor U7498 (N_7498,N_7118,N_6538);
nand U7499 (N_7499,N_6631,N_6712);
nor U7500 (N_7500,N_6554,N_6880);
nor U7501 (N_7501,N_7191,N_6750);
and U7502 (N_7502,N_6504,N_6992);
and U7503 (N_7503,N_6771,N_6828);
nand U7504 (N_7504,N_6663,N_6576);
or U7505 (N_7505,N_7164,N_7188);
nor U7506 (N_7506,N_7166,N_6743);
nor U7507 (N_7507,N_6777,N_6648);
or U7508 (N_7508,N_7000,N_6586);
nor U7509 (N_7509,N_6550,N_6521);
and U7510 (N_7510,N_6874,N_6732);
and U7511 (N_7511,N_6802,N_6752);
nand U7512 (N_7512,N_6637,N_6461);
and U7513 (N_7513,N_6647,N_6781);
nor U7514 (N_7514,N_6446,N_6933);
nor U7515 (N_7515,N_7096,N_6779);
nand U7516 (N_7516,N_6914,N_6585);
nand U7517 (N_7517,N_6572,N_7126);
and U7518 (N_7518,N_6997,N_6821);
nor U7519 (N_7519,N_6866,N_6960);
and U7520 (N_7520,N_7042,N_7063);
and U7521 (N_7521,N_6988,N_6854);
xor U7522 (N_7522,N_7175,N_6826);
nor U7523 (N_7523,N_7147,N_7019);
or U7524 (N_7524,N_6870,N_6460);
nand U7525 (N_7525,N_6856,N_6404);
nor U7526 (N_7526,N_6806,N_6719);
nor U7527 (N_7527,N_7058,N_7172);
nor U7528 (N_7528,N_6717,N_6858);
nand U7529 (N_7529,N_6890,N_6522);
and U7530 (N_7530,N_6964,N_6832);
and U7531 (N_7531,N_6994,N_6766);
nand U7532 (N_7532,N_7078,N_6660);
nand U7533 (N_7533,N_6785,N_6721);
or U7534 (N_7534,N_6814,N_6868);
and U7535 (N_7535,N_7196,N_6470);
and U7536 (N_7536,N_6954,N_6916);
and U7537 (N_7537,N_7176,N_6643);
or U7538 (N_7538,N_7062,N_6587);
and U7539 (N_7539,N_6798,N_6599);
nor U7540 (N_7540,N_6514,N_6795);
nand U7541 (N_7541,N_7081,N_6608);
and U7542 (N_7542,N_6449,N_6873);
nor U7543 (N_7543,N_6943,N_6408);
nand U7544 (N_7544,N_7036,N_6410);
nor U7545 (N_7545,N_7055,N_6793);
nand U7546 (N_7546,N_7122,N_6563);
or U7547 (N_7547,N_6466,N_6407);
and U7548 (N_7548,N_6422,N_6540);
or U7549 (N_7549,N_6859,N_7116);
and U7550 (N_7550,N_7143,N_6709);
and U7551 (N_7551,N_6811,N_7173);
nand U7552 (N_7552,N_6974,N_6596);
and U7553 (N_7553,N_6737,N_6692);
xor U7554 (N_7554,N_6728,N_7067);
or U7555 (N_7555,N_6819,N_6723);
nand U7556 (N_7556,N_6512,N_7021);
or U7557 (N_7557,N_6891,N_7138);
and U7558 (N_7558,N_6654,N_6886);
nor U7559 (N_7559,N_6711,N_6528);
nor U7560 (N_7560,N_6489,N_6506);
nand U7561 (N_7561,N_6541,N_6923);
xnor U7562 (N_7562,N_7190,N_6532);
nand U7563 (N_7563,N_7153,N_7013);
and U7564 (N_7564,N_7120,N_6568);
or U7565 (N_7565,N_6885,N_7044);
nor U7566 (N_7566,N_6716,N_6669);
nand U7567 (N_7567,N_7144,N_6990);
and U7568 (N_7568,N_6546,N_6517);
nor U7569 (N_7569,N_7108,N_6666);
nor U7570 (N_7570,N_6857,N_6952);
and U7571 (N_7571,N_6959,N_6487);
and U7572 (N_7572,N_6936,N_6681);
or U7573 (N_7573,N_7097,N_6981);
nand U7574 (N_7574,N_6918,N_6571);
nor U7575 (N_7575,N_6698,N_6749);
or U7576 (N_7576,N_6588,N_7090);
and U7577 (N_7577,N_7047,N_6670);
nand U7578 (N_7578,N_6975,N_6957);
and U7579 (N_7579,N_6931,N_7092);
nor U7580 (N_7580,N_6765,N_7040);
or U7581 (N_7581,N_6699,N_6809);
and U7582 (N_7582,N_6797,N_7007);
and U7583 (N_7583,N_6942,N_7198);
nor U7584 (N_7584,N_6547,N_6580);
or U7585 (N_7585,N_6626,N_6926);
nand U7586 (N_7586,N_6491,N_7134);
nand U7587 (N_7587,N_6934,N_6545);
or U7588 (N_7588,N_6617,N_6539);
nor U7589 (N_7589,N_7109,N_6741);
nand U7590 (N_7590,N_6673,N_6535);
or U7591 (N_7591,N_6949,N_7084);
and U7592 (N_7592,N_6682,N_6479);
nand U7593 (N_7593,N_6963,N_6801);
or U7594 (N_7594,N_6627,N_6592);
or U7595 (N_7595,N_6492,N_6783);
nand U7596 (N_7596,N_7001,N_7029);
nor U7597 (N_7597,N_6411,N_6887);
or U7598 (N_7598,N_6452,N_6405);
and U7599 (N_7599,N_6560,N_6985);
and U7600 (N_7600,N_7136,N_7094);
or U7601 (N_7601,N_6911,N_6786);
or U7602 (N_7602,N_6542,N_6840);
and U7603 (N_7603,N_6646,N_6680);
and U7604 (N_7604,N_6951,N_6503);
and U7605 (N_7605,N_6789,N_6863);
nand U7606 (N_7606,N_6547,N_7192);
nand U7607 (N_7607,N_6631,N_6793);
and U7608 (N_7608,N_6611,N_6640);
and U7609 (N_7609,N_6454,N_6616);
nor U7610 (N_7610,N_6801,N_6942);
nand U7611 (N_7611,N_6856,N_7050);
or U7612 (N_7612,N_6913,N_6443);
nand U7613 (N_7613,N_6624,N_7151);
nor U7614 (N_7614,N_6549,N_6766);
nand U7615 (N_7615,N_7078,N_6511);
nand U7616 (N_7616,N_6707,N_7107);
and U7617 (N_7617,N_7086,N_6606);
nor U7618 (N_7618,N_6562,N_7172);
nor U7619 (N_7619,N_6418,N_6748);
nor U7620 (N_7620,N_7024,N_6622);
and U7621 (N_7621,N_6897,N_6964);
nand U7622 (N_7622,N_6949,N_6460);
and U7623 (N_7623,N_6563,N_6698);
nand U7624 (N_7624,N_6904,N_6951);
nand U7625 (N_7625,N_7079,N_6719);
and U7626 (N_7626,N_6480,N_7011);
or U7627 (N_7627,N_6948,N_7140);
nand U7628 (N_7628,N_7185,N_6688);
and U7629 (N_7629,N_7022,N_6939);
and U7630 (N_7630,N_6779,N_6751);
nand U7631 (N_7631,N_6722,N_7015);
nand U7632 (N_7632,N_6680,N_6601);
nand U7633 (N_7633,N_7010,N_7122);
or U7634 (N_7634,N_6561,N_6657);
nor U7635 (N_7635,N_6599,N_6659);
and U7636 (N_7636,N_6801,N_6718);
nor U7637 (N_7637,N_7126,N_6980);
or U7638 (N_7638,N_6978,N_6518);
nand U7639 (N_7639,N_6693,N_6414);
and U7640 (N_7640,N_6873,N_6567);
nor U7641 (N_7641,N_6790,N_6744);
or U7642 (N_7642,N_6751,N_6691);
xnor U7643 (N_7643,N_6786,N_7042);
and U7644 (N_7644,N_6720,N_6831);
nand U7645 (N_7645,N_6619,N_7172);
and U7646 (N_7646,N_6449,N_6970);
or U7647 (N_7647,N_6646,N_6644);
and U7648 (N_7648,N_6724,N_6927);
or U7649 (N_7649,N_7141,N_6644);
and U7650 (N_7650,N_6925,N_6955);
nor U7651 (N_7651,N_6771,N_7033);
nor U7652 (N_7652,N_6769,N_6481);
nor U7653 (N_7653,N_7018,N_6901);
nand U7654 (N_7654,N_7104,N_6460);
nor U7655 (N_7655,N_7019,N_6823);
and U7656 (N_7656,N_6925,N_6428);
or U7657 (N_7657,N_7062,N_7043);
nor U7658 (N_7658,N_7051,N_7000);
and U7659 (N_7659,N_6528,N_7156);
nor U7660 (N_7660,N_6971,N_6841);
nand U7661 (N_7661,N_6836,N_6433);
nor U7662 (N_7662,N_6558,N_6612);
and U7663 (N_7663,N_6678,N_7151);
or U7664 (N_7664,N_6709,N_6884);
and U7665 (N_7665,N_7164,N_7013);
and U7666 (N_7666,N_6422,N_6923);
and U7667 (N_7667,N_6780,N_7045);
and U7668 (N_7668,N_6538,N_6446);
and U7669 (N_7669,N_6447,N_6538);
and U7670 (N_7670,N_7004,N_7162);
and U7671 (N_7671,N_6457,N_6731);
or U7672 (N_7672,N_6869,N_6668);
nand U7673 (N_7673,N_7107,N_6935);
nor U7674 (N_7674,N_6918,N_7092);
or U7675 (N_7675,N_6671,N_6768);
nor U7676 (N_7676,N_6877,N_6464);
nand U7677 (N_7677,N_7063,N_6605);
nor U7678 (N_7678,N_6639,N_6847);
nor U7679 (N_7679,N_6899,N_6822);
and U7680 (N_7680,N_6960,N_6676);
and U7681 (N_7681,N_6892,N_6612);
or U7682 (N_7682,N_6788,N_6767);
nand U7683 (N_7683,N_6642,N_7077);
nand U7684 (N_7684,N_6616,N_6713);
nor U7685 (N_7685,N_6461,N_6814);
nand U7686 (N_7686,N_6548,N_7180);
nand U7687 (N_7687,N_6874,N_6748);
nor U7688 (N_7688,N_6834,N_6501);
or U7689 (N_7689,N_6519,N_6805);
and U7690 (N_7690,N_6461,N_6581);
nor U7691 (N_7691,N_6662,N_7001);
nor U7692 (N_7692,N_7008,N_6762);
xnor U7693 (N_7693,N_6706,N_6937);
and U7694 (N_7694,N_7148,N_6971);
and U7695 (N_7695,N_7118,N_6659);
nand U7696 (N_7696,N_6575,N_6467);
nand U7697 (N_7697,N_7033,N_7088);
or U7698 (N_7698,N_6911,N_7047);
nand U7699 (N_7699,N_6550,N_7189);
nand U7700 (N_7700,N_6438,N_6638);
or U7701 (N_7701,N_6905,N_7017);
and U7702 (N_7702,N_6708,N_6402);
nor U7703 (N_7703,N_6542,N_6608);
xor U7704 (N_7704,N_6493,N_7153);
nand U7705 (N_7705,N_6479,N_6463);
or U7706 (N_7706,N_7164,N_6424);
nor U7707 (N_7707,N_6794,N_6749);
and U7708 (N_7708,N_7137,N_6647);
or U7709 (N_7709,N_6459,N_6638);
nand U7710 (N_7710,N_7194,N_6803);
and U7711 (N_7711,N_6796,N_6836);
and U7712 (N_7712,N_6783,N_7036);
and U7713 (N_7713,N_6445,N_6410);
nand U7714 (N_7714,N_7062,N_7159);
or U7715 (N_7715,N_6693,N_7157);
or U7716 (N_7716,N_6658,N_6798);
and U7717 (N_7717,N_6733,N_6742);
or U7718 (N_7718,N_6982,N_6934);
nor U7719 (N_7719,N_7041,N_6964);
nor U7720 (N_7720,N_6858,N_6492);
or U7721 (N_7721,N_6763,N_7137);
and U7722 (N_7722,N_6404,N_6482);
nand U7723 (N_7723,N_7193,N_7161);
nand U7724 (N_7724,N_6615,N_6828);
nor U7725 (N_7725,N_6506,N_6928);
nor U7726 (N_7726,N_6563,N_7129);
or U7727 (N_7727,N_7011,N_6856);
or U7728 (N_7728,N_6905,N_6417);
or U7729 (N_7729,N_6545,N_6484);
nor U7730 (N_7730,N_7006,N_6444);
or U7731 (N_7731,N_6446,N_7036);
nor U7732 (N_7732,N_6625,N_7180);
nor U7733 (N_7733,N_6722,N_6960);
or U7734 (N_7734,N_6633,N_6793);
or U7735 (N_7735,N_6969,N_7004);
or U7736 (N_7736,N_6723,N_6428);
nor U7737 (N_7737,N_6448,N_7186);
and U7738 (N_7738,N_7039,N_6581);
and U7739 (N_7739,N_6881,N_6433);
and U7740 (N_7740,N_7123,N_6804);
nor U7741 (N_7741,N_6426,N_6655);
nand U7742 (N_7742,N_6419,N_7131);
nand U7743 (N_7743,N_6774,N_6972);
nor U7744 (N_7744,N_6709,N_6893);
nor U7745 (N_7745,N_6413,N_6864);
and U7746 (N_7746,N_6414,N_6515);
nor U7747 (N_7747,N_6418,N_6511);
nand U7748 (N_7748,N_6531,N_7065);
nand U7749 (N_7749,N_6577,N_7042);
or U7750 (N_7750,N_6620,N_6818);
nor U7751 (N_7751,N_7023,N_6804);
nor U7752 (N_7752,N_6840,N_6501);
nand U7753 (N_7753,N_7065,N_7052);
nand U7754 (N_7754,N_6797,N_6474);
nor U7755 (N_7755,N_6653,N_6511);
xor U7756 (N_7756,N_7100,N_6574);
and U7757 (N_7757,N_6885,N_6702);
nand U7758 (N_7758,N_6661,N_6850);
nand U7759 (N_7759,N_6729,N_6640);
nand U7760 (N_7760,N_6485,N_6901);
nand U7761 (N_7761,N_7109,N_6403);
nor U7762 (N_7762,N_6555,N_6979);
and U7763 (N_7763,N_7026,N_6553);
and U7764 (N_7764,N_6600,N_6933);
and U7765 (N_7765,N_6474,N_6484);
or U7766 (N_7766,N_7177,N_7009);
and U7767 (N_7767,N_6595,N_6867);
or U7768 (N_7768,N_6699,N_6492);
and U7769 (N_7769,N_6455,N_6807);
and U7770 (N_7770,N_6507,N_7123);
nand U7771 (N_7771,N_6911,N_6823);
and U7772 (N_7772,N_6990,N_6756);
or U7773 (N_7773,N_7125,N_6456);
nand U7774 (N_7774,N_6444,N_7042);
or U7775 (N_7775,N_7027,N_6412);
nand U7776 (N_7776,N_6781,N_6854);
and U7777 (N_7777,N_6695,N_7030);
nand U7778 (N_7778,N_6775,N_6439);
or U7779 (N_7779,N_6702,N_7081);
nand U7780 (N_7780,N_6468,N_6436);
or U7781 (N_7781,N_6841,N_6827);
or U7782 (N_7782,N_7105,N_6494);
nand U7783 (N_7783,N_6466,N_7035);
or U7784 (N_7784,N_6716,N_7160);
or U7785 (N_7785,N_6472,N_6556);
or U7786 (N_7786,N_7197,N_6952);
nor U7787 (N_7787,N_6508,N_6590);
nor U7788 (N_7788,N_7133,N_7149);
and U7789 (N_7789,N_6716,N_6510);
nand U7790 (N_7790,N_6489,N_6991);
nor U7791 (N_7791,N_6450,N_6948);
nor U7792 (N_7792,N_6580,N_6840);
or U7793 (N_7793,N_6539,N_6813);
and U7794 (N_7794,N_7062,N_6475);
xor U7795 (N_7795,N_7154,N_6640);
nor U7796 (N_7796,N_7013,N_7120);
nand U7797 (N_7797,N_6948,N_7029);
and U7798 (N_7798,N_6682,N_7025);
and U7799 (N_7799,N_6800,N_7127);
and U7800 (N_7800,N_7060,N_6849);
nor U7801 (N_7801,N_6567,N_6529);
nor U7802 (N_7802,N_6899,N_7132);
nor U7803 (N_7803,N_6997,N_6695);
or U7804 (N_7804,N_6663,N_6588);
nor U7805 (N_7805,N_6462,N_6705);
and U7806 (N_7806,N_6753,N_6926);
and U7807 (N_7807,N_7129,N_7115);
nand U7808 (N_7808,N_7106,N_7072);
and U7809 (N_7809,N_6452,N_6591);
or U7810 (N_7810,N_6874,N_6677);
nand U7811 (N_7811,N_6578,N_6699);
nand U7812 (N_7812,N_6884,N_6552);
nand U7813 (N_7813,N_7126,N_6988);
nor U7814 (N_7814,N_6475,N_6463);
nor U7815 (N_7815,N_6672,N_6590);
nand U7816 (N_7816,N_6945,N_6416);
nor U7817 (N_7817,N_6430,N_7146);
nor U7818 (N_7818,N_7058,N_6676);
nand U7819 (N_7819,N_7074,N_6506);
nand U7820 (N_7820,N_6832,N_6718);
or U7821 (N_7821,N_6442,N_6705);
and U7822 (N_7822,N_7075,N_7059);
and U7823 (N_7823,N_7182,N_6643);
nor U7824 (N_7824,N_6913,N_6535);
and U7825 (N_7825,N_6726,N_6789);
xor U7826 (N_7826,N_6538,N_7022);
and U7827 (N_7827,N_6796,N_6906);
nor U7828 (N_7828,N_7035,N_6773);
and U7829 (N_7829,N_6745,N_6785);
and U7830 (N_7830,N_6444,N_7137);
or U7831 (N_7831,N_6910,N_6822);
nand U7832 (N_7832,N_6444,N_7005);
or U7833 (N_7833,N_6955,N_6832);
nand U7834 (N_7834,N_6851,N_6789);
and U7835 (N_7835,N_6678,N_6889);
nor U7836 (N_7836,N_7113,N_6485);
nand U7837 (N_7837,N_6724,N_6552);
nor U7838 (N_7838,N_6676,N_6889);
and U7839 (N_7839,N_7080,N_6801);
nand U7840 (N_7840,N_6690,N_6916);
xnor U7841 (N_7841,N_6505,N_6891);
and U7842 (N_7842,N_6981,N_6916);
and U7843 (N_7843,N_6941,N_6801);
nor U7844 (N_7844,N_7066,N_6716);
nor U7845 (N_7845,N_6541,N_6537);
nand U7846 (N_7846,N_7170,N_6932);
nor U7847 (N_7847,N_6774,N_6451);
nor U7848 (N_7848,N_6734,N_6863);
nand U7849 (N_7849,N_6607,N_6864);
and U7850 (N_7850,N_7122,N_7169);
and U7851 (N_7851,N_6975,N_6866);
or U7852 (N_7852,N_6859,N_7074);
or U7853 (N_7853,N_6918,N_6919);
and U7854 (N_7854,N_7119,N_6522);
or U7855 (N_7855,N_6814,N_6491);
and U7856 (N_7856,N_6733,N_6819);
or U7857 (N_7857,N_6713,N_6458);
nand U7858 (N_7858,N_6942,N_6564);
or U7859 (N_7859,N_6958,N_6914);
and U7860 (N_7860,N_6527,N_6661);
or U7861 (N_7861,N_6766,N_6419);
nand U7862 (N_7862,N_7088,N_6577);
or U7863 (N_7863,N_6663,N_7120);
and U7864 (N_7864,N_6582,N_6804);
or U7865 (N_7865,N_6468,N_7147);
nand U7866 (N_7866,N_7134,N_7042);
and U7867 (N_7867,N_6864,N_7160);
and U7868 (N_7868,N_6549,N_7177);
nor U7869 (N_7869,N_7093,N_6437);
nor U7870 (N_7870,N_6789,N_6892);
or U7871 (N_7871,N_6927,N_6818);
or U7872 (N_7872,N_7124,N_6600);
nor U7873 (N_7873,N_6563,N_6410);
and U7874 (N_7874,N_7025,N_6944);
nand U7875 (N_7875,N_6600,N_7039);
nor U7876 (N_7876,N_6402,N_6628);
or U7877 (N_7877,N_6911,N_7114);
nand U7878 (N_7878,N_6724,N_6511);
or U7879 (N_7879,N_6918,N_6668);
or U7880 (N_7880,N_6623,N_6946);
nand U7881 (N_7881,N_6673,N_6973);
nand U7882 (N_7882,N_6655,N_6919);
xor U7883 (N_7883,N_6865,N_6743);
nor U7884 (N_7884,N_6951,N_6403);
nor U7885 (N_7885,N_6446,N_6570);
nand U7886 (N_7886,N_6598,N_7127);
nand U7887 (N_7887,N_6584,N_6712);
xor U7888 (N_7888,N_7146,N_6837);
and U7889 (N_7889,N_7199,N_7100);
nand U7890 (N_7890,N_7150,N_6778);
nor U7891 (N_7891,N_6878,N_6855);
and U7892 (N_7892,N_7116,N_6944);
nor U7893 (N_7893,N_6950,N_6715);
or U7894 (N_7894,N_6674,N_6785);
or U7895 (N_7895,N_6784,N_6637);
or U7896 (N_7896,N_6616,N_6886);
nand U7897 (N_7897,N_6890,N_7063);
nor U7898 (N_7898,N_6717,N_6498);
and U7899 (N_7899,N_6451,N_6874);
nand U7900 (N_7900,N_7091,N_6680);
nor U7901 (N_7901,N_6922,N_6883);
nand U7902 (N_7902,N_6984,N_6432);
nor U7903 (N_7903,N_6748,N_6811);
and U7904 (N_7904,N_7092,N_6809);
nor U7905 (N_7905,N_6641,N_7021);
and U7906 (N_7906,N_6504,N_7025);
and U7907 (N_7907,N_6849,N_6914);
nand U7908 (N_7908,N_6825,N_6854);
nor U7909 (N_7909,N_6890,N_6518);
nor U7910 (N_7910,N_6496,N_6592);
or U7911 (N_7911,N_6655,N_6759);
nor U7912 (N_7912,N_6748,N_7152);
nand U7913 (N_7913,N_6680,N_6550);
nor U7914 (N_7914,N_6644,N_6457);
or U7915 (N_7915,N_6467,N_6745);
nor U7916 (N_7916,N_6863,N_6982);
or U7917 (N_7917,N_6734,N_6402);
nor U7918 (N_7918,N_6600,N_7011);
or U7919 (N_7919,N_6571,N_6793);
nor U7920 (N_7920,N_6909,N_7162);
nor U7921 (N_7921,N_6413,N_6462);
or U7922 (N_7922,N_6408,N_6767);
nor U7923 (N_7923,N_6581,N_6676);
or U7924 (N_7924,N_6728,N_6909);
and U7925 (N_7925,N_6925,N_7035);
and U7926 (N_7926,N_7024,N_6739);
or U7927 (N_7927,N_7113,N_7132);
nand U7928 (N_7928,N_7168,N_7153);
or U7929 (N_7929,N_6587,N_6672);
nor U7930 (N_7930,N_6676,N_7170);
or U7931 (N_7931,N_7186,N_6852);
nand U7932 (N_7932,N_6564,N_7064);
nand U7933 (N_7933,N_6811,N_7065);
nand U7934 (N_7934,N_7117,N_6787);
nor U7935 (N_7935,N_6522,N_6672);
and U7936 (N_7936,N_6938,N_6482);
nand U7937 (N_7937,N_6983,N_7030);
or U7938 (N_7938,N_6934,N_6500);
nor U7939 (N_7939,N_6731,N_6803);
or U7940 (N_7940,N_6730,N_6500);
nor U7941 (N_7941,N_6998,N_6874);
and U7942 (N_7942,N_6465,N_7180);
or U7943 (N_7943,N_7044,N_6716);
nand U7944 (N_7944,N_6593,N_6720);
and U7945 (N_7945,N_6886,N_6450);
nor U7946 (N_7946,N_7137,N_6616);
or U7947 (N_7947,N_6592,N_6758);
nand U7948 (N_7948,N_6423,N_6542);
nand U7949 (N_7949,N_7114,N_7113);
or U7950 (N_7950,N_6865,N_7001);
and U7951 (N_7951,N_6758,N_6993);
and U7952 (N_7952,N_6651,N_6730);
or U7953 (N_7953,N_7106,N_6880);
nor U7954 (N_7954,N_6728,N_6452);
nor U7955 (N_7955,N_6704,N_6706);
or U7956 (N_7956,N_6506,N_6727);
nor U7957 (N_7957,N_6485,N_7047);
and U7958 (N_7958,N_6479,N_7043);
nand U7959 (N_7959,N_6684,N_7034);
and U7960 (N_7960,N_6822,N_7187);
and U7961 (N_7961,N_7139,N_6615);
nor U7962 (N_7962,N_6609,N_6553);
and U7963 (N_7963,N_7019,N_6932);
nand U7964 (N_7964,N_7174,N_6652);
nor U7965 (N_7965,N_6713,N_6829);
and U7966 (N_7966,N_6466,N_7001);
nand U7967 (N_7967,N_6744,N_6954);
nand U7968 (N_7968,N_6637,N_6544);
nor U7969 (N_7969,N_6789,N_6766);
or U7970 (N_7970,N_7194,N_6750);
nand U7971 (N_7971,N_6449,N_6985);
or U7972 (N_7972,N_6595,N_6725);
nand U7973 (N_7973,N_6470,N_6625);
or U7974 (N_7974,N_6470,N_6538);
or U7975 (N_7975,N_7175,N_6741);
and U7976 (N_7976,N_6809,N_6683);
nand U7977 (N_7977,N_7187,N_6513);
xor U7978 (N_7978,N_6485,N_7067);
nand U7979 (N_7979,N_6515,N_7034);
nand U7980 (N_7980,N_6487,N_6879);
nand U7981 (N_7981,N_6971,N_6961);
or U7982 (N_7982,N_7144,N_6773);
or U7983 (N_7983,N_6645,N_6575);
nand U7984 (N_7984,N_6652,N_7020);
and U7985 (N_7985,N_6970,N_6772);
nand U7986 (N_7986,N_6599,N_6727);
nor U7987 (N_7987,N_6996,N_7104);
or U7988 (N_7988,N_7065,N_6933);
nor U7989 (N_7989,N_6689,N_6513);
or U7990 (N_7990,N_6604,N_7085);
nand U7991 (N_7991,N_7149,N_7090);
and U7992 (N_7992,N_6728,N_6520);
nor U7993 (N_7993,N_6600,N_6496);
xor U7994 (N_7994,N_6591,N_6649);
nor U7995 (N_7995,N_7033,N_6662);
or U7996 (N_7996,N_6778,N_6866);
or U7997 (N_7997,N_6565,N_6709);
nand U7998 (N_7998,N_6458,N_6604);
nor U7999 (N_7999,N_7105,N_6641);
nand U8000 (N_8000,N_7462,N_7702);
and U8001 (N_8001,N_7427,N_7251);
and U8002 (N_8002,N_7529,N_7336);
or U8003 (N_8003,N_7925,N_7543);
or U8004 (N_8004,N_7210,N_7709);
or U8005 (N_8005,N_7971,N_7517);
nand U8006 (N_8006,N_7293,N_7376);
or U8007 (N_8007,N_7393,N_7322);
nand U8008 (N_8008,N_7213,N_7843);
and U8009 (N_8009,N_7233,N_7962);
nor U8010 (N_8010,N_7915,N_7568);
nor U8011 (N_8011,N_7435,N_7642);
nand U8012 (N_8012,N_7514,N_7919);
nor U8013 (N_8013,N_7380,N_7283);
or U8014 (N_8014,N_7747,N_7476);
xor U8015 (N_8015,N_7585,N_7533);
or U8016 (N_8016,N_7384,N_7984);
nor U8017 (N_8017,N_7742,N_7878);
and U8018 (N_8018,N_7409,N_7227);
nor U8019 (N_8019,N_7209,N_7350);
and U8020 (N_8020,N_7442,N_7386);
and U8021 (N_8021,N_7626,N_7692);
nand U8022 (N_8022,N_7250,N_7866);
or U8023 (N_8023,N_7707,N_7817);
or U8024 (N_8024,N_7872,N_7601);
and U8025 (N_8025,N_7357,N_7578);
and U8026 (N_8026,N_7847,N_7206);
and U8027 (N_8027,N_7666,N_7657);
nand U8028 (N_8028,N_7965,N_7934);
nand U8029 (N_8029,N_7299,N_7994);
or U8030 (N_8030,N_7257,N_7977);
or U8031 (N_8031,N_7683,N_7445);
and U8032 (N_8032,N_7773,N_7697);
nor U8033 (N_8033,N_7502,N_7289);
and U8034 (N_8034,N_7887,N_7252);
nor U8035 (N_8035,N_7495,N_7775);
or U8036 (N_8036,N_7248,N_7906);
and U8037 (N_8037,N_7733,N_7914);
or U8038 (N_8038,N_7497,N_7216);
nand U8039 (N_8039,N_7649,N_7762);
or U8040 (N_8040,N_7620,N_7602);
and U8041 (N_8041,N_7754,N_7777);
nor U8042 (N_8042,N_7875,N_7761);
or U8043 (N_8043,N_7413,N_7416);
nor U8044 (N_8044,N_7833,N_7218);
nor U8045 (N_8045,N_7629,N_7461);
nand U8046 (N_8046,N_7758,N_7301);
nor U8047 (N_8047,N_7418,N_7896);
and U8048 (N_8048,N_7766,N_7904);
nor U8049 (N_8049,N_7550,N_7411);
nand U8050 (N_8050,N_7610,N_7217);
or U8051 (N_8051,N_7487,N_7600);
xnor U8052 (N_8052,N_7979,N_7499);
and U8053 (N_8053,N_7687,N_7832);
nand U8054 (N_8054,N_7682,N_7716);
or U8055 (N_8055,N_7249,N_7615);
or U8056 (N_8056,N_7563,N_7661);
nand U8057 (N_8057,N_7797,N_7912);
or U8058 (N_8058,N_7272,N_7720);
and U8059 (N_8059,N_7268,N_7963);
and U8060 (N_8060,N_7698,N_7911);
or U8061 (N_8061,N_7735,N_7451);
or U8062 (N_8062,N_7243,N_7907);
nor U8063 (N_8063,N_7638,N_7220);
nor U8064 (N_8064,N_7830,N_7458);
and U8065 (N_8065,N_7814,N_7236);
and U8066 (N_8066,N_7808,N_7894);
nand U8067 (N_8067,N_7329,N_7910);
nor U8068 (N_8068,N_7711,N_7569);
and U8069 (N_8069,N_7799,N_7399);
or U8070 (N_8070,N_7890,N_7996);
nand U8071 (N_8071,N_7245,N_7515);
and U8072 (N_8072,N_7490,N_7860);
or U8073 (N_8073,N_7882,N_7884);
or U8074 (N_8074,N_7549,N_7714);
or U8075 (N_8075,N_7855,N_7946);
or U8076 (N_8076,N_7489,N_7675);
or U8077 (N_8077,N_7653,N_7790);
nor U8078 (N_8078,N_7254,N_7391);
nor U8079 (N_8079,N_7846,N_7603);
nor U8080 (N_8080,N_7659,N_7288);
nor U8081 (N_8081,N_7428,N_7385);
and U8082 (N_8082,N_7483,N_7689);
nand U8083 (N_8083,N_7779,N_7957);
nor U8084 (N_8084,N_7486,N_7313);
nor U8085 (N_8085,N_7794,N_7452);
or U8086 (N_8086,N_7504,N_7985);
nand U8087 (N_8087,N_7595,N_7334);
nand U8088 (N_8088,N_7341,N_7240);
nand U8089 (N_8089,N_7287,N_7787);
nand U8090 (N_8090,N_7640,N_7818);
or U8091 (N_8091,N_7879,N_7410);
and U8092 (N_8092,N_7917,N_7309);
nor U8093 (N_8093,N_7810,N_7852);
nor U8094 (N_8094,N_7656,N_7671);
nand U8095 (N_8095,N_7260,N_7774);
nor U8096 (N_8096,N_7732,N_7567);
or U8097 (N_8097,N_7789,N_7749);
nand U8098 (N_8098,N_7282,N_7223);
nor U8099 (N_8099,N_7317,N_7614);
nor U8100 (N_8100,N_7478,N_7425);
nor U8101 (N_8101,N_7718,N_7538);
nand U8102 (N_8102,N_7966,N_7582);
or U8103 (N_8103,N_7423,N_7304);
and U8104 (N_8104,N_7494,N_7881);
and U8105 (N_8105,N_7953,N_7526);
and U8106 (N_8106,N_7364,N_7997);
or U8107 (N_8107,N_7544,N_7536);
and U8108 (N_8108,N_7838,N_7624);
nand U8109 (N_8109,N_7806,N_7202);
nand U8110 (N_8110,N_7905,N_7854);
or U8111 (N_8111,N_7809,N_7856);
or U8112 (N_8112,N_7553,N_7849);
nand U8113 (N_8113,N_7219,N_7440);
nand U8114 (N_8114,N_7546,N_7715);
nand U8115 (N_8115,N_7510,N_7913);
nor U8116 (N_8116,N_7323,N_7545);
nor U8117 (N_8117,N_7920,N_7331);
nor U8118 (N_8118,N_7883,N_7548);
nor U8119 (N_8119,N_7547,N_7850);
nor U8120 (N_8120,N_7763,N_7297);
nand U8121 (N_8121,N_7347,N_7678);
nand U8122 (N_8122,N_7753,N_7888);
nand U8123 (N_8123,N_7650,N_7400);
nand U8124 (N_8124,N_7672,N_7222);
nor U8125 (N_8125,N_7448,N_7255);
or U8126 (N_8126,N_7505,N_7405);
and U8127 (N_8127,N_7348,N_7314);
or U8128 (N_8128,N_7511,N_7340);
and U8129 (N_8129,N_7555,N_7286);
and U8130 (N_8130,N_7464,N_7613);
and U8131 (N_8131,N_7930,N_7467);
and U8132 (N_8132,N_7951,N_7273);
nor U8133 (N_8133,N_7270,N_7414);
nand U8134 (N_8134,N_7561,N_7319);
nand U8135 (N_8135,N_7475,N_7238);
and U8136 (N_8136,N_7537,N_7802);
and U8137 (N_8137,N_7271,N_7383);
nand U8138 (N_8138,N_7767,N_7598);
or U8139 (N_8139,N_7889,N_7933);
nand U8140 (N_8140,N_7433,N_7279);
and U8141 (N_8141,N_7737,N_7916);
nand U8142 (N_8142,N_7447,N_7812);
and U8143 (N_8143,N_7722,N_7394);
or U8144 (N_8144,N_7738,N_7768);
and U8145 (N_8145,N_7275,N_7646);
nand U8146 (N_8146,N_7530,N_7778);
nor U8147 (N_8147,N_7421,N_7324);
and U8148 (N_8148,N_7803,N_7521);
or U8149 (N_8149,N_7622,N_7221);
or U8150 (N_8150,N_7434,N_7586);
and U8151 (N_8151,N_7205,N_7397);
nor U8152 (N_8152,N_7772,N_7744);
and U8153 (N_8153,N_7891,N_7834);
nor U8154 (N_8154,N_7734,N_7437);
nand U8155 (N_8155,N_7660,N_7353);
or U8156 (N_8156,N_7848,N_7858);
nor U8157 (N_8157,N_7302,N_7988);
and U8158 (N_8158,N_7343,N_7954);
nor U8159 (N_8159,N_7691,N_7577);
or U8160 (N_8160,N_7981,N_7668);
and U8161 (N_8161,N_7457,N_7372);
or U8162 (N_8162,N_7296,N_7793);
or U8163 (N_8163,N_7362,N_7696);
nor U8164 (N_8164,N_7474,N_7520);
and U8165 (N_8165,N_7612,N_7332);
and U8166 (N_8166,N_7300,N_7764);
and U8167 (N_8167,N_7584,N_7215);
and U8168 (N_8168,N_7506,N_7999);
or U8169 (N_8169,N_7728,N_7420);
nand U8170 (N_8170,N_7795,N_7825);
or U8171 (N_8171,N_7375,N_7786);
and U8172 (N_8172,N_7518,N_7315);
nor U8173 (N_8173,N_7992,N_7593);
nor U8174 (N_8174,N_7262,N_7345);
nand U8175 (N_8175,N_7842,N_7226);
and U8176 (N_8176,N_7699,N_7897);
nand U8177 (N_8177,N_7677,N_7611);
and U8178 (N_8178,N_7804,N_7280);
or U8179 (N_8179,N_7701,N_7204);
or U8180 (N_8180,N_7756,N_7588);
and U8181 (N_8181,N_7597,N_7318);
nand U8182 (N_8182,N_7880,N_7676);
or U8183 (N_8183,N_7998,N_7869);
or U8184 (N_8184,N_7960,N_7719);
nand U8185 (N_8185,N_7942,N_7581);
or U8186 (N_8186,N_7899,N_7821);
nand U8187 (N_8187,N_7454,N_7944);
and U8188 (N_8188,N_7508,N_7628);
and U8189 (N_8189,N_7713,N_7378);
and U8190 (N_8190,N_7684,N_7829);
nand U8191 (N_8191,N_7940,N_7616);
or U8192 (N_8192,N_7591,N_7757);
or U8193 (N_8193,N_7704,N_7524);
and U8194 (N_8194,N_7673,N_7415);
or U8195 (N_8195,N_7295,N_7239);
nor U8196 (N_8196,N_7473,N_7583);
nor U8197 (N_8197,N_7573,N_7402);
nor U8198 (N_8198,N_7871,N_7463);
and U8199 (N_8199,N_7377,N_7523);
and U8200 (N_8200,N_7392,N_7532);
nand U8201 (N_8201,N_7358,N_7594);
or U8202 (N_8202,N_7429,N_7864);
and U8203 (N_8203,N_7531,N_7346);
or U8204 (N_8204,N_7827,N_7351);
or U8205 (N_8205,N_7284,N_7308);
or U8206 (N_8206,N_7404,N_7639);
or U8207 (N_8207,N_7658,N_7316);
and U8208 (N_8208,N_7693,N_7498);
and U8209 (N_8209,N_7792,N_7342);
nand U8210 (N_8210,N_7519,N_7516);
nand U8211 (N_8211,N_7551,N_7721);
nand U8212 (N_8212,N_7727,N_7645);
nor U8213 (N_8213,N_7674,N_7471);
or U8214 (N_8214,N_7873,N_7453);
or U8215 (N_8215,N_7496,N_7258);
nor U8216 (N_8216,N_7422,N_7396);
and U8217 (N_8217,N_7253,N_7760);
or U8218 (N_8218,N_7355,N_7264);
or U8219 (N_8219,N_7922,N_7512);
nand U8220 (N_8220,N_7426,N_7886);
nor U8221 (N_8221,N_7401,N_7859);
nand U8222 (N_8222,N_7828,N_7636);
nand U8223 (N_8223,N_7572,N_7559);
or U8224 (N_8224,N_7446,N_7748);
nand U8225 (N_8225,N_7663,N_7726);
nor U8226 (N_8226,N_7755,N_7339);
and U8227 (N_8227,N_7895,N_7836);
nand U8228 (N_8228,N_7522,N_7901);
and U8229 (N_8229,N_7617,N_7439);
and U8230 (N_8230,N_7634,N_7652);
and U8231 (N_8231,N_7667,N_7285);
nand U8232 (N_8232,N_7746,N_7470);
nor U8233 (N_8233,N_7211,N_7924);
or U8234 (N_8234,N_7731,N_7365);
and U8235 (N_8235,N_7443,N_7970);
nand U8236 (N_8236,N_7630,N_7973);
nand U8237 (N_8237,N_7776,N_7811);
nor U8238 (N_8238,N_7867,N_7813);
nand U8239 (N_8239,N_7935,N_7580);
nor U8240 (N_8240,N_7670,N_7281);
nand U8241 (N_8241,N_7203,N_7356);
or U8242 (N_8242,N_7390,N_7900);
or U8243 (N_8243,N_7244,N_7820);
and U8244 (N_8244,N_7961,N_7706);
nand U8245 (N_8245,N_7337,N_7419);
nand U8246 (N_8246,N_7743,N_7633);
or U8247 (N_8247,N_7298,N_7785);
nor U8248 (N_8248,N_7983,N_7228);
or U8249 (N_8249,N_7488,N_7798);
or U8250 (N_8250,N_7407,N_7681);
nor U8251 (N_8251,N_7826,N_7360);
and U8252 (N_8252,N_7751,N_7972);
nor U8253 (N_8253,N_7724,N_7320);
nand U8254 (N_8254,N_7381,N_7840);
or U8255 (N_8255,N_7234,N_7694);
and U8256 (N_8256,N_7592,N_7990);
nor U8257 (N_8257,N_7230,N_7566);
nand U8258 (N_8258,N_7382,N_7807);
and U8259 (N_8259,N_7290,N_7801);
nand U8260 (N_8260,N_7430,N_7625);
and U8261 (N_8261,N_7989,N_7556);
xnor U8262 (N_8262,N_7481,N_7371);
or U8263 (N_8263,N_7441,N_7644);
nand U8264 (N_8264,N_7929,N_7328);
and U8265 (N_8265,N_7480,N_7986);
or U8266 (N_8266,N_7870,N_7740);
or U8267 (N_8267,N_7528,N_7679);
nand U8268 (N_8268,N_7237,N_7403);
and U8269 (N_8269,N_7898,N_7717);
and U8270 (N_8270,N_7857,N_7438);
or U8271 (N_8271,N_7330,N_7712);
nor U8272 (N_8272,N_7389,N_7465);
or U8273 (N_8273,N_7491,N_7741);
or U8274 (N_8274,N_7908,N_7621);
nor U8275 (N_8275,N_7276,N_7609);
nand U8276 (N_8276,N_7853,N_7845);
and U8277 (N_8277,N_7554,N_7831);
or U8278 (N_8278,N_7541,N_7366);
nor U8279 (N_8279,N_7278,N_7321);
nand U8280 (N_8280,N_7589,N_7367);
and U8281 (N_8281,N_7893,N_7501);
and U8282 (N_8282,N_7560,N_7816);
and U8283 (N_8283,N_7225,N_7974);
nand U8284 (N_8284,N_7207,N_7608);
nand U8285 (N_8285,N_7200,N_7931);
or U8286 (N_8286,N_7641,N_7201);
nor U8287 (N_8287,N_7361,N_7306);
nand U8288 (N_8288,N_7466,N_7739);
and U8289 (N_8289,N_7844,N_7686);
nor U8290 (N_8290,N_7647,N_7705);
or U8291 (N_8291,N_7557,N_7752);
and U8292 (N_8292,N_7311,N_7800);
or U8293 (N_8293,N_7771,N_7500);
or U8294 (N_8294,N_7246,N_7267);
or U8295 (N_8295,N_7700,N_7575);
nor U8296 (N_8296,N_7368,N_7780);
nor U8297 (N_8297,N_7662,N_7469);
xnor U8298 (N_8298,N_7269,N_7432);
or U8299 (N_8299,N_7472,N_7379);
nand U8300 (N_8300,N_7680,N_7363);
nand U8301 (N_8301,N_7725,N_7370);
nand U8302 (N_8302,N_7655,N_7948);
nand U8303 (N_8303,N_7412,N_7690);
or U8304 (N_8304,N_7352,N_7325);
nand U8305 (N_8305,N_7937,N_7909);
nor U8306 (N_8306,N_7265,N_7449);
nand U8307 (N_8307,N_7703,N_7214);
and U8308 (N_8308,N_7310,N_7791);
nor U8309 (N_8309,N_7482,N_7605);
nand U8310 (N_8310,N_7835,N_7305);
nand U8311 (N_8311,N_7564,N_7242);
nand U8312 (N_8312,N_7335,N_7261);
nand U8313 (N_8313,N_7623,N_7292);
nor U8314 (N_8314,N_7247,N_7927);
nand U8315 (N_8315,N_7562,N_7333);
nand U8316 (N_8316,N_7995,N_7947);
nor U8317 (N_8317,N_7327,N_7959);
nor U8318 (N_8318,N_7266,N_7664);
nor U8319 (N_8319,N_7326,N_7395);
and U8320 (N_8320,N_7224,N_7941);
and U8321 (N_8321,N_7632,N_7918);
and U8322 (N_8322,N_7688,N_7863);
or U8323 (N_8323,N_7398,N_7710);
nand U8324 (N_8324,N_7839,N_7212);
nor U8325 (N_8325,N_7945,N_7232);
or U8326 (N_8326,N_7263,N_7587);
nor U8327 (N_8327,N_7455,N_7868);
and U8328 (N_8328,N_7669,N_7599);
and U8329 (N_8329,N_7861,N_7955);
or U8330 (N_8330,N_7631,N_7782);
or U8331 (N_8331,N_7876,N_7359);
or U8332 (N_8332,N_7968,N_7431);
or U8333 (N_8333,N_7969,N_7967);
nor U8334 (N_8334,N_7837,N_7665);
or U8335 (N_8335,N_7975,N_7387);
nor U8336 (N_8336,N_7277,N_7750);
nand U8337 (N_8337,N_7241,N_7943);
nor U8338 (N_8338,N_7730,N_7819);
nand U8339 (N_8339,N_7349,N_7374);
nand U8340 (N_8340,N_7877,N_7369);
nand U8341 (N_8341,N_7525,N_7765);
nand U8342 (N_8342,N_7576,N_7408);
and U8343 (N_8343,N_7932,N_7235);
and U8344 (N_8344,N_7492,N_7565);
nor U8345 (N_8345,N_7993,N_7783);
nand U8346 (N_8346,N_7477,N_7815);
nand U8347 (N_8347,N_7208,N_7444);
or U8348 (N_8348,N_7841,N_7862);
or U8349 (N_8349,N_7354,N_7373);
nand U8350 (N_8350,N_7417,N_7851);
and U8351 (N_8351,N_7424,N_7274);
nand U8352 (N_8352,N_7406,N_7823);
nor U8353 (N_8353,N_7651,N_7903);
or U8354 (N_8354,N_7952,N_7604);
or U8355 (N_8355,N_7759,N_7892);
and U8356 (N_8356,N_7745,N_7956);
and U8357 (N_8357,N_7493,N_7643);
or U8358 (N_8358,N_7574,N_7460);
and U8359 (N_8359,N_7484,N_7938);
and U8360 (N_8360,N_7788,N_7540);
and U8361 (N_8361,N_7685,N_7796);
or U8362 (N_8362,N_7294,N_7344);
nand U8363 (N_8363,N_7552,N_7921);
nor U8364 (N_8364,N_7513,N_7618);
nor U8365 (N_8365,N_7822,N_7695);
or U8366 (N_8366,N_7885,N_7936);
nor U8367 (N_8367,N_7509,N_7303);
and U8368 (N_8368,N_7926,N_7527);
or U8369 (N_8369,N_7902,N_7596);
nand U8370 (N_8370,N_7978,N_7991);
nand U8371 (N_8371,N_7964,N_7980);
nand U8372 (N_8372,N_7450,N_7579);
and U8373 (N_8373,N_7503,N_7606);
or U8374 (N_8374,N_7534,N_7619);
nor U8375 (N_8375,N_7958,N_7635);
or U8376 (N_8376,N_7736,N_7231);
nand U8377 (N_8377,N_7648,N_7570);
and U8378 (N_8378,N_7982,N_7571);
or U8379 (N_8379,N_7627,N_7388);
or U8380 (N_8380,N_7542,N_7558);
or U8381 (N_8381,N_7338,N_7229);
nor U8382 (N_8382,N_7874,N_7949);
and U8383 (N_8383,N_7479,N_7708);
nand U8384 (N_8384,N_7923,N_7928);
and U8385 (N_8385,N_7485,N_7939);
nor U8386 (N_8386,N_7259,N_7729);
and U8387 (N_8387,N_7539,N_7507);
nor U8388 (N_8388,N_7824,N_7805);
or U8389 (N_8389,N_7468,N_7312);
and U8390 (N_8390,N_7781,N_7654);
nor U8391 (N_8391,N_7784,N_7256);
or U8392 (N_8392,N_7456,N_7769);
and U8393 (N_8393,N_7307,N_7590);
nor U8394 (N_8394,N_7459,N_7291);
nand U8395 (N_8395,N_7637,N_7723);
nand U8396 (N_8396,N_7987,N_7976);
nor U8397 (N_8397,N_7535,N_7950);
nor U8398 (N_8398,N_7865,N_7436);
nand U8399 (N_8399,N_7770,N_7607);
nand U8400 (N_8400,N_7920,N_7644);
or U8401 (N_8401,N_7510,N_7632);
nand U8402 (N_8402,N_7852,N_7768);
nor U8403 (N_8403,N_7381,N_7750);
and U8404 (N_8404,N_7702,N_7569);
nand U8405 (N_8405,N_7588,N_7212);
xor U8406 (N_8406,N_7767,N_7734);
or U8407 (N_8407,N_7953,N_7923);
nor U8408 (N_8408,N_7572,N_7856);
or U8409 (N_8409,N_7904,N_7686);
nor U8410 (N_8410,N_7895,N_7882);
nand U8411 (N_8411,N_7699,N_7601);
nor U8412 (N_8412,N_7326,N_7409);
or U8413 (N_8413,N_7951,N_7469);
nand U8414 (N_8414,N_7259,N_7882);
nor U8415 (N_8415,N_7965,N_7427);
nor U8416 (N_8416,N_7573,N_7710);
or U8417 (N_8417,N_7785,N_7569);
or U8418 (N_8418,N_7349,N_7994);
nor U8419 (N_8419,N_7425,N_7344);
and U8420 (N_8420,N_7674,N_7501);
nor U8421 (N_8421,N_7924,N_7756);
and U8422 (N_8422,N_7933,N_7841);
nand U8423 (N_8423,N_7454,N_7672);
nor U8424 (N_8424,N_7580,N_7855);
or U8425 (N_8425,N_7424,N_7866);
nor U8426 (N_8426,N_7212,N_7875);
or U8427 (N_8427,N_7790,N_7960);
nand U8428 (N_8428,N_7915,N_7949);
nand U8429 (N_8429,N_7412,N_7578);
nand U8430 (N_8430,N_7991,N_7225);
and U8431 (N_8431,N_7494,N_7243);
nor U8432 (N_8432,N_7233,N_7932);
and U8433 (N_8433,N_7899,N_7703);
and U8434 (N_8434,N_7809,N_7660);
nand U8435 (N_8435,N_7262,N_7794);
nor U8436 (N_8436,N_7788,N_7375);
nand U8437 (N_8437,N_7397,N_7790);
and U8438 (N_8438,N_7999,N_7549);
nand U8439 (N_8439,N_7905,N_7210);
or U8440 (N_8440,N_7630,N_7510);
or U8441 (N_8441,N_7896,N_7687);
nand U8442 (N_8442,N_7348,N_7340);
nand U8443 (N_8443,N_7875,N_7987);
and U8444 (N_8444,N_7771,N_7425);
nor U8445 (N_8445,N_7351,N_7255);
nand U8446 (N_8446,N_7987,N_7884);
and U8447 (N_8447,N_7443,N_7593);
and U8448 (N_8448,N_7996,N_7371);
or U8449 (N_8449,N_7201,N_7448);
or U8450 (N_8450,N_7448,N_7776);
nand U8451 (N_8451,N_7506,N_7501);
nand U8452 (N_8452,N_7272,N_7480);
nor U8453 (N_8453,N_7977,N_7721);
nor U8454 (N_8454,N_7699,N_7435);
nor U8455 (N_8455,N_7573,N_7538);
nand U8456 (N_8456,N_7269,N_7741);
and U8457 (N_8457,N_7906,N_7234);
nor U8458 (N_8458,N_7417,N_7734);
nand U8459 (N_8459,N_7291,N_7259);
nand U8460 (N_8460,N_7314,N_7328);
or U8461 (N_8461,N_7570,N_7906);
and U8462 (N_8462,N_7720,N_7815);
and U8463 (N_8463,N_7268,N_7917);
and U8464 (N_8464,N_7731,N_7209);
nand U8465 (N_8465,N_7702,N_7397);
nor U8466 (N_8466,N_7575,N_7593);
nor U8467 (N_8467,N_7681,N_7471);
nand U8468 (N_8468,N_7219,N_7752);
nand U8469 (N_8469,N_7523,N_7915);
nand U8470 (N_8470,N_7885,N_7368);
nor U8471 (N_8471,N_7878,N_7805);
nor U8472 (N_8472,N_7528,N_7471);
nand U8473 (N_8473,N_7585,N_7307);
or U8474 (N_8474,N_7752,N_7425);
or U8475 (N_8475,N_7510,N_7394);
nand U8476 (N_8476,N_7355,N_7790);
nor U8477 (N_8477,N_7683,N_7338);
nand U8478 (N_8478,N_7431,N_7534);
nand U8479 (N_8479,N_7989,N_7979);
nor U8480 (N_8480,N_7556,N_7760);
nand U8481 (N_8481,N_7889,N_7838);
nor U8482 (N_8482,N_7922,N_7218);
nor U8483 (N_8483,N_7292,N_7279);
nand U8484 (N_8484,N_7635,N_7324);
nor U8485 (N_8485,N_7367,N_7809);
or U8486 (N_8486,N_7235,N_7909);
or U8487 (N_8487,N_7762,N_7771);
and U8488 (N_8488,N_7218,N_7677);
nor U8489 (N_8489,N_7507,N_7421);
nor U8490 (N_8490,N_7985,N_7697);
or U8491 (N_8491,N_7603,N_7434);
nand U8492 (N_8492,N_7685,N_7563);
xor U8493 (N_8493,N_7399,N_7913);
nand U8494 (N_8494,N_7293,N_7753);
nand U8495 (N_8495,N_7489,N_7566);
nand U8496 (N_8496,N_7837,N_7993);
or U8497 (N_8497,N_7984,N_7831);
or U8498 (N_8498,N_7915,N_7356);
and U8499 (N_8499,N_7299,N_7490);
nand U8500 (N_8500,N_7729,N_7781);
nor U8501 (N_8501,N_7958,N_7993);
or U8502 (N_8502,N_7577,N_7985);
and U8503 (N_8503,N_7534,N_7683);
nor U8504 (N_8504,N_7362,N_7386);
nor U8505 (N_8505,N_7857,N_7701);
or U8506 (N_8506,N_7443,N_7633);
nand U8507 (N_8507,N_7616,N_7521);
and U8508 (N_8508,N_7867,N_7686);
or U8509 (N_8509,N_7742,N_7296);
and U8510 (N_8510,N_7218,N_7529);
or U8511 (N_8511,N_7894,N_7943);
nor U8512 (N_8512,N_7243,N_7358);
and U8513 (N_8513,N_7883,N_7774);
nand U8514 (N_8514,N_7841,N_7310);
nor U8515 (N_8515,N_7413,N_7906);
nor U8516 (N_8516,N_7725,N_7301);
xor U8517 (N_8517,N_7945,N_7345);
and U8518 (N_8518,N_7787,N_7829);
or U8519 (N_8519,N_7509,N_7257);
nand U8520 (N_8520,N_7386,N_7890);
and U8521 (N_8521,N_7511,N_7955);
nand U8522 (N_8522,N_7800,N_7462);
and U8523 (N_8523,N_7632,N_7968);
nor U8524 (N_8524,N_7934,N_7639);
or U8525 (N_8525,N_7464,N_7544);
and U8526 (N_8526,N_7214,N_7353);
nor U8527 (N_8527,N_7562,N_7809);
or U8528 (N_8528,N_7276,N_7971);
and U8529 (N_8529,N_7927,N_7556);
nor U8530 (N_8530,N_7399,N_7409);
nor U8531 (N_8531,N_7978,N_7922);
or U8532 (N_8532,N_7879,N_7572);
nor U8533 (N_8533,N_7649,N_7297);
nand U8534 (N_8534,N_7615,N_7422);
nor U8535 (N_8535,N_7916,N_7292);
nor U8536 (N_8536,N_7911,N_7396);
nor U8537 (N_8537,N_7883,N_7253);
and U8538 (N_8538,N_7893,N_7464);
nor U8539 (N_8539,N_7978,N_7918);
nor U8540 (N_8540,N_7740,N_7856);
nor U8541 (N_8541,N_7296,N_7597);
nand U8542 (N_8542,N_7337,N_7346);
nor U8543 (N_8543,N_7693,N_7898);
or U8544 (N_8544,N_7536,N_7982);
nand U8545 (N_8545,N_7501,N_7204);
nand U8546 (N_8546,N_7400,N_7648);
and U8547 (N_8547,N_7959,N_7832);
nor U8548 (N_8548,N_7515,N_7934);
or U8549 (N_8549,N_7452,N_7469);
nand U8550 (N_8550,N_7233,N_7323);
nand U8551 (N_8551,N_7790,N_7938);
nor U8552 (N_8552,N_7780,N_7988);
nand U8553 (N_8553,N_7770,N_7921);
nor U8554 (N_8554,N_7794,N_7757);
nor U8555 (N_8555,N_7862,N_7581);
or U8556 (N_8556,N_7249,N_7501);
or U8557 (N_8557,N_7262,N_7953);
and U8558 (N_8558,N_7299,N_7600);
and U8559 (N_8559,N_7455,N_7878);
nand U8560 (N_8560,N_7916,N_7707);
xor U8561 (N_8561,N_7496,N_7311);
nor U8562 (N_8562,N_7466,N_7821);
or U8563 (N_8563,N_7447,N_7989);
and U8564 (N_8564,N_7890,N_7402);
nor U8565 (N_8565,N_7619,N_7819);
nor U8566 (N_8566,N_7759,N_7980);
and U8567 (N_8567,N_7477,N_7840);
or U8568 (N_8568,N_7410,N_7525);
nor U8569 (N_8569,N_7227,N_7762);
nor U8570 (N_8570,N_7754,N_7682);
or U8571 (N_8571,N_7585,N_7328);
and U8572 (N_8572,N_7842,N_7380);
nand U8573 (N_8573,N_7398,N_7925);
or U8574 (N_8574,N_7424,N_7457);
xnor U8575 (N_8575,N_7728,N_7660);
nand U8576 (N_8576,N_7339,N_7456);
and U8577 (N_8577,N_7472,N_7200);
nor U8578 (N_8578,N_7763,N_7724);
xor U8579 (N_8579,N_7304,N_7342);
and U8580 (N_8580,N_7855,N_7819);
nor U8581 (N_8581,N_7930,N_7453);
or U8582 (N_8582,N_7345,N_7795);
nand U8583 (N_8583,N_7227,N_7445);
or U8584 (N_8584,N_7388,N_7888);
nor U8585 (N_8585,N_7679,N_7422);
and U8586 (N_8586,N_7392,N_7818);
and U8587 (N_8587,N_7521,N_7325);
nand U8588 (N_8588,N_7799,N_7638);
and U8589 (N_8589,N_7531,N_7711);
or U8590 (N_8590,N_7546,N_7312);
or U8591 (N_8591,N_7922,N_7327);
nand U8592 (N_8592,N_7226,N_7837);
nor U8593 (N_8593,N_7604,N_7462);
nand U8594 (N_8594,N_7429,N_7327);
or U8595 (N_8595,N_7457,N_7890);
and U8596 (N_8596,N_7264,N_7353);
and U8597 (N_8597,N_7548,N_7231);
or U8598 (N_8598,N_7774,N_7682);
nand U8599 (N_8599,N_7857,N_7435);
nand U8600 (N_8600,N_7640,N_7956);
and U8601 (N_8601,N_7371,N_7414);
or U8602 (N_8602,N_7761,N_7250);
and U8603 (N_8603,N_7795,N_7454);
nand U8604 (N_8604,N_7757,N_7222);
nor U8605 (N_8605,N_7512,N_7779);
nor U8606 (N_8606,N_7938,N_7475);
or U8607 (N_8607,N_7240,N_7747);
nor U8608 (N_8608,N_7443,N_7791);
nor U8609 (N_8609,N_7200,N_7408);
nand U8610 (N_8610,N_7678,N_7337);
nor U8611 (N_8611,N_7536,N_7397);
or U8612 (N_8612,N_7696,N_7930);
and U8613 (N_8613,N_7341,N_7994);
and U8614 (N_8614,N_7975,N_7860);
and U8615 (N_8615,N_7932,N_7663);
nor U8616 (N_8616,N_7304,N_7622);
and U8617 (N_8617,N_7850,N_7412);
and U8618 (N_8618,N_7808,N_7498);
or U8619 (N_8619,N_7222,N_7607);
nor U8620 (N_8620,N_7696,N_7502);
or U8621 (N_8621,N_7720,N_7812);
nand U8622 (N_8622,N_7970,N_7437);
nand U8623 (N_8623,N_7567,N_7497);
and U8624 (N_8624,N_7754,N_7624);
nand U8625 (N_8625,N_7312,N_7297);
nand U8626 (N_8626,N_7933,N_7362);
or U8627 (N_8627,N_7325,N_7876);
or U8628 (N_8628,N_7678,N_7972);
and U8629 (N_8629,N_7871,N_7974);
or U8630 (N_8630,N_7847,N_7417);
and U8631 (N_8631,N_7539,N_7804);
nand U8632 (N_8632,N_7927,N_7233);
or U8633 (N_8633,N_7267,N_7491);
nand U8634 (N_8634,N_7850,N_7891);
or U8635 (N_8635,N_7923,N_7680);
or U8636 (N_8636,N_7921,N_7480);
and U8637 (N_8637,N_7995,N_7929);
or U8638 (N_8638,N_7390,N_7829);
and U8639 (N_8639,N_7259,N_7956);
or U8640 (N_8640,N_7429,N_7775);
or U8641 (N_8641,N_7579,N_7386);
or U8642 (N_8642,N_7954,N_7275);
nor U8643 (N_8643,N_7508,N_7530);
nand U8644 (N_8644,N_7735,N_7342);
nor U8645 (N_8645,N_7598,N_7576);
nor U8646 (N_8646,N_7318,N_7397);
nor U8647 (N_8647,N_7331,N_7444);
nand U8648 (N_8648,N_7350,N_7867);
nand U8649 (N_8649,N_7610,N_7680);
nor U8650 (N_8650,N_7520,N_7295);
nor U8651 (N_8651,N_7340,N_7231);
nand U8652 (N_8652,N_7580,N_7236);
and U8653 (N_8653,N_7970,N_7346);
or U8654 (N_8654,N_7826,N_7252);
or U8655 (N_8655,N_7582,N_7231);
or U8656 (N_8656,N_7935,N_7524);
xnor U8657 (N_8657,N_7803,N_7518);
and U8658 (N_8658,N_7742,N_7536);
or U8659 (N_8659,N_7219,N_7973);
or U8660 (N_8660,N_7579,N_7841);
or U8661 (N_8661,N_7301,N_7248);
nand U8662 (N_8662,N_7322,N_7879);
nand U8663 (N_8663,N_7887,N_7696);
xor U8664 (N_8664,N_7827,N_7684);
nor U8665 (N_8665,N_7282,N_7503);
and U8666 (N_8666,N_7296,N_7723);
nor U8667 (N_8667,N_7973,N_7492);
or U8668 (N_8668,N_7350,N_7236);
or U8669 (N_8669,N_7449,N_7947);
nor U8670 (N_8670,N_7241,N_7543);
and U8671 (N_8671,N_7693,N_7723);
nand U8672 (N_8672,N_7673,N_7368);
or U8673 (N_8673,N_7669,N_7638);
or U8674 (N_8674,N_7793,N_7672);
and U8675 (N_8675,N_7529,N_7397);
xor U8676 (N_8676,N_7412,N_7693);
nand U8677 (N_8677,N_7553,N_7728);
nor U8678 (N_8678,N_7922,N_7726);
and U8679 (N_8679,N_7866,N_7735);
and U8680 (N_8680,N_7771,N_7263);
nor U8681 (N_8681,N_7588,N_7303);
nand U8682 (N_8682,N_7456,N_7204);
nor U8683 (N_8683,N_7746,N_7691);
nor U8684 (N_8684,N_7763,N_7634);
and U8685 (N_8685,N_7840,N_7357);
nor U8686 (N_8686,N_7468,N_7216);
nor U8687 (N_8687,N_7904,N_7275);
or U8688 (N_8688,N_7504,N_7689);
and U8689 (N_8689,N_7347,N_7884);
nand U8690 (N_8690,N_7238,N_7591);
nand U8691 (N_8691,N_7777,N_7487);
nand U8692 (N_8692,N_7933,N_7524);
nand U8693 (N_8693,N_7247,N_7597);
nor U8694 (N_8694,N_7279,N_7935);
and U8695 (N_8695,N_7988,N_7415);
nor U8696 (N_8696,N_7398,N_7797);
and U8697 (N_8697,N_7400,N_7640);
nor U8698 (N_8698,N_7417,N_7415);
or U8699 (N_8699,N_7772,N_7279);
and U8700 (N_8700,N_7266,N_7919);
nor U8701 (N_8701,N_7852,N_7759);
nor U8702 (N_8702,N_7257,N_7868);
nor U8703 (N_8703,N_7312,N_7307);
nand U8704 (N_8704,N_7504,N_7528);
xnor U8705 (N_8705,N_7382,N_7594);
nor U8706 (N_8706,N_7557,N_7953);
xor U8707 (N_8707,N_7324,N_7248);
or U8708 (N_8708,N_7696,N_7253);
and U8709 (N_8709,N_7218,N_7956);
or U8710 (N_8710,N_7438,N_7534);
or U8711 (N_8711,N_7997,N_7531);
and U8712 (N_8712,N_7218,N_7537);
nand U8713 (N_8713,N_7963,N_7811);
and U8714 (N_8714,N_7792,N_7756);
and U8715 (N_8715,N_7370,N_7213);
nor U8716 (N_8716,N_7705,N_7946);
nor U8717 (N_8717,N_7744,N_7225);
and U8718 (N_8718,N_7265,N_7674);
nor U8719 (N_8719,N_7558,N_7480);
and U8720 (N_8720,N_7923,N_7705);
or U8721 (N_8721,N_7250,N_7733);
nand U8722 (N_8722,N_7862,N_7911);
nor U8723 (N_8723,N_7900,N_7682);
nor U8724 (N_8724,N_7827,N_7990);
nor U8725 (N_8725,N_7550,N_7270);
or U8726 (N_8726,N_7328,N_7709);
and U8727 (N_8727,N_7289,N_7756);
nor U8728 (N_8728,N_7630,N_7656);
and U8729 (N_8729,N_7692,N_7633);
nand U8730 (N_8730,N_7821,N_7219);
or U8731 (N_8731,N_7347,N_7290);
nand U8732 (N_8732,N_7296,N_7609);
and U8733 (N_8733,N_7841,N_7831);
nand U8734 (N_8734,N_7468,N_7203);
nor U8735 (N_8735,N_7387,N_7822);
or U8736 (N_8736,N_7825,N_7870);
and U8737 (N_8737,N_7709,N_7982);
nor U8738 (N_8738,N_7937,N_7510);
and U8739 (N_8739,N_7949,N_7478);
or U8740 (N_8740,N_7434,N_7775);
nand U8741 (N_8741,N_7798,N_7735);
nand U8742 (N_8742,N_7521,N_7675);
and U8743 (N_8743,N_7639,N_7518);
and U8744 (N_8744,N_7248,N_7755);
nand U8745 (N_8745,N_7606,N_7315);
and U8746 (N_8746,N_7411,N_7619);
and U8747 (N_8747,N_7680,N_7919);
nor U8748 (N_8748,N_7914,N_7944);
or U8749 (N_8749,N_7392,N_7810);
or U8750 (N_8750,N_7871,N_7263);
and U8751 (N_8751,N_7860,N_7519);
nand U8752 (N_8752,N_7805,N_7360);
and U8753 (N_8753,N_7677,N_7734);
nor U8754 (N_8754,N_7220,N_7516);
nor U8755 (N_8755,N_7880,N_7592);
and U8756 (N_8756,N_7630,N_7696);
and U8757 (N_8757,N_7586,N_7423);
and U8758 (N_8758,N_7748,N_7584);
nor U8759 (N_8759,N_7860,N_7651);
nand U8760 (N_8760,N_7991,N_7268);
nor U8761 (N_8761,N_7444,N_7323);
and U8762 (N_8762,N_7379,N_7605);
nor U8763 (N_8763,N_7963,N_7258);
and U8764 (N_8764,N_7873,N_7201);
or U8765 (N_8765,N_7385,N_7352);
or U8766 (N_8766,N_7630,N_7769);
or U8767 (N_8767,N_7850,N_7730);
nand U8768 (N_8768,N_7928,N_7806);
or U8769 (N_8769,N_7701,N_7346);
nor U8770 (N_8770,N_7311,N_7418);
nor U8771 (N_8771,N_7335,N_7792);
and U8772 (N_8772,N_7692,N_7554);
nor U8773 (N_8773,N_7343,N_7819);
or U8774 (N_8774,N_7643,N_7766);
nor U8775 (N_8775,N_7539,N_7814);
nor U8776 (N_8776,N_7651,N_7570);
nor U8777 (N_8777,N_7459,N_7486);
or U8778 (N_8778,N_7412,N_7798);
or U8779 (N_8779,N_7647,N_7736);
or U8780 (N_8780,N_7771,N_7811);
nand U8781 (N_8781,N_7226,N_7256);
nand U8782 (N_8782,N_7991,N_7364);
and U8783 (N_8783,N_7972,N_7880);
or U8784 (N_8784,N_7865,N_7262);
or U8785 (N_8785,N_7782,N_7860);
and U8786 (N_8786,N_7666,N_7945);
and U8787 (N_8787,N_7678,N_7255);
or U8788 (N_8788,N_7479,N_7429);
and U8789 (N_8789,N_7577,N_7903);
nor U8790 (N_8790,N_7656,N_7490);
or U8791 (N_8791,N_7780,N_7998);
nor U8792 (N_8792,N_7941,N_7612);
nand U8793 (N_8793,N_7742,N_7315);
and U8794 (N_8794,N_7873,N_7425);
or U8795 (N_8795,N_7770,N_7564);
nor U8796 (N_8796,N_7937,N_7806);
or U8797 (N_8797,N_7655,N_7923);
nand U8798 (N_8798,N_7693,N_7293);
and U8799 (N_8799,N_7907,N_7863);
and U8800 (N_8800,N_8494,N_8362);
nor U8801 (N_8801,N_8190,N_8519);
nand U8802 (N_8802,N_8194,N_8315);
nor U8803 (N_8803,N_8600,N_8500);
nand U8804 (N_8804,N_8419,N_8025);
nor U8805 (N_8805,N_8654,N_8692);
nor U8806 (N_8806,N_8254,N_8711);
nor U8807 (N_8807,N_8133,N_8742);
and U8808 (N_8808,N_8082,N_8202);
nand U8809 (N_8809,N_8203,N_8771);
nand U8810 (N_8810,N_8287,N_8180);
nand U8811 (N_8811,N_8166,N_8724);
nor U8812 (N_8812,N_8551,N_8571);
nand U8813 (N_8813,N_8770,N_8776);
nand U8814 (N_8814,N_8212,N_8487);
xnor U8815 (N_8815,N_8642,N_8789);
and U8816 (N_8816,N_8554,N_8356);
or U8817 (N_8817,N_8174,N_8624);
nand U8818 (N_8818,N_8709,N_8060);
or U8819 (N_8819,N_8697,N_8428);
or U8820 (N_8820,N_8630,N_8491);
nor U8821 (N_8821,N_8458,N_8327);
or U8822 (N_8822,N_8633,N_8220);
and U8823 (N_8823,N_8700,N_8601);
nand U8824 (N_8824,N_8745,N_8749);
nor U8825 (N_8825,N_8499,N_8373);
or U8826 (N_8826,N_8207,N_8296);
or U8827 (N_8827,N_8597,N_8088);
or U8828 (N_8828,N_8734,N_8334);
nand U8829 (N_8829,N_8086,N_8696);
or U8830 (N_8830,N_8503,N_8191);
nor U8831 (N_8831,N_8038,N_8434);
nor U8832 (N_8832,N_8609,N_8274);
or U8833 (N_8833,N_8092,N_8483);
and U8834 (N_8834,N_8746,N_8364);
and U8835 (N_8835,N_8567,N_8306);
nor U8836 (N_8836,N_8637,N_8035);
nor U8837 (N_8837,N_8537,N_8055);
nor U8838 (N_8838,N_8073,N_8546);
nor U8839 (N_8839,N_8393,N_8098);
nand U8840 (N_8840,N_8549,N_8723);
nor U8841 (N_8841,N_8534,N_8740);
or U8842 (N_8842,N_8782,N_8318);
nor U8843 (N_8843,N_8079,N_8282);
nor U8844 (N_8844,N_8460,N_8009);
and U8845 (N_8845,N_8602,N_8784);
nand U8846 (N_8846,N_8096,N_8730);
nand U8847 (N_8847,N_8233,N_8752);
nand U8848 (N_8848,N_8538,N_8014);
or U8849 (N_8849,N_8648,N_8525);
or U8850 (N_8850,N_8066,N_8210);
or U8851 (N_8851,N_8056,N_8660);
and U8852 (N_8852,N_8214,N_8104);
and U8853 (N_8853,N_8024,N_8384);
and U8854 (N_8854,N_8337,N_8271);
nor U8855 (N_8855,N_8012,N_8382);
nor U8856 (N_8856,N_8061,N_8018);
nor U8857 (N_8857,N_8644,N_8392);
nor U8858 (N_8858,N_8559,N_8015);
nand U8859 (N_8859,N_8495,N_8578);
nor U8860 (N_8860,N_8251,N_8353);
and U8861 (N_8861,N_8020,N_8293);
nand U8862 (N_8862,N_8052,N_8478);
and U8863 (N_8863,N_8177,N_8216);
and U8864 (N_8864,N_8276,N_8385);
and U8865 (N_8865,N_8266,N_8242);
nand U8866 (N_8866,N_8744,N_8599);
nand U8867 (N_8867,N_8189,N_8129);
and U8868 (N_8868,N_8774,N_8143);
and U8869 (N_8869,N_8112,N_8232);
nor U8870 (N_8870,N_8077,N_8585);
nor U8871 (N_8871,N_8181,N_8464);
or U8872 (N_8872,N_8344,N_8107);
and U8873 (N_8873,N_8057,N_8629);
nand U8874 (N_8874,N_8354,N_8026);
nor U8875 (N_8875,N_8046,N_8389);
nor U8876 (N_8876,N_8374,N_8037);
and U8877 (N_8877,N_8173,N_8146);
and U8878 (N_8878,N_8067,N_8442);
nor U8879 (N_8879,N_8611,N_8272);
and U8880 (N_8880,N_8668,N_8245);
or U8881 (N_8881,N_8335,N_8726);
and U8882 (N_8882,N_8369,N_8105);
nor U8883 (N_8883,N_8345,N_8541);
nand U8884 (N_8884,N_8323,N_8408);
and U8885 (N_8885,N_8175,N_8050);
nor U8886 (N_8886,N_8339,N_8607);
nor U8887 (N_8887,N_8307,N_8250);
or U8888 (N_8888,N_8132,N_8623);
nor U8889 (N_8889,N_8006,N_8403);
nor U8890 (N_8890,N_8205,N_8610);
and U8891 (N_8891,N_8252,N_8118);
nor U8892 (N_8892,N_8002,N_8729);
nor U8893 (N_8893,N_8506,N_8244);
and U8894 (N_8894,N_8379,N_8588);
nand U8895 (N_8895,N_8168,N_8156);
nor U8896 (N_8896,N_8511,N_8613);
and U8897 (N_8897,N_8063,N_8147);
and U8898 (N_8898,N_8439,N_8301);
or U8899 (N_8899,N_8663,N_8225);
nor U8900 (N_8900,N_8005,N_8000);
or U8901 (N_8901,N_8548,N_8367);
nand U8902 (N_8902,N_8788,N_8594);
nor U8903 (N_8903,N_8447,N_8739);
nor U8904 (N_8904,N_8430,N_8080);
nand U8905 (N_8905,N_8634,N_8192);
and U8906 (N_8906,N_8278,N_8001);
or U8907 (N_8907,N_8641,N_8126);
or U8908 (N_8908,N_8682,N_8703);
and U8909 (N_8909,N_8733,N_8604);
and U8910 (N_8910,N_8451,N_8218);
nor U8911 (N_8911,N_8119,N_8347);
or U8912 (N_8912,N_8671,N_8273);
or U8913 (N_8913,N_8310,N_8256);
or U8914 (N_8914,N_8687,N_8084);
nand U8915 (N_8915,N_8545,N_8440);
nor U8916 (N_8916,N_8110,N_8197);
or U8917 (N_8917,N_8432,N_8477);
nor U8918 (N_8918,N_8170,N_8375);
or U8919 (N_8919,N_8217,N_8198);
and U8920 (N_8920,N_8452,N_8635);
nand U8921 (N_8921,N_8685,N_8593);
or U8922 (N_8922,N_8714,N_8631);
nor U8923 (N_8923,N_8032,N_8155);
or U8924 (N_8924,N_8636,N_8311);
or U8925 (N_8925,N_8275,N_8625);
nand U8926 (N_8926,N_8712,N_8294);
nand U8927 (N_8927,N_8023,N_8200);
nor U8928 (N_8928,N_8341,N_8101);
and U8929 (N_8929,N_8070,N_8386);
nand U8930 (N_8930,N_8680,N_8409);
nand U8931 (N_8931,N_8142,N_8095);
nand U8932 (N_8932,N_8300,N_8580);
and U8933 (N_8933,N_8647,N_8352);
nor U8934 (N_8934,N_8763,N_8078);
or U8935 (N_8935,N_8072,N_8652);
nor U8936 (N_8936,N_8295,N_8003);
nand U8937 (N_8937,N_8441,N_8297);
nor U8938 (N_8938,N_8378,N_8456);
nor U8939 (N_8939,N_8762,N_8532);
nand U8940 (N_8940,N_8258,N_8338);
or U8941 (N_8941,N_8769,N_8484);
nand U8942 (N_8942,N_8526,N_8196);
xnor U8943 (N_8943,N_8397,N_8350);
nor U8944 (N_8944,N_8785,N_8069);
xor U8945 (N_8945,N_8314,N_8667);
or U8946 (N_8946,N_8530,N_8008);
nor U8947 (N_8947,N_8666,N_8372);
nor U8948 (N_8948,N_8791,N_8033);
and U8949 (N_8949,N_8411,N_8777);
or U8950 (N_8950,N_8169,N_8482);
nand U8951 (N_8951,N_8120,N_8376);
nor U8952 (N_8952,N_8627,N_8326);
xnor U8953 (N_8953,N_8358,N_8342);
and U8954 (N_8954,N_8231,N_8405);
or U8955 (N_8955,N_8480,N_8677);
or U8956 (N_8956,N_8649,N_8329);
and U8957 (N_8957,N_8431,N_8725);
nand U8958 (N_8958,N_8330,N_8626);
nand U8959 (N_8959,N_8221,N_8423);
nand U8960 (N_8960,N_8579,N_8658);
and U8961 (N_8961,N_8237,N_8185);
and U8962 (N_8962,N_8135,N_8363);
nor U8963 (N_8963,N_8662,N_8223);
nand U8964 (N_8964,N_8535,N_8243);
and U8965 (N_8965,N_8400,N_8249);
or U8966 (N_8966,N_8760,N_8034);
or U8967 (N_8967,N_8346,N_8312);
nor U8968 (N_8968,N_8794,N_8401);
and U8969 (N_8969,N_8407,N_8246);
nand U8970 (N_8970,N_8463,N_8125);
nor U8971 (N_8971,N_8553,N_8113);
and U8972 (N_8972,N_8091,N_8718);
and U8973 (N_8973,N_8508,N_8435);
or U8974 (N_8974,N_8416,N_8473);
or U8975 (N_8975,N_8558,N_8391);
and U8976 (N_8976,N_8238,N_8333);
nor U8977 (N_8977,N_8563,N_8614);
and U8978 (N_8978,N_8292,N_8094);
nor U8979 (N_8979,N_8542,N_8161);
or U8980 (N_8980,N_8121,N_8608);
nand U8981 (N_8981,N_8544,N_8628);
or U8982 (N_8982,N_8475,N_8468);
nand U8983 (N_8983,N_8493,N_8527);
nand U8984 (N_8984,N_8694,N_8158);
nor U8985 (N_8985,N_8565,N_8427);
nand U8986 (N_8986,N_8188,N_8149);
and U8987 (N_8987,N_8474,N_8016);
nor U8988 (N_8988,N_8162,N_8043);
nor U8989 (N_8989,N_8204,N_8320);
nand U8990 (N_8990,N_8615,N_8612);
xor U8991 (N_8991,N_8085,N_8137);
nor U8992 (N_8992,N_8618,N_8042);
nor U8993 (N_8993,N_8236,N_8365);
nand U8994 (N_8994,N_8028,N_8592);
and U8995 (N_8995,N_8390,N_8768);
and U8996 (N_8996,N_8144,N_8065);
and U8997 (N_8997,N_8522,N_8355);
or U8998 (N_8998,N_8587,N_8651);
or U8999 (N_8999,N_8454,N_8574);
and U9000 (N_9000,N_8255,N_8259);
nand U9001 (N_9001,N_8509,N_8076);
nand U9002 (N_9002,N_8022,N_8781);
nand U9003 (N_9003,N_8450,N_8230);
nand U9004 (N_9004,N_8639,N_8581);
nand U9005 (N_9005,N_8313,N_8701);
and U9006 (N_9006,N_8179,N_8199);
and U9007 (N_9007,N_8343,N_8029);
nor U9008 (N_9008,N_8036,N_8279);
or U9009 (N_9009,N_8524,N_8239);
nand U9010 (N_9010,N_8523,N_8455);
nand U9011 (N_9011,N_8134,N_8421);
and U9012 (N_9012,N_8280,N_8799);
nand U9013 (N_9013,N_8045,N_8415);
or U9014 (N_9014,N_8617,N_8793);
nor U9015 (N_9015,N_8108,N_8741);
nand U9016 (N_9016,N_8340,N_8731);
nor U9017 (N_9017,N_8540,N_8062);
nand U9018 (N_9018,N_8007,N_8253);
and U9019 (N_9019,N_8732,N_8201);
nor U9020 (N_9020,N_8041,N_8620);
and U9021 (N_9021,N_8665,N_8445);
nand U9022 (N_9022,N_8030,N_8426);
nor U9023 (N_9023,N_8673,N_8669);
nor U9024 (N_9024,N_8720,N_8058);
and U9025 (N_9025,N_8303,N_8505);
or U9026 (N_9026,N_8566,N_8176);
nor U9027 (N_9027,N_8235,N_8127);
or U9028 (N_9028,N_8713,N_8324);
and U9029 (N_9029,N_8383,N_8081);
and U9030 (N_9030,N_8750,N_8304);
nor U9031 (N_9031,N_8603,N_8761);
nand U9032 (N_9032,N_8083,N_8674);
nor U9033 (N_9033,N_8257,N_8211);
nor U9034 (N_9034,N_8131,N_8560);
nor U9035 (N_9035,N_8672,N_8591);
or U9036 (N_9036,N_8331,N_8693);
nor U9037 (N_9037,N_8605,N_8160);
and U9038 (N_9038,N_8767,N_8021);
and U9039 (N_9039,N_8520,N_8589);
and U9040 (N_9040,N_8498,N_8321);
or U9041 (N_9041,N_8738,N_8171);
nand U9042 (N_9042,N_8130,N_8074);
nor U9043 (N_9043,N_8691,N_8638);
and U9044 (N_9044,N_8664,N_8470);
and U9045 (N_9045,N_8710,N_8187);
or U9046 (N_9046,N_8429,N_8412);
nand U9047 (N_9047,N_8013,N_8128);
nor U9048 (N_9048,N_8727,N_8695);
nand U9049 (N_9049,N_8690,N_8466);
and U9050 (N_9050,N_8414,N_8717);
nand U9051 (N_9051,N_8780,N_8686);
nor U9052 (N_9052,N_8444,N_8208);
and U9053 (N_9053,N_8163,N_8027);
and U9054 (N_9054,N_8099,N_8462);
and U9055 (N_9055,N_8659,N_8102);
nor U9056 (N_9056,N_8764,N_8319);
or U9057 (N_9057,N_8598,N_8702);
nor U9058 (N_9058,N_8124,N_8247);
and U9059 (N_9059,N_8264,N_8622);
nand U9060 (N_9060,N_8114,N_8795);
and U9061 (N_9061,N_8116,N_8136);
or U9062 (N_9062,N_8182,N_8679);
or U9063 (N_9063,N_8459,N_8512);
and U9064 (N_9064,N_8150,N_8716);
and U9065 (N_9065,N_8516,N_8396);
or U9066 (N_9066,N_8751,N_8681);
nand U9067 (N_9067,N_8504,N_8159);
nor U9068 (N_9068,N_8010,N_8722);
nand U9069 (N_9069,N_8348,N_8766);
and U9070 (N_9070,N_8632,N_8308);
nor U9071 (N_9071,N_8583,N_8241);
xor U9072 (N_9072,N_8621,N_8286);
or U9073 (N_9073,N_8577,N_8465);
nor U9074 (N_9074,N_8172,N_8646);
nor U9075 (N_9075,N_8381,N_8229);
and U9076 (N_9076,N_8436,N_8488);
and U9077 (N_9077,N_8486,N_8469);
or U9078 (N_9078,N_8653,N_8573);
and U9079 (N_9079,N_8284,N_8398);
or U9080 (N_9080,N_8787,N_8796);
or U9081 (N_9081,N_8004,N_8708);
or U9082 (N_9082,N_8550,N_8054);
and U9083 (N_9083,N_8387,N_8675);
nor U9084 (N_9084,N_8786,N_8267);
nand U9085 (N_9085,N_8289,N_8775);
and U9086 (N_9086,N_8209,N_8707);
and U9087 (N_9087,N_8417,N_8048);
or U9088 (N_9088,N_8117,N_8336);
or U9089 (N_9089,N_8684,N_8650);
nand U9090 (N_9090,N_8425,N_8528);
nor U9091 (N_9091,N_8728,N_8316);
or U9092 (N_9092,N_8606,N_8773);
nand U9093 (N_9093,N_8019,N_8655);
nor U9094 (N_9094,N_8476,N_8737);
nand U9095 (N_9095,N_8093,N_8721);
nand U9096 (N_9096,N_8115,N_8446);
or U9097 (N_9097,N_8543,N_8195);
nor U9098 (N_9098,N_8778,N_8049);
nor U9099 (N_9099,N_8492,N_8748);
and U9100 (N_9100,N_8798,N_8268);
or U9101 (N_9101,N_8011,N_8471);
nor U9102 (N_9102,N_8575,N_8290);
and U9103 (N_9103,N_8533,N_8555);
or U9104 (N_9104,N_8075,N_8068);
or U9105 (N_9105,N_8148,N_8394);
nor U9106 (N_9106,N_8413,N_8186);
and U9107 (N_9107,N_8706,N_8406);
nor U9108 (N_9108,N_8228,N_8281);
and U9109 (N_9109,N_8433,N_8402);
or U9110 (N_9110,N_8443,N_8122);
nand U9111 (N_9111,N_8531,N_8502);
and U9112 (N_9112,N_8790,N_8165);
nand U9113 (N_9113,N_8366,N_8288);
and U9114 (N_9114,N_8224,N_8145);
and U9115 (N_9115,N_8497,N_8183);
xnor U9116 (N_9116,N_8564,N_8569);
nor U9117 (N_9117,N_8178,N_8719);
nor U9118 (N_9118,N_8521,N_8472);
nand U9119 (N_9119,N_8557,N_8103);
nor U9120 (N_9120,N_8448,N_8090);
nor U9121 (N_9121,N_8219,N_8699);
and U9122 (N_9122,N_8053,N_8490);
or U9123 (N_9123,N_8418,N_8260);
nor U9124 (N_9124,N_8584,N_8461);
nand U9125 (N_9125,N_8676,N_8064);
nand U9126 (N_9126,N_8582,N_8489);
nand U9127 (N_9127,N_8404,N_8643);
nor U9128 (N_9128,N_8539,N_8689);
or U9129 (N_9129,N_8377,N_8590);
nand U9130 (N_9130,N_8657,N_8517);
nand U9131 (N_9131,N_8265,N_8328);
xnor U9132 (N_9132,N_8051,N_8515);
nor U9133 (N_9133,N_8735,N_8536);
or U9134 (N_9134,N_8507,N_8438);
or U9135 (N_9135,N_8747,N_8262);
nand U9136 (N_9136,N_8704,N_8758);
nand U9137 (N_9137,N_8698,N_8368);
nor U9138 (N_9138,N_8496,N_8305);
and U9139 (N_9139,N_8756,N_8047);
and U9140 (N_9140,N_8283,N_8556);
nand U9141 (N_9141,N_8449,N_8395);
nand U9142 (N_9142,N_8616,N_8595);
or U9143 (N_9143,N_8215,N_8753);
and U9144 (N_9144,N_8510,N_8619);
nand U9145 (N_9145,N_8285,N_8269);
and U9146 (N_9146,N_8106,N_8552);
or U9147 (N_9147,N_8779,N_8164);
nand U9148 (N_9148,N_8437,N_8518);
and U9149 (N_9149,N_8792,N_8457);
or U9150 (N_9150,N_8261,N_8184);
nor U9151 (N_9151,N_8193,N_8705);
or U9152 (N_9152,N_8123,N_8743);
and U9153 (N_9153,N_8772,N_8040);
nor U9154 (N_9154,N_8240,N_8481);
nand U9155 (N_9155,N_8736,N_8370);
or U9156 (N_9156,N_8349,N_8688);
or U9157 (N_9157,N_8453,N_8485);
nand U9158 (N_9158,N_8140,N_8100);
and U9159 (N_9159,N_8332,N_8570);
and U9160 (N_9160,N_8152,N_8568);
nand U9161 (N_9161,N_8754,N_8561);
or U9162 (N_9162,N_8380,N_8765);
and U9163 (N_9163,N_8467,N_8596);
or U9164 (N_9164,N_8797,N_8111);
nand U9165 (N_9165,N_8361,N_8357);
nor U9166 (N_9166,N_8351,N_8501);
nand U9167 (N_9167,N_8325,N_8222);
nor U9168 (N_9168,N_8360,N_8514);
and U9169 (N_9169,N_8154,N_8017);
or U9170 (N_9170,N_8213,N_8388);
or U9171 (N_9171,N_8640,N_8141);
or U9172 (N_9172,N_8031,N_8151);
nor U9173 (N_9173,N_8263,N_8645);
nor U9174 (N_9174,N_8424,N_8138);
nand U9175 (N_9175,N_8757,N_8291);
nor U9176 (N_9176,N_8227,N_8139);
or U9177 (N_9177,N_8270,N_8302);
or U9178 (N_9178,N_8371,N_8087);
or U9179 (N_9179,N_8248,N_8783);
nor U9180 (N_9180,N_8547,N_8759);
nor U9181 (N_9181,N_8299,N_8399);
nor U9182 (N_9182,N_8422,N_8039);
nand U9183 (N_9183,N_8109,N_8586);
nor U9184 (N_9184,N_8097,N_8661);
nor U9185 (N_9185,N_8226,N_8322);
or U9186 (N_9186,N_8157,N_8529);
and U9187 (N_9187,N_8277,N_8670);
nor U9188 (N_9188,N_8715,N_8410);
nor U9189 (N_9189,N_8562,N_8153);
and U9190 (N_9190,N_8089,N_8234);
and U9191 (N_9191,N_8206,N_8576);
or U9192 (N_9192,N_8678,N_8044);
nand U9193 (N_9193,N_8298,N_8167);
and U9194 (N_9194,N_8317,N_8683);
nand U9195 (N_9195,N_8359,N_8309);
and U9196 (N_9196,N_8513,N_8059);
nand U9197 (N_9197,N_8572,N_8755);
nor U9198 (N_9198,N_8071,N_8420);
or U9199 (N_9199,N_8656,N_8479);
nor U9200 (N_9200,N_8416,N_8565);
and U9201 (N_9201,N_8470,N_8082);
or U9202 (N_9202,N_8379,N_8438);
nor U9203 (N_9203,N_8555,N_8783);
nand U9204 (N_9204,N_8674,N_8581);
and U9205 (N_9205,N_8050,N_8474);
nor U9206 (N_9206,N_8672,N_8485);
or U9207 (N_9207,N_8207,N_8795);
or U9208 (N_9208,N_8615,N_8625);
and U9209 (N_9209,N_8076,N_8480);
nor U9210 (N_9210,N_8133,N_8625);
nand U9211 (N_9211,N_8520,N_8263);
nor U9212 (N_9212,N_8315,N_8112);
nand U9213 (N_9213,N_8748,N_8146);
or U9214 (N_9214,N_8697,N_8664);
and U9215 (N_9215,N_8715,N_8197);
and U9216 (N_9216,N_8186,N_8679);
and U9217 (N_9217,N_8328,N_8073);
nand U9218 (N_9218,N_8222,N_8249);
nand U9219 (N_9219,N_8101,N_8090);
and U9220 (N_9220,N_8646,N_8700);
nor U9221 (N_9221,N_8784,N_8614);
and U9222 (N_9222,N_8769,N_8729);
and U9223 (N_9223,N_8029,N_8283);
nor U9224 (N_9224,N_8665,N_8703);
nand U9225 (N_9225,N_8136,N_8143);
nand U9226 (N_9226,N_8238,N_8510);
nand U9227 (N_9227,N_8683,N_8771);
nand U9228 (N_9228,N_8556,N_8478);
and U9229 (N_9229,N_8250,N_8753);
or U9230 (N_9230,N_8388,N_8608);
or U9231 (N_9231,N_8211,N_8743);
or U9232 (N_9232,N_8114,N_8217);
and U9233 (N_9233,N_8649,N_8675);
nand U9234 (N_9234,N_8194,N_8424);
and U9235 (N_9235,N_8712,N_8779);
nor U9236 (N_9236,N_8586,N_8640);
nor U9237 (N_9237,N_8457,N_8650);
nor U9238 (N_9238,N_8314,N_8430);
nor U9239 (N_9239,N_8410,N_8556);
nand U9240 (N_9240,N_8761,N_8657);
nand U9241 (N_9241,N_8240,N_8184);
or U9242 (N_9242,N_8587,N_8731);
and U9243 (N_9243,N_8279,N_8062);
or U9244 (N_9244,N_8450,N_8772);
and U9245 (N_9245,N_8095,N_8031);
or U9246 (N_9246,N_8248,N_8223);
xnor U9247 (N_9247,N_8523,N_8460);
nand U9248 (N_9248,N_8787,N_8408);
nor U9249 (N_9249,N_8090,N_8041);
nor U9250 (N_9250,N_8193,N_8756);
nand U9251 (N_9251,N_8162,N_8668);
nor U9252 (N_9252,N_8638,N_8492);
xnor U9253 (N_9253,N_8594,N_8698);
or U9254 (N_9254,N_8641,N_8282);
nand U9255 (N_9255,N_8505,N_8545);
and U9256 (N_9256,N_8322,N_8789);
or U9257 (N_9257,N_8303,N_8792);
nor U9258 (N_9258,N_8296,N_8178);
nand U9259 (N_9259,N_8258,N_8747);
or U9260 (N_9260,N_8717,N_8166);
nand U9261 (N_9261,N_8086,N_8756);
or U9262 (N_9262,N_8712,N_8342);
nand U9263 (N_9263,N_8088,N_8081);
nand U9264 (N_9264,N_8124,N_8123);
and U9265 (N_9265,N_8391,N_8150);
nor U9266 (N_9266,N_8525,N_8022);
or U9267 (N_9267,N_8378,N_8203);
or U9268 (N_9268,N_8041,N_8709);
or U9269 (N_9269,N_8412,N_8033);
nand U9270 (N_9270,N_8124,N_8750);
or U9271 (N_9271,N_8572,N_8268);
or U9272 (N_9272,N_8526,N_8054);
nand U9273 (N_9273,N_8396,N_8775);
and U9274 (N_9274,N_8329,N_8128);
and U9275 (N_9275,N_8355,N_8310);
or U9276 (N_9276,N_8619,N_8577);
and U9277 (N_9277,N_8303,N_8788);
or U9278 (N_9278,N_8283,N_8132);
and U9279 (N_9279,N_8297,N_8152);
nor U9280 (N_9280,N_8316,N_8627);
and U9281 (N_9281,N_8434,N_8698);
or U9282 (N_9282,N_8400,N_8396);
nand U9283 (N_9283,N_8183,N_8417);
nand U9284 (N_9284,N_8285,N_8530);
and U9285 (N_9285,N_8713,N_8210);
or U9286 (N_9286,N_8261,N_8762);
nor U9287 (N_9287,N_8306,N_8294);
nand U9288 (N_9288,N_8058,N_8131);
nor U9289 (N_9289,N_8476,N_8191);
nand U9290 (N_9290,N_8352,N_8573);
nand U9291 (N_9291,N_8445,N_8748);
or U9292 (N_9292,N_8300,N_8343);
nand U9293 (N_9293,N_8416,N_8634);
nand U9294 (N_9294,N_8263,N_8100);
and U9295 (N_9295,N_8010,N_8237);
nor U9296 (N_9296,N_8067,N_8324);
nand U9297 (N_9297,N_8632,N_8134);
or U9298 (N_9298,N_8598,N_8443);
nand U9299 (N_9299,N_8386,N_8626);
or U9300 (N_9300,N_8647,N_8377);
and U9301 (N_9301,N_8704,N_8150);
nand U9302 (N_9302,N_8070,N_8657);
nand U9303 (N_9303,N_8662,N_8601);
and U9304 (N_9304,N_8510,N_8476);
nand U9305 (N_9305,N_8181,N_8380);
nor U9306 (N_9306,N_8547,N_8489);
nor U9307 (N_9307,N_8483,N_8430);
or U9308 (N_9308,N_8750,N_8289);
and U9309 (N_9309,N_8423,N_8587);
or U9310 (N_9310,N_8737,N_8352);
and U9311 (N_9311,N_8263,N_8014);
or U9312 (N_9312,N_8593,N_8482);
and U9313 (N_9313,N_8144,N_8486);
nand U9314 (N_9314,N_8482,N_8455);
or U9315 (N_9315,N_8642,N_8184);
and U9316 (N_9316,N_8501,N_8528);
nor U9317 (N_9317,N_8618,N_8153);
nand U9318 (N_9318,N_8448,N_8295);
nor U9319 (N_9319,N_8332,N_8101);
or U9320 (N_9320,N_8735,N_8526);
and U9321 (N_9321,N_8137,N_8652);
nand U9322 (N_9322,N_8258,N_8522);
nand U9323 (N_9323,N_8064,N_8697);
or U9324 (N_9324,N_8588,N_8296);
nor U9325 (N_9325,N_8727,N_8176);
nand U9326 (N_9326,N_8333,N_8567);
nor U9327 (N_9327,N_8665,N_8721);
nand U9328 (N_9328,N_8722,N_8377);
nand U9329 (N_9329,N_8447,N_8720);
or U9330 (N_9330,N_8022,N_8166);
nand U9331 (N_9331,N_8024,N_8136);
nor U9332 (N_9332,N_8196,N_8719);
nor U9333 (N_9333,N_8612,N_8132);
or U9334 (N_9334,N_8510,N_8714);
xnor U9335 (N_9335,N_8504,N_8452);
nand U9336 (N_9336,N_8173,N_8058);
or U9337 (N_9337,N_8219,N_8734);
or U9338 (N_9338,N_8235,N_8069);
nor U9339 (N_9339,N_8327,N_8500);
nand U9340 (N_9340,N_8164,N_8758);
nand U9341 (N_9341,N_8359,N_8646);
and U9342 (N_9342,N_8161,N_8315);
xnor U9343 (N_9343,N_8580,N_8491);
and U9344 (N_9344,N_8421,N_8367);
or U9345 (N_9345,N_8754,N_8334);
nor U9346 (N_9346,N_8268,N_8201);
or U9347 (N_9347,N_8298,N_8673);
nand U9348 (N_9348,N_8662,N_8537);
or U9349 (N_9349,N_8527,N_8024);
nand U9350 (N_9350,N_8663,N_8630);
nor U9351 (N_9351,N_8109,N_8320);
nand U9352 (N_9352,N_8769,N_8347);
nor U9353 (N_9353,N_8288,N_8679);
nor U9354 (N_9354,N_8173,N_8354);
nand U9355 (N_9355,N_8510,N_8775);
nor U9356 (N_9356,N_8450,N_8351);
or U9357 (N_9357,N_8566,N_8187);
nand U9358 (N_9358,N_8103,N_8263);
or U9359 (N_9359,N_8204,N_8076);
and U9360 (N_9360,N_8655,N_8772);
nor U9361 (N_9361,N_8734,N_8018);
and U9362 (N_9362,N_8282,N_8460);
nand U9363 (N_9363,N_8127,N_8713);
nand U9364 (N_9364,N_8433,N_8015);
and U9365 (N_9365,N_8562,N_8053);
nor U9366 (N_9366,N_8796,N_8601);
and U9367 (N_9367,N_8307,N_8645);
nor U9368 (N_9368,N_8191,N_8305);
nand U9369 (N_9369,N_8743,N_8016);
or U9370 (N_9370,N_8530,N_8242);
nand U9371 (N_9371,N_8257,N_8285);
and U9372 (N_9372,N_8435,N_8353);
and U9373 (N_9373,N_8045,N_8254);
nor U9374 (N_9374,N_8067,N_8025);
and U9375 (N_9375,N_8208,N_8284);
and U9376 (N_9376,N_8533,N_8396);
nor U9377 (N_9377,N_8011,N_8421);
or U9378 (N_9378,N_8445,N_8560);
nor U9379 (N_9379,N_8060,N_8404);
or U9380 (N_9380,N_8466,N_8350);
nor U9381 (N_9381,N_8631,N_8721);
or U9382 (N_9382,N_8694,N_8094);
and U9383 (N_9383,N_8434,N_8756);
nor U9384 (N_9384,N_8297,N_8485);
or U9385 (N_9385,N_8266,N_8596);
nand U9386 (N_9386,N_8197,N_8714);
and U9387 (N_9387,N_8457,N_8143);
or U9388 (N_9388,N_8646,N_8136);
nor U9389 (N_9389,N_8567,N_8201);
nor U9390 (N_9390,N_8069,N_8726);
or U9391 (N_9391,N_8055,N_8304);
nand U9392 (N_9392,N_8710,N_8325);
nand U9393 (N_9393,N_8485,N_8255);
nand U9394 (N_9394,N_8414,N_8070);
or U9395 (N_9395,N_8648,N_8035);
and U9396 (N_9396,N_8066,N_8590);
nand U9397 (N_9397,N_8394,N_8112);
or U9398 (N_9398,N_8618,N_8145);
nor U9399 (N_9399,N_8257,N_8547);
nand U9400 (N_9400,N_8340,N_8675);
and U9401 (N_9401,N_8580,N_8548);
and U9402 (N_9402,N_8356,N_8532);
or U9403 (N_9403,N_8413,N_8456);
and U9404 (N_9404,N_8040,N_8726);
and U9405 (N_9405,N_8676,N_8322);
and U9406 (N_9406,N_8535,N_8190);
nor U9407 (N_9407,N_8533,N_8236);
nor U9408 (N_9408,N_8438,N_8418);
nand U9409 (N_9409,N_8564,N_8674);
and U9410 (N_9410,N_8517,N_8592);
nand U9411 (N_9411,N_8061,N_8744);
nor U9412 (N_9412,N_8122,N_8548);
nor U9413 (N_9413,N_8091,N_8166);
nor U9414 (N_9414,N_8725,N_8201);
nand U9415 (N_9415,N_8043,N_8638);
and U9416 (N_9416,N_8625,N_8714);
or U9417 (N_9417,N_8617,N_8624);
and U9418 (N_9418,N_8020,N_8784);
or U9419 (N_9419,N_8078,N_8001);
nand U9420 (N_9420,N_8078,N_8534);
or U9421 (N_9421,N_8744,N_8664);
or U9422 (N_9422,N_8487,N_8203);
nand U9423 (N_9423,N_8566,N_8673);
nand U9424 (N_9424,N_8186,N_8395);
nand U9425 (N_9425,N_8114,N_8489);
nor U9426 (N_9426,N_8069,N_8170);
nor U9427 (N_9427,N_8306,N_8325);
nor U9428 (N_9428,N_8024,N_8347);
nand U9429 (N_9429,N_8389,N_8419);
or U9430 (N_9430,N_8765,N_8627);
and U9431 (N_9431,N_8170,N_8626);
and U9432 (N_9432,N_8546,N_8158);
nor U9433 (N_9433,N_8108,N_8776);
or U9434 (N_9434,N_8336,N_8280);
and U9435 (N_9435,N_8555,N_8448);
or U9436 (N_9436,N_8757,N_8231);
or U9437 (N_9437,N_8770,N_8083);
and U9438 (N_9438,N_8263,N_8127);
and U9439 (N_9439,N_8261,N_8004);
xor U9440 (N_9440,N_8333,N_8206);
or U9441 (N_9441,N_8330,N_8252);
or U9442 (N_9442,N_8083,N_8592);
and U9443 (N_9443,N_8242,N_8087);
and U9444 (N_9444,N_8282,N_8449);
nand U9445 (N_9445,N_8115,N_8086);
or U9446 (N_9446,N_8748,N_8325);
and U9447 (N_9447,N_8348,N_8608);
and U9448 (N_9448,N_8781,N_8385);
and U9449 (N_9449,N_8279,N_8659);
or U9450 (N_9450,N_8095,N_8296);
or U9451 (N_9451,N_8587,N_8127);
and U9452 (N_9452,N_8450,N_8631);
and U9453 (N_9453,N_8251,N_8518);
nor U9454 (N_9454,N_8560,N_8093);
nor U9455 (N_9455,N_8407,N_8783);
nor U9456 (N_9456,N_8739,N_8450);
nand U9457 (N_9457,N_8191,N_8038);
and U9458 (N_9458,N_8199,N_8021);
and U9459 (N_9459,N_8397,N_8290);
and U9460 (N_9460,N_8084,N_8503);
nor U9461 (N_9461,N_8105,N_8601);
and U9462 (N_9462,N_8642,N_8469);
and U9463 (N_9463,N_8600,N_8201);
nor U9464 (N_9464,N_8688,N_8664);
xnor U9465 (N_9465,N_8578,N_8151);
nand U9466 (N_9466,N_8111,N_8434);
nand U9467 (N_9467,N_8280,N_8708);
nand U9468 (N_9468,N_8580,N_8365);
or U9469 (N_9469,N_8562,N_8032);
and U9470 (N_9470,N_8164,N_8329);
and U9471 (N_9471,N_8231,N_8071);
or U9472 (N_9472,N_8111,N_8688);
nor U9473 (N_9473,N_8088,N_8588);
nor U9474 (N_9474,N_8674,N_8583);
nand U9475 (N_9475,N_8032,N_8507);
or U9476 (N_9476,N_8421,N_8014);
or U9477 (N_9477,N_8392,N_8575);
nand U9478 (N_9478,N_8156,N_8521);
nor U9479 (N_9479,N_8100,N_8133);
nor U9480 (N_9480,N_8525,N_8328);
nand U9481 (N_9481,N_8463,N_8511);
or U9482 (N_9482,N_8460,N_8098);
xnor U9483 (N_9483,N_8747,N_8465);
nor U9484 (N_9484,N_8589,N_8508);
or U9485 (N_9485,N_8082,N_8229);
or U9486 (N_9486,N_8391,N_8155);
nor U9487 (N_9487,N_8099,N_8566);
nand U9488 (N_9488,N_8455,N_8477);
nor U9489 (N_9489,N_8280,N_8203);
or U9490 (N_9490,N_8767,N_8533);
or U9491 (N_9491,N_8454,N_8649);
nand U9492 (N_9492,N_8247,N_8026);
or U9493 (N_9493,N_8722,N_8263);
and U9494 (N_9494,N_8370,N_8080);
nand U9495 (N_9495,N_8432,N_8731);
nand U9496 (N_9496,N_8126,N_8637);
or U9497 (N_9497,N_8531,N_8159);
or U9498 (N_9498,N_8067,N_8478);
or U9499 (N_9499,N_8790,N_8429);
nor U9500 (N_9500,N_8089,N_8718);
nor U9501 (N_9501,N_8315,N_8231);
or U9502 (N_9502,N_8231,N_8703);
and U9503 (N_9503,N_8245,N_8253);
nand U9504 (N_9504,N_8262,N_8688);
or U9505 (N_9505,N_8643,N_8229);
or U9506 (N_9506,N_8429,N_8413);
nor U9507 (N_9507,N_8127,N_8744);
or U9508 (N_9508,N_8379,N_8448);
and U9509 (N_9509,N_8672,N_8308);
and U9510 (N_9510,N_8515,N_8219);
nand U9511 (N_9511,N_8477,N_8285);
nor U9512 (N_9512,N_8743,N_8666);
nand U9513 (N_9513,N_8239,N_8307);
nor U9514 (N_9514,N_8139,N_8608);
nor U9515 (N_9515,N_8705,N_8468);
nand U9516 (N_9516,N_8743,N_8629);
nand U9517 (N_9517,N_8510,N_8114);
or U9518 (N_9518,N_8018,N_8699);
or U9519 (N_9519,N_8436,N_8377);
nor U9520 (N_9520,N_8350,N_8156);
nand U9521 (N_9521,N_8502,N_8217);
or U9522 (N_9522,N_8619,N_8151);
nand U9523 (N_9523,N_8374,N_8185);
and U9524 (N_9524,N_8096,N_8008);
nand U9525 (N_9525,N_8103,N_8634);
nand U9526 (N_9526,N_8038,N_8104);
or U9527 (N_9527,N_8585,N_8055);
nand U9528 (N_9528,N_8444,N_8031);
nor U9529 (N_9529,N_8605,N_8041);
nor U9530 (N_9530,N_8043,N_8678);
or U9531 (N_9531,N_8265,N_8020);
and U9532 (N_9532,N_8524,N_8368);
or U9533 (N_9533,N_8017,N_8573);
and U9534 (N_9534,N_8390,N_8568);
and U9535 (N_9535,N_8583,N_8770);
nand U9536 (N_9536,N_8467,N_8394);
or U9537 (N_9537,N_8175,N_8477);
nor U9538 (N_9538,N_8216,N_8412);
nor U9539 (N_9539,N_8529,N_8718);
or U9540 (N_9540,N_8668,N_8092);
and U9541 (N_9541,N_8447,N_8165);
or U9542 (N_9542,N_8568,N_8186);
and U9543 (N_9543,N_8133,N_8059);
or U9544 (N_9544,N_8056,N_8765);
nand U9545 (N_9545,N_8346,N_8044);
nand U9546 (N_9546,N_8434,N_8147);
nand U9547 (N_9547,N_8232,N_8210);
nor U9548 (N_9548,N_8518,N_8500);
nor U9549 (N_9549,N_8070,N_8393);
nor U9550 (N_9550,N_8250,N_8607);
and U9551 (N_9551,N_8608,N_8716);
nand U9552 (N_9552,N_8331,N_8578);
or U9553 (N_9553,N_8558,N_8777);
nand U9554 (N_9554,N_8290,N_8550);
or U9555 (N_9555,N_8194,N_8704);
nor U9556 (N_9556,N_8736,N_8642);
nor U9557 (N_9557,N_8546,N_8097);
or U9558 (N_9558,N_8405,N_8690);
nor U9559 (N_9559,N_8351,N_8669);
or U9560 (N_9560,N_8114,N_8276);
and U9561 (N_9561,N_8511,N_8241);
nand U9562 (N_9562,N_8133,N_8148);
nand U9563 (N_9563,N_8138,N_8254);
nor U9564 (N_9564,N_8147,N_8287);
nor U9565 (N_9565,N_8529,N_8565);
or U9566 (N_9566,N_8550,N_8589);
or U9567 (N_9567,N_8363,N_8136);
or U9568 (N_9568,N_8695,N_8442);
nand U9569 (N_9569,N_8529,N_8240);
nor U9570 (N_9570,N_8765,N_8647);
and U9571 (N_9571,N_8434,N_8218);
nand U9572 (N_9572,N_8440,N_8755);
or U9573 (N_9573,N_8680,N_8460);
or U9574 (N_9574,N_8457,N_8551);
or U9575 (N_9575,N_8106,N_8237);
nor U9576 (N_9576,N_8350,N_8140);
nor U9577 (N_9577,N_8580,N_8799);
and U9578 (N_9578,N_8089,N_8236);
nand U9579 (N_9579,N_8738,N_8270);
nor U9580 (N_9580,N_8438,N_8307);
and U9581 (N_9581,N_8536,N_8206);
nor U9582 (N_9582,N_8639,N_8263);
nand U9583 (N_9583,N_8765,N_8288);
or U9584 (N_9584,N_8496,N_8728);
nor U9585 (N_9585,N_8135,N_8291);
or U9586 (N_9586,N_8190,N_8610);
nor U9587 (N_9587,N_8220,N_8165);
nand U9588 (N_9588,N_8332,N_8149);
or U9589 (N_9589,N_8702,N_8722);
nand U9590 (N_9590,N_8781,N_8366);
or U9591 (N_9591,N_8440,N_8017);
or U9592 (N_9592,N_8698,N_8508);
and U9593 (N_9593,N_8716,N_8609);
nand U9594 (N_9594,N_8452,N_8135);
or U9595 (N_9595,N_8580,N_8429);
nand U9596 (N_9596,N_8311,N_8237);
nor U9597 (N_9597,N_8167,N_8390);
and U9598 (N_9598,N_8793,N_8306);
or U9599 (N_9599,N_8333,N_8553);
nor U9600 (N_9600,N_9055,N_9200);
and U9601 (N_9601,N_9023,N_9275);
and U9602 (N_9602,N_9296,N_9422);
nand U9603 (N_9603,N_9056,N_9160);
and U9604 (N_9604,N_9580,N_9110);
and U9605 (N_9605,N_9000,N_9205);
nor U9606 (N_9606,N_9181,N_8911);
nand U9607 (N_9607,N_9093,N_8869);
and U9608 (N_9608,N_9058,N_9236);
or U9609 (N_9609,N_9428,N_9437);
nor U9610 (N_9610,N_9145,N_9177);
and U9611 (N_9611,N_8928,N_9375);
or U9612 (N_9612,N_9231,N_8841);
nand U9613 (N_9613,N_9046,N_9050);
nor U9614 (N_9614,N_9036,N_9596);
and U9615 (N_9615,N_9190,N_9303);
or U9616 (N_9616,N_9116,N_8844);
or U9617 (N_9617,N_8938,N_9455);
and U9618 (N_9618,N_8831,N_9387);
nor U9619 (N_9619,N_8822,N_8860);
nand U9620 (N_9620,N_8919,N_9156);
and U9621 (N_9621,N_9142,N_8840);
nor U9622 (N_9622,N_9026,N_8880);
nand U9623 (N_9623,N_9348,N_9277);
nand U9624 (N_9624,N_9191,N_9176);
nor U9625 (N_9625,N_9589,N_8908);
nor U9626 (N_9626,N_9483,N_9458);
and U9627 (N_9627,N_9328,N_9057);
or U9628 (N_9628,N_9425,N_9140);
nor U9629 (N_9629,N_8990,N_9300);
and U9630 (N_9630,N_8905,N_9249);
or U9631 (N_9631,N_9373,N_9395);
or U9632 (N_9632,N_8848,N_8963);
or U9633 (N_9633,N_8944,N_9529);
and U9634 (N_9634,N_9339,N_9144);
nor U9635 (N_9635,N_9486,N_9267);
and U9636 (N_9636,N_9180,N_9506);
or U9637 (N_9637,N_8981,N_9105);
or U9638 (N_9638,N_9561,N_8940);
nor U9639 (N_9639,N_8918,N_9418);
nor U9640 (N_9640,N_8943,N_9098);
and U9641 (N_9641,N_9208,N_9111);
nand U9642 (N_9642,N_9146,N_9431);
or U9643 (N_9643,N_9376,N_9013);
nand U9644 (N_9644,N_9517,N_9563);
nor U9645 (N_9645,N_9084,N_8900);
or U9646 (N_9646,N_9448,N_9594);
and U9647 (N_9647,N_8913,N_9209);
nor U9648 (N_9648,N_8967,N_9169);
nand U9649 (N_9649,N_9288,N_9312);
and U9650 (N_9650,N_9166,N_9283);
or U9651 (N_9651,N_9578,N_9253);
and U9652 (N_9652,N_9570,N_9310);
nor U9653 (N_9653,N_9149,N_9456);
or U9654 (N_9654,N_9158,N_9281);
and U9655 (N_9655,N_9039,N_9519);
or U9656 (N_9656,N_8916,N_9479);
nand U9657 (N_9657,N_9152,N_9081);
and U9658 (N_9658,N_9393,N_9441);
and U9659 (N_9659,N_9243,N_8932);
and U9660 (N_9660,N_8927,N_9095);
or U9661 (N_9661,N_9014,N_9035);
or U9662 (N_9662,N_9047,N_9223);
and U9663 (N_9663,N_9513,N_9043);
nand U9664 (N_9664,N_9525,N_9193);
nor U9665 (N_9665,N_9510,N_9087);
nand U9666 (N_9666,N_8856,N_9133);
nor U9667 (N_9667,N_9289,N_9385);
or U9668 (N_9668,N_9279,N_8827);
nand U9669 (N_9669,N_9263,N_9357);
nor U9670 (N_9670,N_9558,N_9531);
nand U9671 (N_9671,N_9311,N_8882);
nor U9672 (N_9672,N_9262,N_9031);
and U9673 (N_9673,N_9079,N_8941);
nor U9674 (N_9674,N_9250,N_9413);
or U9675 (N_9675,N_9030,N_9466);
xor U9676 (N_9676,N_9421,N_9521);
and U9677 (N_9677,N_8874,N_9503);
and U9678 (N_9678,N_9259,N_8912);
nand U9679 (N_9679,N_9365,N_9244);
nand U9680 (N_9680,N_9215,N_9196);
nor U9681 (N_9681,N_9576,N_9470);
nand U9682 (N_9682,N_9113,N_8890);
nor U9683 (N_9683,N_9167,N_8846);
and U9684 (N_9684,N_9178,N_9457);
nand U9685 (N_9685,N_8823,N_8865);
and U9686 (N_9686,N_8920,N_9082);
and U9687 (N_9687,N_9439,N_9374);
nor U9688 (N_9688,N_9235,N_9320);
nor U9689 (N_9689,N_9416,N_9528);
and U9690 (N_9690,N_9392,N_9526);
and U9691 (N_9691,N_8946,N_9069);
and U9692 (N_9692,N_9294,N_9543);
and U9693 (N_9693,N_9547,N_8857);
and U9694 (N_9694,N_9153,N_9340);
nor U9695 (N_9695,N_8888,N_9234);
and U9696 (N_9696,N_8804,N_9114);
or U9697 (N_9697,N_9327,N_8934);
or U9698 (N_9698,N_9382,N_9165);
nand U9699 (N_9699,N_9151,N_9171);
or U9700 (N_9700,N_9045,N_8850);
and U9701 (N_9701,N_8942,N_8925);
or U9702 (N_9702,N_8903,N_9060);
or U9703 (N_9703,N_8892,N_9430);
nand U9704 (N_9704,N_9265,N_8962);
nor U9705 (N_9705,N_8839,N_8945);
or U9706 (N_9706,N_9468,N_9390);
nand U9707 (N_9707,N_9398,N_9593);
or U9708 (N_9708,N_9076,N_9257);
nand U9709 (N_9709,N_9012,N_9203);
and U9710 (N_9710,N_8834,N_9505);
nand U9711 (N_9711,N_9371,N_9233);
nand U9712 (N_9712,N_8852,N_9509);
nand U9713 (N_9713,N_9463,N_9366);
nand U9714 (N_9714,N_8838,N_9388);
nand U9715 (N_9715,N_9567,N_9522);
or U9716 (N_9716,N_9029,N_9588);
nor U9717 (N_9717,N_9227,N_9299);
nor U9718 (N_9718,N_8931,N_9112);
nor U9719 (N_9719,N_9564,N_8878);
and U9720 (N_9720,N_8982,N_9332);
nor U9721 (N_9721,N_8847,N_9559);
nor U9722 (N_9722,N_9461,N_9402);
nor U9723 (N_9723,N_9341,N_9285);
or U9724 (N_9724,N_9345,N_8969);
nand U9725 (N_9725,N_9380,N_8876);
nor U9726 (N_9726,N_8817,N_9216);
or U9727 (N_9727,N_9094,N_9063);
nor U9728 (N_9728,N_9117,N_8868);
nor U9729 (N_9729,N_9027,N_8836);
nor U9730 (N_9730,N_9273,N_9099);
or U9731 (N_9731,N_9214,N_9230);
or U9732 (N_9732,N_9305,N_9358);
or U9733 (N_9733,N_9383,N_9286);
and U9734 (N_9734,N_9122,N_9225);
or U9735 (N_9735,N_9183,N_9507);
nand U9736 (N_9736,N_9579,N_9220);
nand U9737 (N_9737,N_9308,N_8801);
nor U9738 (N_9738,N_9555,N_9384);
nand U9739 (N_9739,N_9476,N_8921);
and U9740 (N_9740,N_9092,N_9011);
nor U9741 (N_9741,N_8998,N_9403);
and U9742 (N_9742,N_9571,N_8884);
nor U9743 (N_9743,N_9270,N_8864);
nor U9744 (N_9744,N_9427,N_9417);
or U9745 (N_9745,N_9274,N_9329);
or U9746 (N_9746,N_9173,N_9405);
or U9747 (N_9747,N_9442,N_8898);
nand U9748 (N_9748,N_9239,N_9583);
nand U9749 (N_9749,N_8970,N_8805);
and U9750 (N_9750,N_9297,N_8881);
or U9751 (N_9751,N_9123,N_8997);
nor U9752 (N_9752,N_8914,N_9362);
nand U9753 (N_9753,N_9343,N_9302);
nand U9754 (N_9754,N_9597,N_8809);
nand U9755 (N_9755,N_9005,N_8988);
and U9756 (N_9756,N_9356,N_9246);
or U9757 (N_9757,N_9224,N_9101);
or U9758 (N_9758,N_9467,N_9566);
and U9759 (N_9759,N_9147,N_9293);
nor U9760 (N_9760,N_8964,N_9018);
or U9761 (N_9761,N_9106,N_9445);
nor U9762 (N_9762,N_8872,N_9307);
nand U9763 (N_9763,N_9324,N_9097);
nand U9764 (N_9764,N_8837,N_9034);
or U9765 (N_9765,N_8863,N_9500);
nand U9766 (N_9766,N_9487,N_9434);
nand U9767 (N_9767,N_8845,N_9514);
or U9768 (N_9768,N_9067,N_9040);
and U9769 (N_9769,N_8859,N_9535);
nand U9770 (N_9770,N_8978,N_9022);
and U9771 (N_9771,N_9475,N_9009);
nor U9772 (N_9772,N_8800,N_8951);
and U9773 (N_9773,N_9002,N_9141);
nor U9774 (N_9774,N_9266,N_9548);
or U9775 (N_9775,N_9083,N_9221);
or U9776 (N_9776,N_8915,N_9415);
nand U9777 (N_9777,N_9019,N_9592);
and U9778 (N_9778,N_9462,N_9429);
nand U9779 (N_9779,N_8966,N_8821);
and U9780 (N_9780,N_9194,N_9444);
or U9781 (N_9781,N_9109,N_8842);
and U9782 (N_9782,N_9206,N_9508);
or U9783 (N_9783,N_8955,N_9159);
nand U9784 (N_9784,N_9217,N_8812);
nand U9785 (N_9785,N_9051,N_9070);
nand U9786 (N_9786,N_8957,N_9484);
nand U9787 (N_9787,N_9534,N_9545);
nor U9788 (N_9788,N_9024,N_9091);
or U9789 (N_9789,N_9074,N_8808);
or U9790 (N_9790,N_9512,N_9061);
xnor U9791 (N_9791,N_9541,N_9025);
nor U9792 (N_9792,N_8950,N_8939);
and U9793 (N_9793,N_9021,N_8952);
nand U9794 (N_9794,N_9419,N_8862);
nand U9795 (N_9795,N_8814,N_9459);
xor U9796 (N_9796,N_9586,N_9498);
and U9797 (N_9797,N_9399,N_9549);
nand U9798 (N_9798,N_8871,N_8889);
nand U9799 (N_9799,N_9135,N_9590);
and U9800 (N_9800,N_9477,N_9020);
nor U9801 (N_9801,N_9389,N_9104);
nor U9802 (N_9802,N_8861,N_8853);
and U9803 (N_9803,N_9426,N_9252);
nand U9804 (N_9804,N_9280,N_8989);
or U9805 (N_9805,N_9353,N_8994);
and U9806 (N_9806,N_8985,N_8983);
nor U9807 (N_9807,N_9059,N_9189);
or U9808 (N_9808,N_9359,N_9550);
xor U9809 (N_9809,N_9491,N_8875);
and U9810 (N_9810,N_9049,N_9129);
nor U9811 (N_9811,N_9164,N_9490);
nand U9812 (N_9812,N_9085,N_9408);
or U9813 (N_9813,N_8996,N_9187);
nor U9814 (N_9814,N_9449,N_9068);
nand U9815 (N_9815,N_9179,N_9251);
nand U9816 (N_9816,N_9368,N_9226);
and U9817 (N_9817,N_9086,N_9306);
and U9818 (N_9818,N_9533,N_8896);
or U9819 (N_9819,N_9238,N_9420);
nand U9820 (N_9820,N_9290,N_9482);
or U9821 (N_9821,N_9553,N_9089);
nor U9822 (N_9822,N_9004,N_9041);
nand U9823 (N_9823,N_8979,N_8873);
or U9824 (N_9824,N_8897,N_8886);
or U9825 (N_9825,N_9272,N_8899);
or U9826 (N_9826,N_9492,N_9360);
and U9827 (N_9827,N_9184,N_8980);
nor U9828 (N_9828,N_9044,N_9406);
or U9829 (N_9829,N_9440,N_9443);
and U9830 (N_9830,N_9511,N_8803);
nor U9831 (N_9831,N_9126,N_8811);
xnor U9832 (N_9832,N_9198,N_8849);
or U9833 (N_9833,N_9481,N_9493);
nand U9834 (N_9834,N_8879,N_9473);
and U9835 (N_9835,N_8830,N_9410);
nor U9836 (N_9836,N_9335,N_9572);
and U9837 (N_9837,N_9480,N_8877);
nor U9838 (N_9838,N_8975,N_8977);
nor U9839 (N_9839,N_8991,N_9552);
nand U9840 (N_9840,N_9502,N_9499);
nand U9841 (N_9841,N_9301,N_9066);
or U9842 (N_9842,N_8965,N_9172);
or U9843 (N_9843,N_9207,N_9342);
or U9844 (N_9844,N_9322,N_8923);
nor U9845 (N_9845,N_9378,N_9100);
or U9846 (N_9846,N_9438,N_9396);
nand U9847 (N_9847,N_9315,N_8867);
and U9848 (N_9848,N_9264,N_8807);
or U9849 (N_9849,N_9537,N_8894);
nor U9850 (N_9850,N_9120,N_9520);
nand U9851 (N_9851,N_9271,N_8930);
or U9852 (N_9852,N_8933,N_9530);
nand U9853 (N_9853,N_9573,N_8828);
nor U9854 (N_9854,N_9222,N_9139);
xor U9855 (N_9855,N_9134,N_9218);
nor U9856 (N_9856,N_9075,N_8883);
nor U9857 (N_9857,N_9001,N_8820);
nand U9858 (N_9858,N_9132,N_8929);
or U9859 (N_9859,N_9433,N_9556);
nor U9860 (N_9860,N_9568,N_8833);
nand U9861 (N_9861,N_9407,N_9495);
nor U9862 (N_9862,N_9551,N_9351);
nor U9863 (N_9863,N_8895,N_9137);
nor U9864 (N_9864,N_9228,N_9313);
or U9865 (N_9865,N_8829,N_9210);
or U9866 (N_9866,N_9202,N_9316);
and U9867 (N_9867,N_9115,N_8948);
nor U9868 (N_9868,N_9008,N_9042);
nand U9869 (N_9869,N_9584,N_9527);
and U9870 (N_9870,N_9401,N_9254);
or U9871 (N_9871,N_8947,N_9412);
nor U9872 (N_9872,N_9546,N_9017);
and U9873 (N_9873,N_9245,N_9536);
nor U9874 (N_9874,N_9501,N_9562);
or U9875 (N_9875,N_9212,N_9201);
or U9876 (N_9876,N_8954,N_8937);
nor U9877 (N_9877,N_8953,N_8976);
or U9878 (N_9878,N_9599,N_9454);
and U9879 (N_9879,N_9268,N_9325);
or U9880 (N_9880,N_9240,N_9397);
nor U9881 (N_9881,N_9163,N_9052);
nand U9882 (N_9882,N_9062,N_8825);
nand U9883 (N_9883,N_9336,N_9367);
or U9884 (N_9884,N_9411,N_9326);
nor U9885 (N_9885,N_9372,N_9334);
nand U9886 (N_9886,N_9453,N_9157);
nand U9887 (N_9887,N_9485,N_9595);
nor U9888 (N_9888,N_9331,N_9072);
or U9889 (N_9889,N_9048,N_9295);
nand U9890 (N_9890,N_9028,N_9138);
and U9891 (N_9891,N_9255,N_8906);
or U9892 (N_9892,N_8885,N_9450);
nor U9893 (N_9893,N_9386,N_8858);
nand U9894 (N_9894,N_9304,N_9446);
or U9895 (N_9895,N_9394,N_9287);
nor U9896 (N_9896,N_9037,N_9369);
nor U9897 (N_9897,N_9064,N_9317);
nor U9898 (N_9898,N_9414,N_9554);
or U9899 (N_9899,N_9260,N_9497);
nand U9900 (N_9900,N_9363,N_9565);
nor U9901 (N_9901,N_9078,N_9585);
nand U9902 (N_9902,N_9103,N_8907);
nor U9903 (N_9903,N_9204,N_9435);
nor U9904 (N_9904,N_9472,N_9124);
or U9905 (N_9905,N_9349,N_9003);
and U9906 (N_9906,N_9432,N_8986);
and U9907 (N_9907,N_9436,N_9150);
or U9908 (N_9908,N_8924,N_8902);
nor U9909 (N_9909,N_8887,N_9291);
nor U9910 (N_9910,N_8984,N_9143);
and U9911 (N_9911,N_9096,N_9354);
and U9912 (N_9912,N_9314,N_8909);
or U9913 (N_9913,N_9515,N_9364);
nor U9914 (N_9914,N_8815,N_9333);
or U9915 (N_9915,N_9424,N_9175);
or U9916 (N_9916,N_9319,N_9125);
and U9917 (N_9917,N_9192,N_9460);
or U9918 (N_9918,N_8854,N_9241);
nor U9919 (N_9919,N_8936,N_9577);
or U9920 (N_9920,N_9347,N_9581);
or U9921 (N_9921,N_9195,N_8960);
nor U9922 (N_9922,N_9309,N_9361);
nand U9923 (N_9923,N_9298,N_8935);
or U9924 (N_9924,N_9542,N_9337);
nand U9925 (N_9925,N_9321,N_9155);
nor U9926 (N_9926,N_8993,N_8922);
or U9927 (N_9927,N_8971,N_9127);
nor U9928 (N_9928,N_9465,N_8824);
or U9929 (N_9929,N_9248,N_9409);
nand U9930 (N_9930,N_9350,N_9598);
and U9931 (N_9931,N_9188,N_9488);
and U9932 (N_9932,N_9451,N_9033);
or U9933 (N_9933,N_9524,N_9269);
and U9934 (N_9934,N_8904,N_8910);
and U9935 (N_9935,N_9261,N_9538);
nand U9936 (N_9936,N_8870,N_9540);
nand U9937 (N_9937,N_9102,N_9121);
nor U9938 (N_9938,N_8891,N_8973);
nor U9939 (N_9939,N_9090,N_9557);
nor U9940 (N_9940,N_9007,N_9077);
nand U9941 (N_9941,N_8802,N_9108);
nand U9942 (N_9942,N_9118,N_8968);
or U9943 (N_9943,N_9136,N_8818);
and U9944 (N_9944,N_8972,N_8855);
nor U9945 (N_9945,N_9282,N_9199);
nor U9946 (N_9946,N_8992,N_9080);
or U9947 (N_9947,N_9523,N_8961);
nand U9948 (N_9948,N_9471,N_9379);
nor U9949 (N_9949,N_9284,N_9006);
nor U9950 (N_9950,N_9544,N_9355);
and U9951 (N_9951,N_8832,N_9170);
nor U9952 (N_9952,N_8901,N_9344);
nand U9953 (N_9953,N_9010,N_8956);
and U9954 (N_9954,N_9478,N_9053);
and U9955 (N_9955,N_9197,N_9423);
or U9956 (N_9956,N_9211,N_9400);
or U9957 (N_9957,N_9489,N_8926);
nor U9958 (N_9958,N_9318,N_8893);
nand U9959 (N_9959,N_9496,N_9532);
and U9960 (N_9960,N_9168,N_8819);
nand U9961 (N_9961,N_8851,N_8959);
and U9962 (N_9962,N_9591,N_9032);
nor U9963 (N_9963,N_9276,N_9292);
nand U9964 (N_9964,N_8949,N_8816);
nor U9965 (N_9965,N_9219,N_8995);
or U9966 (N_9966,N_9494,N_9381);
and U9967 (N_9967,N_9474,N_9346);
nor U9968 (N_9968,N_9560,N_9107);
and U9969 (N_9969,N_9073,N_9038);
and U9970 (N_9970,N_9258,N_9575);
and U9971 (N_9971,N_9370,N_8974);
nand U9972 (N_9972,N_9071,N_9154);
or U9973 (N_9973,N_8826,N_9088);
and U9974 (N_9974,N_8917,N_9574);
nor U9975 (N_9975,N_9256,N_8810);
or U9976 (N_9976,N_8866,N_9464);
and U9977 (N_9977,N_8813,N_9587);
nand U9978 (N_9978,N_9582,N_9148);
nor U9979 (N_9979,N_9065,N_9504);
or U9980 (N_9980,N_9015,N_8958);
nor U9981 (N_9981,N_9516,N_9161);
nand U9982 (N_9982,N_9518,N_9391);
nand U9983 (N_9983,N_8835,N_9447);
nand U9984 (N_9984,N_9404,N_9174);
and U9985 (N_9985,N_9452,N_8999);
and U9986 (N_9986,N_9539,N_9130);
or U9987 (N_9987,N_9323,N_9128);
nand U9988 (N_9988,N_9330,N_8843);
or U9989 (N_9989,N_9247,N_9377);
and U9990 (N_9990,N_9185,N_9186);
and U9991 (N_9991,N_9352,N_9016);
nand U9992 (N_9992,N_9278,N_9054);
nor U9993 (N_9993,N_9569,N_9131);
or U9994 (N_9994,N_9232,N_9242);
or U9995 (N_9995,N_9119,N_9213);
nor U9996 (N_9996,N_9162,N_8806);
nand U9997 (N_9997,N_9338,N_9182);
nor U9998 (N_9998,N_9469,N_8987);
nand U9999 (N_9999,N_9229,N_9237);
nand U10000 (N_10000,N_9289,N_9075);
or U10001 (N_10001,N_9491,N_9170);
or U10002 (N_10002,N_9101,N_9400);
or U10003 (N_10003,N_9377,N_8877);
or U10004 (N_10004,N_9448,N_9097);
nand U10005 (N_10005,N_9026,N_9110);
or U10006 (N_10006,N_9041,N_9209);
nand U10007 (N_10007,N_9304,N_9062);
or U10008 (N_10008,N_8949,N_9376);
or U10009 (N_10009,N_8819,N_9365);
and U10010 (N_10010,N_8841,N_9195);
nor U10011 (N_10011,N_9142,N_8921);
and U10012 (N_10012,N_8990,N_8953);
and U10013 (N_10013,N_9146,N_8842);
nand U10014 (N_10014,N_9286,N_9575);
nor U10015 (N_10015,N_8883,N_9193);
or U10016 (N_10016,N_9187,N_8946);
or U10017 (N_10017,N_9072,N_9157);
nand U10018 (N_10018,N_8829,N_9247);
nor U10019 (N_10019,N_8937,N_9050);
nand U10020 (N_10020,N_8879,N_8941);
or U10021 (N_10021,N_9399,N_8890);
or U10022 (N_10022,N_9000,N_9020);
or U10023 (N_10023,N_9000,N_9444);
nor U10024 (N_10024,N_9550,N_8825);
nor U10025 (N_10025,N_9392,N_9097);
or U10026 (N_10026,N_9242,N_9479);
nand U10027 (N_10027,N_9428,N_8848);
nand U10028 (N_10028,N_9556,N_9552);
nor U10029 (N_10029,N_9156,N_9409);
nand U10030 (N_10030,N_8829,N_8974);
or U10031 (N_10031,N_8807,N_8843);
nand U10032 (N_10032,N_9591,N_9192);
nor U10033 (N_10033,N_9123,N_9497);
nor U10034 (N_10034,N_9392,N_8829);
or U10035 (N_10035,N_9129,N_9040);
or U10036 (N_10036,N_8958,N_9584);
and U10037 (N_10037,N_9499,N_9503);
or U10038 (N_10038,N_9161,N_9588);
nor U10039 (N_10039,N_8818,N_9540);
nand U10040 (N_10040,N_9461,N_9151);
nand U10041 (N_10041,N_9192,N_8817);
or U10042 (N_10042,N_9562,N_9067);
nor U10043 (N_10043,N_8925,N_9478);
nor U10044 (N_10044,N_8939,N_9134);
nand U10045 (N_10045,N_9262,N_9181);
and U10046 (N_10046,N_9217,N_9437);
or U10047 (N_10047,N_8986,N_8841);
and U10048 (N_10048,N_8911,N_9060);
nor U10049 (N_10049,N_8878,N_9599);
and U10050 (N_10050,N_8954,N_9090);
nor U10051 (N_10051,N_9371,N_9434);
nor U10052 (N_10052,N_9487,N_9559);
nand U10053 (N_10053,N_9488,N_8992);
nand U10054 (N_10054,N_8889,N_9051);
and U10055 (N_10055,N_9396,N_8956);
and U10056 (N_10056,N_9379,N_9321);
or U10057 (N_10057,N_8937,N_9375);
nor U10058 (N_10058,N_8817,N_9274);
and U10059 (N_10059,N_8851,N_9266);
nor U10060 (N_10060,N_9032,N_9202);
nor U10061 (N_10061,N_9278,N_9106);
or U10062 (N_10062,N_9051,N_9308);
nand U10063 (N_10063,N_9024,N_8950);
and U10064 (N_10064,N_9131,N_8816);
nor U10065 (N_10065,N_9145,N_9208);
nand U10066 (N_10066,N_8986,N_8859);
or U10067 (N_10067,N_9225,N_9117);
nor U10068 (N_10068,N_8800,N_9432);
nor U10069 (N_10069,N_8933,N_8930);
or U10070 (N_10070,N_8908,N_9014);
or U10071 (N_10071,N_9488,N_8966);
nand U10072 (N_10072,N_8994,N_9281);
nor U10073 (N_10073,N_8841,N_8869);
nand U10074 (N_10074,N_9191,N_9505);
and U10075 (N_10075,N_9389,N_8971);
or U10076 (N_10076,N_8944,N_9355);
nor U10077 (N_10077,N_8952,N_8907);
nand U10078 (N_10078,N_9012,N_9135);
or U10079 (N_10079,N_9512,N_8923);
and U10080 (N_10080,N_9540,N_9137);
nand U10081 (N_10081,N_9335,N_8852);
or U10082 (N_10082,N_8961,N_9083);
xnor U10083 (N_10083,N_9055,N_9563);
nand U10084 (N_10084,N_9598,N_8953);
and U10085 (N_10085,N_9395,N_9110);
or U10086 (N_10086,N_9382,N_8874);
or U10087 (N_10087,N_9025,N_9547);
nor U10088 (N_10088,N_8863,N_9522);
xnor U10089 (N_10089,N_8926,N_9573);
nand U10090 (N_10090,N_9029,N_9094);
nor U10091 (N_10091,N_9312,N_9542);
and U10092 (N_10092,N_9488,N_9437);
nand U10093 (N_10093,N_8948,N_9125);
or U10094 (N_10094,N_9527,N_9123);
nand U10095 (N_10095,N_9106,N_9146);
and U10096 (N_10096,N_8920,N_8972);
nor U10097 (N_10097,N_9370,N_9442);
nand U10098 (N_10098,N_8803,N_9524);
nor U10099 (N_10099,N_9317,N_9260);
or U10100 (N_10100,N_8846,N_9517);
nor U10101 (N_10101,N_9343,N_9044);
and U10102 (N_10102,N_9343,N_8895);
xnor U10103 (N_10103,N_9451,N_9585);
nand U10104 (N_10104,N_8890,N_9125);
and U10105 (N_10105,N_9127,N_9318);
nand U10106 (N_10106,N_8856,N_8853);
nand U10107 (N_10107,N_9152,N_9215);
nand U10108 (N_10108,N_9324,N_9238);
and U10109 (N_10109,N_8991,N_9406);
and U10110 (N_10110,N_9457,N_8863);
and U10111 (N_10111,N_9181,N_9441);
nand U10112 (N_10112,N_9288,N_8907);
nand U10113 (N_10113,N_9548,N_8867);
nor U10114 (N_10114,N_9358,N_9485);
nor U10115 (N_10115,N_8800,N_9338);
nand U10116 (N_10116,N_8951,N_9317);
and U10117 (N_10117,N_9354,N_9310);
nand U10118 (N_10118,N_9323,N_9535);
nor U10119 (N_10119,N_8841,N_9023);
nor U10120 (N_10120,N_9106,N_9088);
nor U10121 (N_10121,N_8883,N_9572);
and U10122 (N_10122,N_9497,N_9042);
nand U10123 (N_10123,N_8929,N_9116);
nor U10124 (N_10124,N_8810,N_8950);
nor U10125 (N_10125,N_9352,N_9522);
or U10126 (N_10126,N_9476,N_9345);
and U10127 (N_10127,N_9197,N_9070);
and U10128 (N_10128,N_9209,N_8835);
nand U10129 (N_10129,N_8978,N_9452);
nand U10130 (N_10130,N_9142,N_9285);
nand U10131 (N_10131,N_9360,N_9268);
nor U10132 (N_10132,N_9587,N_9558);
nand U10133 (N_10133,N_9291,N_9086);
nor U10134 (N_10134,N_9510,N_8944);
xnor U10135 (N_10135,N_9332,N_9145);
or U10136 (N_10136,N_9289,N_9586);
or U10137 (N_10137,N_9577,N_9265);
nand U10138 (N_10138,N_9180,N_9173);
or U10139 (N_10139,N_9528,N_8889);
nand U10140 (N_10140,N_9070,N_8800);
and U10141 (N_10141,N_9398,N_9370);
and U10142 (N_10142,N_9174,N_9565);
and U10143 (N_10143,N_9110,N_9253);
and U10144 (N_10144,N_9440,N_9541);
and U10145 (N_10145,N_9023,N_9166);
nand U10146 (N_10146,N_8837,N_9567);
nor U10147 (N_10147,N_8855,N_9435);
and U10148 (N_10148,N_9596,N_9393);
and U10149 (N_10149,N_8833,N_9558);
and U10150 (N_10150,N_9429,N_9508);
and U10151 (N_10151,N_9571,N_9022);
or U10152 (N_10152,N_9479,N_9484);
and U10153 (N_10153,N_9400,N_9337);
or U10154 (N_10154,N_9308,N_9275);
and U10155 (N_10155,N_8805,N_9072);
nor U10156 (N_10156,N_9537,N_9385);
nor U10157 (N_10157,N_9178,N_9174);
nand U10158 (N_10158,N_9451,N_8912);
nor U10159 (N_10159,N_8987,N_9572);
nand U10160 (N_10160,N_9238,N_9297);
or U10161 (N_10161,N_9567,N_8961);
or U10162 (N_10162,N_9271,N_9513);
or U10163 (N_10163,N_9280,N_9159);
nand U10164 (N_10164,N_8959,N_9593);
and U10165 (N_10165,N_9022,N_9360);
or U10166 (N_10166,N_9311,N_9124);
or U10167 (N_10167,N_9566,N_8823);
nor U10168 (N_10168,N_9158,N_9480);
or U10169 (N_10169,N_9205,N_9426);
and U10170 (N_10170,N_9182,N_9234);
or U10171 (N_10171,N_9510,N_9481);
or U10172 (N_10172,N_9225,N_9095);
or U10173 (N_10173,N_8940,N_8962);
or U10174 (N_10174,N_9344,N_9133);
or U10175 (N_10175,N_8965,N_9545);
nand U10176 (N_10176,N_9322,N_9168);
nor U10177 (N_10177,N_8803,N_9175);
or U10178 (N_10178,N_9302,N_8983);
or U10179 (N_10179,N_9453,N_9278);
nor U10180 (N_10180,N_8821,N_8921);
nor U10181 (N_10181,N_9291,N_9460);
nor U10182 (N_10182,N_9198,N_9430);
nor U10183 (N_10183,N_8851,N_9536);
nor U10184 (N_10184,N_8907,N_9555);
and U10185 (N_10185,N_8922,N_9261);
nand U10186 (N_10186,N_9242,N_9129);
or U10187 (N_10187,N_9233,N_9265);
nor U10188 (N_10188,N_9304,N_9031);
nor U10189 (N_10189,N_9097,N_8922);
or U10190 (N_10190,N_8816,N_9213);
and U10191 (N_10191,N_8965,N_8809);
nor U10192 (N_10192,N_8995,N_9410);
or U10193 (N_10193,N_8857,N_9555);
nand U10194 (N_10194,N_9587,N_9407);
and U10195 (N_10195,N_9384,N_9322);
or U10196 (N_10196,N_9103,N_9361);
or U10197 (N_10197,N_9493,N_9516);
nand U10198 (N_10198,N_9395,N_9588);
or U10199 (N_10199,N_9377,N_8846);
nand U10200 (N_10200,N_9022,N_9334);
or U10201 (N_10201,N_9209,N_8897);
or U10202 (N_10202,N_9363,N_9594);
or U10203 (N_10203,N_9321,N_9573);
nand U10204 (N_10204,N_9328,N_9355);
and U10205 (N_10205,N_9303,N_9235);
and U10206 (N_10206,N_9019,N_9052);
nand U10207 (N_10207,N_9146,N_8816);
or U10208 (N_10208,N_9294,N_8826);
nor U10209 (N_10209,N_9140,N_9045);
nand U10210 (N_10210,N_9574,N_9386);
nand U10211 (N_10211,N_8989,N_9596);
or U10212 (N_10212,N_9506,N_8959);
nor U10213 (N_10213,N_9544,N_8843);
and U10214 (N_10214,N_8974,N_9478);
nand U10215 (N_10215,N_9008,N_9453);
nor U10216 (N_10216,N_9127,N_9494);
or U10217 (N_10217,N_8934,N_9030);
nand U10218 (N_10218,N_8926,N_9579);
and U10219 (N_10219,N_8931,N_9332);
nand U10220 (N_10220,N_9207,N_8934);
nand U10221 (N_10221,N_8968,N_9507);
or U10222 (N_10222,N_9571,N_8966);
nor U10223 (N_10223,N_8881,N_9028);
nor U10224 (N_10224,N_9453,N_9524);
and U10225 (N_10225,N_9068,N_9434);
nor U10226 (N_10226,N_9490,N_9027);
nand U10227 (N_10227,N_9483,N_8814);
nor U10228 (N_10228,N_9116,N_9337);
nand U10229 (N_10229,N_9441,N_9175);
or U10230 (N_10230,N_9037,N_9113);
nor U10231 (N_10231,N_9005,N_8838);
and U10232 (N_10232,N_8829,N_9432);
or U10233 (N_10233,N_9444,N_9001);
nand U10234 (N_10234,N_9238,N_9054);
nand U10235 (N_10235,N_9303,N_8884);
nand U10236 (N_10236,N_8877,N_8812);
nand U10237 (N_10237,N_8830,N_8802);
and U10238 (N_10238,N_9371,N_9336);
and U10239 (N_10239,N_8886,N_9026);
or U10240 (N_10240,N_9221,N_9021);
and U10241 (N_10241,N_8921,N_8816);
nand U10242 (N_10242,N_9041,N_8864);
nor U10243 (N_10243,N_9382,N_9376);
nor U10244 (N_10244,N_9463,N_9108);
and U10245 (N_10245,N_9583,N_9159);
nand U10246 (N_10246,N_9306,N_8822);
nor U10247 (N_10247,N_9104,N_9257);
or U10248 (N_10248,N_8849,N_8833);
or U10249 (N_10249,N_9005,N_9479);
or U10250 (N_10250,N_9495,N_9595);
and U10251 (N_10251,N_9527,N_9505);
or U10252 (N_10252,N_9564,N_8830);
and U10253 (N_10253,N_9546,N_9292);
and U10254 (N_10254,N_9102,N_9582);
nand U10255 (N_10255,N_9271,N_9241);
or U10256 (N_10256,N_8978,N_9570);
nor U10257 (N_10257,N_9060,N_9415);
or U10258 (N_10258,N_9427,N_9414);
or U10259 (N_10259,N_8814,N_9479);
nor U10260 (N_10260,N_9415,N_8983);
nor U10261 (N_10261,N_9046,N_8874);
nand U10262 (N_10262,N_9324,N_8876);
or U10263 (N_10263,N_9568,N_9470);
nor U10264 (N_10264,N_9259,N_8812);
and U10265 (N_10265,N_8877,N_8931);
nand U10266 (N_10266,N_9088,N_8856);
and U10267 (N_10267,N_9110,N_8947);
nor U10268 (N_10268,N_9349,N_9363);
nor U10269 (N_10269,N_8916,N_9151);
nor U10270 (N_10270,N_9160,N_9185);
nor U10271 (N_10271,N_9360,N_9468);
or U10272 (N_10272,N_9045,N_9151);
nor U10273 (N_10273,N_9208,N_9559);
or U10274 (N_10274,N_9267,N_9306);
nor U10275 (N_10275,N_9394,N_8914);
and U10276 (N_10276,N_9525,N_9383);
nand U10277 (N_10277,N_9179,N_9529);
nand U10278 (N_10278,N_9163,N_9226);
or U10279 (N_10279,N_9319,N_9334);
nor U10280 (N_10280,N_8880,N_9292);
nor U10281 (N_10281,N_8835,N_9241);
or U10282 (N_10282,N_9164,N_9429);
or U10283 (N_10283,N_8816,N_9250);
or U10284 (N_10284,N_9280,N_9346);
nand U10285 (N_10285,N_9380,N_9569);
nand U10286 (N_10286,N_9315,N_9273);
nor U10287 (N_10287,N_9035,N_8928);
or U10288 (N_10288,N_9332,N_9367);
or U10289 (N_10289,N_9471,N_9469);
or U10290 (N_10290,N_9520,N_9512);
and U10291 (N_10291,N_8991,N_9215);
nand U10292 (N_10292,N_9499,N_8835);
or U10293 (N_10293,N_9361,N_8873);
or U10294 (N_10294,N_9338,N_8883);
and U10295 (N_10295,N_9427,N_8845);
nand U10296 (N_10296,N_9161,N_9567);
nor U10297 (N_10297,N_9291,N_9142);
or U10298 (N_10298,N_9588,N_9511);
nor U10299 (N_10299,N_9280,N_9458);
and U10300 (N_10300,N_9129,N_8992);
nor U10301 (N_10301,N_8832,N_9292);
nand U10302 (N_10302,N_9161,N_9424);
nor U10303 (N_10303,N_9069,N_9271);
nor U10304 (N_10304,N_8858,N_8901);
xnor U10305 (N_10305,N_9244,N_8966);
nor U10306 (N_10306,N_9415,N_9350);
nand U10307 (N_10307,N_8925,N_9120);
nand U10308 (N_10308,N_9360,N_9579);
nor U10309 (N_10309,N_9521,N_9233);
nand U10310 (N_10310,N_8898,N_9446);
nand U10311 (N_10311,N_9202,N_8888);
and U10312 (N_10312,N_9594,N_9503);
nor U10313 (N_10313,N_9522,N_9321);
nor U10314 (N_10314,N_9087,N_8968);
and U10315 (N_10315,N_8930,N_8859);
and U10316 (N_10316,N_8865,N_9159);
nor U10317 (N_10317,N_9067,N_9011);
nand U10318 (N_10318,N_9505,N_9072);
or U10319 (N_10319,N_9041,N_9546);
nand U10320 (N_10320,N_8926,N_9501);
nand U10321 (N_10321,N_9282,N_9437);
nand U10322 (N_10322,N_9096,N_9552);
nor U10323 (N_10323,N_9189,N_8946);
xor U10324 (N_10324,N_9243,N_8938);
nor U10325 (N_10325,N_9046,N_9440);
or U10326 (N_10326,N_9346,N_9294);
nand U10327 (N_10327,N_8913,N_9300);
and U10328 (N_10328,N_9341,N_9315);
and U10329 (N_10329,N_9376,N_9313);
and U10330 (N_10330,N_8998,N_9414);
and U10331 (N_10331,N_9134,N_9075);
nand U10332 (N_10332,N_9016,N_9571);
nor U10333 (N_10333,N_8855,N_9468);
or U10334 (N_10334,N_9230,N_9304);
or U10335 (N_10335,N_9450,N_9331);
and U10336 (N_10336,N_9251,N_8862);
nor U10337 (N_10337,N_8936,N_9472);
nand U10338 (N_10338,N_9245,N_9330);
or U10339 (N_10339,N_9025,N_9497);
and U10340 (N_10340,N_9232,N_9054);
or U10341 (N_10341,N_9270,N_9417);
nand U10342 (N_10342,N_8864,N_9322);
nor U10343 (N_10343,N_9547,N_8930);
or U10344 (N_10344,N_8998,N_8943);
nand U10345 (N_10345,N_9415,N_9435);
and U10346 (N_10346,N_9311,N_9037);
nand U10347 (N_10347,N_9037,N_9443);
nor U10348 (N_10348,N_9119,N_8926);
or U10349 (N_10349,N_9221,N_9464);
nor U10350 (N_10350,N_9508,N_9147);
or U10351 (N_10351,N_9520,N_9208);
and U10352 (N_10352,N_9533,N_9456);
or U10353 (N_10353,N_9428,N_8983);
and U10354 (N_10354,N_9354,N_8816);
or U10355 (N_10355,N_9199,N_9034);
and U10356 (N_10356,N_9597,N_9168);
or U10357 (N_10357,N_8986,N_9099);
nor U10358 (N_10358,N_8920,N_9326);
and U10359 (N_10359,N_9500,N_9049);
or U10360 (N_10360,N_9408,N_8869);
nor U10361 (N_10361,N_9317,N_8816);
nor U10362 (N_10362,N_9038,N_8803);
nand U10363 (N_10363,N_9099,N_9142);
and U10364 (N_10364,N_9191,N_9278);
or U10365 (N_10365,N_9112,N_8814);
or U10366 (N_10366,N_9197,N_9372);
nand U10367 (N_10367,N_9378,N_9589);
nand U10368 (N_10368,N_8913,N_9054);
nand U10369 (N_10369,N_8856,N_9186);
or U10370 (N_10370,N_9536,N_9080);
or U10371 (N_10371,N_9235,N_9130);
nand U10372 (N_10372,N_8914,N_9510);
and U10373 (N_10373,N_9598,N_9090);
nor U10374 (N_10374,N_9488,N_8935);
nor U10375 (N_10375,N_9079,N_9361);
and U10376 (N_10376,N_9209,N_9568);
or U10377 (N_10377,N_9104,N_8802);
nor U10378 (N_10378,N_8885,N_9027);
or U10379 (N_10379,N_8801,N_9415);
and U10380 (N_10380,N_8878,N_9448);
nand U10381 (N_10381,N_9167,N_9050);
or U10382 (N_10382,N_9219,N_8845);
xnor U10383 (N_10383,N_9059,N_9478);
xor U10384 (N_10384,N_8820,N_8889);
nor U10385 (N_10385,N_9279,N_8970);
nand U10386 (N_10386,N_9240,N_9247);
and U10387 (N_10387,N_9403,N_8828);
or U10388 (N_10388,N_8885,N_9554);
xnor U10389 (N_10389,N_9534,N_8946);
nand U10390 (N_10390,N_9220,N_9236);
nand U10391 (N_10391,N_8858,N_8834);
and U10392 (N_10392,N_9142,N_9072);
and U10393 (N_10393,N_8877,N_9417);
or U10394 (N_10394,N_9064,N_9082);
nor U10395 (N_10395,N_8858,N_9512);
and U10396 (N_10396,N_8957,N_8937);
nor U10397 (N_10397,N_8865,N_8812);
or U10398 (N_10398,N_9105,N_8935);
and U10399 (N_10399,N_9526,N_9107);
nand U10400 (N_10400,N_10014,N_9812);
and U10401 (N_10401,N_9660,N_10087);
or U10402 (N_10402,N_10046,N_9750);
nor U10403 (N_10403,N_10126,N_9794);
nand U10404 (N_10404,N_9627,N_9986);
or U10405 (N_10405,N_10124,N_9670);
and U10406 (N_10406,N_9741,N_9976);
and U10407 (N_10407,N_9601,N_9692);
nor U10408 (N_10408,N_10093,N_9697);
and U10409 (N_10409,N_9846,N_10231);
and U10410 (N_10410,N_10163,N_9819);
or U10411 (N_10411,N_9798,N_9771);
or U10412 (N_10412,N_10133,N_10265);
and U10413 (N_10413,N_10106,N_9821);
nor U10414 (N_10414,N_10396,N_9769);
nor U10415 (N_10415,N_9664,N_9895);
or U10416 (N_10416,N_10395,N_10032);
or U10417 (N_10417,N_10342,N_10274);
or U10418 (N_10418,N_10000,N_10140);
nor U10419 (N_10419,N_10115,N_10155);
and U10420 (N_10420,N_9773,N_9731);
and U10421 (N_10421,N_10359,N_9892);
or U10422 (N_10422,N_9837,N_10393);
nand U10423 (N_10423,N_9925,N_10058);
nor U10424 (N_10424,N_9968,N_9981);
and U10425 (N_10425,N_10364,N_9728);
or U10426 (N_10426,N_9839,N_10294);
nor U10427 (N_10427,N_9642,N_9916);
or U10428 (N_10428,N_10045,N_10011);
or U10429 (N_10429,N_10209,N_10268);
nand U10430 (N_10430,N_10034,N_9753);
nor U10431 (N_10431,N_9807,N_10311);
nand U10432 (N_10432,N_9855,N_10355);
nor U10433 (N_10433,N_10105,N_9865);
nor U10434 (N_10434,N_10097,N_9860);
nor U10435 (N_10435,N_9978,N_9936);
or U10436 (N_10436,N_10366,N_9985);
nor U10437 (N_10437,N_10280,N_10299);
nor U10438 (N_10438,N_10263,N_9840);
nand U10439 (N_10439,N_9784,N_9828);
and U10440 (N_10440,N_10232,N_10139);
nor U10441 (N_10441,N_9949,N_10306);
nor U10442 (N_10442,N_9674,N_10394);
or U10443 (N_10443,N_10287,N_10205);
or U10444 (N_10444,N_10259,N_10301);
or U10445 (N_10445,N_10135,N_9706);
or U10446 (N_10446,N_9783,N_9747);
nor U10447 (N_10447,N_9772,N_10138);
or U10448 (N_10448,N_9662,N_10346);
and U10449 (N_10449,N_9938,N_10273);
or U10450 (N_10450,N_9922,N_9680);
and U10451 (N_10451,N_9845,N_9804);
or U10452 (N_10452,N_10389,N_10201);
and U10453 (N_10453,N_9953,N_10196);
or U10454 (N_10454,N_9797,N_9805);
or U10455 (N_10455,N_10085,N_10033);
or U10456 (N_10456,N_10345,N_10023);
nand U10457 (N_10457,N_9746,N_9713);
and U10458 (N_10458,N_9881,N_9708);
nand U10459 (N_10459,N_10242,N_9714);
nor U10460 (N_10460,N_9999,N_9625);
and U10461 (N_10461,N_9904,N_10318);
nor U10462 (N_10462,N_9740,N_9796);
nor U10463 (N_10463,N_10068,N_9979);
or U10464 (N_10464,N_9816,N_10251);
and U10465 (N_10465,N_10199,N_10052);
or U10466 (N_10466,N_10312,N_9624);
or U10467 (N_10467,N_9770,N_10384);
nand U10468 (N_10468,N_10379,N_10088);
and U10469 (N_10469,N_9879,N_9826);
nor U10470 (N_10470,N_10308,N_10149);
or U10471 (N_10471,N_10307,N_10164);
or U10472 (N_10472,N_9891,N_10099);
nor U10473 (N_10473,N_9867,N_10237);
nor U10474 (N_10474,N_10264,N_9951);
or U10475 (N_10475,N_10378,N_10116);
or U10476 (N_10476,N_9665,N_10020);
or U10477 (N_10477,N_10367,N_9945);
nand U10478 (N_10478,N_10112,N_9975);
or U10479 (N_10479,N_10129,N_9727);
nand U10480 (N_10480,N_9899,N_9822);
nand U10481 (N_10481,N_10398,N_9734);
nand U10482 (N_10482,N_10275,N_9795);
or U10483 (N_10483,N_10110,N_9633);
and U10484 (N_10484,N_9813,N_10072);
or U10485 (N_10485,N_10212,N_10240);
or U10486 (N_10486,N_9872,N_9868);
and U10487 (N_10487,N_9913,N_10376);
or U10488 (N_10488,N_10360,N_10067);
nand U10489 (N_10489,N_10385,N_9641);
nor U10490 (N_10490,N_9782,N_10244);
nand U10491 (N_10491,N_9907,N_9705);
nor U10492 (N_10492,N_10066,N_9838);
and U10493 (N_10493,N_9785,N_9956);
nor U10494 (N_10494,N_9737,N_10333);
and U10495 (N_10495,N_10041,N_9668);
nand U10496 (N_10496,N_10062,N_10122);
and U10497 (N_10497,N_10141,N_9751);
nor U10498 (N_10498,N_9995,N_10048);
and U10499 (N_10499,N_9910,N_9791);
or U10500 (N_10500,N_9693,N_10162);
nand U10501 (N_10501,N_9932,N_9656);
and U10502 (N_10502,N_9876,N_10156);
or U10503 (N_10503,N_9924,N_10356);
and U10504 (N_10504,N_9823,N_10173);
nand U10505 (N_10505,N_9767,N_9946);
or U10506 (N_10506,N_10368,N_9632);
or U10507 (N_10507,N_10026,N_10094);
or U10508 (N_10508,N_9612,N_9882);
nor U10509 (N_10509,N_10323,N_10276);
and U10510 (N_10510,N_9998,N_9906);
or U10511 (N_10511,N_9997,N_10193);
nand U10512 (N_10512,N_9960,N_9929);
nor U10513 (N_10513,N_9818,N_9919);
and U10514 (N_10514,N_9673,N_10377);
nor U10515 (N_10515,N_10297,N_10184);
or U10516 (N_10516,N_10006,N_9690);
or U10517 (N_10517,N_10331,N_10392);
and U10518 (N_10518,N_10257,N_9610);
nor U10519 (N_10519,N_10100,N_10019);
and U10520 (N_10520,N_9649,N_10061);
and U10521 (N_10521,N_10245,N_9704);
nand U10522 (N_10522,N_10107,N_9948);
nand U10523 (N_10523,N_10283,N_9659);
nor U10524 (N_10524,N_10317,N_10049);
or U10525 (N_10525,N_9984,N_9699);
and U10526 (N_10526,N_9712,N_10296);
and U10527 (N_10527,N_9736,N_10031);
nand U10528 (N_10528,N_10387,N_9763);
and U10529 (N_10529,N_10008,N_10286);
and U10530 (N_10530,N_9871,N_10213);
nor U10531 (N_10531,N_9824,N_9715);
and U10532 (N_10532,N_9644,N_9702);
nand U10533 (N_10533,N_9792,N_10350);
nand U10534 (N_10534,N_10198,N_10347);
or U10535 (N_10535,N_10260,N_10153);
nor U10536 (N_10536,N_10103,N_10170);
nor U10537 (N_10537,N_9639,N_9917);
xnor U10538 (N_10538,N_9918,N_9745);
nand U10539 (N_10539,N_9732,N_10182);
and U10540 (N_10540,N_9756,N_10168);
and U10541 (N_10541,N_9663,N_10277);
nor U10542 (N_10542,N_9793,N_9754);
xnor U10543 (N_10543,N_10329,N_10254);
and U10544 (N_10544,N_9703,N_10223);
nor U10545 (N_10545,N_9902,N_9829);
or U10546 (N_10546,N_10055,N_10222);
or U10547 (N_10547,N_10202,N_10285);
nand U10548 (N_10548,N_9908,N_10039);
nand U10549 (N_10549,N_10160,N_9629);
nand U10550 (N_10550,N_10047,N_9602);
nor U10551 (N_10551,N_9789,N_9615);
or U10552 (N_10552,N_10130,N_9875);
or U10553 (N_10553,N_9779,N_10091);
nor U10554 (N_10554,N_9677,N_10185);
or U10555 (N_10555,N_9808,N_10146);
nand U10556 (N_10556,N_9764,N_10382);
or U10557 (N_10557,N_10217,N_10148);
and U10558 (N_10558,N_9730,N_10399);
or U10559 (N_10559,N_10235,N_9806);
nand U10560 (N_10560,N_10166,N_10365);
and U10561 (N_10561,N_9983,N_9643);
and U10562 (N_10562,N_9890,N_10239);
or U10563 (N_10563,N_9803,N_9722);
nor U10564 (N_10564,N_9901,N_9992);
nor U10565 (N_10565,N_9810,N_10113);
or U10566 (N_10566,N_10069,N_10241);
or U10567 (N_10567,N_9990,N_9896);
nor U10568 (N_10568,N_10390,N_9646);
or U10569 (N_10569,N_10021,N_9889);
and U10570 (N_10570,N_9980,N_9762);
and U10571 (N_10571,N_9832,N_9851);
and U10572 (N_10572,N_10255,N_9774);
nand U10573 (N_10573,N_10261,N_10322);
or U10574 (N_10574,N_10150,N_9676);
or U10575 (N_10575,N_9620,N_10349);
and U10576 (N_10576,N_10188,N_10338);
nand U10577 (N_10577,N_10336,N_9790);
nand U10578 (N_10578,N_10016,N_10229);
nand U10579 (N_10579,N_9743,N_9850);
nor U10580 (N_10580,N_10314,N_10298);
and U10581 (N_10581,N_10279,N_9631);
nand U10582 (N_10582,N_10340,N_10248);
nor U10583 (N_10583,N_10370,N_9653);
or U10584 (N_10584,N_10042,N_9827);
or U10585 (N_10585,N_10071,N_9621);
and U10586 (N_10586,N_10270,N_10226);
and U10587 (N_10587,N_10343,N_9927);
or U10588 (N_10588,N_9723,N_10079);
nand U10589 (N_10589,N_10169,N_9963);
nand U10590 (N_10590,N_10120,N_10262);
nand U10591 (N_10591,N_9903,N_9954);
nor U10592 (N_10592,N_9761,N_9849);
nand U10593 (N_10593,N_10300,N_10027);
or U10594 (N_10594,N_10330,N_9898);
or U10595 (N_10595,N_9964,N_10288);
nor U10596 (N_10596,N_9930,N_9859);
and U10597 (N_10597,N_10218,N_9969);
nor U10598 (N_10598,N_10167,N_10118);
nor U10599 (N_10599,N_10386,N_10373);
nand U10600 (N_10600,N_10313,N_9884);
nand U10601 (N_10601,N_9669,N_9683);
nor U10602 (N_10602,N_10337,N_10125);
nand U10603 (N_10603,N_9847,N_9623);
and U10604 (N_10604,N_10065,N_10197);
nor U10605 (N_10605,N_9658,N_9700);
and U10606 (N_10606,N_9603,N_10295);
or U10607 (N_10607,N_9637,N_9675);
or U10608 (N_10608,N_9921,N_10243);
or U10609 (N_10609,N_10190,N_10293);
nand U10610 (N_10610,N_9993,N_10381);
or U10611 (N_10611,N_9967,N_9719);
and U10612 (N_10612,N_10136,N_9970);
nor U10613 (N_10613,N_10073,N_10098);
and U10614 (N_10614,N_9681,N_10004);
nand U10615 (N_10615,N_9834,N_10075);
nor U10616 (N_10616,N_9941,N_9848);
and U10617 (N_10617,N_10070,N_9650);
xor U10618 (N_10618,N_9893,N_10187);
or U10619 (N_10619,N_9966,N_10175);
nand U10620 (N_10620,N_9880,N_9852);
or U10621 (N_10621,N_10001,N_9815);
and U10622 (N_10622,N_10238,N_9611);
or U10623 (N_10623,N_10192,N_10171);
xnor U10624 (N_10624,N_10204,N_9934);
or U10625 (N_10625,N_9836,N_10134);
or U10626 (N_10626,N_9900,N_10018);
nor U10627 (N_10627,N_9869,N_9940);
and U10628 (N_10628,N_10210,N_10194);
and U10629 (N_10629,N_9781,N_9842);
and U10630 (N_10630,N_9757,N_9710);
nor U10631 (N_10631,N_10357,N_10207);
or U10632 (N_10632,N_10005,N_9857);
or U10633 (N_10633,N_9691,N_10221);
nand U10634 (N_10634,N_10059,N_10127);
or U10635 (N_10635,N_9698,N_9635);
nor U10636 (N_10636,N_10082,N_10056);
nand U10637 (N_10637,N_10374,N_10319);
and U10638 (N_10638,N_10253,N_10081);
nor U10639 (N_10639,N_10083,N_10315);
nor U10640 (N_10640,N_9802,N_10095);
and U10641 (N_10641,N_9996,N_10054);
nand U10642 (N_10642,N_9614,N_10267);
or U10643 (N_10643,N_10363,N_9942);
and U10644 (N_10644,N_9748,N_10179);
or U10645 (N_10645,N_10353,N_9853);
or U10646 (N_10646,N_10158,N_10348);
nand U10647 (N_10647,N_9630,N_10302);
or U10648 (N_10648,N_9701,N_10024);
nand U10649 (N_10649,N_9923,N_10089);
nor U10650 (N_10650,N_10246,N_9778);
nand U10651 (N_10651,N_10358,N_10284);
nor U10652 (N_10652,N_10015,N_9989);
and U10653 (N_10653,N_9777,N_10316);
nand U10654 (N_10654,N_9817,N_10101);
and U10655 (N_10655,N_10208,N_10269);
and U10656 (N_10656,N_9870,N_10214);
nor U10657 (N_10657,N_10375,N_9688);
nor U10658 (N_10658,N_9655,N_9952);
and U10659 (N_10659,N_9878,N_10352);
or U10660 (N_10660,N_9752,N_9651);
and U10661 (N_10661,N_10211,N_10152);
xnor U10662 (N_10662,N_10290,N_9717);
nand U10663 (N_10663,N_9856,N_9830);
or U10664 (N_10664,N_9607,N_10328);
nor U10665 (N_10665,N_9667,N_10064);
or U10666 (N_10666,N_10178,N_10249);
and U10667 (N_10667,N_10111,N_10234);
and U10668 (N_10668,N_10086,N_10077);
and U10669 (N_10669,N_9962,N_10326);
nand U10670 (N_10670,N_9886,N_10104);
and U10671 (N_10671,N_10050,N_10177);
and U10672 (N_10672,N_10305,N_9866);
or U10673 (N_10673,N_9689,N_10228);
and U10674 (N_10674,N_9605,N_9931);
and U10675 (N_10675,N_9666,N_10051);
nor U10676 (N_10676,N_9638,N_9760);
and U10677 (N_10677,N_9652,N_9874);
and U10678 (N_10678,N_9686,N_9742);
and U10679 (N_10679,N_9622,N_9634);
nand U10680 (N_10680,N_10183,N_9716);
nand U10681 (N_10681,N_9672,N_10161);
and U10682 (N_10682,N_9786,N_10131);
nand U10683 (N_10683,N_9831,N_9604);
nor U10684 (N_10684,N_9987,N_10040);
nand U10685 (N_10685,N_10036,N_10022);
and U10686 (N_10686,N_9654,N_10151);
nand U10687 (N_10687,N_10191,N_9885);
nor U10688 (N_10688,N_9864,N_9613);
or U10689 (N_10689,N_10203,N_10074);
nor U10690 (N_10690,N_10080,N_10291);
or U10691 (N_10691,N_9657,N_9640);
nor U10692 (N_10692,N_10186,N_10137);
nand U10693 (N_10693,N_9974,N_10289);
or U10694 (N_10694,N_9800,N_10303);
nand U10695 (N_10695,N_10320,N_10383);
nor U10696 (N_10696,N_9991,N_10334);
and U10697 (N_10697,N_10002,N_10266);
and U10698 (N_10698,N_9618,N_9729);
nor U10699 (N_10699,N_9726,N_9811);
xnor U10700 (N_10700,N_10195,N_9994);
nor U10701 (N_10701,N_9617,N_9711);
or U10702 (N_10702,N_9733,N_9833);
or U10703 (N_10703,N_10391,N_10339);
and U10704 (N_10704,N_9694,N_10224);
or U10705 (N_10705,N_9724,N_10076);
or U10706 (N_10706,N_10282,N_10325);
and U10707 (N_10707,N_10341,N_9765);
nor U10708 (N_10708,N_10114,N_10258);
nand U10709 (N_10709,N_9950,N_10354);
nor U10710 (N_10710,N_10225,N_10159);
nor U10711 (N_10711,N_9609,N_9973);
and U10712 (N_10712,N_10057,N_9861);
nand U10713 (N_10713,N_10078,N_9707);
and U10714 (N_10714,N_10200,N_9947);
nor U10715 (N_10715,N_10037,N_10092);
and U10716 (N_10716,N_9648,N_9883);
and U10717 (N_10717,N_10121,N_9768);
nand U10718 (N_10718,N_9738,N_10230);
nor U10719 (N_10719,N_9758,N_9933);
or U10720 (N_10720,N_9911,N_9920);
nor U10721 (N_10721,N_9671,N_9626);
or U10722 (N_10722,N_9720,N_10335);
or U10723 (N_10723,N_9854,N_10216);
nand U10724 (N_10724,N_9943,N_9606);
xor U10725 (N_10725,N_10053,N_10028);
or U10726 (N_10726,N_9725,N_10176);
nor U10727 (N_10727,N_10017,N_9647);
nand U10728 (N_10728,N_9971,N_10119);
or U10729 (N_10729,N_10250,N_9958);
nor U10730 (N_10730,N_9961,N_9695);
or U10731 (N_10731,N_9739,N_9939);
nor U10732 (N_10732,N_10351,N_10292);
and U10733 (N_10733,N_10371,N_10108);
or U10734 (N_10734,N_9678,N_10215);
and U10735 (N_10735,N_9843,N_10344);
nand U10736 (N_10736,N_10063,N_10043);
nor U10737 (N_10737,N_10144,N_9928);
nor U10738 (N_10738,N_9759,N_10324);
and U10739 (N_10739,N_9835,N_9600);
nor U10740 (N_10740,N_9888,N_9862);
nor U10741 (N_10741,N_9935,N_10145);
nor U10742 (N_10742,N_9814,N_9776);
nand U10743 (N_10743,N_9863,N_9957);
nor U10744 (N_10744,N_9982,N_9912);
and U10745 (N_10745,N_9897,N_10181);
nand U10746 (N_10746,N_9735,N_10172);
nand U10747 (N_10747,N_9661,N_9628);
nand U10748 (N_10748,N_9645,N_10132);
nor U10749 (N_10749,N_10109,N_9721);
nor U10750 (N_10750,N_9944,N_9780);
nand U10751 (N_10751,N_10012,N_10233);
or U10752 (N_10752,N_9915,N_10272);
nand U10753 (N_10753,N_10165,N_10030);
nor U10754 (N_10754,N_9718,N_9844);
nor U10755 (N_10755,N_9766,N_9696);
or U10756 (N_10756,N_9905,N_10369);
or U10757 (N_10757,N_10096,N_10060);
nor U10758 (N_10758,N_10010,N_10227);
and U10759 (N_10759,N_10397,N_9709);
nand U10760 (N_10760,N_9955,N_10361);
nand U10761 (N_10761,N_9820,N_9858);
or U10762 (N_10762,N_10206,N_10102);
and U10763 (N_10763,N_10220,N_9775);
or U10764 (N_10764,N_10332,N_10321);
nor U10765 (N_10765,N_10128,N_10025);
and U10766 (N_10766,N_9937,N_9887);
or U10767 (N_10767,N_9685,N_10157);
or U10768 (N_10768,N_10029,N_9825);
and U10769 (N_10769,N_9959,N_10013);
nor U10770 (N_10770,N_9972,N_9684);
nor U10771 (N_10771,N_10147,N_9619);
and U10772 (N_10772,N_9977,N_9809);
and U10773 (N_10773,N_10388,N_9788);
nor U10774 (N_10774,N_10278,N_10174);
and U10775 (N_10775,N_9877,N_10154);
nand U10776 (N_10776,N_9787,N_10123);
or U10777 (N_10777,N_10007,N_9873);
and U10778 (N_10778,N_9841,N_10380);
or U10779 (N_10779,N_9926,N_10009);
or U10780 (N_10780,N_10309,N_10044);
and U10781 (N_10781,N_10219,N_10236);
and U10782 (N_10782,N_9914,N_10247);
nor U10783 (N_10783,N_10143,N_10281);
and U10784 (N_10784,N_9616,N_10304);
nand U10785 (N_10785,N_9687,N_10327);
and U10786 (N_10786,N_9965,N_10271);
or U10787 (N_10787,N_9988,N_10310);
or U10788 (N_10788,N_10372,N_10362);
nand U10789 (N_10789,N_9636,N_10003);
nor U10790 (N_10790,N_10256,N_9682);
or U10791 (N_10791,N_9744,N_9801);
or U10792 (N_10792,N_10090,N_9799);
nand U10793 (N_10793,N_9755,N_10180);
nor U10794 (N_10794,N_10252,N_9894);
nand U10795 (N_10795,N_9679,N_9909);
nand U10796 (N_10796,N_9749,N_10189);
nor U10797 (N_10797,N_10035,N_10084);
and U10798 (N_10798,N_9608,N_10038);
nand U10799 (N_10799,N_10117,N_10142);
and U10800 (N_10800,N_9789,N_10251);
nor U10801 (N_10801,N_9891,N_10385);
or U10802 (N_10802,N_9902,N_9833);
or U10803 (N_10803,N_10346,N_10263);
and U10804 (N_10804,N_9917,N_10167);
nor U10805 (N_10805,N_9819,N_9902);
or U10806 (N_10806,N_9976,N_10164);
nor U10807 (N_10807,N_9823,N_10304);
nor U10808 (N_10808,N_9786,N_10337);
nand U10809 (N_10809,N_9767,N_10008);
and U10810 (N_10810,N_10152,N_10118);
or U10811 (N_10811,N_10314,N_10377);
or U10812 (N_10812,N_10276,N_10384);
or U10813 (N_10813,N_10323,N_10034);
and U10814 (N_10814,N_9754,N_10295);
nand U10815 (N_10815,N_10016,N_9936);
or U10816 (N_10816,N_9675,N_9684);
or U10817 (N_10817,N_10144,N_10316);
nor U10818 (N_10818,N_9716,N_9685);
and U10819 (N_10819,N_10250,N_9990);
nor U10820 (N_10820,N_10000,N_9978);
nor U10821 (N_10821,N_10297,N_9837);
or U10822 (N_10822,N_9693,N_9932);
and U10823 (N_10823,N_9738,N_10122);
nor U10824 (N_10824,N_10041,N_10183);
or U10825 (N_10825,N_9609,N_10308);
and U10826 (N_10826,N_10353,N_9684);
nor U10827 (N_10827,N_10259,N_9997);
or U10828 (N_10828,N_9766,N_9801);
and U10829 (N_10829,N_10253,N_10336);
nor U10830 (N_10830,N_10127,N_9755);
nor U10831 (N_10831,N_9958,N_10302);
or U10832 (N_10832,N_10017,N_10084);
nand U10833 (N_10833,N_10264,N_10345);
nand U10834 (N_10834,N_9611,N_9969);
xnor U10835 (N_10835,N_9933,N_9679);
nand U10836 (N_10836,N_9793,N_9617);
nand U10837 (N_10837,N_10307,N_10269);
nand U10838 (N_10838,N_10113,N_9841);
nand U10839 (N_10839,N_9962,N_9984);
nor U10840 (N_10840,N_9855,N_9837);
nand U10841 (N_10841,N_10180,N_10398);
nor U10842 (N_10842,N_10297,N_9859);
or U10843 (N_10843,N_9910,N_9646);
and U10844 (N_10844,N_10301,N_9803);
nand U10845 (N_10845,N_9709,N_10079);
or U10846 (N_10846,N_10121,N_10147);
nand U10847 (N_10847,N_9773,N_10180);
nand U10848 (N_10848,N_10156,N_9891);
nand U10849 (N_10849,N_9663,N_9961);
nor U10850 (N_10850,N_10366,N_9758);
or U10851 (N_10851,N_9893,N_9615);
or U10852 (N_10852,N_9602,N_9653);
nor U10853 (N_10853,N_9984,N_9740);
xnor U10854 (N_10854,N_9747,N_9936);
nor U10855 (N_10855,N_9971,N_9836);
nor U10856 (N_10856,N_9671,N_9926);
or U10857 (N_10857,N_9734,N_10167);
nand U10858 (N_10858,N_10117,N_9882);
and U10859 (N_10859,N_10007,N_9953);
and U10860 (N_10860,N_10332,N_10065);
and U10861 (N_10861,N_10269,N_10354);
nand U10862 (N_10862,N_10261,N_10110);
nand U10863 (N_10863,N_9815,N_10245);
and U10864 (N_10864,N_9910,N_9743);
or U10865 (N_10865,N_9774,N_10120);
nand U10866 (N_10866,N_10096,N_9822);
or U10867 (N_10867,N_9691,N_9733);
nor U10868 (N_10868,N_10163,N_10269);
or U10869 (N_10869,N_10004,N_10229);
nor U10870 (N_10870,N_9799,N_9864);
and U10871 (N_10871,N_10062,N_9694);
or U10872 (N_10872,N_10295,N_9984);
and U10873 (N_10873,N_9650,N_9950);
and U10874 (N_10874,N_10071,N_9875);
nor U10875 (N_10875,N_10012,N_10292);
or U10876 (N_10876,N_9841,N_10219);
nor U10877 (N_10877,N_9702,N_9923);
or U10878 (N_10878,N_9687,N_10066);
nand U10879 (N_10879,N_10112,N_10395);
or U10880 (N_10880,N_9985,N_10016);
or U10881 (N_10881,N_10200,N_9659);
and U10882 (N_10882,N_9880,N_10005);
nand U10883 (N_10883,N_9957,N_10151);
or U10884 (N_10884,N_9638,N_10143);
nand U10885 (N_10885,N_10312,N_10102);
nor U10886 (N_10886,N_10097,N_9874);
and U10887 (N_10887,N_10205,N_10238);
nand U10888 (N_10888,N_9785,N_10393);
or U10889 (N_10889,N_9623,N_10379);
or U10890 (N_10890,N_10286,N_9723);
nor U10891 (N_10891,N_10024,N_10151);
nand U10892 (N_10892,N_9672,N_10197);
and U10893 (N_10893,N_10394,N_9637);
nand U10894 (N_10894,N_9819,N_9687);
nand U10895 (N_10895,N_10161,N_10392);
nor U10896 (N_10896,N_10069,N_9902);
nor U10897 (N_10897,N_10046,N_9880);
and U10898 (N_10898,N_9841,N_9809);
and U10899 (N_10899,N_10212,N_9842);
or U10900 (N_10900,N_9663,N_9666);
nand U10901 (N_10901,N_10206,N_9746);
and U10902 (N_10902,N_9726,N_9971);
and U10903 (N_10903,N_9846,N_10099);
xor U10904 (N_10904,N_9970,N_10124);
or U10905 (N_10905,N_9731,N_9763);
or U10906 (N_10906,N_10227,N_9708);
nand U10907 (N_10907,N_9615,N_9624);
or U10908 (N_10908,N_9721,N_9634);
nor U10909 (N_10909,N_9891,N_9988);
and U10910 (N_10910,N_9896,N_10083);
and U10911 (N_10911,N_10388,N_10096);
and U10912 (N_10912,N_9908,N_10244);
and U10913 (N_10913,N_9648,N_10355);
nor U10914 (N_10914,N_10072,N_10229);
or U10915 (N_10915,N_9885,N_9917);
nor U10916 (N_10916,N_10177,N_9928);
and U10917 (N_10917,N_10269,N_10135);
and U10918 (N_10918,N_10131,N_9646);
or U10919 (N_10919,N_9994,N_10291);
nand U10920 (N_10920,N_10159,N_10346);
nor U10921 (N_10921,N_10379,N_10166);
and U10922 (N_10922,N_9839,N_10030);
nand U10923 (N_10923,N_10302,N_10313);
or U10924 (N_10924,N_9637,N_10097);
or U10925 (N_10925,N_9807,N_10171);
and U10926 (N_10926,N_10148,N_9822);
nor U10927 (N_10927,N_10397,N_9775);
and U10928 (N_10928,N_9829,N_9640);
nor U10929 (N_10929,N_9736,N_10030);
nand U10930 (N_10930,N_9828,N_10155);
or U10931 (N_10931,N_9692,N_10179);
nand U10932 (N_10932,N_9642,N_9917);
nor U10933 (N_10933,N_9663,N_9632);
and U10934 (N_10934,N_9876,N_9929);
nand U10935 (N_10935,N_10291,N_9706);
nor U10936 (N_10936,N_9822,N_10348);
or U10937 (N_10937,N_9824,N_10399);
nor U10938 (N_10938,N_9898,N_10018);
nand U10939 (N_10939,N_10074,N_10242);
nand U10940 (N_10940,N_9722,N_9935);
and U10941 (N_10941,N_9751,N_10239);
nand U10942 (N_10942,N_10096,N_9617);
or U10943 (N_10943,N_9603,N_10270);
nand U10944 (N_10944,N_9966,N_10215);
nand U10945 (N_10945,N_10055,N_10096);
or U10946 (N_10946,N_10287,N_10137);
nand U10947 (N_10947,N_10029,N_10031);
nor U10948 (N_10948,N_10140,N_10176);
nand U10949 (N_10949,N_10353,N_10136);
nand U10950 (N_10950,N_10068,N_9787);
and U10951 (N_10951,N_10045,N_9643);
or U10952 (N_10952,N_10150,N_10091);
xnor U10953 (N_10953,N_10024,N_9969);
nor U10954 (N_10954,N_10285,N_9643);
nand U10955 (N_10955,N_9752,N_10319);
nor U10956 (N_10956,N_10173,N_9646);
and U10957 (N_10957,N_9994,N_9849);
nor U10958 (N_10958,N_9807,N_9681);
nor U10959 (N_10959,N_9737,N_10171);
and U10960 (N_10960,N_10077,N_9876);
and U10961 (N_10961,N_9789,N_10217);
nand U10962 (N_10962,N_9895,N_10210);
nand U10963 (N_10963,N_10112,N_10299);
nand U10964 (N_10964,N_10063,N_10039);
or U10965 (N_10965,N_9824,N_9991);
nand U10966 (N_10966,N_9725,N_10171);
or U10967 (N_10967,N_10009,N_10119);
nor U10968 (N_10968,N_10270,N_10064);
nand U10969 (N_10969,N_9919,N_9750);
and U10970 (N_10970,N_9728,N_10265);
or U10971 (N_10971,N_10279,N_10363);
nand U10972 (N_10972,N_10144,N_10295);
nand U10973 (N_10973,N_10261,N_9765);
and U10974 (N_10974,N_10242,N_10231);
nand U10975 (N_10975,N_9624,N_9707);
and U10976 (N_10976,N_9917,N_9871);
nor U10977 (N_10977,N_9763,N_10178);
nand U10978 (N_10978,N_10169,N_10392);
or U10979 (N_10979,N_10298,N_9691);
and U10980 (N_10980,N_10120,N_10263);
nor U10981 (N_10981,N_9935,N_9645);
nor U10982 (N_10982,N_10394,N_10142);
nor U10983 (N_10983,N_10109,N_9724);
nand U10984 (N_10984,N_9999,N_9607);
nor U10985 (N_10985,N_10382,N_9858);
nor U10986 (N_10986,N_10269,N_9915);
nand U10987 (N_10987,N_10202,N_10333);
and U10988 (N_10988,N_9880,N_10059);
and U10989 (N_10989,N_10162,N_10348);
nor U10990 (N_10990,N_9926,N_10081);
and U10991 (N_10991,N_10381,N_9777);
nor U10992 (N_10992,N_10134,N_10384);
nand U10993 (N_10993,N_10275,N_10251);
or U10994 (N_10994,N_9914,N_9996);
nor U10995 (N_10995,N_9761,N_10391);
or U10996 (N_10996,N_10205,N_9700);
nand U10997 (N_10997,N_9790,N_10121);
and U10998 (N_10998,N_10280,N_9961);
nand U10999 (N_10999,N_9825,N_9637);
or U11000 (N_11000,N_9756,N_9779);
and U11001 (N_11001,N_10315,N_9753);
nor U11002 (N_11002,N_10004,N_10224);
nand U11003 (N_11003,N_10298,N_9928);
nand U11004 (N_11004,N_10261,N_9779);
or U11005 (N_11005,N_10005,N_10026);
nand U11006 (N_11006,N_9672,N_10080);
nor U11007 (N_11007,N_10053,N_10054);
and U11008 (N_11008,N_9899,N_9691);
nand U11009 (N_11009,N_10220,N_10091);
nand U11010 (N_11010,N_10025,N_9675);
or U11011 (N_11011,N_10327,N_10264);
or U11012 (N_11012,N_10104,N_9660);
nor U11013 (N_11013,N_10272,N_10035);
nor U11014 (N_11014,N_9838,N_9675);
or U11015 (N_11015,N_9614,N_9945);
nand U11016 (N_11016,N_9961,N_9694);
and U11017 (N_11017,N_10104,N_10207);
and U11018 (N_11018,N_9696,N_10261);
nor U11019 (N_11019,N_9653,N_10059);
or U11020 (N_11020,N_10309,N_10084);
nor U11021 (N_11021,N_9684,N_10093);
or U11022 (N_11022,N_10005,N_9744);
and U11023 (N_11023,N_10388,N_9783);
and U11024 (N_11024,N_9933,N_9960);
nor U11025 (N_11025,N_10200,N_9650);
and U11026 (N_11026,N_10093,N_10388);
nor U11027 (N_11027,N_9875,N_9648);
or U11028 (N_11028,N_9744,N_9813);
and U11029 (N_11029,N_10282,N_10222);
or U11030 (N_11030,N_9673,N_9912);
and U11031 (N_11031,N_10318,N_9973);
and U11032 (N_11032,N_10216,N_9687);
or U11033 (N_11033,N_9856,N_9932);
nor U11034 (N_11034,N_9921,N_10109);
nand U11035 (N_11035,N_10089,N_9960);
nor U11036 (N_11036,N_9854,N_9891);
xor U11037 (N_11037,N_10352,N_10200);
nand U11038 (N_11038,N_9834,N_10085);
nor U11039 (N_11039,N_9871,N_9956);
and U11040 (N_11040,N_9767,N_9943);
or U11041 (N_11041,N_10119,N_10012);
and U11042 (N_11042,N_10283,N_9953);
nand U11043 (N_11043,N_10075,N_10158);
nor U11044 (N_11044,N_10241,N_10082);
or U11045 (N_11045,N_10028,N_9881);
and U11046 (N_11046,N_10171,N_10338);
nor U11047 (N_11047,N_10292,N_9776);
nor U11048 (N_11048,N_10066,N_10089);
xnor U11049 (N_11049,N_10003,N_9856);
nor U11050 (N_11050,N_10335,N_9785);
nand U11051 (N_11051,N_10058,N_10289);
or U11052 (N_11052,N_10135,N_9899);
or U11053 (N_11053,N_9822,N_9853);
or U11054 (N_11054,N_9741,N_10323);
nand U11055 (N_11055,N_10291,N_9708);
nor U11056 (N_11056,N_9790,N_9750);
nand U11057 (N_11057,N_9689,N_9982);
nor U11058 (N_11058,N_9886,N_10326);
nor U11059 (N_11059,N_10085,N_10239);
nand U11060 (N_11060,N_10112,N_10394);
nor U11061 (N_11061,N_9785,N_9848);
and U11062 (N_11062,N_10072,N_10080);
and U11063 (N_11063,N_9647,N_9740);
and U11064 (N_11064,N_10334,N_9685);
nand U11065 (N_11065,N_10298,N_9732);
and U11066 (N_11066,N_9799,N_9757);
nor U11067 (N_11067,N_10013,N_10212);
nor U11068 (N_11068,N_9622,N_9944);
or U11069 (N_11069,N_9847,N_10100);
or U11070 (N_11070,N_10393,N_9911);
nor U11071 (N_11071,N_9917,N_9790);
nand U11072 (N_11072,N_10235,N_10133);
nor U11073 (N_11073,N_9780,N_10286);
nand U11074 (N_11074,N_9766,N_10015);
and U11075 (N_11075,N_10253,N_10006);
nor U11076 (N_11076,N_9855,N_10163);
or U11077 (N_11077,N_10385,N_9982);
nand U11078 (N_11078,N_10038,N_9818);
and U11079 (N_11079,N_10118,N_10108);
nand U11080 (N_11080,N_9980,N_9775);
nand U11081 (N_11081,N_9944,N_9773);
and U11082 (N_11082,N_10368,N_10096);
nand U11083 (N_11083,N_9794,N_10175);
nor U11084 (N_11084,N_9924,N_9603);
or U11085 (N_11085,N_10241,N_9721);
or U11086 (N_11086,N_9746,N_10229);
and U11087 (N_11087,N_9660,N_10036);
or U11088 (N_11088,N_10305,N_10189);
nor U11089 (N_11089,N_9603,N_9753);
nand U11090 (N_11090,N_10129,N_9742);
nor U11091 (N_11091,N_10005,N_10351);
or U11092 (N_11092,N_9798,N_9679);
nor U11093 (N_11093,N_10057,N_9993);
nand U11094 (N_11094,N_9830,N_9695);
or U11095 (N_11095,N_9635,N_9743);
nand U11096 (N_11096,N_10174,N_10324);
nor U11097 (N_11097,N_9654,N_9705);
nor U11098 (N_11098,N_9863,N_10161);
and U11099 (N_11099,N_10228,N_9609);
and U11100 (N_11100,N_9928,N_10074);
nor U11101 (N_11101,N_10196,N_9608);
and U11102 (N_11102,N_10008,N_9929);
nand U11103 (N_11103,N_10285,N_10085);
nand U11104 (N_11104,N_9817,N_10371);
or U11105 (N_11105,N_10393,N_9732);
nor U11106 (N_11106,N_9817,N_10123);
nand U11107 (N_11107,N_9895,N_9697);
and U11108 (N_11108,N_10095,N_10246);
and U11109 (N_11109,N_9878,N_10164);
nand U11110 (N_11110,N_10140,N_10390);
nand U11111 (N_11111,N_9785,N_9663);
and U11112 (N_11112,N_9737,N_10228);
or U11113 (N_11113,N_9835,N_10253);
nor U11114 (N_11114,N_9810,N_10326);
or U11115 (N_11115,N_9682,N_10011);
nor U11116 (N_11116,N_9913,N_10398);
nand U11117 (N_11117,N_10152,N_9977);
nor U11118 (N_11118,N_10307,N_9720);
or U11119 (N_11119,N_9891,N_9814);
or U11120 (N_11120,N_9709,N_10278);
nand U11121 (N_11121,N_9699,N_9987);
or U11122 (N_11122,N_10094,N_9798);
xor U11123 (N_11123,N_10241,N_9922);
nor U11124 (N_11124,N_9958,N_9637);
or U11125 (N_11125,N_9761,N_9787);
or U11126 (N_11126,N_9771,N_9777);
nor U11127 (N_11127,N_9671,N_10123);
nor U11128 (N_11128,N_9993,N_9888);
nor U11129 (N_11129,N_10301,N_10244);
or U11130 (N_11130,N_9696,N_10357);
and U11131 (N_11131,N_9873,N_10303);
nand U11132 (N_11132,N_9825,N_9737);
and U11133 (N_11133,N_9819,N_10010);
nand U11134 (N_11134,N_9765,N_10377);
nand U11135 (N_11135,N_9735,N_10021);
nand U11136 (N_11136,N_9878,N_10351);
or U11137 (N_11137,N_9832,N_10186);
nand U11138 (N_11138,N_10243,N_9895);
and U11139 (N_11139,N_9736,N_10287);
and U11140 (N_11140,N_10336,N_10045);
and U11141 (N_11141,N_9746,N_10022);
and U11142 (N_11142,N_9929,N_10205);
or U11143 (N_11143,N_9747,N_9746);
or U11144 (N_11144,N_10219,N_10112);
and U11145 (N_11145,N_9767,N_9869);
or U11146 (N_11146,N_10208,N_9618);
nor U11147 (N_11147,N_10241,N_10126);
nor U11148 (N_11148,N_10201,N_10244);
and U11149 (N_11149,N_10007,N_9615);
nand U11150 (N_11150,N_10337,N_10247);
nor U11151 (N_11151,N_10241,N_9763);
nor U11152 (N_11152,N_10172,N_9825);
nand U11153 (N_11153,N_10269,N_9677);
and U11154 (N_11154,N_9896,N_10133);
nand U11155 (N_11155,N_9615,N_10228);
or U11156 (N_11156,N_10107,N_10372);
nor U11157 (N_11157,N_9864,N_9645);
nor U11158 (N_11158,N_10023,N_9823);
and U11159 (N_11159,N_10073,N_9864);
nor U11160 (N_11160,N_9853,N_10214);
nor U11161 (N_11161,N_10071,N_10059);
or U11162 (N_11162,N_9978,N_9845);
or U11163 (N_11163,N_9971,N_10010);
and U11164 (N_11164,N_10013,N_9813);
nand U11165 (N_11165,N_9693,N_10084);
or U11166 (N_11166,N_10076,N_9695);
or U11167 (N_11167,N_10268,N_9995);
nand U11168 (N_11168,N_10149,N_10002);
or U11169 (N_11169,N_10236,N_10118);
nand U11170 (N_11170,N_10099,N_9724);
and U11171 (N_11171,N_9606,N_9936);
xnor U11172 (N_11172,N_10322,N_9808);
nand U11173 (N_11173,N_9836,N_10016);
or U11174 (N_11174,N_9896,N_9907);
or U11175 (N_11175,N_9929,N_10028);
and U11176 (N_11176,N_10024,N_10183);
nor U11177 (N_11177,N_10357,N_9682);
and U11178 (N_11178,N_9907,N_9942);
and U11179 (N_11179,N_9622,N_10049);
nor U11180 (N_11180,N_10291,N_10133);
nand U11181 (N_11181,N_9799,N_10318);
or U11182 (N_11182,N_9849,N_9679);
nor U11183 (N_11183,N_9686,N_9977);
or U11184 (N_11184,N_9726,N_10146);
or U11185 (N_11185,N_10113,N_9661);
nor U11186 (N_11186,N_9963,N_10050);
or U11187 (N_11187,N_10217,N_9893);
nor U11188 (N_11188,N_9825,N_10338);
and U11189 (N_11189,N_9937,N_9640);
or U11190 (N_11190,N_9649,N_10331);
nor U11191 (N_11191,N_9768,N_10206);
nor U11192 (N_11192,N_10391,N_9662);
nor U11193 (N_11193,N_9780,N_10053);
nand U11194 (N_11194,N_9744,N_9714);
and U11195 (N_11195,N_10343,N_9663);
nor U11196 (N_11196,N_9701,N_10135);
or U11197 (N_11197,N_9864,N_10359);
or U11198 (N_11198,N_9990,N_10273);
or U11199 (N_11199,N_10383,N_10122);
nor U11200 (N_11200,N_10559,N_10568);
nor U11201 (N_11201,N_10666,N_10806);
nor U11202 (N_11202,N_11173,N_10723);
or U11203 (N_11203,N_11007,N_11114);
nand U11204 (N_11204,N_10580,N_10824);
and U11205 (N_11205,N_10887,N_10965);
nand U11206 (N_11206,N_10602,N_10859);
or U11207 (N_11207,N_10505,N_10698);
nand U11208 (N_11208,N_10810,N_11148);
or U11209 (N_11209,N_11073,N_11181);
nand U11210 (N_11210,N_10593,N_10402);
and U11211 (N_11211,N_10491,N_10823);
and U11212 (N_11212,N_10769,N_10653);
nor U11213 (N_11213,N_11140,N_10622);
nor U11214 (N_11214,N_11196,N_10743);
and U11215 (N_11215,N_10672,N_10554);
nor U11216 (N_11216,N_10456,N_11195);
nand U11217 (N_11217,N_10676,N_11055);
and U11218 (N_11218,N_10684,N_10889);
and U11219 (N_11219,N_10663,N_10601);
or U11220 (N_11220,N_10725,N_10413);
nand U11221 (N_11221,N_10520,N_10801);
nand U11222 (N_11222,N_10641,N_10635);
nor U11223 (N_11223,N_10944,N_10691);
nand U11224 (N_11224,N_11092,N_11040);
or U11225 (N_11225,N_11070,N_10951);
nor U11226 (N_11226,N_10667,N_10862);
nand U11227 (N_11227,N_10938,N_10523);
and U11228 (N_11228,N_11194,N_11011);
nand U11229 (N_11229,N_11042,N_10976);
and U11230 (N_11230,N_10940,N_10713);
nand U11231 (N_11231,N_10752,N_10606);
and U11232 (N_11232,N_10816,N_10910);
nand U11233 (N_11233,N_10758,N_11032);
and U11234 (N_11234,N_10902,N_10675);
and U11235 (N_11235,N_11090,N_11163);
nand U11236 (N_11236,N_10891,N_10754);
nand U11237 (N_11237,N_11013,N_10953);
nor U11238 (N_11238,N_10613,N_10884);
nor U11239 (N_11239,N_10971,N_11096);
nand U11240 (N_11240,N_10818,N_10681);
nor U11241 (N_11241,N_10646,N_10843);
and U11242 (N_11242,N_10524,N_10893);
nand U11243 (N_11243,N_11156,N_10868);
nand U11244 (N_11244,N_10642,N_10920);
and U11245 (N_11245,N_10917,N_10746);
nand U11246 (N_11246,N_10848,N_10756);
nor U11247 (N_11247,N_11034,N_11121);
nor U11248 (N_11248,N_10650,N_11087);
nor U11249 (N_11249,N_10931,N_11144);
and U11250 (N_11250,N_10620,N_10738);
or U11251 (N_11251,N_11113,N_10498);
and U11252 (N_11252,N_11190,N_10897);
nor U11253 (N_11253,N_10423,N_11037);
xor U11254 (N_11254,N_10531,N_10945);
nand U11255 (N_11255,N_10793,N_10452);
and U11256 (N_11256,N_11115,N_10429);
or U11257 (N_11257,N_10730,N_10831);
or U11258 (N_11258,N_10465,N_11175);
and U11259 (N_11259,N_10728,N_10934);
or U11260 (N_11260,N_10797,N_11160);
and U11261 (N_11261,N_10710,N_10670);
or U11262 (N_11262,N_10608,N_10538);
or U11263 (N_11263,N_11157,N_11149);
nor U11264 (N_11264,N_10655,N_10913);
nor U11265 (N_11265,N_10790,N_10566);
and U11266 (N_11266,N_10814,N_10533);
nand U11267 (N_11267,N_10584,N_10490);
nand U11268 (N_11268,N_10478,N_11048);
and U11269 (N_11269,N_10495,N_10749);
and U11270 (N_11270,N_10428,N_10509);
nor U11271 (N_11271,N_10853,N_11005);
nor U11272 (N_11272,N_10909,N_10841);
nand U11273 (N_11273,N_11107,N_10536);
and U11274 (N_11274,N_10729,N_10718);
nand U11275 (N_11275,N_11057,N_10407);
nor U11276 (N_11276,N_10677,N_10694);
nor U11277 (N_11277,N_11162,N_10585);
or U11278 (N_11278,N_10786,N_10547);
and U11279 (N_11279,N_10532,N_10764);
nand U11280 (N_11280,N_11008,N_11147);
nor U11281 (N_11281,N_10832,N_10974);
or U11282 (N_11282,N_10419,N_10783);
and U11283 (N_11283,N_10851,N_10789);
or U11284 (N_11284,N_11120,N_10665);
and U11285 (N_11285,N_11052,N_11061);
nor U11286 (N_11286,N_11025,N_10846);
nand U11287 (N_11287,N_10686,N_10594);
or U11288 (N_11288,N_11091,N_10855);
nand U11289 (N_11289,N_11085,N_10412);
nor U11290 (N_11290,N_11118,N_10401);
or U11291 (N_11291,N_10486,N_10682);
nor U11292 (N_11292,N_10502,N_10581);
or U11293 (N_11293,N_10572,N_10624);
and U11294 (N_11294,N_10527,N_10599);
nor U11295 (N_11295,N_10869,N_11150);
nor U11296 (N_11296,N_10946,N_10956);
nor U11297 (N_11297,N_10575,N_10437);
or U11298 (N_11298,N_10448,N_11129);
and U11299 (N_11299,N_11179,N_10629);
nor U11300 (N_11300,N_10453,N_10949);
and U11301 (N_11301,N_11093,N_10717);
nand U11302 (N_11302,N_11003,N_11063);
nand U11303 (N_11303,N_10709,N_10493);
or U11304 (N_11304,N_10741,N_10430);
and U11305 (N_11305,N_10800,N_10455);
or U11306 (N_11306,N_10778,N_10739);
and U11307 (N_11307,N_10432,N_10995);
nand U11308 (N_11308,N_10903,N_10883);
and U11309 (N_11309,N_10745,N_11192);
or U11310 (N_11310,N_11026,N_10640);
or U11311 (N_11311,N_10591,N_11119);
xnor U11312 (N_11312,N_10583,N_10632);
nand U11313 (N_11313,N_11044,N_10551);
or U11314 (N_11314,N_10444,N_10664);
or U11315 (N_11315,N_11176,N_11064);
nor U11316 (N_11316,N_10701,N_10898);
and U11317 (N_11317,N_10659,N_11078);
nor U11318 (N_11318,N_11006,N_11095);
nand U11319 (N_11319,N_11153,N_11111);
or U11320 (N_11320,N_10481,N_10757);
and U11321 (N_11321,N_10431,N_10529);
nor U11322 (N_11322,N_11009,N_10708);
and U11323 (N_11323,N_10464,N_11030);
nand U11324 (N_11324,N_10886,N_10919);
nand U11325 (N_11325,N_11143,N_10535);
and U11326 (N_11326,N_10497,N_11101);
or U11327 (N_11327,N_10712,N_11123);
and U11328 (N_11328,N_10427,N_11075);
or U11329 (N_11329,N_11130,N_10929);
or U11330 (N_11330,N_10522,N_10807);
and U11331 (N_11331,N_11184,N_10703);
nand U11332 (N_11332,N_10454,N_10611);
or U11333 (N_11333,N_11116,N_10834);
and U11334 (N_11334,N_10612,N_10623);
and U11335 (N_11335,N_10751,N_10982);
or U11336 (N_11336,N_10403,N_10857);
nand U11337 (N_11337,N_11098,N_11188);
xnor U11338 (N_11338,N_11014,N_10827);
nor U11339 (N_11339,N_11000,N_10406);
nand U11340 (N_11340,N_10589,N_10962);
and U11341 (N_11341,N_10469,N_11083);
nand U11342 (N_11342,N_10459,N_10442);
and U11343 (N_11343,N_11178,N_10922);
nand U11344 (N_11344,N_10879,N_11109);
nand U11345 (N_11345,N_10711,N_10901);
or U11346 (N_11346,N_10519,N_10685);
nand U11347 (N_11347,N_10918,N_10961);
and U11348 (N_11348,N_10617,N_10908);
or U11349 (N_11349,N_10933,N_10417);
nand U11350 (N_11350,N_10802,N_11043);
nor U11351 (N_11351,N_10947,N_11062);
or U11352 (N_11352,N_10721,N_10492);
xor U11353 (N_11353,N_10979,N_11038);
nor U11354 (N_11354,N_10876,N_10537);
nand U11355 (N_11355,N_10496,N_10578);
and U11356 (N_11356,N_10528,N_10614);
or U11357 (N_11357,N_10610,N_10470);
and U11358 (N_11358,N_10792,N_11161);
and U11359 (N_11359,N_11127,N_10542);
nand U11360 (N_11360,N_11158,N_10959);
and U11361 (N_11361,N_10992,N_10768);
and U11362 (N_11362,N_11145,N_11185);
nor U11363 (N_11363,N_10815,N_10760);
nand U11364 (N_11364,N_11125,N_10759);
or U11365 (N_11365,N_10636,N_10451);
or U11366 (N_11366,N_11047,N_10467);
nand U11367 (N_11367,N_10942,N_10480);
nand U11368 (N_11368,N_11106,N_10443);
nor U11369 (N_11369,N_10939,N_10514);
and U11370 (N_11370,N_10744,N_10915);
nand U11371 (N_11371,N_10557,N_11135);
nand U11372 (N_11372,N_10870,N_10424);
or U11373 (N_11373,N_10895,N_10967);
nand U11374 (N_11374,N_10411,N_11050);
nand U11375 (N_11375,N_10704,N_10461);
or U11376 (N_11376,N_10726,N_10488);
or U11377 (N_11377,N_10626,N_11060);
nand U11378 (N_11378,N_10863,N_10660);
nand U11379 (N_11379,N_11152,N_11079);
nand U11380 (N_11380,N_11132,N_11141);
nand U11381 (N_11381,N_10852,N_10410);
nand U11382 (N_11382,N_10516,N_10991);
or U11383 (N_11383,N_10925,N_10963);
and U11384 (N_11384,N_10926,N_10560);
nor U11385 (N_11385,N_11051,N_10668);
and U11386 (N_11386,N_10647,N_10872);
nor U11387 (N_11387,N_10860,N_10742);
nand U11388 (N_11388,N_10702,N_10564);
or U11389 (N_11389,N_10927,N_11080);
and U11390 (N_11390,N_11069,N_11108);
or U11391 (N_11391,N_10540,N_10878);
or U11392 (N_11392,N_10795,N_10700);
and U11393 (N_11393,N_10981,N_10999);
nand U11394 (N_11394,N_10472,N_11198);
and U11395 (N_11395,N_10501,N_10762);
nand U11396 (N_11396,N_10874,N_10798);
nor U11397 (N_11397,N_10994,N_10658);
or U11398 (N_11398,N_11021,N_10761);
nor U11399 (N_11399,N_10534,N_10662);
or U11400 (N_11400,N_11053,N_10777);
nor U11401 (N_11401,N_10780,N_10936);
nand U11402 (N_11402,N_10871,N_11104);
nand U11403 (N_11403,N_10914,N_10479);
nor U11404 (N_11404,N_11159,N_10861);
or U11405 (N_11405,N_10881,N_11049);
nand U11406 (N_11406,N_10805,N_10696);
and U11407 (N_11407,N_10548,N_11019);
and U11408 (N_11408,N_11010,N_10794);
and U11409 (N_11409,N_10955,N_10784);
and U11410 (N_11410,N_10485,N_11137);
or U11411 (N_11411,N_10899,N_10421);
or U11412 (N_11412,N_10799,N_11122);
nand U11413 (N_11413,N_11187,N_10673);
nand U11414 (N_11414,N_10625,N_10733);
nand U11415 (N_11415,N_10724,N_10838);
and U11416 (N_11416,N_10577,N_10693);
and U11417 (N_11417,N_11031,N_10638);
nor U11418 (N_11418,N_11142,N_10924);
nand U11419 (N_11419,N_10621,N_11099);
nor U11420 (N_11420,N_10517,N_10867);
or U11421 (N_11421,N_11133,N_11165);
nor U11422 (N_11422,N_10634,N_10458);
nand U11423 (N_11423,N_10513,N_10661);
and U11424 (N_11424,N_10678,N_10449);
or U11425 (N_11425,N_11084,N_10989);
nor U11426 (N_11426,N_10828,N_11169);
or U11427 (N_11427,N_10541,N_10969);
nand U11428 (N_11428,N_10445,N_11033);
nor U11429 (N_11429,N_10582,N_11066);
or U11430 (N_11430,N_10980,N_11059);
nor U11431 (N_11431,N_10836,N_10890);
nor U11432 (N_11432,N_10494,N_10657);
nand U11433 (N_11433,N_10719,N_10482);
or U11434 (N_11434,N_10787,N_10607);
nand U11435 (N_11435,N_10996,N_11199);
nand U11436 (N_11436,N_10574,N_10483);
nand U11437 (N_11437,N_10715,N_10839);
nor U11438 (N_11438,N_10561,N_11002);
or U11439 (N_11439,N_10986,N_10811);
or U11440 (N_11440,N_11186,N_11071);
and U11441 (N_11441,N_11136,N_11017);
nand U11442 (N_11442,N_10615,N_11012);
nand U11443 (N_11443,N_10714,N_10952);
or U11444 (N_11444,N_10735,N_10829);
nand U11445 (N_11445,N_10819,N_10425);
nor U11446 (N_11446,N_11054,N_10690);
or U11447 (N_11447,N_10770,N_11029);
or U11448 (N_11448,N_10512,N_11004);
or U11449 (N_11449,N_10679,N_10987);
and U11450 (N_11450,N_10434,N_10556);
nor U11451 (N_11451,N_10555,N_10567);
or U11452 (N_11452,N_10825,N_10750);
or U11453 (N_11453,N_10408,N_10603);
nor U11454 (N_11454,N_10618,N_10779);
or U11455 (N_11455,N_10985,N_11089);
nand U11456 (N_11456,N_10404,N_11097);
or U11457 (N_11457,N_10854,N_10518);
nor U11458 (N_11458,N_10821,N_10426);
nor U11459 (N_11459,N_10616,N_10562);
or U11460 (N_11460,N_11068,N_11046);
and U11461 (N_11461,N_10695,N_10935);
nand U11462 (N_11462,N_10900,N_10774);
or U11463 (N_11463,N_10888,N_10643);
nand U11464 (N_11464,N_11027,N_10771);
and U11465 (N_11465,N_11022,N_10896);
nor U11466 (N_11466,N_10446,N_10569);
or U11467 (N_11467,N_10484,N_10511);
nand U11468 (N_11468,N_10648,N_10782);
and U11469 (N_11469,N_11105,N_10877);
or U11470 (N_11470,N_11082,N_10579);
and U11471 (N_11471,N_10705,N_10968);
and U11472 (N_11472,N_10791,N_11100);
nor U11473 (N_11473,N_10983,N_10950);
or U11474 (N_11474,N_10573,N_10652);
and U11475 (N_11475,N_11088,N_10553);
or U11476 (N_11476,N_11128,N_10639);
or U11477 (N_11477,N_10627,N_10439);
nor U11478 (N_11478,N_10748,N_11045);
nand U11479 (N_11479,N_10804,N_10858);
and U11480 (N_11480,N_10587,N_10978);
nor U11481 (N_11481,N_11086,N_10865);
and U11482 (N_11482,N_10476,N_11072);
nand U11483 (N_11483,N_10438,N_10803);
and U11484 (N_11484,N_10781,N_10977);
and U11485 (N_11485,N_10414,N_10904);
nor U11486 (N_11486,N_10409,N_10563);
or U11487 (N_11487,N_10785,N_11191);
and U11488 (N_11488,N_10833,N_11039);
and U11489 (N_11489,N_10500,N_10948);
and U11490 (N_11490,N_10630,N_11058);
or U11491 (N_11491,N_10507,N_11065);
and U11492 (N_11492,N_10549,N_11134);
nor U11493 (N_11493,N_10775,N_10973);
nand U11494 (N_11494,N_11126,N_10740);
nand U11495 (N_11495,N_10477,N_10656);
or U11496 (N_11496,N_10958,N_11001);
nor U11497 (N_11497,N_10755,N_11124);
or U11498 (N_11498,N_10960,N_10707);
nand U11499 (N_11499,N_10609,N_10916);
and U11500 (N_11500,N_11035,N_11177);
nor U11501 (N_11501,N_11197,N_10975);
nor U11502 (N_11502,N_10813,N_10683);
or U11503 (N_11503,N_10911,N_10737);
or U11504 (N_11504,N_10543,N_10812);
nand U11505 (N_11505,N_11074,N_10418);
nand U11506 (N_11506,N_10586,N_10689);
nand U11507 (N_11507,N_10474,N_11016);
nor U11508 (N_11508,N_11024,N_10436);
or U11509 (N_11509,N_10966,N_10595);
nor U11510 (N_11510,N_11112,N_10687);
or U11511 (N_11511,N_10720,N_10400);
nor U11512 (N_11512,N_11171,N_10840);
nand U11513 (N_11513,N_10849,N_11102);
nand U11514 (N_11514,N_10637,N_11170);
nor U11515 (N_11515,N_10984,N_10435);
nand U11516 (N_11516,N_10850,N_10928);
nor U11517 (N_11517,N_10466,N_10471);
or U11518 (N_11518,N_10415,N_10510);
nor U11519 (N_11519,N_10592,N_10450);
and U11520 (N_11520,N_11183,N_10463);
nand U11521 (N_11521,N_10504,N_10565);
nor U11522 (N_11522,N_11146,N_10732);
nor U11523 (N_11523,N_10796,N_10882);
and U11524 (N_11524,N_10697,N_10550);
nand U11525 (N_11525,N_10930,N_10998);
nor U11526 (N_11526,N_10788,N_11155);
nand U11527 (N_11527,N_10526,N_10837);
nand U11528 (N_11528,N_10521,N_10880);
or U11529 (N_11529,N_10590,N_10628);
nor U11530 (N_11530,N_10416,N_10923);
nand U11531 (N_11531,N_10604,N_10885);
or U11532 (N_11532,N_10826,N_10441);
nor U11533 (N_11533,N_10722,N_10649);
nor U11534 (N_11534,N_10468,N_10907);
nor U11535 (N_11535,N_10835,N_10866);
and U11536 (N_11536,N_10506,N_10530);
nand U11537 (N_11537,N_10912,N_10763);
nor U11538 (N_11538,N_11131,N_11028);
and U11539 (N_11539,N_10440,N_10447);
xnor U11540 (N_11540,N_11103,N_10892);
and U11541 (N_11541,N_10921,N_10460);
nor U11542 (N_11542,N_10864,N_10773);
nor U11543 (N_11543,N_10766,N_11020);
nand U11544 (N_11544,N_10767,N_11180);
nor U11545 (N_11545,N_10906,N_10957);
or U11546 (N_11546,N_11036,N_11151);
nor U11547 (N_11547,N_11138,N_10808);
nor U11548 (N_11548,N_11015,N_10651);
and U11549 (N_11549,N_10731,N_11168);
or U11550 (N_11550,N_10597,N_10422);
and U11551 (N_11551,N_10558,N_10736);
nand U11552 (N_11552,N_10988,N_10576);
nor U11553 (N_11553,N_10894,N_10932);
nand U11554 (N_11554,N_10644,N_11189);
nand U11555 (N_11555,N_10845,N_11094);
nand U11556 (N_11556,N_11154,N_11166);
nor U11557 (N_11557,N_10964,N_10954);
and U11558 (N_11558,N_10747,N_10475);
nor U11559 (N_11559,N_10539,N_11182);
or U11560 (N_11560,N_10457,N_10544);
and U11561 (N_11561,N_10820,N_10552);
nand U11562 (N_11562,N_11076,N_10598);
nor U11563 (N_11563,N_10645,N_10844);
or U11564 (N_11564,N_10420,N_10588);
nand U11565 (N_11565,N_10633,N_10716);
nor U11566 (N_11566,N_10856,N_10706);
nor U11567 (N_11567,N_10674,N_10462);
nand U11568 (N_11568,N_10993,N_10692);
nor U11569 (N_11569,N_10515,N_10619);
nor U11570 (N_11570,N_11193,N_10941);
nand U11571 (N_11571,N_11056,N_10822);
nor U11572 (N_11572,N_10943,N_10847);
nand U11573 (N_11573,N_10997,N_10817);
or U11574 (N_11574,N_10499,N_10830);
nand U11575 (N_11575,N_10508,N_10842);
nand U11576 (N_11576,N_10525,N_11174);
or U11577 (N_11577,N_10753,N_10503);
nor U11578 (N_11578,N_10809,N_10734);
nor U11579 (N_11579,N_11023,N_10688);
nor U11580 (N_11580,N_10680,N_11139);
and U11581 (N_11581,N_10727,N_10905);
nand U11582 (N_11582,N_10545,N_10654);
and U11583 (N_11583,N_11110,N_10776);
nor U11584 (N_11584,N_11081,N_11167);
nor U11585 (N_11585,N_10487,N_10405);
nand U11586 (N_11586,N_10669,N_11077);
nor U11587 (N_11587,N_10473,N_10489);
nand U11588 (N_11588,N_10605,N_10546);
or U11589 (N_11589,N_10970,N_11067);
nor U11590 (N_11590,N_11018,N_11164);
or U11591 (N_11591,N_11172,N_10433);
nor U11592 (N_11592,N_10596,N_10873);
nor U11593 (N_11593,N_10570,N_10990);
or U11594 (N_11594,N_10772,N_11041);
nand U11595 (N_11595,N_10937,N_11117);
nand U11596 (N_11596,N_10765,N_10875);
nand U11597 (N_11597,N_10600,N_10671);
nor U11598 (N_11598,N_10571,N_10699);
or U11599 (N_11599,N_10972,N_10631);
nor U11600 (N_11600,N_11177,N_10997);
nor U11601 (N_11601,N_11072,N_10660);
and U11602 (N_11602,N_10839,N_10549);
or U11603 (N_11603,N_10964,N_11180);
nand U11604 (N_11604,N_10587,N_10628);
or U11605 (N_11605,N_11016,N_10412);
nand U11606 (N_11606,N_11118,N_10826);
nor U11607 (N_11607,N_10750,N_10603);
and U11608 (N_11608,N_10669,N_10620);
nor U11609 (N_11609,N_11019,N_10897);
nand U11610 (N_11610,N_10575,N_10489);
or U11611 (N_11611,N_10924,N_11099);
or U11612 (N_11612,N_11169,N_10910);
xnor U11613 (N_11613,N_10667,N_11097);
nor U11614 (N_11614,N_10497,N_10618);
nor U11615 (N_11615,N_10786,N_10779);
nand U11616 (N_11616,N_10873,N_11189);
and U11617 (N_11617,N_10654,N_10787);
nand U11618 (N_11618,N_10871,N_11072);
or U11619 (N_11619,N_10478,N_10839);
and U11620 (N_11620,N_10663,N_10907);
nand U11621 (N_11621,N_11188,N_11122);
nand U11622 (N_11622,N_10873,N_11009);
or U11623 (N_11623,N_10951,N_10708);
and U11624 (N_11624,N_10884,N_11004);
or U11625 (N_11625,N_10589,N_10630);
and U11626 (N_11626,N_10409,N_11124);
or U11627 (N_11627,N_10657,N_10713);
nor U11628 (N_11628,N_10649,N_10892);
or U11629 (N_11629,N_10887,N_10706);
or U11630 (N_11630,N_10443,N_10619);
nand U11631 (N_11631,N_10525,N_10945);
nor U11632 (N_11632,N_10929,N_10408);
nor U11633 (N_11633,N_10426,N_10819);
nand U11634 (N_11634,N_10644,N_10955);
and U11635 (N_11635,N_10738,N_10544);
xor U11636 (N_11636,N_10891,N_10544);
or U11637 (N_11637,N_10813,N_10805);
nor U11638 (N_11638,N_10770,N_10568);
and U11639 (N_11639,N_10710,N_11162);
xor U11640 (N_11640,N_10900,N_10922);
and U11641 (N_11641,N_11057,N_11155);
and U11642 (N_11642,N_10628,N_10627);
and U11643 (N_11643,N_10540,N_10582);
and U11644 (N_11644,N_10604,N_11156);
nor U11645 (N_11645,N_10690,N_11042);
nand U11646 (N_11646,N_10816,N_11173);
or U11647 (N_11647,N_10874,N_10572);
or U11648 (N_11648,N_10559,N_10877);
nand U11649 (N_11649,N_10545,N_10957);
or U11650 (N_11650,N_10952,N_10497);
or U11651 (N_11651,N_10447,N_10936);
or U11652 (N_11652,N_11165,N_11017);
nor U11653 (N_11653,N_10941,N_10830);
nor U11654 (N_11654,N_11151,N_10448);
and U11655 (N_11655,N_11098,N_10526);
and U11656 (N_11656,N_10922,N_10721);
or U11657 (N_11657,N_10685,N_11160);
nor U11658 (N_11658,N_10660,N_10956);
nand U11659 (N_11659,N_10553,N_10868);
or U11660 (N_11660,N_10821,N_10520);
or U11661 (N_11661,N_10606,N_10704);
and U11662 (N_11662,N_10877,N_10684);
nor U11663 (N_11663,N_10668,N_10407);
and U11664 (N_11664,N_10450,N_10692);
nor U11665 (N_11665,N_10946,N_10905);
or U11666 (N_11666,N_10789,N_10463);
and U11667 (N_11667,N_10879,N_10715);
nand U11668 (N_11668,N_10841,N_10677);
or U11669 (N_11669,N_11074,N_10841);
and U11670 (N_11670,N_10561,N_10631);
nand U11671 (N_11671,N_10859,N_10976);
nand U11672 (N_11672,N_11162,N_11053);
and U11673 (N_11673,N_11000,N_11013);
nor U11674 (N_11674,N_11070,N_10523);
or U11675 (N_11675,N_10828,N_10665);
nor U11676 (N_11676,N_10516,N_10469);
nand U11677 (N_11677,N_10884,N_10970);
or U11678 (N_11678,N_11067,N_10871);
nand U11679 (N_11679,N_10532,N_10617);
and U11680 (N_11680,N_10557,N_10699);
nand U11681 (N_11681,N_10743,N_10963);
and U11682 (N_11682,N_10958,N_10981);
or U11683 (N_11683,N_10979,N_11086);
nand U11684 (N_11684,N_10723,N_11010);
and U11685 (N_11685,N_10450,N_10936);
or U11686 (N_11686,N_10965,N_10625);
nand U11687 (N_11687,N_10797,N_11181);
and U11688 (N_11688,N_10519,N_10998);
and U11689 (N_11689,N_10703,N_10543);
or U11690 (N_11690,N_10546,N_10917);
or U11691 (N_11691,N_10676,N_10967);
xor U11692 (N_11692,N_11057,N_11095);
and U11693 (N_11693,N_11095,N_11044);
nor U11694 (N_11694,N_10682,N_10797);
xor U11695 (N_11695,N_10614,N_11023);
and U11696 (N_11696,N_11095,N_11181);
or U11697 (N_11697,N_10747,N_10825);
or U11698 (N_11698,N_10695,N_11129);
and U11699 (N_11699,N_11049,N_10570);
and U11700 (N_11700,N_10591,N_10564);
or U11701 (N_11701,N_11056,N_10436);
nor U11702 (N_11702,N_10979,N_10492);
nand U11703 (N_11703,N_10647,N_11024);
or U11704 (N_11704,N_10928,N_10988);
or U11705 (N_11705,N_10563,N_10460);
or U11706 (N_11706,N_10971,N_10650);
or U11707 (N_11707,N_10935,N_11178);
or U11708 (N_11708,N_10725,N_10882);
nand U11709 (N_11709,N_10999,N_10941);
or U11710 (N_11710,N_11133,N_10750);
xor U11711 (N_11711,N_10447,N_10597);
nor U11712 (N_11712,N_11116,N_10721);
nor U11713 (N_11713,N_10542,N_11049);
nand U11714 (N_11714,N_11099,N_10987);
or U11715 (N_11715,N_10845,N_11082);
nand U11716 (N_11716,N_10509,N_10610);
nor U11717 (N_11717,N_11136,N_10798);
or U11718 (N_11718,N_10846,N_10719);
nor U11719 (N_11719,N_10968,N_10626);
and U11720 (N_11720,N_10732,N_10617);
nor U11721 (N_11721,N_11176,N_10403);
nor U11722 (N_11722,N_11026,N_11187);
nor U11723 (N_11723,N_10560,N_11174);
nor U11724 (N_11724,N_10834,N_10415);
nor U11725 (N_11725,N_10765,N_11179);
nor U11726 (N_11726,N_10573,N_10871);
or U11727 (N_11727,N_10838,N_10946);
or U11728 (N_11728,N_11073,N_10789);
nor U11729 (N_11729,N_10920,N_11074);
nor U11730 (N_11730,N_10618,N_10486);
nand U11731 (N_11731,N_10872,N_10760);
and U11732 (N_11732,N_11178,N_10501);
nor U11733 (N_11733,N_10918,N_11145);
nand U11734 (N_11734,N_10766,N_11151);
xor U11735 (N_11735,N_10833,N_10918);
nand U11736 (N_11736,N_10583,N_10741);
or U11737 (N_11737,N_10751,N_10945);
nand U11738 (N_11738,N_10693,N_10889);
and U11739 (N_11739,N_11124,N_10537);
and U11740 (N_11740,N_10883,N_11019);
nor U11741 (N_11741,N_10614,N_10982);
nor U11742 (N_11742,N_10683,N_10436);
or U11743 (N_11743,N_11020,N_11162);
or U11744 (N_11744,N_10875,N_10564);
nor U11745 (N_11745,N_10470,N_10800);
nand U11746 (N_11746,N_10814,N_10991);
and U11747 (N_11747,N_11058,N_10870);
nor U11748 (N_11748,N_10779,N_10530);
nand U11749 (N_11749,N_10865,N_11108);
or U11750 (N_11750,N_10944,N_10820);
nand U11751 (N_11751,N_10523,N_11079);
nand U11752 (N_11752,N_10449,N_11144);
nor U11753 (N_11753,N_11016,N_10413);
and U11754 (N_11754,N_10813,N_10633);
nand U11755 (N_11755,N_11079,N_10411);
nor U11756 (N_11756,N_10512,N_10788);
or U11757 (N_11757,N_10900,N_11110);
and U11758 (N_11758,N_10407,N_10751);
and U11759 (N_11759,N_11102,N_10420);
and U11760 (N_11760,N_10680,N_11106);
nand U11761 (N_11761,N_10629,N_10949);
or U11762 (N_11762,N_10750,N_10506);
nor U11763 (N_11763,N_11064,N_10621);
nor U11764 (N_11764,N_10633,N_10788);
nor U11765 (N_11765,N_10403,N_10813);
nand U11766 (N_11766,N_10966,N_10490);
and U11767 (N_11767,N_10740,N_10944);
nor U11768 (N_11768,N_10683,N_11106);
or U11769 (N_11769,N_11166,N_10807);
and U11770 (N_11770,N_11089,N_10400);
or U11771 (N_11771,N_10796,N_10763);
nand U11772 (N_11772,N_10826,N_10674);
nand U11773 (N_11773,N_10849,N_10425);
and U11774 (N_11774,N_10850,N_10605);
nand U11775 (N_11775,N_10824,N_10643);
nand U11776 (N_11776,N_10433,N_10803);
nor U11777 (N_11777,N_10890,N_10914);
nor U11778 (N_11778,N_10829,N_10698);
nor U11779 (N_11779,N_11170,N_10596);
nand U11780 (N_11780,N_10600,N_11127);
nor U11781 (N_11781,N_11166,N_11116);
nand U11782 (N_11782,N_10858,N_10576);
nand U11783 (N_11783,N_10759,N_10915);
nor U11784 (N_11784,N_10591,N_10752);
or U11785 (N_11785,N_10600,N_10707);
nand U11786 (N_11786,N_10713,N_10835);
and U11787 (N_11787,N_10998,N_10630);
nand U11788 (N_11788,N_10724,N_10831);
or U11789 (N_11789,N_10420,N_10751);
or U11790 (N_11790,N_10497,N_11039);
and U11791 (N_11791,N_10875,N_11158);
nand U11792 (N_11792,N_10712,N_10590);
and U11793 (N_11793,N_10779,N_10731);
nand U11794 (N_11794,N_10750,N_11095);
nor U11795 (N_11795,N_11164,N_11021);
nor U11796 (N_11796,N_10619,N_11048);
and U11797 (N_11797,N_10402,N_11189);
and U11798 (N_11798,N_11130,N_10427);
nor U11799 (N_11799,N_11145,N_10514);
and U11800 (N_11800,N_11132,N_10895);
and U11801 (N_11801,N_10715,N_10870);
and U11802 (N_11802,N_10478,N_10948);
nor U11803 (N_11803,N_11044,N_10748);
nand U11804 (N_11804,N_10936,N_10966);
nand U11805 (N_11805,N_10971,N_10812);
nor U11806 (N_11806,N_10755,N_10486);
and U11807 (N_11807,N_10880,N_10969);
or U11808 (N_11808,N_10512,N_11196);
nor U11809 (N_11809,N_10978,N_10540);
nor U11810 (N_11810,N_10637,N_11006);
nor U11811 (N_11811,N_11017,N_11194);
and U11812 (N_11812,N_10488,N_11150);
and U11813 (N_11813,N_10676,N_10874);
or U11814 (N_11814,N_11054,N_10714);
nor U11815 (N_11815,N_10506,N_10565);
and U11816 (N_11816,N_10562,N_10941);
and U11817 (N_11817,N_10592,N_10990);
nand U11818 (N_11818,N_10431,N_11083);
nand U11819 (N_11819,N_10910,N_10594);
nor U11820 (N_11820,N_10476,N_10473);
nand U11821 (N_11821,N_10709,N_10968);
and U11822 (N_11822,N_11055,N_10433);
or U11823 (N_11823,N_11170,N_10425);
and U11824 (N_11824,N_10455,N_10559);
nand U11825 (N_11825,N_10426,N_10561);
xor U11826 (N_11826,N_10475,N_10448);
or U11827 (N_11827,N_10507,N_10553);
or U11828 (N_11828,N_10859,N_10655);
and U11829 (N_11829,N_10723,N_10532);
or U11830 (N_11830,N_10429,N_10440);
nor U11831 (N_11831,N_10704,N_10456);
or U11832 (N_11832,N_11038,N_10514);
or U11833 (N_11833,N_11149,N_11125);
or U11834 (N_11834,N_10810,N_11013);
nand U11835 (N_11835,N_10926,N_10704);
and U11836 (N_11836,N_11117,N_10721);
nand U11837 (N_11837,N_10906,N_10602);
and U11838 (N_11838,N_10609,N_10686);
nand U11839 (N_11839,N_10706,N_10842);
and U11840 (N_11840,N_10721,N_10972);
nand U11841 (N_11841,N_10996,N_10815);
nand U11842 (N_11842,N_11102,N_10487);
nand U11843 (N_11843,N_10540,N_10771);
nand U11844 (N_11844,N_10607,N_10881);
nor U11845 (N_11845,N_10480,N_10895);
or U11846 (N_11846,N_10416,N_10984);
nand U11847 (N_11847,N_10615,N_10544);
and U11848 (N_11848,N_10587,N_10769);
nor U11849 (N_11849,N_10900,N_10793);
nor U11850 (N_11850,N_10505,N_10810);
and U11851 (N_11851,N_10844,N_10791);
and U11852 (N_11852,N_10417,N_11045);
or U11853 (N_11853,N_10508,N_10459);
nor U11854 (N_11854,N_10684,N_10660);
nor U11855 (N_11855,N_11081,N_11097);
nor U11856 (N_11856,N_10710,N_10768);
nor U11857 (N_11857,N_10464,N_10425);
nor U11858 (N_11858,N_11128,N_11144);
or U11859 (N_11859,N_10642,N_10728);
and U11860 (N_11860,N_11078,N_10496);
nor U11861 (N_11861,N_11027,N_10960);
nand U11862 (N_11862,N_10408,N_10638);
and U11863 (N_11863,N_10656,N_10439);
nor U11864 (N_11864,N_10882,N_11072);
nand U11865 (N_11865,N_10622,N_10530);
nand U11866 (N_11866,N_10567,N_10779);
nor U11867 (N_11867,N_10438,N_10817);
nor U11868 (N_11868,N_10790,N_10614);
nand U11869 (N_11869,N_10509,N_10825);
and U11870 (N_11870,N_10749,N_11199);
or U11871 (N_11871,N_10690,N_10679);
or U11872 (N_11872,N_10496,N_11128);
nand U11873 (N_11873,N_10526,N_10905);
nand U11874 (N_11874,N_10618,N_11151);
nor U11875 (N_11875,N_10606,N_10874);
and U11876 (N_11876,N_11060,N_10587);
nor U11877 (N_11877,N_10929,N_10875);
nand U11878 (N_11878,N_10815,N_10938);
and U11879 (N_11879,N_10635,N_10563);
and U11880 (N_11880,N_10559,N_10481);
nor U11881 (N_11881,N_10703,N_10795);
or U11882 (N_11882,N_10537,N_10902);
nand U11883 (N_11883,N_10456,N_10820);
nor U11884 (N_11884,N_10898,N_10548);
and U11885 (N_11885,N_11179,N_10786);
or U11886 (N_11886,N_10639,N_10682);
nor U11887 (N_11887,N_11179,N_10691);
nand U11888 (N_11888,N_10748,N_10875);
or U11889 (N_11889,N_10652,N_10420);
nand U11890 (N_11890,N_10867,N_10593);
and U11891 (N_11891,N_10525,N_10732);
nor U11892 (N_11892,N_10868,N_10985);
or U11893 (N_11893,N_10922,N_10647);
nand U11894 (N_11894,N_11030,N_10454);
or U11895 (N_11895,N_10509,N_10898);
nand U11896 (N_11896,N_11106,N_10859);
or U11897 (N_11897,N_10692,N_10502);
nor U11898 (N_11898,N_11068,N_10927);
nor U11899 (N_11899,N_11053,N_10563);
nor U11900 (N_11900,N_11067,N_11145);
and U11901 (N_11901,N_10673,N_10883);
and U11902 (N_11902,N_10745,N_10934);
and U11903 (N_11903,N_11120,N_10849);
and U11904 (N_11904,N_10446,N_11115);
and U11905 (N_11905,N_10635,N_10982);
or U11906 (N_11906,N_10662,N_10654);
nand U11907 (N_11907,N_10963,N_10503);
nand U11908 (N_11908,N_10789,N_10587);
or U11909 (N_11909,N_11095,N_10649);
nand U11910 (N_11910,N_10891,N_10774);
nor U11911 (N_11911,N_10844,N_10924);
and U11912 (N_11912,N_11069,N_10520);
or U11913 (N_11913,N_10880,N_10733);
nand U11914 (N_11914,N_10613,N_10725);
nand U11915 (N_11915,N_10500,N_10904);
or U11916 (N_11916,N_10450,N_11000);
or U11917 (N_11917,N_10697,N_10846);
or U11918 (N_11918,N_10581,N_10409);
nor U11919 (N_11919,N_10889,N_10997);
and U11920 (N_11920,N_10483,N_10582);
nand U11921 (N_11921,N_10843,N_10830);
nor U11922 (N_11922,N_10780,N_11134);
or U11923 (N_11923,N_11153,N_10742);
or U11924 (N_11924,N_10533,N_10893);
or U11925 (N_11925,N_10903,N_11035);
nor U11926 (N_11926,N_10782,N_11019);
nor U11927 (N_11927,N_10824,N_11086);
nand U11928 (N_11928,N_10480,N_11078);
nand U11929 (N_11929,N_10738,N_10803);
nor U11930 (N_11930,N_10708,N_10548);
or U11931 (N_11931,N_10417,N_10607);
or U11932 (N_11932,N_11040,N_11002);
nor U11933 (N_11933,N_11001,N_10465);
or U11934 (N_11934,N_10664,N_10885);
nor U11935 (N_11935,N_11162,N_10596);
and U11936 (N_11936,N_10450,N_10845);
and U11937 (N_11937,N_10675,N_10904);
and U11938 (N_11938,N_11049,N_10893);
nor U11939 (N_11939,N_10607,N_10573);
nor U11940 (N_11940,N_11049,N_10571);
or U11941 (N_11941,N_11009,N_10763);
or U11942 (N_11942,N_10739,N_10832);
or U11943 (N_11943,N_11016,N_11007);
or U11944 (N_11944,N_11038,N_10493);
nand U11945 (N_11945,N_10558,N_10702);
xor U11946 (N_11946,N_10478,N_10697);
nor U11947 (N_11947,N_10934,N_10599);
nand U11948 (N_11948,N_10896,N_10644);
or U11949 (N_11949,N_11069,N_10405);
or U11950 (N_11950,N_10458,N_10977);
or U11951 (N_11951,N_10783,N_10812);
and U11952 (N_11952,N_10431,N_10729);
or U11953 (N_11953,N_10467,N_10462);
or U11954 (N_11954,N_10610,N_11040);
or U11955 (N_11955,N_10451,N_10572);
and U11956 (N_11956,N_10758,N_10413);
or U11957 (N_11957,N_10529,N_10856);
and U11958 (N_11958,N_10656,N_10734);
xnor U11959 (N_11959,N_10952,N_10471);
nand U11960 (N_11960,N_10655,N_10814);
nand U11961 (N_11961,N_10671,N_10913);
or U11962 (N_11962,N_10484,N_10500);
xor U11963 (N_11963,N_11114,N_10647);
nor U11964 (N_11964,N_10513,N_10528);
nand U11965 (N_11965,N_11134,N_10888);
nor U11966 (N_11966,N_10625,N_11119);
or U11967 (N_11967,N_10629,N_10973);
or U11968 (N_11968,N_10961,N_11169);
or U11969 (N_11969,N_10826,N_11047);
or U11970 (N_11970,N_10864,N_10844);
nor U11971 (N_11971,N_10647,N_10909);
and U11972 (N_11972,N_11020,N_10580);
nand U11973 (N_11973,N_10521,N_11018);
or U11974 (N_11974,N_11183,N_10455);
nand U11975 (N_11975,N_10698,N_10926);
or U11976 (N_11976,N_10429,N_10897);
nand U11977 (N_11977,N_10523,N_11056);
nand U11978 (N_11978,N_11123,N_10795);
and U11979 (N_11979,N_11178,N_11110);
nand U11980 (N_11980,N_10647,N_10945);
and U11981 (N_11981,N_10577,N_10824);
or U11982 (N_11982,N_10597,N_10429);
and U11983 (N_11983,N_10423,N_11157);
nor U11984 (N_11984,N_11172,N_11090);
nand U11985 (N_11985,N_11082,N_10649);
nor U11986 (N_11986,N_10769,N_10676);
xor U11987 (N_11987,N_10736,N_10500);
or U11988 (N_11988,N_10998,N_10418);
or U11989 (N_11989,N_11131,N_10969);
or U11990 (N_11990,N_11119,N_10980);
or U11991 (N_11991,N_10837,N_10897);
nor U11992 (N_11992,N_10747,N_10736);
nor U11993 (N_11993,N_10636,N_10967);
and U11994 (N_11994,N_11018,N_10578);
nand U11995 (N_11995,N_10591,N_10489);
nand U11996 (N_11996,N_10985,N_11115);
nor U11997 (N_11997,N_10539,N_11087);
nand U11998 (N_11998,N_11024,N_10541);
or U11999 (N_11999,N_10744,N_10617);
or U12000 (N_12000,N_11299,N_11801);
nor U12001 (N_12001,N_11469,N_11525);
or U12002 (N_12002,N_11845,N_11473);
nor U12003 (N_12003,N_11269,N_11673);
nand U12004 (N_12004,N_11694,N_11701);
or U12005 (N_12005,N_11758,N_11677);
or U12006 (N_12006,N_11558,N_11867);
and U12007 (N_12007,N_11715,N_11557);
nor U12008 (N_12008,N_11748,N_11272);
nand U12009 (N_12009,N_11807,N_11967);
nand U12010 (N_12010,N_11309,N_11571);
xor U12011 (N_12011,N_11518,N_11257);
nor U12012 (N_12012,N_11608,N_11850);
and U12013 (N_12013,N_11851,N_11654);
or U12014 (N_12014,N_11592,N_11780);
nand U12015 (N_12015,N_11337,N_11759);
nand U12016 (N_12016,N_11708,N_11392);
or U12017 (N_12017,N_11636,N_11515);
or U12018 (N_12018,N_11933,N_11374);
and U12019 (N_12019,N_11767,N_11745);
nor U12020 (N_12020,N_11951,N_11735);
nand U12021 (N_12021,N_11600,N_11455);
or U12022 (N_12022,N_11417,N_11800);
or U12023 (N_12023,N_11764,N_11976);
nor U12024 (N_12024,N_11832,N_11458);
and U12025 (N_12025,N_11591,N_11354);
nand U12026 (N_12026,N_11603,N_11233);
or U12027 (N_12027,N_11516,N_11884);
xnor U12028 (N_12028,N_11987,N_11485);
nor U12029 (N_12029,N_11679,N_11754);
nand U12030 (N_12030,N_11366,N_11419);
or U12031 (N_12031,N_11833,N_11998);
and U12032 (N_12032,N_11903,N_11864);
nor U12033 (N_12033,N_11830,N_11357);
nor U12034 (N_12034,N_11385,N_11956);
and U12035 (N_12035,N_11983,N_11364);
nand U12036 (N_12036,N_11295,N_11939);
or U12037 (N_12037,N_11893,N_11911);
nand U12038 (N_12038,N_11883,N_11649);
or U12039 (N_12039,N_11925,N_11323);
and U12040 (N_12040,N_11420,N_11245);
nor U12041 (N_12041,N_11293,N_11820);
nor U12042 (N_12042,N_11443,N_11535);
nor U12043 (N_12043,N_11424,N_11502);
or U12044 (N_12044,N_11457,N_11888);
or U12045 (N_12045,N_11260,N_11234);
and U12046 (N_12046,N_11235,N_11493);
and U12047 (N_12047,N_11492,N_11796);
nand U12048 (N_12048,N_11853,N_11210);
and U12049 (N_12049,N_11223,N_11786);
and U12050 (N_12050,N_11330,N_11549);
nor U12051 (N_12051,N_11988,N_11497);
xor U12052 (N_12052,N_11878,N_11769);
and U12053 (N_12053,N_11824,N_11686);
nand U12054 (N_12054,N_11952,N_11938);
nand U12055 (N_12055,N_11890,N_11248);
or U12056 (N_12056,N_11746,N_11844);
nand U12057 (N_12057,N_11537,N_11669);
or U12058 (N_12058,N_11821,N_11563);
nor U12059 (N_12059,N_11719,N_11478);
and U12060 (N_12060,N_11255,N_11924);
or U12061 (N_12061,N_11504,N_11705);
nand U12062 (N_12062,N_11740,N_11437);
or U12063 (N_12063,N_11281,N_11509);
nand U12064 (N_12064,N_11250,N_11781);
nor U12065 (N_12065,N_11348,N_11852);
nand U12066 (N_12066,N_11367,N_11476);
or U12067 (N_12067,N_11288,N_11263);
or U12068 (N_12068,N_11662,N_11750);
or U12069 (N_12069,N_11962,N_11201);
xor U12070 (N_12070,N_11533,N_11810);
nor U12071 (N_12071,N_11660,N_11401);
nand U12072 (N_12072,N_11847,N_11658);
nand U12073 (N_12073,N_11283,N_11427);
nor U12074 (N_12074,N_11463,N_11752);
or U12075 (N_12075,N_11287,N_11728);
nand U12076 (N_12076,N_11363,N_11615);
nor U12077 (N_12077,N_11991,N_11241);
or U12078 (N_12078,N_11650,N_11266);
nor U12079 (N_12079,N_11731,N_11441);
or U12080 (N_12080,N_11477,N_11564);
xor U12081 (N_12081,N_11400,N_11913);
or U12082 (N_12082,N_11739,N_11904);
nand U12083 (N_12083,N_11944,N_11655);
nor U12084 (N_12084,N_11702,N_11928);
and U12085 (N_12085,N_11433,N_11683);
nand U12086 (N_12086,N_11247,N_11232);
and U12087 (N_12087,N_11804,N_11413);
nor U12088 (N_12088,N_11303,N_11953);
nand U12089 (N_12089,N_11256,N_11465);
nand U12090 (N_12090,N_11484,N_11858);
nor U12091 (N_12091,N_11547,N_11560);
nor U12092 (N_12092,N_11506,N_11816);
or U12093 (N_12093,N_11430,N_11787);
nor U12094 (N_12094,N_11803,N_11588);
or U12095 (N_12095,N_11582,N_11992);
nor U12096 (N_12096,N_11579,N_11342);
and U12097 (N_12097,N_11320,N_11448);
and U12098 (N_12098,N_11665,N_11369);
nor U12099 (N_12099,N_11524,N_11207);
nand U12100 (N_12100,N_11755,N_11865);
nand U12101 (N_12101,N_11545,N_11859);
nand U12102 (N_12102,N_11877,N_11365);
nand U12103 (N_12103,N_11813,N_11325);
or U12104 (N_12104,N_11438,N_11959);
or U12105 (N_12105,N_11934,N_11494);
or U12106 (N_12106,N_11301,N_11598);
or U12107 (N_12107,N_11499,N_11627);
and U12108 (N_12108,N_11411,N_11912);
nand U12109 (N_12109,N_11559,N_11450);
nand U12110 (N_12110,N_11467,N_11874);
nor U12111 (N_12111,N_11838,N_11202);
or U12112 (N_12112,N_11379,N_11707);
nand U12113 (N_12113,N_11989,N_11773);
nand U12114 (N_12114,N_11611,N_11723);
nand U12115 (N_12115,N_11872,N_11425);
and U12116 (N_12116,N_11416,N_11397);
nand U12117 (N_12117,N_11358,N_11968);
and U12118 (N_12118,N_11936,N_11927);
nor U12119 (N_12119,N_11355,N_11575);
or U12120 (N_12120,N_11314,N_11870);
or U12121 (N_12121,N_11652,N_11335);
nor U12122 (N_12122,N_11389,N_11561);
and U12123 (N_12123,N_11251,N_11866);
nor U12124 (N_12124,N_11242,N_11880);
and U12125 (N_12125,N_11979,N_11405);
and U12126 (N_12126,N_11311,N_11788);
nand U12127 (N_12127,N_11646,N_11380);
or U12128 (N_12128,N_11921,N_11324);
xnor U12129 (N_12129,N_11664,N_11666);
nor U12130 (N_12130,N_11902,N_11737);
nand U12131 (N_12131,N_11729,N_11923);
and U12132 (N_12132,N_11698,N_11586);
nand U12133 (N_12133,N_11344,N_11971);
nor U12134 (N_12134,N_11640,N_11969);
and U12135 (N_12135,N_11790,N_11648);
nand U12136 (N_12136,N_11602,N_11327);
or U12137 (N_12137,N_11753,N_11595);
or U12138 (N_12138,N_11584,N_11695);
nor U12139 (N_12139,N_11244,N_11583);
and U12140 (N_12140,N_11929,N_11328);
nand U12141 (N_12141,N_11580,N_11625);
nor U12142 (N_12142,N_11633,N_11846);
and U12143 (N_12143,N_11200,N_11262);
and U12144 (N_12144,N_11490,N_11548);
nand U12145 (N_12145,N_11208,N_11520);
or U12146 (N_12146,N_11970,N_11749);
or U12147 (N_12147,N_11697,N_11390);
and U12148 (N_12148,N_11512,N_11205);
nand U12149 (N_12149,N_11229,N_11534);
nor U12150 (N_12150,N_11356,N_11487);
nor U12151 (N_12151,N_11577,N_11370);
and U12152 (N_12152,N_11578,N_11727);
nor U12153 (N_12153,N_11763,N_11222);
nand U12154 (N_12154,N_11860,N_11892);
nor U12155 (N_12155,N_11213,N_11285);
and U12156 (N_12156,N_11896,N_11218);
and U12157 (N_12157,N_11814,N_11840);
nor U12158 (N_12158,N_11453,N_11553);
nor U12159 (N_12159,N_11291,N_11239);
or U12160 (N_12160,N_11491,N_11774);
or U12161 (N_12161,N_11460,N_11961);
and U12162 (N_12162,N_11542,N_11212);
and U12163 (N_12163,N_11641,N_11604);
nand U12164 (N_12164,N_11576,N_11797);
nand U12165 (N_12165,N_11624,N_11556);
nor U12166 (N_12166,N_11990,N_11711);
and U12167 (N_12167,N_11947,N_11514);
nand U12168 (N_12168,N_11415,N_11696);
nor U12169 (N_12169,N_11862,N_11435);
and U12170 (N_12170,N_11606,N_11307);
nor U12171 (N_12171,N_11521,N_11778);
nor U12172 (N_12172,N_11730,N_11206);
nor U12173 (N_12173,N_11368,N_11724);
nand U12174 (N_12174,N_11720,N_11926);
or U12175 (N_12175,N_11551,N_11217);
or U12176 (N_12176,N_11498,N_11289);
nand U12177 (N_12177,N_11802,N_11446);
and U12178 (N_12178,N_11805,N_11350);
nor U12179 (N_12179,N_11265,N_11891);
or U12180 (N_12180,N_11326,N_11985);
and U12181 (N_12181,N_11734,N_11981);
or U12182 (N_12182,N_11294,N_11334);
nand U12183 (N_12183,N_11538,N_11343);
nor U12184 (N_12184,N_11993,N_11554);
nor U12185 (N_12185,N_11541,N_11345);
or U12186 (N_12186,N_11622,N_11569);
and U12187 (N_12187,N_11676,N_11612);
and U12188 (N_12188,N_11259,N_11657);
nand U12189 (N_12189,N_11261,N_11974);
or U12190 (N_12190,N_11230,N_11587);
nand U12191 (N_12191,N_11359,N_11589);
nor U12192 (N_12192,N_11226,N_11889);
nand U12193 (N_12193,N_11274,N_11529);
nor U12194 (N_12194,N_11333,N_11918);
nor U12195 (N_12195,N_11381,N_11744);
and U12196 (N_12196,N_11388,N_11732);
nand U12197 (N_12197,N_11211,N_11237);
or U12198 (N_12198,N_11378,N_11596);
and U12199 (N_12199,N_11312,N_11482);
and U12200 (N_12200,N_11680,N_11687);
or U12201 (N_12201,N_11225,N_11428);
or U12202 (N_12202,N_11815,N_11496);
nand U12203 (N_12203,N_11656,N_11619);
and U12204 (N_12204,N_11812,N_11631);
nor U12205 (N_12205,N_11887,N_11785);
nand U12206 (N_12206,N_11422,N_11318);
nor U12207 (N_12207,N_11826,N_11886);
and U12208 (N_12208,N_11643,N_11672);
nor U12209 (N_12209,N_11329,N_11562);
nand U12210 (N_12210,N_11882,N_11937);
or U12211 (N_12211,N_11278,N_11224);
and U12212 (N_12212,N_11614,N_11965);
nand U12213 (N_12213,N_11331,N_11638);
nor U12214 (N_12214,N_11771,N_11500);
or U12215 (N_12215,N_11372,N_11308);
nor U12216 (N_12216,N_11900,N_11338);
and U12217 (N_12217,N_11404,N_11645);
and U12218 (N_12218,N_11620,N_11336);
nor U12219 (N_12219,N_11565,N_11907);
nand U12220 (N_12220,N_11818,N_11834);
nand U12221 (N_12221,N_11945,N_11943);
and U12222 (N_12222,N_11635,N_11402);
nand U12223 (N_12223,N_11352,N_11382);
or U12224 (N_12224,N_11670,N_11517);
and U12225 (N_12225,N_11827,N_11470);
nand U12226 (N_12226,N_11546,N_11957);
and U12227 (N_12227,N_11848,N_11973);
nand U12228 (N_12228,N_11948,N_11488);
and U12229 (N_12229,N_11667,N_11616);
nand U12230 (N_12230,N_11462,N_11637);
and U12231 (N_12231,N_11733,N_11710);
nor U12232 (N_12232,N_11383,N_11568);
nor U12233 (N_12233,N_11501,N_11572);
nand U12234 (N_12234,N_11914,N_11340);
nand U12235 (N_12235,N_11980,N_11747);
and U12236 (N_12236,N_11941,N_11240);
nand U12237 (N_12237,N_11837,N_11573);
nand U12238 (N_12238,N_11714,N_11618);
nor U12239 (N_12239,N_11445,N_11935);
nor U12240 (N_12240,N_11270,N_11316);
and U12241 (N_12241,N_11811,N_11214);
and U12242 (N_12242,N_11332,N_11699);
or U12243 (N_12243,N_11439,N_11647);
nor U12244 (N_12244,N_11671,N_11854);
and U12245 (N_12245,N_11204,N_11339);
nand U12246 (N_12246,N_11298,N_11915);
and U12247 (N_12247,N_11599,N_11607);
and U12248 (N_12248,N_11597,N_11403);
and U12249 (N_12249,N_11609,N_11682);
nand U12250 (N_12250,N_11958,N_11977);
and U12251 (N_12251,N_11271,N_11685);
nand U12252 (N_12252,N_11258,N_11267);
or U12253 (N_12253,N_11955,N_11601);
nand U12254 (N_12254,N_11431,N_11806);
nand U12255 (N_12255,N_11661,N_11489);
and U12256 (N_12256,N_11362,N_11984);
nand U12257 (N_12257,N_11628,N_11203);
nand U12258 (N_12258,N_11505,N_11508);
nor U12259 (N_12259,N_11319,N_11550);
nand U12260 (N_12260,N_11282,N_11447);
xor U12261 (N_12261,N_11995,N_11290);
and U12262 (N_12262,N_11280,N_11898);
and U12263 (N_12263,N_11444,N_11279);
nor U12264 (N_12264,N_11651,N_11304);
nand U12265 (N_12265,N_11238,N_11297);
nor U12266 (N_12266,N_11770,N_11653);
nand U12267 (N_12267,N_11906,N_11527);
or U12268 (N_12268,N_11585,N_11963);
nor U12269 (N_12269,N_11442,N_11613);
xnor U12270 (N_12270,N_11522,N_11808);
and U12271 (N_12271,N_11684,N_11227);
or U12272 (N_12272,N_11691,N_11775);
nand U12273 (N_12273,N_11881,N_11885);
nor U12274 (N_12274,N_11373,N_11982);
nor U12275 (N_12275,N_11253,N_11794);
nand U12276 (N_12276,N_11451,N_11414);
nor U12277 (N_12277,N_11454,N_11766);
nor U12278 (N_12278,N_11986,N_11570);
nor U12279 (N_12279,N_11429,N_11756);
or U12280 (N_12280,N_11581,N_11789);
nor U12281 (N_12281,N_11709,N_11706);
or U12282 (N_12282,N_11408,N_11317);
or U12283 (N_12283,N_11922,N_11792);
and U12284 (N_12284,N_11975,N_11386);
and U12285 (N_12285,N_11341,N_11371);
nand U12286 (N_12286,N_11966,N_11793);
nor U12287 (N_12287,N_11964,N_11639);
nor U12288 (N_12288,N_11879,N_11762);
and U12289 (N_12289,N_11784,N_11736);
or U12290 (N_12290,N_11481,N_11276);
nand U12291 (N_12291,N_11346,N_11871);
nand U12292 (N_12292,N_11856,N_11432);
nor U12293 (N_12293,N_11668,N_11249);
nand U12294 (N_12294,N_11574,N_11817);
nand U12295 (N_12295,N_11940,N_11632);
nor U12296 (N_12296,N_11321,N_11799);
nor U12297 (N_12297,N_11690,N_11423);
nor U12298 (N_12298,N_11776,N_11868);
nand U12299 (N_12299,N_11306,N_11917);
nor U12300 (N_12300,N_11209,N_11910);
nor U12301 (N_12301,N_11978,N_11519);
nor U12302 (N_12302,N_11539,N_11349);
or U12303 (N_12303,N_11216,N_11839);
and U12304 (N_12304,N_11757,N_11531);
nand U12305 (N_12305,N_11930,N_11828);
and U12306 (N_12306,N_11809,N_11296);
nand U12307 (N_12307,N_11836,N_11721);
nor U12308 (N_12308,N_11268,N_11741);
nor U12309 (N_12309,N_11946,N_11421);
and U12310 (N_12310,N_11899,N_11264);
nor U12311 (N_12311,N_11566,N_11782);
or U12312 (N_12312,N_11543,N_11452);
and U12313 (N_12313,N_11742,N_11972);
and U12314 (N_12314,N_11221,N_11876);
or U12315 (N_12315,N_11722,N_11725);
and U12316 (N_12316,N_11693,N_11440);
or U12317 (N_12317,N_11610,N_11920);
and U12318 (N_12318,N_11475,N_11310);
nor U12319 (N_12319,N_11456,N_11406);
or U12320 (N_12320,N_11219,N_11841);
nor U12321 (N_12321,N_11396,N_11617);
nand U12322 (N_12322,N_11875,N_11393);
and U12323 (N_12323,N_11712,N_11916);
nor U12324 (N_12324,N_11526,N_11302);
nor U12325 (N_12325,N_11630,N_11300);
and U12326 (N_12326,N_11426,N_11954);
nor U12327 (N_12327,N_11642,N_11399);
nand U12328 (N_12328,N_11384,N_11873);
nor U12329 (N_12329,N_11688,N_11459);
and U12330 (N_12330,N_11623,N_11777);
nor U12331 (N_12331,N_11252,N_11798);
nand U12332 (N_12332,N_11908,N_11387);
nand U12333 (N_12333,N_11464,N_11663);
nor U12334 (N_12334,N_11919,N_11700);
or U12335 (N_12335,N_11243,N_11761);
nand U12336 (N_12336,N_11552,N_11472);
and U12337 (N_12337,N_11305,N_11743);
nor U12338 (N_12338,N_11825,N_11996);
nand U12339 (N_12339,N_11468,N_11905);
and U12340 (N_12340,N_11949,N_11674);
or U12341 (N_12341,N_11277,N_11829);
and U12342 (N_12342,N_11461,N_11360);
and U12343 (N_12343,N_11689,N_11412);
or U12344 (N_12344,N_11760,N_11855);
or U12345 (N_12345,N_11997,N_11449);
nand U12346 (N_12346,N_11254,N_11292);
nand U12347 (N_12347,N_11536,N_11483);
nand U12348 (N_12348,N_11897,N_11895);
nor U12349 (N_12349,N_11849,N_11823);
nor U12350 (N_12350,N_11284,N_11495);
and U12351 (N_12351,N_11718,N_11474);
nand U12352 (N_12352,N_11713,N_11391);
or U12353 (N_12353,N_11626,N_11351);
nand U12354 (N_12354,N_11772,N_11377);
nor U12355 (N_12355,N_11418,N_11842);
nand U12356 (N_12356,N_11681,N_11479);
and U12357 (N_12357,N_11822,N_11831);
nor U12358 (N_12358,N_11703,N_11932);
or U12359 (N_12359,N_11960,N_11644);
nor U12360 (N_12360,N_11395,N_11894);
and U12361 (N_12361,N_11909,N_11942);
and U12362 (N_12362,N_11594,N_11523);
nand U12363 (N_12363,N_11738,N_11791);
and U12364 (N_12364,N_11220,N_11315);
and U12365 (N_12365,N_11795,N_11634);
nor U12366 (N_12366,N_11704,N_11322);
nand U12367 (N_12367,N_11931,N_11510);
or U12368 (N_12368,N_11353,N_11273);
nor U12369 (N_12369,N_11361,N_11434);
and U12370 (N_12370,N_11863,N_11228);
and U12371 (N_12371,N_11950,N_11629);
or U12372 (N_12372,N_11567,N_11236);
nor U12373 (N_12373,N_11590,N_11751);
nand U12374 (N_12374,N_11275,N_11675);
xnor U12375 (N_12375,N_11768,N_11286);
and U12376 (N_12376,N_11716,N_11466);
nand U12377 (N_12377,N_11835,N_11765);
nor U12378 (N_12378,N_11869,N_11659);
and U12379 (N_12379,N_11605,N_11528);
or U12380 (N_12380,N_11503,N_11394);
nand U12381 (N_12381,N_11901,N_11215);
or U12382 (N_12382,N_11313,N_11779);
nand U12383 (N_12383,N_11783,N_11375);
and U12384 (N_12384,N_11398,N_11376);
nand U12385 (N_12385,N_11593,N_11544);
and U12386 (N_12386,N_11726,N_11480);
nand U12387 (N_12387,N_11513,N_11717);
and U12388 (N_12388,N_11555,N_11471);
nand U12389 (N_12389,N_11407,N_11999);
or U12390 (N_12390,N_11994,N_11843);
nand U12391 (N_12391,N_11861,N_11678);
nor U12392 (N_12392,N_11409,N_11347);
nand U12393 (N_12393,N_11511,N_11692);
and U12394 (N_12394,N_11819,N_11246);
and U12395 (N_12395,N_11436,N_11486);
nor U12396 (N_12396,N_11857,N_11530);
or U12397 (N_12397,N_11231,N_11621);
or U12398 (N_12398,N_11532,N_11410);
nor U12399 (N_12399,N_11540,N_11507);
or U12400 (N_12400,N_11750,N_11484);
nor U12401 (N_12401,N_11410,N_11731);
and U12402 (N_12402,N_11896,N_11322);
or U12403 (N_12403,N_11466,N_11729);
and U12404 (N_12404,N_11204,N_11243);
or U12405 (N_12405,N_11579,N_11521);
and U12406 (N_12406,N_11344,N_11927);
nor U12407 (N_12407,N_11387,N_11723);
nor U12408 (N_12408,N_11330,N_11308);
nor U12409 (N_12409,N_11923,N_11966);
nor U12410 (N_12410,N_11781,N_11370);
nand U12411 (N_12411,N_11401,N_11857);
nand U12412 (N_12412,N_11911,N_11606);
nor U12413 (N_12413,N_11771,N_11889);
and U12414 (N_12414,N_11766,N_11649);
nand U12415 (N_12415,N_11210,N_11725);
or U12416 (N_12416,N_11953,N_11726);
and U12417 (N_12417,N_11568,N_11665);
or U12418 (N_12418,N_11906,N_11400);
and U12419 (N_12419,N_11599,N_11529);
or U12420 (N_12420,N_11992,N_11237);
nor U12421 (N_12421,N_11439,N_11999);
or U12422 (N_12422,N_11827,N_11220);
or U12423 (N_12423,N_11792,N_11633);
nor U12424 (N_12424,N_11886,N_11360);
and U12425 (N_12425,N_11272,N_11715);
nor U12426 (N_12426,N_11882,N_11927);
and U12427 (N_12427,N_11601,N_11250);
xnor U12428 (N_12428,N_11210,N_11341);
and U12429 (N_12429,N_11894,N_11587);
nand U12430 (N_12430,N_11965,N_11992);
or U12431 (N_12431,N_11402,N_11479);
nor U12432 (N_12432,N_11772,N_11886);
and U12433 (N_12433,N_11822,N_11367);
nand U12434 (N_12434,N_11617,N_11470);
and U12435 (N_12435,N_11604,N_11566);
and U12436 (N_12436,N_11975,N_11277);
nor U12437 (N_12437,N_11750,N_11225);
nand U12438 (N_12438,N_11862,N_11264);
or U12439 (N_12439,N_11306,N_11245);
nand U12440 (N_12440,N_11833,N_11284);
and U12441 (N_12441,N_11329,N_11909);
xor U12442 (N_12442,N_11204,N_11837);
or U12443 (N_12443,N_11898,N_11259);
or U12444 (N_12444,N_11768,N_11512);
nand U12445 (N_12445,N_11588,N_11430);
nand U12446 (N_12446,N_11656,N_11308);
and U12447 (N_12447,N_11630,N_11220);
and U12448 (N_12448,N_11306,N_11476);
nand U12449 (N_12449,N_11805,N_11840);
or U12450 (N_12450,N_11547,N_11829);
nor U12451 (N_12451,N_11928,N_11985);
and U12452 (N_12452,N_11674,N_11293);
and U12453 (N_12453,N_11805,N_11780);
nor U12454 (N_12454,N_11577,N_11276);
and U12455 (N_12455,N_11732,N_11855);
or U12456 (N_12456,N_11332,N_11274);
nor U12457 (N_12457,N_11609,N_11426);
or U12458 (N_12458,N_11763,N_11363);
nand U12459 (N_12459,N_11776,N_11652);
and U12460 (N_12460,N_11435,N_11712);
and U12461 (N_12461,N_11228,N_11385);
and U12462 (N_12462,N_11801,N_11514);
or U12463 (N_12463,N_11367,N_11649);
and U12464 (N_12464,N_11473,N_11604);
or U12465 (N_12465,N_11295,N_11471);
and U12466 (N_12466,N_11498,N_11265);
nand U12467 (N_12467,N_11668,N_11860);
nor U12468 (N_12468,N_11963,N_11571);
and U12469 (N_12469,N_11262,N_11248);
nor U12470 (N_12470,N_11642,N_11590);
nor U12471 (N_12471,N_11677,N_11696);
and U12472 (N_12472,N_11959,N_11743);
and U12473 (N_12473,N_11271,N_11268);
nand U12474 (N_12474,N_11204,N_11892);
or U12475 (N_12475,N_11390,N_11662);
nand U12476 (N_12476,N_11205,N_11501);
nand U12477 (N_12477,N_11776,N_11244);
nor U12478 (N_12478,N_11679,N_11927);
nor U12479 (N_12479,N_11804,N_11275);
or U12480 (N_12480,N_11627,N_11811);
or U12481 (N_12481,N_11837,N_11217);
and U12482 (N_12482,N_11696,N_11447);
nand U12483 (N_12483,N_11471,N_11760);
or U12484 (N_12484,N_11795,N_11901);
and U12485 (N_12485,N_11938,N_11507);
and U12486 (N_12486,N_11999,N_11251);
and U12487 (N_12487,N_11903,N_11274);
or U12488 (N_12488,N_11859,N_11543);
xor U12489 (N_12489,N_11834,N_11415);
nor U12490 (N_12490,N_11954,N_11773);
or U12491 (N_12491,N_11976,N_11515);
nand U12492 (N_12492,N_11878,N_11639);
nand U12493 (N_12493,N_11649,N_11467);
nand U12494 (N_12494,N_11379,N_11731);
nand U12495 (N_12495,N_11784,N_11888);
and U12496 (N_12496,N_11292,N_11963);
nor U12497 (N_12497,N_11654,N_11591);
nand U12498 (N_12498,N_11356,N_11354);
nand U12499 (N_12499,N_11400,N_11998);
nor U12500 (N_12500,N_11576,N_11795);
nand U12501 (N_12501,N_11394,N_11785);
nand U12502 (N_12502,N_11536,N_11801);
nand U12503 (N_12503,N_11330,N_11273);
nor U12504 (N_12504,N_11274,N_11700);
nor U12505 (N_12505,N_11284,N_11949);
nor U12506 (N_12506,N_11382,N_11403);
or U12507 (N_12507,N_11701,N_11853);
nand U12508 (N_12508,N_11601,N_11548);
and U12509 (N_12509,N_11250,N_11318);
and U12510 (N_12510,N_11508,N_11991);
or U12511 (N_12511,N_11445,N_11283);
or U12512 (N_12512,N_11905,N_11657);
nand U12513 (N_12513,N_11698,N_11543);
and U12514 (N_12514,N_11743,N_11255);
nand U12515 (N_12515,N_11868,N_11318);
nor U12516 (N_12516,N_11923,N_11751);
nor U12517 (N_12517,N_11592,N_11325);
nand U12518 (N_12518,N_11761,N_11318);
or U12519 (N_12519,N_11229,N_11903);
xnor U12520 (N_12520,N_11565,N_11695);
nor U12521 (N_12521,N_11647,N_11889);
and U12522 (N_12522,N_11412,N_11245);
nor U12523 (N_12523,N_11583,N_11846);
or U12524 (N_12524,N_11415,N_11717);
and U12525 (N_12525,N_11677,N_11561);
nor U12526 (N_12526,N_11992,N_11757);
and U12527 (N_12527,N_11874,N_11937);
or U12528 (N_12528,N_11889,N_11696);
or U12529 (N_12529,N_11703,N_11717);
nand U12530 (N_12530,N_11943,N_11452);
nand U12531 (N_12531,N_11667,N_11393);
nor U12532 (N_12532,N_11421,N_11294);
and U12533 (N_12533,N_11831,N_11941);
or U12534 (N_12534,N_11950,N_11489);
nand U12535 (N_12535,N_11597,N_11902);
and U12536 (N_12536,N_11761,N_11568);
xor U12537 (N_12537,N_11657,N_11296);
nor U12538 (N_12538,N_11662,N_11987);
nand U12539 (N_12539,N_11541,N_11659);
nor U12540 (N_12540,N_11380,N_11288);
and U12541 (N_12541,N_11521,N_11992);
and U12542 (N_12542,N_11494,N_11763);
xnor U12543 (N_12543,N_11532,N_11342);
nand U12544 (N_12544,N_11944,N_11694);
or U12545 (N_12545,N_11744,N_11331);
nor U12546 (N_12546,N_11247,N_11555);
and U12547 (N_12547,N_11891,N_11282);
nor U12548 (N_12548,N_11884,N_11353);
and U12549 (N_12549,N_11664,N_11458);
or U12550 (N_12550,N_11466,N_11557);
nor U12551 (N_12551,N_11478,N_11503);
nand U12552 (N_12552,N_11966,N_11761);
or U12553 (N_12553,N_11227,N_11601);
nand U12554 (N_12554,N_11515,N_11960);
and U12555 (N_12555,N_11732,N_11598);
nor U12556 (N_12556,N_11895,N_11806);
nor U12557 (N_12557,N_11679,N_11747);
and U12558 (N_12558,N_11479,N_11563);
or U12559 (N_12559,N_11754,N_11716);
nand U12560 (N_12560,N_11694,N_11275);
nand U12561 (N_12561,N_11906,N_11705);
nor U12562 (N_12562,N_11277,N_11982);
or U12563 (N_12563,N_11776,N_11855);
nor U12564 (N_12564,N_11200,N_11202);
nor U12565 (N_12565,N_11528,N_11723);
or U12566 (N_12566,N_11404,N_11969);
nand U12567 (N_12567,N_11572,N_11560);
nand U12568 (N_12568,N_11447,N_11441);
nor U12569 (N_12569,N_11584,N_11526);
nor U12570 (N_12570,N_11342,N_11254);
and U12571 (N_12571,N_11207,N_11639);
xnor U12572 (N_12572,N_11553,N_11686);
or U12573 (N_12573,N_11367,N_11753);
nand U12574 (N_12574,N_11548,N_11772);
and U12575 (N_12575,N_11810,N_11355);
nand U12576 (N_12576,N_11259,N_11294);
nand U12577 (N_12577,N_11484,N_11989);
nor U12578 (N_12578,N_11704,N_11392);
nor U12579 (N_12579,N_11524,N_11817);
or U12580 (N_12580,N_11219,N_11437);
nand U12581 (N_12581,N_11977,N_11448);
and U12582 (N_12582,N_11351,N_11263);
xnor U12583 (N_12583,N_11916,N_11615);
or U12584 (N_12584,N_11632,N_11783);
nor U12585 (N_12585,N_11965,N_11353);
nor U12586 (N_12586,N_11634,N_11299);
and U12587 (N_12587,N_11969,N_11405);
nor U12588 (N_12588,N_11422,N_11254);
nor U12589 (N_12589,N_11263,N_11444);
nand U12590 (N_12590,N_11998,N_11700);
or U12591 (N_12591,N_11584,N_11724);
nand U12592 (N_12592,N_11854,N_11222);
nand U12593 (N_12593,N_11654,N_11408);
and U12594 (N_12594,N_11658,N_11796);
nand U12595 (N_12595,N_11675,N_11837);
nand U12596 (N_12596,N_11691,N_11664);
and U12597 (N_12597,N_11703,N_11462);
and U12598 (N_12598,N_11573,N_11791);
or U12599 (N_12599,N_11778,N_11503);
nand U12600 (N_12600,N_11385,N_11963);
nor U12601 (N_12601,N_11265,N_11812);
and U12602 (N_12602,N_11765,N_11924);
nor U12603 (N_12603,N_11617,N_11564);
nand U12604 (N_12604,N_11255,N_11963);
xor U12605 (N_12605,N_11244,N_11788);
and U12606 (N_12606,N_11755,N_11674);
nor U12607 (N_12607,N_11277,N_11624);
or U12608 (N_12608,N_11684,N_11481);
and U12609 (N_12609,N_11769,N_11583);
or U12610 (N_12610,N_11482,N_11369);
or U12611 (N_12611,N_11969,N_11214);
nand U12612 (N_12612,N_11599,N_11566);
or U12613 (N_12613,N_11479,N_11664);
or U12614 (N_12614,N_11838,N_11953);
nand U12615 (N_12615,N_11699,N_11363);
or U12616 (N_12616,N_11319,N_11333);
nand U12617 (N_12617,N_11889,N_11322);
or U12618 (N_12618,N_11673,N_11689);
or U12619 (N_12619,N_11974,N_11625);
and U12620 (N_12620,N_11737,N_11647);
and U12621 (N_12621,N_11872,N_11200);
nand U12622 (N_12622,N_11460,N_11283);
nand U12623 (N_12623,N_11232,N_11223);
nor U12624 (N_12624,N_11430,N_11481);
or U12625 (N_12625,N_11281,N_11571);
xnor U12626 (N_12626,N_11243,N_11699);
or U12627 (N_12627,N_11904,N_11209);
or U12628 (N_12628,N_11977,N_11481);
nand U12629 (N_12629,N_11654,N_11838);
and U12630 (N_12630,N_11666,N_11371);
or U12631 (N_12631,N_11913,N_11766);
or U12632 (N_12632,N_11608,N_11982);
nand U12633 (N_12633,N_11297,N_11345);
nand U12634 (N_12634,N_11972,N_11903);
nor U12635 (N_12635,N_11696,N_11382);
or U12636 (N_12636,N_11595,N_11665);
nor U12637 (N_12637,N_11883,N_11291);
or U12638 (N_12638,N_11512,N_11266);
nand U12639 (N_12639,N_11534,N_11745);
nor U12640 (N_12640,N_11228,N_11474);
or U12641 (N_12641,N_11354,N_11468);
or U12642 (N_12642,N_11456,N_11349);
nand U12643 (N_12643,N_11426,N_11583);
nand U12644 (N_12644,N_11246,N_11468);
xor U12645 (N_12645,N_11236,N_11741);
and U12646 (N_12646,N_11600,N_11598);
or U12647 (N_12647,N_11878,N_11750);
nand U12648 (N_12648,N_11824,N_11412);
or U12649 (N_12649,N_11846,N_11318);
nand U12650 (N_12650,N_11519,N_11466);
or U12651 (N_12651,N_11830,N_11506);
and U12652 (N_12652,N_11598,N_11512);
or U12653 (N_12653,N_11935,N_11313);
nand U12654 (N_12654,N_11767,N_11934);
and U12655 (N_12655,N_11930,N_11745);
nor U12656 (N_12656,N_11708,N_11557);
nand U12657 (N_12657,N_11938,N_11832);
nand U12658 (N_12658,N_11220,N_11995);
nand U12659 (N_12659,N_11909,N_11275);
or U12660 (N_12660,N_11207,N_11541);
or U12661 (N_12661,N_11367,N_11946);
and U12662 (N_12662,N_11749,N_11406);
or U12663 (N_12663,N_11433,N_11350);
or U12664 (N_12664,N_11449,N_11276);
or U12665 (N_12665,N_11570,N_11346);
nor U12666 (N_12666,N_11541,N_11951);
nor U12667 (N_12667,N_11805,N_11822);
or U12668 (N_12668,N_11688,N_11318);
nor U12669 (N_12669,N_11297,N_11636);
and U12670 (N_12670,N_11780,N_11366);
or U12671 (N_12671,N_11590,N_11857);
nor U12672 (N_12672,N_11697,N_11643);
or U12673 (N_12673,N_11774,N_11854);
and U12674 (N_12674,N_11348,N_11546);
nand U12675 (N_12675,N_11726,N_11971);
or U12676 (N_12676,N_11930,N_11419);
nand U12677 (N_12677,N_11768,N_11350);
nor U12678 (N_12678,N_11811,N_11246);
nor U12679 (N_12679,N_11536,N_11475);
and U12680 (N_12680,N_11593,N_11397);
nor U12681 (N_12681,N_11884,N_11378);
nand U12682 (N_12682,N_11576,N_11965);
nand U12683 (N_12683,N_11604,N_11401);
nor U12684 (N_12684,N_11620,N_11510);
nor U12685 (N_12685,N_11397,N_11797);
or U12686 (N_12686,N_11453,N_11841);
nand U12687 (N_12687,N_11369,N_11667);
and U12688 (N_12688,N_11935,N_11293);
and U12689 (N_12689,N_11920,N_11622);
nand U12690 (N_12690,N_11327,N_11829);
nor U12691 (N_12691,N_11812,N_11804);
nand U12692 (N_12692,N_11674,N_11445);
and U12693 (N_12693,N_11629,N_11445);
nand U12694 (N_12694,N_11978,N_11449);
nor U12695 (N_12695,N_11465,N_11829);
nand U12696 (N_12696,N_11842,N_11998);
and U12697 (N_12697,N_11930,N_11670);
nor U12698 (N_12698,N_11380,N_11371);
and U12699 (N_12699,N_11872,N_11716);
and U12700 (N_12700,N_11604,N_11292);
and U12701 (N_12701,N_11588,N_11366);
nand U12702 (N_12702,N_11734,N_11538);
or U12703 (N_12703,N_11859,N_11835);
xnor U12704 (N_12704,N_11776,N_11604);
or U12705 (N_12705,N_11489,N_11774);
nor U12706 (N_12706,N_11407,N_11553);
or U12707 (N_12707,N_11855,N_11474);
and U12708 (N_12708,N_11440,N_11515);
nor U12709 (N_12709,N_11309,N_11454);
nor U12710 (N_12710,N_11385,N_11416);
or U12711 (N_12711,N_11559,N_11627);
nor U12712 (N_12712,N_11757,N_11210);
or U12713 (N_12713,N_11200,N_11221);
nor U12714 (N_12714,N_11821,N_11880);
and U12715 (N_12715,N_11802,N_11245);
or U12716 (N_12716,N_11469,N_11289);
nor U12717 (N_12717,N_11243,N_11600);
or U12718 (N_12718,N_11758,N_11628);
and U12719 (N_12719,N_11254,N_11395);
nand U12720 (N_12720,N_11713,N_11537);
nor U12721 (N_12721,N_11969,N_11484);
nor U12722 (N_12722,N_11910,N_11377);
and U12723 (N_12723,N_11753,N_11681);
nor U12724 (N_12724,N_11898,N_11580);
nand U12725 (N_12725,N_11853,N_11474);
nand U12726 (N_12726,N_11964,N_11987);
or U12727 (N_12727,N_11585,N_11459);
nand U12728 (N_12728,N_11406,N_11403);
and U12729 (N_12729,N_11514,N_11774);
nand U12730 (N_12730,N_11269,N_11319);
or U12731 (N_12731,N_11928,N_11368);
nand U12732 (N_12732,N_11770,N_11377);
or U12733 (N_12733,N_11679,N_11764);
and U12734 (N_12734,N_11723,N_11788);
or U12735 (N_12735,N_11307,N_11321);
or U12736 (N_12736,N_11922,N_11390);
or U12737 (N_12737,N_11480,N_11789);
or U12738 (N_12738,N_11664,N_11563);
and U12739 (N_12739,N_11214,N_11848);
or U12740 (N_12740,N_11785,N_11710);
nand U12741 (N_12741,N_11320,N_11467);
nor U12742 (N_12742,N_11803,N_11602);
nand U12743 (N_12743,N_11326,N_11661);
and U12744 (N_12744,N_11939,N_11469);
nand U12745 (N_12745,N_11754,N_11693);
and U12746 (N_12746,N_11745,N_11945);
nor U12747 (N_12747,N_11631,N_11390);
and U12748 (N_12748,N_11334,N_11472);
nor U12749 (N_12749,N_11796,N_11235);
nand U12750 (N_12750,N_11442,N_11503);
nor U12751 (N_12751,N_11664,N_11221);
xnor U12752 (N_12752,N_11436,N_11740);
or U12753 (N_12753,N_11659,N_11769);
and U12754 (N_12754,N_11897,N_11474);
nand U12755 (N_12755,N_11956,N_11785);
and U12756 (N_12756,N_11513,N_11278);
nand U12757 (N_12757,N_11584,N_11646);
nand U12758 (N_12758,N_11843,N_11959);
or U12759 (N_12759,N_11593,N_11940);
and U12760 (N_12760,N_11943,N_11395);
and U12761 (N_12761,N_11440,N_11340);
or U12762 (N_12762,N_11991,N_11470);
nor U12763 (N_12763,N_11358,N_11616);
and U12764 (N_12764,N_11224,N_11403);
nor U12765 (N_12765,N_11249,N_11587);
and U12766 (N_12766,N_11396,N_11572);
nor U12767 (N_12767,N_11570,N_11684);
or U12768 (N_12768,N_11865,N_11241);
or U12769 (N_12769,N_11657,N_11236);
nor U12770 (N_12770,N_11885,N_11481);
nand U12771 (N_12771,N_11854,N_11643);
or U12772 (N_12772,N_11324,N_11249);
nand U12773 (N_12773,N_11285,N_11845);
or U12774 (N_12774,N_11380,N_11881);
or U12775 (N_12775,N_11766,N_11494);
nand U12776 (N_12776,N_11241,N_11456);
nor U12777 (N_12777,N_11362,N_11569);
nor U12778 (N_12778,N_11579,N_11540);
nand U12779 (N_12779,N_11927,N_11967);
or U12780 (N_12780,N_11908,N_11822);
xor U12781 (N_12781,N_11895,N_11887);
nor U12782 (N_12782,N_11918,N_11520);
or U12783 (N_12783,N_11421,N_11522);
and U12784 (N_12784,N_11418,N_11785);
nor U12785 (N_12785,N_11951,N_11844);
nand U12786 (N_12786,N_11631,N_11491);
and U12787 (N_12787,N_11736,N_11711);
nor U12788 (N_12788,N_11955,N_11312);
and U12789 (N_12789,N_11969,N_11745);
or U12790 (N_12790,N_11750,N_11214);
nor U12791 (N_12791,N_11866,N_11864);
or U12792 (N_12792,N_11234,N_11551);
nand U12793 (N_12793,N_11704,N_11809);
and U12794 (N_12794,N_11842,N_11564);
or U12795 (N_12795,N_11305,N_11587);
or U12796 (N_12796,N_11426,N_11914);
nor U12797 (N_12797,N_11819,N_11922);
nand U12798 (N_12798,N_11866,N_11915);
or U12799 (N_12799,N_11210,N_11922);
nor U12800 (N_12800,N_12197,N_12083);
nand U12801 (N_12801,N_12268,N_12235);
nand U12802 (N_12802,N_12708,N_12711);
and U12803 (N_12803,N_12211,N_12581);
nor U12804 (N_12804,N_12342,N_12443);
or U12805 (N_12805,N_12042,N_12469);
nand U12806 (N_12806,N_12769,N_12272);
and U12807 (N_12807,N_12509,N_12670);
nand U12808 (N_12808,N_12321,N_12075);
or U12809 (N_12809,N_12672,N_12363);
and U12810 (N_12810,N_12775,N_12455);
nor U12811 (N_12811,N_12101,N_12104);
and U12812 (N_12812,N_12088,N_12512);
nor U12813 (N_12813,N_12229,N_12753);
or U12814 (N_12814,N_12430,N_12442);
nand U12815 (N_12815,N_12242,N_12511);
nor U12816 (N_12816,N_12464,N_12515);
or U12817 (N_12817,N_12137,N_12221);
nand U12818 (N_12818,N_12749,N_12326);
nand U12819 (N_12819,N_12517,N_12444);
and U12820 (N_12820,N_12699,N_12159);
or U12821 (N_12821,N_12752,N_12562);
and U12822 (N_12822,N_12791,N_12662);
or U12823 (N_12823,N_12693,N_12480);
nor U12824 (N_12824,N_12608,N_12356);
and U12825 (N_12825,N_12317,N_12239);
nor U12826 (N_12826,N_12015,N_12592);
nand U12827 (N_12827,N_12647,N_12679);
nor U12828 (N_12828,N_12723,N_12384);
or U12829 (N_12829,N_12357,N_12583);
nor U12830 (N_12830,N_12489,N_12566);
or U12831 (N_12831,N_12387,N_12352);
nand U12832 (N_12832,N_12278,N_12161);
and U12833 (N_12833,N_12270,N_12709);
nor U12834 (N_12834,N_12358,N_12234);
and U12835 (N_12835,N_12308,N_12668);
nand U12836 (N_12836,N_12786,N_12702);
nor U12837 (N_12837,N_12284,N_12025);
and U12838 (N_12838,N_12605,N_12418);
and U12839 (N_12839,N_12790,N_12386);
and U12840 (N_12840,N_12434,N_12655);
nand U12841 (N_12841,N_12334,N_12466);
or U12842 (N_12842,N_12764,N_12189);
and U12843 (N_12843,N_12733,N_12425);
and U12844 (N_12844,N_12779,N_12119);
nor U12845 (N_12845,N_12617,N_12461);
and U12846 (N_12846,N_12126,N_12459);
nor U12847 (N_12847,N_12000,N_12666);
or U12848 (N_12848,N_12732,N_12404);
and U12849 (N_12849,N_12663,N_12660);
and U12850 (N_12850,N_12479,N_12378);
and U12851 (N_12851,N_12661,N_12540);
or U12852 (N_12852,N_12586,N_12493);
nand U12853 (N_12853,N_12241,N_12324);
or U12854 (N_12854,N_12615,N_12701);
and U12855 (N_12855,N_12522,N_12628);
nor U12856 (N_12856,N_12422,N_12105);
nor U12857 (N_12857,N_12194,N_12738);
nand U12858 (N_12858,N_12001,N_12499);
or U12859 (N_12859,N_12123,N_12223);
and U12860 (N_12860,N_12618,N_12591);
nor U12861 (N_12861,N_12669,N_12501);
or U12862 (N_12862,N_12040,N_12406);
and U12863 (N_12863,N_12488,N_12081);
nand U12864 (N_12864,N_12058,N_12680);
nor U12865 (N_12865,N_12755,N_12012);
nand U12866 (N_12866,N_12758,N_12788);
nand U12867 (N_12867,N_12068,N_12539);
nor U12868 (N_12868,N_12286,N_12623);
or U12869 (N_12869,N_12022,N_12392);
nand U12870 (N_12870,N_12307,N_12237);
nand U12871 (N_12871,N_12649,N_12742);
nand U12872 (N_12872,N_12627,N_12041);
nor U12873 (N_12873,N_12465,N_12259);
and U12874 (N_12874,N_12759,N_12207);
and U12875 (N_12875,N_12298,N_12637);
nand U12876 (N_12876,N_12247,N_12062);
or U12877 (N_12877,N_12158,N_12181);
nand U12878 (N_12878,N_12588,N_12500);
and U12879 (N_12879,N_12431,N_12141);
nor U12880 (N_12880,N_12118,N_12044);
or U12881 (N_12881,N_12034,N_12651);
and U12882 (N_12882,N_12129,N_12082);
and U12883 (N_12883,N_12671,N_12110);
nand U12884 (N_12884,N_12593,N_12257);
nor U12885 (N_12885,N_12557,N_12027);
and U12886 (N_12886,N_12565,N_12178);
nor U12887 (N_12887,N_12611,N_12139);
nor U12888 (N_12888,N_12458,N_12125);
and U12889 (N_12889,N_12604,N_12339);
or U12890 (N_12890,N_12589,N_12633);
nor U12891 (N_12891,N_12282,N_12658);
and U12892 (N_12892,N_12408,N_12302);
or U12893 (N_12893,N_12399,N_12361);
nand U12894 (N_12894,N_12198,N_12559);
and U12895 (N_12895,N_12255,N_12398);
nor U12896 (N_12896,N_12403,N_12228);
or U12897 (N_12897,N_12251,N_12024);
nor U12898 (N_12898,N_12736,N_12787);
and U12899 (N_12899,N_12173,N_12016);
or U12900 (N_12900,N_12560,N_12706);
or U12901 (N_12901,N_12319,N_12396);
nor U12902 (N_12902,N_12536,N_12724);
and U12903 (N_12903,N_12776,N_12799);
or U12904 (N_12904,N_12745,N_12164);
nand U12905 (N_12905,N_12681,N_12697);
and U12906 (N_12906,N_12312,N_12383);
nand U12907 (N_12907,N_12475,N_12478);
nand U12908 (N_12908,N_12071,N_12541);
nand U12909 (N_12909,N_12160,N_12544);
and U12910 (N_12910,N_12320,N_12574);
nor U12911 (N_12911,N_12549,N_12543);
nor U12912 (N_12912,N_12518,N_12714);
and U12913 (N_12913,N_12630,N_12698);
nor U12914 (N_12914,N_12756,N_12219);
and U12915 (N_12915,N_12380,N_12254);
nor U12916 (N_12916,N_12009,N_12740);
nor U12917 (N_12917,N_12305,N_12086);
and U12918 (N_12918,N_12303,N_12166);
nor U12919 (N_12919,N_12797,N_12322);
or U12920 (N_12920,N_12638,N_12196);
or U12921 (N_12921,N_12631,N_12148);
nor U12922 (N_12922,N_12460,N_12610);
nand U12923 (N_12923,N_12453,N_12603);
and U12924 (N_12924,N_12297,N_12765);
or U12925 (N_12925,N_12664,N_12429);
or U12926 (N_12926,N_12098,N_12252);
and U12927 (N_12927,N_12503,N_12747);
nor U12928 (N_12928,N_12550,N_12450);
nand U12929 (N_12929,N_12304,N_12175);
nor U12930 (N_12930,N_12188,N_12644);
nor U12931 (N_12931,N_12057,N_12411);
and U12932 (N_12932,N_12463,N_12011);
nand U12933 (N_12933,N_12351,N_12064);
and U12934 (N_12934,N_12620,N_12705);
and U12935 (N_12935,N_12177,N_12066);
nor U12936 (N_12936,N_12156,N_12013);
nor U12937 (N_12937,N_12632,N_12224);
or U12938 (N_12938,N_12353,N_12438);
nor U12939 (N_12939,N_12032,N_12625);
nand U12940 (N_12940,N_12120,N_12529);
or U12941 (N_12941,N_12199,N_12147);
nor U12942 (N_12942,N_12486,N_12548);
or U12943 (N_12943,N_12523,N_12629);
nor U12944 (N_12944,N_12420,N_12341);
nor U12945 (N_12945,N_12067,N_12744);
nand U12946 (N_12946,N_12564,N_12760);
nand U12947 (N_12947,N_12505,N_12172);
xor U12948 (N_12948,N_12472,N_12323);
nand U12949 (N_12949,N_12456,N_12279);
nor U12950 (N_12950,N_12214,N_12613);
or U12951 (N_12951,N_12180,N_12263);
nand U12952 (N_12952,N_12401,N_12531);
and U12953 (N_12953,N_12296,N_12468);
and U12954 (N_12954,N_12416,N_12004);
nand U12955 (N_12955,N_12739,N_12439);
and U12956 (N_12956,N_12454,N_12641);
nor U12957 (N_12957,N_12191,N_12171);
nor U12958 (N_12958,N_12354,N_12691);
and U12959 (N_12959,N_12793,N_12155);
nand U12960 (N_12960,N_12579,N_12570);
nand U12961 (N_12961,N_12275,N_12049);
and U12962 (N_12962,N_12021,N_12682);
nor U12963 (N_12963,N_12367,N_12743);
nor U12964 (N_12964,N_12130,N_12785);
nand U12965 (N_12965,N_12528,N_12291);
and U12966 (N_12966,N_12375,N_12766);
nand U12967 (N_12967,N_12345,N_12093);
nand U12968 (N_12968,N_12726,N_12794);
and U12969 (N_12969,N_12530,N_12372);
nand U12970 (N_12970,N_12212,N_12645);
nor U12971 (N_12971,N_12400,N_12571);
and U12972 (N_12972,N_12169,N_12193);
nor U12973 (N_12973,N_12048,N_12133);
nand U12974 (N_12974,N_12731,N_12167);
or U12975 (N_12975,N_12216,N_12267);
nand U12976 (N_12976,N_12325,N_12763);
or U12977 (N_12977,N_12287,N_12673);
nand U12978 (N_12978,N_12773,N_12634);
and U12979 (N_12979,N_12572,N_12561);
and U12980 (N_12980,N_12165,N_12264);
nor U12981 (N_12981,N_12768,N_12294);
nor U12982 (N_12982,N_12762,N_12423);
or U12983 (N_12983,N_12084,N_12407);
or U12984 (N_12984,N_12721,N_12195);
nand U12985 (N_12985,N_12245,N_12151);
or U12986 (N_12986,N_12778,N_12598);
and U12987 (N_12987,N_12428,N_12240);
and U12988 (N_12988,N_12132,N_12421);
or U12989 (N_12989,N_12265,N_12606);
and U12990 (N_12990,N_12149,N_12507);
or U12991 (N_12991,N_12694,N_12782);
and U12992 (N_12992,N_12366,N_12446);
xnor U12993 (N_12993,N_12232,N_12185);
nor U12994 (N_12994,N_12692,N_12192);
nor U12995 (N_12995,N_12236,N_12654);
nand U12996 (N_12996,N_12121,N_12646);
nor U12997 (N_12997,N_12514,N_12359);
nand U12998 (N_12998,N_12371,N_12470);
nand U12999 (N_12999,N_12678,N_12784);
and U13000 (N_13000,N_12639,N_12316);
and U13001 (N_13001,N_12092,N_12152);
nand U13002 (N_13002,N_12487,N_12640);
nor U13003 (N_13003,N_12220,N_12700);
nand U13004 (N_13004,N_12017,N_12145);
nand U13005 (N_13005,N_12602,N_12094);
nand U13006 (N_13006,N_12447,N_12377);
nor U13007 (N_13007,N_12696,N_12533);
and U13008 (N_13008,N_12269,N_12204);
nand U13009 (N_13009,N_12520,N_12656);
and U13010 (N_13010,N_12767,N_12689);
and U13011 (N_13011,N_12715,N_12657);
or U13012 (N_13012,N_12619,N_12186);
and U13013 (N_13013,N_12626,N_12360);
and U13014 (N_13014,N_12491,N_12210);
nand U13015 (N_13015,N_12445,N_12055);
nand U13016 (N_13016,N_12770,N_12525);
or U13017 (N_13017,N_12532,N_12737);
nor U13018 (N_13018,N_12233,N_12329);
nor U13019 (N_13019,N_12607,N_12340);
or U13020 (N_13020,N_12652,N_12362);
nand U13021 (N_13021,N_12643,N_12440);
or U13022 (N_13022,N_12248,N_12496);
or U13023 (N_13023,N_12222,N_12558);
and U13024 (N_13024,N_12290,N_12409);
nand U13025 (N_13025,N_12402,N_12748);
or U13026 (N_13026,N_12449,N_12281);
or U13027 (N_13027,N_12348,N_12005);
nand U13028 (N_13028,N_12484,N_12215);
or U13029 (N_13029,N_12476,N_12047);
nand U13030 (N_13030,N_12551,N_12033);
nor U13031 (N_13031,N_12609,N_12018);
or U13032 (N_13032,N_12650,N_12538);
and U13033 (N_13033,N_12154,N_12474);
nor U13034 (N_13034,N_12096,N_12332);
and U13035 (N_13035,N_12718,N_12039);
nand U13036 (N_13036,N_12246,N_12136);
and U13037 (N_13037,N_12575,N_12006);
nor U13038 (N_13038,N_12335,N_12299);
nor U13039 (N_13039,N_12107,N_12771);
xor U13040 (N_13040,N_12261,N_12381);
or U13041 (N_13041,N_12382,N_12684);
or U13042 (N_13042,N_12163,N_12338);
or U13043 (N_13043,N_12410,N_12028);
nor U13044 (N_13044,N_12677,N_12053);
and U13045 (N_13045,N_12050,N_12546);
nand U13046 (N_13046,N_12276,N_12783);
or U13047 (N_13047,N_12208,N_12170);
and U13048 (N_13048,N_12614,N_12201);
nand U13049 (N_13049,N_12508,N_12757);
or U13050 (N_13050,N_12457,N_12433);
and U13051 (N_13051,N_12412,N_12209);
nand U13052 (N_13052,N_12318,N_12131);
nor U13053 (N_13053,N_12035,N_12330);
and U13054 (N_13054,N_12687,N_12648);
and U13055 (N_13055,N_12238,N_12087);
nand U13056 (N_13056,N_12369,N_12725);
nor U13057 (N_13057,N_12249,N_12060);
nor U13058 (N_13058,N_12002,N_12676);
nor U13059 (N_13059,N_12056,N_12492);
nand U13060 (N_13060,N_12043,N_12502);
nor U13061 (N_13061,N_12590,N_12576);
nand U13062 (N_13062,N_12622,N_12621);
and U13063 (N_13063,N_12497,N_12616);
and U13064 (N_13064,N_12280,N_12485);
or U13065 (N_13065,N_12054,N_12124);
or U13066 (N_13066,N_12010,N_12095);
nand U13067 (N_13067,N_12097,N_12331);
nor U13068 (N_13068,N_12162,N_12707);
nand U13069 (N_13069,N_12309,N_12003);
or U13070 (N_13070,N_12059,N_12206);
nand U13071 (N_13071,N_12665,N_12019);
or U13072 (N_13072,N_12350,N_12168);
or U13073 (N_13073,N_12713,N_12079);
and U13074 (N_13074,N_12601,N_12070);
nor U13075 (N_13075,N_12688,N_12435);
or U13076 (N_13076,N_12274,N_12547);
or U13077 (N_13077,N_12498,N_12537);
nand U13078 (N_13078,N_12419,N_12683);
and U13079 (N_13079,N_12080,N_12596);
and U13080 (N_13080,N_12138,N_12150);
nand U13081 (N_13081,N_12355,N_12065);
nor U13082 (N_13082,N_12253,N_12052);
and U13083 (N_13083,N_12277,N_12471);
nand U13084 (N_13084,N_12300,N_12527);
nand U13085 (N_13085,N_12008,N_12462);
or U13086 (N_13086,N_12481,N_12792);
and U13087 (N_13087,N_12504,N_12516);
and U13088 (N_13088,N_12580,N_12182);
nor U13089 (N_13089,N_12311,N_12552);
nor U13090 (N_13090,N_12127,N_12072);
and U13091 (N_13091,N_12063,N_12573);
nand U13092 (N_13092,N_12183,N_12395);
nand U13093 (N_13093,N_12069,N_12031);
or U13094 (N_13094,N_12102,N_12751);
nand U13095 (N_13095,N_12202,N_12283);
nor U13096 (N_13096,N_12686,N_12437);
nor U13097 (N_13097,N_12327,N_12336);
nand U13098 (N_13098,N_12675,N_12143);
or U13099 (N_13099,N_12730,N_12563);
and U13100 (N_13100,N_12370,N_12521);
and U13101 (N_13101,N_12077,N_12624);
and U13102 (N_13102,N_12385,N_12256);
or U13103 (N_13103,N_12347,N_12535);
or U13104 (N_13104,N_12142,N_12100);
and U13105 (N_13105,N_12146,N_12111);
or U13106 (N_13106,N_12599,N_12467);
nand U13107 (N_13107,N_12494,N_12727);
and U13108 (N_13108,N_12781,N_12519);
nand U13109 (N_13109,N_12122,N_12260);
nand U13110 (N_13110,N_12720,N_12789);
nor U13111 (N_13111,N_12587,N_12436);
or U13112 (N_13112,N_12293,N_12754);
or U13113 (N_13113,N_12685,N_12289);
and U13114 (N_13114,N_12427,N_12441);
nor U13115 (N_13115,N_12337,N_12513);
nor U13116 (N_13116,N_12258,N_12078);
nand U13117 (N_13117,N_12200,N_12405);
or U13118 (N_13118,N_12116,N_12365);
xnor U13119 (N_13119,N_12712,N_12734);
or U13120 (N_13120,N_12584,N_12424);
or U13121 (N_13121,N_12076,N_12719);
nand U13122 (N_13122,N_12038,N_12451);
nor U13123 (N_13123,N_12556,N_12091);
and U13124 (N_13124,N_12750,N_12314);
xnor U13125 (N_13125,N_12577,N_12482);
and U13126 (N_13126,N_12328,N_12271);
or U13127 (N_13127,N_12205,N_12448);
nand U13128 (N_13128,N_12397,N_12642);
nand U13129 (N_13129,N_12176,N_12452);
and U13130 (N_13130,N_12099,N_12379);
or U13131 (N_13131,N_12542,N_12495);
nand U13132 (N_13132,N_12554,N_12426);
or U13133 (N_13133,N_12594,N_12716);
and U13134 (N_13134,N_12343,N_12746);
and U13135 (N_13135,N_12761,N_12288);
or U13136 (N_13136,N_12295,N_12568);
and U13137 (N_13137,N_12413,N_12157);
nand U13138 (N_13138,N_12243,N_12089);
nand U13139 (N_13139,N_12373,N_12226);
or U13140 (N_13140,N_12510,N_12710);
or U13141 (N_13141,N_12029,N_12569);
and U13142 (N_13142,N_12273,N_12140);
and U13143 (N_13143,N_12073,N_12777);
nand U13144 (N_13144,N_12128,N_12106);
nand U13145 (N_13145,N_12112,N_12780);
and U13146 (N_13146,N_12704,N_12477);
or U13147 (N_13147,N_12153,N_12225);
and U13148 (N_13148,N_12795,N_12026);
nor U13149 (N_13149,N_12250,N_12483);
xor U13150 (N_13150,N_12595,N_12600);
and U13151 (N_13151,N_12717,N_12774);
nand U13152 (N_13152,N_12115,N_12203);
nor U13153 (N_13153,N_12389,N_12285);
nor U13154 (N_13154,N_12364,N_12635);
or U13155 (N_13155,N_12313,N_12374);
nand U13156 (N_13156,N_12187,N_12703);
nand U13157 (N_13157,N_12114,N_12722);
and U13158 (N_13158,N_12653,N_12230);
and U13159 (N_13159,N_12585,N_12578);
or U13160 (N_13160,N_12023,N_12037);
or U13161 (N_13161,N_12414,N_12090);
or U13162 (N_13162,N_12526,N_12134);
nand U13163 (N_13163,N_12695,N_12393);
and U13164 (N_13164,N_12582,N_12555);
or U13165 (N_13165,N_12333,N_12227);
nand U13166 (N_13166,N_12014,N_12074);
and U13167 (N_13167,N_12674,N_12534);
nor U13168 (N_13168,N_12553,N_12190);
and U13169 (N_13169,N_12415,N_12113);
nor U13170 (N_13170,N_12741,N_12612);
nor U13171 (N_13171,N_12796,N_12368);
nand U13172 (N_13172,N_12597,N_12390);
or U13173 (N_13173,N_12545,N_12524);
and U13174 (N_13174,N_12117,N_12490);
nor U13175 (N_13175,N_12030,N_12184);
and U13176 (N_13176,N_12346,N_12391);
nor U13177 (N_13177,N_12292,N_12798);
nor U13178 (N_13178,N_12262,N_12667);
and U13179 (N_13179,N_12244,N_12306);
and U13180 (N_13180,N_12007,N_12144);
nand U13181 (N_13181,N_12728,N_12301);
or U13182 (N_13182,N_12109,N_12217);
or U13183 (N_13183,N_12266,N_12659);
or U13184 (N_13184,N_12729,N_12473);
nand U13185 (N_13185,N_12394,N_12310);
and U13186 (N_13186,N_12690,N_12085);
nand U13187 (N_13187,N_12772,N_12045);
nand U13188 (N_13188,N_12432,N_12231);
or U13189 (N_13189,N_12506,N_12103);
and U13190 (N_13190,N_12179,N_12051);
nor U13191 (N_13191,N_12417,N_12020);
or U13192 (N_13192,N_12376,N_12135);
nor U13193 (N_13193,N_12636,N_12735);
or U13194 (N_13194,N_12567,N_12108);
nand U13195 (N_13195,N_12036,N_12213);
or U13196 (N_13196,N_12388,N_12174);
nand U13197 (N_13197,N_12349,N_12315);
nor U13198 (N_13198,N_12061,N_12344);
and U13199 (N_13199,N_12218,N_12046);
or U13200 (N_13200,N_12396,N_12259);
nor U13201 (N_13201,N_12081,N_12772);
nand U13202 (N_13202,N_12015,N_12173);
nand U13203 (N_13203,N_12164,N_12727);
or U13204 (N_13204,N_12493,N_12744);
or U13205 (N_13205,N_12433,N_12265);
or U13206 (N_13206,N_12614,N_12792);
nand U13207 (N_13207,N_12696,N_12265);
nor U13208 (N_13208,N_12110,N_12448);
and U13209 (N_13209,N_12289,N_12096);
and U13210 (N_13210,N_12365,N_12051);
or U13211 (N_13211,N_12708,N_12783);
and U13212 (N_13212,N_12502,N_12562);
nand U13213 (N_13213,N_12647,N_12694);
or U13214 (N_13214,N_12215,N_12581);
nor U13215 (N_13215,N_12264,N_12071);
or U13216 (N_13216,N_12724,N_12089);
nor U13217 (N_13217,N_12777,N_12719);
xnor U13218 (N_13218,N_12624,N_12643);
and U13219 (N_13219,N_12365,N_12248);
nor U13220 (N_13220,N_12658,N_12026);
and U13221 (N_13221,N_12699,N_12262);
nor U13222 (N_13222,N_12743,N_12486);
and U13223 (N_13223,N_12015,N_12416);
nand U13224 (N_13224,N_12640,N_12774);
and U13225 (N_13225,N_12756,N_12013);
nor U13226 (N_13226,N_12222,N_12263);
nand U13227 (N_13227,N_12365,N_12221);
and U13228 (N_13228,N_12320,N_12541);
nor U13229 (N_13229,N_12204,N_12038);
or U13230 (N_13230,N_12658,N_12258);
nor U13231 (N_13231,N_12285,N_12414);
nand U13232 (N_13232,N_12108,N_12427);
or U13233 (N_13233,N_12081,N_12034);
nand U13234 (N_13234,N_12484,N_12475);
or U13235 (N_13235,N_12497,N_12718);
nand U13236 (N_13236,N_12431,N_12559);
nand U13237 (N_13237,N_12593,N_12403);
nand U13238 (N_13238,N_12252,N_12776);
or U13239 (N_13239,N_12391,N_12550);
nor U13240 (N_13240,N_12796,N_12111);
nand U13241 (N_13241,N_12667,N_12544);
or U13242 (N_13242,N_12599,N_12277);
nor U13243 (N_13243,N_12005,N_12477);
nor U13244 (N_13244,N_12555,N_12651);
nand U13245 (N_13245,N_12631,N_12413);
nand U13246 (N_13246,N_12303,N_12144);
and U13247 (N_13247,N_12628,N_12604);
nand U13248 (N_13248,N_12617,N_12479);
nand U13249 (N_13249,N_12181,N_12682);
or U13250 (N_13250,N_12146,N_12119);
and U13251 (N_13251,N_12169,N_12037);
nand U13252 (N_13252,N_12450,N_12405);
nor U13253 (N_13253,N_12383,N_12227);
nand U13254 (N_13254,N_12494,N_12206);
nand U13255 (N_13255,N_12132,N_12426);
nand U13256 (N_13256,N_12158,N_12052);
nand U13257 (N_13257,N_12791,N_12575);
nor U13258 (N_13258,N_12618,N_12029);
or U13259 (N_13259,N_12333,N_12549);
nor U13260 (N_13260,N_12220,N_12023);
nor U13261 (N_13261,N_12596,N_12533);
and U13262 (N_13262,N_12542,N_12742);
and U13263 (N_13263,N_12603,N_12797);
and U13264 (N_13264,N_12189,N_12577);
nor U13265 (N_13265,N_12114,N_12431);
nand U13266 (N_13266,N_12798,N_12675);
and U13267 (N_13267,N_12689,N_12543);
or U13268 (N_13268,N_12501,N_12046);
nor U13269 (N_13269,N_12484,N_12180);
nor U13270 (N_13270,N_12686,N_12243);
nor U13271 (N_13271,N_12679,N_12772);
and U13272 (N_13272,N_12558,N_12157);
and U13273 (N_13273,N_12301,N_12713);
nand U13274 (N_13274,N_12025,N_12019);
and U13275 (N_13275,N_12562,N_12618);
xnor U13276 (N_13276,N_12739,N_12703);
nand U13277 (N_13277,N_12469,N_12765);
and U13278 (N_13278,N_12668,N_12033);
or U13279 (N_13279,N_12414,N_12653);
or U13280 (N_13280,N_12559,N_12565);
or U13281 (N_13281,N_12311,N_12326);
and U13282 (N_13282,N_12600,N_12596);
or U13283 (N_13283,N_12458,N_12469);
and U13284 (N_13284,N_12363,N_12000);
or U13285 (N_13285,N_12555,N_12427);
nand U13286 (N_13286,N_12212,N_12201);
and U13287 (N_13287,N_12035,N_12296);
nor U13288 (N_13288,N_12019,N_12539);
and U13289 (N_13289,N_12515,N_12458);
or U13290 (N_13290,N_12047,N_12448);
nor U13291 (N_13291,N_12686,N_12598);
and U13292 (N_13292,N_12139,N_12462);
nor U13293 (N_13293,N_12766,N_12465);
and U13294 (N_13294,N_12042,N_12354);
nand U13295 (N_13295,N_12059,N_12691);
and U13296 (N_13296,N_12208,N_12710);
or U13297 (N_13297,N_12187,N_12624);
or U13298 (N_13298,N_12353,N_12338);
or U13299 (N_13299,N_12767,N_12633);
nand U13300 (N_13300,N_12043,N_12328);
nand U13301 (N_13301,N_12195,N_12312);
nand U13302 (N_13302,N_12158,N_12647);
nand U13303 (N_13303,N_12774,N_12682);
and U13304 (N_13304,N_12462,N_12742);
and U13305 (N_13305,N_12234,N_12454);
or U13306 (N_13306,N_12212,N_12256);
nand U13307 (N_13307,N_12440,N_12414);
or U13308 (N_13308,N_12329,N_12038);
nor U13309 (N_13309,N_12430,N_12086);
and U13310 (N_13310,N_12712,N_12207);
and U13311 (N_13311,N_12468,N_12533);
or U13312 (N_13312,N_12213,N_12061);
nor U13313 (N_13313,N_12619,N_12327);
or U13314 (N_13314,N_12102,N_12137);
nand U13315 (N_13315,N_12761,N_12577);
nand U13316 (N_13316,N_12731,N_12448);
and U13317 (N_13317,N_12503,N_12735);
or U13318 (N_13318,N_12377,N_12779);
and U13319 (N_13319,N_12138,N_12377);
or U13320 (N_13320,N_12222,N_12737);
nand U13321 (N_13321,N_12562,N_12521);
or U13322 (N_13322,N_12341,N_12086);
and U13323 (N_13323,N_12694,N_12605);
or U13324 (N_13324,N_12283,N_12127);
nor U13325 (N_13325,N_12119,N_12037);
nand U13326 (N_13326,N_12230,N_12539);
nor U13327 (N_13327,N_12406,N_12445);
nor U13328 (N_13328,N_12425,N_12373);
nand U13329 (N_13329,N_12501,N_12056);
or U13330 (N_13330,N_12427,N_12731);
nand U13331 (N_13331,N_12381,N_12524);
nor U13332 (N_13332,N_12486,N_12061);
nor U13333 (N_13333,N_12002,N_12467);
nor U13334 (N_13334,N_12402,N_12064);
nor U13335 (N_13335,N_12370,N_12438);
and U13336 (N_13336,N_12633,N_12522);
nand U13337 (N_13337,N_12626,N_12359);
nor U13338 (N_13338,N_12513,N_12558);
or U13339 (N_13339,N_12614,N_12353);
or U13340 (N_13340,N_12236,N_12322);
nor U13341 (N_13341,N_12619,N_12407);
nor U13342 (N_13342,N_12184,N_12363);
nor U13343 (N_13343,N_12780,N_12573);
nor U13344 (N_13344,N_12647,N_12783);
and U13345 (N_13345,N_12090,N_12769);
nand U13346 (N_13346,N_12748,N_12300);
and U13347 (N_13347,N_12485,N_12071);
or U13348 (N_13348,N_12112,N_12068);
or U13349 (N_13349,N_12040,N_12431);
nand U13350 (N_13350,N_12510,N_12413);
nand U13351 (N_13351,N_12555,N_12654);
and U13352 (N_13352,N_12239,N_12664);
and U13353 (N_13353,N_12302,N_12568);
nor U13354 (N_13354,N_12583,N_12759);
and U13355 (N_13355,N_12545,N_12627);
or U13356 (N_13356,N_12541,N_12740);
nand U13357 (N_13357,N_12061,N_12681);
or U13358 (N_13358,N_12426,N_12545);
and U13359 (N_13359,N_12182,N_12622);
nor U13360 (N_13360,N_12362,N_12635);
nor U13361 (N_13361,N_12154,N_12463);
nand U13362 (N_13362,N_12324,N_12261);
and U13363 (N_13363,N_12136,N_12310);
and U13364 (N_13364,N_12719,N_12773);
or U13365 (N_13365,N_12234,N_12495);
nor U13366 (N_13366,N_12403,N_12234);
nor U13367 (N_13367,N_12441,N_12277);
or U13368 (N_13368,N_12037,N_12721);
nor U13369 (N_13369,N_12411,N_12033);
nand U13370 (N_13370,N_12013,N_12346);
nor U13371 (N_13371,N_12548,N_12238);
nor U13372 (N_13372,N_12029,N_12785);
nor U13373 (N_13373,N_12679,N_12525);
and U13374 (N_13374,N_12796,N_12692);
and U13375 (N_13375,N_12744,N_12753);
or U13376 (N_13376,N_12707,N_12204);
and U13377 (N_13377,N_12380,N_12409);
or U13378 (N_13378,N_12039,N_12633);
nor U13379 (N_13379,N_12271,N_12245);
and U13380 (N_13380,N_12097,N_12684);
nor U13381 (N_13381,N_12264,N_12713);
nand U13382 (N_13382,N_12637,N_12473);
or U13383 (N_13383,N_12548,N_12154);
nand U13384 (N_13384,N_12107,N_12531);
and U13385 (N_13385,N_12333,N_12533);
nand U13386 (N_13386,N_12152,N_12381);
nor U13387 (N_13387,N_12229,N_12746);
nor U13388 (N_13388,N_12265,N_12236);
nor U13389 (N_13389,N_12571,N_12133);
nor U13390 (N_13390,N_12448,N_12759);
nor U13391 (N_13391,N_12194,N_12783);
nor U13392 (N_13392,N_12500,N_12695);
and U13393 (N_13393,N_12792,N_12757);
and U13394 (N_13394,N_12127,N_12517);
and U13395 (N_13395,N_12354,N_12054);
nor U13396 (N_13396,N_12345,N_12194);
nand U13397 (N_13397,N_12345,N_12491);
nor U13398 (N_13398,N_12113,N_12326);
and U13399 (N_13399,N_12679,N_12004);
xor U13400 (N_13400,N_12760,N_12407);
nand U13401 (N_13401,N_12482,N_12747);
or U13402 (N_13402,N_12231,N_12277);
xnor U13403 (N_13403,N_12172,N_12073);
or U13404 (N_13404,N_12635,N_12773);
xor U13405 (N_13405,N_12117,N_12743);
or U13406 (N_13406,N_12620,N_12617);
nand U13407 (N_13407,N_12032,N_12505);
nor U13408 (N_13408,N_12320,N_12235);
nand U13409 (N_13409,N_12059,N_12581);
nand U13410 (N_13410,N_12743,N_12792);
nor U13411 (N_13411,N_12563,N_12545);
nor U13412 (N_13412,N_12651,N_12209);
or U13413 (N_13413,N_12456,N_12284);
or U13414 (N_13414,N_12238,N_12286);
and U13415 (N_13415,N_12164,N_12189);
or U13416 (N_13416,N_12141,N_12168);
nand U13417 (N_13417,N_12658,N_12368);
xor U13418 (N_13418,N_12594,N_12232);
nor U13419 (N_13419,N_12771,N_12529);
nand U13420 (N_13420,N_12762,N_12732);
nor U13421 (N_13421,N_12198,N_12346);
nor U13422 (N_13422,N_12583,N_12247);
or U13423 (N_13423,N_12692,N_12408);
nand U13424 (N_13424,N_12540,N_12673);
nand U13425 (N_13425,N_12241,N_12480);
and U13426 (N_13426,N_12654,N_12452);
nand U13427 (N_13427,N_12648,N_12030);
nor U13428 (N_13428,N_12416,N_12332);
nand U13429 (N_13429,N_12568,N_12107);
or U13430 (N_13430,N_12370,N_12356);
nand U13431 (N_13431,N_12709,N_12737);
nor U13432 (N_13432,N_12764,N_12237);
and U13433 (N_13433,N_12776,N_12350);
and U13434 (N_13434,N_12039,N_12536);
nor U13435 (N_13435,N_12242,N_12090);
nand U13436 (N_13436,N_12405,N_12372);
nor U13437 (N_13437,N_12473,N_12538);
nand U13438 (N_13438,N_12454,N_12154);
or U13439 (N_13439,N_12000,N_12144);
and U13440 (N_13440,N_12745,N_12540);
nand U13441 (N_13441,N_12190,N_12548);
nor U13442 (N_13442,N_12707,N_12717);
and U13443 (N_13443,N_12294,N_12193);
nor U13444 (N_13444,N_12543,N_12028);
and U13445 (N_13445,N_12102,N_12591);
or U13446 (N_13446,N_12098,N_12531);
and U13447 (N_13447,N_12227,N_12073);
nand U13448 (N_13448,N_12222,N_12231);
or U13449 (N_13449,N_12210,N_12377);
or U13450 (N_13450,N_12190,N_12793);
or U13451 (N_13451,N_12165,N_12466);
nor U13452 (N_13452,N_12633,N_12025);
nand U13453 (N_13453,N_12761,N_12424);
or U13454 (N_13454,N_12289,N_12733);
nand U13455 (N_13455,N_12096,N_12505);
and U13456 (N_13456,N_12300,N_12205);
or U13457 (N_13457,N_12292,N_12118);
or U13458 (N_13458,N_12350,N_12492);
or U13459 (N_13459,N_12552,N_12773);
and U13460 (N_13460,N_12463,N_12160);
nand U13461 (N_13461,N_12747,N_12682);
nor U13462 (N_13462,N_12097,N_12738);
and U13463 (N_13463,N_12239,N_12793);
nor U13464 (N_13464,N_12209,N_12641);
xor U13465 (N_13465,N_12010,N_12316);
nor U13466 (N_13466,N_12312,N_12660);
or U13467 (N_13467,N_12472,N_12713);
or U13468 (N_13468,N_12640,N_12410);
and U13469 (N_13469,N_12603,N_12026);
nor U13470 (N_13470,N_12603,N_12211);
nand U13471 (N_13471,N_12343,N_12190);
and U13472 (N_13472,N_12459,N_12726);
nand U13473 (N_13473,N_12166,N_12544);
or U13474 (N_13474,N_12395,N_12216);
or U13475 (N_13475,N_12762,N_12568);
nor U13476 (N_13476,N_12562,N_12685);
nor U13477 (N_13477,N_12748,N_12237);
nor U13478 (N_13478,N_12789,N_12561);
and U13479 (N_13479,N_12040,N_12383);
nand U13480 (N_13480,N_12354,N_12637);
nand U13481 (N_13481,N_12514,N_12190);
and U13482 (N_13482,N_12798,N_12120);
nand U13483 (N_13483,N_12400,N_12650);
or U13484 (N_13484,N_12065,N_12729);
nor U13485 (N_13485,N_12560,N_12558);
or U13486 (N_13486,N_12026,N_12696);
nand U13487 (N_13487,N_12144,N_12027);
nor U13488 (N_13488,N_12739,N_12635);
or U13489 (N_13489,N_12354,N_12034);
and U13490 (N_13490,N_12460,N_12324);
nor U13491 (N_13491,N_12277,N_12355);
nand U13492 (N_13492,N_12239,N_12395);
nand U13493 (N_13493,N_12361,N_12024);
or U13494 (N_13494,N_12725,N_12337);
and U13495 (N_13495,N_12662,N_12130);
nor U13496 (N_13496,N_12729,N_12580);
nand U13497 (N_13497,N_12096,N_12756);
nand U13498 (N_13498,N_12155,N_12049);
nor U13499 (N_13499,N_12344,N_12177);
or U13500 (N_13500,N_12555,N_12202);
and U13501 (N_13501,N_12282,N_12436);
nand U13502 (N_13502,N_12734,N_12203);
nor U13503 (N_13503,N_12538,N_12178);
or U13504 (N_13504,N_12589,N_12544);
nor U13505 (N_13505,N_12300,N_12371);
or U13506 (N_13506,N_12764,N_12262);
nand U13507 (N_13507,N_12607,N_12618);
nand U13508 (N_13508,N_12528,N_12193);
and U13509 (N_13509,N_12717,N_12337);
nor U13510 (N_13510,N_12718,N_12480);
nor U13511 (N_13511,N_12061,N_12657);
nand U13512 (N_13512,N_12492,N_12145);
nor U13513 (N_13513,N_12337,N_12735);
nand U13514 (N_13514,N_12036,N_12673);
nor U13515 (N_13515,N_12107,N_12795);
or U13516 (N_13516,N_12663,N_12341);
or U13517 (N_13517,N_12181,N_12559);
nor U13518 (N_13518,N_12449,N_12257);
and U13519 (N_13519,N_12541,N_12035);
nor U13520 (N_13520,N_12476,N_12760);
nor U13521 (N_13521,N_12314,N_12389);
nor U13522 (N_13522,N_12036,N_12789);
and U13523 (N_13523,N_12290,N_12522);
and U13524 (N_13524,N_12425,N_12792);
or U13525 (N_13525,N_12141,N_12774);
or U13526 (N_13526,N_12438,N_12721);
or U13527 (N_13527,N_12338,N_12753);
and U13528 (N_13528,N_12391,N_12459);
or U13529 (N_13529,N_12113,N_12465);
and U13530 (N_13530,N_12458,N_12606);
nor U13531 (N_13531,N_12005,N_12131);
nor U13532 (N_13532,N_12739,N_12456);
xor U13533 (N_13533,N_12306,N_12694);
and U13534 (N_13534,N_12106,N_12694);
or U13535 (N_13535,N_12660,N_12647);
nand U13536 (N_13536,N_12492,N_12518);
nand U13537 (N_13537,N_12623,N_12554);
or U13538 (N_13538,N_12195,N_12065);
nand U13539 (N_13539,N_12045,N_12359);
nand U13540 (N_13540,N_12716,N_12080);
or U13541 (N_13541,N_12542,N_12069);
nand U13542 (N_13542,N_12084,N_12424);
and U13543 (N_13543,N_12151,N_12001);
or U13544 (N_13544,N_12717,N_12228);
or U13545 (N_13545,N_12483,N_12074);
nand U13546 (N_13546,N_12063,N_12230);
and U13547 (N_13547,N_12133,N_12614);
nand U13548 (N_13548,N_12275,N_12641);
and U13549 (N_13549,N_12721,N_12394);
or U13550 (N_13550,N_12506,N_12623);
or U13551 (N_13551,N_12215,N_12118);
nand U13552 (N_13552,N_12067,N_12698);
or U13553 (N_13553,N_12000,N_12081);
and U13554 (N_13554,N_12084,N_12536);
xor U13555 (N_13555,N_12725,N_12794);
or U13556 (N_13556,N_12470,N_12746);
nor U13557 (N_13557,N_12193,N_12013);
or U13558 (N_13558,N_12508,N_12474);
or U13559 (N_13559,N_12068,N_12598);
or U13560 (N_13560,N_12187,N_12116);
nor U13561 (N_13561,N_12455,N_12432);
and U13562 (N_13562,N_12404,N_12543);
nand U13563 (N_13563,N_12505,N_12371);
and U13564 (N_13564,N_12626,N_12488);
and U13565 (N_13565,N_12477,N_12071);
nand U13566 (N_13566,N_12269,N_12678);
and U13567 (N_13567,N_12088,N_12463);
and U13568 (N_13568,N_12144,N_12308);
and U13569 (N_13569,N_12150,N_12285);
nand U13570 (N_13570,N_12222,N_12134);
nand U13571 (N_13571,N_12624,N_12524);
nand U13572 (N_13572,N_12375,N_12417);
and U13573 (N_13573,N_12668,N_12407);
or U13574 (N_13574,N_12443,N_12617);
nand U13575 (N_13575,N_12454,N_12507);
or U13576 (N_13576,N_12283,N_12493);
or U13577 (N_13577,N_12245,N_12111);
and U13578 (N_13578,N_12436,N_12640);
and U13579 (N_13579,N_12156,N_12000);
or U13580 (N_13580,N_12518,N_12356);
nand U13581 (N_13581,N_12039,N_12180);
and U13582 (N_13582,N_12269,N_12572);
nand U13583 (N_13583,N_12486,N_12608);
nand U13584 (N_13584,N_12517,N_12286);
and U13585 (N_13585,N_12010,N_12221);
nand U13586 (N_13586,N_12069,N_12318);
or U13587 (N_13587,N_12386,N_12008);
nand U13588 (N_13588,N_12349,N_12763);
nor U13589 (N_13589,N_12757,N_12277);
or U13590 (N_13590,N_12313,N_12785);
and U13591 (N_13591,N_12138,N_12163);
or U13592 (N_13592,N_12789,N_12386);
and U13593 (N_13593,N_12359,N_12380);
and U13594 (N_13594,N_12099,N_12308);
nor U13595 (N_13595,N_12122,N_12346);
nor U13596 (N_13596,N_12048,N_12714);
nand U13597 (N_13597,N_12112,N_12093);
nand U13598 (N_13598,N_12629,N_12626);
nand U13599 (N_13599,N_12799,N_12135);
nor U13600 (N_13600,N_13469,N_12832);
nor U13601 (N_13601,N_12906,N_13039);
or U13602 (N_13602,N_13449,N_13382);
xor U13603 (N_13603,N_12817,N_12897);
nand U13604 (N_13604,N_13306,N_12875);
and U13605 (N_13605,N_13145,N_13074);
or U13606 (N_13606,N_13002,N_13336);
and U13607 (N_13607,N_13439,N_12911);
and U13608 (N_13608,N_13094,N_13089);
nand U13609 (N_13609,N_12929,N_12956);
or U13610 (N_13610,N_13305,N_13506);
nor U13611 (N_13611,N_12950,N_13071);
or U13612 (N_13612,N_13377,N_13205);
nor U13613 (N_13613,N_13058,N_13433);
and U13614 (N_13614,N_13418,N_13076);
or U13615 (N_13615,N_13151,N_13133);
or U13616 (N_13616,N_13226,N_13582);
nor U13617 (N_13617,N_13011,N_13533);
nor U13618 (N_13618,N_13148,N_12974);
and U13619 (N_13619,N_13276,N_13060);
and U13620 (N_13620,N_12936,N_13153);
nand U13621 (N_13621,N_13102,N_13188);
nor U13622 (N_13622,N_13190,N_13373);
nor U13623 (N_13623,N_13405,N_13375);
and U13624 (N_13624,N_13480,N_13477);
and U13625 (N_13625,N_13195,N_13494);
nand U13626 (N_13626,N_13444,N_13157);
nor U13627 (N_13627,N_12989,N_12846);
nand U13628 (N_13628,N_12914,N_13108);
or U13629 (N_13629,N_13220,N_12941);
nor U13630 (N_13630,N_12899,N_12807);
and U13631 (N_13631,N_13465,N_13257);
and U13632 (N_13632,N_13374,N_13558);
or U13633 (N_13633,N_13458,N_13202);
nand U13634 (N_13634,N_13097,N_13595);
nor U13635 (N_13635,N_13378,N_13163);
nand U13636 (N_13636,N_12963,N_12959);
or U13637 (N_13637,N_12841,N_13473);
nand U13638 (N_13638,N_12852,N_13292);
and U13639 (N_13639,N_12858,N_13553);
or U13640 (N_13640,N_13347,N_13580);
and U13641 (N_13641,N_13491,N_13571);
or U13642 (N_13642,N_13046,N_13550);
nor U13643 (N_13643,N_13057,N_12812);
nand U13644 (N_13644,N_13345,N_13495);
nand U13645 (N_13645,N_13036,N_12982);
nand U13646 (N_13646,N_12973,N_13112);
nor U13647 (N_13647,N_13001,N_12831);
and U13648 (N_13648,N_13185,N_13173);
nor U13649 (N_13649,N_13370,N_12979);
and U13650 (N_13650,N_13169,N_13243);
nand U13651 (N_13651,N_12993,N_13399);
nor U13652 (N_13652,N_13517,N_13474);
or U13653 (N_13653,N_12946,N_13056);
nor U13654 (N_13654,N_12928,N_13197);
nand U13655 (N_13655,N_13274,N_12940);
and U13656 (N_13656,N_13519,N_13260);
nand U13657 (N_13657,N_13155,N_13263);
and U13658 (N_13658,N_13103,N_12879);
and U13659 (N_13659,N_13514,N_13597);
nor U13660 (N_13660,N_13438,N_13249);
or U13661 (N_13661,N_13028,N_12876);
and U13662 (N_13662,N_13338,N_13177);
nand U13663 (N_13663,N_13532,N_13122);
nor U13664 (N_13664,N_13525,N_12919);
nand U13665 (N_13665,N_13037,N_13181);
or U13666 (N_13666,N_12826,N_13326);
or U13667 (N_13667,N_13222,N_13049);
nand U13668 (N_13668,N_13352,N_13124);
nand U13669 (N_13669,N_13587,N_13068);
or U13670 (N_13670,N_13584,N_13107);
and U13671 (N_13671,N_13271,N_13518);
or U13672 (N_13672,N_12964,N_13476);
or U13673 (N_13673,N_13441,N_13266);
nor U13674 (N_13674,N_12883,N_13383);
nor U13675 (N_13675,N_13238,N_13515);
and U13676 (N_13676,N_12996,N_13052);
or U13677 (N_13677,N_13023,N_12834);
and U13678 (N_13678,N_13388,N_13219);
nor U13679 (N_13679,N_13556,N_13273);
nor U13680 (N_13680,N_13093,N_12909);
or U13681 (N_13681,N_12872,N_13363);
and U13682 (N_13682,N_13174,N_13579);
or U13683 (N_13683,N_13530,N_13161);
nand U13684 (N_13684,N_12965,N_13420);
nor U13685 (N_13685,N_13411,N_13229);
nand U13686 (N_13686,N_13047,N_12819);
nor U13687 (N_13687,N_13258,N_12983);
nor U13688 (N_13688,N_13406,N_12984);
or U13689 (N_13689,N_13078,N_13077);
nor U13690 (N_13690,N_13537,N_12967);
and U13691 (N_13691,N_13470,N_12844);
and U13692 (N_13692,N_13536,N_13212);
nand U13693 (N_13693,N_13261,N_13455);
or U13694 (N_13694,N_12981,N_13315);
nor U13695 (N_13695,N_13164,N_13072);
nor U13696 (N_13696,N_13282,N_13129);
nand U13697 (N_13697,N_13483,N_13593);
xor U13698 (N_13698,N_13127,N_12925);
and U13699 (N_13699,N_13138,N_12930);
nor U13700 (N_13700,N_13291,N_13310);
and U13701 (N_13701,N_12961,N_13198);
or U13702 (N_13702,N_12887,N_13030);
and U13703 (N_13703,N_12994,N_13193);
nor U13704 (N_13704,N_13268,N_13064);
or U13705 (N_13705,N_13371,N_13069);
nor U13706 (N_13706,N_12801,N_13095);
nand U13707 (N_13707,N_13296,N_13423);
or U13708 (N_13708,N_13445,N_13490);
nand U13709 (N_13709,N_13385,N_13351);
and U13710 (N_13710,N_13572,N_13568);
nor U13711 (N_13711,N_12836,N_13355);
or U13712 (N_13712,N_12847,N_12820);
or U13713 (N_13713,N_13115,N_13005);
nand U13714 (N_13714,N_13502,N_13029);
and U13715 (N_13715,N_13430,N_12856);
nand U13716 (N_13716,N_13573,N_13019);
and U13717 (N_13717,N_13534,N_13557);
nand U13718 (N_13718,N_13496,N_13548);
nand U13719 (N_13719,N_12802,N_13365);
xor U13720 (N_13720,N_12874,N_13114);
or U13721 (N_13721,N_12860,N_13403);
or U13722 (N_13722,N_13464,N_12823);
nor U13723 (N_13723,N_12999,N_13589);
or U13724 (N_13724,N_13009,N_13234);
nand U13725 (N_13725,N_13309,N_13203);
nand U13726 (N_13726,N_13538,N_13179);
nor U13727 (N_13727,N_12962,N_13516);
or U13728 (N_13728,N_12885,N_12977);
nand U13729 (N_13729,N_13436,N_13443);
nand U13730 (N_13730,N_13435,N_13528);
nand U13731 (N_13731,N_13280,N_12873);
or U13732 (N_13732,N_13492,N_12896);
nand U13733 (N_13733,N_13225,N_12995);
nor U13734 (N_13734,N_13098,N_13171);
and U13735 (N_13735,N_13182,N_13394);
nand U13736 (N_13736,N_12842,N_13594);
and U13737 (N_13737,N_13105,N_12953);
and U13738 (N_13738,N_12815,N_13462);
or U13739 (N_13739,N_13442,N_13467);
nand U13740 (N_13740,N_13279,N_13563);
or U13741 (N_13741,N_13017,N_13505);
and U13742 (N_13742,N_13520,N_13313);
and U13743 (N_13743,N_13307,N_13410);
or U13744 (N_13744,N_13531,N_13397);
nand U13745 (N_13745,N_13241,N_13487);
and U13746 (N_13746,N_13488,N_13246);
or U13747 (N_13747,N_13040,N_13081);
nand U13748 (N_13748,N_13523,N_13269);
and U13749 (N_13749,N_13484,N_13390);
nor U13750 (N_13750,N_12969,N_12934);
nand U13751 (N_13751,N_13468,N_13143);
or U13752 (N_13752,N_13192,N_13301);
nor U13753 (N_13753,N_13343,N_13598);
nand U13754 (N_13754,N_13284,N_12881);
or U13755 (N_13755,N_13239,N_13547);
or U13756 (N_13756,N_13250,N_13569);
nand U13757 (N_13757,N_13475,N_13543);
or U13758 (N_13758,N_13456,N_13278);
nand U13759 (N_13759,N_13391,N_13059);
or U13760 (N_13760,N_13576,N_12990);
nor U13761 (N_13761,N_12866,N_12884);
nor U13762 (N_13762,N_13025,N_12833);
and U13763 (N_13763,N_12827,N_13293);
and U13764 (N_13764,N_12809,N_13228);
nor U13765 (N_13765,N_13581,N_12918);
and U13766 (N_13766,N_13327,N_12870);
nand U13767 (N_13767,N_13311,N_13508);
nand U13768 (N_13768,N_13073,N_12931);
and U13769 (N_13769,N_12900,N_13044);
nand U13770 (N_13770,N_13522,N_13366);
nand U13771 (N_13771,N_13575,N_13004);
and U13772 (N_13772,N_12935,N_13413);
and U13773 (N_13773,N_13409,N_13350);
nand U13774 (N_13774,N_13223,N_13554);
nor U13775 (N_13775,N_13245,N_12835);
nor U13776 (N_13776,N_12895,N_13006);
nor U13777 (N_13777,N_12840,N_13312);
and U13778 (N_13778,N_13051,N_12912);
or U13779 (N_13779,N_13175,N_13207);
nand U13780 (N_13780,N_13578,N_13450);
and U13781 (N_13781,N_12943,N_12904);
or U13782 (N_13782,N_12971,N_13401);
and U13783 (N_13783,N_13404,N_12988);
nor U13784 (N_13784,N_13369,N_13559);
nand U13785 (N_13785,N_13116,N_13135);
nor U13786 (N_13786,N_12976,N_13204);
or U13787 (N_13787,N_13299,N_12932);
or U13788 (N_13788,N_13552,N_13574);
or U13789 (N_13789,N_13147,N_13214);
and U13790 (N_13790,N_13139,N_13591);
nand U13791 (N_13791,N_13294,N_13539);
nor U13792 (N_13792,N_12814,N_13248);
and U13793 (N_13793,N_12893,N_13083);
and U13794 (N_13794,N_13217,N_13482);
nand U13795 (N_13795,N_13067,N_13199);
xor U13796 (N_13796,N_13170,N_13070);
nand U13797 (N_13797,N_12803,N_13564);
nand U13798 (N_13798,N_13026,N_13437);
or U13799 (N_13799,N_13149,N_13407);
or U13800 (N_13800,N_13334,N_13331);
and U13801 (N_13801,N_12838,N_13416);
or U13802 (N_13802,N_13168,N_13141);
nor U13803 (N_13803,N_13372,N_13144);
and U13804 (N_13804,N_12920,N_12938);
or U13805 (N_13805,N_12902,N_13429);
or U13806 (N_13806,N_12978,N_13131);
or U13807 (N_13807,N_13189,N_13440);
nand U13808 (N_13808,N_13463,N_13230);
and U13809 (N_13809,N_13165,N_13194);
or U13810 (N_13810,N_13562,N_13038);
and U13811 (N_13811,N_12987,N_13035);
and U13812 (N_13812,N_12947,N_12954);
and U13813 (N_13813,N_13275,N_13590);
nand U13814 (N_13814,N_13201,N_13288);
or U13815 (N_13815,N_13412,N_13592);
nor U13816 (N_13816,N_13356,N_13360);
or U13817 (N_13817,N_13446,N_13513);
nand U13818 (N_13818,N_13196,N_12980);
nor U13819 (N_13819,N_13459,N_12960);
or U13820 (N_13820,N_13050,N_12958);
xnor U13821 (N_13821,N_13066,N_13362);
or U13822 (N_13822,N_13478,N_13498);
nor U13823 (N_13823,N_13020,N_13493);
and U13824 (N_13824,N_12891,N_13330);
nand U13825 (N_13825,N_13027,N_13134);
or U13826 (N_13826,N_12921,N_12926);
and U13827 (N_13827,N_12949,N_12972);
nand U13828 (N_13828,N_13392,N_13111);
nor U13829 (N_13829,N_13048,N_13158);
and U13830 (N_13830,N_12944,N_13191);
and U13831 (N_13831,N_12937,N_13024);
and U13832 (N_13832,N_13320,N_13332);
nand U13833 (N_13833,N_12882,N_13585);
and U13834 (N_13834,N_13289,N_13256);
nand U13835 (N_13835,N_12966,N_13216);
nand U13836 (N_13836,N_13396,N_13504);
nor U13837 (N_13837,N_13252,N_12849);
and U13838 (N_13838,N_13361,N_13259);
nor U13839 (N_13839,N_13546,N_13113);
nand U13840 (N_13840,N_13460,N_12915);
and U13841 (N_13841,N_12818,N_12992);
or U13842 (N_13842,N_13422,N_13224);
nand U13843 (N_13843,N_13100,N_12888);
nor U13844 (N_13844,N_13032,N_12865);
or U13845 (N_13845,N_13298,N_13099);
or U13846 (N_13846,N_13453,N_13542);
or U13847 (N_13847,N_13221,N_13080);
and U13848 (N_13848,N_13079,N_13096);
nand U13849 (N_13849,N_13142,N_13346);
nand U13850 (N_13850,N_13128,N_12851);
nor U13851 (N_13851,N_12864,N_13088);
and U13852 (N_13852,N_13152,N_13267);
or U13853 (N_13853,N_12952,N_13075);
and U13854 (N_13854,N_12843,N_12892);
nor U13855 (N_13855,N_13120,N_13053);
nor U13856 (N_13856,N_13290,N_12828);
or U13857 (N_13857,N_13324,N_13596);
or U13858 (N_13858,N_12862,N_13337);
and U13859 (N_13859,N_13384,N_13014);
nor U13860 (N_13860,N_12901,N_12825);
xnor U13861 (N_13861,N_13018,N_13321);
nor U13862 (N_13862,N_12933,N_12800);
or U13863 (N_13863,N_13535,N_13570);
nand U13864 (N_13864,N_13130,N_13215);
or U13865 (N_13865,N_13526,N_13244);
and U13866 (N_13866,N_13090,N_13387);
or U13867 (N_13867,N_13354,N_12886);
or U13868 (N_13868,N_13395,N_13092);
and U13869 (N_13869,N_13031,N_13325);
nand U13870 (N_13870,N_13457,N_13187);
nand U13871 (N_13871,N_13417,N_13277);
nor U13872 (N_13872,N_13472,N_13156);
and U13873 (N_13873,N_13400,N_13063);
or U13874 (N_13874,N_13479,N_13357);
and U13875 (N_13875,N_13398,N_12877);
nand U13876 (N_13876,N_12871,N_13428);
nand U13877 (N_13877,N_12811,N_13297);
and U13878 (N_13878,N_12848,N_13551);
nor U13879 (N_13879,N_13447,N_12927);
nand U13880 (N_13880,N_13461,N_13527);
nand U13881 (N_13881,N_13389,N_13167);
or U13882 (N_13882,N_13233,N_12804);
or U13883 (N_13883,N_12822,N_12970);
nand U13884 (N_13884,N_13583,N_13184);
nand U13885 (N_13885,N_13426,N_12942);
nand U13886 (N_13886,N_13242,N_13489);
nand U13887 (N_13887,N_13335,N_13328);
nand U13888 (N_13888,N_13454,N_13264);
nor U13889 (N_13889,N_12821,N_13255);
or U13890 (N_13890,N_12986,N_12878);
and U13891 (N_13891,N_12913,N_13016);
nand U13892 (N_13892,N_13281,N_13588);
and U13893 (N_13893,N_13010,N_13555);
or U13894 (N_13894,N_13367,N_13507);
nor U13895 (N_13895,N_13414,N_13524);
nand U13896 (N_13896,N_13132,N_12998);
nor U13897 (N_13897,N_12985,N_13510);
nor U13898 (N_13898,N_13376,N_13062);
nor U13899 (N_13899,N_13265,N_12957);
or U13900 (N_13900,N_13379,N_13566);
or U13901 (N_13901,N_13211,N_13034);
nor U13902 (N_13902,N_13380,N_13349);
or U13903 (N_13903,N_13364,N_12910);
and U13904 (N_13904,N_13000,N_13237);
and U13905 (N_13905,N_12867,N_13486);
or U13906 (N_13906,N_12839,N_13159);
nand U13907 (N_13907,N_13393,N_13300);
nand U13908 (N_13908,N_13541,N_13186);
nand U13909 (N_13909,N_13432,N_13353);
and U13910 (N_13910,N_12855,N_13270);
nor U13911 (N_13911,N_13125,N_12924);
nor U13912 (N_13912,N_12908,N_13381);
or U13913 (N_13913,N_12863,N_13421);
nand U13914 (N_13914,N_12854,N_12951);
nor U13915 (N_13915,N_13304,N_13065);
and U13916 (N_13916,N_13323,N_13283);
and U13917 (N_13917,N_13082,N_13425);
or U13918 (N_13918,N_13340,N_13358);
nand U13919 (N_13919,N_12939,N_12948);
or U13920 (N_13920,N_13431,N_12917);
nor U13921 (N_13921,N_12880,N_13232);
and U13922 (N_13922,N_13545,N_13021);
nand U13923 (N_13923,N_12810,N_13121);
or U13924 (N_13924,N_13316,N_13287);
nor U13925 (N_13925,N_13015,N_13109);
nand U13926 (N_13926,N_13448,N_13150);
and U13927 (N_13927,N_13117,N_12903);
and U13928 (N_13928,N_13160,N_13424);
nand U13929 (N_13929,N_13471,N_12850);
nand U13930 (N_13930,N_13285,N_13511);
nand U13931 (N_13931,N_13303,N_12845);
or U13932 (N_13932,N_13013,N_13126);
nand U13933 (N_13933,N_13500,N_13368);
or U13934 (N_13934,N_13419,N_12853);
nor U13935 (N_13935,N_12806,N_13033);
or U13936 (N_13936,N_13162,N_13042);
or U13937 (N_13937,N_13586,N_13272);
nand U13938 (N_13938,N_13045,N_12894);
nor U13939 (N_13939,N_13227,N_12868);
nor U13940 (N_13940,N_12975,N_13118);
and U13941 (N_13941,N_13560,N_13521);
or U13942 (N_13942,N_12869,N_13434);
or U13943 (N_13943,N_13251,N_13344);
or U13944 (N_13944,N_13104,N_13087);
nor U13945 (N_13945,N_12955,N_13577);
nor U13946 (N_13946,N_13322,N_13061);
or U13947 (N_13947,N_12907,N_13084);
or U13948 (N_13948,N_13235,N_13086);
or U13949 (N_13949,N_12889,N_13180);
or U13950 (N_13950,N_13166,N_13339);
or U13951 (N_13951,N_13481,N_13561);
or U13952 (N_13952,N_13043,N_13286);
or U13953 (N_13953,N_13240,N_12824);
nand U13954 (N_13954,N_13497,N_12890);
nor U13955 (N_13955,N_13247,N_13236);
nor U13956 (N_13956,N_13302,N_13209);
or U13957 (N_13957,N_13402,N_13567);
and U13958 (N_13958,N_13106,N_13342);
or U13959 (N_13959,N_12968,N_13022);
nor U13960 (N_13960,N_13178,N_12923);
nor U13961 (N_13961,N_13308,N_13540);
nor U13962 (N_13962,N_13599,N_13253);
and U13963 (N_13963,N_13466,N_12916);
and U13964 (N_13964,N_13254,N_12813);
and U13965 (N_13965,N_13172,N_13509);
or U13966 (N_13966,N_13110,N_13341);
or U13967 (N_13967,N_13154,N_13231);
and U13968 (N_13968,N_13208,N_13262);
or U13969 (N_13969,N_13295,N_13101);
or U13970 (N_13970,N_13136,N_13318);
nand U13971 (N_13971,N_13140,N_13427);
and U13972 (N_13972,N_13415,N_13512);
nand U13973 (N_13973,N_13012,N_12808);
or U13974 (N_13974,N_12857,N_12837);
nor U13975 (N_13975,N_13146,N_12830);
and U13976 (N_13976,N_13085,N_13054);
or U13977 (N_13977,N_13176,N_13544);
nand U13978 (N_13978,N_13359,N_12829);
nor U13979 (N_13979,N_12816,N_13210);
or U13980 (N_13980,N_13008,N_13206);
or U13981 (N_13981,N_13333,N_13529);
nand U13982 (N_13982,N_13319,N_13501);
nand U13983 (N_13983,N_13452,N_13329);
nor U13984 (N_13984,N_13317,N_13119);
and U13985 (N_13985,N_12861,N_13408);
nor U13986 (N_13986,N_13137,N_12922);
or U13987 (N_13987,N_13183,N_13451);
and U13988 (N_13988,N_13503,N_13200);
nand U13989 (N_13989,N_13003,N_13499);
or U13990 (N_13990,N_13348,N_12991);
nor U13991 (N_13991,N_12905,N_12805);
nand U13992 (N_13992,N_13055,N_13549);
nor U13993 (N_13993,N_13213,N_12997);
nor U13994 (N_13994,N_12859,N_12945);
nor U13995 (N_13995,N_13218,N_13041);
nor U13996 (N_13996,N_13123,N_13485);
and U13997 (N_13997,N_13091,N_13007);
nor U13998 (N_13998,N_13386,N_13565);
and U13999 (N_13999,N_12898,N_13314);
or U14000 (N_14000,N_13478,N_13097);
nor U14001 (N_14001,N_13165,N_13137);
and U14002 (N_14002,N_13402,N_12978);
nor U14003 (N_14003,N_12841,N_13126);
or U14004 (N_14004,N_13262,N_13079);
and U14005 (N_14005,N_13247,N_13252);
and U14006 (N_14006,N_13022,N_12813);
and U14007 (N_14007,N_13535,N_13418);
and U14008 (N_14008,N_12984,N_12891);
nor U14009 (N_14009,N_13438,N_13330);
nor U14010 (N_14010,N_13594,N_13511);
or U14011 (N_14011,N_13583,N_12904);
and U14012 (N_14012,N_13573,N_13174);
nand U14013 (N_14013,N_13457,N_13113);
nand U14014 (N_14014,N_13583,N_12996);
or U14015 (N_14015,N_13092,N_13188);
nor U14016 (N_14016,N_13120,N_13057);
nor U14017 (N_14017,N_13058,N_13049);
or U14018 (N_14018,N_13262,N_13401);
nand U14019 (N_14019,N_12823,N_13566);
nand U14020 (N_14020,N_13440,N_12944);
and U14021 (N_14021,N_13140,N_12867);
or U14022 (N_14022,N_13149,N_12882);
or U14023 (N_14023,N_13288,N_13318);
nand U14024 (N_14024,N_12802,N_13387);
or U14025 (N_14025,N_12801,N_12803);
and U14026 (N_14026,N_12904,N_13485);
or U14027 (N_14027,N_13078,N_12831);
and U14028 (N_14028,N_13091,N_13245);
nor U14029 (N_14029,N_13270,N_12972);
nand U14030 (N_14030,N_13164,N_13145);
and U14031 (N_14031,N_13395,N_12945);
nor U14032 (N_14032,N_13597,N_13078);
nor U14033 (N_14033,N_13385,N_13121);
nand U14034 (N_14034,N_13003,N_12836);
nand U14035 (N_14035,N_12976,N_13587);
nand U14036 (N_14036,N_13535,N_13556);
xor U14037 (N_14037,N_12931,N_13466);
or U14038 (N_14038,N_13078,N_13107);
nor U14039 (N_14039,N_12928,N_13482);
and U14040 (N_14040,N_13425,N_12944);
nor U14041 (N_14041,N_13523,N_13333);
or U14042 (N_14042,N_12859,N_12981);
or U14043 (N_14043,N_13193,N_13268);
or U14044 (N_14044,N_12805,N_13315);
or U14045 (N_14045,N_13305,N_13485);
nand U14046 (N_14046,N_13566,N_12815);
nand U14047 (N_14047,N_12859,N_13207);
nand U14048 (N_14048,N_12886,N_13236);
nor U14049 (N_14049,N_13143,N_13001);
nand U14050 (N_14050,N_12859,N_12964);
or U14051 (N_14051,N_13544,N_13430);
and U14052 (N_14052,N_12913,N_13219);
and U14053 (N_14053,N_13410,N_13278);
and U14054 (N_14054,N_12929,N_13122);
and U14055 (N_14055,N_12870,N_12983);
or U14056 (N_14056,N_13567,N_12810);
or U14057 (N_14057,N_13521,N_13299);
nor U14058 (N_14058,N_13523,N_12866);
nand U14059 (N_14059,N_12832,N_12948);
or U14060 (N_14060,N_13366,N_13426);
nor U14061 (N_14061,N_13494,N_13316);
nor U14062 (N_14062,N_12864,N_13124);
nand U14063 (N_14063,N_13088,N_13087);
nor U14064 (N_14064,N_13514,N_12969);
nand U14065 (N_14065,N_13596,N_13291);
nand U14066 (N_14066,N_12927,N_13372);
and U14067 (N_14067,N_12823,N_13234);
and U14068 (N_14068,N_12831,N_13296);
nor U14069 (N_14069,N_13230,N_13029);
nor U14070 (N_14070,N_12997,N_12898);
nand U14071 (N_14071,N_13243,N_13529);
nand U14072 (N_14072,N_12939,N_13593);
or U14073 (N_14073,N_12848,N_13089);
and U14074 (N_14074,N_13005,N_13323);
or U14075 (N_14075,N_13328,N_13543);
and U14076 (N_14076,N_12901,N_13457);
or U14077 (N_14077,N_13598,N_13134);
or U14078 (N_14078,N_13117,N_13293);
nand U14079 (N_14079,N_13123,N_13543);
xnor U14080 (N_14080,N_12891,N_13258);
nand U14081 (N_14081,N_13264,N_12941);
nand U14082 (N_14082,N_13324,N_13042);
nor U14083 (N_14083,N_13357,N_12906);
nor U14084 (N_14084,N_13114,N_13048);
nand U14085 (N_14085,N_12994,N_13261);
nand U14086 (N_14086,N_12937,N_12813);
nor U14087 (N_14087,N_13196,N_13261);
xnor U14088 (N_14088,N_13252,N_13138);
nand U14089 (N_14089,N_12853,N_13415);
and U14090 (N_14090,N_13386,N_13167);
nor U14091 (N_14091,N_12879,N_13523);
nor U14092 (N_14092,N_13257,N_12985);
nor U14093 (N_14093,N_13051,N_13198);
nor U14094 (N_14094,N_13557,N_13502);
and U14095 (N_14095,N_13235,N_13263);
nor U14096 (N_14096,N_13264,N_13115);
nand U14097 (N_14097,N_13255,N_12979);
nand U14098 (N_14098,N_13164,N_12870);
and U14099 (N_14099,N_13048,N_12925);
and U14100 (N_14100,N_12917,N_12934);
or U14101 (N_14101,N_12846,N_12844);
nor U14102 (N_14102,N_12866,N_13593);
nor U14103 (N_14103,N_12987,N_13193);
nor U14104 (N_14104,N_12939,N_13255);
and U14105 (N_14105,N_13189,N_12994);
and U14106 (N_14106,N_13052,N_13285);
and U14107 (N_14107,N_13066,N_13268);
and U14108 (N_14108,N_13178,N_13073);
and U14109 (N_14109,N_12959,N_12949);
and U14110 (N_14110,N_13290,N_13444);
or U14111 (N_14111,N_13470,N_13096);
or U14112 (N_14112,N_13273,N_13262);
nand U14113 (N_14113,N_13178,N_12952);
nor U14114 (N_14114,N_13233,N_13365);
nor U14115 (N_14115,N_13296,N_13384);
nand U14116 (N_14116,N_12974,N_12998);
nor U14117 (N_14117,N_13180,N_13554);
and U14118 (N_14118,N_13291,N_13124);
nor U14119 (N_14119,N_13410,N_12930);
nand U14120 (N_14120,N_13222,N_12985);
and U14121 (N_14121,N_13064,N_13366);
nor U14122 (N_14122,N_13201,N_13228);
nor U14123 (N_14123,N_12937,N_12896);
nand U14124 (N_14124,N_12975,N_13019);
and U14125 (N_14125,N_13177,N_13303);
or U14126 (N_14126,N_13289,N_12864);
nand U14127 (N_14127,N_13346,N_13306);
and U14128 (N_14128,N_13146,N_13260);
or U14129 (N_14129,N_13198,N_12866);
nor U14130 (N_14130,N_13364,N_13142);
or U14131 (N_14131,N_13125,N_13245);
nand U14132 (N_14132,N_13053,N_13086);
nand U14133 (N_14133,N_12965,N_13188);
and U14134 (N_14134,N_13289,N_13387);
nor U14135 (N_14135,N_13138,N_13106);
nand U14136 (N_14136,N_12957,N_13072);
nand U14137 (N_14137,N_13391,N_13592);
nor U14138 (N_14138,N_13057,N_12958);
and U14139 (N_14139,N_12909,N_12989);
and U14140 (N_14140,N_13285,N_13134);
nand U14141 (N_14141,N_13513,N_13305);
and U14142 (N_14142,N_13412,N_13032);
nand U14143 (N_14143,N_12937,N_13283);
nor U14144 (N_14144,N_13425,N_13420);
nand U14145 (N_14145,N_13540,N_13165);
nand U14146 (N_14146,N_13323,N_12864);
nand U14147 (N_14147,N_12948,N_13026);
and U14148 (N_14148,N_13086,N_12985);
or U14149 (N_14149,N_12965,N_13551);
or U14150 (N_14150,N_13138,N_13147);
and U14151 (N_14151,N_12944,N_12856);
or U14152 (N_14152,N_13428,N_13016);
and U14153 (N_14153,N_13408,N_13287);
xor U14154 (N_14154,N_13581,N_12994);
nor U14155 (N_14155,N_13390,N_13000);
nor U14156 (N_14156,N_13241,N_13544);
and U14157 (N_14157,N_12845,N_13116);
and U14158 (N_14158,N_13335,N_13222);
nor U14159 (N_14159,N_13454,N_13354);
nand U14160 (N_14160,N_13336,N_13165);
or U14161 (N_14161,N_13298,N_13310);
and U14162 (N_14162,N_13483,N_13232);
nand U14163 (N_14163,N_13101,N_13160);
nand U14164 (N_14164,N_13289,N_13160);
nor U14165 (N_14165,N_13138,N_13570);
nand U14166 (N_14166,N_13417,N_13093);
xor U14167 (N_14167,N_12952,N_12872);
or U14168 (N_14168,N_13438,N_13106);
and U14169 (N_14169,N_12984,N_13221);
nand U14170 (N_14170,N_13185,N_13480);
or U14171 (N_14171,N_13066,N_13312);
or U14172 (N_14172,N_13178,N_13261);
nand U14173 (N_14173,N_13089,N_13238);
nor U14174 (N_14174,N_13293,N_12812);
or U14175 (N_14175,N_13411,N_13439);
or U14176 (N_14176,N_12956,N_13068);
nor U14177 (N_14177,N_13476,N_13012);
nand U14178 (N_14178,N_13542,N_13551);
xnor U14179 (N_14179,N_13361,N_13025);
nor U14180 (N_14180,N_12867,N_13376);
and U14181 (N_14181,N_13434,N_13127);
or U14182 (N_14182,N_13021,N_13034);
nor U14183 (N_14183,N_13462,N_13123);
and U14184 (N_14184,N_13232,N_13159);
or U14185 (N_14185,N_13295,N_13034);
or U14186 (N_14186,N_12905,N_13385);
nor U14187 (N_14187,N_13526,N_13148);
and U14188 (N_14188,N_13498,N_13442);
nand U14189 (N_14189,N_12815,N_13056);
or U14190 (N_14190,N_13388,N_12992);
nand U14191 (N_14191,N_13283,N_12810);
or U14192 (N_14192,N_13019,N_13575);
nand U14193 (N_14193,N_12981,N_13155);
nand U14194 (N_14194,N_13061,N_13543);
nand U14195 (N_14195,N_13532,N_13129);
nor U14196 (N_14196,N_13324,N_12916);
nand U14197 (N_14197,N_13368,N_12931);
xnor U14198 (N_14198,N_13289,N_13227);
or U14199 (N_14199,N_12972,N_13262);
or U14200 (N_14200,N_13021,N_13184);
or U14201 (N_14201,N_13596,N_12851);
nand U14202 (N_14202,N_13112,N_12935);
or U14203 (N_14203,N_13184,N_13508);
and U14204 (N_14204,N_13417,N_13159);
nor U14205 (N_14205,N_12847,N_13323);
and U14206 (N_14206,N_13008,N_13436);
xor U14207 (N_14207,N_13275,N_13452);
nor U14208 (N_14208,N_13335,N_12843);
xor U14209 (N_14209,N_12962,N_12822);
and U14210 (N_14210,N_13540,N_13265);
and U14211 (N_14211,N_13554,N_13037);
nand U14212 (N_14212,N_12954,N_13046);
and U14213 (N_14213,N_13112,N_13137);
nand U14214 (N_14214,N_13054,N_13317);
and U14215 (N_14215,N_13284,N_13060);
nor U14216 (N_14216,N_13135,N_13305);
nand U14217 (N_14217,N_13113,N_13340);
nor U14218 (N_14218,N_13233,N_12918);
nand U14219 (N_14219,N_13385,N_12866);
or U14220 (N_14220,N_13486,N_13055);
nand U14221 (N_14221,N_12884,N_13350);
nand U14222 (N_14222,N_13287,N_13327);
and U14223 (N_14223,N_13551,N_12985);
nand U14224 (N_14224,N_13587,N_13306);
nand U14225 (N_14225,N_12965,N_13305);
and U14226 (N_14226,N_12832,N_13281);
nand U14227 (N_14227,N_13014,N_13586);
and U14228 (N_14228,N_12894,N_12818);
nand U14229 (N_14229,N_13039,N_12871);
or U14230 (N_14230,N_12925,N_12986);
and U14231 (N_14231,N_13205,N_12819);
nor U14232 (N_14232,N_13479,N_13534);
and U14233 (N_14233,N_12842,N_13461);
nor U14234 (N_14234,N_13250,N_12943);
nand U14235 (N_14235,N_13037,N_13166);
or U14236 (N_14236,N_13083,N_13263);
nand U14237 (N_14237,N_13514,N_13041);
and U14238 (N_14238,N_13593,N_12819);
nor U14239 (N_14239,N_13419,N_13202);
and U14240 (N_14240,N_13488,N_12825);
nor U14241 (N_14241,N_13128,N_13122);
nor U14242 (N_14242,N_13100,N_12990);
and U14243 (N_14243,N_12905,N_13254);
nor U14244 (N_14244,N_12844,N_13592);
nor U14245 (N_14245,N_13172,N_13169);
nor U14246 (N_14246,N_13471,N_13524);
nor U14247 (N_14247,N_12845,N_13202);
or U14248 (N_14248,N_13422,N_12986);
nand U14249 (N_14249,N_13523,N_12990);
nor U14250 (N_14250,N_13199,N_13393);
nor U14251 (N_14251,N_13089,N_13105);
and U14252 (N_14252,N_13570,N_13075);
xnor U14253 (N_14253,N_13299,N_13055);
nor U14254 (N_14254,N_13417,N_13342);
or U14255 (N_14255,N_12876,N_13358);
nand U14256 (N_14256,N_13213,N_13259);
nand U14257 (N_14257,N_12966,N_13380);
or U14258 (N_14258,N_13591,N_13396);
or U14259 (N_14259,N_13281,N_13001);
nand U14260 (N_14260,N_13450,N_13499);
nor U14261 (N_14261,N_13375,N_12806);
and U14262 (N_14262,N_13269,N_13068);
nor U14263 (N_14263,N_13094,N_13282);
nor U14264 (N_14264,N_13031,N_13265);
nor U14265 (N_14265,N_13408,N_12921);
nor U14266 (N_14266,N_13277,N_13251);
or U14267 (N_14267,N_12959,N_13278);
nand U14268 (N_14268,N_13221,N_13110);
nand U14269 (N_14269,N_13228,N_12898);
and U14270 (N_14270,N_13293,N_13322);
and U14271 (N_14271,N_13307,N_12908);
nand U14272 (N_14272,N_13480,N_13228);
nor U14273 (N_14273,N_13555,N_13497);
or U14274 (N_14274,N_13519,N_12812);
or U14275 (N_14275,N_12967,N_12973);
or U14276 (N_14276,N_13489,N_12896);
or U14277 (N_14277,N_12837,N_12976);
or U14278 (N_14278,N_12803,N_13445);
nor U14279 (N_14279,N_12834,N_12849);
nand U14280 (N_14280,N_12835,N_13422);
nand U14281 (N_14281,N_13012,N_13595);
nand U14282 (N_14282,N_13460,N_13186);
and U14283 (N_14283,N_13233,N_13167);
and U14284 (N_14284,N_13224,N_13443);
and U14285 (N_14285,N_13083,N_12959);
nor U14286 (N_14286,N_13417,N_12837);
nand U14287 (N_14287,N_13336,N_13061);
or U14288 (N_14288,N_13443,N_13266);
nor U14289 (N_14289,N_12899,N_13191);
or U14290 (N_14290,N_13444,N_13097);
nand U14291 (N_14291,N_13069,N_13210);
and U14292 (N_14292,N_12803,N_12996);
or U14293 (N_14293,N_13144,N_12958);
or U14294 (N_14294,N_12813,N_12878);
nand U14295 (N_14295,N_13350,N_12889);
nand U14296 (N_14296,N_13195,N_13315);
nand U14297 (N_14297,N_13457,N_13106);
nand U14298 (N_14298,N_13503,N_13309);
and U14299 (N_14299,N_13324,N_13171);
nor U14300 (N_14300,N_13139,N_12948);
nand U14301 (N_14301,N_12872,N_12926);
or U14302 (N_14302,N_13027,N_13227);
nor U14303 (N_14303,N_13523,N_13497);
nand U14304 (N_14304,N_13240,N_13100);
or U14305 (N_14305,N_13422,N_12819);
nor U14306 (N_14306,N_13119,N_13591);
and U14307 (N_14307,N_13018,N_12987);
nand U14308 (N_14308,N_13051,N_13177);
nand U14309 (N_14309,N_13384,N_13563);
nor U14310 (N_14310,N_13255,N_13578);
nor U14311 (N_14311,N_13067,N_13078);
nand U14312 (N_14312,N_13246,N_13467);
or U14313 (N_14313,N_13251,N_13555);
nor U14314 (N_14314,N_13179,N_12902);
nand U14315 (N_14315,N_13128,N_13426);
or U14316 (N_14316,N_12922,N_12938);
or U14317 (N_14317,N_13453,N_12877);
nand U14318 (N_14318,N_13229,N_13008);
nor U14319 (N_14319,N_13205,N_13416);
and U14320 (N_14320,N_13122,N_13392);
or U14321 (N_14321,N_12924,N_13158);
and U14322 (N_14322,N_13403,N_13501);
or U14323 (N_14323,N_13514,N_13237);
or U14324 (N_14324,N_13136,N_13393);
nor U14325 (N_14325,N_13158,N_13457);
and U14326 (N_14326,N_13201,N_13526);
and U14327 (N_14327,N_12803,N_12922);
and U14328 (N_14328,N_12985,N_13282);
or U14329 (N_14329,N_13557,N_12808);
nor U14330 (N_14330,N_12805,N_12910);
or U14331 (N_14331,N_12903,N_12891);
nor U14332 (N_14332,N_13048,N_13028);
or U14333 (N_14333,N_13477,N_13552);
or U14334 (N_14334,N_12890,N_13593);
or U14335 (N_14335,N_12933,N_12812);
or U14336 (N_14336,N_13422,N_13185);
nor U14337 (N_14337,N_13211,N_13586);
and U14338 (N_14338,N_13415,N_13232);
nor U14339 (N_14339,N_13529,N_13321);
nand U14340 (N_14340,N_13125,N_13167);
nand U14341 (N_14341,N_13358,N_12821);
nand U14342 (N_14342,N_13132,N_13210);
nor U14343 (N_14343,N_12909,N_12836);
nand U14344 (N_14344,N_13525,N_12916);
and U14345 (N_14345,N_12844,N_13093);
or U14346 (N_14346,N_13331,N_12827);
and U14347 (N_14347,N_13274,N_13013);
or U14348 (N_14348,N_13288,N_13084);
and U14349 (N_14349,N_13181,N_13395);
or U14350 (N_14350,N_13062,N_12901);
or U14351 (N_14351,N_12939,N_13416);
or U14352 (N_14352,N_13506,N_13308);
nand U14353 (N_14353,N_12963,N_12962);
nor U14354 (N_14354,N_13539,N_13153);
and U14355 (N_14355,N_13316,N_13363);
or U14356 (N_14356,N_12827,N_12996);
nand U14357 (N_14357,N_13293,N_13471);
nand U14358 (N_14358,N_13112,N_13298);
nand U14359 (N_14359,N_12993,N_12982);
or U14360 (N_14360,N_13225,N_13106);
xnor U14361 (N_14361,N_13042,N_13003);
or U14362 (N_14362,N_13124,N_13515);
and U14363 (N_14363,N_13148,N_12803);
or U14364 (N_14364,N_13446,N_12929);
or U14365 (N_14365,N_13309,N_12884);
or U14366 (N_14366,N_13585,N_13596);
and U14367 (N_14367,N_13300,N_13491);
and U14368 (N_14368,N_12823,N_13425);
nand U14369 (N_14369,N_13024,N_13246);
nand U14370 (N_14370,N_13096,N_12966);
nand U14371 (N_14371,N_12878,N_12882);
or U14372 (N_14372,N_12998,N_13285);
and U14373 (N_14373,N_13101,N_12854);
or U14374 (N_14374,N_12875,N_13066);
nor U14375 (N_14375,N_13318,N_13510);
and U14376 (N_14376,N_13025,N_13043);
nor U14377 (N_14377,N_12847,N_12946);
nand U14378 (N_14378,N_13276,N_13229);
nor U14379 (N_14379,N_13128,N_13190);
and U14380 (N_14380,N_13501,N_13572);
nand U14381 (N_14381,N_13359,N_12996);
nand U14382 (N_14382,N_13497,N_13598);
xor U14383 (N_14383,N_13396,N_12954);
nor U14384 (N_14384,N_12892,N_13536);
and U14385 (N_14385,N_13323,N_13231);
nand U14386 (N_14386,N_13065,N_13399);
nand U14387 (N_14387,N_13576,N_13361);
and U14388 (N_14388,N_12892,N_13503);
nor U14389 (N_14389,N_12835,N_13523);
and U14390 (N_14390,N_13423,N_13191);
nand U14391 (N_14391,N_13165,N_13546);
or U14392 (N_14392,N_13165,N_13400);
nand U14393 (N_14393,N_13255,N_13216);
nand U14394 (N_14394,N_13508,N_12860);
or U14395 (N_14395,N_13310,N_12918);
nand U14396 (N_14396,N_13283,N_13432);
nand U14397 (N_14397,N_13097,N_13324);
and U14398 (N_14398,N_13199,N_13410);
or U14399 (N_14399,N_13217,N_13211);
nand U14400 (N_14400,N_14325,N_13803);
and U14401 (N_14401,N_14027,N_14048);
or U14402 (N_14402,N_14378,N_14081);
or U14403 (N_14403,N_13649,N_14067);
nor U14404 (N_14404,N_14074,N_14220);
or U14405 (N_14405,N_14221,N_13915);
nor U14406 (N_14406,N_14046,N_13745);
and U14407 (N_14407,N_13815,N_13938);
and U14408 (N_14408,N_13642,N_14098);
or U14409 (N_14409,N_14391,N_14372);
nand U14410 (N_14410,N_13710,N_13684);
nor U14411 (N_14411,N_14056,N_14135);
nand U14412 (N_14412,N_14241,N_14269);
or U14413 (N_14413,N_13676,N_14266);
or U14414 (N_14414,N_13919,N_13601);
or U14415 (N_14415,N_14084,N_13709);
and U14416 (N_14416,N_14304,N_14394);
nand U14417 (N_14417,N_13814,N_14293);
or U14418 (N_14418,N_14340,N_14308);
or U14419 (N_14419,N_14077,N_13848);
and U14420 (N_14420,N_14109,N_14256);
or U14421 (N_14421,N_13858,N_14363);
or U14422 (N_14422,N_13847,N_14037);
nand U14423 (N_14423,N_14367,N_13944);
and U14424 (N_14424,N_14319,N_14019);
nor U14425 (N_14425,N_13740,N_13977);
and U14426 (N_14426,N_14263,N_14150);
or U14427 (N_14427,N_14085,N_13708);
nand U14428 (N_14428,N_14195,N_13764);
nor U14429 (N_14429,N_13648,N_13725);
and U14430 (N_14430,N_13687,N_14217);
and U14431 (N_14431,N_13742,N_13747);
or U14432 (N_14432,N_13974,N_13822);
and U14433 (N_14433,N_13975,N_14021);
nor U14434 (N_14434,N_13630,N_13972);
nand U14435 (N_14435,N_14318,N_14274);
and U14436 (N_14436,N_13653,N_14291);
or U14437 (N_14437,N_14247,N_14213);
and U14438 (N_14438,N_13806,N_13827);
or U14439 (N_14439,N_13800,N_13786);
or U14440 (N_14440,N_13668,N_13777);
nor U14441 (N_14441,N_14347,N_13624);
nor U14442 (N_14442,N_14159,N_14317);
and U14443 (N_14443,N_13783,N_14038);
nand U14444 (N_14444,N_14113,N_14285);
nand U14445 (N_14445,N_13970,N_14301);
nor U14446 (N_14446,N_14128,N_14232);
and U14447 (N_14447,N_13850,N_14359);
and U14448 (N_14448,N_14315,N_13669);
and U14449 (N_14449,N_13730,N_14013);
and U14450 (N_14450,N_13695,N_13646);
and U14451 (N_14451,N_14354,N_13962);
or U14452 (N_14452,N_14193,N_13785);
nand U14453 (N_14453,N_14160,N_13690);
nor U14454 (N_14454,N_14306,N_13634);
nor U14455 (N_14455,N_13771,N_14351);
or U14456 (N_14456,N_13600,N_13776);
nand U14457 (N_14457,N_14146,N_14239);
nor U14458 (N_14458,N_14370,N_14130);
nor U14459 (N_14459,N_14222,N_13888);
nor U14460 (N_14460,N_13914,N_14083);
nand U14461 (N_14461,N_13950,N_13656);
and U14462 (N_14462,N_13895,N_14395);
nor U14463 (N_14463,N_13818,N_13907);
nor U14464 (N_14464,N_13920,N_14052);
nand U14465 (N_14465,N_13635,N_13908);
or U14466 (N_14466,N_14396,N_13799);
nor U14467 (N_14467,N_14248,N_13942);
and U14468 (N_14468,N_13623,N_13791);
or U14469 (N_14469,N_14384,N_13704);
nor U14470 (N_14470,N_14070,N_14287);
and U14471 (N_14471,N_14258,N_13992);
nor U14472 (N_14472,N_13715,N_13660);
or U14473 (N_14473,N_13901,N_14211);
nand U14474 (N_14474,N_14186,N_14179);
nand U14475 (N_14475,N_14334,N_13645);
nor U14476 (N_14476,N_14259,N_14358);
and U14477 (N_14477,N_14024,N_13606);
or U14478 (N_14478,N_13863,N_13658);
or U14479 (N_14479,N_13963,N_13775);
nor U14480 (N_14480,N_14022,N_13774);
or U14481 (N_14481,N_14377,N_14339);
and U14482 (N_14482,N_13906,N_14235);
and U14483 (N_14483,N_14245,N_13654);
nor U14484 (N_14484,N_14071,N_13918);
nand U14485 (N_14485,N_14264,N_13767);
or U14486 (N_14486,N_14086,N_14393);
nand U14487 (N_14487,N_14194,N_14151);
nor U14488 (N_14488,N_13940,N_14397);
nand U14489 (N_14489,N_14092,N_14348);
and U14490 (N_14490,N_14234,N_13813);
nand U14491 (N_14491,N_13766,N_14107);
xnor U14492 (N_14492,N_13788,N_14337);
or U14493 (N_14493,N_13714,N_13861);
or U14494 (N_14494,N_13639,N_14373);
nor U14495 (N_14495,N_13770,N_13955);
nand U14496 (N_14496,N_14157,N_14224);
or U14497 (N_14497,N_13926,N_14023);
or U14498 (N_14498,N_13947,N_14271);
nand U14499 (N_14499,N_13867,N_13967);
or U14500 (N_14500,N_14129,N_13825);
nand U14501 (N_14501,N_14254,N_13820);
nand U14502 (N_14502,N_14229,N_13986);
or U14503 (N_14503,N_13757,N_14161);
or U14504 (N_14504,N_13719,N_13762);
nor U14505 (N_14505,N_14294,N_14177);
nand U14506 (N_14506,N_14163,N_14345);
nand U14507 (N_14507,N_13885,N_13670);
nor U14508 (N_14508,N_13697,N_13741);
and U14509 (N_14509,N_14366,N_14261);
nor U14510 (N_14510,N_14117,N_13664);
and U14511 (N_14511,N_13923,N_13989);
nand U14512 (N_14512,N_13969,N_14008);
nor U14513 (N_14513,N_13769,N_13994);
or U14514 (N_14514,N_14126,N_14143);
nand U14515 (N_14515,N_14356,N_13904);
or U14516 (N_14516,N_13807,N_14200);
and U14517 (N_14517,N_13722,N_14277);
and U14518 (N_14518,N_13675,N_14093);
and U14519 (N_14519,N_13717,N_14145);
or U14520 (N_14520,N_14360,N_13931);
or U14521 (N_14521,N_14243,N_14114);
nand U14522 (N_14522,N_14281,N_14167);
nor U14523 (N_14523,N_13765,N_13759);
or U14524 (N_14524,N_14132,N_14399);
and U14525 (N_14525,N_13968,N_14064);
nor U14526 (N_14526,N_14355,N_14004);
and U14527 (N_14527,N_13711,N_13781);
nand U14528 (N_14528,N_13935,N_14270);
or U14529 (N_14529,N_14025,N_13981);
and U14530 (N_14530,N_13737,N_14119);
nand U14531 (N_14531,N_14329,N_13958);
and U14532 (N_14532,N_13622,N_13726);
nand U14533 (N_14533,N_14171,N_13638);
and U14534 (N_14534,N_14326,N_14058);
nor U14535 (N_14535,N_14127,N_14267);
or U14536 (N_14536,N_13846,N_13749);
nor U14537 (N_14537,N_13988,N_14342);
nor U14538 (N_14538,N_14050,N_13841);
and U14539 (N_14539,N_13753,N_14047);
nor U14540 (N_14540,N_13934,N_13853);
or U14541 (N_14541,N_13641,N_13933);
or U14542 (N_14542,N_13971,N_14196);
or U14543 (N_14543,N_14230,N_14014);
and U14544 (N_14544,N_14244,N_13787);
nor U14545 (N_14545,N_14204,N_14072);
nor U14546 (N_14546,N_13666,N_13680);
or U14547 (N_14547,N_13812,N_14283);
and U14548 (N_14548,N_14189,N_13864);
and U14549 (N_14549,N_14231,N_14218);
or U14550 (N_14550,N_14296,N_13804);
or U14551 (N_14551,N_13712,N_14298);
nor U14552 (N_14552,N_13945,N_14011);
and U14553 (N_14553,N_13637,N_14180);
and U14554 (N_14554,N_14252,N_13921);
nand U14555 (N_14555,N_14103,N_13999);
nor U14556 (N_14556,N_13924,N_13862);
nor U14557 (N_14557,N_14152,N_14147);
and U14558 (N_14558,N_13796,N_13889);
or U14559 (N_14559,N_14295,N_13881);
nor U14560 (N_14560,N_13723,N_14102);
nor U14561 (N_14561,N_14068,N_13916);
nor U14562 (N_14562,N_14066,N_14034);
nor U14563 (N_14563,N_14346,N_13801);
nor U14564 (N_14564,N_14182,N_13845);
or U14565 (N_14565,N_13874,N_14307);
and U14566 (N_14566,N_13677,N_13625);
nand U14567 (N_14567,N_13689,N_13706);
nand U14568 (N_14568,N_14279,N_13602);
xor U14569 (N_14569,N_14108,N_13898);
and U14570 (N_14570,N_13844,N_14133);
nand U14571 (N_14571,N_14238,N_13707);
nor U14572 (N_14572,N_13629,N_13903);
nand U14573 (N_14573,N_14015,N_14349);
or U14574 (N_14574,N_13748,N_14062);
or U14575 (N_14575,N_14139,N_14185);
and U14576 (N_14576,N_13946,N_13936);
nand U14577 (N_14577,N_13868,N_14089);
nor U14578 (N_14578,N_14018,N_14344);
nor U14579 (N_14579,N_14090,N_13836);
or U14580 (N_14580,N_14289,N_14330);
nor U14581 (N_14581,N_13982,N_14389);
or U14582 (N_14582,N_14202,N_13976);
nor U14583 (N_14583,N_13896,N_14206);
and U14584 (N_14584,N_14225,N_14327);
nand U14585 (N_14585,N_13832,N_13829);
or U14586 (N_14586,N_14026,N_14000);
or U14587 (N_14587,N_14110,N_14375);
nand U14588 (N_14588,N_14138,N_14361);
or U14589 (N_14589,N_13893,N_13713);
nor U14590 (N_14590,N_13611,N_14164);
or U14591 (N_14591,N_13732,N_13692);
and U14592 (N_14592,N_13911,N_14112);
nor U14593 (N_14593,N_13855,N_13842);
nor U14594 (N_14594,N_13790,N_14055);
nor U14595 (N_14595,N_13939,N_13949);
nor U14596 (N_14596,N_13773,N_13609);
and U14597 (N_14597,N_13973,N_13752);
nor U14598 (N_14598,N_14197,N_14191);
or U14599 (N_14599,N_13808,N_14380);
or U14600 (N_14600,N_14388,N_13905);
or U14601 (N_14601,N_14369,N_13961);
nand U14602 (N_14602,N_14060,N_14175);
or U14603 (N_14603,N_14237,N_14041);
nand U14604 (N_14604,N_13652,N_14385);
and U14605 (N_14605,N_14332,N_13951);
nor U14606 (N_14606,N_13912,N_13834);
nand U14607 (N_14607,N_14005,N_13763);
or U14608 (N_14608,N_14212,N_14299);
and U14609 (N_14609,N_14278,N_14120);
nor U14610 (N_14610,N_13626,N_13884);
nand U14611 (N_14611,N_13852,N_14268);
nor U14612 (N_14612,N_14106,N_14124);
and U14613 (N_14613,N_13702,N_13984);
nand U14614 (N_14614,N_13672,N_13686);
nand U14615 (N_14615,N_14311,N_14115);
and U14616 (N_14616,N_14242,N_13631);
nand U14617 (N_14617,N_14273,N_13816);
nor U14618 (N_14618,N_13794,N_14379);
or U14619 (N_14619,N_13917,N_14309);
or U14620 (N_14620,N_13691,N_13835);
and U14621 (N_14621,N_14168,N_13819);
nand U14622 (N_14622,N_14350,N_14031);
nand U14623 (N_14623,N_13760,N_13805);
nand U14624 (N_14624,N_14383,N_14216);
nor U14625 (N_14625,N_14331,N_14272);
nor U14626 (N_14626,N_14039,N_13925);
or U14627 (N_14627,N_14003,N_14097);
nand U14628 (N_14628,N_14170,N_13880);
and U14629 (N_14629,N_13838,N_14249);
xor U14630 (N_14630,N_13849,N_14134);
nor U14631 (N_14631,N_14040,N_14105);
and U14632 (N_14632,N_14290,N_13734);
or U14633 (N_14633,N_14096,N_14017);
nand U14634 (N_14634,N_14007,N_14228);
and U14635 (N_14635,N_14044,N_13985);
or U14636 (N_14636,N_14250,N_13733);
or U14637 (N_14637,N_14313,N_13746);
and U14638 (N_14638,N_13612,N_13768);
nor U14639 (N_14639,N_13633,N_14343);
and U14640 (N_14640,N_14032,N_13698);
or U14641 (N_14641,N_13987,N_13650);
or U14642 (N_14642,N_14045,N_13833);
nor U14643 (N_14643,N_13681,N_13887);
nor U14644 (N_14644,N_14036,N_13727);
or U14645 (N_14645,N_14076,N_13618);
nor U14646 (N_14646,N_13954,N_14257);
or U14647 (N_14647,N_14226,N_13952);
nand U14648 (N_14648,N_13736,N_14364);
nor U14649 (N_14649,N_13703,N_14155);
or U14650 (N_14650,N_14276,N_13610);
nor U14651 (N_14651,N_13795,N_13941);
nand U14652 (N_14652,N_13739,N_14053);
nand U14653 (N_14653,N_14136,N_14288);
nor U14654 (N_14654,N_13922,N_13657);
or U14655 (N_14655,N_14174,N_13671);
or U14656 (N_14656,N_13632,N_14374);
nor U14657 (N_14657,N_13964,N_14284);
or U14658 (N_14658,N_13857,N_13688);
nor U14659 (N_14659,N_14001,N_13810);
nor U14660 (N_14660,N_13866,N_13882);
nor U14661 (N_14661,N_13929,N_14240);
nand U14662 (N_14662,N_14321,N_14148);
or U14663 (N_14663,N_13661,N_14122);
nand U14664 (N_14664,N_13754,N_13683);
nand U14665 (N_14665,N_13843,N_14265);
or U14666 (N_14666,N_14149,N_13651);
nor U14667 (N_14667,N_14020,N_13655);
nand U14668 (N_14668,N_14116,N_13854);
or U14669 (N_14669,N_13802,N_13621);
or U14670 (N_14670,N_13897,N_13628);
or U14671 (N_14671,N_13705,N_13724);
nand U14672 (N_14672,N_14075,N_14357);
and U14673 (N_14673,N_13830,N_13721);
and U14674 (N_14674,N_14292,N_14286);
or U14675 (N_14675,N_13701,N_14312);
or U14676 (N_14676,N_14169,N_14121);
and U14677 (N_14677,N_13678,N_13948);
and U14678 (N_14678,N_13615,N_14322);
or U14679 (N_14679,N_14338,N_13729);
nand U14680 (N_14680,N_13797,N_14390);
nand U14681 (N_14681,N_14201,N_13910);
or U14682 (N_14682,N_14303,N_13662);
nand U14683 (N_14683,N_14335,N_14009);
nor U14684 (N_14684,N_13870,N_13909);
nor U14685 (N_14685,N_14323,N_13674);
nor U14686 (N_14686,N_14215,N_13667);
nand U14687 (N_14687,N_13761,N_14156);
nand U14688 (N_14688,N_14310,N_14251);
nand U14689 (N_14689,N_13605,N_13983);
or U14690 (N_14690,N_13607,N_14029);
nor U14691 (N_14691,N_14333,N_14183);
and U14692 (N_14692,N_13828,N_13859);
or U14693 (N_14693,N_13860,N_13957);
nor U14694 (N_14694,N_14381,N_13891);
and U14695 (N_14695,N_14371,N_13735);
xor U14696 (N_14696,N_14324,N_13798);
nand U14697 (N_14697,N_14280,N_13682);
nor U14698 (N_14698,N_13956,N_13694);
and U14699 (N_14699,N_13991,N_13876);
or U14700 (N_14700,N_13731,N_13643);
nand U14701 (N_14701,N_13998,N_14398);
or U14702 (N_14702,N_13751,N_14198);
nand U14703 (N_14703,N_13640,N_14203);
nand U14704 (N_14704,N_14341,N_14236);
nand U14705 (N_14705,N_14051,N_14049);
and U14706 (N_14706,N_14188,N_13756);
and U14707 (N_14707,N_13890,N_13943);
nand U14708 (N_14708,N_13793,N_13995);
nand U14709 (N_14709,N_14208,N_13960);
nor U14710 (N_14710,N_14178,N_13792);
and U14711 (N_14711,N_13738,N_14302);
nor U14712 (N_14712,N_13636,N_14207);
nor U14713 (N_14713,N_14219,N_13840);
nand U14714 (N_14714,N_14141,N_13693);
nor U14715 (N_14715,N_13604,N_13879);
nor U14716 (N_14716,N_14382,N_13620);
or U14717 (N_14717,N_14028,N_13700);
or U14718 (N_14718,N_13892,N_14316);
and U14719 (N_14719,N_14192,N_14227);
or U14720 (N_14720,N_14153,N_14035);
and U14721 (N_14721,N_13779,N_14140);
and U14722 (N_14722,N_13869,N_13953);
nor U14723 (N_14723,N_13959,N_13673);
or U14724 (N_14724,N_13619,N_14118);
nand U14725 (N_14725,N_13979,N_14006);
nand U14726 (N_14726,N_13644,N_13930);
or U14727 (N_14727,N_14165,N_14314);
nor U14728 (N_14728,N_14078,N_14069);
nor U14729 (N_14729,N_14205,N_14073);
and U14730 (N_14730,N_14387,N_14101);
nand U14731 (N_14731,N_13663,N_13718);
nor U14732 (N_14732,N_13780,N_14091);
nor U14733 (N_14733,N_13647,N_14082);
or U14734 (N_14734,N_13856,N_14173);
nor U14735 (N_14735,N_13616,N_14099);
nor U14736 (N_14736,N_13809,N_13824);
nor U14737 (N_14737,N_14386,N_13873);
and U14738 (N_14738,N_13990,N_14255);
nand U14739 (N_14739,N_13877,N_14088);
nand U14740 (N_14740,N_14376,N_14057);
nand U14741 (N_14741,N_14154,N_14353);
or U14742 (N_14742,N_13716,N_13980);
or U14743 (N_14743,N_14320,N_14368);
nor U14744 (N_14744,N_14214,N_13886);
or U14745 (N_14745,N_13817,N_13996);
and U14746 (N_14746,N_14095,N_14166);
nor U14747 (N_14747,N_13789,N_14260);
and U14748 (N_14748,N_13743,N_14030);
nor U14749 (N_14749,N_13627,N_14144);
or U14750 (N_14750,N_13883,N_13965);
and U14751 (N_14751,N_14063,N_13837);
or U14752 (N_14752,N_14365,N_13603);
and U14753 (N_14753,N_14162,N_14137);
nand U14754 (N_14754,N_13811,N_13608);
and U14755 (N_14755,N_14209,N_14305);
and U14756 (N_14756,N_14275,N_13839);
nor U14757 (N_14757,N_14125,N_14043);
and U14758 (N_14758,N_13966,N_14172);
and U14759 (N_14759,N_14223,N_13831);
nand U14760 (N_14760,N_14328,N_14282);
or U14761 (N_14761,N_14094,N_14199);
nand U14762 (N_14762,N_14079,N_13865);
and U14763 (N_14763,N_13871,N_13928);
nor U14764 (N_14764,N_14336,N_14065);
or U14765 (N_14765,N_14297,N_13937);
nand U14766 (N_14766,N_13872,N_14392);
nand U14767 (N_14767,N_13900,N_13851);
or U14768 (N_14768,N_14246,N_13978);
and U14769 (N_14769,N_13894,N_13665);
nand U14770 (N_14770,N_13784,N_14190);
nand U14771 (N_14771,N_14233,N_13728);
nor U14772 (N_14772,N_13913,N_13878);
and U14773 (N_14773,N_13782,N_14352);
or U14774 (N_14774,N_14033,N_13932);
and U14775 (N_14775,N_13613,N_13699);
and U14776 (N_14776,N_14184,N_13902);
nor U14777 (N_14777,N_13755,N_14042);
nor U14778 (N_14778,N_14059,N_14016);
or U14779 (N_14779,N_14061,N_14087);
and U14780 (N_14780,N_13823,N_14158);
and U14781 (N_14781,N_14080,N_13659);
nor U14782 (N_14782,N_14210,N_14142);
nor U14783 (N_14783,N_14262,N_13772);
nor U14784 (N_14784,N_14012,N_13685);
and U14785 (N_14785,N_14187,N_13750);
and U14786 (N_14786,N_13758,N_14123);
or U14787 (N_14787,N_13899,N_13696);
nor U14788 (N_14788,N_14100,N_13826);
nor U14789 (N_14789,N_13927,N_14253);
nand U14790 (N_14790,N_13997,N_13614);
or U14791 (N_14791,N_13875,N_14176);
nand U14792 (N_14792,N_14362,N_14131);
nor U14793 (N_14793,N_13744,N_14010);
nand U14794 (N_14794,N_13720,N_13778);
and U14795 (N_14795,N_14111,N_13617);
xor U14796 (N_14796,N_13679,N_13993);
nand U14797 (N_14797,N_14181,N_14054);
and U14798 (N_14798,N_14300,N_14104);
nand U14799 (N_14799,N_13821,N_14002);
xor U14800 (N_14800,N_14053,N_13866);
and U14801 (N_14801,N_13950,N_14301);
nor U14802 (N_14802,N_13893,N_13685);
nor U14803 (N_14803,N_14049,N_14158);
nor U14804 (N_14804,N_13603,N_13912);
and U14805 (N_14805,N_14044,N_13680);
nand U14806 (N_14806,N_13601,N_14129);
or U14807 (N_14807,N_14196,N_13998);
nand U14808 (N_14808,N_14270,N_13618);
nor U14809 (N_14809,N_13831,N_13781);
nand U14810 (N_14810,N_13926,N_14366);
and U14811 (N_14811,N_13791,N_13617);
and U14812 (N_14812,N_13857,N_14031);
nand U14813 (N_14813,N_14066,N_13893);
and U14814 (N_14814,N_13861,N_13625);
and U14815 (N_14815,N_13825,N_14164);
and U14816 (N_14816,N_14124,N_13846);
nor U14817 (N_14817,N_14268,N_13707);
nor U14818 (N_14818,N_14364,N_14373);
or U14819 (N_14819,N_14106,N_14162);
nand U14820 (N_14820,N_13806,N_13898);
nand U14821 (N_14821,N_14140,N_14049);
nand U14822 (N_14822,N_14058,N_13634);
nand U14823 (N_14823,N_13994,N_14219);
and U14824 (N_14824,N_13610,N_13922);
nand U14825 (N_14825,N_13722,N_14101);
or U14826 (N_14826,N_13873,N_13817);
and U14827 (N_14827,N_14172,N_13672);
xor U14828 (N_14828,N_13906,N_13817);
nor U14829 (N_14829,N_13805,N_13675);
nor U14830 (N_14830,N_14251,N_14243);
nor U14831 (N_14831,N_14215,N_14218);
nor U14832 (N_14832,N_13990,N_14269);
or U14833 (N_14833,N_14196,N_13953);
nand U14834 (N_14834,N_13782,N_14373);
or U14835 (N_14835,N_14381,N_14339);
nor U14836 (N_14836,N_13847,N_13743);
nand U14837 (N_14837,N_14149,N_13623);
nor U14838 (N_14838,N_14390,N_13773);
nor U14839 (N_14839,N_13698,N_14177);
or U14840 (N_14840,N_14168,N_13805);
or U14841 (N_14841,N_13715,N_13665);
and U14842 (N_14842,N_14043,N_14253);
nand U14843 (N_14843,N_14373,N_13778);
nor U14844 (N_14844,N_14188,N_14156);
and U14845 (N_14845,N_13914,N_13656);
nor U14846 (N_14846,N_13830,N_13926);
nor U14847 (N_14847,N_13746,N_14100);
nand U14848 (N_14848,N_13799,N_13821);
or U14849 (N_14849,N_13601,N_13723);
or U14850 (N_14850,N_13854,N_13807);
or U14851 (N_14851,N_14295,N_14256);
or U14852 (N_14852,N_14357,N_13916);
and U14853 (N_14853,N_13670,N_13676);
nor U14854 (N_14854,N_14325,N_13809);
nand U14855 (N_14855,N_14171,N_14331);
and U14856 (N_14856,N_14266,N_13917);
nor U14857 (N_14857,N_13865,N_13974);
and U14858 (N_14858,N_14386,N_14361);
nand U14859 (N_14859,N_13731,N_14009);
or U14860 (N_14860,N_13761,N_14312);
or U14861 (N_14861,N_14293,N_14008);
nor U14862 (N_14862,N_14230,N_14234);
or U14863 (N_14863,N_13963,N_13726);
and U14864 (N_14864,N_13925,N_14141);
nor U14865 (N_14865,N_13901,N_14380);
or U14866 (N_14866,N_13924,N_14397);
or U14867 (N_14867,N_14152,N_14087);
or U14868 (N_14868,N_14041,N_13673);
or U14869 (N_14869,N_13897,N_13639);
nor U14870 (N_14870,N_13891,N_13845);
or U14871 (N_14871,N_14068,N_13860);
or U14872 (N_14872,N_13798,N_14077);
or U14873 (N_14873,N_14152,N_14226);
and U14874 (N_14874,N_14233,N_13732);
nand U14875 (N_14875,N_13801,N_14215);
or U14876 (N_14876,N_13950,N_13759);
or U14877 (N_14877,N_13811,N_14058);
nand U14878 (N_14878,N_14101,N_13655);
nor U14879 (N_14879,N_13779,N_13921);
nor U14880 (N_14880,N_14092,N_13915);
nand U14881 (N_14881,N_13853,N_14179);
or U14882 (N_14882,N_14164,N_14110);
nand U14883 (N_14883,N_14035,N_13697);
and U14884 (N_14884,N_14092,N_13882);
nor U14885 (N_14885,N_13677,N_14000);
and U14886 (N_14886,N_13881,N_14104);
nor U14887 (N_14887,N_14112,N_13780);
and U14888 (N_14888,N_14179,N_13970);
and U14889 (N_14889,N_14190,N_13858);
and U14890 (N_14890,N_14351,N_14173);
nand U14891 (N_14891,N_13696,N_13990);
or U14892 (N_14892,N_13813,N_13810);
nor U14893 (N_14893,N_13736,N_14360);
nand U14894 (N_14894,N_13838,N_14027);
or U14895 (N_14895,N_13919,N_14127);
and U14896 (N_14896,N_13770,N_13686);
nor U14897 (N_14897,N_14211,N_14222);
and U14898 (N_14898,N_13991,N_14394);
nand U14899 (N_14899,N_13698,N_13997);
and U14900 (N_14900,N_14262,N_14098);
nand U14901 (N_14901,N_13899,N_13629);
or U14902 (N_14902,N_14170,N_14393);
and U14903 (N_14903,N_14183,N_14012);
and U14904 (N_14904,N_14236,N_14339);
and U14905 (N_14905,N_14144,N_14044);
and U14906 (N_14906,N_13609,N_13757);
nand U14907 (N_14907,N_13802,N_14334);
or U14908 (N_14908,N_14098,N_13793);
or U14909 (N_14909,N_13805,N_13753);
nor U14910 (N_14910,N_13994,N_14163);
or U14911 (N_14911,N_14293,N_13693);
or U14912 (N_14912,N_13797,N_13792);
nor U14913 (N_14913,N_14034,N_13705);
nor U14914 (N_14914,N_13678,N_14244);
nor U14915 (N_14915,N_14324,N_13680);
or U14916 (N_14916,N_14074,N_14065);
nand U14917 (N_14917,N_14261,N_14057);
or U14918 (N_14918,N_13804,N_13743);
nand U14919 (N_14919,N_13839,N_14395);
and U14920 (N_14920,N_13649,N_13840);
or U14921 (N_14921,N_13714,N_14043);
nor U14922 (N_14922,N_14276,N_13629);
nor U14923 (N_14923,N_14358,N_13863);
nor U14924 (N_14924,N_13934,N_14356);
nor U14925 (N_14925,N_13797,N_14135);
nand U14926 (N_14926,N_14358,N_13708);
nor U14927 (N_14927,N_13890,N_13836);
and U14928 (N_14928,N_13751,N_14012);
nor U14929 (N_14929,N_14228,N_13814);
nor U14930 (N_14930,N_13986,N_14241);
nand U14931 (N_14931,N_13787,N_13970);
or U14932 (N_14932,N_14193,N_13700);
xnor U14933 (N_14933,N_13622,N_14330);
and U14934 (N_14934,N_13988,N_13684);
nor U14935 (N_14935,N_14296,N_14372);
and U14936 (N_14936,N_14218,N_13895);
and U14937 (N_14937,N_13963,N_14012);
nand U14938 (N_14938,N_13759,N_13654);
or U14939 (N_14939,N_13860,N_13759);
or U14940 (N_14940,N_14101,N_13716);
and U14941 (N_14941,N_14085,N_14184);
or U14942 (N_14942,N_14154,N_13829);
and U14943 (N_14943,N_13771,N_14164);
and U14944 (N_14944,N_14321,N_14244);
nor U14945 (N_14945,N_13752,N_14061);
xor U14946 (N_14946,N_13955,N_14117);
and U14947 (N_14947,N_13923,N_14330);
and U14948 (N_14948,N_14357,N_14059);
or U14949 (N_14949,N_13813,N_14215);
nand U14950 (N_14950,N_14253,N_13813);
nand U14951 (N_14951,N_14308,N_13908);
or U14952 (N_14952,N_14216,N_14126);
or U14953 (N_14953,N_13972,N_14380);
nor U14954 (N_14954,N_14380,N_14390);
nand U14955 (N_14955,N_13694,N_14068);
or U14956 (N_14956,N_13623,N_13689);
nor U14957 (N_14957,N_13644,N_14280);
and U14958 (N_14958,N_14282,N_13718);
and U14959 (N_14959,N_13795,N_14109);
or U14960 (N_14960,N_13701,N_14357);
nor U14961 (N_14961,N_14085,N_13850);
nand U14962 (N_14962,N_14295,N_14241);
and U14963 (N_14963,N_14008,N_14287);
nand U14964 (N_14964,N_14233,N_13608);
nor U14965 (N_14965,N_14034,N_13641);
or U14966 (N_14966,N_13942,N_14222);
and U14967 (N_14967,N_13729,N_14197);
and U14968 (N_14968,N_14157,N_14374);
nand U14969 (N_14969,N_14354,N_13897);
nor U14970 (N_14970,N_13822,N_14334);
nor U14971 (N_14971,N_14114,N_13822);
nand U14972 (N_14972,N_14396,N_14219);
or U14973 (N_14973,N_14087,N_13814);
nand U14974 (N_14974,N_13900,N_13665);
nor U14975 (N_14975,N_14373,N_14269);
nor U14976 (N_14976,N_14198,N_13901);
or U14977 (N_14977,N_13652,N_13842);
or U14978 (N_14978,N_14142,N_13632);
nand U14979 (N_14979,N_14157,N_14358);
nand U14980 (N_14980,N_14091,N_14154);
nand U14981 (N_14981,N_13870,N_14005);
nand U14982 (N_14982,N_13881,N_14052);
nor U14983 (N_14983,N_13795,N_13607);
nand U14984 (N_14984,N_13794,N_13927);
or U14985 (N_14985,N_13785,N_13728);
nand U14986 (N_14986,N_14248,N_13762);
nand U14987 (N_14987,N_14289,N_14343);
nor U14988 (N_14988,N_14333,N_14351);
nor U14989 (N_14989,N_14368,N_14043);
nand U14990 (N_14990,N_13626,N_13693);
nor U14991 (N_14991,N_13613,N_13824);
nand U14992 (N_14992,N_14037,N_13753);
nand U14993 (N_14993,N_14136,N_13912);
nor U14994 (N_14994,N_13661,N_14074);
or U14995 (N_14995,N_14003,N_13672);
or U14996 (N_14996,N_13739,N_13906);
nor U14997 (N_14997,N_13830,N_14089);
or U14998 (N_14998,N_14114,N_14379);
and U14999 (N_14999,N_13933,N_14253);
or U15000 (N_15000,N_13865,N_13778);
or U15001 (N_15001,N_14093,N_14133);
nand U15002 (N_15002,N_13628,N_14313);
and U15003 (N_15003,N_14269,N_14086);
or U15004 (N_15004,N_14059,N_13699);
nand U15005 (N_15005,N_13990,N_13833);
and U15006 (N_15006,N_13886,N_13862);
nand U15007 (N_15007,N_13984,N_13611);
and U15008 (N_15008,N_14258,N_13672);
or U15009 (N_15009,N_13867,N_14307);
nor U15010 (N_15010,N_13907,N_13825);
nor U15011 (N_15011,N_13606,N_14347);
nand U15012 (N_15012,N_13904,N_13646);
nand U15013 (N_15013,N_13963,N_14204);
nor U15014 (N_15014,N_13642,N_14287);
or U15015 (N_15015,N_13940,N_14278);
or U15016 (N_15016,N_14085,N_14293);
nor U15017 (N_15017,N_14204,N_13608);
nor U15018 (N_15018,N_13943,N_14177);
nand U15019 (N_15019,N_14195,N_13793);
and U15020 (N_15020,N_13607,N_14038);
and U15021 (N_15021,N_13626,N_13794);
nor U15022 (N_15022,N_14268,N_14354);
nand U15023 (N_15023,N_13641,N_13992);
and U15024 (N_15024,N_14281,N_14038);
or U15025 (N_15025,N_13815,N_13768);
nor U15026 (N_15026,N_14171,N_14280);
nand U15027 (N_15027,N_14293,N_14218);
nand U15028 (N_15028,N_14293,N_13716);
and U15029 (N_15029,N_14333,N_13840);
nor U15030 (N_15030,N_14290,N_14264);
or U15031 (N_15031,N_13749,N_13844);
xor U15032 (N_15032,N_13688,N_13715);
or U15033 (N_15033,N_14308,N_13779);
and U15034 (N_15034,N_13889,N_13662);
or U15035 (N_15035,N_13914,N_13678);
and U15036 (N_15036,N_13847,N_13749);
nand U15037 (N_15037,N_14205,N_14262);
or U15038 (N_15038,N_14399,N_14386);
nor U15039 (N_15039,N_13715,N_14190);
nand U15040 (N_15040,N_13967,N_14394);
or U15041 (N_15041,N_13816,N_14100);
nand U15042 (N_15042,N_13635,N_14205);
and U15043 (N_15043,N_14240,N_14008);
and U15044 (N_15044,N_13720,N_14279);
and U15045 (N_15045,N_13647,N_14139);
or U15046 (N_15046,N_14044,N_14289);
nor U15047 (N_15047,N_13601,N_14079);
and U15048 (N_15048,N_14104,N_13769);
and U15049 (N_15049,N_14157,N_13606);
and U15050 (N_15050,N_13662,N_14242);
or U15051 (N_15051,N_13996,N_13668);
nand U15052 (N_15052,N_13828,N_14358);
or U15053 (N_15053,N_13843,N_14150);
nor U15054 (N_15054,N_14194,N_14230);
nand U15055 (N_15055,N_13614,N_13730);
and U15056 (N_15056,N_13756,N_14168);
nand U15057 (N_15057,N_14194,N_14241);
nor U15058 (N_15058,N_14273,N_14262);
and U15059 (N_15059,N_14197,N_13750);
nor U15060 (N_15060,N_13873,N_14129);
nand U15061 (N_15061,N_14011,N_14155);
nor U15062 (N_15062,N_14365,N_13946);
nand U15063 (N_15063,N_13994,N_14107);
nand U15064 (N_15064,N_13707,N_13675);
nor U15065 (N_15065,N_13712,N_13784);
or U15066 (N_15066,N_13972,N_13870);
nand U15067 (N_15067,N_14180,N_13623);
or U15068 (N_15068,N_14074,N_13615);
nand U15069 (N_15069,N_13841,N_14219);
nor U15070 (N_15070,N_13716,N_13776);
nand U15071 (N_15071,N_13633,N_13610);
xor U15072 (N_15072,N_14289,N_13906);
or U15073 (N_15073,N_14285,N_13774);
or U15074 (N_15074,N_13760,N_14296);
nor U15075 (N_15075,N_13790,N_14016);
and U15076 (N_15076,N_14399,N_14158);
nor U15077 (N_15077,N_14077,N_13922);
and U15078 (N_15078,N_13765,N_14123);
and U15079 (N_15079,N_14009,N_14152);
and U15080 (N_15080,N_14385,N_14032);
nand U15081 (N_15081,N_14216,N_14049);
nand U15082 (N_15082,N_13842,N_14033);
nand U15083 (N_15083,N_13990,N_13960);
nand U15084 (N_15084,N_13995,N_14197);
nor U15085 (N_15085,N_13628,N_13811);
or U15086 (N_15086,N_13951,N_13835);
or U15087 (N_15087,N_14007,N_14332);
or U15088 (N_15088,N_13848,N_14361);
nand U15089 (N_15089,N_13984,N_13795);
nand U15090 (N_15090,N_13888,N_13909);
and U15091 (N_15091,N_14147,N_14176);
and U15092 (N_15092,N_13661,N_13694);
or U15093 (N_15093,N_13657,N_14392);
nor U15094 (N_15094,N_13737,N_13697);
and U15095 (N_15095,N_14222,N_14276);
or U15096 (N_15096,N_13694,N_14330);
and U15097 (N_15097,N_14010,N_13977);
nor U15098 (N_15098,N_13776,N_13748);
or U15099 (N_15099,N_14197,N_13784);
nand U15100 (N_15100,N_13619,N_14132);
nor U15101 (N_15101,N_13946,N_14267);
or U15102 (N_15102,N_13956,N_13930);
nand U15103 (N_15103,N_14275,N_14346);
and U15104 (N_15104,N_13923,N_13726);
and U15105 (N_15105,N_14267,N_14285);
or U15106 (N_15106,N_13998,N_14098);
nand U15107 (N_15107,N_14276,N_14253);
or U15108 (N_15108,N_14080,N_13848);
nor U15109 (N_15109,N_14094,N_13705);
nand U15110 (N_15110,N_14048,N_14370);
or U15111 (N_15111,N_13632,N_14328);
nor U15112 (N_15112,N_13623,N_14382);
nand U15113 (N_15113,N_13855,N_13862);
and U15114 (N_15114,N_14214,N_13754);
nand U15115 (N_15115,N_13687,N_13922);
nor U15116 (N_15116,N_13928,N_14033);
and U15117 (N_15117,N_14274,N_13691);
and U15118 (N_15118,N_14064,N_14170);
nor U15119 (N_15119,N_14277,N_14092);
nand U15120 (N_15120,N_13814,N_13737);
nand U15121 (N_15121,N_13604,N_13749);
nand U15122 (N_15122,N_14280,N_13716);
and U15123 (N_15123,N_14015,N_14123);
nand U15124 (N_15124,N_14003,N_14163);
nand U15125 (N_15125,N_13965,N_14080);
nor U15126 (N_15126,N_13729,N_14383);
nand U15127 (N_15127,N_13730,N_14055);
and U15128 (N_15128,N_13744,N_14236);
and U15129 (N_15129,N_14245,N_14049);
nand U15130 (N_15130,N_13835,N_13767);
and U15131 (N_15131,N_14011,N_14229);
or U15132 (N_15132,N_14178,N_13603);
or U15133 (N_15133,N_14194,N_13793);
nor U15134 (N_15134,N_14300,N_13681);
or U15135 (N_15135,N_14386,N_13967);
or U15136 (N_15136,N_13908,N_13961);
or U15137 (N_15137,N_14374,N_13759);
and U15138 (N_15138,N_13974,N_13667);
nand U15139 (N_15139,N_13608,N_14025);
nand U15140 (N_15140,N_14250,N_13624);
nor U15141 (N_15141,N_14391,N_13693);
and U15142 (N_15142,N_13868,N_14274);
and U15143 (N_15143,N_14376,N_13883);
and U15144 (N_15144,N_14161,N_14157);
and U15145 (N_15145,N_13902,N_14295);
and U15146 (N_15146,N_13951,N_14397);
nand U15147 (N_15147,N_13620,N_14156);
or U15148 (N_15148,N_13671,N_13682);
nor U15149 (N_15149,N_13735,N_14017);
nor U15150 (N_15150,N_14187,N_13781);
nor U15151 (N_15151,N_13756,N_14258);
and U15152 (N_15152,N_14383,N_13892);
and U15153 (N_15153,N_14391,N_13703);
and U15154 (N_15154,N_14193,N_13882);
nand U15155 (N_15155,N_14076,N_13896);
or U15156 (N_15156,N_13761,N_13656);
and U15157 (N_15157,N_14025,N_13649);
or U15158 (N_15158,N_14051,N_13776);
nor U15159 (N_15159,N_13886,N_14098);
or U15160 (N_15160,N_14287,N_13945);
and U15161 (N_15161,N_13601,N_14180);
nand U15162 (N_15162,N_13851,N_13610);
nor U15163 (N_15163,N_14225,N_14265);
nand U15164 (N_15164,N_14201,N_14207);
or U15165 (N_15165,N_13910,N_14058);
nor U15166 (N_15166,N_13803,N_13703);
nor U15167 (N_15167,N_14397,N_13747);
and U15168 (N_15168,N_13705,N_13804);
nor U15169 (N_15169,N_13840,N_14029);
and U15170 (N_15170,N_14256,N_13806);
nand U15171 (N_15171,N_14085,N_13624);
or U15172 (N_15172,N_13750,N_13758);
nand U15173 (N_15173,N_13686,N_13791);
or U15174 (N_15174,N_14390,N_14119);
nand U15175 (N_15175,N_14199,N_13722);
and U15176 (N_15176,N_14076,N_13714);
and U15177 (N_15177,N_13842,N_14264);
nor U15178 (N_15178,N_14238,N_13696);
nand U15179 (N_15179,N_13625,N_14085);
or U15180 (N_15180,N_14264,N_14286);
and U15181 (N_15181,N_13753,N_13779);
and U15182 (N_15182,N_14064,N_14328);
nand U15183 (N_15183,N_13784,N_13725);
nor U15184 (N_15184,N_13739,N_14200);
nand U15185 (N_15185,N_14305,N_13783);
or U15186 (N_15186,N_13974,N_13658);
nand U15187 (N_15187,N_14095,N_13955);
nor U15188 (N_15188,N_14298,N_13615);
and U15189 (N_15189,N_14204,N_14030);
and U15190 (N_15190,N_14256,N_13972);
xor U15191 (N_15191,N_14089,N_14283);
and U15192 (N_15192,N_13810,N_13619);
nand U15193 (N_15193,N_14053,N_14033);
nor U15194 (N_15194,N_13958,N_13841);
nor U15195 (N_15195,N_13886,N_13813);
or U15196 (N_15196,N_14178,N_13703);
or U15197 (N_15197,N_13845,N_14257);
nor U15198 (N_15198,N_14049,N_14162);
nor U15199 (N_15199,N_14051,N_13666);
nor U15200 (N_15200,N_14500,N_14727);
nand U15201 (N_15201,N_14568,N_14878);
nor U15202 (N_15202,N_14803,N_15115);
nor U15203 (N_15203,N_14760,N_15055);
nand U15204 (N_15204,N_14444,N_14574);
or U15205 (N_15205,N_14520,N_14653);
or U15206 (N_15206,N_14449,N_15099);
nand U15207 (N_15207,N_14741,N_14692);
or U15208 (N_15208,N_14994,N_14590);
or U15209 (N_15209,N_14579,N_14557);
or U15210 (N_15210,N_14804,N_14441);
or U15211 (N_15211,N_14596,N_14640);
nand U15212 (N_15212,N_14863,N_14756);
nand U15213 (N_15213,N_14715,N_15067);
nand U15214 (N_15214,N_15134,N_14573);
nand U15215 (N_15215,N_14890,N_14752);
and U15216 (N_15216,N_14602,N_14676);
nor U15217 (N_15217,N_15191,N_15151);
or U15218 (N_15218,N_15053,N_14838);
nand U15219 (N_15219,N_14896,N_14782);
nand U15220 (N_15220,N_14543,N_14980);
and U15221 (N_15221,N_14469,N_14758);
and U15222 (N_15222,N_14660,N_14981);
and U15223 (N_15223,N_14502,N_14612);
nand U15224 (N_15224,N_15188,N_14928);
nand U15225 (N_15225,N_14737,N_14765);
nor U15226 (N_15226,N_15157,N_14996);
or U15227 (N_15227,N_14569,N_15068);
or U15228 (N_15228,N_14824,N_14535);
nand U15229 (N_15229,N_15036,N_14817);
nor U15230 (N_15230,N_15193,N_14932);
or U15231 (N_15231,N_14903,N_14806);
and U15232 (N_15232,N_14443,N_14982);
or U15233 (N_15233,N_14517,N_14632);
nand U15234 (N_15234,N_15081,N_14537);
and U15235 (N_15235,N_14889,N_14914);
or U15236 (N_15236,N_14467,N_14807);
or U15237 (N_15237,N_15167,N_14948);
or U15238 (N_15238,N_14839,N_14603);
nor U15239 (N_15239,N_14910,N_14462);
nor U15240 (N_15240,N_14565,N_14563);
nor U15241 (N_15241,N_15077,N_14691);
nor U15242 (N_15242,N_15040,N_15039);
or U15243 (N_15243,N_14466,N_14822);
nand U15244 (N_15244,N_14470,N_14965);
nand U15245 (N_15245,N_15025,N_14987);
or U15246 (N_15246,N_15139,N_14472);
and U15247 (N_15247,N_15061,N_14908);
nand U15248 (N_15248,N_14915,N_15083);
nor U15249 (N_15249,N_14954,N_14417);
nor U15250 (N_15250,N_14882,N_14551);
nor U15251 (N_15251,N_14595,N_14798);
nand U15252 (N_15252,N_14825,N_14820);
or U15253 (N_15253,N_14944,N_14591);
nand U15254 (N_15254,N_14459,N_14518);
nor U15255 (N_15255,N_15108,N_14841);
nor U15256 (N_15256,N_14924,N_14753);
and U15257 (N_15257,N_14904,N_14522);
or U15258 (N_15258,N_14962,N_15159);
nor U15259 (N_15259,N_14463,N_14643);
and U15260 (N_15260,N_15003,N_14983);
nor U15261 (N_15261,N_14990,N_15112);
and U15262 (N_15262,N_15042,N_14668);
and U15263 (N_15263,N_14770,N_15072);
or U15264 (N_15264,N_14821,N_14431);
nor U15265 (N_15265,N_14750,N_15073);
or U15266 (N_15266,N_14402,N_14546);
and U15267 (N_15267,N_14702,N_14625);
nor U15268 (N_15268,N_14508,N_14687);
nor U15269 (N_15269,N_14411,N_14641);
nand U15270 (N_15270,N_14634,N_14891);
and U15271 (N_15271,N_14425,N_15132);
nor U15272 (N_15272,N_14456,N_14902);
or U15273 (N_15273,N_14626,N_15175);
nor U15274 (N_15274,N_14638,N_14706);
nor U15275 (N_15275,N_15044,N_14859);
or U15276 (N_15276,N_14974,N_14696);
or U15277 (N_15277,N_15030,N_14805);
and U15278 (N_15278,N_15095,N_15001);
and U15279 (N_15279,N_15093,N_15023);
and U15280 (N_15280,N_14482,N_14658);
and U15281 (N_15281,N_14724,N_14869);
or U15282 (N_15282,N_14480,N_14471);
nand U15283 (N_15283,N_14585,N_15172);
nor U15284 (N_15284,N_15084,N_14465);
or U15285 (N_15285,N_14736,N_14645);
and U15286 (N_15286,N_14986,N_14504);
and U15287 (N_15287,N_14850,N_15153);
nor U15288 (N_15288,N_14652,N_14498);
and U15289 (N_15289,N_14671,N_14515);
xor U15290 (N_15290,N_15104,N_14985);
nand U15291 (N_15291,N_14420,N_14777);
nand U15292 (N_15292,N_14588,N_14792);
nor U15293 (N_15293,N_14661,N_15190);
or U15294 (N_15294,N_14826,N_14672);
nor U15295 (N_15295,N_14647,N_14446);
nand U15296 (N_15296,N_15179,N_15165);
nor U15297 (N_15297,N_14966,N_15018);
nor U15298 (N_15298,N_14969,N_14973);
nor U15299 (N_15299,N_14992,N_14607);
nand U15300 (N_15300,N_14938,N_14450);
nand U15301 (N_15301,N_14561,N_14552);
or U15302 (N_15302,N_14527,N_14766);
nor U15303 (N_15303,N_14485,N_15079);
and U15304 (N_15304,N_14418,N_14873);
or U15305 (N_15305,N_14440,N_15140);
and U15306 (N_15306,N_14707,N_14955);
or U15307 (N_15307,N_14454,N_15103);
nand U15308 (N_15308,N_14490,N_14748);
and U15309 (N_15309,N_15074,N_14744);
nand U15310 (N_15310,N_15135,N_14587);
nand U15311 (N_15311,N_14559,N_14649);
or U15312 (N_15312,N_15120,N_14830);
and U15313 (N_15313,N_15002,N_15124);
and U15314 (N_15314,N_14633,N_15090);
or U15315 (N_15315,N_14534,N_14494);
and U15316 (N_15316,N_14870,N_14808);
and U15317 (N_15317,N_14790,N_14922);
nor U15318 (N_15318,N_14430,N_14679);
nand U15319 (N_15319,N_14959,N_14894);
and U15320 (N_15320,N_15060,N_15008);
nor U15321 (N_15321,N_14503,N_14725);
and U15322 (N_15322,N_14414,N_15184);
and U15323 (N_15323,N_14913,N_14867);
nor U15324 (N_15324,N_14438,N_15071);
nor U15325 (N_15325,N_14723,N_15037);
or U15326 (N_15326,N_14769,N_14428);
nor U15327 (N_15327,N_14422,N_14495);
nand U15328 (N_15328,N_14875,N_14678);
and U15329 (N_15329,N_14631,N_14989);
and U15330 (N_15330,N_15075,N_14593);
or U15331 (N_15331,N_15088,N_14709);
or U15332 (N_15332,N_15106,N_14885);
or U15333 (N_15333,N_14476,N_14917);
or U15334 (N_15334,N_14510,N_14564);
nor U15335 (N_15335,N_14815,N_14762);
and U15336 (N_15336,N_14683,N_14993);
nor U15337 (N_15337,N_15102,N_14613);
nand U15338 (N_15338,N_14542,N_14720);
and U15339 (N_15339,N_14560,N_14555);
nand U15340 (N_15340,N_14621,N_14615);
and U15341 (N_15341,N_14572,N_14868);
xnor U15342 (N_15342,N_14541,N_14710);
nand U15343 (N_15343,N_14733,N_14916);
nand U15344 (N_15344,N_14995,N_14481);
or U15345 (N_15345,N_14478,N_14599);
or U15346 (N_15346,N_14496,N_15000);
nand U15347 (N_15347,N_14623,N_14856);
nand U15348 (N_15348,N_15187,N_15035);
and U15349 (N_15349,N_14403,N_15137);
nand U15350 (N_15350,N_15130,N_14905);
and U15351 (N_15351,N_14881,N_14968);
nand U15352 (N_15352,N_14434,N_15101);
xor U15353 (N_15353,N_14688,N_14547);
nand U15354 (N_15354,N_15051,N_15062);
nor U15355 (N_15355,N_14637,N_14909);
nand U15356 (N_15356,N_14519,N_14943);
nand U15357 (N_15357,N_14600,N_14899);
and U15358 (N_15358,N_14785,N_14664);
nand U15359 (N_15359,N_15082,N_14415);
and U15360 (N_15360,N_14852,N_15136);
and U15361 (N_15361,N_14705,N_14700);
and U15362 (N_15362,N_14442,N_14473);
or U15363 (N_15363,N_14963,N_15152);
or U15364 (N_15364,N_14594,N_14605);
nor U15365 (N_15365,N_14616,N_14492);
nor U15366 (N_15366,N_14505,N_14728);
and U15367 (N_15367,N_14920,N_14578);
or U15368 (N_15368,N_14703,N_14684);
or U15369 (N_15369,N_14864,N_15141);
and U15370 (N_15370,N_14521,N_14925);
and U15371 (N_15371,N_14988,N_15015);
nor U15372 (N_15372,N_14536,N_14892);
and U15373 (N_15373,N_15007,N_14501);
or U15374 (N_15374,N_14774,N_14732);
or U15375 (N_15375,N_14712,N_14975);
nand U15376 (N_15376,N_14775,N_14836);
nand U15377 (N_15377,N_14796,N_14718);
or U15378 (N_15378,N_14639,N_15066);
nor U15379 (N_15379,N_15195,N_14675);
or U15380 (N_15380,N_14862,N_15024);
and U15381 (N_15381,N_14432,N_14749);
nor U15382 (N_15382,N_14998,N_15004);
nor U15383 (N_15383,N_15078,N_14512);
nor U15384 (N_15384,N_15125,N_14934);
nor U15385 (N_15385,N_14538,N_14754);
or U15386 (N_15386,N_14942,N_15100);
or U15387 (N_15387,N_15047,N_14423);
nand U15388 (N_15388,N_15183,N_15026);
and U15389 (N_15389,N_14514,N_14642);
and U15390 (N_15390,N_14818,N_15138);
nor U15391 (N_15391,N_15022,N_14907);
nand U15392 (N_15392,N_14738,N_14970);
nor U15393 (N_15393,N_14961,N_14735);
and U15394 (N_15394,N_14606,N_15017);
and U15395 (N_15395,N_14483,N_14813);
nor U15396 (N_15396,N_14567,N_14947);
or U15397 (N_15397,N_14648,N_14939);
and U15398 (N_15398,N_15057,N_14513);
or U15399 (N_15399,N_14693,N_15176);
nor U15400 (N_15400,N_14949,N_15189);
nor U15401 (N_15401,N_14831,N_14845);
nand U15402 (N_15402,N_14898,N_14577);
or U15403 (N_15403,N_15194,N_14529);
nor U15404 (N_15404,N_14722,N_15052);
nor U15405 (N_15405,N_14837,N_14767);
nand U15406 (N_15406,N_15021,N_14719);
or U15407 (N_15407,N_14582,N_15177);
and U15408 (N_15408,N_14400,N_14778);
nand U15409 (N_15409,N_15064,N_14657);
nand U15410 (N_15410,N_15043,N_14779);
and U15411 (N_15411,N_14698,N_14620);
nor U15412 (N_15412,N_14636,N_14714);
and U15413 (N_15413,N_15121,N_15110);
or U15414 (N_15414,N_15063,N_14933);
or U15415 (N_15415,N_14865,N_14419);
nor U15416 (N_15416,N_14776,N_14751);
nand U15417 (N_15417,N_15109,N_15196);
and U15418 (N_15418,N_14608,N_14405);
and U15419 (N_15419,N_14956,N_14911);
and U15420 (N_15420,N_14835,N_14584);
or U15421 (N_15421,N_15016,N_15059);
or U15422 (N_15422,N_15180,N_14789);
and U15423 (N_15423,N_15005,N_14999);
nor U15424 (N_15424,N_15092,N_14819);
or U15425 (N_15425,N_14946,N_15186);
nor U15426 (N_15426,N_14435,N_14516);
or U15427 (N_15427,N_14964,N_15028);
or U15428 (N_15428,N_15034,N_14656);
nor U15429 (N_15429,N_14912,N_14528);
and U15430 (N_15430,N_14477,N_14953);
nand U15431 (N_15431,N_14935,N_14544);
nor U15432 (N_15432,N_14524,N_14893);
and U15433 (N_15433,N_14655,N_14461);
or U15434 (N_15434,N_14701,N_15085);
or U15435 (N_15435,N_14740,N_15070);
nor U15436 (N_15436,N_14877,N_14879);
or U15437 (N_15437,N_14834,N_14458);
or U15438 (N_15438,N_14493,N_14763);
and U15439 (N_15439,N_14548,N_14848);
nand U15440 (N_15440,N_14931,N_14950);
nand U15441 (N_15441,N_15197,N_14445);
or U15442 (N_15442,N_14618,N_15006);
or U15443 (N_15443,N_14854,N_14876);
and U15444 (N_15444,N_14704,N_15012);
nand U15445 (N_15445,N_14971,N_14833);
nand U15446 (N_15446,N_14629,N_14486);
nand U15447 (N_15447,N_14853,N_14901);
nand U15448 (N_15448,N_14952,N_14977);
nand U15449 (N_15449,N_15147,N_14457);
nand U15450 (N_15450,N_14930,N_14690);
nor U15451 (N_15451,N_14554,N_14523);
nor U15452 (N_15452,N_14829,N_14844);
or U15453 (N_15453,N_15020,N_14598);
nand U15454 (N_15454,N_14880,N_14491);
and U15455 (N_15455,N_14426,N_14976);
nand U15456 (N_15456,N_14888,N_14866);
and U15457 (N_15457,N_15114,N_14791);
nor U15458 (N_15458,N_14611,N_14787);
and U15459 (N_15459,N_14746,N_14812);
nor U15460 (N_15460,N_15166,N_14886);
or U15461 (N_15461,N_14436,N_15198);
and U15462 (N_15462,N_14566,N_15192);
nand U15463 (N_15463,N_14646,N_15168);
nor U15464 (N_15464,N_14682,N_14583);
nor U15465 (N_15465,N_14525,N_15148);
nor U15466 (N_15466,N_15116,N_14797);
or U15467 (N_15467,N_14858,N_15164);
nand U15468 (N_15468,N_15123,N_14871);
nor U15469 (N_15469,N_14951,N_14699);
or U15470 (N_15470,N_14780,N_14681);
nor U15471 (N_15471,N_15169,N_14451);
and U15472 (N_15472,N_15076,N_15050);
nand U15473 (N_15473,N_14972,N_14439);
nand U15474 (N_15474,N_14526,N_14918);
nand U15475 (N_15475,N_15119,N_15128);
or U15476 (N_15476,N_14919,N_14883);
or U15477 (N_15477,N_14757,N_14739);
and U15478 (N_15478,N_14810,N_14497);
nor U15479 (N_15479,N_14530,N_14800);
and U15480 (N_15480,N_14967,N_15041);
nand U15481 (N_15481,N_14764,N_15019);
and U15482 (N_15482,N_14558,N_14743);
nor U15483 (N_15483,N_15185,N_14689);
nand U15484 (N_15484,N_14447,N_15118);
nor U15485 (N_15485,N_14673,N_15046);
or U15486 (N_15486,N_14921,N_14539);
nand U15487 (N_15487,N_15032,N_14427);
nand U15488 (N_15488,N_14487,N_14571);
nand U15489 (N_15489,N_14695,N_14589);
nand U15490 (N_15490,N_14540,N_14771);
or U15491 (N_15491,N_14957,N_14827);
nand U15492 (N_15492,N_14711,N_14624);
and U15493 (N_15493,N_14406,N_14416);
nand U15494 (N_15494,N_15156,N_14786);
and U15495 (N_15495,N_15117,N_14874);
nand U15496 (N_15496,N_15027,N_14861);
nor U15497 (N_15497,N_14906,N_14697);
nor U15498 (N_15498,N_15144,N_14960);
nor U15499 (N_15499,N_14828,N_15097);
nand U15500 (N_15500,N_14816,N_14694);
or U15501 (N_15501,N_14475,N_14460);
nor U15502 (N_15502,N_14991,N_14452);
and U15503 (N_15503,N_15143,N_14549);
nand U15504 (N_15504,N_14978,N_14772);
nand U15505 (N_15505,N_14506,N_14669);
nor U15506 (N_15506,N_14408,N_14670);
nand U15507 (N_15507,N_14936,N_14562);
nand U15508 (N_15508,N_15163,N_14793);
nor U15509 (N_15509,N_15173,N_14545);
or U15510 (N_15510,N_14433,N_14761);
nand U15511 (N_15511,N_15048,N_15031);
nand U15512 (N_15512,N_14811,N_14958);
and U15513 (N_15513,N_14644,N_14437);
and U15514 (N_15514,N_14884,N_14840);
or U15515 (N_15515,N_14412,N_14628);
and U15516 (N_15516,N_14601,N_15127);
and U15517 (N_15517,N_15154,N_14677);
nand U15518 (N_15518,N_14650,N_15111);
nor U15519 (N_15519,N_14499,N_14759);
or U15520 (N_15520,N_14842,N_14531);
and U15521 (N_15521,N_14407,N_14468);
and U15522 (N_15522,N_15107,N_15011);
or U15523 (N_15523,N_14489,N_14849);
or U15524 (N_15524,N_15181,N_14799);
nand U15525 (N_15525,N_15014,N_14855);
or U15526 (N_15526,N_15199,N_14851);
nand U15527 (N_15527,N_15096,N_14474);
and U15528 (N_15528,N_14507,N_14708);
nand U15529 (N_15529,N_15150,N_14509);
and U15530 (N_15530,N_14941,N_15122);
or U15531 (N_15531,N_14667,N_14556);
nor U15532 (N_15532,N_14843,N_15098);
nand U15533 (N_15533,N_14617,N_14897);
nand U15534 (N_15534,N_15094,N_14666);
nand U15535 (N_15535,N_14635,N_15131);
nor U15536 (N_15536,N_14900,N_15160);
nor U15537 (N_15537,N_15065,N_14570);
and U15538 (N_15538,N_14610,N_14413);
nand U15539 (N_15539,N_14597,N_14622);
nor U15540 (N_15540,N_15133,N_15129);
or U15541 (N_15541,N_14424,N_15009);
nand U15542 (N_15542,N_15149,N_14453);
nor U15543 (N_15543,N_14627,N_14686);
nor U15544 (N_15544,N_14581,N_14926);
or U15545 (N_15545,N_15089,N_14783);
nor U15546 (N_15546,N_15171,N_14665);
or U15547 (N_15547,N_14680,N_14745);
or U15548 (N_15548,N_15142,N_15069);
or U15549 (N_15549,N_14464,N_14742);
nand U15550 (N_15550,N_14604,N_14488);
and U15551 (N_15551,N_15113,N_14788);
and U15552 (N_15552,N_14659,N_15126);
and U15553 (N_15553,N_14619,N_15080);
nand U15554 (N_15554,N_14455,N_15145);
and U15555 (N_15555,N_14794,N_14979);
nor U15556 (N_15556,N_15158,N_14575);
nor U15557 (N_15557,N_14795,N_14984);
or U15558 (N_15558,N_14823,N_15010);
nor U15559 (N_15559,N_15182,N_15045);
and U15560 (N_15560,N_14929,N_14895);
and U15561 (N_15561,N_15091,N_14409);
and U15562 (N_15562,N_14685,N_15038);
nor U15563 (N_15563,N_14747,N_14802);
nor U15564 (N_15564,N_14609,N_14662);
nand U15565 (N_15565,N_14773,N_14410);
or U15566 (N_15566,N_14729,N_14404);
nand U15567 (N_15567,N_14713,N_15162);
nand U15568 (N_15568,N_15174,N_14533);
nand U15569 (N_15569,N_15029,N_14651);
nor U15570 (N_15570,N_14674,N_14927);
nor U15571 (N_15571,N_14401,N_15058);
nand U15572 (N_15572,N_14532,N_15178);
and U15573 (N_15573,N_14717,N_14630);
nand U15574 (N_15574,N_15170,N_14586);
and U15575 (N_15575,N_15146,N_14768);
and U15576 (N_15576,N_14654,N_14721);
nand U15577 (N_15577,N_14814,N_15086);
nor U15578 (N_15578,N_15155,N_14429);
and U15579 (N_15579,N_14448,N_14592);
nand U15580 (N_15580,N_14550,N_15049);
or U15581 (N_15581,N_14937,N_14997);
and U15582 (N_15582,N_15056,N_14872);
and U15583 (N_15583,N_14940,N_14731);
nor U15584 (N_15584,N_14809,N_15105);
nand U15585 (N_15585,N_14887,N_14847);
nor U15586 (N_15586,N_14663,N_14421);
and U15587 (N_15587,N_15013,N_14801);
or U15588 (N_15588,N_14576,N_14945);
and U15589 (N_15589,N_14860,N_14484);
nor U15590 (N_15590,N_14553,N_14716);
nand U15591 (N_15591,N_14784,N_15087);
and U15592 (N_15592,N_15054,N_14857);
nor U15593 (N_15593,N_14511,N_14832);
or U15594 (N_15594,N_14730,N_14614);
or U15595 (N_15595,N_14734,N_14781);
or U15596 (N_15596,N_14846,N_14726);
nor U15597 (N_15597,N_15161,N_14923);
and U15598 (N_15598,N_14479,N_15033);
and U15599 (N_15599,N_14755,N_14580);
and U15600 (N_15600,N_14822,N_14433);
and U15601 (N_15601,N_14958,N_15070);
nand U15602 (N_15602,N_14969,N_14453);
nand U15603 (N_15603,N_15178,N_14491);
nor U15604 (N_15604,N_14941,N_14994);
nand U15605 (N_15605,N_14401,N_14565);
and U15606 (N_15606,N_14711,N_14419);
nand U15607 (N_15607,N_14677,N_14894);
and U15608 (N_15608,N_14779,N_14674);
nand U15609 (N_15609,N_15080,N_15105);
nand U15610 (N_15610,N_14988,N_14724);
nor U15611 (N_15611,N_14401,N_15123);
nand U15612 (N_15612,N_15044,N_14647);
nand U15613 (N_15613,N_15067,N_14495);
or U15614 (N_15614,N_14756,N_14554);
and U15615 (N_15615,N_14539,N_15130);
or U15616 (N_15616,N_14448,N_14717);
or U15617 (N_15617,N_15097,N_14530);
nor U15618 (N_15618,N_14966,N_14958);
nand U15619 (N_15619,N_14534,N_14834);
nand U15620 (N_15620,N_15103,N_15195);
or U15621 (N_15621,N_15039,N_14835);
nor U15622 (N_15622,N_14785,N_14407);
or U15623 (N_15623,N_14623,N_14786);
or U15624 (N_15624,N_14697,N_14445);
nor U15625 (N_15625,N_14989,N_14737);
or U15626 (N_15626,N_14853,N_14764);
nand U15627 (N_15627,N_14796,N_14459);
or U15628 (N_15628,N_14929,N_14539);
and U15629 (N_15629,N_14638,N_14802);
and U15630 (N_15630,N_14772,N_15111);
nand U15631 (N_15631,N_14797,N_15040);
or U15632 (N_15632,N_14941,N_14503);
and U15633 (N_15633,N_14764,N_14861);
nand U15634 (N_15634,N_14615,N_14628);
nor U15635 (N_15635,N_14625,N_15037);
or U15636 (N_15636,N_14860,N_14921);
nand U15637 (N_15637,N_14832,N_14587);
or U15638 (N_15638,N_14842,N_14818);
or U15639 (N_15639,N_15177,N_14485);
and U15640 (N_15640,N_14726,N_14679);
nand U15641 (N_15641,N_15192,N_14632);
nand U15642 (N_15642,N_14812,N_14792);
nor U15643 (N_15643,N_14488,N_14663);
or U15644 (N_15644,N_15162,N_14714);
nor U15645 (N_15645,N_14848,N_14946);
nor U15646 (N_15646,N_14887,N_14458);
and U15647 (N_15647,N_15042,N_15029);
nor U15648 (N_15648,N_15136,N_14434);
or U15649 (N_15649,N_15161,N_14591);
or U15650 (N_15650,N_14401,N_14615);
or U15651 (N_15651,N_14628,N_14577);
or U15652 (N_15652,N_15036,N_14996);
nand U15653 (N_15653,N_14418,N_15153);
or U15654 (N_15654,N_15032,N_14474);
or U15655 (N_15655,N_14882,N_14894);
and U15656 (N_15656,N_14425,N_14924);
and U15657 (N_15657,N_14737,N_14508);
or U15658 (N_15658,N_14592,N_15060);
nand U15659 (N_15659,N_14767,N_15021);
nor U15660 (N_15660,N_14408,N_14756);
nand U15661 (N_15661,N_15128,N_15166);
or U15662 (N_15662,N_14473,N_14909);
xnor U15663 (N_15663,N_15092,N_14910);
and U15664 (N_15664,N_14593,N_14632);
nor U15665 (N_15665,N_14546,N_14451);
nor U15666 (N_15666,N_14675,N_14948);
or U15667 (N_15667,N_14559,N_15132);
or U15668 (N_15668,N_14564,N_14843);
and U15669 (N_15669,N_14633,N_15026);
or U15670 (N_15670,N_14411,N_14795);
or U15671 (N_15671,N_14534,N_14428);
nand U15672 (N_15672,N_14451,N_14507);
and U15673 (N_15673,N_14807,N_14437);
nand U15674 (N_15674,N_14755,N_14912);
nand U15675 (N_15675,N_14679,N_15193);
nor U15676 (N_15676,N_15029,N_15126);
nand U15677 (N_15677,N_14659,N_14525);
or U15678 (N_15678,N_15057,N_14980);
or U15679 (N_15679,N_14747,N_15088);
or U15680 (N_15680,N_14691,N_14971);
and U15681 (N_15681,N_14488,N_14932);
nand U15682 (N_15682,N_14947,N_14813);
nor U15683 (N_15683,N_14919,N_14633);
nor U15684 (N_15684,N_14816,N_15166);
or U15685 (N_15685,N_15075,N_14651);
and U15686 (N_15686,N_14561,N_14450);
nor U15687 (N_15687,N_14648,N_14485);
nor U15688 (N_15688,N_14701,N_14531);
nor U15689 (N_15689,N_14727,N_14868);
or U15690 (N_15690,N_14992,N_14704);
nor U15691 (N_15691,N_14694,N_14855);
or U15692 (N_15692,N_14507,N_15156);
or U15693 (N_15693,N_14891,N_14639);
nor U15694 (N_15694,N_15106,N_14510);
and U15695 (N_15695,N_15053,N_14853);
nor U15696 (N_15696,N_15034,N_14542);
or U15697 (N_15697,N_14701,N_14418);
or U15698 (N_15698,N_15008,N_14652);
and U15699 (N_15699,N_14933,N_14827);
and U15700 (N_15700,N_15079,N_14439);
nor U15701 (N_15701,N_15199,N_14924);
or U15702 (N_15702,N_14523,N_15023);
and U15703 (N_15703,N_14434,N_15195);
nand U15704 (N_15704,N_14455,N_14482);
nor U15705 (N_15705,N_14699,N_14636);
or U15706 (N_15706,N_14668,N_15133);
or U15707 (N_15707,N_14500,N_14437);
and U15708 (N_15708,N_15007,N_14642);
or U15709 (N_15709,N_14819,N_14646);
nand U15710 (N_15710,N_14845,N_14971);
nand U15711 (N_15711,N_14993,N_14414);
and U15712 (N_15712,N_14877,N_15013);
nor U15713 (N_15713,N_15185,N_14585);
nor U15714 (N_15714,N_14517,N_14886);
or U15715 (N_15715,N_15104,N_14813);
or U15716 (N_15716,N_14746,N_14634);
or U15717 (N_15717,N_14691,N_14588);
and U15718 (N_15718,N_14653,N_14958);
or U15719 (N_15719,N_14747,N_14637);
or U15720 (N_15720,N_15166,N_14529);
or U15721 (N_15721,N_14914,N_14906);
and U15722 (N_15722,N_14968,N_15074);
or U15723 (N_15723,N_14783,N_15125);
nand U15724 (N_15724,N_14484,N_15128);
nor U15725 (N_15725,N_14440,N_14483);
nor U15726 (N_15726,N_15089,N_14571);
or U15727 (N_15727,N_14690,N_14870);
or U15728 (N_15728,N_14646,N_14814);
nand U15729 (N_15729,N_14527,N_14674);
and U15730 (N_15730,N_14904,N_14535);
or U15731 (N_15731,N_14573,N_14969);
and U15732 (N_15732,N_14477,N_14684);
nor U15733 (N_15733,N_15045,N_14451);
nor U15734 (N_15734,N_14614,N_14566);
xor U15735 (N_15735,N_14682,N_15039);
and U15736 (N_15736,N_14547,N_14458);
nand U15737 (N_15737,N_14633,N_14935);
nand U15738 (N_15738,N_14713,N_14801);
and U15739 (N_15739,N_14916,N_14584);
nand U15740 (N_15740,N_15061,N_14943);
nor U15741 (N_15741,N_14765,N_15136);
and U15742 (N_15742,N_14789,N_15168);
nand U15743 (N_15743,N_14693,N_14980);
or U15744 (N_15744,N_14948,N_14635);
nand U15745 (N_15745,N_15081,N_14767);
and U15746 (N_15746,N_14609,N_15087);
and U15747 (N_15747,N_14425,N_14616);
nand U15748 (N_15748,N_14428,N_14680);
and U15749 (N_15749,N_14970,N_14962);
or U15750 (N_15750,N_14845,N_14514);
nor U15751 (N_15751,N_14871,N_14728);
or U15752 (N_15752,N_14836,N_14883);
and U15753 (N_15753,N_15077,N_14640);
or U15754 (N_15754,N_15040,N_14967);
and U15755 (N_15755,N_14465,N_14894);
nand U15756 (N_15756,N_14893,N_14859);
nor U15757 (N_15757,N_14985,N_14673);
nor U15758 (N_15758,N_14625,N_14509);
nand U15759 (N_15759,N_14601,N_15099);
or U15760 (N_15760,N_14731,N_14554);
or U15761 (N_15761,N_14476,N_15032);
nor U15762 (N_15762,N_14950,N_14546);
xnor U15763 (N_15763,N_14837,N_15010);
and U15764 (N_15764,N_14742,N_14954);
and U15765 (N_15765,N_14452,N_14411);
nand U15766 (N_15766,N_14728,N_14714);
and U15767 (N_15767,N_14443,N_14878);
and U15768 (N_15768,N_15168,N_14634);
nor U15769 (N_15769,N_14643,N_14873);
and U15770 (N_15770,N_14452,N_14509);
and U15771 (N_15771,N_15108,N_14819);
nor U15772 (N_15772,N_15009,N_14449);
nand U15773 (N_15773,N_14943,N_15157);
nand U15774 (N_15774,N_15000,N_14984);
or U15775 (N_15775,N_14883,N_15080);
nand U15776 (N_15776,N_14481,N_14815);
and U15777 (N_15777,N_14743,N_15168);
nor U15778 (N_15778,N_14866,N_14750);
or U15779 (N_15779,N_14906,N_15082);
or U15780 (N_15780,N_14492,N_14847);
and U15781 (N_15781,N_14619,N_14864);
or U15782 (N_15782,N_14977,N_14773);
or U15783 (N_15783,N_14868,N_14944);
nor U15784 (N_15784,N_14990,N_14974);
nand U15785 (N_15785,N_15151,N_14490);
nand U15786 (N_15786,N_14850,N_14557);
nor U15787 (N_15787,N_14950,N_14697);
or U15788 (N_15788,N_14923,N_14746);
nor U15789 (N_15789,N_15028,N_14785);
and U15790 (N_15790,N_14408,N_14652);
nor U15791 (N_15791,N_14861,N_15023);
and U15792 (N_15792,N_14797,N_14487);
nand U15793 (N_15793,N_14502,N_15071);
nor U15794 (N_15794,N_14682,N_14703);
nand U15795 (N_15795,N_15134,N_14795);
nor U15796 (N_15796,N_14492,N_14522);
nand U15797 (N_15797,N_14541,N_14671);
or U15798 (N_15798,N_14547,N_15058);
or U15799 (N_15799,N_14924,N_14609);
or U15800 (N_15800,N_14685,N_14658);
or U15801 (N_15801,N_15190,N_15081);
or U15802 (N_15802,N_14423,N_15003);
and U15803 (N_15803,N_15064,N_15061);
nand U15804 (N_15804,N_15110,N_14592);
nor U15805 (N_15805,N_14936,N_15087);
or U15806 (N_15806,N_14905,N_14870);
and U15807 (N_15807,N_14859,N_15026);
or U15808 (N_15808,N_14779,N_14505);
nand U15809 (N_15809,N_15015,N_14510);
nor U15810 (N_15810,N_15038,N_15134);
and U15811 (N_15811,N_14917,N_15128);
nor U15812 (N_15812,N_14993,N_14673);
nand U15813 (N_15813,N_14978,N_14530);
or U15814 (N_15814,N_14659,N_15084);
or U15815 (N_15815,N_15050,N_14489);
nor U15816 (N_15816,N_14576,N_14440);
and U15817 (N_15817,N_15110,N_14844);
and U15818 (N_15818,N_14970,N_15136);
nor U15819 (N_15819,N_15168,N_14464);
or U15820 (N_15820,N_14441,N_14976);
nand U15821 (N_15821,N_14894,N_15078);
nand U15822 (N_15822,N_15159,N_14845);
nor U15823 (N_15823,N_15068,N_14650);
and U15824 (N_15824,N_14869,N_14553);
nor U15825 (N_15825,N_14596,N_14695);
and U15826 (N_15826,N_15092,N_14673);
and U15827 (N_15827,N_14865,N_15122);
or U15828 (N_15828,N_14987,N_14751);
or U15829 (N_15829,N_14627,N_15082);
nor U15830 (N_15830,N_14997,N_14416);
nor U15831 (N_15831,N_14688,N_14943);
nand U15832 (N_15832,N_15057,N_14809);
and U15833 (N_15833,N_14540,N_14413);
or U15834 (N_15834,N_14879,N_14779);
and U15835 (N_15835,N_14562,N_14827);
nand U15836 (N_15836,N_15184,N_15165);
nor U15837 (N_15837,N_14689,N_14992);
nand U15838 (N_15838,N_14985,N_14814);
and U15839 (N_15839,N_15113,N_14897);
nand U15840 (N_15840,N_14413,N_15105);
and U15841 (N_15841,N_14861,N_14727);
or U15842 (N_15842,N_14510,N_14505);
and U15843 (N_15843,N_14645,N_14856);
nor U15844 (N_15844,N_15169,N_14645);
and U15845 (N_15845,N_14712,N_14648);
nor U15846 (N_15846,N_14908,N_14825);
or U15847 (N_15847,N_15018,N_14981);
nand U15848 (N_15848,N_14673,N_14674);
nand U15849 (N_15849,N_15168,N_14750);
nor U15850 (N_15850,N_14656,N_14630);
nor U15851 (N_15851,N_15095,N_14766);
nor U15852 (N_15852,N_15165,N_14425);
and U15853 (N_15853,N_15153,N_14724);
or U15854 (N_15854,N_15132,N_15198);
and U15855 (N_15855,N_15025,N_14543);
or U15856 (N_15856,N_14989,N_14951);
and U15857 (N_15857,N_14724,N_14502);
and U15858 (N_15858,N_14715,N_15027);
and U15859 (N_15859,N_14551,N_14567);
nor U15860 (N_15860,N_15124,N_14495);
or U15861 (N_15861,N_14727,N_15187);
nand U15862 (N_15862,N_14811,N_15122);
nand U15863 (N_15863,N_14815,N_14456);
and U15864 (N_15864,N_14921,N_14847);
or U15865 (N_15865,N_14585,N_14996);
or U15866 (N_15866,N_14616,N_15182);
and U15867 (N_15867,N_14985,N_14674);
nand U15868 (N_15868,N_14721,N_14884);
nor U15869 (N_15869,N_14824,N_14633);
nor U15870 (N_15870,N_14441,N_14930);
or U15871 (N_15871,N_14531,N_15058);
nand U15872 (N_15872,N_14827,N_14526);
or U15873 (N_15873,N_14615,N_14532);
nand U15874 (N_15874,N_14870,N_15197);
nor U15875 (N_15875,N_14928,N_14799);
and U15876 (N_15876,N_14863,N_14961);
or U15877 (N_15877,N_14779,N_14823);
nand U15878 (N_15878,N_14652,N_15004);
and U15879 (N_15879,N_14714,N_14581);
and U15880 (N_15880,N_15031,N_14997);
nor U15881 (N_15881,N_14685,N_14690);
nor U15882 (N_15882,N_14438,N_15081);
nor U15883 (N_15883,N_14546,N_14831);
nor U15884 (N_15884,N_14427,N_15135);
nor U15885 (N_15885,N_14711,N_15173);
nand U15886 (N_15886,N_15154,N_15129);
nand U15887 (N_15887,N_14477,N_14701);
and U15888 (N_15888,N_15079,N_14479);
nand U15889 (N_15889,N_14742,N_14674);
nor U15890 (N_15890,N_14962,N_15024);
and U15891 (N_15891,N_14461,N_15199);
or U15892 (N_15892,N_14888,N_14572);
nand U15893 (N_15893,N_14453,N_15181);
nor U15894 (N_15894,N_14644,N_15043);
and U15895 (N_15895,N_15045,N_14994);
and U15896 (N_15896,N_15044,N_15088);
or U15897 (N_15897,N_14831,N_14729);
and U15898 (N_15898,N_14862,N_14500);
or U15899 (N_15899,N_14964,N_14949);
and U15900 (N_15900,N_14552,N_14405);
or U15901 (N_15901,N_14431,N_14845);
or U15902 (N_15902,N_15035,N_14559);
nand U15903 (N_15903,N_14982,N_15155);
and U15904 (N_15904,N_14790,N_14882);
or U15905 (N_15905,N_14503,N_14909);
nand U15906 (N_15906,N_15148,N_14739);
or U15907 (N_15907,N_14688,N_14843);
nand U15908 (N_15908,N_14417,N_14709);
nand U15909 (N_15909,N_14513,N_14956);
and U15910 (N_15910,N_14896,N_15038);
nand U15911 (N_15911,N_15114,N_14959);
nor U15912 (N_15912,N_14936,N_15105);
and U15913 (N_15913,N_14597,N_14562);
or U15914 (N_15914,N_15102,N_15191);
nand U15915 (N_15915,N_14453,N_14806);
nor U15916 (N_15916,N_15157,N_14606);
nand U15917 (N_15917,N_14890,N_15181);
and U15918 (N_15918,N_14681,N_14454);
and U15919 (N_15919,N_14935,N_15089);
nand U15920 (N_15920,N_14658,N_14674);
nor U15921 (N_15921,N_14960,N_15104);
or U15922 (N_15922,N_14548,N_14764);
and U15923 (N_15923,N_14968,N_14708);
nand U15924 (N_15924,N_15079,N_14623);
or U15925 (N_15925,N_15087,N_15111);
nand U15926 (N_15926,N_14975,N_14414);
nand U15927 (N_15927,N_14859,N_14553);
nand U15928 (N_15928,N_15035,N_14653);
and U15929 (N_15929,N_14565,N_14494);
and U15930 (N_15930,N_14409,N_14922);
or U15931 (N_15931,N_14602,N_15041);
nor U15932 (N_15932,N_14560,N_14841);
nand U15933 (N_15933,N_14492,N_14932);
or U15934 (N_15934,N_14549,N_14507);
and U15935 (N_15935,N_14956,N_15088);
and U15936 (N_15936,N_14870,N_14484);
or U15937 (N_15937,N_14447,N_15024);
nor U15938 (N_15938,N_14960,N_14635);
or U15939 (N_15939,N_14852,N_14520);
and U15940 (N_15940,N_14978,N_14851);
and U15941 (N_15941,N_14617,N_14703);
and U15942 (N_15942,N_14755,N_14886);
and U15943 (N_15943,N_14774,N_15038);
or U15944 (N_15944,N_14599,N_14936);
nand U15945 (N_15945,N_14805,N_14883);
or U15946 (N_15946,N_15094,N_14694);
nor U15947 (N_15947,N_14760,N_15187);
xnor U15948 (N_15948,N_15039,N_14976);
nor U15949 (N_15949,N_14720,N_15191);
or U15950 (N_15950,N_15039,N_14772);
or U15951 (N_15951,N_14843,N_14718);
or U15952 (N_15952,N_14859,N_15092);
nand U15953 (N_15953,N_14870,N_15022);
nor U15954 (N_15954,N_14433,N_14599);
nor U15955 (N_15955,N_14514,N_14988);
nand U15956 (N_15956,N_15051,N_14683);
nor U15957 (N_15957,N_14752,N_14949);
nor U15958 (N_15958,N_14801,N_14756);
or U15959 (N_15959,N_14415,N_14691);
nand U15960 (N_15960,N_14698,N_15047);
and U15961 (N_15961,N_14553,N_14717);
and U15962 (N_15962,N_15179,N_14456);
or U15963 (N_15963,N_14853,N_14526);
and U15964 (N_15964,N_15010,N_15034);
and U15965 (N_15965,N_14814,N_15179);
nor U15966 (N_15966,N_15163,N_15119);
nor U15967 (N_15967,N_14847,N_14507);
nor U15968 (N_15968,N_14490,N_15012);
nand U15969 (N_15969,N_15197,N_15180);
and U15970 (N_15970,N_15159,N_15147);
or U15971 (N_15971,N_15084,N_14525);
nand U15972 (N_15972,N_14585,N_14918);
nor U15973 (N_15973,N_14697,N_15161);
nor U15974 (N_15974,N_14464,N_14460);
nand U15975 (N_15975,N_14850,N_14955);
nand U15976 (N_15976,N_14585,N_14859);
and U15977 (N_15977,N_14429,N_15009);
nand U15978 (N_15978,N_14438,N_14852);
nand U15979 (N_15979,N_14749,N_14527);
nand U15980 (N_15980,N_14954,N_14824);
and U15981 (N_15981,N_14652,N_14747);
xor U15982 (N_15982,N_14732,N_14455);
nand U15983 (N_15983,N_15121,N_14576);
and U15984 (N_15984,N_14906,N_14602);
nor U15985 (N_15985,N_14879,N_14863);
nor U15986 (N_15986,N_15055,N_14527);
nand U15987 (N_15987,N_14443,N_14730);
nor U15988 (N_15988,N_14714,N_14448);
or U15989 (N_15989,N_14605,N_14926);
and U15990 (N_15990,N_14751,N_14446);
or U15991 (N_15991,N_15127,N_14479);
or U15992 (N_15992,N_14894,N_14892);
and U15993 (N_15993,N_15020,N_14775);
or U15994 (N_15994,N_14688,N_15062);
and U15995 (N_15995,N_14816,N_15107);
and U15996 (N_15996,N_14465,N_14854);
or U15997 (N_15997,N_14589,N_15084);
nor U15998 (N_15998,N_14533,N_14949);
and U15999 (N_15999,N_14851,N_15114);
and U16000 (N_16000,N_15520,N_15701);
and U16001 (N_16001,N_15274,N_15319);
nand U16002 (N_16002,N_15236,N_15551);
or U16003 (N_16003,N_15597,N_15289);
and U16004 (N_16004,N_15860,N_15892);
nand U16005 (N_16005,N_15910,N_15834);
or U16006 (N_16006,N_15502,N_15880);
nor U16007 (N_16007,N_15667,N_15848);
nor U16008 (N_16008,N_15463,N_15496);
xnor U16009 (N_16009,N_15385,N_15991);
or U16010 (N_16010,N_15664,N_15838);
nor U16011 (N_16011,N_15392,N_15321);
and U16012 (N_16012,N_15317,N_15789);
nor U16013 (N_16013,N_15883,N_15347);
nor U16014 (N_16014,N_15654,N_15921);
and U16015 (N_16015,N_15332,N_15453);
nand U16016 (N_16016,N_15526,N_15490);
nand U16017 (N_16017,N_15420,N_15872);
and U16018 (N_16018,N_15300,N_15607);
or U16019 (N_16019,N_15975,N_15574);
nand U16020 (N_16020,N_15955,N_15229);
xor U16021 (N_16021,N_15686,N_15590);
nor U16022 (N_16022,N_15690,N_15458);
nor U16023 (N_16023,N_15234,N_15292);
or U16024 (N_16024,N_15823,N_15613);
or U16025 (N_16025,N_15889,N_15969);
nor U16026 (N_16026,N_15312,N_15800);
and U16027 (N_16027,N_15916,N_15581);
or U16028 (N_16028,N_15986,N_15459);
and U16029 (N_16029,N_15753,N_15330);
or U16030 (N_16030,N_15402,N_15573);
or U16031 (N_16031,N_15617,N_15666);
or U16032 (N_16032,N_15736,N_15863);
or U16033 (N_16033,N_15315,N_15530);
and U16034 (N_16034,N_15318,N_15498);
nor U16035 (N_16035,N_15412,N_15846);
nor U16036 (N_16036,N_15564,N_15596);
or U16037 (N_16037,N_15480,N_15956);
nand U16038 (N_16038,N_15235,N_15741);
and U16039 (N_16039,N_15216,N_15288);
nor U16040 (N_16040,N_15746,N_15757);
or U16041 (N_16041,N_15772,N_15454);
nor U16042 (N_16042,N_15905,N_15250);
or U16043 (N_16043,N_15864,N_15541);
and U16044 (N_16044,N_15255,N_15243);
and U16045 (N_16045,N_15219,N_15637);
nand U16046 (N_16046,N_15380,N_15728);
and U16047 (N_16047,N_15710,N_15427);
nand U16048 (N_16048,N_15777,N_15430);
nand U16049 (N_16049,N_15951,N_15485);
and U16050 (N_16050,N_15529,N_15985);
nor U16051 (N_16051,N_15922,N_15796);
and U16052 (N_16052,N_15875,N_15499);
nor U16053 (N_16053,N_15363,N_15466);
or U16054 (N_16054,N_15641,N_15578);
or U16055 (N_16055,N_15351,N_15546);
and U16056 (N_16056,N_15553,N_15394);
nand U16057 (N_16057,N_15675,N_15437);
and U16058 (N_16058,N_15791,N_15333);
nor U16059 (N_16059,N_15718,N_15349);
nand U16060 (N_16060,N_15859,N_15781);
or U16061 (N_16061,N_15784,N_15649);
or U16062 (N_16062,N_15805,N_15411);
and U16063 (N_16063,N_15543,N_15409);
nand U16064 (N_16064,N_15750,N_15388);
and U16065 (N_16065,N_15215,N_15565);
and U16066 (N_16066,N_15579,N_15837);
nor U16067 (N_16067,N_15395,N_15900);
or U16068 (N_16068,N_15888,N_15920);
and U16069 (N_16069,N_15345,N_15893);
nor U16070 (N_16070,N_15524,N_15803);
nor U16071 (N_16071,N_15595,N_15337);
or U16072 (N_16072,N_15311,N_15704);
and U16073 (N_16073,N_15301,N_15972);
nor U16074 (N_16074,N_15493,N_15720);
nor U16075 (N_16075,N_15907,N_15536);
or U16076 (N_16076,N_15958,N_15810);
or U16077 (N_16077,N_15782,N_15850);
or U16078 (N_16078,N_15712,N_15685);
or U16079 (N_16079,N_15725,N_15677);
and U16080 (N_16080,N_15627,N_15625);
nor U16081 (N_16081,N_15906,N_15523);
or U16082 (N_16082,N_15545,N_15946);
and U16083 (N_16083,N_15995,N_15731);
or U16084 (N_16084,N_15623,N_15534);
or U16085 (N_16085,N_15949,N_15687);
and U16086 (N_16086,N_15276,N_15818);
nor U16087 (N_16087,N_15362,N_15861);
nor U16088 (N_16088,N_15372,N_15811);
nor U16089 (N_16089,N_15689,N_15851);
or U16090 (N_16090,N_15809,N_15778);
nor U16091 (N_16091,N_15299,N_15447);
or U16092 (N_16092,N_15483,N_15615);
or U16093 (N_16093,N_15239,N_15223);
or U16094 (N_16094,N_15305,N_15929);
or U16095 (N_16095,N_15976,N_15397);
or U16096 (N_16096,N_15484,N_15729);
nand U16097 (N_16097,N_15714,N_15220);
and U16098 (N_16098,N_15237,N_15918);
and U16099 (N_16099,N_15267,N_15455);
nand U16100 (N_16100,N_15924,N_15899);
or U16101 (N_16101,N_15342,N_15793);
or U16102 (N_16102,N_15228,N_15282);
nand U16103 (N_16103,N_15503,N_15592);
and U16104 (N_16104,N_15399,N_15703);
and U16105 (N_16105,N_15618,N_15540);
nand U16106 (N_16106,N_15797,N_15568);
or U16107 (N_16107,N_15877,N_15304);
nor U16108 (N_16108,N_15417,N_15759);
and U16109 (N_16109,N_15711,N_15908);
and U16110 (N_16110,N_15205,N_15435);
or U16111 (N_16111,N_15962,N_15386);
and U16112 (N_16112,N_15843,N_15383);
or U16113 (N_16113,N_15896,N_15914);
or U16114 (N_16114,N_15936,N_15754);
nand U16115 (N_16115,N_15683,N_15945);
nand U16116 (N_16116,N_15230,N_15659);
nor U16117 (N_16117,N_15436,N_15602);
nand U16118 (N_16118,N_15381,N_15488);
xor U16119 (N_16119,N_15290,N_15751);
and U16120 (N_16120,N_15295,N_15462);
and U16121 (N_16121,N_15773,N_15377);
or U16122 (N_16122,N_15978,N_15240);
nand U16123 (N_16123,N_15375,N_15531);
nor U16124 (N_16124,N_15770,N_15213);
or U16125 (N_16125,N_15702,N_15355);
and U16126 (N_16126,N_15482,N_15248);
nor U16127 (N_16127,N_15933,N_15376);
or U16128 (N_16128,N_15519,N_15218);
nor U16129 (N_16129,N_15616,N_15422);
and U16130 (N_16130,N_15472,N_15280);
and U16131 (N_16131,N_15525,N_15365);
and U16132 (N_16132,N_15768,N_15651);
nor U16133 (N_16133,N_15259,N_15960);
nor U16134 (N_16134,N_15571,N_15478);
nor U16135 (N_16135,N_15238,N_15890);
nor U16136 (N_16136,N_15293,N_15698);
or U16137 (N_16137,N_15373,N_15360);
or U16138 (N_16138,N_15987,N_15650);
or U16139 (N_16139,N_15585,N_15981);
nor U16140 (N_16140,N_15895,N_15854);
nor U16141 (N_16141,N_15604,N_15210);
nand U16142 (N_16142,N_15467,N_15494);
and U16143 (N_16143,N_15507,N_15994);
nand U16144 (N_16144,N_15857,N_15973);
nand U16145 (N_16145,N_15721,N_15771);
nor U16146 (N_16146,N_15856,N_15790);
nor U16147 (N_16147,N_15628,N_15251);
nor U16148 (N_16148,N_15971,N_15737);
nand U16149 (N_16149,N_15652,N_15325);
and U16150 (N_16150,N_15302,N_15416);
nor U16151 (N_16151,N_15217,N_15897);
nand U16152 (N_16152,N_15456,N_15272);
and U16153 (N_16153,N_15434,N_15776);
nand U16154 (N_16154,N_15513,N_15634);
nor U16155 (N_16155,N_15879,N_15461);
or U16156 (N_16156,N_15418,N_15947);
nor U16157 (N_16157,N_15682,N_15886);
nor U16158 (N_16158,N_15479,N_15569);
and U16159 (N_16159,N_15726,N_15799);
and U16160 (N_16160,N_15727,N_15323);
and U16161 (N_16161,N_15827,N_15369);
nor U16162 (N_16162,N_15817,N_15473);
nor U16163 (N_16163,N_15780,N_15779);
nor U16164 (N_16164,N_15925,N_15887);
and U16165 (N_16165,N_15999,N_15764);
and U16166 (N_16166,N_15849,N_15491);
nand U16167 (N_16167,N_15277,N_15979);
or U16168 (N_16168,N_15841,N_15425);
nor U16169 (N_16169,N_15669,N_15765);
and U16170 (N_16170,N_15593,N_15405);
nor U16171 (N_16171,N_15752,N_15917);
or U16172 (N_16172,N_15357,N_15928);
nand U16173 (N_16173,N_15258,N_15723);
and U16174 (N_16174,N_15705,N_15224);
and U16175 (N_16175,N_15672,N_15242);
nand U16176 (N_16176,N_15716,N_15644);
nand U16177 (N_16177,N_15855,N_15885);
and U16178 (N_16178,N_15819,N_15443);
and U16179 (N_16179,N_15265,N_15606);
or U16180 (N_16180,N_15839,N_15594);
nand U16181 (N_16181,N_15948,N_15264);
nor U16182 (N_16182,N_15655,N_15661);
nand U16183 (N_16183,N_15798,N_15582);
xor U16184 (N_16184,N_15967,N_15694);
or U16185 (N_16185,N_15440,N_15474);
nand U16186 (N_16186,N_15983,N_15774);
or U16187 (N_16187,N_15927,N_15470);
and U16188 (N_16188,N_15953,N_15642);
nand U16189 (N_16189,N_15679,N_15533);
nor U16190 (N_16190,N_15674,N_15204);
or U16191 (N_16191,N_15518,N_15510);
and U16192 (N_16192,N_15471,N_15477);
and U16193 (N_16193,N_15400,N_15214);
and U16194 (N_16194,N_15423,N_15743);
nand U16195 (N_16195,N_15469,N_15329);
nor U16196 (N_16196,N_15419,N_15283);
or U16197 (N_16197,N_15629,N_15867);
or U16198 (N_16198,N_15207,N_15268);
and U16199 (N_16199,N_15598,N_15465);
or U16200 (N_16200,N_15206,N_15424);
or U16201 (N_16201,N_15308,N_15665);
nand U16202 (N_16202,N_15869,N_15403);
nand U16203 (N_16203,N_15339,N_15586);
nor U16204 (N_16204,N_15306,N_15605);
and U16205 (N_16205,N_15662,N_15587);
and U16206 (N_16206,N_15278,N_15847);
nand U16207 (N_16207,N_15415,N_15610);
or U16208 (N_16208,N_15824,N_15309);
nand U16209 (N_16209,N_15515,N_15816);
and U16210 (N_16210,N_15445,N_15387);
or U16211 (N_16211,N_15747,N_15733);
nor U16212 (N_16212,N_15912,N_15954);
or U16213 (N_16213,N_15648,N_15919);
and U16214 (N_16214,N_15835,N_15639);
nor U16215 (N_16215,N_15748,N_15670);
nor U16216 (N_16216,N_15366,N_15556);
nand U16217 (N_16217,N_15766,N_15575);
nand U16218 (N_16218,N_15433,N_15338);
nand U16219 (N_16219,N_15275,N_15744);
nand U16220 (N_16220,N_15451,N_15930);
and U16221 (N_16221,N_15539,N_15364);
nand U16222 (N_16222,N_15614,N_15944);
or U16223 (N_16223,N_15635,N_15547);
or U16224 (N_16224,N_15426,N_15506);
nand U16225 (N_16225,N_15512,N_15732);
and U16226 (N_16226,N_15550,N_15915);
or U16227 (N_16227,N_15671,N_15787);
and U16228 (N_16228,N_15699,N_15891);
and U16229 (N_16229,N_15783,N_15911);
nand U16230 (N_16230,N_15350,N_15331);
nor U16231 (N_16231,N_15609,N_15566);
nor U16232 (N_16232,N_15840,N_15990);
and U16233 (N_16233,N_15697,N_15996);
nor U16234 (N_16234,N_15865,N_15576);
and U16235 (N_16235,N_15830,N_15354);
or U16236 (N_16236,N_15314,N_15821);
and U16237 (N_16237,N_15882,N_15624);
nand U16238 (N_16238,N_15583,N_15619);
nand U16239 (N_16239,N_15923,N_15769);
nand U16240 (N_16240,N_15495,N_15442);
and U16241 (N_16241,N_15486,N_15457);
or U16242 (N_16242,N_15735,N_15942);
nor U16243 (N_16243,N_15233,N_15438);
or U16244 (N_16244,N_15562,N_15646);
nor U16245 (N_16245,N_15208,N_15707);
or U16246 (N_16246,N_15804,N_15468);
nor U16247 (N_16247,N_15501,N_15678);
and U16248 (N_16248,N_15358,N_15656);
nor U16249 (N_16249,N_15414,N_15448);
nor U16250 (N_16250,N_15352,N_15738);
nand U16251 (N_16251,N_15421,N_15952);
and U16252 (N_16252,N_15998,N_15441);
and U16253 (N_16253,N_15831,N_15226);
or U16254 (N_16254,N_15298,N_15633);
and U16255 (N_16255,N_15505,N_15511);
or U16256 (N_16256,N_15684,N_15970);
or U16257 (N_16257,N_15313,N_15901);
or U16258 (N_16258,N_15866,N_15262);
or U16259 (N_16259,N_15935,N_15601);
and U16260 (N_16260,N_15695,N_15567);
or U16261 (N_16261,N_15252,N_15977);
nand U16262 (N_16262,N_15706,N_15842);
nand U16263 (N_16263,N_15761,N_15367);
nor U16264 (N_16264,N_15621,N_15563);
nand U16265 (N_16265,N_15795,N_15868);
nand U16266 (N_16266,N_15446,N_15963);
nand U16267 (N_16267,N_15432,N_15813);
and U16268 (N_16268,N_15227,N_15269);
nor U16269 (N_16269,N_15584,N_15989);
nor U16270 (N_16270,N_15965,N_15500);
nand U16271 (N_16271,N_15904,N_15320);
nor U16272 (N_16272,N_15257,N_15961);
nand U16273 (N_16273,N_15808,N_15361);
or U16274 (N_16274,N_15263,N_15353);
nand U16275 (N_16275,N_15926,N_15786);
nor U16276 (N_16276,N_15212,N_15241);
nor U16277 (N_16277,N_15871,N_15833);
or U16278 (N_16278,N_15222,N_15335);
and U16279 (N_16279,N_15504,N_15755);
nand U16280 (N_16280,N_15608,N_15807);
or U16281 (N_16281,N_15244,N_15984);
or U16282 (N_16282,N_15231,N_15591);
nor U16283 (N_16283,N_15481,N_15407);
nor U16284 (N_16284,N_15340,N_15806);
nand U16285 (N_16285,N_15246,N_15862);
nand U16286 (N_16286,N_15371,N_15344);
nor U16287 (N_16287,N_15284,N_15894);
and U16288 (N_16288,N_15663,N_15202);
nor U16289 (N_16289,N_15555,N_15476);
nor U16290 (N_16290,N_15626,N_15832);
and U16291 (N_16291,N_15374,N_15647);
nor U16292 (N_16292,N_15903,N_15898);
nor U16293 (N_16293,N_15802,N_15941);
and U16294 (N_16294,N_15561,N_15742);
nand U16295 (N_16295,N_15393,N_15508);
nand U16296 (N_16296,N_15988,N_15291);
nor U16297 (N_16297,N_15668,N_15296);
nor U16298 (N_16298,N_15964,N_15792);
or U16299 (N_16299,N_15532,N_15396);
or U16300 (N_16300,N_15696,N_15836);
or U16301 (N_16301,N_15391,N_15700);
nor U16302 (N_16302,N_15788,N_15909);
nor U16303 (N_16303,N_15286,N_15611);
and U16304 (N_16304,N_15548,N_15521);
nand U16305 (N_16305,N_15825,N_15401);
or U16306 (N_16306,N_15870,N_15558);
or U16307 (N_16307,N_15815,N_15572);
nor U16308 (N_16308,N_15559,N_15509);
nand U16309 (N_16309,N_15211,N_15873);
nand U16310 (N_16310,N_15640,N_15968);
nand U16311 (N_16311,N_15516,N_15537);
xnor U16312 (N_16312,N_15767,N_15260);
nor U16313 (N_16313,N_15724,N_15858);
or U16314 (N_16314,N_15636,N_15620);
nand U16315 (N_16315,N_15382,N_15577);
and U16316 (N_16316,N_15599,N_15356);
and U16317 (N_16317,N_15271,N_15938);
and U16318 (N_16318,N_15785,N_15939);
and U16319 (N_16319,N_15874,N_15913);
xor U16320 (N_16320,N_15643,N_15359);
nand U16321 (N_16321,N_15535,N_15389);
nand U16322 (N_16322,N_15822,N_15254);
nand U16323 (N_16323,N_15232,N_15801);
nor U16324 (N_16324,N_15343,N_15326);
and U16325 (N_16325,N_15273,N_15570);
nor U16326 (N_16326,N_15221,N_15514);
and U16327 (N_16327,N_15413,N_15630);
nor U16328 (N_16328,N_15209,N_15876);
and U16329 (N_16329,N_15464,N_15631);
nor U16330 (N_16330,N_15982,N_15980);
xor U16331 (N_16331,N_15554,N_15406);
and U16332 (N_16332,N_15253,N_15398);
nor U16333 (N_16333,N_15730,N_15557);
nor U16334 (N_16334,N_15688,N_15829);
nor U16335 (N_16335,N_15449,N_15522);
nand U16336 (N_16336,N_15845,N_15814);
nand U16337 (N_16337,N_15713,N_15297);
or U16338 (N_16338,N_15294,N_15739);
or U16339 (N_16339,N_15487,N_15715);
and U16340 (N_16340,N_15997,N_15327);
or U16341 (N_16341,N_15826,N_15762);
or U16342 (N_16342,N_15680,N_15932);
nor U16343 (N_16343,N_15950,N_15307);
nor U16344 (N_16344,N_15722,N_15256);
and U16345 (N_16345,N_15603,N_15937);
and U16346 (N_16346,N_15316,N_15303);
and U16347 (N_16347,N_15709,N_15622);
and U16348 (N_16348,N_15660,N_15760);
and U16349 (N_16349,N_15341,N_15681);
nor U16350 (N_16350,N_15589,N_15653);
nor U16351 (N_16351,N_15600,N_15287);
and U16352 (N_16352,N_15475,N_15719);
xnor U16353 (N_16353,N_15517,N_15708);
nand U16354 (N_16354,N_15245,N_15612);
nand U16355 (N_16355,N_15758,N_15756);
and U16356 (N_16356,N_15200,N_15657);
and U16357 (N_16357,N_15692,N_15673);
or U16358 (N_16358,N_15428,N_15270);
and U16359 (N_16359,N_15538,N_15544);
and U16360 (N_16360,N_15812,N_15429);
nor U16361 (N_16361,N_15931,N_15370);
and U16362 (N_16362,N_15884,N_15378);
nor U16363 (N_16363,N_15645,N_15878);
xnor U16364 (N_16364,N_15279,N_15310);
and U16365 (N_16365,N_15740,N_15247);
and U16366 (N_16366,N_15632,N_15549);
nor U16367 (N_16367,N_15201,N_15959);
nor U16368 (N_16368,N_15404,N_15763);
nor U16369 (N_16369,N_15285,N_15384);
nand U16370 (N_16370,N_15691,N_15328);
nand U16371 (N_16371,N_15368,N_15431);
and U16372 (N_16372,N_15452,N_15693);
and U16373 (N_16373,N_15820,N_15460);
nand U16374 (N_16374,N_15966,N_15322);
nor U16375 (N_16375,N_15444,N_15734);
nand U16376 (N_16376,N_15390,N_15334);
and U16377 (N_16377,N_15992,N_15560);
and U16378 (N_16378,N_15492,N_15450);
nand U16379 (N_16379,N_15410,N_15638);
nand U16380 (N_16380,N_15658,N_15993);
or U16381 (N_16381,N_15852,N_15902);
nor U16382 (N_16382,N_15881,N_15528);
and U16383 (N_16383,N_15261,N_15580);
nor U16384 (N_16384,N_15957,N_15676);
nor U16385 (N_16385,N_15717,N_15828);
or U16386 (N_16386,N_15281,N_15408);
and U16387 (N_16387,N_15943,N_15249);
nor U16388 (N_16388,N_15552,N_15225);
nand U16389 (N_16389,N_15324,N_15853);
and U16390 (N_16390,N_15745,N_15588);
or U16391 (N_16391,N_15203,N_15527);
nand U16392 (N_16392,N_15379,N_15348);
nor U16393 (N_16393,N_15775,N_15934);
and U16394 (N_16394,N_15346,N_15439);
nor U16395 (N_16395,N_15974,N_15336);
nor U16396 (N_16396,N_15542,N_15940);
nor U16397 (N_16397,N_15794,N_15844);
nor U16398 (N_16398,N_15266,N_15749);
nor U16399 (N_16399,N_15489,N_15497);
nand U16400 (N_16400,N_15523,N_15900);
and U16401 (N_16401,N_15334,N_15684);
and U16402 (N_16402,N_15517,N_15813);
nor U16403 (N_16403,N_15766,N_15731);
or U16404 (N_16404,N_15291,N_15408);
or U16405 (N_16405,N_15245,N_15293);
nor U16406 (N_16406,N_15345,N_15767);
and U16407 (N_16407,N_15483,N_15640);
nor U16408 (N_16408,N_15471,N_15676);
nor U16409 (N_16409,N_15914,N_15227);
nand U16410 (N_16410,N_15644,N_15351);
or U16411 (N_16411,N_15665,N_15678);
nor U16412 (N_16412,N_15689,N_15452);
and U16413 (N_16413,N_15821,N_15410);
and U16414 (N_16414,N_15883,N_15588);
and U16415 (N_16415,N_15960,N_15720);
and U16416 (N_16416,N_15805,N_15920);
nor U16417 (N_16417,N_15843,N_15670);
nand U16418 (N_16418,N_15716,N_15994);
and U16419 (N_16419,N_15506,N_15572);
and U16420 (N_16420,N_15816,N_15475);
nand U16421 (N_16421,N_15441,N_15319);
nor U16422 (N_16422,N_15546,N_15935);
or U16423 (N_16423,N_15866,N_15888);
nand U16424 (N_16424,N_15853,N_15704);
and U16425 (N_16425,N_15735,N_15325);
nand U16426 (N_16426,N_15299,N_15632);
nand U16427 (N_16427,N_15648,N_15300);
or U16428 (N_16428,N_15874,N_15766);
or U16429 (N_16429,N_15361,N_15428);
nor U16430 (N_16430,N_15945,N_15248);
nor U16431 (N_16431,N_15464,N_15343);
or U16432 (N_16432,N_15858,N_15930);
or U16433 (N_16433,N_15498,N_15493);
nor U16434 (N_16434,N_15991,N_15497);
nand U16435 (N_16435,N_15239,N_15737);
and U16436 (N_16436,N_15333,N_15489);
nand U16437 (N_16437,N_15294,N_15206);
and U16438 (N_16438,N_15721,N_15744);
and U16439 (N_16439,N_15275,N_15202);
nor U16440 (N_16440,N_15806,N_15974);
or U16441 (N_16441,N_15676,N_15411);
and U16442 (N_16442,N_15483,N_15498);
or U16443 (N_16443,N_15895,N_15429);
nor U16444 (N_16444,N_15313,N_15534);
and U16445 (N_16445,N_15461,N_15573);
nor U16446 (N_16446,N_15236,N_15699);
nand U16447 (N_16447,N_15470,N_15693);
nand U16448 (N_16448,N_15559,N_15285);
nor U16449 (N_16449,N_15600,N_15224);
and U16450 (N_16450,N_15789,N_15460);
or U16451 (N_16451,N_15864,N_15933);
nor U16452 (N_16452,N_15471,N_15757);
and U16453 (N_16453,N_15382,N_15364);
or U16454 (N_16454,N_15566,N_15219);
nand U16455 (N_16455,N_15834,N_15891);
nor U16456 (N_16456,N_15564,N_15780);
and U16457 (N_16457,N_15935,N_15337);
nor U16458 (N_16458,N_15782,N_15835);
or U16459 (N_16459,N_15254,N_15935);
or U16460 (N_16460,N_15590,N_15577);
or U16461 (N_16461,N_15566,N_15642);
nand U16462 (N_16462,N_15226,N_15477);
or U16463 (N_16463,N_15238,N_15599);
nor U16464 (N_16464,N_15920,N_15377);
and U16465 (N_16465,N_15590,N_15266);
or U16466 (N_16466,N_15413,N_15357);
or U16467 (N_16467,N_15574,N_15424);
nand U16468 (N_16468,N_15411,N_15773);
and U16469 (N_16469,N_15228,N_15545);
nand U16470 (N_16470,N_15982,N_15438);
nand U16471 (N_16471,N_15345,N_15586);
nand U16472 (N_16472,N_15904,N_15978);
and U16473 (N_16473,N_15772,N_15424);
nor U16474 (N_16474,N_15572,N_15230);
or U16475 (N_16475,N_15723,N_15590);
nor U16476 (N_16476,N_15665,N_15340);
nand U16477 (N_16477,N_15218,N_15728);
nor U16478 (N_16478,N_15230,N_15672);
nor U16479 (N_16479,N_15706,N_15922);
or U16480 (N_16480,N_15230,N_15475);
or U16481 (N_16481,N_15646,N_15753);
or U16482 (N_16482,N_15335,N_15404);
or U16483 (N_16483,N_15718,N_15763);
nor U16484 (N_16484,N_15451,N_15589);
nor U16485 (N_16485,N_15348,N_15893);
or U16486 (N_16486,N_15900,N_15404);
or U16487 (N_16487,N_15819,N_15227);
nor U16488 (N_16488,N_15923,N_15637);
nor U16489 (N_16489,N_15836,N_15523);
nand U16490 (N_16490,N_15568,N_15540);
and U16491 (N_16491,N_15527,N_15633);
and U16492 (N_16492,N_15947,N_15813);
and U16493 (N_16493,N_15397,N_15408);
nor U16494 (N_16494,N_15367,N_15803);
and U16495 (N_16495,N_15756,N_15598);
or U16496 (N_16496,N_15311,N_15732);
or U16497 (N_16497,N_15631,N_15902);
or U16498 (N_16498,N_15337,N_15806);
and U16499 (N_16499,N_15985,N_15437);
or U16500 (N_16500,N_15399,N_15417);
and U16501 (N_16501,N_15326,N_15926);
and U16502 (N_16502,N_15211,N_15731);
and U16503 (N_16503,N_15571,N_15554);
and U16504 (N_16504,N_15210,N_15439);
nand U16505 (N_16505,N_15414,N_15447);
and U16506 (N_16506,N_15212,N_15387);
and U16507 (N_16507,N_15738,N_15876);
and U16508 (N_16508,N_15765,N_15434);
and U16509 (N_16509,N_15333,N_15855);
nand U16510 (N_16510,N_15328,N_15476);
or U16511 (N_16511,N_15985,N_15664);
nor U16512 (N_16512,N_15612,N_15516);
and U16513 (N_16513,N_15810,N_15742);
nand U16514 (N_16514,N_15598,N_15678);
xnor U16515 (N_16515,N_15566,N_15561);
nor U16516 (N_16516,N_15494,N_15509);
and U16517 (N_16517,N_15938,N_15709);
and U16518 (N_16518,N_15646,N_15421);
or U16519 (N_16519,N_15950,N_15679);
or U16520 (N_16520,N_15310,N_15215);
nand U16521 (N_16521,N_15556,N_15649);
and U16522 (N_16522,N_15434,N_15263);
nor U16523 (N_16523,N_15456,N_15312);
and U16524 (N_16524,N_15987,N_15626);
nor U16525 (N_16525,N_15485,N_15692);
nor U16526 (N_16526,N_15502,N_15268);
or U16527 (N_16527,N_15459,N_15561);
or U16528 (N_16528,N_15828,N_15420);
nor U16529 (N_16529,N_15986,N_15595);
and U16530 (N_16530,N_15408,N_15811);
or U16531 (N_16531,N_15555,N_15991);
nand U16532 (N_16532,N_15891,N_15503);
and U16533 (N_16533,N_15463,N_15475);
and U16534 (N_16534,N_15792,N_15799);
nand U16535 (N_16535,N_15910,N_15757);
nor U16536 (N_16536,N_15798,N_15707);
and U16537 (N_16537,N_15436,N_15633);
or U16538 (N_16538,N_15482,N_15731);
nor U16539 (N_16539,N_15649,N_15393);
and U16540 (N_16540,N_15582,N_15558);
nor U16541 (N_16541,N_15849,N_15972);
nand U16542 (N_16542,N_15277,N_15690);
nor U16543 (N_16543,N_15517,N_15281);
nand U16544 (N_16544,N_15483,N_15635);
and U16545 (N_16545,N_15311,N_15207);
nor U16546 (N_16546,N_15673,N_15685);
or U16547 (N_16547,N_15977,N_15853);
or U16548 (N_16548,N_15302,N_15439);
or U16549 (N_16549,N_15291,N_15959);
nor U16550 (N_16550,N_15422,N_15412);
nand U16551 (N_16551,N_15317,N_15544);
xor U16552 (N_16552,N_15296,N_15405);
and U16553 (N_16553,N_15676,N_15332);
nand U16554 (N_16554,N_15462,N_15891);
nand U16555 (N_16555,N_15678,N_15387);
nor U16556 (N_16556,N_15358,N_15528);
and U16557 (N_16557,N_15789,N_15857);
nor U16558 (N_16558,N_15244,N_15404);
nor U16559 (N_16559,N_15495,N_15593);
nor U16560 (N_16560,N_15984,N_15608);
and U16561 (N_16561,N_15390,N_15720);
or U16562 (N_16562,N_15604,N_15954);
nand U16563 (N_16563,N_15686,N_15379);
or U16564 (N_16564,N_15311,N_15926);
or U16565 (N_16565,N_15801,N_15396);
nor U16566 (N_16566,N_15204,N_15617);
or U16567 (N_16567,N_15846,N_15901);
nor U16568 (N_16568,N_15268,N_15242);
or U16569 (N_16569,N_15881,N_15599);
nor U16570 (N_16570,N_15765,N_15631);
or U16571 (N_16571,N_15805,N_15545);
or U16572 (N_16572,N_15703,N_15920);
nand U16573 (N_16573,N_15323,N_15249);
or U16574 (N_16574,N_15987,N_15484);
nor U16575 (N_16575,N_15829,N_15853);
xnor U16576 (N_16576,N_15224,N_15740);
nand U16577 (N_16577,N_15753,N_15922);
nor U16578 (N_16578,N_15942,N_15907);
and U16579 (N_16579,N_15855,N_15615);
nor U16580 (N_16580,N_15281,N_15828);
nor U16581 (N_16581,N_15366,N_15310);
nor U16582 (N_16582,N_15659,N_15341);
or U16583 (N_16583,N_15674,N_15741);
nand U16584 (N_16584,N_15711,N_15747);
nand U16585 (N_16585,N_15360,N_15201);
nand U16586 (N_16586,N_15607,N_15600);
or U16587 (N_16587,N_15749,N_15204);
xnor U16588 (N_16588,N_15630,N_15752);
nand U16589 (N_16589,N_15877,N_15312);
or U16590 (N_16590,N_15715,N_15683);
nand U16591 (N_16591,N_15860,N_15671);
nor U16592 (N_16592,N_15421,N_15885);
or U16593 (N_16593,N_15393,N_15402);
nor U16594 (N_16594,N_15597,N_15442);
xnor U16595 (N_16595,N_15983,N_15902);
or U16596 (N_16596,N_15232,N_15215);
or U16597 (N_16597,N_15817,N_15710);
or U16598 (N_16598,N_15753,N_15232);
nand U16599 (N_16599,N_15939,N_15895);
nand U16600 (N_16600,N_15258,N_15771);
nor U16601 (N_16601,N_15419,N_15402);
and U16602 (N_16602,N_15643,N_15451);
nor U16603 (N_16603,N_15299,N_15244);
nor U16604 (N_16604,N_15393,N_15258);
or U16605 (N_16605,N_15746,N_15954);
nor U16606 (N_16606,N_15465,N_15642);
nor U16607 (N_16607,N_15506,N_15488);
and U16608 (N_16608,N_15486,N_15610);
and U16609 (N_16609,N_15634,N_15389);
nor U16610 (N_16610,N_15390,N_15699);
nor U16611 (N_16611,N_15885,N_15414);
nor U16612 (N_16612,N_15670,N_15554);
nand U16613 (N_16613,N_15326,N_15919);
or U16614 (N_16614,N_15727,N_15809);
nor U16615 (N_16615,N_15476,N_15801);
and U16616 (N_16616,N_15544,N_15769);
and U16617 (N_16617,N_15370,N_15599);
and U16618 (N_16618,N_15600,N_15552);
nand U16619 (N_16619,N_15505,N_15996);
and U16620 (N_16620,N_15917,N_15264);
nand U16621 (N_16621,N_15883,N_15684);
and U16622 (N_16622,N_15502,N_15482);
and U16623 (N_16623,N_15309,N_15657);
nor U16624 (N_16624,N_15240,N_15675);
and U16625 (N_16625,N_15777,N_15786);
and U16626 (N_16626,N_15801,N_15502);
or U16627 (N_16627,N_15436,N_15475);
or U16628 (N_16628,N_15728,N_15376);
nand U16629 (N_16629,N_15518,N_15694);
and U16630 (N_16630,N_15987,N_15793);
and U16631 (N_16631,N_15901,N_15428);
nand U16632 (N_16632,N_15234,N_15988);
nand U16633 (N_16633,N_15909,N_15445);
nand U16634 (N_16634,N_15656,N_15772);
or U16635 (N_16635,N_15379,N_15432);
nor U16636 (N_16636,N_15606,N_15655);
nor U16637 (N_16637,N_15938,N_15898);
or U16638 (N_16638,N_15778,N_15773);
nand U16639 (N_16639,N_15945,N_15888);
nand U16640 (N_16640,N_15314,N_15931);
nand U16641 (N_16641,N_15510,N_15805);
nor U16642 (N_16642,N_15665,N_15795);
nand U16643 (N_16643,N_15785,N_15370);
nor U16644 (N_16644,N_15954,N_15246);
xor U16645 (N_16645,N_15867,N_15486);
nand U16646 (N_16646,N_15583,N_15670);
or U16647 (N_16647,N_15247,N_15272);
nand U16648 (N_16648,N_15486,N_15412);
nand U16649 (N_16649,N_15553,N_15314);
nand U16650 (N_16650,N_15475,N_15261);
or U16651 (N_16651,N_15632,N_15883);
or U16652 (N_16652,N_15841,N_15216);
nor U16653 (N_16653,N_15344,N_15743);
or U16654 (N_16654,N_15265,N_15777);
or U16655 (N_16655,N_15230,N_15848);
nand U16656 (N_16656,N_15610,N_15398);
nand U16657 (N_16657,N_15460,N_15717);
and U16658 (N_16658,N_15692,N_15856);
and U16659 (N_16659,N_15486,N_15360);
nand U16660 (N_16660,N_15238,N_15749);
nand U16661 (N_16661,N_15652,N_15679);
nand U16662 (N_16662,N_15910,N_15704);
nand U16663 (N_16663,N_15305,N_15956);
and U16664 (N_16664,N_15318,N_15846);
nand U16665 (N_16665,N_15471,N_15296);
nor U16666 (N_16666,N_15984,N_15686);
nand U16667 (N_16667,N_15410,N_15782);
nor U16668 (N_16668,N_15849,N_15576);
nor U16669 (N_16669,N_15304,N_15369);
nand U16670 (N_16670,N_15513,N_15328);
nand U16671 (N_16671,N_15500,N_15748);
xnor U16672 (N_16672,N_15768,N_15892);
and U16673 (N_16673,N_15968,N_15860);
or U16674 (N_16674,N_15886,N_15208);
nor U16675 (N_16675,N_15414,N_15526);
or U16676 (N_16676,N_15384,N_15681);
nor U16677 (N_16677,N_15591,N_15594);
nand U16678 (N_16678,N_15346,N_15795);
nand U16679 (N_16679,N_15389,N_15332);
and U16680 (N_16680,N_15616,N_15551);
nand U16681 (N_16681,N_15564,N_15597);
or U16682 (N_16682,N_15280,N_15380);
nor U16683 (N_16683,N_15207,N_15460);
or U16684 (N_16684,N_15249,N_15800);
or U16685 (N_16685,N_15291,N_15788);
or U16686 (N_16686,N_15694,N_15201);
nor U16687 (N_16687,N_15601,N_15468);
or U16688 (N_16688,N_15396,N_15391);
and U16689 (N_16689,N_15633,N_15662);
nand U16690 (N_16690,N_15922,N_15656);
nor U16691 (N_16691,N_15977,N_15444);
nand U16692 (N_16692,N_15789,N_15610);
or U16693 (N_16693,N_15859,N_15539);
nor U16694 (N_16694,N_15283,N_15472);
nor U16695 (N_16695,N_15610,N_15890);
nand U16696 (N_16696,N_15223,N_15965);
nor U16697 (N_16697,N_15606,N_15414);
nor U16698 (N_16698,N_15868,N_15867);
and U16699 (N_16699,N_15887,N_15489);
or U16700 (N_16700,N_15263,N_15400);
nor U16701 (N_16701,N_15914,N_15659);
and U16702 (N_16702,N_15964,N_15573);
nand U16703 (N_16703,N_15448,N_15312);
or U16704 (N_16704,N_15793,N_15878);
nor U16705 (N_16705,N_15987,N_15692);
or U16706 (N_16706,N_15291,N_15844);
and U16707 (N_16707,N_15966,N_15400);
nand U16708 (N_16708,N_15517,N_15794);
nor U16709 (N_16709,N_15909,N_15937);
nand U16710 (N_16710,N_15654,N_15440);
nor U16711 (N_16711,N_15245,N_15231);
nor U16712 (N_16712,N_15341,N_15286);
or U16713 (N_16713,N_15401,N_15312);
and U16714 (N_16714,N_15263,N_15449);
nand U16715 (N_16715,N_15735,N_15366);
nand U16716 (N_16716,N_15763,N_15330);
or U16717 (N_16717,N_15790,N_15712);
nand U16718 (N_16718,N_15680,N_15210);
or U16719 (N_16719,N_15831,N_15622);
nand U16720 (N_16720,N_15915,N_15316);
or U16721 (N_16721,N_15953,N_15374);
nor U16722 (N_16722,N_15557,N_15330);
or U16723 (N_16723,N_15773,N_15506);
nand U16724 (N_16724,N_15889,N_15428);
and U16725 (N_16725,N_15256,N_15475);
and U16726 (N_16726,N_15673,N_15393);
nor U16727 (N_16727,N_15495,N_15519);
nand U16728 (N_16728,N_15306,N_15529);
nor U16729 (N_16729,N_15491,N_15527);
or U16730 (N_16730,N_15877,N_15300);
and U16731 (N_16731,N_15378,N_15650);
nand U16732 (N_16732,N_15902,N_15273);
or U16733 (N_16733,N_15648,N_15828);
nor U16734 (N_16734,N_15421,N_15708);
nand U16735 (N_16735,N_15575,N_15451);
and U16736 (N_16736,N_15312,N_15241);
and U16737 (N_16737,N_15625,N_15778);
or U16738 (N_16738,N_15768,N_15811);
nor U16739 (N_16739,N_15866,N_15480);
or U16740 (N_16740,N_15419,N_15981);
nand U16741 (N_16741,N_15694,N_15937);
and U16742 (N_16742,N_15311,N_15878);
and U16743 (N_16743,N_15852,N_15940);
and U16744 (N_16744,N_15838,N_15970);
and U16745 (N_16745,N_15741,N_15621);
nand U16746 (N_16746,N_15379,N_15383);
or U16747 (N_16747,N_15380,N_15482);
or U16748 (N_16748,N_15945,N_15339);
and U16749 (N_16749,N_15238,N_15868);
nor U16750 (N_16750,N_15796,N_15369);
or U16751 (N_16751,N_15999,N_15493);
nor U16752 (N_16752,N_15330,N_15634);
and U16753 (N_16753,N_15528,N_15772);
nand U16754 (N_16754,N_15518,N_15451);
and U16755 (N_16755,N_15513,N_15652);
nor U16756 (N_16756,N_15550,N_15945);
or U16757 (N_16757,N_15288,N_15384);
nand U16758 (N_16758,N_15284,N_15646);
nor U16759 (N_16759,N_15546,N_15337);
or U16760 (N_16760,N_15722,N_15595);
nand U16761 (N_16761,N_15480,N_15847);
and U16762 (N_16762,N_15347,N_15853);
and U16763 (N_16763,N_15227,N_15683);
or U16764 (N_16764,N_15308,N_15778);
nand U16765 (N_16765,N_15624,N_15785);
and U16766 (N_16766,N_15434,N_15551);
or U16767 (N_16767,N_15323,N_15402);
or U16768 (N_16768,N_15535,N_15455);
or U16769 (N_16769,N_15782,N_15967);
and U16770 (N_16770,N_15647,N_15445);
and U16771 (N_16771,N_15913,N_15401);
and U16772 (N_16772,N_15870,N_15813);
nor U16773 (N_16773,N_15888,N_15925);
or U16774 (N_16774,N_15251,N_15906);
nor U16775 (N_16775,N_15662,N_15428);
nor U16776 (N_16776,N_15652,N_15621);
nor U16777 (N_16777,N_15540,N_15676);
nand U16778 (N_16778,N_15527,N_15365);
nor U16779 (N_16779,N_15396,N_15776);
and U16780 (N_16780,N_15278,N_15936);
nand U16781 (N_16781,N_15889,N_15461);
nor U16782 (N_16782,N_15449,N_15925);
nand U16783 (N_16783,N_15431,N_15818);
nand U16784 (N_16784,N_15535,N_15680);
nand U16785 (N_16785,N_15429,N_15865);
or U16786 (N_16786,N_15718,N_15430);
or U16787 (N_16787,N_15254,N_15752);
nor U16788 (N_16788,N_15264,N_15379);
or U16789 (N_16789,N_15921,N_15885);
or U16790 (N_16790,N_15231,N_15737);
and U16791 (N_16791,N_15354,N_15773);
nor U16792 (N_16792,N_15886,N_15579);
or U16793 (N_16793,N_15224,N_15237);
nand U16794 (N_16794,N_15471,N_15805);
nor U16795 (N_16795,N_15283,N_15226);
and U16796 (N_16796,N_15872,N_15930);
or U16797 (N_16797,N_15640,N_15735);
and U16798 (N_16798,N_15445,N_15569);
and U16799 (N_16799,N_15231,N_15292);
or U16800 (N_16800,N_16549,N_16755);
nand U16801 (N_16801,N_16408,N_16345);
nand U16802 (N_16802,N_16750,N_16541);
nand U16803 (N_16803,N_16438,N_16735);
nand U16804 (N_16804,N_16448,N_16537);
nand U16805 (N_16805,N_16210,N_16275);
nand U16806 (N_16806,N_16709,N_16294);
nand U16807 (N_16807,N_16002,N_16258);
nor U16808 (N_16808,N_16401,N_16336);
or U16809 (N_16809,N_16502,N_16024);
or U16810 (N_16810,N_16256,N_16273);
or U16811 (N_16811,N_16638,N_16053);
nor U16812 (N_16812,N_16089,N_16375);
nand U16813 (N_16813,N_16251,N_16607);
nand U16814 (N_16814,N_16324,N_16550);
nand U16815 (N_16815,N_16070,N_16492);
or U16816 (N_16816,N_16392,N_16429);
and U16817 (N_16817,N_16302,N_16621);
and U16818 (N_16818,N_16741,N_16241);
or U16819 (N_16819,N_16214,N_16304);
and U16820 (N_16820,N_16376,N_16413);
or U16821 (N_16821,N_16087,N_16091);
nand U16822 (N_16822,N_16298,N_16516);
or U16823 (N_16823,N_16104,N_16022);
and U16824 (N_16824,N_16487,N_16268);
nand U16825 (N_16825,N_16523,N_16416);
and U16826 (N_16826,N_16309,N_16675);
nor U16827 (N_16827,N_16546,N_16643);
nand U16828 (N_16828,N_16757,N_16035);
nor U16829 (N_16829,N_16235,N_16605);
or U16830 (N_16830,N_16146,N_16283);
and U16831 (N_16831,N_16797,N_16548);
nor U16832 (N_16832,N_16059,N_16759);
or U16833 (N_16833,N_16494,N_16719);
and U16834 (N_16834,N_16027,N_16667);
xnor U16835 (N_16835,N_16303,N_16028);
nand U16836 (N_16836,N_16721,N_16430);
and U16837 (N_16837,N_16185,N_16247);
or U16838 (N_16838,N_16432,N_16468);
or U16839 (N_16839,N_16318,N_16535);
nor U16840 (N_16840,N_16503,N_16533);
and U16841 (N_16841,N_16019,N_16680);
nand U16842 (N_16842,N_16579,N_16493);
nor U16843 (N_16843,N_16219,N_16152);
nor U16844 (N_16844,N_16658,N_16103);
and U16845 (N_16845,N_16061,N_16124);
nor U16846 (N_16846,N_16562,N_16459);
and U16847 (N_16847,N_16161,N_16334);
and U16848 (N_16848,N_16718,N_16566);
nand U16849 (N_16849,N_16062,N_16505);
nand U16850 (N_16850,N_16526,N_16326);
nand U16851 (N_16851,N_16199,N_16005);
and U16852 (N_16852,N_16159,N_16598);
and U16853 (N_16853,N_16099,N_16329);
nor U16854 (N_16854,N_16398,N_16726);
and U16855 (N_16855,N_16732,N_16385);
and U16856 (N_16856,N_16204,N_16120);
or U16857 (N_16857,N_16007,N_16637);
nor U16858 (N_16858,N_16601,N_16572);
nor U16859 (N_16859,N_16313,N_16282);
nor U16860 (N_16860,N_16001,N_16631);
nand U16861 (N_16861,N_16754,N_16292);
nand U16862 (N_16862,N_16047,N_16195);
nor U16863 (N_16863,N_16011,N_16397);
and U16864 (N_16864,N_16236,N_16540);
and U16865 (N_16865,N_16229,N_16069);
nor U16866 (N_16866,N_16246,N_16362);
nand U16867 (N_16867,N_16350,N_16702);
or U16868 (N_16868,N_16696,N_16349);
nand U16869 (N_16869,N_16288,N_16181);
or U16870 (N_16870,N_16421,N_16271);
and U16871 (N_16871,N_16173,N_16434);
and U16872 (N_16872,N_16232,N_16046);
and U16873 (N_16873,N_16188,N_16426);
or U16874 (N_16874,N_16386,N_16372);
or U16875 (N_16875,N_16354,N_16048);
or U16876 (N_16876,N_16427,N_16619);
and U16877 (N_16877,N_16064,N_16593);
nor U16878 (N_16878,N_16636,N_16314);
nor U16879 (N_16879,N_16629,N_16100);
or U16880 (N_16880,N_16690,N_16399);
and U16881 (N_16881,N_16583,N_16093);
or U16882 (N_16882,N_16641,N_16012);
nor U16883 (N_16883,N_16708,N_16633);
nor U16884 (N_16884,N_16435,N_16685);
and U16885 (N_16885,N_16003,N_16105);
and U16886 (N_16886,N_16267,N_16769);
nor U16887 (N_16887,N_16114,N_16649);
nand U16888 (N_16888,N_16361,N_16163);
nand U16889 (N_16889,N_16652,N_16119);
or U16890 (N_16890,N_16728,N_16058);
or U16891 (N_16891,N_16265,N_16166);
or U16892 (N_16892,N_16575,N_16151);
nand U16893 (N_16893,N_16238,N_16066);
nor U16894 (N_16894,N_16739,N_16196);
nand U16895 (N_16895,N_16230,N_16520);
nand U16896 (N_16896,N_16514,N_16014);
or U16897 (N_16897,N_16194,N_16457);
nor U16898 (N_16898,N_16560,N_16691);
or U16899 (N_16899,N_16594,N_16076);
and U16900 (N_16900,N_16369,N_16351);
nor U16901 (N_16901,N_16308,N_16772);
or U16902 (N_16902,N_16664,N_16272);
nor U16903 (N_16903,N_16297,N_16080);
and U16904 (N_16904,N_16600,N_16259);
nor U16905 (N_16905,N_16559,N_16316);
nor U16906 (N_16906,N_16711,N_16679);
or U16907 (N_16907,N_16176,N_16556);
or U16908 (N_16908,N_16625,N_16443);
and U16909 (N_16909,N_16131,N_16720);
nor U16910 (N_16910,N_16142,N_16244);
xor U16911 (N_16911,N_16618,N_16578);
nand U16912 (N_16912,N_16422,N_16778);
or U16913 (N_16913,N_16333,N_16261);
or U16914 (N_16914,N_16057,N_16522);
nor U16915 (N_16915,N_16228,N_16032);
nor U16916 (N_16916,N_16604,N_16111);
and U16917 (N_16917,N_16464,N_16175);
nor U16918 (N_16918,N_16642,N_16130);
or U16919 (N_16919,N_16786,N_16359);
or U16920 (N_16920,N_16731,N_16060);
and U16921 (N_16921,N_16155,N_16542);
and U16922 (N_16922,N_16323,N_16306);
and U16923 (N_16923,N_16133,N_16410);
xor U16924 (N_16924,N_16678,N_16123);
or U16925 (N_16925,N_16599,N_16231);
and U16926 (N_16926,N_16743,N_16178);
or U16927 (N_16927,N_16050,N_16092);
nand U16928 (N_16928,N_16332,N_16337);
nand U16929 (N_16929,N_16781,N_16084);
or U16930 (N_16930,N_16446,N_16669);
and U16931 (N_16931,N_16738,N_16191);
nand U16932 (N_16932,N_16474,N_16248);
nand U16933 (N_16933,N_16668,N_16545);
nor U16934 (N_16934,N_16041,N_16703);
or U16935 (N_16935,N_16499,N_16149);
nor U16936 (N_16936,N_16409,N_16209);
nor U16937 (N_16937,N_16543,N_16379);
nor U16938 (N_16938,N_16775,N_16000);
nand U16939 (N_16939,N_16747,N_16277);
and U16940 (N_16940,N_16798,N_16608);
nand U16941 (N_16941,N_16179,N_16138);
or U16942 (N_16942,N_16673,N_16164);
or U16943 (N_16943,N_16102,N_16697);
and U16944 (N_16944,N_16029,N_16097);
nand U16945 (N_16945,N_16733,N_16752);
xor U16946 (N_16946,N_16490,N_16167);
nor U16947 (N_16947,N_16687,N_16215);
nor U16948 (N_16948,N_16192,N_16407);
nor U16949 (N_16949,N_16193,N_16026);
or U16950 (N_16950,N_16476,N_16383);
nor U16951 (N_16951,N_16758,N_16237);
nor U16952 (N_16952,N_16170,N_16539);
and U16953 (N_16953,N_16683,N_16287);
nand U16954 (N_16954,N_16016,N_16343);
or U16955 (N_16955,N_16420,N_16730);
nor U16956 (N_16956,N_16141,N_16063);
nand U16957 (N_16957,N_16472,N_16122);
nor U16958 (N_16958,N_16473,N_16394);
and U16959 (N_16959,N_16441,N_16112);
nand U16960 (N_16960,N_16582,N_16322);
nor U16961 (N_16961,N_16727,N_16686);
and U16962 (N_16962,N_16342,N_16634);
or U16963 (N_16963,N_16065,N_16190);
nor U16964 (N_16964,N_16544,N_16762);
nand U16965 (N_16965,N_16495,N_16653);
or U16966 (N_16966,N_16239,N_16144);
nand U16967 (N_16967,N_16714,N_16305);
and U16968 (N_16968,N_16617,N_16347);
or U16969 (N_16969,N_16234,N_16094);
nor U16970 (N_16970,N_16651,N_16475);
and U16971 (N_16971,N_16320,N_16040);
and U16972 (N_16972,N_16554,N_16736);
nand U16973 (N_16973,N_16281,N_16143);
and U16974 (N_16974,N_16612,N_16371);
nor U16975 (N_16975,N_16116,N_16025);
or U16976 (N_16976,N_16782,N_16174);
and U16977 (N_16977,N_16460,N_16467);
nor U16978 (N_16978,N_16716,N_16201);
and U16979 (N_16979,N_16341,N_16573);
and U16980 (N_16980,N_16425,N_16513);
and U16981 (N_16981,N_16074,N_16626);
or U16982 (N_16982,N_16036,N_16682);
nand U16983 (N_16983,N_16646,N_16411);
nand U16984 (N_16984,N_16623,N_16712);
nor U16985 (N_16985,N_16761,N_16722);
nand U16986 (N_16986,N_16213,N_16156);
or U16987 (N_16987,N_16037,N_16603);
nor U16988 (N_16988,N_16574,N_16158);
nor U16989 (N_16989,N_16510,N_16627);
nor U16990 (N_16990,N_16734,N_16795);
nor U16991 (N_16991,N_16746,N_16455);
nand U16992 (N_16992,N_16307,N_16291);
xor U16993 (N_16993,N_16364,N_16796);
and U16994 (N_16994,N_16588,N_16663);
nor U16995 (N_16995,N_16374,N_16278);
or U16996 (N_16996,N_16462,N_16216);
and U16997 (N_16997,N_16134,N_16445);
nand U16998 (N_16998,N_16504,N_16498);
xor U16999 (N_16999,N_16205,N_16515);
nand U17000 (N_17000,N_16373,N_16034);
and U17001 (N_17001,N_16260,N_16676);
or U17002 (N_17002,N_16128,N_16404);
nand U17003 (N_17003,N_16480,N_16269);
and U17004 (N_17004,N_16452,N_16787);
nor U17005 (N_17005,N_16530,N_16381);
or U17006 (N_17006,N_16095,N_16115);
or U17007 (N_17007,N_16671,N_16224);
nand U17008 (N_17008,N_16052,N_16140);
nand U17009 (N_17009,N_16565,N_16107);
nand U17010 (N_17010,N_16039,N_16577);
or U17011 (N_17011,N_16776,N_16589);
nand U17012 (N_17012,N_16129,N_16299);
nor U17013 (N_17013,N_16483,N_16713);
and U17014 (N_17014,N_16370,N_16774);
xnor U17015 (N_17015,N_16551,N_16295);
nand U17016 (N_17016,N_16558,N_16531);
nand U17017 (N_17017,N_16528,N_16169);
and U17018 (N_17018,N_16581,N_16681);
nor U17019 (N_17019,N_16512,N_16279);
nor U17020 (N_17020,N_16606,N_16098);
and U17021 (N_17021,N_16110,N_16406);
nand U17022 (N_17022,N_16444,N_16628);
nand U17023 (N_17023,N_16249,N_16742);
and U17024 (N_17024,N_16763,N_16339);
nor U17025 (N_17025,N_16765,N_16262);
and U17026 (N_17026,N_16317,N_16729);
or U17027 (N_17027,N_16132,N_16799);
and U17028 (N_17028,N_16180,N_16447);
or U17029 (N_17029,N_16597,N_16055);
nand U17030 (N_17030,N_16771,N_16698);
and U17031 (N_17031,N_16610,N_16616);
nor U17032 (N_17032,N_16072,N_16365);
nand U17033 (N_17033,N_16276,N_16009);
nand U17034 (N_17034,N_16699,N_16078);
nor U17035 (N_17035,N_16783,N_16335);
nor U17036 (N_17036,N_16118,N_16596);
and U17037 (N_17037,N_16785,N_16766);
nor U17038 (N_17038,N_16491,N_16356);
or U17039 (N_17039,N_16745,N_16650);
or U17040 (N_17040,N_16358,N_16218);
and U17041 (N_17041,N_16200,N_16075);
and U17042 (N_17042,N_16773,N_16154);
or U17043 (N_17043,N_16033,N_16454);
and U17044 (N_17044,N_16684,N_16564);
and U17045 (N_17045,N_16353,N_16252);
or U17046 (N_17046,N_16437,N_16451);
nand U17047 (N_17047,N_16340,N_16568);
and U17048 (N_17048,N_16428,N_16534);
or U17049 (N_17049,N_16157,N_16760);
or U17050 (N_17050,N_16160,N_16348);
and U17051 (N_17051,N_16693,N_16552);
or U17052 (N_17052,N_16255,N_16296);
or U17053 (N_17053,N_16384,N_16366);
nand U17054 (N_17054,N_16378,N_16021);
and U17055 (N_17055,N_16139,N_16784);
xor U17056 (N_17056,N_16109,N_16580);
nor U17057 (N_17057,N_16183,N_16792);
nand U17058 (N_17058,N_16590,N_16789);
and U17059 (N_17059,N_16496,N_16670);
nand U17060 (N_17060,N_16486,N_16688);
or U17061 (N_17061,N_16780,N_16082);
or U17062 (N_17062,N_16511,N_16478);
nor U17063 (N_17063,N_16700,N_16477);
and U17064 (N_17064,N_16790,N_16672);
nand U17065 (N_17065,N_16624,N_16660);
nand U17066 (N_17066,N_16471,N_16640);
or U17067 (N_17067,N_16657,N_16042);
nor U17068 (N_17068,N_16764,N_16587);
or U17069 (N_17069,N_16088,N_16327);
and U17070 (N_17070,N_16031,N_16479);
nand U17071 (N_17071,N_16225,N_16440);
and U17072 (N_17072,N_16484,N_16655);
and U17073 (N_17073,N_16096,N_16442);
or U17074 (N_17074,N_16217,N_16701);
or U17075 (N_17075,N_16692,N_16485);
and U17076 (N_17076,N_16274,N_16644);
nor U17077 (N_17077,N_16538,N_16312);
nor U17078 (N_17078,N_16125,N_16257);
nand U17079 (N_17079,N_16419,N_16101);
or U17080 (N_17080,N_16004,N_16632);
and U17081 (N_17081,N_16010,N_16223);
and U17082 (N_17082,N_16013,N_16553);
nor U17083 (N_17083,N_16389,N_16396);
or U17084 (N_17084,N_16767,N_16233);
nor U17085 (N_17085,N_16630,N_16054);
and U17086 (N_17086,N_16137,N_16266);
nor U17087 (N_17087,N_16507,N_16744);
nor U17088 (N_17088,N_16519,N_16254);
nor U17089 (N_17089,N_16635,N_16794);
nand U17090 (N_17090,N_16162,N_16221);
and U17091 (N_17091,N_16212,N_16319);
nand U17092 (N_17092,N_16108,N_16749);
and U17093 (N_17093,N_16020,N_16777);
nand U17094 (N_17094,N_16186,N_16240);
nand U17095 (N_17095,N_16456,N_16659);
nor U17096 (N_17096,N_16330,N_16211);
nand U17097 (N_17097,N_16208,N_16517);
and U17098 (N_17098,N_16038,N_16250);
nor U17099 (N_17099,N_16595,N_16226);
and U17100 (N_17100,N_16352,N_16725);
nand U17101 (N_17101,N_16424,N_16622);
or U17102 (N_17102,N_16068,N_16536);
nor U17103 (N_17103,N_16245,N_16506);
or U17104 (N_17104,N_16049,N_16338);
nand U17105 (N_17105,N_16051,N_16400);
and U17106 (N_17106,N_16723,N_16044);
or U17107 (N_17107,N_16740,N_16083);
nor U17108 (N_17108,N_16015,N_16045);
and U17109 (N_17109,N_16666,N_16465);
nand U17110 (N_17110,N_16086,N_16591);
nand U17111 (N_17111,N_16242,N_16207);
and U17112 (N_17112,N_16331,N_16592);
or U17113 (N_17113,N_16325,N_16301);
or U17114 (N_17114,N_16018,N_16390);
nor U17115 (N_17115,N_16586,N_16368);
or U17116 (N_17116,N_16469,N_16647);
nor U17117 (N_17117,N_16751,N_16439);
or U17118 (N_17118,N_16008,N_16253);
nor U17119 (N_17119,N_16023,N_16017);
and U17120 (N_17120,N_16508,N_16470);
nor U17121 (N_17121,N_16363,N_16584);
and U17122 (N_17122,N_16532,N_16656);
nor U17123 (N_17123,N_16187,N_16357);
or U17124 (N_17124,N_16521,N_16222);
nand U17125 (N_17125,N_16395,N_16321);
or U17126 (N_17126,N_16661,N_16576);
nor U17127 (N_17127,N_16529,N_16753);
nand U17128 (N_17128,N_16615,N_16127);
nand U17129 (N_17129,N_16768,N_16418);
and U17130 (N_17130,N_16563,N_16135);
nor U17131 (N_17131,N_16189,N_16360);
nor U17132 (N_17132,N_16184,N_16662);
or U17133 (N_17133,N_16449,N_16756);
or U17134 (N_17134,N_16150,N_16415);
nand U17135 (N_17135,N_16177,N_16171);
nor U17136 (N_17136,N_16412,N_16525);
nand U17137 (N_17137,N_16488,N_16770);
nand U17138 (N_17138,N_16518,N_16466);
nor U17139 (N_17139,N_16270,N_16620);
nor U17140 (N_17140,N_16106,N_16524);
and U17141 (N_17141,N_16489,N_16639);
or U17142 (N_17142,N_16677,N_16220);
nand U17143 (N_17143,N_16117,N_16147);
nand U17144 (N_17144,N_16706,N_16355);
and U17145 (N_17145,N_16609,N_16090);
and U17146 (N_17146,N_16431,N_16264);
nor U17147 (N_17147,N_16153,N_16056);
nand U17148 (N_17148,N_16715,N_16463);
or U17149 (N_17149,N_16284,N_16293);
or U17150 (N_17150,N_16547,N_16121);
or U17151 (N_17151,N_16085,N_16570);
or U17152 (N_17152,N_16500,N_16694);
and U17153 (N_17153,N_16388,N_16433);
or U17154 (N_17154,N_16748,N_16481);
or U17155 (N_17155,N_16067,N_16206);
and U17156 (N_17156,N_16614,N_16285);
nand U17157 (N_17157,N_16695,N_16779);
nor U17158 (N_17158,N_16689,N_16145);
nand U17159 (N_17159,N_16346,N_16665);
or U17160 (N_17160,N_16280,N_16263);
and U17161 (N_17161,N_16344,N_16203);
and U17162 (N_17162,N_16571,N_16509);
and U17163 (N_17163,N_16328,N_16788);
and U17164 (N_17164,N_16289,N_16081);
or U17165 (N_17165,N_16453,N_16710);
and U17166 (N_17166,N_16405,N_16414);
nor U17167 (N_17167,N_16417,N_16707);
or U17168 (N_17168,N_16705,N_16793);
nor U17169 (N_17169,N_16561,N_16202);
and U17170 (N_17170,N_16450,N_16030);
nor U17171 (N_17171,N_16458,N_16391);
and U17172 (N_17172,N_16077,N_16645);
nand U17173 (N_17173,N_16300,N_16602);
xnor U17174 (N_17174,N_16674,N_16403);
nand U17175 (N_17175,N_16071,N_16073);
nand U17176 (N_17176,N_16290,N_16402);
and U17177 (N_17177,N_16286,N_16497);
nand U17178 (N_17178,N_16585,N_16613);
nand U17179 (N_17179,N_16182,N_16557);
nand U17180 (N_17180,N_16382,N_16311);
and U17181 (N_17181,N_16126,N_16165);
or U17182 (N_17182,N_16654,N_16227);
nand U17183 (N_17183,N_16611,N_16567);
nor U17184 (N_17184,N_16393,N_16501);
and U17185 (N_17185,N_16043,N_16243);
and U17186 (N_17186,N_16377,N_16168);
or U17187 (N_17187,N_16315,N_16555);
and U17188 (N_17188,N_16527,N_16310);
and U17189 (N_17189,N_16148,N_16136);
nor U17190 (N_17190,N_16461,N_16423);
or U17191 (N_17191,N_16704,N_16648);
and U17192 (N_17192,N_16724,N_16387);
nand U17193 (N_17193,N_16737,N_16569);
or U17194 (N_17194,N_16172,N_16367);
or U17195 (N_17195,N_16380,N_16006);
and U17196 (N_17196,N_16079,N_16791);
and U17197 (N_17197,N_16436,N_16717);
and U17198 (N_17198,N_16113,N_16197);
nand U17199 (N_17199,N_16482,N_16198);
and U17200 (N_17200,N_16046,N_16478);
or U17201 (N_17201,N_16228,N_16765);
and U17202 (N_17202,N_16724,N_16124);
and U17203 (N_17203,N_16183,N_16237);
or U17204 (N_17204,N_16559,N_16767);
nand U17205 (N_17205,N_16616,N_16108);
and U17206 (N_17206,N_16068,N_16788);
nor U17207 (N_17207,N_16090,N_16033);
or U17208 (N_17208,N_16661,N_16251);
xor U17209 (N_17209,N_16104,N_16236);
nand U17210 (N_17210,N_16212,N_16219);
or U17211 (N_17211,N_16234,N_16190);
or U17212 (N_17212,N_16134,N_16361);
nand U17213 (N_17213,N_16791,N_16326);
nand U17214 (N_17214,N_16755,N_16522);
nand U17215 (N_17215,N_16226,N_16150);
nand U17216 (N_17216,N_16642,N_16638);
and U17217 (N_17217,N_16085,N_16463);
nor U17218 (N_17218,N_16547,N_16409);
or U17219 (N_17219,N_16462,N_16591);
and U17220 (N_17220,N_16051,N_16488);
nor U17221 (N_17221,N_16629,N_16217);
nor U17222 (N_17222,N_16589,N_16353);
and U17223 (N_17223,N_16307,N_16127);
nand U17224 (N_17224,N_16342,N_16313);
or U17225 (N_17225,N_16783,N_16411);
or U17226 (N_17226,N_16794,N_16417);
or U17227 (N_17227,N_16121,N_16080);
or U17228 (N_17228,N_16031,N_16762);
nor U17229 (N_17229,N_16031,N_16149);
nand U17230 (N_17230,N_16373,N_16580);
and U17231 (N_17231,N_16340,N_16391);
or U17232 (N_17232,N_16419,N_16621);
nor U17233 (N_17233,N_16242,N_16185);
and U17234 (N_17234,N_16645,N_16225);
nor U17235 (N_17235,N_16230,N_16699);
or U17236 (N_17236,N_16214,N_16437);
nand U17237 (N_17237,N_16195,N_16352);
and U17238 (N_17238,N_16240,N_16766);
and U17239 (N_17239,N_16377,N_16107);
nand U17240 (N_17240,N_16724,N_16319);
and U17241 (N_17241,N_16769,N_16496);
and U17242 (N_17242,N_16661,N_16520);
nand U17243 (N_17243,N_16488,N_16235);
and U17244 (N_17244,N_16635,N_16450);
xnor U17245 (N_17245,N_16443,N_16162);
and U17246 (N_17246,N_16574,N_16795);
nor U17247 (N_17247,N_16084,N_16502);
or U17248 (N_17248,N_16216,N_16724);
nand U17249 (N_17249,N_16489,N_16620);
nand U17250 (N_17250,N_16604,N_16297);
nand U17251 (N_17251,N_16598,N_16322);
and U17252 (N_17252,N_16762,N_16357);
and U17253 (N_17253,N_16632,N_16340);
or U17254 (N_17254,N_16664,N_16713);
and U17255 (N_17255,N_16326,N_16724);
and U17256 (N_17256,N_16406,N_16326);
nand U17257 (N_17257,N_16607,N_16410);
nor U17258 (N_17258,N_16088,N_16259);
nor U17259 (N_17259,N_16342,N_16431);
nand U17260 (N_17260,N_16567,N_16517);
nand U17261 (N_17261,N_16191,N_16390);
or U17262 (N_17262,N_16154,N_16384);
and U17263 (N_17263,N_16171,N_16349);
and U17264 (N_17264,N_16566,N_16178);
nor U17265 (N_17265,N_16054,N_16136);
nand U17266 (N_17266,N_16522,N_16013);
nand U17267 (N_17267,N_16005,N_16461);
nand U17268 (N_17268,N_16325,N_16713);
nor U17269 (N_17269,N_16549,N_16005);
nor U17270 (N_17270,N_16003,N_16555);
nand U17271 (N_17271,N_16403,N_16449);
and U17272 (N_17272,N_16605,N_16586);
nand U17273 (N_17273,N_16236,N_16556);
nand U17274 (N_17274,N_16409,N_16556);
and U17275 (N_17275,N_16699,N_16040);
and U17276 (N_17276,N_16329,N_16044);
nand U17277 (N_17277,N_16104,N_16517);
and U17278 (N_17278,N_16494,N_16575);
nand U17279 (N_17279,N_16381,N_16320);
or U17280 (N_17280,N_16051,N_16243);
or U17281 (N_17281,N_16734,N_16466);
nor U17282 (N_17282,N_16349,N_16701);
nor U17283 (N_17283,N_16641,N_16706);
and U17284 (N_17284,N_16220,N_16122);
nor U17285 (N_17285,N_16630,N_16115);
nand U17286 (N_17286,N_16164,N_16200);
nor U17287 (N_17287,N_16003,N_16706);
or U17288 (N_17288,N_16710,N_16709);
and U17289 (N_17289,N_16128,N_16000);
nor U17290 (N_17290,N_16131,N_16748);
nand U17291 (N_17291,N_16695,N_16428);
nand U17292 (N_17292,N_16041,N_16381);
nand U17293 (N_17293,N_16481,N_16515);
nand U17294 (N_17294,N_16309,N_16039);
or U17295 (N_17295,N_16639,N_16514);
and U17296 (N_17296,N_16061,N_16055);
or U17297 (N_17297,N_16742,N_16767);
nor U17298 (N_17298,N_16502,N_16407);
nand U17299 (N_17299,N_16172,N_16432);
and U17300 (N_17300,N_16621,N_16041);
nor U17301 (N_17301,N_16314,N_16509);
xnor U17302 (N_17302,N_16751,N_16749);
and U17303 (N_17303,N_16659,N_16394);
nor U17304 (N_17304,N_16041,N_16758);
nand U17305 (N_17305,N_16739,N_16756);
and U17306 (N_17306,N_16450,N_16419);
nor U17307 (N_17307,N_16052,N_16656);
nand U17308 (N_17308,N_16266,N_16032);
xor U17309 (N_17309,N_16384,N_16605);
nor U17310 (N_17310,N_16557,N_16689);
and U17311 (N_17311,N_16452,N_16021);
and U17312 (N_17312,N_16109,N_16331);
nor U17313 (N_17313,N_16303,N_16241);
or U17314 (N_17314,N_16439,N_16258);
or U17315 (N_17315,N_16668,N_16445);
xnor U17316 (N_17316,N_16711,N_16185);
and U17317 (N_17317,N_16475,N_16102);
nand U17318 (N_17318,N_16694,N_16586);
nand U17319 (N_17319,N_16173,N_16146);
and U17320 (N_17320,N_16725,N_16323);
nor U17321 (N_17321,N_16737,N_16200);
or U17322 (N_17322,N_16726,N_16721);
nand U17323 (N_17323,N_16779,N_16425);
nor U17324 (N_17324,N_16245,N_16048);
nor U17325 (N_17325,N_16077,N_16566);
or U17326 (N_17326,N_16754,N_16773);
and U17327 (N_17327,N_16076,N_16299);
nand U17328 (N_17328,N_16348,N_16245);
and U17329 (N_17329,N_16376,N_16121);
and U17330 (N_17330,N_16735,N_16041);
and U17331 (N_17331,N_16637,N_16286);
and U17332 (N_17332,N_16296,N_16463);
nand U17333 (N_17333,N_16681,N_16268);
nor U17334 (N_17334,N_16116,N_16776);
and U17335 (N_17335,N_16196,N_16599);
nor U17336 (N_17336,N_16401,N_16691);
nor U17337 (N_17337,N_16483,N_16773);
nor U17338 (N_17338,N_16612,N_16296);
and U17339 (N_17339,N_16623,N_16656);
and U17340 (N_17340,N_16107,N_16739);
and U17341 (N_17341,N_16434,N_16300);
and U17342 (N_17342,N_16631,N_16699);
or U17343 (N_17343,N_16678,N_16434);
and U17344 (N_17344,N_16161,N_16699);
nor U17345 (N_17345,N_16480,N_16794);
nor U17346 (N_17346,N_16156,N_16617);
and U17347 (N_17347,N_16747,N_16469);
nand U17348 (N_17348,N_16784,N_16399);
nand U17349 (N_17349,N_16532,N_16205);
or U17350 (N_17350,N_16707,N_16389);
nor U17351 (N_17351,N_16755,N_16402);
and U17352 (N_17352,N_16776,N_16697);
nor U17353 (N_17353,N_16590,N_16179);
nand U17354 (N_17354,N_16684,N_16716);
nand U17355 (N_17355,N_16532,N_16482);
nand U17356 (N_17356,N_16400,N_16348);
or U17357 (N_17357,N_16241,N_16334);
nor U17358 (N_17358,N_16447,N_16755);
nor U17359 (N_17359,N_16103,N_16392);
and U17360 (N_17360,N_16321,N_16209);
nor U17361 (N_17361,N_16047,N_16718);
nor U17362 (N_17362,N_16710,N_16767);
or U17363 (N_17363,N_16014,N_16652);
nor U17364 (N_17364,N_16671,N_16013);
nand U17365 (N_17365,N_16079,N_16488);
nor U17366 (N_17366,N_16761,N_16550);
or U17367 (N_17367,N_16671,N_16120);
nor U17368 (N_17368,N_16008,N_16004);
or U17369 (N_17369,N_16600,N_16493);
and U17370 (N_17370,N_16654,N_16559);
and U17371 (N_17371,N_16076,N_16085);
nor U17372 (N_17372,N_16312,N_16613);
and U17373 (N_17373,N_16188,N_16435);
xnor U17374 (N_17374,N_16096,N_16689);
nor U17375 (N_17375,N_16391,N_16444);
and U17376 (N_17376,N_16140,N_16636);
and U17377 (N_17377,N_16288,N_16725);
or U17378 (N_17378,N_16734,N_16700);
nand U17379 (N_17379,N_16174,N_16662);
and U17380 (N_17380,N_16158,N_16594);
or U17381 (N_17381,N_16089,N_16532);
nor U17382 (N_17382,N_16351,N_16399);
nand U17383 (N_17383,N_16169,N_16731);
nand U17384 (N_17384,N_16549,N_16383);
nor U17385 (N_17385,N_16655,N_16625);
nor U17386 (N_17386,N_16002,N_16010);
or U17387 (N_17387,N_16124,N_16281);
and U17388 (N_17388,N_16437,N_16594);
and U17389 (N_17389,N_16370,N_16470);
and U17390 (N_17390,N_16752,N_16691);
or U17391 (N_17391,N_16534,N_16170);
nand U17392 (N_17392,N_16127,N_16310);
nor U17393 (N_17393,N_16084,N_16523);
and U17394 (N_17394,N_16163,N_16585);
nor U17395 (N_17395,N_16569,N_16425);
or U17396 (N_17396,N_16640,N_16368);
and U17397 (N_17397,N_16409,N_16579);
nor U17398 (N_17398,N_16142,N_16461);
or U17399 (N_17399,N_16243,N_16441);
nor U17400 (N_17400,N_16478,N_16788);
nor U17401 (N_17401,N_16412,N_16748);
nor U17402 (N_17402,N_16509,N_16190);
and U17403 (N_17403,N_16716,N_16078);
nor U17404 (N_17404,N_16442,N_16764);
and U17405 (N_17405,N_16172,N_16152);
nor U17406 (N_17406,N_16036,N_16354);
or U17407 (N_17407,N_16562,N_16036);
nor U17408 (N_17408,N_16511,N_16057);
and U17409 (N_17409,N_16588,N_16063);
nand U17410 (N_17410,N_16530,N_16612);
nand U17411 (N_17411,N_16607,N_16397);
nand U17412 (N_17412,N_16276,N_16012);
and U17413 (N_17413,N_16368,N_16399);
and U17414 (N_17414,N_16467,N_16199);
and U17415 (N_17415,N_16664,N_16303);
nand U17416 (N_17416,N_16496,N_16542);
and U17417 (N_17417,N_16444,N_16513);
nor U17418 (N_17418,N_16700,N_16711);
or U17419 (N_17419,N_16798,N_16315);
and U17420 (N_17420,N_16635,N_16749);
or U17421 (N_17421,N_16374,N_16063);
nand U17422 (N_17422,N_16065,N_16448);
or U17423 (N_17423,N_16767,N_16107);
nand U17424 (N_17424,N_16776,N_16683);
and U17425 (N_17425,N_16753,N_16356);
and U17426 (N_17426,N_16376,N_16128);
nand U17427 (N_17427,N_16169,N_16412);
or U17428 (N_17428,N_16465,N_16097);
nor U17429 (N_17429,N_16103,N_16029);
and U17430 (N_17430,N_16086,N_16612);
or U17431 (N_17431,N_16174,N_16383);
or U17432 (N_17432,N_16704,N_16363);
and U17433 (N_17433,N_16402,N_16164);
nand U17434 (N_17434,N_16215,N_16213);
or U17435 (N_17435,N_16313,N_16624);
nor U17436 (N_17436,N_16727,N_16201);
or U17437 (N_17437,N_16787,N_16020);
nor U17438 (N_17438,N_16286,N_16147);
nand U17439 (N_17439,N_16460,N_16009);
nor U17440 (N_17440,N_16125,N_16538);
nor U17441 (N_17441,N_16386,N_16257);
and U17442 (N_17442,N_16295,N_16179);
nand U17443 (N_17443,N_16653,N_16155);
nor U17444 (N_17444,N_16452,N_16283);
nor U17445 (N_17445,N_16242,N_16254);
and U17446 (N_17446,N_16377,N_16179);
nor U17447 (N_17447,N_16106,N_16381);
nor U17448 (N_17448,N_16653,N_16507);
and U17449 (N_17449,N_16301,N_16235);
nor U17450 (N_17450,N_16211,N_16168);
nor U17451 (N_17451,N_16570,N_16407);
and U17452 (N_17452,N_16224,N_16203);
nand U17453 (N_17453,N_16407,N_16670);
and U17454 (N_17454,N_16514,N_16543);
nor U17455 (N_17455,N_16245,N_16400);
and U17456 (N_17456,N_16376,N_16633);
and U17457 (N_17457,N_16426,N_16217);
and U17458 (N_17458,N_16318,N_16216);
nor U17459 (N_17459,N_16356,N_16528);
or U17460 (N_17460,N_16227,N_16789);
and U17461 (N_17461,N_16563,N_16756);
or U17462 (N_17462,N_16151,N_16788);
nand U17463 (N_17463,N_16464,N_16624);
and U17464 (N_17464,N_16794,N_16060);
and U17465 (N_17465,N_16279,N_16488);
and U17466 (N_17466,N_16770,N_16478);
or U17467 (N_17467,N_16547,N_16157);
and U17468 (N_17468,N_16236,N_16385);
and U17469 (N_17469,N_16405,N_16382);
nor U17470 (N_17470,N_16569,N_16522);
nand U17471 (N_17471,N_16138,N_16247);
nand U17472 (N_17472,N_16585,N_16210);
and U17473 (N_17473,N_16199,N_16383);
nor U17474 (N_17474,N_16504,N_16355);
nor U17475 (N_17475,N_16379,N_16582);
and U17476 (N_17476,N_16445,N_16765);
or U17477 (N_17477,N_16152,N_16681);
or U17478 (N_17478,N_16122,N_16272);
and U17479 (N_17479,N_16532,N_16568);
nor U17480 (N_17480,N_16598,N_16291);
and U17481 (N_17481,N_16327,N_16682);
and U17482 (N_17482,N_16720,N_16438);
and U17483 (N_17483,N_16359,N_16182);
and U17484 (N_17484,N_16571,N_16086);
nand U17485 (N_17485,N_16374,N_16283);
nand U17486 (N_17486,N_16666,N_16438);
nand U17487 (N_17487,N_16645,N_16670);
nand U17488 (N_17488,N_16480,N_16373);
nand U17489 (N_17489,N_16180,N_16756);
nand U17490 (N_17490,N_16537,N_16668);
nand U17491 (N_17491,N_16313,N_16275);
or U17492 (N_17492,N_16189,N_16696);
or U17493 (N_17493,N_16201,N_16468);
xnor U17494 (N_17494,N_16424,N_16334);
or U17495 (N_17495,N_16363,N_16133);
or U17496 (N_17496,N_16428,N_16596);
nor U17497 (N_17497,N_16675,N_16398);
and U17498 (N_17498,N_16794,N_16213);
nor U17499 (N_17499,N_16319,N_16545);
nor U17500 (N_17500,N_16410,N_16505);
or U17501 (N_17501,N_16658,N_16568);
or U17502 (N_17502,N_16073,N_16631);
or U17503 (N_17503,N_16172,N_16427);
nor U17504 (N_17504,N_16320,N_16294);
nor U17505 (N_17505,N_16376,N_16123);
nor U17506 (N_17506,N_16012,N_16470);
and U17507 (N_17507,N_16168,N_16043);
or U17508 (N_17508,N_16417,N_16601);
nand U17509 (N_17509,N_16240,N_16271);
or U17510 (N_17510,N_16695,N_16671);
or U17511 (N_17511,N_16459,N_16056);
nand U17512 (N_17512,N_16105,N_16247);
or U17513 (N_17513,N_16409,N_16691);
and U17514 (N_17514,N_16163,N_16611);
nand U17515 (N_17515,N_16638,N_16212);
and U17516 (N_17516,N_16368,N_16301);
and U17517 (N_17517,N_16758,N_16054);
and U17518 (N_17518,N_16006,N_16201);
and U17519 (N_17519,N_16467,N_16133);
and U17520 (N_17520,N_16792,N_16362);
nand U17521 (N_17521,N_16377,N_16398);
or U17522 (N_17522,N_16502,N_16646);
nor U17523 (N_17523,N_16530,N_16230);
or U17524 (N_17524,N_16031,N_16093);
nand U17525 (N_17525,N_16531,N_16387);
nand U17526 (N_17526,N_16594,N_16254);
or U17527 (N_17527,N_16479,N_16205);
and U17528 (N_17528,N_16484,N_16463);
nand U17529 (N_17529,N_16406,N_16019);
nand U17530 (N_17530,N_16605,N_16277);
nand U17531 (N_17531,N_16493,N_16624);
nor U17532 (N_17532,N_16198,N_16454);
nor U17533 (N_17533,N_16593,N_16008);
nand U17534 (N_17534,N_16181,N_16456);
nand U17535 (N_17535,N_16058,N_16091);
and U17536 (N_17536,N_16445,N_16702);
nand U17537 (N_17537,N_16374,N_16124);
or U17538 (N_17538,N_16047,N_16611);
or U17539 (N_17539,N_16640,N_16275);
nor U17540 (N_17540,N_16695,N_16723);
nand U17541 (N_17541,N_16026,N_16495);
and U17542 (N_17542,N_16736,N_16506);
nor U17543 (N_17543,N_16470,N_16248);
nor U17544 (N_17544,N_16194,N_16565);
nand U17545 (N_17545,N_16342,N_16488);
nand U17546 (N_17546,N_16110,N_16413);
nand U17547 (N_17547,N_16221,N_16213);
or U17548 (N_17548,N_16752,N_16089);
nand U17549 (N_17549,N_16166,N_16478);
nand U17550 (N_17550,N_16701,N_16263);
nand U17551 (N_17551,N_16445,N_16259);
nor U17552 (N_17552,N_16602,N_16785);
or U17553 (N_17553,N_16193,N_16646);
or U17554 (N_17554,N_16745,N_16020);
nand U17555 (N_17555,N_16074,N_16685);
nand U17556 (N_17556,N_16154,N_16411);
or U17557 (N_17557,N_16186,N_16611);
nand U17558 (N_17558,N_16065,N_16147);
nor U17559 (N_17559,N_16030,N_16146);
and U17560 (N_17560,N_16371,N_16357);
or U17561 (N_17561,N_16348,N_16111);
or U17562 (N_17562,N_16230,N_16601);
nor U17563 (N_17563,N_16639,N_16447);
and U17564 (N_17564,N_16729,N_16195);
and U17565 (N_17565,N_16009,N_16301);
nand U17566 (N_17566,N_16089,N_16698);
and U17567 (N_17567,N_16613,N_16462);
or U17568 (N_17568,N_16308,N_16381);
or U17569 (N_17569,N_16008,N_16112);
nand U17570 (N_17570,N_16378,N_16430);
nor U17571 (N_17571,N_16558,N_16485);
or U17572 (N_17572,N_16140,N_16082);
and U17573 (N_17573,N_16346,N_16769);
and U17574 (N_17574,N_16286,N_16683);
nand U17575 (N_17575,N_16138,N_16094);
or U17576 (N_17576,N_16131,N_16753);
nand U17577 (N_17577,N_16700,N_16187);
nor U17578 (N_17578,N_16258,N_16446);
and U17579 (N_17579,N_16764,N_16364);
nor U17580 (N_17580,N_16436,N_16676);
or U17581 (N_17581,N_16248,N_16205);
and U17582 (N_17582,N_16493,N_16245);
nand U17583 (N_17583,N_16749,N_16023);
and U17584 (N_17584,N_16331,N_16496);
nor U17585 (N_17585,N_16302,N_16237);
nand U17586 (N_17586,N_16355,N_16076);
nor U17587 (N_17587,N_16520,N_16627);
and U17588 (N_17588,N_16726,N_16421);
and U17589 (N_17589,N_16162,N_16441);
nand U17590 (N_17590,N_16238,N_16480);
or U17591 (N_17591,N_16487,N_16400);
or U17592 (N_17592,N_16735,N_16670);
or U17593 (N_17593,N_16762,N_16192);
nor U17594 (N_17594,N_16775,N_16223);
or U17595 (N_17595,N_16683,N_16153);
or U17596 (N_17596,N_16044,N_16377);
and U17597 (N_17597,N_16576,N_16377);
nor U17598 (N_17598,N_16375,N_16386);
nand U17599 (N_17599,N_16279,N_16077);
and U17600 (N_17600,N_16894,N_17548);
nand U17601 (N_17601,N_17020,N_16863);
and U17602 (N_17602,N_16915,N_17064);
nor U17603 (N_17603,N_17093,N_16841);
nor U17604 (N_17604,N_16805,N_16869);
nand U17605 (N_17605,N_17431,N_16905);
and U17606 (N_17606,N_17155,N_16909);
nand U17607 (N_17607,N_17165,N_17081);
and U17608 (N_17608,N_17398,N_17530);
and U17609 (N_17609,N_17354,N_17090);
and U17610 (N_17610,N_17535,N_17433);
nand U17611 (N_17611,N_17338,N_17108);
nand U17612 (N_17612,N_17510,N_17067);
nand U17613 (N_17613,N_16828,N_17505);
nand U17614 (N_17614,N_17286,N_16997);
nor U17615 (N_17615,N_17170,N_17021);
nand U17616 (N_17616,N_17047,N_17477);
and U17617 (N_17617,N_17357,N_17464);
nand U17618 (N_17618,N_16867,N_16939);
nor U17619 (N_17619,N_16810,N_17340);
or U17620 (N_17620,N_17399,N_17308);
nand U17621 (N_17621,N_17434,N_16891);
or U17622 (N_17622,N_16975,N_16836);
or U17623 (N_17623,N_17251,N_17330);
nor U17624 (N_17624,N_17045,N_17305);
nor U17625 (N_17625,N_17373,N_17413);
nand U17626 (N_17626,N_17134,N_17185);
or U17627 (N_17627,N_17551,N_16953);
or U17628 (N_17628,N_17270,N_17011);
and U17629 (N_17629,N_17313,N_17521);
or U17630 (N_17630,N_17365,N_16801);
and U17631 (N_17631,N_17391,N_17219);
or U17632 (N_17632,N_17426,N_16812);
nand U17633 (N_17633,N_17417,N_17578);
nor U17634 (N_17634,N_17389,N_17010);
nor U17635 (N_17635,N_16901,N_17002);
and U17636 (N_17636,N_17545,N_17161);
and U17637 (N_17637,N_17440,N_17425);
or U17638 (N_17638,N_17173,N_17188);
nand U17639 (N_17639,N_17329,N_17175);
nor U17640 (N_17640,N_17544,N_17282);
or U17641 (N_17641,N_16806,N_17240);
nor U17642 (N_17642,N_17557,N_16896);
nor U17643 (N_17643,N_16946,N_17301);
or U17644 (N_17644,N_16897,N_16804);
nand U17645 (N_17645,N_17590,N_17446);
and U17646 (N_17646,N_17414,N_17350);
and U17647 (N_17647,N_17547,N_17005);
nand U17648 (N_17648,N_17153,N_17152);
and U17649 (N_17649,N_17517,N_17035);
or U17650 (N_17650,N_16999,N_17042);
or U17651 (N_17651,N_17129,N_17393);
nor U17652 (N_17652,N_17197,N_17546);
or U17653 (N_17653,N_16855,N_16852);
nor U17654 (N_17654,N_16994,N_16914);
or U17655 (N_17655,N_16960,N_17019);
nor U17656 (N_17656,N_17369,N_17052);
and U17657 (N_17657,N_17363,N_17043);
or U17658 (N_17658,N_17111,N_17589);
nand U17659 (N_17659,N_16974,N_17157);
and U17660 (N_17660,N_17407,N_16827);
or U17661 (N_17661,N_17514,N_17271);
and U17662 (N_17662,N_16954,N_17281);
nor U17663 (N_17663,N_17083,N_17349);
nor U17664 (N_17664,N_16964,N_17242);
or U17665 (N_17665,N_17495,N_17216);
and U17666 (N_17666,N_16961,N_17506);
nor U17667 (N_17667,N_17420,N_17563);
nor U17668 (N_17668,N_16814,N_17279);
and U17669 (N_17669,N_16957,N_17015);
nand U17670 (N_17670,N_16990,N_16979);
nand U17671 (N_17671,N_17125,N_16929);
or U17672 (N_17672,N_16969,N_17418);
or U17673 (N_17673,N_17117,N_17204);
nor U17674 (N_17674,N_17581,N_17124);
or U17675 (N_17675,N_17387,N_16923);
or U17676 (N_17676,N_17068,N_16919);
or U17677 (N_17677,N_17004,N_17381);
nor U17678 (N_17678,N_17296,N_17574);
nor U17679 (N_17679,N_17230,N_17226);
or U17680 (N_17680,N_17583,N_17362);
or U17681 (N_17681,N_16913,N_17238);
and U17682 (N_17682,N_17562,N_17411);
and U17683 (N_17683,N_17056,N_16985);
nor U17684 (N_17684,N_17423,N_17118);
or U17685 (N_17685,N_16887,N_17499);
and U17686 (N_17686,N_16912,N_17333);
nor U17687 (N_17687,N_17508,N_17497);
or U17688 (N_17688,N_17409,N_17579);
and U17689 (N_17689,N_17375,N_17335);
nand U17690 (N_17690,N_16924,N_17177);
nand U17691 (N_17691,N_17538,N_17038);
nor U17692 (N_17692,N_17202,N_17438);
nand U17693 (N_17693,N_17311,N_17353);
or U17694 (N_17694,N_16819,N_16821);
and U17695 (N_17695,N_17140,N_16983);
nor U17696 (N_17696,N_17540,N_16881);
xor U17697 (N_17697,N_17086,N_16883);
or U17698 (N_17698,N_16949,N_17323);
or U17699 (N_17699,N_17267,N_17364);
and U17700 (N_17700,N_17189,N_16968);
and U17701 (N_17701,N_16947,N_17284);
xnor U17702 (N_17702,N_17253,N_17077);
or U17703 (N_17703,N_17490,N_17156);
nor U17704 (N_17704,N_17534,N_17494);
nor U17705 (N_17705,N_17442,N_17231);
or U17706 (N_17706,N_16832,N_17303);
or U17707 (N_17707,N_16933,N_16966);
nand U17708 (N_17708,N_17080,N_17565);
nand U17709 (N_17709,N_17130,N_17057);
nand U17710 (N_17710,N_17037,N_17554);
nor U17711 (N_17711,N_17229,N_17537);
nor U17712 (N_17712,N_17332,N_17556);
or U17713 (N_17713,N_17082,N_17212);
nor U17714 (N_17714,N_17447,N_17249);
nor U17715 (N_17715,N_17151,N_17261);
and U17716 (N_17716,N_17314,N_17103);
or U17717 (N_17717,N_16856,N_17192);
nand U17718 (N_17718,N_16973,N_16996);
nand U17719 (N_17719,N_17050,N_16965);
or U17720 (N_17720,N_17444,N_17377);
nor U17721 (N_17721,N_17481,N_17529);
or U17722 (N_17722,N_16958,N_16831);
nor U17723 (N_17723,N_17078,N_17048);
and U17724 (N_17724,N_17098,N_17351);
and U17725 (N_17725,N_16847,N_17252);
or U17726 (N_17726,N_17123,N_16845);
nor U17727 (N_17727,N_17044,N_17553);
nand U17728 (N_17728,N_16921,N_17408);
nand U17729 (N_17729,N_17183,N_17254);
nor U17730 (N_17730,N_17588,N_17541);
or U17731 (N_17731,N_17273,N_17312);
or U17732 (N_17732,N_17450,N_16907);
or U17733 (N_17733,N_17516,N_17193);
nand U17734 (N_17734,N_16844,N_17033);
nand U17735 (N_17735,N_17030,N_17525);
and U17736 (N_17736,N_17594,N_17416);
nand U17737 (N_17737,N_17248,N_17009);
nand U17738 (N_17738,N_16925,N_16818);
and U17739 (N_17739,N_17327,N_16868);
or U17740 (N_17740,N_17582,N_17214);
and U17741 (N_17741,N_17572,N_16934);
and U17742 (N_17742,N_17451,N_17287);
and U17743 (N_17743,N_16858,N_17384);
and U17744 (N_17744,N_17424,N_16888);
or U17745 (N_17745,N_17519,N_17336);
nand U17746 (N_17746,N_17550,N_17470);
nand U17747 (N_17747,N_17441,N_17022);
nand U17748 (N_17748,N_17075,N_17055);
and U17749 (N_17749,N_17573,N_16916);
nor U17750 (N_17750,N_17070,N_16835);
nor U17751 (N_17751,N_17133,N_17000);
and U17752 (N_17752,N_17106,N_16864);
or U17753 (N_17753,N_17298,N_16943);
or U17754 (N_17754,N_16976,N_17127);
nand U17755 (N_17755,N_17272,N_17250);
and U17756 (N_17756,N_16865,N_17396);
nor U17757 (N_17757,N_17569,N_17536);
nand U17758 (N_17758,N_17302,N_17091);
or U17759 (N_17759,N_17243,N_16952);
and U17760 (N_17760,N_17207,N_17258);
nor U17761 (N_17761,N_17361,N_17315);
and U17762 (N_17762,N_16808,N_17454);
nor U17763 (N_17763,N_16991,N_17213);
nand U17764 (N_17764,N_16850,N_17241);
nor U17765 (N_17765,N_16816,N_16838);
nor U17766 (N_17766,N_17233,N_16935);
nor U17767 (N_17767,N_17345,N_17113);
or U17768 (N_17768,N_16911,N_17294);
or U17769 (N_17769,N_17162,N_17116);
nor U17770 (N_17770,N_17120,N_17085);
and U17771 (N_17771,N_17266,N_16826);
xor U17772 (N_17772,N_17568,N_16848);
and U17773 (N_17773,N_16842,N_17458);
or U17774 (N_17774,N_17386,N_16833);
nand U17775 (N_17775,N_17346,N_17491);
and U17776 (N_17776,N_17006,N_17184);
nor U17777 (N_17777,N_17208,N_17217);
nand U17778 (N_17778,N_17316,N_17366);
nor U17779 (N_17779,N_17533,N_17283);
nand U17780 (N_17780,N_17264,N_17360);
nand U17781 (N_17781,N_17419,N_16902);
and U17782 (N_17782,N_17370,N_17112);
nand U17783 (N_17783,N_16857,N_17092);
nor U17784 (N_17784,N_16959,N_17065);
or U17785 (N_17785,N_17235,N_17169);
nor U17786 (N_17786,N_17144,N_17257);
and U17787 (N_17787,N_16930,N_17147);
or U17788 (N_17788,N_17174,N_17527);
and U17789 (N_17789,N_16886,N_17379);
nand U17790 (N_17790,N_17017,N_17460);
and U17791 (N_17791,N_17228,N_17376);
and U17792 (N_17792,N_17058,N_17001);
or U17793 (N_17793,N_16803,N_17584);
and U17794 (N_17794,N_17392,N_16899);
nor U17795 (N_17795,N_16989,N_17559);
and U17796 (N_17796,N_16846,N_17522);
nor U17797 (N_17797,N_17580,N_17307);
nor U17798 (N_17798,N_16984,N_17060);
or U17799 (N_17799,N_17148,N_17164);
nand U17800 (N_17800,N_17181,N_17105);
and U17801 (N_17801,N_17088,N_17206);
and U17802 (N_17802,N_17437,N_17406);
nor U17803 (N_17803,N_16937,N_17131);
and U17804 (N_17804,N_17455,N_17263);
and U17805 (N_17805,N_17289,N_17593);
nor U17806 (N_17806,N_17100,N_17459);
or U17807 (N_17807,N_17107,N_17430);
or U17808 (N_17808,N_17475,N_17507);
and U17809 (N_17809,N_16840,N_17500);
nand U17810 (N_17810,N_17319,N_17049);
or U17811 (N_17811,N_17515,N_16876);
nor U17812 (N_17812,N_17154,N_17489);
or U17813 (N_17813,N_16938,N_17223);
nand U17814 (N_17814,N_17160,N_16922);
or U17815 (N_17815,N_17293,N_17528);
nor U17816 (N_17816,N_16906,N_17291);
and U17817 (N_17817,N_16843,N_17385);
or U17818 (N_17818,N_17415,N_16931);
and U17819 (N_17819,N_17520,N_17566);
nor U17820 (N_17820,N_16853,N_17278);
nand U17821 (N_17821,N_17585,N_17089);
nor U17822 (N_17822,N_17462,N_16870);
and U17823 (N_17823,N_16977,N_17421);
nor U17824 (N_17824,N_17026,N_16903);
or U17825 (N_17825,N_17542,N_16825);
or U17826 (N_17826,N_17403,N_17549);
or U17827 (N_17827,N_17150,N_17493);
and U17828 (N_17828,N_17472,N_17171);
nor U17829 (N_17829,N_17110,N_17115);
xor U17830 (N_17830,N_17136,N_16967);
and U17831 (N_17831,N_17275,N_17575);
nand U17832 (N_17832,N_17102,N_17180);
or U17833 (N_17833,N_17040,N_17095);
and U17834 (N_17834,N_17503,N_16940);
and U17835 (N_17835,N_17003,N_17269);
and U17836 (N_17836,N_17355,N_17167);
and U17837 (N_17837,N_17178,N_17059);
and U17838 (N_17838,N_16972,N_17555);
xor U17839 (N_17839,N_17288,N_17410);
nor U17840 (N_17840,N_17467,N_16978);
nand U17841 (N_17841,N_17039,N_17471);
nor U17842 (N_17842,N_17227,N_17496);
nor U17843 (N_17843,N_17591,N_16860);
nor U17844 (N_17844,N_17586,N_16908);
nand U17845 (N_17845,N_17378,N_16802);
or U17846 (N_17846,N_17318,N_16962);
nor U17847 (N_17847,N_16859,N_17259);
and U17848 (N_17848,N_17199,N_17331);
nand U17849 (N_17849,N_17244,N_17076);
nor U17850 (N_17850,N_17029,N_17492);
and U17851 (N_17851,N_17461,N_16932);
nor U17852 (N_17852,N_16874,N_16880);
and U17853 (N_17853,N_16820,N_16877);
nor U17854 (N_17854,N_17518,N_17448);
nor U17855 (N_17855,N_17439,N_17277);
or U17856 (N_17856,N_17334,N_17232);
and U17857 (N_17857,N_16884,N_17163);
nor U17858 (N_17858,N_16995,N_17394);
nand U17859 (N_17859,N_16817,N_17488);
or U17860 (N_17860,N_16834,N_16981);
nand U17861 (N_17861,N_17428,N_17066);
nor U17862 (N_17862,N_17074,N_17126);
nand U17863 (N_17863,N_16822,N_17402);
nand U17864 (N_17864,N_17201,N_17145);
nor U17865 (N_17865,N_17452,N_17560);
nor U17866 (N_17866,N_17342,N_17141);
nor U17867 (N_17867,N_16993,N_16854);
and U17868 (N_17868,N_17449,N_17036);
nor U17869 (N_17869,N_17187,N_17482);
nor U17870 (N_17870,N_17007,N_17457);
nand U17871 (N_17871,N_17501,N_17079);
nand U17872 (N_17872,N_17062,N_17096);
nand U17873 (N_17873,N_17051,N_17587);
nand U17874 (N_17874,N_17290,N_17466);
nand U17875 (N_17875,N_16879,N_17436);
nor U17876 (N_17876,N_16941,N_17328);
or U17877 (N_17877,N_17285,N_17498);
or U17878 (N_17878,N_16849,N_17485);
or U17879 (N_17879,N_17429,N_16988);
and U17880 (N_17880,N_16829,N_17337);
nand U17881 (N_17881,N_16927,N_17094);
or U17882 (N_17882,N_17143,N_17128);
nor U17883 (N_17883,N_16900,N_17324);
and U17884 (N_17884,N_17368,N_17225);
or U17885 (N_17885,N_16987,N_17073);
nor U17886 (N_17886,N_17432,N_16944);
nand U17887 (N_17887,N_17292,N_16873);
or U17888 (N_17888,N_17195,N_16878);
and U17889 (N_17889,N_16861,N_16971);
nor U17890 (N_17890,N_17028,N_17513);
nor U17891 (N_17891,N_17320,N_17310);
or U17892 (N_17892,N_17260,N_16811);
and U17893 (N_17893,N_16951,N_17237);
or U17894 (N_17894,N_16885,N_17325);
nor U17895 (N_17895,N_17061,N_17570);
nor U17896 (N_17896,N_17597,N_16809);
or U17897 (N_17897,N_17531,N_17158);
nand U17898 (N_17898,N_17599,N_17478);
nor U17899 (N_17899,N_17168,N_17159);
and U17900 (N_17900,N_17023,N_17063);
or U17901 (N_17901,N_16918,N_17191);
and U17902 (N_17902,N_17222,N_17256);
nand U17903 (N_17903,N_17194,N_17309);
nor U17904 (N_17904,N_17138,N_17139);
and U17905 (N_17905,N_17395,N_17255);
nor U17906 (N_17906,N_17018,N_17317);
nor U17907 (N_17907,N_16815,N_16926);
nor U17908 (N_17908,N_17046,N_16875);
or U17909 (N_17909,N_17179,N_17245);
nor U17910 (N_17910,N_16895,N_17109);
or U17911 (N_17911,N_16986,N_16936);
or U17912 (N_17912,N_16862,N_17072);
nor U17913 (N_17913,N_17476,N_16982);
nor U17914 (N_17914,N_17196,N_17479);
nor U17915 (N_17915,N_17347,N_17469);
nand U17916 (N_17916,N_17166,N_16830);
nor U17917 (N_17917,N_16898,N_17246);
nor U17918 (N_17918,N_17182,N_16970);
or U17919 (N_17919,N_17119,N_17262);
nor U17920 (N_17920,N_16892,N_17247);
and U17921 (N_17921,N_17224,N_17146);
or U17922 (N_17922,N_17465,N_16839);
and U17923 (N_17923,N_17211,N_17132);
nand U17924 (N_17924,N_16866,N_17084);
nand U17925 (N_17925,N_17343,N_17567);
and U17926 (N_17926,N_17380,N_17435);
and U17927 (N_17927,N_17234,N_16950);
or U17928 (N_17928,N_17512,N_17382);
nand U17929 (N_17929,N_17504,N_17532);
or U17930 (N_17930,N_17304,N_17473);
nor U17931 (N_17931,N_17405,N_16904);
and U17932 (N_17932,N_17480,N_17592);
nand U17933 (N_17933,N_17558,N_17215);
nor U17934 (N_17934,N_17321,N_16823);
nand U17935 (N_17935,N_16942,N_17295);
nand U17936 (N_17936,N_17268,N_17552);
nor U17937 (N_17937,N_17099,N_17390);
or U17938 (N_17938,N_17571,N_17221);
nor U17939 (N_17939,N_16824,N_17326);
and U17940 (N_17940,N_17486,N_17524);
nor U17941 (N_17941,N_17265,N_17135);
nand U17942 (N_17942,N_17356,N_17359);
and U17943 (N_17943,N_17299,N_16917);
nand U17944 (N_17944,N_17383,N_17012);
or U17945 (N_17945,N_17463,N_17236);
nand U17946 (N_17946,N_17210,N_17577);
or U17947 (N_17947,N_17203,N_16893);
xor U17948 (N_17948,N_17374,N_17031);
nand U17949 (N_17949,N_17422,N_17027);
or U17950 (N_17950,N_17596,N_17509);
or U17951 (N_17951,N_17025,N_17564);
nor U17952 (N_17952,N_17348,N_17276);
nor U17953 (N_17953,N_17474,N_17200);
and U17954 (N_17954,N_17322,N_17300);
and U17955 (N_17955,N_17190,N_16871);
and U17956 (N_17956,N_17397,N_17352);
or U17957 (N_17957,N_17523,N_17024);
nor U17958 (N_17958,N_16800,N_17539);
nand U17959 (N_17959,N_17511,N_17032);
or U17960 (N_17960,N_17186,N_17595);
nor U17961 (N_17961,N_17137,N_17014);
nand U17962 (N_17962,N_17205,N_16920);
and U17963 (N_17963,N_17487,N_16851);
and U17964 (N_17964,N_17274,N_17388);
nor U17965 (N_17965,N_16890,N_16948);
and U17966 (N_17966,N_16945,N_17502);
xnor U17967 (N_17967,N_17453,N_17114);
nor U17968 (N_17968,N_17404,N_17209);
nor U17969 (N_17969,N_17339,N_17483);
nand U17970 (N_17970,N_17543,N_16889);
or U17971 (N_17971,N_17053,N_17054);
and U17972 (N_17972,N_17445,N_17401);
or U17973 (N_17973,N_17097,N_17598);
nand U17974 (N_17974,N_16882,N_17121);
nand U17975 (N_17975,N_17372,N_17358);
and U17976 (N_17976,N_16992,N_17013);
or U17977 (N_17977,N_17427,N_17069);
or U17978 (N_17978,N_17087,N_16998);
nand U17979 (N_17979,N_17561,N_16813);
or U17980 (N_17980,N_17239,N_17198);
nand U17981 (N_17981,N_16963,N_17456);
xor U17982 (N_17982,N_17412,N_16807);
and U17983 (N_17983,N_17172,N_17297);
and U17984 (N_17984,N_17220,N_16872);
nand U17985 (N_17985,N_17367,N_16956);
or U17986 (N_17986,N_17218,N_17142);
or U17987 (N_17987,N_17526,N_17101);
or U17988 (N_17988,N_16980,N_17484);
nor U17989 (N_17989,N_17400,N_17041);
or U17990 (N_17990,N_17443,N_17280);
nand U17991 (N_17991,N_16928,N_17341);
nand U17992 (N_17992,N_17344,N_17149);
nand U17993 (N_17993,N_17576,N_17104);
nor U17994 (N_17994,N_17122,N_17371);
nor U17995 (N_17995,N_17016,N_17176);
nand U17996 (N_17996,N_16910,N_16837);
nand U17997 (N_17997,N_17071,N_17034);
or U17998 (N_17998,N_16955,N_17468);
nor U17999 (N_17999,N_17306,N_17008);
nor U18000 (N_18000,N_17471,N_17519);
or U18001 (N_18001,N_17328,N_17351);
nor U18002 (N_18002,N_17140,N_16976);
and U18003 (N_18003,N_17137,N_17195);
and U18004 (N_18004,N_17438,N_17535);
and U18005 (N_18005,N_16938,N_17337);
or U18006 (N_18006,N_17382,N_16984);
or U18007 (N_18007,N_17182,N_17366);
nand U18008 (N_18008,N_17185,N_17147);
nor U18009 (N_18009,N_17322,N_17210);
and U18010 (N_18010,N_17366,N_17370);
or U18011 (N_18011,N_17143,N_17479);
or U18012 (N_18012,N_16937,N_16971);
nor U18013 (N_18013,N_17158,N_16858);
or U18014 (N_18014,N_16927,N_17214);
and U18015 (N_18015,N_16926,N_17526);
or U18016 (N_18016,N_16955,N_16810);
and U18017 (N_18017,N_17311,N_16847);
and U18018 (N_18018,N_16967,N_17323);
or U18019 (N_18019,N_17510,N_17113);
nor U18020 (N_18020,N_17231,N_17514);
and U18021 (N_18021,N_17445,N_17385);
or U18022 (N_18022,N_17275,N_17019);
nand U18023 (N_18023,N_17078,N_17464);
nand U18024 (N_18024,N_17061,N_17139);
or U18025 (N_18025,N_17203,N_17181);
nand U18026 (N_18026,N_16954,N_17386);
and U18027 (N_18027,N_17480,N_17134);
nand U18028 (N_18028,N_16867,N_17456);
or U18029 (N_18029,N_17570,N_17436);
nand U18030 (N_18030,N_17158,N_17302);
and U18031 (N_18031,N_17469,N_16934);
and U18032 (N_18032,N_17099,N_17231);
nor U18033 (N_18033,N_17223,N_17160);
nand U18034 (N_18034,N_17369,N_17095);
and U18035 (N_18035,N_17303,N_17551);
or U18036 (N_18036,N_17494,N_17591);
and U18037 (N_18037,N_17338,N_17205);
nand U18038 (N_18038,N_17408,N_17505);
or U18039 (N_18039,N_17258,N_17276);
and U18040 (N_18040,N_17051,N_17350);
and U18041 (N_18041,N_16940,N_17483);
or U18042 (N_18042,N_16963,N_17329);
and U18043 (N_18043,N_17133,N_17404);
nor U18044 (N_18044,N_17515,N_16861);
or U18045 (N_18045,N_17220,N_17147);
and U18046 (N_18046,N_17325,N_17123);
and U18047 (N_18047,N_16959,N_17172);
or U18048 (N_18048,N_17470,N_17469);
nand U18049 (N_18049,N_16821,N_17175);
nand U18050 (N_18050,N_17480,N_17418);
nor U18051 (N_18051,N_17450,N_17150);
nor U18052 (N_18052,N_16975,N_17538);
and U18053 (N_18053,N_17325,N_16877);
and U18054 (N_18054,N_17284,N_17370);
or U18055 (N_18055,N_17491,N_17594);
and U18056 (N_18056,N_17196,N_17014);
nor U18057 (N_18057,N_17403,N_16880);
or U18058 (N_18058,N_17530,N_17585);
or U18059 (N_18059,N_17481,N_17087);
nor U18060 (N_18060,N_17210,N_17506);
or U18061 (N_18061,N_17123,N_17249);
or U18062 (N_18062,N_17103,N_17209);
nand U18063 (N_18063,N_16963,N_17375);
and U18064 (N_18064,N_17270,N_16882);
nor U18065 (N_18065,N_17239,N_16823);
or U18066 (N_18066,N_17246,N_16880);
nor U18067 (N_18067,N_16892,N_17420);
or U18068 (N_18068,N_17143,N_17017);
and U18069 (N_18069,N_17138,N_17552);
or U18070 (N_18070,N_16852,N_16902);
xor U18071 (N_18071,N_17071,N_17499);
or U18072 (N_18072,N_17175,N_17520);
and U18073 (N_18073,N_17270,N_17231);
or U18074 (N_18074,N_17007,N_16931);
nand U18075 (N_18075,N_17297,N_16831);
nor U18076 (N_18076,N_17313,N_17216);
nand U18077 (N_18077,N_17205,N_17579);
and U18078 (N_18078,N_16879,N_16887);
nor U18079 (N_18079,N_16836,N_16823);
nor U18080 (N_18080,N_17545,N_17579);
and U18081 (N_18081,N_17477,N_17481);
and U18082 (N_18082,N_17287,N_17081);
nor U18083 (N_18083,N_17421,N_16897);
nor U18084 (N_18084,N_17473,N_16808);
and U18085 (N_18085,N_17343,N_17056);
and U18086 (N_18086,N_17076,N_16807);
and U18087 (N_18087,N_17479,N_17409);
nor U18088 (N_18088,N_17167,N_17409);
nor U18089 (N_18089,N_17080,N_17562);
or U18090 (N_18090,N_17397,N_17538);
nor U18091 (N_18091,N_17173,N_17132);
nand U18092 (N_18092,N_17331,N_17229);
or U18093 (N_18093,N_16967,N_17178);
or U18094 (N_18094,N_17114,N_17583);
nor U18095 (N_18095,N_17378,N_17115);
xnor U18096 (N_18096,N_16977,N_16835);
and U18097 (N_18097,N_17379,N_16875);
and U18098 (N_18098,N_17173,N_17398);
nor U18099 (N_18099,N_17468,N_17456);
nor U18100 (N_18100,N_17287,N_16947);
nand U18101 (N_18101,N_17465,N_17482);
nand U18102 (N_18102,N_17449,N_17197);
nor U18103 (N_18103,N_17076,N_16906);
nand U18104 (N_18104,N_16823,N_17205);
or U18105 (N_18105,N_17419,N_17256);
and U18106 (N_18106,N_16896,N_17523);
or U18107 (N_18107,N_17477,N_16880);
nor U18108 (N_18108,N_17031,N_17253);
nand U18109 (N_18109,N_16854,N_17390);
and U18110 (N_18110,N_17325,N_16937);
or U18111 (N_18111,N_17427,N_17362);
or U18112 (N_18112,N_16902,N_16800);
nand U18113 (N_18113,N_17596,N_17105);
nand U18114 (N_18114,N_17030,N_17018);
nor U18115 (N_18115,N_16941,N_17534);
nand U18116 (N_18116,N_17126,N_17236);
nand U18117 (N_18117,N_17235,N_17061);
nor U18118 (N_18118,N_17263,N_17599);
nand U18119 (N_18119,N_16999,N_17352);
nand U18120 (N_18120,N_17563,N_17520);
or U18121 (N_18121,N_17094,N_17361);
and U18122 (N_18122,N_16902,N_17188);
or U18123 (N_18123,N_17279,N_17432);
nand U18124 (N_18124,N_17425,N_17030);
or U18125 (N_18125,N_16974,N_17467);
or U18126 (N_18126,N_17072,N_16819);
or U18127 (N_18127,N_17106,N_17394);
or U18128 (N_18128,N_17576,N_16890);
nor U18129 (N_18129,N_17030,N_16812);
nor U18130 (N_18130,N_17037,N_17547);
and U18131 (N_18131,N_17368,N_17121);
nor U18132 (N_18132,N_17266,N_16981);
nand U18133 (N_18133,N_17202,N_17220);
nand U18134 (N_18134,N_17107,N_16975);
and U18135 (N_18135,N_17035,N_17520);
nand U18136 (N_18136,N_17015,N_17188);
nand U18137 (N_18137,N_16817,N_17069);
or U18138 (N_18138,N_17267,N_17233);
nand U18139 (N_18139,N_16935,N_17153);
nand U18140 (N_18140,N_17536,N_16821);
nand U18141 (N_18141,N_16981,N_17367);
and U18142 (N_18142,N_17063,N_17198);
nand U18143 (N_18143,N_17320,N_17286);
nand U18144 (N_18144,N_17331,N_17441);
nand U18145 (N_18145,N_17272,N_17369);
nor U18146 (N_18146,N_16933,N_17343);
or U18147 (N_18147,N_17576,N_16968);
nand U18148 (N_18148,N_17430,N_17029);
nand U18149 (N_18149,N_17493,N_17499);
nor U18150 (N_18150,N_17096,N_17352);
nand U18151 (N_18151,N_17414,N_17364);
nand U18152 (N_18152,N_16815,N_17431);
and U18153 (N_18153,N_16887,N_16909);
nand U18154 (N_18154,N_17063,N_17238);
nor U18155 (N_18155,N_17040,N_17182);
and U18156 (N_18156,N_17328,N_16904);
nor U18157 (N_18157,N_16910,N_17364);
nand U18158 (N_18158,N_16803,N_17165);
and U18159 (N_18159,N_17075,N_16862);
nor U18160 (N_18160,N_17175,N_16844);
and U18161 (N_18161,N_17369,N_17068);
nand U18162 (N_18162,N_17491,N_17362);
and U18163 (N_18163,N_17199,N_17181);
nand U18164 (N_18164,N_17588,N_17355);
nor U18165 (N_18165,N_17255,N_17245);
and U18166 (N_18166,N_16986,N_17114);
nor U18167 (N_18167,N_17523,N_17100);
nand U18168 (N_18168,N_17363,N_17031);
nand U18169 (N_18169,N_17345,N_17076);
and U18170 (N_18170,N_17404,N_17286);
and U18171 (N_18171,N_16934,N_17180);
nand U18172 (N_18172,N_17470,N_17343);
and U18173 (N_18173,N_17256,N_17129);
nor U18174 (N_18174,N_17444,N_16967);
nand U18175 (N_18175,N_17053,N_17171);
and U18176 (N_18176,N_16830,N_17239);
or U18177 (N_18177,N_16909,N_17584);
nor U18178 (N_18178,N_17426,N_16856);
and U18179 (N_18179,N_16915,N_17101);
nand U18180 (N_18180,N_16987,N_16941);
and U18181 (N_18181,N_17558,N_17454);
and U18182 (N_18182,N_17204,N_17490);
nor U18183 (N_18183,N_16811,N_17018);
or U18184 (N_18184,N_17005,N_17292);
nand U18185 (N_18185,N_17451,N_17079);
or U18186 (N_18186,N_17394,N_17056);
nor U18187 (N_18187,N_17188,N_17493);
or U18188 (N_18188,N_17224,N_16898);
nand U18189 (N_18189,N_17502,N_17464);
or U18190 (N_18190,N_17204,N_17356);
nand U18191 (N_18191,N_17382,N_17117);
nand U18192 (N_18192,N_17384,N_17546);
and U18193 (N_18193,N_17398,N_17283);
or U18194 (N_18194,N_17210,N_17588);
or U18195 (N_18195,N_17414,N_16825);
nand U18196 (N_18196,N_17005,N_17414);
nand U18197 (N_18197,N_17334,N_17092);
nor U18198 (N_18198,N_17538,N_17035);
and U18199 (N_18199,N_17213,N_16802);
nor U18200 (N_18200,N_17569,N_16915);
nor U18201 (N_18201,N_17328,N_17218);
or U18202 (N_18202,N_17175,N_16914);
nor U18203 (N_18203,N_17019,N_17108);
and U18204 (N_18204,N_17415,N_16950);
and U18205 (N_18205,N_17010,N_17251);
nor U18206 (N_18206,N_17143,N_17309);
nor U18207 (N_18207,N_17284,N_17577);
and U18208 (N_18208,N_17007,N_17519);
or U18209 (N_18209,N_16853,N_17214);
or U18210 (N_18210,N_17398,N_17464);
nor U18211 (N_18211,N_16854,N_17040);
and U18212 (N_18212,N_16955,N_16892);
nor U18213 (N_18213,N_16920,N_17293);
nor U18214 (N_18214,N_17402,N_17186);
and U18215 (N_18215,N_16851,N_17401);
or U18216 (N_18216,N_17095,N_17454);
or U18217 (N_18217,N_17598,N_17232);
nand U18218 (N_18218,N_16940,N_17278);
and U18219 (N_18219,N_17587,N_17512);
and U18220 (N_18220,N_17254,N_17491);
and U18221 (N_18221,N_17185,N_17393);
and U18222 (N_18222,N_17111,N_16988);
nand U18223 (N_18223,N_16818,N_16809);
or U18224 (N_18224,N_17538,N_17469);
nor U18225 (N_18225,N_17006,N_17559);
and U18226 (N_18226,N_17197,N_17261);
or U18227 (N_18227,N_17311,N_17512);
nand U18228 (N_18228,N_17513,N_17038);
or U18229 (N_18229,N_17469,N_17392);
nor U18230 (N_18230,N_17101,N_17413);
or U18231 (N_18231,N_17475,N_17281);
nor U18232 (N_18232,N_17053,N_17233);
or U18233 (N_18233,N_17018,N_17481);
nand U18234 (N_18234,N_17215,N_17462);
nor U18235 (N_18235,N_17411,N_17330);
nand U18236 (N_18236,N_17306,N_16882);
nor U18237 (N_18237,N_17249,N_17121);
xor U18238 (N_18238,N_17423,N_17517);
or U18239 (N_18239,N_17246,N_17452);
nor U18240 (N_18240,N_17032,N_16876);
nor U18241 (N_18241,N_16945,N_17190);
or U18242 (N_18242,N_16872,N_17551);
nor U18243 (N_18243,N_17134,N_17165);
or U18244 (N_18244,N_17214,N_17502);
nor U18245 (N_18245,N_17575,N_17365);
nand U18246 (N_18246,N_16930,N_17374);
and U18247 (N_18247,N_17283,N_16850);
and U18248 (N_18248,N_17132,N_17197);
and U18249 (N_18249,N_17274,N_17467);
or U18250 (N_18250,N_17414,N_17521);
nor U18251 (N_18251,N_16878,N_17569);
nor U18252 (N_18252,N_17373,N_17448);
or U18253 (N_18253,N_16894,N_16878);
nor U18254 (N_18254,N_17205,N_17379);
and U18255 (N_18255,N_17279,N_17119);
nand U18256 (N_18256,N_17506,N_17384);
nor U18257 (N_18257,N_17071,N_16898);
and U18258 (N_18258,N_17437,N_17533);
nor U18259 (N_18259,N_17336,N_17287);
or U18260 (N_18260,N_17511,N_16944);
nor U18261 (N_18261,N_17165,N_17404);
or U18262 (N_18262,N_16951,N_17165);
nor U18263 (N_18263,N_16973,N_17439);
and U18264 (N_18264,N_16965,N_17205);
and U18265 (N_18265,N_17495,N_17512);
or U18266 (N_18266,N_17367,N_17023);
or U18267 (N_18267,N_17261,N_17316);
nand U18268 (N_18268,N_16966,N_17048);
nand U18269 (N_18269,N_16983,N_17338);
xnor U18270 (N_18270,N_16883,N_17335);
nor U18271 (N_18271,N_17495,N_16999);
and U18272 (N_18272,N_17069,N_16991);
nor U18273 (N_18273,N_17464,N_17034);
nand U18274 (N_18274,N_17083,N_17416);
and U18275 (N_18275,N_16959,N_17176);
or U18276 (N_18276,N_16815,N_17440);
and U18277 (N_18277,N_17101,N_17340);
and U18278 (N_18278,N_17332,N_16873);
or U18279 (N_18279,N_16901,N_17003);
and U18280 (N_18280,N_17143,N_17319);
nand U18281 (N_18281,N_17277,N_17159);
or U18282 (N_18282,N_17554,N_16803);
nand U18283 (N_18283,N_16856,N_17487);
and U18284 (N_18284,N_17317,N_17432);
or U18285 (N_18285,N_17045,N_17465);
nor U18286 (N_18286,N_17038,N_17170);
nand U18287 (N_18287,N_17541,N_17045);
and U18288 (N_18288,N_17137,N_17113);
nand U18289 (N_18289,N_17368,N_17551);
nand U18290 (N_18290,N_17127,N_16867);
nor U18291 (N_18291,N_16862,N_17203);
nor U18292 (N_18292,N_17195,N_17016);
nor U18293 (N_18293,N_17173,N_17475);
nand U18294 (N_18294,N_16825,N_17225);
nand U18295 (N_18295,N_17524,N_17136);
nor U18296 (N_18296,N_17218,N_17085);
nor U18297 (N_18297,N_17218,N_17480);
nor U18298 (N_18298,N_17388,N_17024);
and U18299 (N_18299,N_17084,N_17040);
or U18300 (N_18300,N_17137,N_16866);
or U18301 (N_18301,N_17167,N_16949);
or U18302 (N_18302,N_17251,N_17421);
and U18303 (N_18303,N_17254,N_17184);
or U18304 (N_18304,N_17342,N_17123);
and U18305 (N_18305,N_17151,N_16901);
nand U18306 (N_18306,N_17569,N_17036);
nand U18307 (N_18307,N_17225,N_16912);
or U18308 (N_18308,N_17430,N_17128);
nor U18309 (N_18309,N_17316,N_17003);
nor U18310 (N_18310,N_17331,N_17360);
or U18311 (N_18311,N_16805,N_17403);
or U18312 (N_18312,N_16915,N_17438);
nand U18313 (N_18313,N_17150,N_17123);
nor U18314 (N_18314,N_17350,N_17098);
nand U18315 (N_18315,N_17195,N_17363);
and U18316 (N_18316,N_17488,N_17168);
or U18317 (N_18317,N_17525,N_17443);
or U18318 (N_18318,N_17121,N_17450);
nand U18319 (N_18319,N_17387,N_17425);
nor U18320 (N_18320,N_16947,N_17204);
or U18321 (N_18321,N_17083,N_17313);
nor U18322 (N_18322,N_17538,N_17507);
nand U18323 (N_18323,N_17141,N_17343);
and U18324 (N_18324,N_16994,N_16831);
and U18325 (N_18325,N_17316,N_17597);
nor U18326 (N_18326,N_17195,N_17516);
or U18327 (N_18327,N_17480,N_16942);
nor U18328 (N_18328,N_17453,N_16911);
nand U18329 (N_18329,N_17244,N_17022);
nor U18330 (N_18330,N_17179,N_17156);
and U18331 (N_18331,N_17255,N_17439);
nor U18332 (N_18332,N_17116,N_17358);
nand U18333 (N_18333,N_17369,N_17380);
nand U18334 (N_18334,N_17011,N_17266);
nand U18335 (N_18335,N_16998,N_17115);
nor U18336 (N_18336,N_17155,N_16842);
nor U18337 (N_18337,N_16975,N_17030);
nor U18338 (N_18338,N_17153,N_17332);
nor U18339 (N_18339,N_17028,N_17338);
nand U18340 (N_18340,N_17084,N_16815);
and U18341 (N_18341,N_17003,N_17089);
nand U18342 (N_18342,N_17200,N_17217);
nor U18343 (N_18343,N_17375,N_17249);
and U18344 (N_18344,N_17445,N_17342);
nor U18345 (N_18345,N_17006,N_17385);
or U18346 (N_18346,N_17017,N_16986);
xor U18347 (N_18347,N_17081,N_17190);
nand U18348 (N_18348,N_17581,N_16901);
or U18349 (N_18349,N_17308,N_17544);
nor U18350 (N_18350,N_17252,N_17569);
nand U18351 (N_18351,N_16817,N_17068);
or U18352 (N_18352,N_17285,N_17065);
or U18353 (N_18353,N_17075,N_17337);
or U18354 (N_18354,N_16914,N_17138);
nor U18355 (N_18355,N_16948,N_17308);
nand U18356 (N_18356,N_17451,N_17384);
and U18357 (N_18357,N_17524,N_17399);
and U18358 (N_18358,N_17399,N_17572);
or U18359 (N_18359,N_17595,N_16831);
nand U18360 (N_18360,N_17170,N_17079);
or U18361 (N_18361,N_16832,N_17482);
nor U18362 (N_18362,N_17369,N_16809);
or U18363 (N_18363,N_17236,N_17430);
and U18364 (N_18364,N_17038,N_16834);
nand U18365 (N_18365,N_17575,N_17593);
and U18366 (N_18366,N_17147,N_16909);
or U18367 (N_18367,N_17391,N_17305);
nand U18368 (N_18368,N_17003,N_17520);
nand U18369 (N_18369,N_17483,N_16851);
nand U18370 (N_18370,N_17124,N_17348);
or U18371 (N_18371,N_17470,N_17357);
nand U18372 (N_18372,N_17257,N_17128);
nand U18373 (N_18373,N_17190,N_17183);
and U18374 (N_18374,N_17117,N_17192);
nand U18375 (N_18375,N_16994,N_17191);
nand U18376 (N_18376,N_17223,N_16942);
nor U18377 (N_18377,N_17086,N_17320);
or U18378 (N_18378,N_16973,N_17435);
and U18379 (N_18379,N_17449,N_17446);
and U18380 (N_18380,N_17418,N_16805);
and U18381 (N_18381,N_17104,N_17455);
nand U18382 (N_18382,N_17146,N_16859);
and U18383 (N_18383,N_16910,N_17478);
or U18384 (N_18384,N_17522,N_17104);
and U18385 (N_18385,N_17385,N_17519);
and U18386 (N_18386,N_17036,N_17046);
nor U18387 (N_18387,N_17323,N_17069);
and U18388 (N_18388,N_17437,N_17482);
or U18389 (N_18389,N_17561,N_17203);
nor U18390 (N_18390,N_17117,N_17143);
or U18391 (N_18391,N_17488,N_17495);
and U18392 (N_18392,N_16974,N_17305);
nor U18393 (N_18393,N_17329,N_17023);
and U18394 (N_18394,N_17372,N_17183);
or U18395 (N_18395,N_17524,N_17471);
nor U18396 (N_18396,N_16927,N_17455);
nand U18397 (N_18397,N_17292,N_17018);
nor U18398 (N_18398,N_16906,N_17193);
nand U18399 (N_18399,N_17288,N_17189);
and U18400 (N_18400,N_17964,N_17995);
and U18401 (N_18401,N_17919,N_17647);
and U18402 (N_18402,N_17634,N_17806);
nor U18403 (N_18403,N_17715,N_17688);
nand U18404 (N_18404,N_17887,N_18016);
nand U18405 (N_18405,N_18387,N_17819);
nor U18406 (N_18406,N_18166,N_18118);
and U18407 (N_18407,N_17623,N_17920);
nor U18408 (N_18408,N_17693,N_17968);
nand U18409 (N_18409,N_17924,N_17639);
nand U18410 (N_18410,N_17845,N_17657);
or U18411 (N_18411,N_17949,N_17654);
or U18412 (N_18412,N_18019,N_17916);
nand U18413 (N_18413,N_18229,N_17703);
and U18414 (N_18414,N_18033,N_17977);
and U18415 (N_18415,N_18189,N_18073);
nand U18416 (N_18416,N_17840,N_17954);
nor U18417 (N_18417,N_18060,N_17883);
and U18418 (N_18418,N_18212,N_17926);
nand U18419 (N_18419,N_17874,N_18323);
nor U18420 (N_18420,N_18059,N_18285);
and U18421 (N_18421,N_18273,N_17791);
nor U18422 (N_18422,N_18268,N_18025);
or U18423 (N_18423,N_17927,N_17979);
nand U18424 (N_18424,N_17793,N_17700);
or U18425 (N_18425,N_17865,N_18051);
and U18426 (N_18426,N_17767,N_17910);
and U18427 (N_18427,N_17640,N_18041);
nor U18428 (N_18428,N_18047,N_17904);
or U18429 (N_18429,N_18175,N_17690);
and U18430 (N_18430,N_17712,N_18252);
or U18431 (N_18431,N_18356,N_17875);
nor U18432 (N_18432,N_17808,N_17967);
and U18433 (N_18433,N_17901,N_18042);
and U18434 (N_18434,N_17831,N_17627);
and U18435 (N_18435,N_18143,N_18005);
nand U18436 (N_18436,N_18048,N_17776);
and U18437 (N_18437,N_18030,N_18181);
nor U18438 (N_18438,N_18104,N_18077);
nand U18439 (N_18439,N_17983,N_18319);
and U18440 (N_18440,N_17706,N_17822);
nor U18441 (N_18441,N_18293,N_17947);
nor U18442 (N_18442,N_17721,N_18138);
nand U18443 (N_18443,N_17679,N_17913);
and U18444 (N_18444,N_17827,N_18239);
and U18445 (N_18445,N_17963,N_18271);
nor U18446 (N_18446,N_17873,N_17771);
or U18447 (N_18447,N_18053,N_18159);
nor U18448 (N_18448,N_17992,N_18313);
or U18449 (N_18449,N_18103,N_17761);
nand U18450 (N_18450,N_17989,N_17660);
or U18451 (N_18451,N_18262,N_17600);
and U18452 (N_18452,N_18187,N_18330);
or U18453 (N_18453,N_17773,N_18193);
and U18454 (N_18454,N_18378,N_18282);
nor U18455 (N_18455,N_17757,N_17998);
nor U18456 (N_18456,N_17820,N_17815);
nor U18457 (N_18457,N_18327,N_18375);
or U18458 (N_18458,N_17956,N_18297);
nor U18459 (N_18459,N_18287,N_17922);
nor U18460 (N_18460,N_18192,N_17974);
and U18461 (N_18461,N_18312,N_17925);
and U18462 (N_18462,N_18288,N_17689);
nand U18463 (N_18463,N_18370,N_17986);
and U18464 (N_18464,N_17809,N_17710);
or U18465 (N_18465,N_17980,N_18004);
or U18466 (N_18466,N_18217,N_18165);
nor U18467 (N_18467,N_18055,N_18334);
nand U18468 (N_18468,N_18173,N_18219);
and U18469 (N_18469,N_17948,N_17976);
nand U18470 (N_18470,N_17718,N_17866);
and U18471 (N_18471,N_18183,N_18379);
or U18472 (N_18472,N_17663,N_18160);
or U18473 (N_18473,N_17928,N_18167);
or U18474 (N_18474,N_17863,N_18302);
and U18475 (N_18475,N_17763,N_18084);
and U18476 (N_18476,N_18069,N_18298);
or U18477 (N_18477,N_18200,N_18054);
nor U18478 (N_18478,N_17881,N_17655);
and U18479 (N_18479,N_18266,N_17959);
and U18480 (N_18480,N_18354,N_17936);
and U18481 (N_18481,N_17629,N_17635);
or U18482 (N_18482,N_18342,N_18010);
nor U18483 (N_18483,N_18249,N_18206);
or U18484 (N_18484,N_18202,N_18106);
nand U18485 (N_18485,N_18326,N_18315);
and U18486 (N_18486,N_17841,N_18345);
or U18487 (N_18487,N_17962,N_18117);
nand U18488 (N_18488,N_17902,N_18329);
and U18489 (N_18489,N_18256,N_18348);
nor U18490 (N_18490,N_18180,N_17732);
or U18491 (N_18491,N_18038,N_17966);
nand U18492 (N_18492,N_18093,N_17944);
nor U18493 (N_18493,N_18322,N_17691);
nand U18494 (N_18494,N_17993,N_17911);
or U18495 (N_18495,N_18110,N_17669);
nand U18496 (N_18496,N_18132,N_18336);
nand U18497 (N_18497,N_18260,N_17886);
or U18498 (N_18498,N_18254,N_17682);
nor U18499 (N_18499,N_17641,N_17683);
or U18500 (N_18500,N_17929,N_18109);
nand U18501 (N_18501,N_17839,N_17788);
or U18502 (N_18502,N_17803,N_17770);
nand U18503 (N_18503,N_17651,N_17906);
nor U18504 (N_18504,N_17960,N_18082);
and U18505 (N_18505,N_17969,N_17858);
nor U18506 (N_18506,N_18352,N_18362);
and U18507 (N_18507,N_18098,N_18365);
or U18508 (N_18508,N_17996,N_17662);
nor U18509 (N_18509,N_18368,N_17991);
nor U18510 (N_18510,N_17664,N_18203);
nand U18511 (N_18511,N_18179,N_18294);
and U18512 (N_18512,N_18140,N_17801);
or U18513 (N_18513,N_18220,N_17988);
nor U18514 (N_18514,N_17725,N_18095);
nor U18515 (N_18515,N_18191,N_17751);
and U18516 (N_18516,N_18049,N_17946);
nor U18517 (N_18517,N_18119,N_17722);
nand U18518 (N_18518,N_18000,N_17782);
or U18519 (N_18519,N_17987,N_17970);
and U18520 (N_18520,N_18307,N_17608);
and U18521 (N_18521,N_18246,N_18150);
or U18522 (N_18522,N_18035,N_18242);
nand U18523 (N_18523,N_17617,N_18014);
or U18524 (N_18524,N_18225,N_17792);
nand U18525 (N_18525,N_17642,N_17610);
nand U18526 (N_18526,N_17898,N_17879);
and U18527 (N_18527,N_17734,N_17632);
nand U18528 (N_18528,N_18341,N_18208);
nor U18529 (N_18529,N_18338,N_17885);
nand U18530 (N_18530,N_18332,N_18218);
and U18531 (N_18531,N_17878,N_18320);
or U18532 (N_18532,N_17785,N_17882);
nor U18533 (N_18533,N_17807,N_18331);
or U18534 (N_18534,N_17935,N_17685);
or U18535 (N_18535,N_17674,N_18376);
nor U18536 (N_18536,N_18137,N_18278);
nand U18537 (N_18537,N_17832,N_18009);
nor U18538 (N_18538,N_18300,N_18351);
and U18539 (N_18539,N_17951,N_18318);
nor U18540 (N_18540,N_17726,N_18359);
and U18541 (N_18541,N_17978,N_17802);
nor U18542 (N_18542,N_18089,N_18064);
or U18543 (N_18543,N_18096,N_18090);
nor U18544 (N_18544,N_18008,N_18176);
nor U18545 (N_18545,N_18099,N_18258);
or U18546 (N_18546,N_18074,N_17643);
or U18547 (N_18547,N_17851,N_18255);
or U18548 (N_18548,N_18028,N_17799);
nand U18549 (N_18549,N_18155,N_17838);
and U18550 (N_18550,N_17915,N_18066);
and U18551 (N_18551,N_18102,N_18304);
nand U18552 (N_18552,N_17934,N_18321);
nor U18553 (N_18553,N_18032,N_18280);
or U18554 (N_18554,N_17736,N_17621);
nand U18555 (N_18555,N_18396,N_18152);
and U18556 (N_18556,N_17783,N_18068);
nand U18557 (N_18557,N_17649,N_17638);
nor U18558 (N_18558,N_18100,N_17772);
and U18559 (N_18559,N_17730,N_18210);
and U18560 (N_18560,N_17733,N_18349);
nand U18561 (N_18561,N_17945,N_17766);
nand U18562 (N_18562,N_17900,N_18039);
nor U18563 (N_18563,N_17680,N_17894);
or U18564 (N_18564,N_17787,N_17869);
or U18565 (N_18565,N_17931,N_17990);
nor U18566 (N_18566,N_17686,N_18314);
nor U18567 (N_18567,N_17699,N_17756);
and U18568 (N_18568,N_18395,N_17798);
and U18569 (N_18569,N_17932,N_18353);
and U18570 (N_18570,N_17661,N_18339);
nor U18571 (N_18571,N_18381,N_17637);
nand U18572 (N_18572,N_17880,N_17645);
or U18573 (N_18573,N_17613,N_18147);
nand U18574 (N_18574,N_18094,N_18083);
or U18575 (N_18575,N_18107,N_18158);
and U18576 (N_18576,N_17846,N_18316);
or U18577 (N_18577,N_17941,N_18394);
and U18578 (N_18578,N_18299,N_17855);
nor U18579 (N_18579,N_18034,N_18305);
or U18580 (N_18580,N_17912,N_18283);
nand U18581 (N_18581,N_17835,N_18245);
nor U18582 (N_18582,N_17850,N_17626);
or U18583 (N_18583,N_18131,N_17716);
and U18584 (N_18584,N_18156,N_18020);
and U18585 (N_18585,N_18006,N_18071);
or U18586 (N_18586,N_17895,N_17687);
and U18587 (N_18587,N_17695,N_18186);
and U18588 (N_18588,N_18002,N_18178);
or U18589 (N_18589,N_17981,N_18373);
nor U18590 (N_18590,N_18129,N_18018);
and U18591 (N_18591,N_18328,N_18024);
or U18592 (N_18592,N_17602,N_17797);
or U18593 (N_18593,N_18289,N_18162);
nor U18594 (N_18594,N_17950,N_18228);
and U18595 (N_18595,N_17940,N_17701);
and U18596 (N_18596,N_17777,N_18235);
nand U18597 (N_18597,N_17888,N_17917);
nor U18598 (N_18598,N_18236,N_18044);
nand U18599 (N_18599,N_18295,N_18311);
nor U18600 (N_18600,N_17742,N_17921);
nand U18601 (N_18601,N_17707,N_18075);
or U18602 (N_18602,N_18013,N_17681);
nand U18603 (N_18603,N_18061,N_18086);
nand U18604 (N_18604,N_17868,N_18374);
nand U18605 (N_18605,N_17648,N_18325);
or U18606 (N_18606,N_18301,N_18309);
nand U18607 (N_18607,N_17823,N_17975);
or U18608 (N_18608,N_17739,N_17755);
nand U18609 (N_18609,N_17909,N_18015);
or U18610 (N_18610,N_17728,N_17752);
nand U18611 (N_18611,N_18080,N_17867);
or U18612 (N_18612,N_17658,N_18134);
or U18613 (N_18613,N_18031,N_18393);
nor U18614 (N_18614,N_18275,N_17899);
or U18615 (N_18615,N_17942,N_17829);
nor U18616 (N_18616,N_18123,N_18324);
or U18617 (N_18617,N_17816,N_18270);
nor U18618 (N_18618,N_18250,N_18174);
or U18619 (N_18619,N_18386,N_18363);
or U18620 (N_18620,N_17903,N_17746);
or U18621 (N_18621,N_18241,N_18108);
nor U18622 (N_18622,N_18171,N_17708);
or U18623 (N_18623,N_18052,N_17741);
nand U18624 (N_18624,N_18230,N_18023);
or U18625 (N_18625,N_18392,N_17790);
or U18626 (N_18626,N_17644,N_18358);
nor U18627 (N_18627,N_18172,N_18292);
nor U18628 (N_18628,N_17620,N_17709);
nand U18629 (N_18629,N_18036,N_17619);
xor U18630 (N_18630,N_17818,N_18136);
and U18631 (N_18631,N_18390,N_18269);
or U18632 (N_18632,N_18072,N_18177);
or U18633 (N_18633,N_17844,N_17631);
and U18634 (N_18634,N_17836,N_17982);
nor U18635 (N_18635,N_17666,N_17854);
or U18636 (N_18636,N_17696,N_18306);
and U18637 (N_18637,N_17675,N_18046);
and U18638 (N_18638,N_17817,N_18204);
nand U18639 (N_18639,N_18265,N_18383);
and U18640 (N_18640,N_17859,N_17952);
or U18641 (N_18641,N_17953,N_18146);
nand U18642 (N_18642,N_17625,N_17656);
nand U18643 (N_18643,N_18397,N_18058);
nand U18644 (N_18644,N_17830,N_17694);
and U18645 (N_18645,N_17748,N_17872);
nand U18646 (N_18646,N_17786,N_18276);
or U18647 (N_18647,N_18380,N_17719);
or U18648 (N_18648,N_18284,N_17667);
nand U18649 (N_18649,N_18221,N_18201);
nand U18650 (N_18650,N_17889,N_18227);
or U18651 (N_18651,N_17857,N_17697);
or U18652 (N_18652,N_18057,N_17938);
xnor U18653 (N_18653,N_18149,N_17814);
or U18654 (N_18654,N_17826,N_17764);
nand U18655 (N_18655,N_17671,N_17957);
nor U18656 (N_18656,N_17765,N_17636);
or U18657 (N_18657,N_18065,N_17612);
and U18658 (N_18658,N_17896,N_18251);
nand U18659 (N_18659,N_18022,N_18385);
and U18660 (N_18660,N_17955,N_17923);
nand U18661 (N_18661,N_18085,N_17628);
or U18662 (N_18662,N_17884,N_18233);
nand U18663 (N_18663,N_17743,N_17775);
or U18664 (N_18664,N_18040,N_18120);
nor U18665 (N_18665,N_17713,N_18238);
or U18666 (N_18666,N_17828,N_17738);
nand U18667 (N_18667,N_18169,N_18125);
nor U18668 (N_18668,N_17673,N_17837);
or U18669 (N_18669,N_18286,N_17652);
nand U18670 (N_18670,N_18111,N_17781);
and U18671 (N_18671,N_17961,N_17760);
or U18672 (N_18672,N_17714,N_18114);
and U18673 (N_18673,N_18092,N_17754);
and U18674 (N_18674,N_18113,N_17630);
nor U18675 (N_18675,N_17762,N_18398);
nor U18676 (N_18676,N_17744,N_18340);
nor U18677 (N_18677,N_18122,N_18237);
nand U18678 (N_18678,N_17862,N_18012);
nand U18679 (N_18679,N_17665,N_18190);
nor U18680 (N_18680,N_17759,N_18377);
nor U18681 (N_18681,N_18127,N_17821);
nor U18682 (N_18682,N_18115,N_17615);
and U18683 (N_18683,N_17824,N_18003);
and U18684 (N_18684,N_17603,N_18357);
nand U18685 (N_18685,N_17812,N_18011);
or U18686 (N_18686,N_17745,N_17605);
nor U18687 (N_18687,N_18369,N_18164);
and U18688 (N_18688,N_18372,N_18141);
or U18689 (N_18689,N_17908,N_17624);
nand U18690 (N_18690,N_17930,N_17842);
nor U18691 (N_18691,N_17794,N_18343);
or U18692 (N_18692,N_18081,N_17972);
nand U18693 (N_18693,N_17618,N_18244);
and U18694 (N_18694,N_18001,N_18253);
nand U18695 (N_18695,N_17811,N_17753);
and U18696 (N_18696,N_17834,N_17729);
or U18697 (N_18697,N_18124,N_17668);
nand U18698 (N_18698,N_18399,N_18196);
nand U18699 (N_18699,N_17737,N_18105);
and U18700 (N_18700,N_18272,N_17847);
or U18701 (N_18701,N_18303,N_18088);
and U18702 (N_18702,N_17779,N_18198);
nand U18703 (N_18703,N_17870,N_18333);
nor U18704 (N_18704,N_18026,N_18223);
and U18705 (N_18705,N_17892,N_17800);
or U18706 (N_18706,N_17804,N_17705);
or U18707 (N_18707,N_18214,N_18317);
nor U18708 (N_18708,N_18366,N_18037);
nand U18709 (N_18709,N_18335,N_18211);
or U18710 (N_18710,N_18185,N_18027);
nor U18711 (N_18711,N_18222,N_17650);
or U18712 (N_18712,N_18281,N_18050);
or U18713 (N_18713,N_18391,N_17758);
nand U18714 (N_18714,N_18168,N_18184);
nand U18715 (N_18715,N_18205,N_18101);
and U18716 (N_18716,N_18267,N_17877);
or U18717 (N_18717,N_18135,N_18367);
nor U18718 (N_18718,N_18388,N_18079);
nand U18719 (N_18719,N_17973,N_17860);
or U18720 (N_18720,N_17653,N_17864);
and U18721 (N_18721,N_18063,N_18207);
and U18722 (N_18722,N_18151,N_18153);
or U18723 (N_18723,N_18232,N_18070);
or U18724 (N_18724,N_17825,N_17609);
nand U18725 (N_18725,N_17810,N_17891);
nand U18726 (N_18726,N_17678,N_18360);
nand U18727 (N_18727,N_18170,N_18290);
nor U18728 (N_18728,N_17997,N_18154);
and U18729 (N_18729,N_18361,N_18384);
and U18730 (N_18730,N_18209,N_17780);
nand U18731 (N_18731,N_18195,N_18263);
nand U18732 (N_18732,N_18142,N_18078);
or U18733 (N_18733,N_18163,N_17907);
nor U18734 (N_18734,N_17659,N_17774);
or U18735 (N_18735,N_17717,N_17965);
and U18736 (N_18736,N_18045,N_17805);
or U18737 (N_18737,N_17994,N_17852);
nand U18738 (N_18738,N_18133,N_17702);
nor U18739 (N_18739,N_18043,N_17843);
xor U18740 (N_18740,N_17604,N_18243);
nor U18741 (N_18741,N_18182,N_18247);
or U18742 (N_18742,N_18296,N_18112);
nor U18743 (N_18743,N_18274,N_17723);
and U18744 (N_18744,N_17813,N_18261);
or U18745 (N_18745,N_18257,N_17769);
nand U18746 (N_18746,N_18234,N_17670);
and U18747 (N_18747,N_17893,N_17622);
or U18748 (N_18748,N_18355,N_17897);
or U18749 (N_18749,N_17848,N_18224);
nor U18750 (N_18750,N_17985,N_18116);
nor U18751 (N_18751,N_17749,N_18121);
and U18752 (N_18752,N_17853,N_17943);
nor U18753 (N_18753,N_17784,N_18188);
and U18754 (N_18754,N_17720,N_18148);
nor U18755 (N_18755,N_18007,N_18291);
nand U18756 (N_18756,N_18161,N_18264);
nand U18757 (N_18757,N_18226,N_18259);
and U18758 (N_18758,N_17735,N_17905);
and U18759 (N_18759,N_18389,N_18215);
and U18760 (N_18760,N_18056,N_18216);
and U18761 (N_18761,N_17939,N_18067);
nor U18762 (N_18762,N_18097,N_18248);
and U18763 (N_18763,N_17731,N_17684);
nor U18764 (N_18764,N_17611,N_17849);
or U18765 (N_18765,N_17933,N_17796);
xor U18766 (N_18766,N_18199,N_18087);
nand U18767 (N_18767,N_18310,N_17876);
nand U18768 (N_18768,N_17698,N_17740);
and U18769 (N_18769,N_17676,N_17747);
nand U18770 (N_18770,N_18130,N_17711);
or U18771 (N_18771,N_18017,N_17914);
nor U18772 (N_18772,N_17768,N_18145);
or U18773 (N_18773,N_18364,N_17778);
nor U18774 (N_18774,N_17918,N_17704);
or U18775 (N_18775,N_18213,N_18346);
and U18776 (N_18776,N_18197,N_18157);
nor U18777 (N_18777,N_18021,N_18347);
nand U18778 (N_18778,N_17999,N_17607);
and U18779 (N_18779,N_18091,N_17672);
nand U18780 (N_18780,N_18371,N_17724);
nor U18781 (N_18781,N_17890,N_18308);
or U18782 (N_18782,N_18344,N_17856);
nor U18783 (N_18783,N_17833,N_18337);
or U18784 (N_18784,N_17677,N_17601);
nor U18785 (N_18785,N_17646,N_18240);
nand U18786 (N_18786,N_17614,N_17871);
nor U18787 (N_18787,N_18126,N_17789);
nand U18788 (N_18788,N_18062,N_17692);
nor U18789 (N_18789,N_17984,N_18231);
nor U18790 (N_18790,N_17861,N_18139);
or U18791 (N_18791,N_17971,N_17606);
nor U18792 (N_18792,N_18279,N_18382);
or U18793 (N_18793,N_18029,N_17616);
nor U18794 (N_18794,N_18194,N_17958);
nor U18795 (N_18795,N_18277,N_17633);
nor U18796 (N_18796,N_18128,N_18144);
nand U18797 (N_18797,N_17795,N_17727);
or U18798 (N_18798,N_17937,N_17750);
and U18799 (N_18799,N_18350,N_18076);
and U18800 (N_18800,N_18091,N_18350);
nand U18801 (N_18801,N_18304,N_17866);
or U18802 (N_18802,N_18107,N_18163);
and U18803 (N_18803,N_17699,N_17843);
and U18804 (N_18804,N_18143,N_17774);
nor U18805 (N_18805,N_17933,N_17884);
nand U18806 (N_18806,N_18385,N_17919);
or U18807 (N_18807,N_17955,N_17753);
nor U18808 (N_18808,N_17760,N_18219);
or U18809 (N_18809,N_18050,N_18378);
nand U18810 (N_18810,N_18247,N_18096);
nor U18811 (N_18811,N_18170,N_17969);
nor U18812 (N_18812,N_18359,N_18198);
nand U18813 (N_18813,N_18373,N_18203);
and U18814 (N_18814,N_17996,N_17672);
or U18815 (N_18815,N_17761,N_17661);
and U18816 (N_18816,N_18078,N_17858);
nand U18817 (N_18817,N_17769,N_17736);
and U18818 (N_18818,N_17771,N_18292);
nand U18819 (N_18819,N_18131,N_17974);
and U18820 (N_18820,N_18051,N_18002);
or U18821 (N_18821,N_18160,N_18127);
nor U18822 (N_18822,N_17639,N_18355);
and U18823 (N_18823,N_18252,N_18169);
or U18824 (N_18824,N_17622,N_17713);
nand U18825 (N_18825,N_18367,N_17995);
nand U18826 (N_18826,N_17645,N_18139);
or U18827 (N_18827,N_17845,N_18215);
xor U18828 (N_18828,N_18300,N_17796);
and U18829 (N_18829,N_17659,N_18149);
and U18830 (N_18830,N_18058,N_17908);
nor U18831 (N_18831,N_17641,N_18089);
nand U18832 (N_18832,N_18210,N_18150);
or U18833 (N_18833,N_17991,N_17954);
nor U18834 (N_18834,N_17887,N_18040);
or U18835 (N_18835,N_18257,N_18240);
nor U18836 (N_18836,N_17864,N_18213);
nor U18837 (N_18837,N_17993,N_18381);
nand U18838 (N_18838,N_17976,N_18267);
nor U18839 (N_18839,N_17870,N_18129);
and U18840 (N_18840,N_17976,N_17665);
nor U18841 (N_18841,N_17687,N_18297);
or U18842 (N_18842,N_17675,N_18293);
and U18843 (N_18843,N_17642,N_18070);
nand U18844 (N_18844,N_18168,N_18378);
or U18845 (N_18845,N_17630,N_18008);
and U18846 (N_18846,N_17750,N_17798);
and U18847 (N_18847,N_18170,N_17623);
or U18848 (N_18848,N_18114,N_17905);
nor U18849 (N_18849,N_18101,N_17729);
or U18850 (N_18850,N_17903,N_18000);
xor U18851 (N_18851,N_17915,N_17779);
nand U18852 (N_18852,N_17827,N_18044);
nor U18853 (N_18853,N_17684,N_17997);
or U18854 (N_18854,N_17803,N_18199);
or U18855 (N_18855,N_18001,N_18268);
nor U18856 (N_18856,N_17934,N_18218);
nand U18857 (N_18857,N_18016,N_18142);
nor U18858 (N_18858,N_18367,N_17702);
nor U18859 (N_18859,N_17796,N_17995);
nand U18860 (N_18860,N_17634,N_18338);
or U18861 (N_18861,N_18053,N_17818);
and U18862 (N_18862,N_18005,N_18315);
and U18863 (N_18863,N_17744,N_17784);
nor U18864 (N_18864,N_18338,N_17636);
nand U18865 (N_18865,N_17700,N_17770);
and U18866 (N_18866,N_18370,N_18240);
nor U18867 (N_18867,N_18381,N_17839);
or U18868 (N_18868,N_18353,N_18289);
or U18869 (N_18869,N_18190,N_18291);
or U18870 (N_18870,N_18335,N_17606);
nor U18871 (N_18871,N_17803,N_18282);
and U18872 (N_18872,N_17610,N_17689);
or U18873 (N_18873,N_17751,N_18347);
or U18874 (N_18874,N_17717,N_18086);
xnor U18875 (N_18875,N_17839,N_18230);
nand U18876 (N_18876,N_18306,N_17735);
and U18877 (N_18877,N_17840,N_18010);
nor U18878 (N_18878,N_17910,N_18210);
or U18879 (N_18879,N_18176,N_18387);
nand U18880 (N_18880,N_17624,N_18122);
nand U18881 (N_18881,N_18356,N_17943);
nor U18882 (N_18882,N_18095,N_18187);
nor U18883 (N_18883,N_18281,N_17851);
or U18884 (N_18884,N_17716,N_17773);
nand U18885 (N_18885,N_18262,N_18108);
and U18886 (N_18886,N_17994,N_18175);
nor U18887 (N_18887,N_18392,N_17871);
and U18888 (N_18888,N_17916,N_18330);
nand U18889 (N_18889,N_17671,N_18055);
xnor U18890 (N_18890,N_17929,N_18061);
or U18891 (N_18891,N_18160,N_18308);
nand U18892 (N_18892,N_18352,N_18005);
nand U18893 (N_18893,N_18167,N_17967);
nand U18894 (N_18894,N_18150,N_17637);
or U18895 (N_18895,N_17800,N_17770);
or U18896 (N_18896,N_18288,N_17739);
or U18897 (N_18897,N_17696,N_17930);
or U18898 (N_18898,N_17613,N_17780);
and U18899 (N_18899,N_17808,N_18196);
or U18900 (N_18900,N_18270,N_18220);
nor U18901 (N_18901,N_17990,N_18322);
and U18902 (N_18902,N_18212,N_17739);
nand U18903 (N_18903,N_18373,N_18248);
or U18904 (N_18904,N_17761,N_18122);
or U18905 (N_18905,N_17636,N_17785);
nor U18906 (N_18906,N_17684,N_17712);
or U18907 (N_18907,N_18070,N_18034);
nor U18908 (N_18908,N_18304,N_18014);
and U18909 (N_18909,N_18190,N_17855);
nor U18910 (N_18910,N_17709,N_17949);
nor U18911 (N_18911,N_17961,N_17790);
nand U18912 (N_18912,N_17687,N_17905);
nor U18913 (N_18913,N_17656,N_18289);
and U18914 (N_18914,N_18169,N_18217);
nor U18915 (N_18915,N_18056,N_18325);
nand U18916 (N_18916,N_17757,N_17659);
and U18917 (N_18917,N_17670,N_18341);
or U18918 (N_18918,N_18001,N_17940);
nand U18919 (N_18919,N_17662,N_17641);
or U18920 (N_18920,N_17979,N_18178);
or U18921 (N_18921,N_18138,N_17630);
or U18922 (N_18922,N_17738,N_17915);
and U18923 (N_18923,N_17976,N_18363);
nand U18924 (N_18924,N_17862,N_17736);
or U18925 (N_18925,N_17630,N_17891);
nand U18926 (N_18926,N_18141,N_18214);
and U18927 (N_18927,N_18128,N_18110);
or U18928 (N_18928,N_18004,N_18375);
and U18929 (N_18929,N_18274,N_18013);
nand U18930 (N_18930,N_18211,N_18285);
and U18931 (N_18931,N_17721,N_18184);
and U18932 (N_18932,N_18185,N_18280);
nand U18933 (N_18933,N_17886,N_17724);
or U18934 (N_18934,N_18221,N_18133);
nor U18935 (N_18935,N_18086,N_17944);
or U18936 (N_18936,N_18213,N_18254);
xor U18937 (N_18937,N_17734,N_18353);
nand U18938 (N_18938,N_17838,N_17726);
nor U18939 (N_18939,N_18037,N_18047);
xnor U18940 (N_18940,N_17964,N_17945);
nand U18941 (N_18941,N_18099,N_18220);
nor U18942 (N_18942,N_18072,N_17756);
nor U18943 (N_18943,N_18046,N_18175);
nand U18944 (N_18944,N_17731,N_17772);
nand U18945 (N_18945,N_18259,N_18156);
or U18946 (N_18946,N_18342,N_17914);
or U18947 (N_18947,N_18312,N_17699);
or U18948 (N_18948,N_18198,N_17786);
and U18949 (N_18949,N_18348,N_18091);
nor U18950 (N_18950,N_18283,N_18279);
nand U18951 (N_18951,N_18268,N_18205);
nand U18952 (N_18952,N_18303,N_17609);
or U18953 (N_18953,N_18075,N_18340);
or U18954 (N_18954,N_17992,N_17939);
nor U18955 (N_18955,N_18251,N_17994);
or U18956 (N_18956,N_18246,N_18229);
or U18957 (N_18957,N_17822,N_18056);
or U18958 (N_18958,N_17812,N_17601);
or U18959 (N_18959,N_17935,N_18028);
or U18960 (N_18960,N_17775,N_18145);
nand U18961 (N_18961,N_17883,N_17876);
and U18962 (N_18962,N_18158,N_17951);
and U18963 (N_18963,N_18351,N_17744);
xor U18964 (N_18964,N_17859,N_17772);
nor U18965 (N_18965,N_18039,N_18235);
nor U18966 (N_18966,N_18335,N_17700);
and U18967 (N_18967,N_17802,N_18010);
nor U18968 (N_18968,N_18227,N_18396);
nand U18969 (N_18969,N_18239,N_18014);
nand U18970 (N_18970,N_18068,N_17888);
nand U18971 (N_18971,N_17656,N_18303);
or U18972 (N_18972,N_17715,N_17895);
nor U18973 (N_18973,N_17813,N_18026);
nand U18974 (N_18974,N_18346,N_17826);
or U18975 (N_18975,N_17952,N_18101);
and U18976 (N_18976,N_17629,N_18093);
nor U18977 (N_18977,N_17910,N_18203);
and U18978 (N_18978,N_17677,N_17733);
and U18979 (N_18979,N_18337,N_17869);
nand U18980 (N_18980,N_17969,N_18066);
nor U18981 (N_18981,N_17825,N_17928);
nor U18982 (N_18982,N_17692,N_18340);
nor U18983 (N_18983,N_17755,N_18232);
nand U18984 (N_18984,N_18290,N_18153);
nand U18985 (N_18985,N_17826,N_18188);
and U18986 (N_18986,N_17947,N_17904);
nor U18987 (N_18987,N_17988,N_17634);
nor U18988 (N_18988,N_18221,N_17806);
or U18989 (N_18989,N_17904,N_17878);
nor U18990 (N_18990,N_18192,N_18087);
nand U18991 (N_18991,N_17627,N_17642);
nor U18992 (N_18992,N_17809,N_17791);
nand U18993 (N_18993,N_18293,N_17815);
nor U18994 (N_18994,N_18193,N_18195);
nand U18995 (N_18995,N_17805,N_18006);
nand U18996 (N_18996,N_17967,N_18373);
xor U18997 (N_18997,N_18050,N_17719);
nor U18998 (N_18998,N_17668,N_18189);
or U18999 (N_18999,N_18052,N_17812);
and U19000 (N_19000,N_17641,N_18005);
and U19001 (N_19001,N_18228,N_17709);
nand U19002 (N_19002,N_17848,N_18299);
or U19003 (N_19003,N_18114,N_17788);
nor U19004 (N_19004,N_17793,N_18377);
nand U19005 (N_19005,N_17676,N_17631);
nor U19006 (N_19006,N_18381,N_18181);
and U19007 (N_19007,N_18286,N_18348);
and U19008 (N_19008,N_18029,N_17807);
or U19009 (N_19009,N_18368,N_18245);
or U19010 (N_19010,N_18084,N_17800);
and U19011 (N_19011,N_18350,N_17690);
or U19012 (N_19012,N_18174,N_17849);
or U19013 (N_19013,N_17927,N_17729);
or U19014 (N_19014,N_18216,N_17922);
nand U19015 (N_19015,N_17796,N_18043);
and U19016 (N_19016,N_18189,N_18254);
nor U19017 (N_19017,N_18079,N_17951);
nand U19018 (N_19018,N_18229,N_18160);
xnor U19019 (N_19019,N_17808,N_18238);
nor U19020 (N_19020,N_18270,N_18330);
nand U19021 (N_19021,N_18289,N_17755);
nor U19022 (N_19022,N_17677,N_17785);
or U19023 (N_19023,N_17930,N_17899);
and U19024 (N_19024,N_17658,N_17662);
and U19025 (N_19025,N_17893,N_17806);
and U19026 (N_19026,N_17749,N_18185);
nand U19027 (N_19027,N_17627,N_17779);
nor U19028 (N_19028,N_18270,N_18077);
nand U19029 (N_19029,N_17739,N_18331);
nor U19030 (N_19030,N_18070,N_18175);
nor U19031 (N_19031,N_17886,N_18326);
nand U19032 (N_19032,N_18171,N_18154);
nand U19033 (N_19033,N_17674,N_17788);
nor U19034 (N_19034,N_18369,N_18051);
and U19035 (N_19035,N_18276,N_17707);
or U19036 (N_19036,N_17788,N_17603);
and U19037 (N_19037,N_18124,N_18290);
nand U19038 (N_19038,N_18272,N_17909);
nand U19039 (N_19039,N_17976,N_18228);
or U19040 (N_19040,N_17744,N_18032);
and U19041 (N_19041,N_17784,N_17999);
nand U19042 (N_19042,N_17981,N_18341);
nor U19043 (N_19043,N_17918,N_18354);
nand U19044 (N_19044,N_18260,N_18114);
and U19045 (N_19045,N_18371,N_18057);
nand U19046 (N_19046,N_17963,N_17814);
and U19047 (N_19047,N_18051,N_17729);
nor U19048 (N_19048,N_17770,N_17779);
or U19049 (N_19049,N_18170,N_17922);
or U19050 (N_19050,N_18060,N_18148);
and U19051 (N_19051,N_17701,N_18078);
or U19052 (N_19052,N_17668,N_17832);
nand U19053 (N_19053,N_18370,N_17858);
and U19054 (N_19054,N_17883,N_17673);
and U19055 (N_19055,N_18191,N_17938);
nand U19056 (N_19056,N_17802,N_18069);
nand U19057 (N_19057,N_18172,N_17934);
or U19058 (N_19058,N_17711,N_17772);
or U19059 (N_19059,N_17727,N_18206);
and U19060 (N_19060,N_17807,N_18186);
or U19061 (N_19061,N_17696,N_18232);
nand U19062 (N_19062,N_18367,N_17906);
or U19063 (N_19063,N_18297,N_17914);
nor U19064 (N_19064,N_17924,N_17991);
or U19065 (N_19065,N_18360,N_17885);
nor U19066 (N_19066,N_17877,N_18315);
and U19067 (N_19067,N_18164,N_18225);
nand U19068 (N_19068,N_17783,N_17650);
nand U19069 (N_19069,N_17928,N_18253);
nand U19070 (N_19070,N_18338,N_17783);
or U19071 (N_19071,N_17829,N_17803);
and U19072 (N_19072,N_17742,N_17799);
and U19073 (N_19073,N_18255,N_18300);
or U19074 (N_19074,N_17886,N_17808);
or U19075 (N_19075,N_18216,N_17761);
xnor U19076 (N_19076,N_18039,N_18194);
nor U19077 (N_19077,N_17668,N_17634);
nand U19078 (N_19078,N_17803,N_17995);
nand U19079 (N_19079,N_17936,N_17618);
and U19080 (N_19080,N_17976,N_18270);
nand U19081 (N_19081,N_18042,N_17678);
and U19082 (N_19082,N_18338,N_18361);
nand U19083 (N_19083,N_17761,N_17977);
or U19084 (N_19084,N_18024,N_17809);
nor U19085 (N_19085,N_18266,N_18292);
nand U19086 (N_19086,N_18360,N_17897);
nor U19087 (N_19087,N_17704,N_18039);
and U19088 (N_19088,N_18372,N_18133);
nor U19089 (N_19089,N_18371,N_17838);
and U19090 (N_19090,N_18194,N_17782);
nor U19091 (N_19091,N_18253,N_18068);
nand U19092 (N_19092,N_18060,N_17811);
or U19093 (N_19093,N_18395,N_18362);
and U19094 (N_19094,N_18106,N_17871);
or U19095 (N_19095,N_18178,N_17742);
or U19096 (N_19096,N_18292,N_17911);
nor U19097 (N_19097,N_17920,N_17653);
or U19098 (N_19098,N_17667,N_18281);
or U19099 (N_19099,N_18092,N_17657);
nor U19100 (N_19100,N_18333,N_17764);
nand U19101 (N_19101,N_18201,N_17680);
xnor U19102 (N_19102,N_17781,N_17934);
nand U19103 (N_19103,N_18153,N_18014);
nand U19104 (N_19104,N_17634,N_17990);
nand U19105 (N_19105,N_17604,N_17744);
or U19106 (N_19106,N_17763,N_18302);
nand U19107 (N_19107,N_18329,N_18225);
or U19108 (N_19108,N_17618,N_17666);
or U19109 (N_19109,N_17747,N_18312);
nand U19110 (N_19110,N_17669,N_17886);
and U19111 (N_19111,N_17997,N_18298);
or U19112 (N_19112,N_18354,N_18379);
or U19113 (N_19113,N_18329,N_17975);
and U19114 (N_19114,N_17699,N_17814);
nor U19115 (N_19115,N_17873,N_17691);
nand U19116 (N_19116,N_18066,N_18225);
nor U19117 (N_19117,N_18187,N_18247);
nand U19118 (N_19118,N_17698,N_18184);
and U19119 (N_19119,N_18073,N_18336);
nor U19120 (N_19120,N_18131,N_18133);
and U19121 (N_19121,N_17826,N_18193);
nor U19122 (N_19122,N_17992,N_17910);
nor U19123 (N_19123,N_18040,N_17819);
nor U19124 (N_19124,N_18141,N_17928);
nor U19125 (N_19125,N_18127,N_18181);
and U19126 (N_19126,N_17646,N_17772);
nand U19127 (N_19127,N_18030,N_17776);
and U19128 (N_19128,N_17774,N_17847);
or U19129 (N_19129,N_18357,N_17683);
and U19130 (N_19130,N_18125,N_18150);
nand U19131 (N_19131,N_17843,N_18354);
nor U19132 (N_19132,N_18277,N_18363);
nand U19133 (N_19133,N_17652,N_18201);
nand U19134 (N_19134,N_17915,N_18132);
nor U19135 (N_19135,N_17993,N_17831);
and U19136 (N_19136,N_18362,N_18317);
nand U19137 (N_19137,N_18122,N_17746);
nor U19138 (N_19138,N_18021,N_18239);
nor U19139 (N_19139,N_18019,N_18205);
or U19140 (N_19140,N_18215,N_17636);
nor U19141 (N_19141,N_17763,N_17729);
nor U19142 (N_19142,N_17655,N_17950);
nand U19143 (N_19143,N_17731,N_17600);
and U19144 (N_19144,N_17899,N_18265);
or U19145 (N_19145,N_17954,N_17909);
nand U19146 (N_19146,N_17924,N_18167);
nor U19147 (N_19147,N_18059,N_17830);
or U19148 (N_19148,N_18327,N_18283);
or U19149 (N_19149,N_18092,N_17632);
nand U19150 (N_19150,N_18090,N_17637);
or U19151 (N_19151,N_17718,N_18188);
and U19152 (N_19152,N_18315,N_18216);
nand U19153 (N_19153,N_18388,N_18051);
nand U19154 (N_19154,N_17792,N_17832);
and U19155 (N_19155,N_17797,N_18377);
nor U19156 (N_19156,N_18141,N_18150);
and U19157 (N_19157,N_17855,N_18255);
nor U19158 (N_19158,N_18220,N_17974);
nor U19159 (N_19159,N_18005,N_18102);
and U19160 (N_19160,N_18366,N_18261);
nand U19161 (N_19161,N_18109,N_18006);
nor U19162 (N_19162,N_18087,N_18023);
nor U19163 (N_19163,N_18269,N_17986);
and U19164 (N_19164,N_17643,N_17927);
or U19165 (N_19165,N_18052,N_18157);
nor U19166 (N_19166,N_18285,N_18172);
or U19167 (N_19167,N_18113,N_17942);
or U19168 (N_19168,N_18211,N_18274);
or U19169 (N_19169,N_18257,N_18085);
nor U19170 (N_19170,N_18127,N_17709);
nor U19171 (N_19171,N_17790,N_18267);
and U19172 (N_19172,N_17712,N_17645);
nor U19173 (N_19173,N_18120,N_18304);
or U19174 (N_19174,N_18227,N_17707);
nand U19175 (N_19175,N_18228,N_18320);
nor U19176 (N_19176,N_18279,N_18095);
nor U19177 (N_19177,N_18036,N_18143);
nand U19178 (N_19178,N_17835,N_17744);
nand U19179 (N_19179,N_17853,N_17994);
or U19180 (N_19180,N_17631,N_18095);
nor U19181 (N_19181,N_17667,N_18085);
nor U19182 (N_19182,N_17972,N_17987);
nand U19183 (N_19183,N_18344,N_18082);
nand U19184 (N_19184,N_18202,N_18358);
or U19185 (N_19185,N_17910,N_18283);
or U19186 (N_19186,N_17616,N_17996);
nand U19187 (N_19187,N_17969,N_17601);
nand U19188 (N_19188,N_17716,N_17987);
or U19189 (N_19189,N_18363,N_18046);
nor U19190 (N_19190,N_18309,N_17983);
nand U19191 (N_19191,N_17778,N_18319);
nand U19192 (N_19192,N_17972,N_18121);
or U19193 (N_19193,N_18044,N_18053);
or U19194 (N_19194,N_17601,N_17660);
or U19195 (N_19195,N_17853,N_17795);
or U19196 (N_19196,N_17737,N_18081);
and U19197 (N_19197,N_18326,N_18394);
nor U19198 (N_19198,N_17818,N_18246);
nand U19199 (N_19199,N_17626,N_18052);
and U19200 (N_19200,N_18916,N_18689);
nand U19201 (N_19201,N_18735,N_19070);
or U19202 (N_19202,N_18640,N_18774);
nand U19203 (N_19203,N_18754,N_18747);
and U19204 (N_19204,N_19041,N_19069);
or U19205 (N_19205,N_18732,N_18554);
or U19206 (N_19206,N_18792,N_18587);
nand U19207 (N_19207,N_18626,N_18543);
nand U19208 (N_19208,N_19164,N_18548);
or U19209 (N_19209,N_19184,N_18571);
nor U19210 (N_19210,N_18863,N_19096);
or U19211 (N_19211,N_18716,N_18615);
and U19212 (N_19212,N_18831,N_19007);
xor U19213 (N_19213,N_18421,N_19124);
or U19214 (N_19214,N_18468,N_18429);
nand U19215 (N_19215,N_18785,N_18847);
and U19216 (N_19216,N_19154,N_18676);
and U19217 (N_19217,N_19165,N_18550);
and U19218 (N_19218,N_18555,N_18857);
and U19219 (N_19219,N_19040,N_18565);
nor U19220 (N_19220,N_18400,N_18599);
nand U19221 (N_19221,N_18406,N_19052);
or U19222 (N_19222,N_18845,N_18422);
nor U19223 (N_19223,N_18466,N_18434);
or U19224 (N_19224,N_19121,N_18741);
nor U19225 (N_19225,N_18883,N_18808);
and U19226 (N_19226,N_18632,N_18670);
nor U19227 (N_19227,N_18749,N_19162);
nor U19228 (N_19228,N_18909,N_19123);
nand U19229 (N_19229,N_18534,N_18974);
or U19230 (N_19230,N_18625,N_18842);
and U19231 (N_19231,N_19144,N_19075);
nand U19232 (N_19232,N_18979,N_19112);
nor U19233 (N_19233,N_19054,N_19066);
and U19234 (N_19234,N_18603,N_18743);
nand U19235 (N_19235,N_18506,N_18728);
or U19236 (N_19236,N_19183,N_19025);
and U19237 (N_19237,N_18494,N_18514);
xnor U19238 (N_19238,N_18901,N_18800);
nor U19239 (N_19239,N_18585,N_18451);
and U19240 (N_19240,N_18899,N_18556);
and U19241 (N_19241,N_18870,N_18773);
nor U19242 (N_19242,N_18865,N_18660);
nand U19243 (N_19243,N_19093,N_18493);
and U19244 (N_19244,N_18944,N_18456);
nor U19245 (N_19245,N_18699,N_18614);
and U19246 (N_19246,N_19005,N_18923);
nor U19247 (N_19247,N_18520,N_18746);
nor U19248 (N_19248,N_18873,N_19171);
nand U19249 (N_19249,N_18634,N_18818);
nor U19250 (N_19250,N_18824,N_18907);
and U19251 (N_19251,N_18673,N_19017);
nor U19252 (N_19252,N_19181,N_19085);
or U19253 (N_19253,N_19035,N_18991);
xnor U19254 (N_19254,N_19147,N_18665);
or U19255 (N_19255,N_19145,N_18450);
nor U19256 (N_19256,N_19026,N_18521);
or U19257 (N_19257,N_18533,N_18612);
nor U19258 (N_19258,N_18681,N_18410);
and U19259 (N_19259,N_19081,N_18874);
and U19260 (N_19260,N_18758,N_18940);
nand U19261 (N_19261,N_18569,N_18969);
nor U19262 (N_19262,N_19047,N_18581);
nor U19263 (N_19263,N_18639,N_18545);
and U19264 (N_19264,N_18577,N_18481);
and U19265 (N_19265,N_19033,N_18678);
and U19266 (N_19266,N_18935,N_18621);
or U19267 (N_19267,N_18835,N_18862);
or U19268 (N_19268,N_18697,N_18557);
or U19269 (N_19269,N_19125,N_18685);
nand U19270 (N_19270,N_19021,N_18775);
xor U19271 (N_19271,N_18996,N_18801);
or U19272 (N_19272,N_18837,N_18489);
nor U19273 (N_19273,N_19191,N_19051);
or U19274 (N_19274,N_18423,N_19114);
or U19275 (N_19275,N_18963,N_18522);
and U19276 (N_19276,N_18441,N_18849);
nor U19277 (N_19277,N_19119,N_18932);
xnor U19278 (N_19278,N_19100,N_19042);
and U19279 (N_19279,N_18720,N_18449);
nor U19280 (N_19280,N_19107,N_18913);
and U19281 (N_19281,N_19101,N_18627);
nor U19282 (N_19282,N_18787,N_19126);
nand U19283 (N_19283,N_18680,N_18455);
nor U19284 (N_19284,N_18498,N_18496);
nand U19285 (N_19285,N_18814,N_18630);
nor U19286 (N_19286,N_18579,N_18917);
and U19287 (N_19287,N_18443,N_18420);
nand U19288 (N_19288,N_18440,N_18897);
nand U19289 (N_19289,N_18624,N_18582);
and U19290 (N_19290,N_19089,N_19088);
and U19291 (N_19291,N_19142,N_18834);
and U19292 (N_19292,N_18851,N_18971);
or U19293 (N_19293,N_18575,N_18675);
nand U19294 (N_19294,N_18714,N_19030);
nand U19295 (N_19295,N_18731,N_18852);
or U19296 (N_19296,N_18633,N_18433);
and U19297 (N_19297,N_18461,N_18515);
and U19298 (N_19298,N_18967,N_18962);
nand U19299 (N_19299,N_19060,N_19168);
and U19300 (N_19300,N_19055,N_19079);
nand U19301 (N_19301,N_19149,N_18813);
nor U19302 (N_19302,N_18791,N_18952);
nand U19303 (N_19303,N_18649,N_19132);
and U19304 (N_19304,N_18957,N_18998);
nand U19305 (N_19305,N_19151,N_18536);
and U19306 (N_19306,N_18667,N_18715);
and U19307 (N_19307,N_18478,N_19053);
or U19308 (N_19308,N_18797,N_18964);
nor U19309 (N_19309,N_18495,N_18644);
nand U19310 (N_19310,N_18419,N_19086);
nand U19311 (N_19311,N_19062,N_18475);
and U19312 (N_19312,N_18802,N_18447);
or U19313 (N_19313,N_18896,N_18472);
nand U19314 (N_19314,N_18929,N_18799);
nor U19315 (N_19315,N_18620,N_18505);
nand U19316 (N_19316,N_18884,N_18822);
or U19317 (N_19317,N_18994,N_18497);
nand U19318 (N_19318,N_18700,N_18658);
nor U19319 (N_19319,N_18954,N_18558);
nand U19320 (N_19320,N_18807,N_18942);
nor U19321 (N_19321,N_19048,N_18958);
and U19322 (N_19322,N_18803,N_19128);
nor U19323 (N_19323,N_18580,N_18961);
and U19324 (N_19324,N_18938,N_18510);
nor U19325 (N_19325,N_18753,N_18442);
nand U19326 (N_19326,N_18826,N_18539);
nor U19327 (N_19327,N_18424,N_18618);
and U19328 (N_19328,N_18764,N_18823);
and U19329 (N_19329,N_19068,N_18972);
nor U19330 (N_19330,N_18610,N_19039);
nand U19331 (N_19331,N_18476,N_18462);
nor U19332 (N_19332,N_18647,N_19167);
nand U19333 (N_19333,N_18866,N_18927);
and U19334 (N_19334,N_19049,N_18409);
and U19335 (N_19335,N_19141,N_18708);
nand U19336 (N_19336,N_18730,N_18888);
or U19337 (N_19337,N_18759,N_19058);
nand U19338 (N_19338,N_18672,N_18605);
nand U19339 (N_19339,N_19152,N_19120);
nand U19340 (N_19340,N_18578,N_18815);
or U19341 (N_19341,N_18993,N_19158);
and U19342 (N_19342,N_19190,N_18693);
or U19343 (N_19343,N_18487,N_18805);
nand U19344 (N_19344,N_19178,N_18637);
nand U19345 (N_19345,N_19194,N_18454);
or U19346 (N_19346,N_18457,N_18717);
and U19347 (N_19347,N_18418,N_18525);
or U19348 (N_19348,N_18950,N_18491);
nand U19349 (N_19349,N_19139,N_19076);
and U19350 (N_19350,N_18524,N_18904);
or U19351 (N_19351,N_18628,N_18987);
and U19352 (N_19352,N_18878,N_19027);
or U19353 (N_19353,N_18893,N_18982);
and U19354 (N_19354,N_18513,N_18919);
and U19355 (N_19355,N_19138,N_18407);
and U19356 (N_19356,N_18793,N_18947);
nand U19357 (N_19357,N_18425,N_18934);
nand U19358 (N_19358,N_18654,N_18984);
nand U19359 (N_19359,N_18782,N_18761);
xnor U19360 (N_19360,N_18794,N_19180);
and U19361 (N_19361,N_18756,N_19187);
nor U19362 (N_19362,N_18684,N_18414);
and U19363 (N_19363,N_18609,N_18978);
and U19364 (N_19364,N_18776,N_18464);
nor U19365 (N_19365,N_18903,N_18674);
xnor U19366 (N_19366,N_18920,N_18894);
or U19367 (N_19367,N_18981,N_18540);
or U19368 (N_19368,N_18733,N_18825);
nand U19369 (N_19369,N_18829,N_18483);
and U19370 (N_19370,N_18530,N_19022);
xor U19371 (N_19371,N_18566,N_18943);
or U19372 (N_19372,N_18868,N_18860);
and U19373 (N_19373,N_18711,N_18688);
or U19374 (N_19374,N_19135,N_18918);
nand U19375 (N_19375,N_18588,N_19045);
or U19376 (N_19376,N_18959,N_18526);
nand U19377 (N_19377,N_18703,N_18473);
nor U19378 (N_19378,N_18821,N_18788);
nand U19379 (N_19379,N_18692,N_18739);
or U19380 (N_19380,N_18854,N_18986);
nor U19381 (N_19381,N_18480,N_19077);
or U19382 (N_19382,N_19153,N_18740);
nand U19383 (N_19383,N_18698,N_19078);
nor U19384 (N_19384,N_19161,N_19185);
nor U19385 (N_19385,N_19199,N_18501);
or U19386 (N_19386,N_18936,N_19074);
or U19387 (N_19387,N_18643,N_18819);
and U19388 (N_19388,N_18767,N_19110);
nor U19389 (N_19389,N_18405,N_18606);
nor U19390 (N_19390,N_18502,N_18855);
nand U19391 (N_19391,N_18709,N_18768);
and U19392 (N_19392,N_19080,N_18995);
nor U19393 (N_19393,N_18437,N_18836);
or U19394 (N_19394,N_18504,N_18560);
nand U19395 (N_19395,N_18645,N_18727);
or U19396 (N_19396,N_18623,N_18912);
and U19397 (N_19397,N_18417,N_18930);
and U19398 (N_19398,N_18511,N_18786);
nand U19399 (N_19399,N_18762,N_18482);
nand U19400 (N_19400,N_19065,N_18766);
nor U19401 (N_19401,N_19002,N_18980);
nor U19402 (N_19402,N_18751,N_18474);
nor U19403 (N_19403,N_18646,N_18838);
nand U19404 (N_19404,N_18563,N_18611);
and U19405 (N_19405,N_18895,N_18622);
and U19406 (N_19406,N_18902,N_18436);
and U19407 (N_19407,N_19032,N_18535);
nand U19408 (N_19408,N_18547,N_18701);
nand U19409 (N_19409,N_18507,N_18401);
nor U19410 (N_19410,N_18721,N_18945);
or U19411 (N_19411,N_19038,N_19166);
xor U19412 (N_19412,N_18820,N_18772);
or U19413 (N_19413,N_18850,N_19175);
nor U19414 (N_19414,N_18789,N_18973);
nor U19415 (N_19415,N_19163,N_18691);
and U19416 (N_19416,N_18882,N_18778);
or U19417 (N_19417,N_19133,N_18816);
or U19418 (N_19418,N_18544,N_18949);
or U19419 (N_19419,N_19134,N_18617);
nor U19420 (N_19420,N_18983,N_18430);
xnor U19421 (N_19421,N_19091,N_18593);
nand U19422 (N_19422,N_18413,N_18806);
nor U19423 (N_19423,N_18886,N_18867);
and U19424 (N_19424,N_18553,N_18718);
nand U19425 (N_19425,N_18584,N_18435);
nand U19426 (N_19426,N_18592,N_18830);
nor U19427 (N_19427,N_18948,N_18607);
or U19428 (N_19428,N_19043,N_18900);
and U19429 (N_19429,N_18908,N_18404);
nand U19430 (N_19430,N_19198,N_18428);
nand U19431 (N_19431,N_18402,N_18997);
or U19432 (N_19432,N_18976,N_19136);
nand U19433 (N_19433,N_18570,N_18891);
and U19434 (N_19434,N_19176,N_18928);
or U19435 (N_19435,N_18999,N_18532);
or U19436 (N_19436,N_18519,N_18887);
and U19437 (N_19437,N_18613,N_18966);
or U19438 (N_19438,N_19015,N_18469);
or U19439 (N_19439,N_18629,N_19189);
nor U19440 (N_19440,N_18517,N_18828);
and U19441 (N_19441,N_18859,N_18704);
nand U19442 (N_19442,N_18713,N_19008);
or U19443 (N_19443,N_19020,N_18885);
and U19444 (N_19444,N_19192,N_19109);
nand U19445 (N_19445,N_18953,N_18573);
nor U19446 (N_19446,N_18696,N_18541);
and U19447 (N_19447,N_19001,N_19061);
or U19448 (N_19448,N_18542,N_18869);
and U19449 (N_19449,N_18687,N_18784);
nor U19450 (N_19450,N_18926,N_19087);
and U19451 (N_19451,N_19098,N_18661);
and U19452 (N_19452,N_18910,N_18677);
and U19453 (N_19453,N_18780,N_18990);
or U19454 (N_19454,N_18567,N_18529);
or U19455 (N_19455,N_19018,N_18439);
nand U19456 (N_19456,N_19067,N_18911);
nand U19457 (N_19457,N_18551,N_18712);
xnor U19458 (N_19458,N_18906,N_19082);
nor U19459 (N_19459,N_18537,N_18937);
and U19460 (N_19460,N_18662,N_18889);
or U19461 (N_19461,N_19102,N_18683);
and U19462 (N_19462,N_18757,N_19105);
and U19463 (N_19463,N_19140,N_18856);
nand U19464 (N_19464,N_18832,N_18748);
nor U19465 (N_19465,N_18956,N_19177);
and U19466 (N_19466,N_19160,N_19195);
or U19467 (N_19467,N_18531,N_18452);
and U19468 (N_19468,N_19072,N_19186);
or U19469 (N_19469,N_19083,N_18528);
and U19470 (N_19470,N_19004,N_18479);
nor U19471 (N_19471,N_18561,N_19012);
nand U19472 (N_19472,N_18933,N_18760);
or U19473 (N_19473,N_19044,N_18922);
or U19474 (N_19474,N_18559,N_19174);
nor U19475 (N_19475,N_18871,N_18989);
and U19476 (N_19476,N_19108,N_18594);
and U19477 (N_19477,N_18568,N_19057);
and U19478 (N_19478,N_18946,N_18695);
nor U19479 (N_19479,N_18583,N_18686);
and U19480 (N_19480,N_18729,N_18795);
and U19481 (N_19481,N_18426,N_18722);
nand U19482 (N_19482,N_18931,N_18552);
or U19483 (N_19483,N_18486,N_19116);
or U19484 (N_19484,N_18460,N_19092);
or U19485 (N_19485,N_18427,N_18671);
nor U19486 (N_19486,N_18641,N_18589);
and U19487 (N_19487,N_19113,N_18653);
and U19488 (N_19488,N_18527,N_18951);
xnor U19489 (N_19489,N_18985,N_18635);
or U19490 (N_19490,N_19146,N_18655);
and U19491 (N_19491,N_19031,N_18771);
nor U19492 (N_19492,N_18898,N_18988);
nor U19493 (N_19493,N_18872,N_18459);
nand U19494 (N_19494,N_18445,N_18488);
nor U19495 (N_19495,N_19143,N_18719);
nor U19496 (N_19496,N_18745,N_19099);
or U19497 (N_19497,N_18642,N_19011);
or U19498 (N_19498,N_18765,N_19129);
nor U19499 (N_19499,N_18861,N_18652);
nor U19500 (N_19500,N_18516,N_18467);
or U19501 (N_19501,N_19071,N_18992);
nand U19502 (N_19502,N_19019,N_18518);
or U19503 (N_19503,N_18651,N_18710);
and U19504 (N_19504,N_18669,N_18848);
nor U19505 (N_19505,N_19159,N_19056);
or U19506 (N_19506,N_19155,N_18839);
and U19507 (N_19507,N_19046,N_18875);
nor U19508 (N_19508,N_18833,N_18500);
nand U19509 (N_19509,N_19137,N_18790);
nand U19510 (N_19510,N_18939,N_19169);
or U19511 (N_19511,N_19090,N_18858);
nor U19512 (N_19512,N_19173,N_18596);
and U19513 (N_19513,N_18604,N_18809);
and U19514 (N_19514,N_18512,N_19003);
or U19515 (N_19515,N_19130,N_19118);
and U19516 (N_19516,N_18650,N_18879);
or U19517 (N_19517,N_18656,N_18586);
nand U19518 (N_19518,N_18890,N_19037);
nand U19519 (N_19519,N_18490,N_19063);
nand U19520 (N_19520,N_18742,N_18600);
nor U19521 (N_19521,N_18960,N_18549);
nand U19522 (N_19522,N_19115,N_18755);
nor U19523 (N_19523,N_18590,N_18881);
and U19524 (N_19524,N_19172,N_18707);
nand U19525 (N_19525,N_18602,N_18779);
or U19526 (N_19526,N_18477,N_18905);
nand U19527 (N_19527,N_18804,N_18432);
nand U19528 (N_19528,N_19009,N_18448);
and U19529 (N_19529,N_19014,N_18458);
and U19530 (N_19530,N_18817,N_18892);
nand U19531 (N_19531,N_18664,N_19150);
or U19532 (N_19532,N_18638,N_19016);
nand U19533 (N_19533,N_18827,N_18914);
nand U19534 (N_19534,N_18723,N_18574);
nor U19535 (N_19535,N_18444,N_18864);
nor U19536 (N_19536,N_19073,N_18763);
nor U19537 (N_19537,N_18463,N_19148);
and U19538 (N_19538,N_18597,N_18416);
and U19539 (N_19539,N_18941,N_18744);
or U19540 (N_19540,N_18925,N_18608);
nor U19541 (N_19541,N_18415,N_19034);
or U19542 (N_19542,N_18705,N_18843);
xnor U19543 (N_19543,N_18619,N_18812);
and U19544 (N_19544,N_18564,N_18915);
nand U19545 (N_19545,N_18595,N_18453);
or U19546 (N_19546,N_19010,N_18783);
nand U19547 (N_19547,N_18648,N_18798);
nor U19548 (N_19548,N_18657,N_19028);
and U19549 (N_19549,N_18663,N_19106);
or U19550 (N_19550,N_18738,N_19013);
or U19551 (N_19551,N_18770,N_19188);
or U19552 (N_19552,N_18598,N_19111);
nor U19553 (N_19553,N_19095,N_18499);
nor U19554 (N_19554,N_18616,N_18734);
or U19555 (N_19555,N_18492,N_18538);
nand U19556 (N_19556,N_19094,N_18636);
nand U19557 (N_19557,N_18796,N_18706);
or U19558 (N_19558,N_18503,N_19023);
or U19559 (N_19559,N_19193,N_18659);
nor U19560 (N_19560,N_19024,N_19064);
nor U19561 (N_19561,N_18726,N_19006);
nand U19562 (N_19562,N_18725,N_18438);
nand U19563 (N_19563,N_18668,N_18572);
nor U19564 (N_19564,N_18781,N_18471);
nand U19565 (N_19565,N_18601,N_18546);
or U19566 (N_19566,N_18841,N_18576);
and U19567 (N_19567,N_18465,N_18508);
and U19568 (N_19568,N_18968,N_18750);
and U19569 (N_19569,N_18484,N_18470);
nand U19570 (N_19570,N_18408,N_19170);
and U19571 (N_19571,N_19122,N_18412);
nor U19572 (N_19572,N_19029,N_18977);
nand U19573 (N_19573,N_18690,N_18840);
or U19574 (N_19574,N_19000,N_18877);
nand U19575 (N_19575,N_19117,N_19157);
and U19576 (N_19576,N_19036,N_18679);
and U19577 (N_19577,N_19103,N_18562);
and U19578 (N_19578,N_18876,N_18411);
nand U19579 (N_19579,N_19050,N_18811);
nor U19580 (N_19580,N_19131,N_19197);
and U19581 (N_19581,N_18810,N_18403);
nor U19582 (N_19582,N_18523,N_19084);
nand U19583 (N_19583,N_18737,N_18682);
xor U19584 (N_19584,N_19127,N_18694);
nor U19585 (N_19585,N_18880,N_18724);
nor U19586 (N_19586,N_19104,N_18921);
or U19587 (N_19587,N_19196,N_19097);
or U19588 (N_19588,N_18431,N_18970);
nand U19589 (N_19589,N_18446,N_19059);
and U19590 (N_19590,N_18975,N_18752);
nor U19591 (N_19591,N_19179,N_19182);
nor U19592 (N_19592,N_18769,N_18844);
nor U19593 (N_19593,N_18955,N_18666);
or U19594 (N_19594,N_18853,N_18485);
nor U19595 (N_19595,N_18591,N_18736);
or U19596 (N_19596,N_18965,N_18702);
or U19597 (N_19597,N_18777,N_18631);
or U19598 (N_19598,N_18509,N_18924);
or U19599 (N_19599,N_19156,N_18846);
nand U19600 (N_19600,N_18735,N_18988);
and U19601 (N_19601,N_18532,N_19195);
and U19602 (N_19602,N_18405,N_19150);
nand U19603 (N_19603,N_19050,N_18768);
nor U19604 (N_19604,N_18853,N_19100);
and U19605 (N_19605,N_18408,N_19037);
nor U19606 (N_19606,N_19195,N_19140);
and U19607 (N_19607,N_19176,N_18634);
or U19608 (N_19608,N_19131,N_18845);
or U19609 (N_19609,N_19042,N_19052);
or U19610 (N_19610,N_19126,N_18615);
nand U19611 (N_19611,N_18537,N_18413);
nor U19612 (N_19612,N_19030,N_18625);
nor U19613 (N_19613,N_18509,N_18414);
nand U19614 (N_19614,N_18946,N_18709);
nor U19615 (N_19615,N_19116,N_18690);
nor U19616 (N_19616,N_18411,N_18925);
nor U19617 (N_19617,N_18959,N_18576);
nor U19618 (N_19618,N_18624,N_18809);
or U19619 (N_19619,N_19068,N_18790);
or U19620 (N_19620,N_18668,N_18918);
and U19621 (N_19621,N_18906,N_18579);
or U19622 (N_19622,N_18524,N_18454);
nand U19623 (N_19623,N_18806,N_18913);
nor U19624 (N_19624,N_18474,N_18857);
and U19625 (N_19625,N_18566,N_18738);
nor U19626 (N_19626,N_19060,N_18457);
or U19627 (N_19627,N_18421,N_18556);
nand U19628 (N_19628,N_19087,N_19084);
nand U19629 (N_19629,N_18754,N_18412);
or U19630 (N_19630,N_18984,N_19137);
or U19631 (N_19631,N_18892,N_18454);
nand U19632 (N_19632,N_18725,N_18745);
nor U19633 (N_19633,N_18924,N_18471);
and U19634 (N_19634,N_18469,N_18636);
nand U19635 (N_19635,N_18519,N_18547);
or U19636 (N_19636,N_18759,N_18423);
and U19637 (N_19637,N_18430,N_19067);
nor U19638 (N_19638,N_18703,N_19108);
nor U19639 (N_19639,N_19038,N_18419);
and U19640 (N_19640,N_19060,N_18870);
nor U19641 (N_19641,N_18751,N_18673);
or U19642 (N_19642,N_18549,N_19041);
nand U19643 (N_19643,N_19015,N_18437);
nand U19644 (N_19644,N_18779,N_18486);
nor U19645 (N_19645,N_18516,N_19029);
or U19646 (N_19646,N_18956,N_19166);
or U19647 (N_19647,N_18968,N_19184);
and U19648 (N_19648,N_18862,N_19109);
or U19649 (N_19649,N_18633,N_18758);
and U19650 (N_19650,N_19031,N_18789);
nor U19651 (N_19651,N_18547,N_18679);
or U19652 (N_19652,N_18781,N_18982);
nor U19653 (N_19653,N_19109,N_18694);
nand U19654 (N_19654,N_18980,N_18667);
or U19655 (N_19655,N_18904,N_18908);
nor U19656 (N_19656,N_18546,N_18653);
and U19657 (N_19657,N_18442,N_18637);
nor U19658 (N_19658,N_18869,N_18502);
nand U19659 (N_19659,N_19025,N_18743);
nor U19660 (N_19660,N_18956,N_18668);
nor U19661 (N_19661,N_18504,N_18762);
and U19662 (N_19662,N_18575,N_18697);
and U19663 (N_19663,N_19126,N_18475);
and U19664 (N_19664,N_18781,N_19169);
and U19665 (N_19665,N_18875,N_18407);
and U19666 (N_19666,N_18615,N_18408);
nand U19667 (N_19667,N_19048,N_18757);
nand U19668 (N_19668,N_19086,N_18409);
and U19669 (N_19669,N_19125,N_18971);
or U19670 (N_19670,N_18694,N_18627);
nor U19671 (N_19671,N_18759,N_18496);
and U19672 (N_19672,N_18747,N_19041);
and U19673 (N_19673,N_18929,N_18904);
nand U19674 (N_19674,N_18408,N_19150);
nor U19675 (N_19675,N_18484,N_19022);
nor U19676 (N_19676,N_18845,N_18550);
nand U19677 (N_19677,N_18570,N_19066);
and U19678 (N_19678,N_18807,N_18745);
nor U19679 (N_19679,N_18699,N_18912);
and U19680 (N_19680,N_18817,N_18987);
and U19681 (N_19681,N_18714,N_18509);
or U19682 (N_19682,N_19066,N_18704);
nor U19683 (N_19683,N_19180,N_18582);
nand U19684 (N_19684,N_19063,N_18781);
nor U19685 (N_19685,N_18699,N_19137);
nor U19686 (N_19686,N_18866,N_18731);
nor U19687 (N_19687,N_18735,N_18967);
or U19688 (N_19688,N_18900,N_18958);
or U19689 (N_19689,N_18683,N_19080);
nor U19690 (N_19690,N_18752,N_18527);
nand U19691 (N_19691,N_18419,N_18983);
or U19692 (N_19692,N_18533,N_19159);
or U19693 (N_19693,N_18415,N_18471);
nand U19694 (N_19694,N_18426,N_18444);
and U19695 (N_19695,N_19121,N_19177);
nor U19696 (N_19696,N_18448,N_19153);
or U19697 (N_19697,N_18767,N_19094);
and U19698 (N_19698,N_18729,N_19092);
or U19699 (N_19699,N_18986,N_19029);
or U19700 (N_19700,N_18989,N_18745);
or U19701 (N_19701,N_18974,N_18792);
nand U19702 (N_19702,N_18963,N_18951);
nand U19703 (N_19703,N_18732,N_18931);
and U19704 (N_19704,N_19093,N_18762);
and U19705 (N_19705,N_19167,N_19041);
and U19706 (N_19706,N_19044,N_19008);
nor U19707 (N_19707,N_18841,N_18865);
nand U19708 (N_19708,N_18733,N_18403);
and U19709 (N_19709,N_18894,N_18730);
nor U19710 (N_19710,N_19056,N_19154);
nand U19711 (N_19711,N_18565,N_18504);
and U19712 (N_19712,N_18910,N_18815);
or U19713 (N_19713,N_18786,N_18605);
and U19714 (N_19714,N_18831,N_18742);
or U19715 (N_19715,N_18904,N_18486);
nor U19716 (N_19716,N_18709,N_18575);
nor U19717 (N_19717,N_19100,N_18958);
and U19718 (N_19718,N_18642,N_18692);
and U19719 (N_19719,N_18402,N_19047);
nor U19720 (N_19720,N_18854,N_18719);
or U19721 (N_19721,N_18925,N_18753);
and U19722 (N_19722,N_18707,N_19104);
or U19723 (N_19723,N_18853,N_18456);
nor U19724 (N_19724,N_19110,N_18622);
nand U19725 (N_19725,N_18459,N_18737);
or U19726 (N_19726,N_18731,N_19044);
and U19727 (N_19727,N_18724,N_18681);
or U19728 (N_19728,N_18782,N_18656);
nor U19729 (N_19729,N_18849,N_18857);
or U19730 (N_19730,N_19170,N_19173);
nor U19731 (N_19731,N_18517,N_18974);
nor U19732 (N_19732,N_19188,N_18864);
nand U19733 (N_19733,N_18759,N_18563);
nand U19734 (N_19734,N_18793,N_18554);
or U19735 (N_19735,N_18522,N_19031);
nor U19736 (N_19736,N_19180,N_18581);
nor U19737 (N_19737,N_19021,N_18901);
nor U19738 (N_19738,N_18812,N_19195);
nor U19739 (N_19739,N_18527,N_18790);
and U19740 (N_19740,N_18483,N_18442);
nand U19741 (N_19741,N_18504,N_18751);
nand U19742 (N_19742,N_18646,N_18903);
nor U19743 (N_19743,N_18752,N_18670);
and U19744 (N_19744,N_19185,N_18578);
and U19745 (N_19745,N_18565,N_19178);
or U19746 (N_19746,N_18432,N_19187);
nand U19747 (N_19747,N_19134,N_18665);
nor U19748 (N_19748,N_18900,N_19090);
nor U19749 (N_19749,N_18623,N_18526);
nand U19750 (N_19750,N_18606,N_18636);
nand U19751 (N_19751,N_19014,N_19082);
or U19752 (N_19752,N_18799,N_18638);
nand U19753 (N_19753,N_18458,N_19067);
and U19754 (N_19754,N_18618,N_18694);
or U19755 (N_19755,N_19001,N_18703);
or U19756 (N_19756,N_19174,N_18939);
or U19757 (N_19757,N_19123,N_19150);
nand U19758 (N_19758,N_18521,N_19039);
nand U19759 (N_19759,N_18763,N_18439);
or U19760 (N_19760,N_18596,N_18595);
nand U19761 (N_19761,N_18446,N_19157);
and U19762 (N_19762,N_18877,N_19136);
or U19763 (N_19763,N_18992,N_18827);
nand U19764 (N_19764,N_18776,N_18411);
and U19765 (N_19765,N_19045,N_18778);
nor U19766 (N_19766,N_19062,N_18533);
nor U19767 (N_19767,N_18816,N_18627);
or U19768 (N_19768,N_18898,N_18423);
nor U19769 (N_19769,N_19049,N_19180);
nand U19770 (N_19770,N_19027,N_18614);
nor U19771 (N_19771,N_18586,N_18949);
or U19772 (N_19772,N_18750,N_18900);
and U19773 (N_19773,N_19100,N_18830);
nand U19774 (N_19774,N_18493,N_18961);
nor U19775 (N_19775,N_19139,N_18403);
nor U19776 (N_19776,N_18597,N_18420);
nand U19777 (N_19777,N_18794,N_18673);
and U19778 (N_19778,N_18959,N_18967);
or U19779 (N_19779,N_19122,N_18409);
and U19780 (N_19780,N_18880,N_18531);
and U19781 (N_19781,N_18786,N_19130);
or U19782 (N_19782,N_18968,N_18840);
nor U19783 (N_19783,N_18455,N_18673);
nor U19784 (N_19784,N_18908,N_19156);
nor U19785 (N_19785,N_18830,N_18845);
nor U19786 (N_19786,N_18898,N_18425);
nor U19787 (N_19787,N_19008,N_18785);
nand U19788 (N_19788,N_18623,N_18501);
and U19789 (N_19789,N_18935,N_19172);
or U19790 (N_19790,N_18608,N_18879);
nor U19791 (N_19791,N_18601,N_18429);
xnor U19792 (N_19792,N_18948,N_18968);
nand U19793 (N_19793,N_18516,N_18582);
or U19794 (N_19794,N_19049,N_18486);
and U19795 (N_19795,N_18502,N_18884);
and U19796 (N_19796,N_18625,N_19105);
nor U19797 (N_19797,N_18855,N_18969);
or U19798 (N_19798,N_19143,N_18582);
nand U19799 (N_19799,N_18688,N_18858);
and U19800 (N_19800,N_19051,N_19027);
or U19801 (N_19801,N_18456,N_19088);
or U19802 (N_19802,N_18629,N_18678);
or U19803 (N_19803,N_18996,N_18598);
nand U19804 (N_19804,N_18787,N_19072);
nor U19805 (N_19805,N_18834,N_18690);
nor U19806 (N_19806,N_18782,N_18853);
or U19807 (N_19807,N_19045,N_18981);
and U19808 (N_19808,N_18934,N_18925);
or U19809 (N_19809,N_18831,N_18602);
or U19810 (N_19810,N_19034,N_19126);
nor U19811 (N_19811,N_18537,N_18443);
nand U19812 (N_19812,N_19054,N_19042);
nand U19813 (N_19813,N_18882,N_18990);
and U19814 (N_19814,N_18867,N_18834);
nand U19815 (N_19815,N_18816,N_18538);
and U19816 (N_19816,N_18436,N_18818);
nand U19817 (N_19817,N_18420,N_19068);
and U19818 (N_19818,N_18611,N_18778);
nor U19819 (N_19819,N_18623,N_18967);
and U19820 (N_19820,N_18911,N_18868);
and U19821 (N_19821,N_18884,N_18741);
and U19822 (N_19822,N_18944,N_19178);
nand U19823 (N_19823,N_18480,N_18673);
and U19824 (N_19824,N_18918,N_18591);
or U19825 (N_19825,N_18448,N_18433);
nand U19826 (N_19826,N_19035,N_18797);
and U19827 (N_19827,N_18669,N_18821);
and U19828 (N_19828,N_18800,N_19083);
nand U19829 (N_19829,N_18886,N_18511);
nor U19830 (N_19830,N_18803,N_18707);
or U19831 (N_19831,N_18874,N_18784);
nand U19832 (N_19832,N_18538,N_18969);
nor U19833 (N_19833,N_19157,N_18812);
and U19834 (N_19834,N_18839,N_18590);
nor U19835 (N_19835,N_18766,N_18978);
and U19836 (N_19836,N_18407,N_19105);
or U19837 (N_19837,N_18407,N_19158);
or U19838 (N_19838,N_18432,N_18845);
nand U19839 (N_19839,N_18809,N_19016);
and U19840 (N_19840,N_18718,N_18777);
xnor U19841 (N_19841,N_18950,N_18552);
or U19842 (N_19842,N_19026,N_18839);
nor U19843 (N_19843,N_18468,N_18915);
or U19844 (N_19844,N_19179,N_19144);
nor U19845 (N_19845,N_18443,N_18885);
nor U19846 (N_19846,N_19122,N_18841);
nand U19847 (N_19847,N_18500,N_18703);
and U19848 (N_19848,N_18722,N_18916);
xnor U19849 (N_19849,N_18615,N_18956);
and U19850 (N_19850,N_18979,N_19170);
nand U19851 (N_19851,N_19058,N_18627);
and U19852 (N_19852,N_18671,N_18666);
or U19853 (N_19853,N_18985,N_18525);
and U19854 (N_19854,N_19190,N_18836);
and U19855 (N_19855,N_18493,N_19192);
nor U19856 (N_19856,N_18719,N_18676);
and U19857 (N_19857,N_19023,N_18575);
or U19858 (N_19858,N_19164,N_19097);
nor U19859 (N_19859,N_18696,N_18493);
or U19860 (N_19860,N_18877,N_19063);
or U19861 (N_19861,N_18932,N_18667);
nand U19862 (N_19862,N_18530,N_18800);
nor U19863 (N_19863,N_18806,N_19166);
nand U19864 (N_19864,N_18426,N_19102);
or U19865 (N_19865,N_18780,N_18925);
nor U19866 (N_19866,N_19090,N_18668);
or U19867 (N_19867,N_18647,N_18983);
nor U19868 (N_19868,N_18665,N_18801);
nor U19869 (N_19869,N_18832,N_18522);
and U19870 (N_19870,N_19036,N_18783);
nor U19871 (N_19871,N_19058,N_19031);
or U19872 (N_19872,N_19138,N_19015);
nand U19873 (N_19873,N_19078,N_18570);
nand U19874 (N_19874,N_18414,N_18464);
or U19875 (N_19875,N_18787,N_18755);
nand U19876 (N_19876,N_18525,N_18809);
nor U19877 (N_19877,N_18696,N_19176);
nand U19878 (N_19878,N_18624,N_18644);
and U19879 (N_19879,N_18415,N_19115);
xnor U19880 (N_19880,N_18426,N_19095);
or U19881 (N_19881,N_18726,N_18933);
nor U19882 (N_19882,N_18567,N_18485);
nand U19883 (N_19883,N_18990,N_18531);
nand U19884 (N_19884,N_18650,N_18506);
nor U19885 (N_19885,N_18500,N_19053);
or U19886 (N_19886,N_18809,N_18515);
and U19887 (N_19887,N_18857,N_18611);
or U19888 (N_19888,N_18922,N_18497);
nand U19889 (N_19889,N_18432,N_18869);
nor U19890 (N_19890,N_19072,N_19091);
nand U19891 (N_19891,N_18868,N_18567);
or U19892 (N_19892,N_18584,N_18480);
or U19893 (N_19893,N_19141,N_18476);
or U19894 (N_19894,N_19098,N_18927);
nand U19895 (N_19895,N_18623,N_18990);
nor U19896 (N_19896,N_18844,N_18608);
and U19897 (N_19897,N_18661,N_19078);
or U19898 (N_19898,N_18647,N_18871);
nand U19899 (N_19899,N_18570,N_19124);
and U19900 (N_19900,N_18575,N_19184);
or U19901 (N_19901,N_19199,N_18749);
nor U19902 (N_19902,N_19069,N_19022);
nor U19903 (N_19903,N_18802,N_19079);
nor U19904 (N_19904,N_18995,N_18758);
nand U19905 (N_19905,N_18964,N_19197);
nor U19906 (N_19906,N_19124,N_19194);
nor U19907 (N_19907,N_18639,N_18922);
nor U19908 (N_19908,N_18570,N_18840);
nand U19909 (N_19909,N_19001,N_18405);
or U19910 (N_19910,N_18530,N_19132);
and U19911 (N_19911,N_18619,N_18609);
or U19912 (N_19912,N_19147,N_18466);
or U19913 (N_19913,N_19196,N_19162);
nor U19914 (N_19914,N_18537,N_19139);
or U19915 (N_19915,N_18518,N_19089);
and U19916 (N_19916,N_19140,N_18592);
or U19917 (N_19917,N_18847,N_18931);
nor U19918 (N_19918,N_19126,N_18762);
or U19919 (N_19919,N_18533,N_18679);
or U19920 (N_19920,N_18411,N_18850);
or U19921 (N_19921,N_18939,N_19108);
and U19922 (N_19922,N_18703,N_18926);
nor U19923 (N_19923,N_18728,N_18566);
nand U19924 (N_19924,N_19144,N_19122);
and U19925 (N_19925,N_19011,N_19130);
or U19926 (N_19926,N_18598,N_18787);
nor U19927 (N_19927,N_18527,N_18992);
or U19928 (N_19928,N_19078,N_18427);
nor U19929 (N_19929,N_19019,N_18544);
nor U19930 (N_19930,N_18617,N_18898);
nor U19931 (N_19931,N_18685,N_18861);
or U19932 (N_19932,N_18545,N_18908);
or U19933 (N_19933,N_18932,N_18886);
or U19934 (N_19934,N_18433,N_18781);
or U19935 (N_19935,N_18951,N_19074);
or U19936 (N_19936,N_18812,N_18411);
or U19937 (N_19937,N_18611,N_19196);
and U19938 (N_19938,N_18930,N_18576);
nand U19939 (N_19939,N_18461,N_18866);
and U19940 (N_19940,N_19070,N_18891);
and U19941 (N_19941,N_19137,N_18484);
or U19942 (N_19942,N_19090,N_18749);
and U19943 (N_19943,N_18946,N_18793);
nand U19944 (N_19944,N_19039,N_18477);
nor U19945 (N_19945,N_18572,N_19184);
and U19946 (N_19946,N_19076,N_18719);
nor U19947 (N_19947,N_18550,N_18935);
and U19948 (N_19948,N_18441,N_19142);
nor U19949 (N_19949,N_19074,N_18797);
nor U19950 (N_19950,N_19196,N_18635);
nand U19951 (N_19951,N_18655,N_18445);
nor U19952 (N_19952,N_18572,N_18813);
and U19953 (N_19953,N_18512,N_18503);
or U19954 (N_19954,N_18870,N_19009);
and U19955 (N_19955,N_18636,N_18615);
nand U19956 (N_19956,N_18504,N_18679);
and U19957 (N_19957,N_18712,N_18442);
or U19958 (N_19958,N_18944,N_18838);
and U19959 (N_19959,N_18859,N_19099);
nand U19960 (N_19960,N_18498,N_19106);
and U19961 (N_19961,N_19171,N_18500);
and U19962 (N_19962,N_19105,N_18648);
nand U19963 (N_19963,N_18879,N_18485);
nor U19964 (N_19964,N_18563,N_18627);
and U19965 (N_19965,N_18458,N_18988);
xor U19966 (N_19966,N_19074,N_18756);
or U19967 (N_19967,N_19143,N_18857);
or U19968 (N_19968,N_18677,N_18965);
nand U19969 (N_19969,N_18874,N_18533);
nor U19970 (N_19970,N_18445,N_18465);
nor U19971 (N_19971,N_18661,N_18523);
nand U19972 (N_19972,N_18917,N_18618);
and U19973 (N_19973,N_18410,N_18596);
nor U19974 (N_19974,N_18943,N_18674);
or U19975 (N_19975,N_18732,N_18897);
nor U19976 (N_19976,N_18505,N_19033);
or U19977 (N_19977,N_18841,N_18477);
nand U19978 (N_19978,N_18984,N_18677);
nor U19979 (N_19979,N_18764,N_19106);
or U19980 (N_19980,N_18465,N_18609);
nand U19981 (N_19981,N_18704,N_18402);
nor U19982 (N_19982,N_18644,N_19025);
nand U19983 (N_19983,N_18474,N_18883);
nor U19984 (N_19984,N_18617,N_18495);
and U19985 (N_19985,N_18755,N_18753);
nand U19986 (N_19986,N_18428,N_19102);
nand U19987 (N_19987,N_18576,N_19178);
and U19988 (N_19988,N_18950,N_18705);
nor U19989 (N_19989,N_18682,N_19057);
and U19990 (N_19990,N_18483,N_18906);
nor U19991 (N_19991,N_18937,N_18564);
or U19992 (N_19992,N_18779,N_19056);
nor U19993 (N_19993,N_18706,N_18520);
nor U19994 (N_19994,N_19119,N_18837);
and U19995 (N_19995,N_18437,N_18954);
nand U19996 (N_19996,N_18721,N_19153);
nor U19997 (N_19997,N_18563,N_18935);
and U19998 (N_19998,N_18760,N_18742);
and U19999 (N_19999,N_18611,N_18764);
nand UO_0 (O_0,N_19338,N_19618);
nor UO_1 (O_1,N_19461,N_19918);
or UO_2 (O_2,N_19814,N_19352);
or UO_3 (O_3,N_19438,N_19307);
or UO_4 (O_4,N_19981,N_19697);
nand UO_5 (O_5,N_19721,N_19774);
or UO_6 (O_6,N_19512,N_19544);
and UO_7 (O_7,N_19932,N_19910);
nor UO_8 (O_8,N_19747,N_19773);
and UO_9 (O_9,N_19841,N_19432);
and UO_10 (O_10,N_19764,N_19920);
nand UO_11 (O_11,N_19681,N_19299);
nor UO_12 (O_12,N_19771,N_19958);
nor UO_13 (O_13,N_19809,N_19431);
or UO_14 (O_14,N_19703,N_19762);
or UO_15 (O_15,N_19673,N_19353);
nor UO_16 (O_16,N_19374,N_19200);
or UO_17 (O_17,N_19689,N_19882);
or UO_18 (O_18,N_19948,N_19643);
and UO_19 (O_19,N_19530,N_19381);
nor UO_20 (O_20,N_19439,N_19331);
or UO_21 (O_21,N_19633,N_19532);
nand UO_22 (O_22,N_19852,N_19785);
nor UO_23 (O_23,N_19607,N_19952);
nor UO_24 (O_24,N_19207,N_19216);
nand UO_25 (O_25,N_19498,N_19940);
nand UO_26 (O_26,N_19237,N_19434);
xnor UO_27 (O_27,N_19997,N_19863);
nor UO_28 (O_28,N_19848,N_19558);
or UO_29 (O_29,N_19402,N_19684);
and UO_30 (O_30,N_19383,N_19449);
nor UO_31 (O_31,N_19407,N_19750);
nor UO_32 (O_32,N_19358,N_19692);
or UO_33 (O_33,N_19775,N_19202);
and UO_34 (O_34,N_19741,N_19453);
nand UO_35 (O_35,N_19411,N_19536);
and UO_36 (O_36,N_19610,N_19831);
or UO_37 (O_37,N_19266,N_19350);
and UO_38 (O_38,N_19788,N_19570);
and UO_39 (O_39,N_19351,N_19529);
or UO_40 (O_40,N_19626,N_19543);
or UO_41 (O_41,N_19826,N_19465);
nand UO_42 (O_42,N_19317,N_19445);
nor UO_43 (O_43,N_19225,N_19608);
and UO_44 (O_44,N_19746,N_19421);
or UO_45 (O_45,N_19575,N_19221);
nor UO_46 (O_46,N_19694,N_19794);
nor UO_47 (O_47,N_19339,N_19629);
or UO_48 (O_48,N_19611,N_19229);
and UO_49 (O_49,N_19399,N_19691);
nor UO_50 (O_50,N_19325,N_19740);
xnor UO_51 (O_51,N_19437,N_19564);
nor UO_52 (O_52,N_19735,N_19727);
and UO_53 (O_53,N_19376,N_19938);
or UO_54 (O_54,N_19466,N_19479);
nor UO_55 (O_55,N_19447,N_19685);
and UO_56 (O_56,N_19667,N_19913);
and UO_57 (O_57,N_19666,N_19586);
xnor UO_58 (O_58,N_19969,N_19895);
or UO_59 (O_59,N_19812,N_19556);
and UO_60 (O_60,N_19683,N_19894);
and UO_61 (O_61,N_19855,N_19241);
and UO_62 (O_62,N_19695,N_19429);
and UO_63 (O_63,N_19323,N_19985);
and UO_64 (O_64,N_19600,N_19640);
nand UO_65 (O_65,N_19395,N_19250);
nand UO_66 (O_66,N_19451,N_19968);
nand UO_67 (O_67,N_19763,N_19336);
or UO_68 (O_68,N_19550,N_19373);
nor UO_69 (O_69,N_19546,N_19527);
and UO_70 (O_70,N_19833,N_19239);
nor UO_71 (O_71,N_19375,N_19211);
or UO_72 (O_72,N_19597,N_19859);
nor UO_73 (O_73,N_19242,N_19287);
and UO_74 (O_74,N_19810,N_19356);
or UO_75 (O_75,N_19616,N_19518);
nand UO_76 (O_76,N_19561,N_19917);
nor UO_77 (O_77,N_19269,N_19423);
nor UO_78 (O_78,N_19568,N_19717);
or UO_79 (O_79,N_19332,N_19819);
or UO_80 (O_80,N_19672,N_19631);
nor UO_81 (O_81,N_19410,N_19401);
or UO_82 (O_82,N_19502,N_19319);
and UO_83 (O_83,N_19745,N_19496);
or UO_84 (O_84,N_19405,N_19582);
or UO_85 (O_85,N_19776,N_19247);
nand UO_86 (O_86,N_19845,N_19452);
and UO_87 (O_87,N_19382,N_19286);
nand UO_88 (O_88,N_19253,N_19791);
and UO_89 (O_89,N_19680,N_19892);
nand UO_90 (O_90,N_19223,N_19738);
or UO_91 (O_91,N_19906,N_19951);
or UO_92 (O_92,N_19973,N_19688);
or UO_93 (O_93,N_19276,N_19379);
or UO_94 (O_94,N_19385,N_19988);
and UO_95 (O_95,N_19494,N_19240);
nand UO_96 (O_96,N_19283,N_19909);
and UO_97 (O_97,N_19469,N_19843);
nand UO_98 (O_98,N_19728,N_19823);
or UO_99 (O_99,N_19921,N_19765);
and UO_100 (O_100,N_19871,N_19285);
nor UO_101 (O_101,N_19712,N_19228);
and UO_102 (O_102,N_19937,N_19598);
and UO_103 (O_103,N_19982,N_19653);
or UO_104 (O_104,N_19236,N_19998);
nor UO_105 (O_105,N_19244,N_19210);
nand UO_106 (O_106,N_19368,N_19330);
and UO_107 (O_107,N_19388,N_19959);
or UO_108 (O_108,N_19687,N_19294);
or UO_109 (O_109,N_19567,N_19475);
nand UO_110 (O_110,N_19856,N_19533);
or UO_111 (O_111,N_19208,N_19357);
nor UO_112 (O_112,N_19448,N_19671);
xnor UO_113 (O_113,N_19866,N_19961);
or UO_114 (O_114,N_19457,N_19813);
or UO_115 (O_115,N_19908,N_19898);
or UO_116 (O_116,N_19682,N_19566);
nor UO_117 (O_117,N_19359,N_19486);
and UO_118 (O_118,N_19398,N_19679);
and UO_119 (O_119,N_19621,N_19590);
and UO_120 (O_120,N_19657,N_19493);
nor UO_121 (O_121,N_19989,N_19542);
nor UO_122 (O_122,N_19880,N_19537);
nor UO_123 (O_123,N_19509,N_19301);
or UO_124 (O_124,N_19868,N_19329);
or UO_125 (O_125,N_19847,N_19589);
nor UO_126 (O_126,N_19950,N_19955);
nand UO_127 (O_127,N_19815,N_19730);
and UO_128 (O_128,N_19779,N_19510);
nand UO_129 (O_129,N_19574,N_19651);
nand UO_130 (O_130,N_19525,N_19949);
or UO_131 (O_131,N_19974,N_19637);
or UO_132 (O_132,N_19860,N_19713);
nand UO_133 (O_133,N_19613,N_19770);
nand UO_134 (O_134,N_19956,N_19280);
or UO_135 (O_135,N_19739,N_19450);
nand UO_136 (O_136,N_19425,N_19553);
and UO_137 (O_137,N_19484,N_19252);
nand UO_138 (O_138,N_19977,N_19471);
nor UO_139 (O_139,N_19214,N_19840);
and UO_140 (O_140,N_19964,N_19805);
and UO_141 (O_141,N_19534,N_19768);
nand UO_142 (O_142,N_19372,N_19404);
nor UO_143 (O_143,N_19473,N_19944);
nor UO_144 (O_144,N_19737,N_19715);
and UO_145 (O_145,N_19295,N_19842);
or UO_146 (O_146,N_19234,N_19227);
and UO_147 (O_147,N_19936,N_19251);
or UO_148 (O_148,N_19665,N_19522);
and UO_149 (O_149,N_19702,N_19369);
nand UO_150 (O_150,N_19321,N_19462);
xor UO_151 (O_151,N_19606,N_19886);
nand UO_152 (O_152,N_19263,N_19261);
nor UO_153 (O_153,N_19226,N_19675);
nand UO_154 (O_154,N_19203,N_19857);
xor UO_155 (O_155,N_19719,N_19535);
nand UO_156 (O_156,N_19878,N_19858);
and UO_157 (O_157,N_19264,N_19443);
nor UO_158 (O_158,N_19759,N_19693);
nand UO_159 (O_159,N_19464,N_19980);
or UO_160 (O_160,N_19901,N_19889);
nand UO_161 (O_161,N_19274,N_19806);
and UO_162 (O_162,N_19864,N_19624);
and UO_163 (O_163,N_19990,N_19930);
and UO_164 (O_164,N_19839,N_19408);
and UO_165 (O_165,N_19515,N_19658);
and UO_166 (O_166,N_19259,N_19736);
nor UO_167 (O_167,N_19309,N_19914);
nor UO_168 (O_168,N_19361,N_19634);
nor UO_169 (O_169,N_19232,N_19347);
nand UO_170 (O_170,N_19994,N_19881);
nor UO_171 (O_171,N_19965,N_19504);
or UO_172 (O_172,N_19853,N_19472);
and UO_173 (O_173,N_19348,N_19639);
nand UO_174 (O_174,N_19904,N_19931);
nor UO_175 (O_175,N_19460,N_19476);
or UO_176 (O_176,N_19732,N_19816);
nor UO_177 (O_177,N_19862,N_19370);
and UO_178 (O_178,N_19322,N_19867);
nor UO_179 (O_179,N_19418,N_19844);
nand UO_180 (O_180,N_19755,N_19340);
nor UO_181 (O_181,N_19846,N_19400);
nand UO_182 (O_182,N_19344,N_19896);
or UO_183 (O_183,N_19617,N_19463);
and UO_184 (O_184,N_19632,N_19213);
nor UO_185 (O_185,N_19828,N_19824);
and UO_186 (O_186,N_19403,N_19686);
nand UO_187 (O_187,N_19209,N_19492);
or UO_188 (O_188,N_19726,N_19258);
nor UO_189 (O_189,N_19291,N_19387);
nand UO_190 (O_190,N_19754,N_19939);
nor UO_191 (O_191,N_19677,N_19579);
and UO_192 (O_192,N_19716,N_19678);
and UO_193 (O_193,N_19333,N_19326);
nor UO_194 (O_194,N_19507,N_19419);
and UO_195 (O_195,N_19636,N_19619);
nor UO_196 (O_196,N_19396,N_19524);
and UO_197 (O_197,N_19659,N_19832);
and UO_198 (O_198,N_19560,N_19327);
and UO_199 (O_199,N_19335,N_19924);
nor UO_200 (O_200,N_19531,N_19976);
or UO_201 (O_201,N_19623,N_19707);
and UO_202 (O_202,N_19305,N_19792);
nor UO_203 (O_203,N_19829,N_19706);
or UO_204 (O_204,N_19834,N_19497);
or UO_205 (O_205,N_19899,N_19999);
nand UO_206 (O_206,N_19354,N_19346);
and UO_207 (O_207,N_19793,N_19987);
and UO_208 (O_208,N_19238,N_19934);
and UO_209 (O_209,N_19729,N_19341);
nor UO_210 (O_210,N_19945,N_19800);
or UO_211 (O_211,N_19212,N_19386);
or UO_212 (O_212,N_19435,N_19430);
nor UO_213 (O_213,N_19569,N_19915);
or UO_214 (O_214,N_19257,N_19478);
or UO_215 (O_215,N_19433,N_19320);
nand UO_216 (O_216,N_19778,N_19797);
or UO_217 (O_217,N_19912,N_19282);
nand UO_218 (O_218,N_19483,N_19345);
and UO_219 (O_219,N_19256,N_19708);
nand UO_220 (O_220,N_19267,N_19663);
or UO_221 (O_221,N_19477,N_19907);
nand UO_222 (O_222,N_19565,N_19316);
and UO_223 (O_223,N_19393,N_19487);
nor UO_224 (O_224,N_19722,N_19514);
nand UO_225 (O_225,N_19397,N_19647);
or UO_226 (O_226,N_19204,N_19377);
nor UO_227 (O_227,N_19442,N_19887);
nand UO_228 (O_228,N_19709,N_19668);
nand UO_229 (O_229,N_19260,N_19300);
nand UO_230 (O_230,N_19235,N_19662);
or UO_231 (O_231,N_19482,N_19270);
nor UO_232 (O_232,N_19983,N_19869);
nand UO_233 (O_233,N_19620,N_19519);
nor UO_234 (O_234,N_19772,N_19748);
and UO_235 (O_235,N_19986,N_19246);
or UO_236 (O_236,N_19262,N_19935);
and UO_237 (O_237,N_19704,N_19562);
nor UO_238 (O_238,N_19872,N_19281);
nand UO_239 (O_239,N_19585,N_19766);
and UO_240 (O_240,N_19355,N_19803);
and UO_241 (O_241,N_19578,N_19539);
nor UO_242 (O_242,N_19314,N_19308);
nor UO_243 (O_243,N_19576,N_19441);
nor UO_244 (O_244,N_19919,N_19865);
nor UO_245 (O_245,N_19362,N_19495);
xnor UO_246 (O_246,N_19718,N_19470);
nand UO_247 (O_247,N_19724,N_19723);
and UO_248 (O_248,N_19655,N_19777);
nand UO_249 (O_249,N_19960,N_19962);
nor UO_250 (O_250,N_19409,N_19851);
and UO_251 (O_251,N_19415,N_19818);
and UO_252 (O_252,N_19584,N_19807);
nor UO_253 (O_253,N_19583,N_19516);
and UO_254 (O_254,N_19874,N_19966);
and UO_255 (O_255,N_19787,N_19389);
and UO_256 (O_256,N_19459,N_19557);
nor UO_257 (O_257,N_19233,N_19273);
and UO_258 (O_258,N_19652,N_19641);
nand UO_259 (O_259,N_19916,N_19897);
or UO_260 (O_260,N_19893,N_19753);
nor UO_261 (O_261,N_19523,N_19946);
or UO_262 (O_262,N_19628,N_19268);
nor UO_263 (O_263,N_19364,N_19751);
nand UO_264 (O_264,N_19972,N_19861);
nor UO_265 (O_265,N_19649,N_19888);
nor UO_266 (O_266,N_19521,N_19784);
or UO_267 (O_267,N_19601,N_19627);
nor UO_268 (O_268,N_19749,N_19954);
nor UO_269 (O_269,N_19885,N_19277);
and UO_270 (O_270,N_19547,N_19849);
nand UO_271 (O_271,N_19548,N_19508);
nand UO_272 (O_272,N_19603,N_19656);
nor UO_273 (O_273,N_19789,N_19201);
and UO_274 (O_274,N_19324,N_19761);
or UO_275 (O_275,N_19925,N_19363);
and UO_276 (O_276,N_19947,N_19436);
nor UO_277 (O_277,N_19555,N_19625);
and UO_278 (O_278,N_19455,N_19995);
or UO_279 (O_279,N_19752,N_19406);
nor UO_280 (O_280,N_19310,N_19481);
and UO_281 (O_281,N_19614,N_19661);
nand UO_282 (O_282,N_19854,N_19979);
or UO_283 (O_283,N_19725,N_19271);
or UO_284 (O_284,N_19249,N_19838);
or UO_285 (O_285,N_19343,N_19905);
or UO_286 (O_286,N_19798,N_19334);
nor UO_287 (O_287,N_19313,N_19743);
and UO_288 (O_288,N_19541,N_19890);
nand UO_289 (O_289,N_19390,N_19206);
nand UO_290 (O_290,N_19540,N_19922);
nor UO_291 (O_291,N_19581,N_19366);
nand UO_292 (O_292,N_19664,N_19231);
nand UO_293 (O_293,N_19414,N_19394);
or UO_294 (O_294,N_19837,N_19474);
nor UO_295 (O_295,N_19699,N_19255);
nand UO_296 (O_296,N_19417,N_19392);
or UO_297 (O_297,N_19714,N_19489);
nor UO_298 (O_298,N_19219,N_19248);
and UO_299 (O_299,N_19733,N_19505);
nand UO_300 (O_300,N_19923,N_19500);
nand UO_301 (O_301,N_19520,N_19337);
or UO_302 (O_302,N_19422,N_19488);
or UO_303 (O_303,N_19420,N_19278);
or UO_304 (O_304,N_19942,N_19468);
and UO_305 (O_305,N_19304,N_19825);
or UO_306 (O_306,N_19911,N_19424);
or UO_307 (O_307,N_19289,N_19467);
and UO_308 (O_308,N_19485,N_19349);
and UO_309 (O_309,N_19758,N_19821);
nor UO_310 (O_310,N_19941,N_19205);
nor UO_311 (O_311,N_19593,N_19676);
nand UO_312 (O_312,N_19594,N_19275);
nor UO_313 (O_313,N_19644,N_19587);
or UO_314 (O_314,N_19780,N_19552);
and UO_315 (O_315,N_19757,N_19298);
and UO_316 (O_316,N_19224,N_19710);
and UO_317 (O_317,N_19660,N_19360);
or UO_318 (O_318,N_19595,N_19744);
nand UO_319 (O_319,N_19836,N_19230);
nor UO_320 (O_320,N_19572,N_19967);
or UO_321 (O_321,N_19879,N_19440);
nand UO_322 (O_322,N_19491,N_19991);
nand UO_323 (O_323,N_19705,N_19254);
nor UO_324 (O_324,N_19975,N_19303);
and UO_325 (O_325,N_19284,N_19220);
or UO_326 (O_326,N_19596,N_19311);
and UO_327 (O_327,N_19517,N_19279);
and UO_328 (O_328,N_19963,N_19883);
or UO_329 (O_329,N_19698,N_19850);
xor UO_330 (O_330,N_19312,N_19996);
nand UO_331 (O_331,N_19795,N_19992);
nand UO_332 (O_332,N_19731,N_19215);
nand UO_333 (O_333,N_19884,N_19571);
nor UO_334 (O_334,N_19297,N_19622);
or UO_335 (O_335,N_19526,N_19957);
nor UO_336 (O_336,N_19559,N_19444);
nand UO_337 (O_337,N_19302,N_19769);
and UO_338 (O_338,N_19384,N_19528);
nor UO_339 (O_339,N_19767,N_19416);
nand UO_340 (O_340,N_19783,N_19635);
and UO_341 (O_341,N_19480,N_19782);
and UO_342 (O_342,N_19588,N_19808);
nor UO_343 (O_343,N_19820,N_19943);
or UO_344 (O_344,N_19760,N_19427);
nor UO_345 (O_345,N_19877,N_19612);
nor UO_346 (O_346,N_19218,N_19978);
nand UO_347 (O_347,N_19245,N_19993);
or UO_348 (O_348,N_19501,N_19563);
nand UO_349 (O_349,N_19630,N_19545);
nor UO_350 (O_350,N_19700,N_19876);
or UO_351 (O_351,N_19902,N_19822);
nor UO_352 (O_352,N_19875,N_19927);
nor UO_353 (O_353,N_19827,N_19506);
or UO_354 (O_354,N_19293,N_19511);
nor UO_355 (O_355,N_19645,N_19591);
nand UO_356 (O_356,N_19953,N_19642);
nor UO_357 (O_357,N_19426,N_19873);
nand UO_358 (O_358,N_19378,N_19801);
or UO_359 (O_359,N_19391,N_19243);
nor UO_360 (O_360,N_19292,N_19650);
nand UO_361 (O_361,N_19900,N_19781);
nand UO_362 (O_362,N_19638,N_19288);
xor UO_363 (O_363,N_19674,N_19971);
and UO_364 (O_364,N_19577,N_19811);
nor UO_365 (O_365,N_19367,N_19830);
or UO_366 (O_366,N_19646,N_19669);
and UO_367 (O_367,N_19296,N_19551);
or UO_368 (O_368,N_19933,N_19318);
and UO_369 (O_369,N_19615,N_19742);
nand UO_370 (O_370,N_19573,N_19428);
and UO_371 (O_371,N_19456,N_19580);
nor UO_372 (O_372,N_19928,N_19592);
or UO_373 (O_373,N_19599,N_19696);
or UO_374 (O_374,N_19891,N_19538);
or UO_375 (O_375,N_19654,N_19217);
or UO_376 (O_376,N_19648,N_19380);
and UO_377 (O_377,N_19602,N_19835);
nor UO_378 (O_378,N_19670,N_19817);
nor UO_379 (O_379,N_19458,N_19734);
and UO_380 (O_380,N_19756,N_19701);
nor UO_381 (O_381,N_19690,N_19604);
or UO_382 (O_382,N_19786,N_19984);
or UO_383 (O_383,N_19371,N_19454);
nand UO_384 (O_384,N_19903,N_19222);
nor UO_385 (O_385,N_19413,N_19804);
or UO_386 (O_386,N_19446,N_19315);
and UO_387 (O_387,N_19790,N_19870);
and UO_388 (O_388,N_19499,N_19272);
nor UO_389 (O_389,N_19265,N_19711);
and UO_390 (O_390,N_19513,N_19412);
or UO_391 (O_391,N_19796,N_19554);
nor UO_392 (O_392,N_19926,N_19970);
or UO_393 (O_393,N_19503,N_19609);
nor UO_394 (O_394,N_19342,N_19720);
and UO_395 (O_395,N_19328,N_19365);
and UO_396 (O_396,N_19490,N_19929);
nand UO_397 (O_397,N_19306,N_19605);
or UO_398 (O_398,N_19799,N_19549);
and UO_399 (O_399,N_19802,N_19290);
and UO_400 (O_400,N_19724,N_19991);
or UO_401 (O_401,N_19725,N_19342);
nor UO_402 (O_402,N_19371,N_19257);
nor UO_403 (O_403,N_19796,N_19456);
and UO_404 (O_404,N_19825,N_19735);
nand UO_405 (O_405,N_19803,N_19705);
nor UO_406 (O_406,N_19470,N_19214);
nand UO_407 (O_407,N_19972,N_19657);
nor UO_408 (O_408,N_19500,N_19435);
and UO_409 (O_409,N_19587,N_19571);
nand UO_410 (O_410,N_19458,N_19779);
nand UO_411 (O_411,N_19528,N_19981);
or UO_412 (O_412,N_19975,N_19299);
and UO_413 (O_413,N_19872,N_19477);
xor UO_414 (O_414,N_19755,N_19553);
nand UO_415 (O_415,N_19930,N_19631);
nand UO_416 (O_416,N_19748,N_19893);
or UO_417 (O_417,N_19693,N_19812);
nor UO_418 (O_418,N_19892,N_19814);
nand UO_419 (O_419,N_19833,N_19949);
and UO_420 (O_420,N_19766,N_19777);
xor UO_421 (O_421,N_19320,N_19299);
nor UO_422 (O_422,N_19288,N_19697);
nor UO_423 (O_423,N_19308,N_19887);
and UO_424 (O_424,N_19305,N_19370);
xor UO_425 (O_425,N_19488,N_19460);
or UO_426 (O_426,N_19255,N_19706);
and UO_427 (O_427,N_19619,N_19662);
nand UO_428 (O_428,N_19360,N_19824);
nand UO_429 (O_429,N_19464,N_19782);
or UO_430 (O_430,N_19349,N_19703);
and UO_431 (O_431,N_19839,N_19580);
nand UO_432 (O_432,N_19514,N_19361);
nand UO_433 (O_433,N_19935,N_19264);
and UO_434 (O_434,N_19410,N_19221);
or UO_435 (O_435,N_19938,N_19348);
nand UO_436 (O_436,N_19473,N_19684);
nand UO_437 (O_437,N_19978,N_19616);
or UO_438 (O_438,N_19771,N_19528);
and UO_439 (O_439,N_19201,N_19586);
and UO_440 (O_440,N_19240,N_19790);
or UO_441 (O_441,N_19805,N_19326);
and UO_442 (O_442,N_19760,N_19749);
or UO_443 (O_443,N_19767,N_19325);
nor UO_444 (O_444,N_19493,N_19756);
or UO_445 (O_445,N_19492,N_19681);
or UO_446 (O_446,N_19853,N_19463);
and UO_447 (O_447,N_19928,N_19417);
nand UO_448 (O_448,N_19707,N_19348);
nor UO_449 (O_449,N_19608,N_19411);
and UO_450 (O_450,N_19909,N_19218);
and UO_451 (O_451,N_19500,N_19660);
or UO_452 (O_452,N_19630,N_19440);
or UO_453 (O_453,N_19451,N_19687);
nor UO_454 (O_454,N_19395,N_19257);
or UO_455 (O_455,N_19988,N_19746);
nor UO_456 (O_456,N_19906,N_19699);
nor UO_457 (O_457,N_19636,N_19672);
and UO_458 (O_458,N_19345,N_19880);
or UO_459 (O_459,N_19858,N_19396);
or UO_460 (O_460,N_19732,N_19537);
nand UO_461 (O_461,N_19419,N_19726);
nand UO_462 (O_462,N_19638,N_19907);
and UO_463 (O_463,N_19596,N_19975);
or UO_464 (O_464,N_19360,N_19866);
nor UO_465 (O_465,N_19977,N_19293);
nand UO_466 (O_466,N_19273,N_19232);
nor UO_467 (O_467,N_19269,N_19503);
nor UO_468 (O_468,N_19747,N_19466);
nor UO_469 (O_469,N_19939,N_19362);
or UO_470 (O_470,N_19309,N_19267);
or UO_471 (O_471,N_19667,N_19977);
nand UO_472 (O_472,N_19609,N_19671);
and UO_473 (O_473,N_19774,N_19571);
and UO_474 (O_474,N_19840,N_19282);
and UO_475 (O_475,N_19300,N_19918);
or UO_476 (O_476,N_19787,N_19425);
nand UO_477 (O_477,N_19766,N_19224);
nor UO_478 (O_478,N_19675,N_19246);
or UO_479 (O_479,N_19747,N_19673);
and UO_480 (O_480,N_19873,N_19279);
or UO_481 (O_481,N_19682,N_19661);
nor UO_482 (O_482,N_19825,N_19363);
or UO_483 (O_483,N_19737,N_19460);
nor UO_484 (O_484,N_19817,N_19969);
nor UO_485 (O_485,N_19361,N_19353);
or UO_486 (O_486,N_19839,N_19594);
nand UO_487 (O_487,N_19801,N_19896);
and UO_488 (O_488,N_19768,N_19928);
and UO_489 (O_489,N_19697,N_19358);
nand UO_490 (O_490,N_19933,N_19842);
or UO_491 (O_491,N_19703,N_19875);
nor UO_492 (O_492,N_19841,N_19842);
or UO_493 (O_493,N_19753,N_19650);
and UO_494 (O_494,N_19807,N_19495);
nand UO_495 (O_495,N_19345,N_19669);
nor UO_496 (O_496,N_19576,N_19496);
nand UO_497 (O_497,N_19559,N_19404);
nand UO_498 (O_498,N_19530,N_19603);
nand UO_499 (O_499,N_19716,N_19765);
or UO_500 (O_500,N_19276,N_19951);
or UO_501 (O_501,N_19201,N_19304);
nand UO_502 (O_502,N_19445,N_19640);
or UO_503 (O_503,N_19389,N_19683);
nand UO_504 (O_504,N_19513,N_19859);
and UO_505 (O_505,N_19788,N_19977);
nand UO_506 (O_506,N_19801,N_19200);
nor UO_507 (O_507,N_19417,N_19637);
or UO_508 (O_508,N_19325,N_19987);
or UO_509 (O_509,N_19479,N_19846);
and UO_510 (O_510,N_19504,N_19922);
or UO_511 (O_511,N_19548,N_19247);
and UO_512 (O_512,N_19337,N_19355);
nand UO_513 (O_513,N_19725,N_19662);
or UO_514 (O_514,N_19628,N_19712);
nand UO_515 (O_515,N_19530,N_19489);
and UO_516 (O_516,N_19769,N_19608);
or UO_517 (O_517,N_19565,N_19761);
nand UO_518 (O_518,N_19296,N_19730);
nor UO_519 (O_519,N_19897,N_19914);
or UO_520 (O_520,N_19207,N_19723);
or UO_521 (O_521,N_19521,N_19529);
nor UO_522 (O_522,N_19268,N_19378);
nand UO_523 (O_523,N_19730,N_19763);
or UO_524 (O_524,N_19717,N_19581);
nor UO_525 (O_525,N_19878,N_19574);
nand UO_526 (O_526,N_19577,N_19761);
or UO_527 (O_527,N_19533,N_19246);
nor UO_528 (O_528,N_19840,N_19314);
nor UO_529 (O_529,N_19282,N_19372);
or UO_530 (O_530,N_19290,N_19536);
nor UO_531 (O_531,N_19402,N_19586);
nand UO_532 (O_532,N_19466,N_19874);
nand UO_533 (O_533,N_19946,N_19699);
nor UO_534 (O_534,N_19304,N_19718);
or UO_535 (O_535,N_19928,N_19720);
nor UO_536 (O_536,N_19651,N_19799);
nor UO_537 (O_537,N_19682,N_19623);
nor UO_538 (O_538,N_19624,N_19551);
and UO_539 (O_539,N_19399,N_19684);
nor UO_540 (O_540,N_19887,N_19413);
nor UO_541 (O_541,N_19305,N_19663);
and UO_542 (O_542,N_19662,N_19350);
nor UO_543 (O_543,N_19732,N_19573);
or UO_544 (O_544,N_19470,N_19795);
or UO_545 (O_545,N_19244,N_19711);
nor UO_546 (O_546,N_19570,N_19706);
nor UO_547 (O_547,N_19773,N_19393);
or UO_548 (O_548,N_19790,N_19399);
nor UO_549 (O_549,N_19362,N_19308);
nor UO_550 (O_550,N_19645,N_19513);
and UO_551 (O_551,N_19311,N_19381);
and UO_552 (O_552,N_19650,N_19956);
nor UO_553 (O_553,N_19904,N_19691);
or UO_554 (O_554,N_19952,N_19973);
and UO_555 (O_555,N_19657,N_19442);
nor UO_556 (O_556,N_19518,N_19865);
nor UO_557 (O_557,N_19871,N_19347);
nor UO_558 (O_558,N_19714,N_19602);
nor UO_559 (O_559,N_19809,N_19254);
nor UO_560 (O_560,N_19406,N_19202);
nor UO_561 (O_561,N_19446,N_19580);
and UO_562 (O_562,N_19667,N_19319);
and UO_563 (O_563,N_19924,N_19353);
nand UO_564 (O_564,N_19827,N_19535);
nor UO_565 (O_565,N_19798,N_19552);
or UO_566 (O_566,N_19844,N_19458);
nand UO_567 (O_567,N_19861,N_19545);
nand UO_568 (O_568,N_19348,N_19688);
xor UO_569 (O_569,N_19610,N_19295);
nand UO_570 (O_570,N_19770,N_19515);
and UO_571 (O_571,N_19516,N_19895);
and UO_572 (O_572,N_19755,N_19965);
or UO_573 (O_573,N_19808,N_19596);
and UO_574 (O_574,N_19613,N_19264);
nor UO_575 (O_575,N_19275,N_19856);
nand UO_576 (O_576,N_19235,N_19931);
or UO_577 (O_577,N_19997,N_19717);
nand UO_578 (O_578,N_19275,N_19954);
nand UO_579 (O_579,N_19690,N_19740);
nor UO_580 (O_580,N_19716,N_19411);
and UO_581 (O_581,N_19653,N_19958);
nor UO_582 (O_582,N_19513,N_19635);
nand UO_583 (O_583,N_19314,N_19927);
or UO_584 (O_584,N_19754,N_19654);
and UO_585 (O_585,N_19458,N_19878);
and UO_586 (O_586,N_19806,N_19253);
nand UO_587 (O_587,N_19621,N_19807);
or UO_588 (O_588,N_19500,N_19559);
nand UO_589 (O_589,N_19997,N_19256);
xor UO_590 (O_590,N_19602,N_19823);
nor UO_591 (O_591,N_19661,N_19444);
nand UO_592 (O_592,N_19272,N_19870);
or UO_593 (O_593,N_19227,N_19944);
xnor UO_594 (O_594,N_19567,N_19466);
and UO_595 (O_595,N_19957,N_19699);
nor UO_596 (O_596,N_19453,N_19299);
nand UO_597 (O_597,N_19738,N_19702);
xnor UO_598 (O_598,N_19526,N_19691);
nor UO_599 (O_599,N_19282,N_19737);
nand UO_600 (O_600,N_19873,N_19892);
or UO_601 (O_601,N_19529,N_19723);
nand UO_602 (O_602,N_19533,N_19848);
nor UO_603 (O_603,N_19226,N_19512);
nor UO_604 (O_604,N_19453,N_19672);
and UO_605 (O_605,N_19978,N_19217);
or UO_606 (O_606,N_19746,N_19570);
or UO_607 (O_607,N_19575,N_19802);
nor UO_608 (O_608,N_19291,N_19654);
nor UO_609 (O_609,N_19355,N_19402);
nand UO_610 (O_610,N_19562,N_19469);
nand UO_611 (O_611,N_19646,N_19330);
or UO_612 (O_612,N_19912,N_19582);
nand UO_613 (O_613,N_19406,N_19682);
nand UO_614 (O_614,N_19425,N_19333);
xnor UO_615 (O_615,N_19944,N_19994);
and UO_616 (O_616,N_19340,N_19961);
nand UO_617 (O_617,N_19811,N_19244);
nand UO_618 (O_618,N_19536,N_19919);
or UO_619 (O_619,N_19765,N_19633);
nor UO_620 (O_620,N_19514,N_19835);
and UO_621 (O_621,N_19596,N_19259);
or UO_622 (O_622,N_19389,N_19967);
or UO_623 (O_623,N_19603,N_19749);
nand UO_624 (O_624,N_19485,N_19505);
or UO_625 (O_625,N_19450,N_19836);
or UO_626 (O_626,N_19972,N_19896);
and UO_627 (O_627,N_19767,N_19300);
and UO_628 (O_628,N_19644,N_19410);
nand UO_629 (O_629,N_19323,N_19220);
nor UO_630 (O_630,N_19989,N_19783);
nand UO_631 (O_631,N_19654,N_19812);
nor UO_632 (O_632,N_19842,N_19720);
nor UO_633 (O_633,N_19795,N_19449);
nand UO_634 (O_634,N_19586,N_19709);
and UO_635 (O_635,N_19398,N_19612);
nor UO_636 (O_636,N_19965,N_19229);
nand UO_637 (O_637,N_19566,N_19752);
or UO_638 (O_638,N_19382,N_19823);
nor UO_639 (O_639,N_19710,N_19630);
or UO_640 (O_640,N_19201,N_19784);
and UO_641 (O_641,N_19463,N_19854);
nand UO_642 (O_642,N_19762,N_19420);
or UO_643 (O_643,N_19966,N_19577);
nor UO_644 (O_644,N_19399,N_19441);
nor UO_645 (O_645,N_19273,N_19676);
or UO_646 (O_646,N_19719,N_19735);
nand UO_647 (O_647,N_19862,N_19740);
nor UO_648 (O_648,N_19473,N_19457);
or UO_649 (O_649,N_19353,N_19656);
and UO_650 (O_650,N_19938,N_19414);
nand UO_651 (O_651,N_19429,N_19675);
nor UO_652 (O_652,N_19986,N_19515);
nor UO_653 (O_653,N_19623,N_19869);
nand UO_654 (O_654,N_19648,N_19368);
nand UO_655 (O_655,N_19205,N_19569);
nor UO_656 (O_656,N_19431,N_19616);
or UO_657 (O_657,N_19815,N_19729);
nor UO_658 (O_658,N_19524,N_19287);
nor UO_659 (O_659,N_19260,N_19399);
and UO_660 (O_660,N_19663,N_19973);
and UO_661 (O_661,N_19379,N_19696);
nor UO_662 (O_662,N_19243,N_19838);
or UO_663 (O_663,N_19897,N_19676);
nor UO_664 (O_664,N_19485,N_19345);
nor UO_665 (O_665,N_19527,N_19435);
nor UO_666 (O_666,N_19644,N_19571);
nor UO_667 (O_667,N_19286,N_19471);
nand UO_668 (O_668,N_19485,N_19915);
nor UO_669 (O_669,N_19418,N_19667);
nor UO_670 (O_670,N_19605,N_19664);
or UO_671 (O_671,N_19751,N_19444);
and UO_672 (O_672,N_19534,N_19955);
or UO_673 (O_673,N_19359,N_19847);
nor UO_674 (O_674,N_19536,N_19789);
or UO_675 (O_675,N_19958,N_19749);
nor UO_676 (O_676,N_19271,N_19219);
nor UO_677 (O_677,N_19714,N_19831);
or UO_678 (O_678,N_19385,N_19953);
nand UO_679 (O_679,N_19972,N_19819);
or UO_680 (O_680,N_19900,N_19647);
nand UO_681 (O_681,N_19727,N_19626);
and UO_682 (O_682,N_19364,N_19594);
nor UO_683 (O_683,N_19383,N_19385);
or UO_684 (O_684,N_19590,N_19783);
and UO_685 (O_685,N_19256,N_19989);
or UO_686 (O_686,N_19309,N_19751);
nor UO_687 (O_687,N_19613,N_19424);
nor UO_688 (O_688,N_19358,N_19539);
or UO_689 (O_689,N_19401,N_19248);
nand UO_690 (O_690,N_19607,N_19506);
and UO_691 (O_691,N_19683,N_19328);
and UO_692 (O_692,N_19828,N_19426);
and UO_693 (O_693,N_19331,N_19540);
and UO_694 (O_694,N_19510,N_19200);
or UO_695 (O_695,N_19352,N_19312);
and UO_696 (O_696,N_19899,N_19945);
or UO_697 (O_697,N_19612,N_19466);
nand UO_698 (O_698,N_19925,N_19352);
or UO_699 (O_699,N_19341,N_19941);
or UO_700 (O_700,N_19596,N_19884);
nor UO_701 (O_701,N_19243,N_19248);
nor UO_702 (O_702,N_19814,N_19598);
or UO_703 (O_703,N_19490,N_19964);
nand UO_704 (O_704,N_19898,N_19949);
nand UO_705 (O_705,N_19463,N_19879);
nand UO_706 (O_706,N_19883,N_19377);
and UO_707 (O_707,N_19406,N_19237);
nand UO_708 (O_708,N_19431,N_19686);
and UO_709 (O_709,N_19201,N_19718);
and UO_710 (O_710,N_19429,N_19300);
or UO_711 (O_711,N_19881,N_19953);
and UO_712 (O_712,N_19791,N_19778);
and UO_713 (O_713,N_19414,N_19952);
nor UO_714 (O_714,N_19255,N_19412);
nor UO_715 (O_715,N_19538,N_19765);
and UO_716 (O_716,N_19266,N_19360);
and UO_717 (O_717,N_19236,N_19572);
nor UO_718 (O_718,N_19374,N_19275);
and UO_719 (O_719,N_19339,N_19526);
and UO_720 (O_720,N_19613,N_19489);
or UO_721 (O_721,N_19468,N_19469);
nand UO_722 (O_722,N_19378,N_19508);
and UO_723 (O_723,N_19548,N_19946);
nor UO_724 (O_724,N_19241,N_19853);
nor UO_725 (O_725,N_19247,N_19900);
or UO_726 (O_726,N_19728,N_19987);
nand UO_727 (O_727,N_19658,N_19573);
and UO_728 (O_728,N_19387,N_19700);
nand UO_729 (O_729,N_19285,N_19595);
nand UO_730 (O_730,N_19275,N_19421);
and UO_731 (O_731,N_19332,N_19745);
nand UO_732 (O_732,N_19422,N_19476);
nand UO_733 (O_733,N_19898,N_19381);
or UO_734 (O_734,N_19852,N_19251);
or UO_735 (O_735,N_19566,N_19739);
and UO_736 (O_736,N_19704,N_19869);
nor UO_737 (O_737,N_19928,N_19597);
and UO_738 (O_738,N_19629,N_19816);
and UO_739 (O_739,N_19990,N_19764);
nor UO_740 (O_740,N_19919,N_19810);
and UO_741 (O_741,N_19733,N_19612);
and UO_742 (O_742,N_19802,N_19640);
nand UO_743 (O_743,N_19323,N_19247);
or UO_744 (O_744,N_19377,N_19988);
nand UO_745 (O_745,N_19441,N_19221);
or UO_746 (O_746,N_19570,N_19202);
or UO_747 (O_747,N_19495,N_19519);
nor UO_748 (O_748,N_19665,N_19363);
nor UO_749 (O_749,N_19870,N_19851);
and UO_750 (O_750,N_19439,N_19607);
nand UO_751 (O_751,N_19812,N_19731);
nor UO_752 (O_752,N_19566,N_19993);
nand UO_753 (O_753,N_19734,N_19437);
or UO_754 (O_754,N_19965,N_19985);
nand UO_755 (O_755,N_19243,N_19533);
nor UO_756 (O_756,N_19763,N_19791);
nor UO_757 (O_757,N_19678,N_19352);
nor UO_758 (O_758,N_19925,N_19622);
nor UO_759 (O_759,N_19434,N_19479);
and UO_760 (O_760,N_19517,N_19858);
xnor UO_761 (O_761,N_19692,N_19209);
and UO_762 (O_762,N_19782,N_19351);
nand UO_763 (O_763,N_19321,N_19430);
nor UO_764 (O_764,N_19424,N_19627);
or UO_765 (O_765,N_19317,N_19833);
and UO_766 (O_766,N_19269,N_19312);
or UO_767 (O_767,N_19991,N_19477);
nand UO_768 (O_768,N_19572,N_19664);
and UO_769 (O_769,N_19579,N_19733);
nor UO_770 (O_770,N_19994,N_19731);
or UO_771 (O_771,N_19212,N_19965);
or UO_772 (O_772,N_19992,N_19752);
and UO_773 (O_773,N_19624,N_19214);
nor UO_774 (O_774,N_19519,N_19539);
nand UO_775 (O_775,N_19790,N_19928);
or UO_776 (O_776,N_19871,N_19785);
or UO_777 (O_777,N_19532,N_19729);
or UO_778 (O_778,N_19354,N_19410);
nand UO_779 (O_779,N_19690,N_19203);
nor UO_780 (O_780,N_19618,N_19666);
xor UO_781 (O_781,N_19237,N_19307);
nand UO_782 (O_782,N_19809,N_19948);
nand UO_783 (O_783,N_19364,N_19724);
and UO_784 (O_784,N_19418,N_19244);
and UO_785 (O_785,N_19373,N_19756);
nand UO_786 (O_786,N_19272,N_19662);
nor UO_787 (O_787,N_19229,N_19475);
or UO_788 (O_788,N_19660,N_19602);
and UO_789 (O_789,N_19556,N_19277);
or UO_790 (O_790,N_19549,N_19713);
and UO_791 (O_791,N_19437,N_19682);
or UO_792 (O_792,N_19213,N_19503);
or UO_793 (O_793,N_19889,N_19347);
nor UO_794 (O_794,N_19683,N_19289);
nor UO_795 (O_795,N_19508,N_19941);
and UO_796 (O_796,N_19213,N_19773);
nor UO_797 (O_797,N_19563,N_19420);
nand UO_798 (O_798,N_19318,N_19275);
and UO_799 (O_799,N_19368,N_19886);
nand UO_800 (O_800,N_19822,N_19659);
or UO_801 (O_801,N_19692,N_19232);
and UO_802 (O_802,N_19331,N_19840);
and UO_803 (O_803,N_19222,N_19691);
nand UO_804 (O_804,N_19382,N_19348);
or UO_805 (O_805,N_19422,N_19851);
nand UO_806 (O_806,N_19255,N_19278);
nor UO_807 (O_807,N_19289,N_19868);
and UO_808 (O_808,N_19374,N_19814);
nand UO_809 (O_809,N_19953,N_19391);
or UO_810 (O_810,N_19357,N_19481);
nor UO_811 (O_811,N_19889,N_19617);
nor UO_812 (O_812,N_19690,N_19891);
nand UO_813 (O_813,N_19290,N_19945);
and UO_814 (O_814,N_19502,N_19899);
nand UO_815 (O_815,N_19927,N_19800);
nor UO_816 (O_816,N_19219,N_19790);
and UO_817 (O_817,N_19990,N_19382);
nor UO_818 (O_818,N_19316,N_19902);
nor UO_819 (O_819,N_19403,N_19525);
or UO_820 (O_820,N_19636,N_19807);
and UO_821 (O_821,N_19862,N_19816);
or UO_822 (O_822,N_19260,N_19860);
nor UO_823 (O_823,N_19328,N_19950);
and UO_824 (O_824,N_19576,N_19241);
or UO_825 (O_825,N_19601,N_19488);
and UO_826 (O_826,N_19680,N_19295);
nor UO_827 (O_827,N_19657,N_19785);
and UO_828 (O_828,N_19908,N_19414);
nor UO_829 (O_829,N_19227,N_19257);
nor UO_830 (O_830,N_19347,N_19920);
nand UO_831 (O_831,N_19600,N_19267);
nor UO_832 (O_832,N_19855,N_19771);
and UO_833 (O_833,N_19292,N_19389);
xor UO_834 (O_834,N_19742,N_19690);
nor UO_835 (O_835,N_19376,N_19568);
nand UO_836 (O_836,N_19246,N_19264);
nand UO_837 (O_837,N_19737,N_19379);
or UO_838 (O_838,N_19586,N_19877);
or UO_839 (O_839,N_19520,N_19363);
and UO_840 (O_840,N_19860,N_19475);
or UO_841 (O_841,N_19426,N_19664);
or UO_842 (O_842,N_19336,N_19714);
nand UO_843 (O_843,N_19686,N_19311);
nor UO_844 (O_844,N_19288,N_19613);
nand UO_845 (O_845,N_19567,N_19318);
and UO_846 (O_846,N_19992,N_19430);
nand UO_847 (O_847,N_19488,N_19902);
nor UO_848 (O_848,N_19585,N_19650);
nand UO_849 (O_849,N_19398,N_19282);
or UO_850 (O_850,N_19540,N_19955);
and UO_851 (O_851,N_19645,N_19619);
nor UO_852 (O_852,N_19809,N_19868);
and UO_853 (O_853,N_19481,N_19852);
nor UO_854 (O_854,N_19260,N_19213);
and UO_855 (O_855,N_19260,N_19238);
nor UO_856 (O_856,N_19225,N_19720);
or UO_857 (O_857,N_19804,N_19837);
or UO_858 (O_858,N_19885,N_19499);
nor UO_859 (O_859,N_19580,N_19448);
nor UO_860 (O_860,N_19444,N_19793);
nor UO_861 (O_861,N_19236,N_19419);
and UO_862 (O_862,N_19933,N_19415);
nand UO_863 (O_863,N_19460,N_19665);
nand UO_864 (O_864,N_19955,N_19370);
and UO_865 (O_865,N_19365,N_19698);
or UO_866 (O_866,N_19378,N_19394);
nand UO_867 (O_867,N_19780,N_19938);
and UO_868 (O_868,N_19297,N_19723);
and UO_869 (O_869,N_19563,N_19723);
nand UO_870 (O_870,N_19425,N_19409);
nand UO_871 (O_871,N_19813,N_19652);
nor UO_872 (O_872,N_19480,N_19671);
or UO_873 (O_873,N_19212,N_19242);
nand UO_874 (O_874,N_19296,N_19307);
and UO_875 (O_875,N_19635,N_19632);
nor UO_876 (O_876,N_19897,N_19617);
nor UO_877 (O_877,N_19497,N_19737);
and UO_878 (O_878,N_19396,N_19319);
or UO_879 (O_879,N_19835,N_19948);
and UO_880 (O_880,N_19921,N_19494);
and UO_881 (O_881,N_19388,N_19326);
nand UO_882 (O_882,N_19404,N_19412);
and UO_883 (O_883,N_19365,N_19587);
nand UO_884 (O_884,N_19410,N_19295);
or UO_885 (O_885,N_19288,N_19973);
nand UO_886 (O_886,N_19736,N_19380);
nand UO_887 (O_887,N_19759,N_19872);
nor UO_888 (O_888,N_19995,N_19765);
nor UO_889 (O_889,N_19578,N_19860);
and UO_890 (O_890,N_19594,N_19573);
nor UO_891 (O_891,N_19731,N_19935);
and UO_892 (O_892,N_19879,N_19930);
nand UO_893 (O_893,N_19285,N_19924);
and UO_894 (O_894,N_19793,N_19327);
nand UO_895 (O_895,N_19893,N_19462);
or UO_896 (O_896,N_19239,N_19550);
and UO_897 (O_897,N_19283,N_19962);
or UO_898 (O_898,N_19707,N_19303);
nor UO_899 (O_899,N_19782,N_19950);
nor UO_900 (O_900,N_19327,N_19483);
and UO_901 (O_901,N_19871,N_19445);
nor UO_902 (O_902,N_19681,N_19810);
and UO_903 (O_903,N_19490,N_19852);
and UO_904 (O_904,N_19852,N_19892);
nand UO_905 (O_905,N_19822,N_19804);
and UO_906 (O_906,N_19398,N_19803);
and UO_907 (O_907,N_19687,N_19501);
nor UO_908 (O_908,N_19283,N_19752);
nand UO_909 (O_909,N_19480,N_19987);
nor UO_910 (O_910,N_19212,N_19534);
or UO_911 (O_911,N_19543,N_19589);
or UO_912 (O_912,N_19639,N_19890);
or UO_913 (O_913,N_19258,N_19729);
nand UO_914 (O_914,N_19982,N_19345);
nand UO_915 (O_915,N_19536,N_19292);
nand UO_916 (O_916,N_19792,N_19972);
or UO_917 (O_917,N_19305,N_19977);
nor UO_918 (O_918,N_19361,N_19690);
or UO_919 (O_919,N_19806,N_19221);
nand UO_920 (O_920,N_19320,N_19755);
nor UO_921 (O_921,N_19226,N_19818);
and UO_922 (O_922,N_19593,N_19229);
or UO_923 (O_923,N_19216,N_19514);
nor UO_924 (O_924,N_19616,N_19606);
nor UO_925 (O_925,N_19874,N_19448);
or UO_926 (O_926,N_19629,N_19432);
and UO_927 (O_927,N_19531,N_19319);
or UO_928 (O_928,N_19978,N_19726);
nand UO_929 (O_929,N_19704,N_19650);
nand UO_930 (O_930,N_19994,N_19239);
or UO_931 (O_931,N_19571,N_19728);
or UO_932 (O_932,N_19575,N_19346);
nor UO_933 (O_933,N_19901,N_19721);
nor UO_934 (O_934,N_19332,N_19711);
or UO_935 (O_935,N_19692,N_19835);
nor UO_936 (O_936,N_19728,N_19721);
and UO_937 (O_937,N_19249,N_19957);
nand UO_938 (O_938,N_19493,N_19790);
or UO_939 (O_939,N_19631,N_19245);
or UO_940 (O_940,N_19247,N_19882);
or UO_941 (O_941,N_19986,N_19602);
nand UO_942 (O_942,N_19413,N_19417);
and UO_943 (O_943,N_19269,N_19239);
nor UO_944 (O_944,N_19567,N_19564);
or UO_945 (O_945,N_19770,N_19721);
nor UO_946 (O_946,N_19694,N_19825);
and UO_947 (O_947,N_19284,N_19829);
nand UO_948 (O_948,N_19378,N_19670);
or UO_949 (O_949,N_19679,N_19946);
nand UO_950 (O_950,N_19797,N_19335);
nor UO_951 (O_951,N_19798,N_19293);
or UO_952 (O_952,N_19209,N_19726);
and UO_953 (O_953,N_19914,N_19316);
and UO_954 (O_954,N_19529,N_19672);
and UO_955 (O_955,N_19923,N_19433);
or UO_956 (O_956,N_19897,N_19742);
and UO_957 (O_957,N_19838,N_19636);
nand UO_958 (O_958,N_19634,N_19289);
and UO_959 (O_959,N_19564,N_19949);
or UO_960 (O_960,N_19447,N_19637);
nand UO_961 (O_961,N_19314,N_19389);
nand UO_962 (O_962,N_19673,N_19997);
or UO_963 (O_963,N_19380,N_19728);
and UO_964 (O_964,N_19755,N_19788);
nor UO_965 (O_965,N_19650,N_19212);
and UO_966 (O_966,N_19274,N_19835);
and UO_967 (O_967,N_19509,N_19630);
nand UO_968 (O_968,N_19710,N_19998);
nand UO_969 (O_969,N_19862,N_19667);
nand UO_970 (O_970,N_19850,N_19978);
nor UO_971 (O_971,N_19912,N_19839);
nor UO_972 (O_972,N_19694,N_19423);
nor UO_973 (O_973,N_19527,N_19273);
or UO_974 (O_974,N_19958,N_19849);
and UO_975 (O_975,N_19686,N_19756);
nand UO_976 (O_976,N_19995,N_19519);
and UO_977 (O_977,N_19471,N_19229);
nand UO_978 (O_978,N_19255,N_19927);
nor UO_979 (O_979,N_19495,N_19469);
and UO_980 (O_980,N_19409,N_19353);
or UO_981 (O_981,N_19911,N_19647);
and UO_982 (O_982,N_19478,N_19785);
and UO_983 (O_983,N_19736,N_19956);
and UO_984 (O_984,N_19461,N_19689);
nor UO_985 (O_985,N_19798,N_19280);
nor UO_986 (O_986,N_19513,N_19637);
nand UO_987 (O_987,N_19610,N_19279);
and UO_988 (O_988,N_19556,N_19661);
nand UO_989 (O_989,N_19854,N_19439);
or UO_990 (O_990,N_19253,N_19352);
and UO_991 (O_991,N_19887,N_19799);
nor UO_992 (O_992,N_19439,N_19646);
or UO_993 (O_993,N_19403,N_19741);
and UO_994 (O_994,N_19279,N_19607);
nor UO_995 (O_995,N_19690,N_19923);
or UO_996 (O_996,N_19710,N_19202);
or UO_997 (O_997,N_19984,N_19365);
and UO_998 (O_998,N_19211,N_19830);
or UO_999 (O_999,N_19539,N_19911);
nand UO_1000 (O_1000,N_19886,N_19830);
nand UO_1001 (O_1001,N_19238,N_19332);
nand UO_1002 (O_1002,N_19257,N_19398);
or UO_1003 (O_1003,N_19477,N_19511);
and UO_1004 (O_1004,N_19864,N_19522);
and UO_1005 (O_1005,N_19791,N_19922);
and UO_1006 (O_1006,N_19711,N_19467);
nor UO_1007 (O_1007,N_19440,N_19438);
nand UO_1008 (O_1008,N_19281,N_19934);
or UO_1009 (O_1009,N_19496,N_19657);
nand UO_1010 (O_1010,N_19863,N_19666);
nor UO_1011 (O_1011,N_19504,N_19348);
nor UO_1012 (O_1012,N_19707,N_19518);
and UO_1013 (O_1013,N_19841,N_19229);
nand UO_1014 (O_1014,N_19343,N_19413);
and UO_1015 (O_1015,N_19667,N_19857);
nand UO_1016 (O_1016,N_19772,N_19369);
and UO_1017 (O_1017,N_19490,N_19501);
or UO_1018 (O_1018,N_19482,N_19462);
and UO_1019 (O_1019,N_19913,N_19523);
nor UO_1020 (O_1020,N_19498,N_19245);
nor UO_1021 (O_1021,N_19395,N_19295);
nor UO_1022 (O_1022,N_19885,N_19317);
nor UO_1023 (O_1023,N_19724,N_19462);
nor UO_1024 (O_1024,N_19436,N_19786);
nand UO_1025 (O_1025,N_19267,N_19291);
nand UO_1026 (O_1026,N_19898,N_19543);
nand UO_1027 (O_1027,N_19287,N_19310);
and UO_1028 (O_1028,N_19751,N_19796);
nor UO_1029 (O_1029,N_19618,N_19340);
nor UO_1030 (O_1030,N_19402,N_19459);
nor UO_1031 (O_1031,N_19321,N_19850);
and UO_1032 (O_1032,N_19956,N_19667);
or UO_1033 (O_1033,N_19568,N_19768);
and UO_1034 (O_1034,N_19540,N_19771);
nand UO_1035 (O_1035,N_19486,N_19341);
or UO_1036 (O_1036,N_19989,N_19847);
and UO_1037 (O_1037,N_19977,N_19456);
nor UO_1038 (O_1038,N_19654,N_19916);
nand UO_1039 (O_1039,N_19324,N_19657);
or UO_1040 (O_1040,N_19534,N_19569);
nor UO_1041 (O_1041,N_19468,N_19907);
and UO_1042 (O_1042,N_19573,N_19311);
nand UO_1043 (O_1043,N_19451,N_19203);
nor UO_1044 (O_1044,N_19379,N_19714);
nand UO_1045 (O_1045,N_19588,N_19256);
nand UO_1046 (O_1046,N_19547,N_19359);
nand UO_1047 (O_1047,N_19807,N_19887);
nand UO_1048 (O_1048,N_19743,N_19762);
and UO_1049 (O_1049,N_19206,N_19852);
and UO_1050 (O_1050,N_19511,N_19668);
nor UO_1051 (O_1051,N_19798,N_19672);
nand UO_1052 (O_1052,N_19700,N_19671);
nand UO_1053 (O_1053,N_19722,N_19446);
and UO_1054 (O_1054,N_19267,N_19250);
nand UO_1055 (O_1055,N_19372,N_19681);
or UO_1056 (O_1056,N_19358,N_19519);
nand UO_1057 (O_1057,N_19216,N_19302);
nand UO_1058 (O_1058,N_19237,N_19599);
and UO_1059 (O_1059,N_19608,N_19571);
and UO_1060 (O_1060,N_19969,N_19761);
and UO_1061 (O_1061,N_19435,N_19366);
nor UO_1062 (O_1062,N_19540,N_19912);
nor UO_1063 (O_1063,N_19673,N_19961);
nand UO_1064 (O_1064,N_19965,N_19499);
nor UO_1065 (O_1065,N_19417,N_19257);
or UO_1066 (O_1066,N_19622,N_19788);
nor UO_1067 (O_1067,N_19218,N_19543);
nor UO_1068 (O_1068,N_19409,N_19349);
nor UO_1069 (O_1069,N_19360,N_19677);
and UO_1070 (O_1070,N_19825,N_19512);
or UO_1071 (O_1071,N_19422,N_19503);
nand UO_1072 (O_1072,N_19325,N_19209);
and UO_1073 (O_1073,N_19532,N_19206);
nor UO_1074 (O_1074,N_19640,N_19609);
nand UO_1075 (O_1075,N_19970,N_19777);
and UO_1076 (O_1076,N_19273,N_19834);
or UO_1077 (O_1077,N_19657,N_19344);
nor UO_1078 (O_1078,N_19379,N_19694);
xnor UO_1079 (O_1079,N_19468,N_19755);
nor UO_1080 (O_1080,N_19884,N_19430);
and UO_1081 (O_1081,N_19730,N_19958);
or UO_1082 (O_1082,N_19875,N_19258);
and UO_1083 (O_1083,N_19582,N_19771);
nor UO_1084 (O_1084,N_19533,N_19313);
nor UO_1085 (O_1085,N_19352,N_19326);
and UO_1086 (O_1086,N_19429,N_19459);
nor UO_1087 (O_1087,N_19754,N_19963);
xor UO_1088 (O_1088,N_19846,N_19305);
nor UO_1089 (O_1089,N_19494,N_19482);
nand UO_1090 (O_1090,N_19545,N_19958);
and UO_1091 (O_1091,N_19210,N_19248);
or UO_1092 (O_1092,N_19974,N_19416);
nand UO_1093 (O_1093,N_19851,N_19513);
and UO_1094 (O_1094,N_19758,N_19354);
nand UO_1095 (O_1095,N_19904,N_19496);
and UO_1096 (O_1096,N_19562,N_19777);
and UO_1097 (O_1097,N_19713,N_19724);
nand UO_1098 (O_1098,N_19831,N_19373);
nor UO_1099 (O_1099,N_19708,N_19812);
or UO_1100 (O_1100,N_19506,N_19278);
or UO_1101 (O_1101,N_19437,N_19554);
and UO_1102 (O_1102,N_19942,N_19478);
nor UO_1103 (O_1103,N_19556,N_19878);
nand UO_1104 (O_1104,N_19878,N_19266);
or UO_1105 (O_1105,N_19526,N_19822);
and UO_1106 (O_1106,N_19967,N_19581);
nor UO_1107 (O_1107,N_19856,N_19650);
and UO_1108 (O_1108,N_19514,N_19358);
or UO_1109 (O_1109,N_19731,N_19313);
and UO_1110 (O_1110,N_19807,N_19388);
and UO_1111 (O_1111,N_19843,N_19228);
nand UO_1112 (O_1112,N_19419,N_19242);
and UO_1113 (O_1113,N_19423,N_19219);
and UO_1114 (O_1114,N_19376,N_19203);
nand UO_1115 (O_1115,N_19398,N_19802);
or UO_1116 (O_1116,N_19352,N_19469);
and UO_1117 (O_1117,N_19713,N_19474);
and UO_1118 (O_1118,N_19421,N_19943);
nor UO_1119 (O_1119,N_19899,N_19599);
nand UO_1120 (O_1120,N_19681,N_19882);
and UO_1121 (O_1121,N_19335,N_19806);
nor UO_1122 (O_1122,N_19275,N_19753);
and UO_1123 (O_1123,N_19602,N_19216);
and UO_1124 (O_1124,N_19521,N_19308);
and UO_1125 (O_1125,N_19421,N_19485);
nand UO_1126 (O_1126,N_19849,N_19968);
and UO_1127 (O_1127,N_19986,N_19918);
nor UO_1128 (O_1128,N_19361,N_19259);
nand UO_1129 (O_1129,N_19621,N_19928);
and UO_1130 (O_1130,N_19251,N_19946);
or UO_1131 (O_1131,N_19398,N_19303);
or UO_1132 (O_1132,N_19309,N_19417);
and UO_1133 (O_1133,N_19246,N_19320);
or UO_1134 (O_1134,N_19894,N_19701);
and UO_1135 (O_1135,N_19662,N_19553);
and UO_1136 (O_1136,N_19772,N_19802);
or UO_1137 (O_1137,N_19456,N_19863);
and UO_1138 (O_1138,N_19255,N_19899);
nor UO_1139 (O_1139,N_19513,N_19302);
or UO_1140 (O_1140,N_19257,N_19387);
nor UO_1141 (O_1141,N_19864,N_19660);
nand UO_1142 (O_1142,N_19490,N_19796);
and UO_1143 (O_1143,N_19205,N_19555);
nor UO_1144 (O_1144,N_19486,N_19669);
and UO_1145 (O_1145,N_19346,N_19288);
nor UO_1146 (O_1146,N_19365,N_19412);
nor UO_1147 (O_1147,N_19994,N_19559);
or UO_1148 (O_1148,N_19857,N_19768);
nand UO_1149 (O_1149,N_19615,N_19542);
nand UO_1150 (O_1150,N_19788,N_19292);
nand UO_1151 (O_1151,N_19305,N_19853);
nor UO_1152 (O_1152,N_19825,N_19753);
nor UO_1153 (O_1153,N_19668,N_19866);
and UO_1154 (O_1154,N_19452,N_19466);
or UO_1155 (O_1155,N_19467,N_19327);
and UO_1156 (O_1156,N_19421,N_19634);
or UO_1157 (O_1157,N_19948,N_19580);
xor UO_1158 (O_1158,N_19269,N_19691);
or UO_1159 (O_1159,N_19803,N_19892);
nor UO_1160 (O_1160,N_19243,N_19671);
and UO_1161 (O_1161,N_19525,N_19569);
and UO_1162 (O_1162,N_19781,N_19854);
xor UO_1163 (O_1163,N_19884,N_19502);
nor UO_1164 (O_1164,N_19776,N_19700);
nor UO_1165 (O_1165,N_19335,N_19234);
and UO_1166 (O_1166,N_19382,N_19322);
or UO_1167 (O_1167,N_19505,N_19370);
and UO_1168 (O_1168,N_19667,N_19619);
nand UO_1169 (O_1169,N_19865,N_19802);
nand UO_1170 (O_1170,N_19464,N_19443);
or UO_1171 (O_1171,N_19822,N_19533);
nand UO_1172 (O_1172,N_19260,N_19994);
or UO_1173 (O_1173,N_19365,N_19287);
and UO_1174 (O_1174,N_19619,N_19341);
and UO_1175 (O_1175,N_19287,N_19875);
nor UO_1176 (O_1176,N_19661,N_19330);
nand UO_1177 (O_1177,N_19981,N_19510);
nor UO_1178 (O_1178,N_19468,N_19309);
nand UO_1179 (O_1179,N_19723,N_19482);
and UO_1180 (O_1180,N_19286,N_19577);
nor UO_1181 (O_1181,N_19394,N_19907);
and UO_1182 (O_1182,N_19448,N_19915);
or UO_1183 (O_1183,N_19875,N_19901);
and UO_1184 (O_1184,N_19440,N_19911);
and UO_1185 (O_1185,N_19256,N_19211);
or UO_1186 (O_1186,N_19268,N_19287);
and UO_1187 (O_1187,N_19242,N_19330);
nor UO_1188 (O_1188,N_19753,N_19849);
or UO_1189 (O_1189,N_19550,N_19500);
and UO_1190 (O_1190,N_19742,N_19529);
nand UO_1191 (O_1191,N_19632,N_19955);
nand UO_1192 (O_1192,N_19415,N_19635);
nor UO_1193 (O_1193,N_19504,N_19644);
nand UO_1194 (O_1194,N_19549,N_19995);
nand UO_1195 (O_1195,N_19650,N_19845);
nor UO_1196 (O_1196,N_19577,N_19200);
nand UO_1197 (O_1197,N_19887,N_19605);
and UO_1198 (O_1198,N_19897,N_19229);
or UO_1199 (O_1199,N_19217,N_19375);
nor UO_1200 (O_1200,N_19307,N_19865);
or UO_1201 (O_1201,N_19731,N_19945);
or UO_1202 (O_1202,N_19240,N_19250);
or UO_1203 (O_1203,N_19780,N_19709);
and UO_1204 (O_1204,N_19725,N_19674);
or UO_1205 (O_1205,N_19207,N_19699);
nand UO_1206 (O_1206,N_19681,N_19945);
nor UO_1207 (O_1207,N_19714,N_19317);
or UO_1208 (O_1208,N_19471,N_19698);
nand UO_1209 (O_1209,N_19695,N_19604);
and UO_1210 (O_1210,N_19783,N_19586);
and UO_1211 (O_1211,N_19666,N_19415);
or UO_1212 (O_1212,N_19669,N_19467);
or UO_1213 (O_1213,N_19713,N_19556);
nor UO_1214 (O_1214,N_19558,N_19811);
nor UO_1215 (O_1215,N_19452,N_19595);
nor UO_1216 (O_1216,N_19360,N_19656);
xnor UO_1217 (O_1217,N_19874,N_19224);
or UO_1218 (O_1218,N_19967,N_19402);
nand UO_1219 (O_1219,N_19992,N_19693);
and UO_1220 (O_1220,N_19310,N_19245);
or UO_1221 (O_1221,N_19323,N_19337);
nor UO_1222 (O_1222,N_19909,N_19690);
or UO_1223 (O_1223,N_19417,N_19613);
nand UO_1224 (O_1224,N_19612,N_19903);
or UO_1225 (O_1225,N_19398,N_19675);
nand UO_1226 (O_1226,N_19258,N_19601);
nand UO_1227 (O_1227,N_19515,N_19269);
nor UO_1228 (O_1228,N_19554,N_19785);
and UO_1229 (O_1229,N_19389,N_19476);
or UO_1230 (O_1230,N_19313,N_19262);
or UO_1231 (O_1231,N_19778,N_19269);
or UO_1232 (O_1232,N_19994,N_19675);
or UO_1233 (O_1233,N_19332,N_19702);
and UO_1234 (O_1234,N_19733,N_19864);
and UO_1235 (O_1235,N_19482,N_19929);
nor UO_1236 (O_1236,N_19677,N_19388);
nand UO_1237 (O_1237,N_19763,N_19444);
or UO_1238 (O_1238,N_19885,N_19293);
nor UO_1239 (O_1239,N_19527,N_19541);
nor UO_1240 (O_1240,N_19997,N_19787);
and UO_1241 (O_1241,N_19974,N_19883);
nor UO_1242 (O_1242,N_19427,N_19387);
and UO_1243 (O_1243,N_19245,N_19772);
and UO_1244 (O_1244,N_19568,N_19319);
or UO_1245 (O_1245,N_19806,N_19821);
or UO_1246 (O_1246,N_19237,N_19412);
or UO_1247 (O_1247,N_19346,N_19463);
nand UO_1248 (O_1248,N_19452,N_19228);
nand UO_1249 (O_1249,N_19536,N_19891);
or UO_1250 (O_1250,N_19212,N_19807);
nor UO_1251 (O_1251,N_19460,N_19214);
nand UO_1252 (O_1252,N_19817,N_19404);
or UO_1253 (O_1253,N_19664,N_19845);
nand UO_1254 (O_1254,N_19567,N_19558);
nand UO_1255 (O_1255,N_19911,N_19530);
nand UO_1256 (O_1256,N_19522,N_19731);
or UO_1257 (O_1257,N_19939,N_19895);
or UO_1258 (O_1258,N_19223,N_19402);
nor UO_1259 (O_1259,N_19325,N_19931);
xor UO_1260 (O_1260,N_19568,N_19902);
nor UO_1261 (O_1261,N_19880,N_19418);
and UO_1262 (O_1262,N_19544,N_19809);
nor UO_1263 (O_1263,N_19521,N_19590);
nand UO_1264 (O_1264,N_19858,N_19734);
nand UO_1265 (O_1265,N_19505,N_19266);
and UO_1266 (O_1266,N_19817,N_19375);
nor UO_1267 (O_1267,N_19987,N_19803);
and UO_1268 (O_1268,N_19223,N_19551);
and UO_1269 (O_1269,N_19637,N_19917);
nor UO_1270 (O_1270,N_19951,N_19769);
nor UO_1271 (O_1271,N_19566,N_19660);
nand UO_1272 (O_1272,N_19570,N_19383);
or UO_1273 (O_1273,N_19965,N_19737);
or UO_1274 (O_1274,N_19638,N_19440);
nor UO_1275 (O_1275,N_19713,N_19619);
nor UO_1276 (O_1276,N_19567,N_19739);
and UO_1277 (O_1277,N_19684,N_19318);
and UO_1278 (O_1278,N_19943,N_19937);
or UO_1279 (O_1279,N_19808,N_19747);
nand UO_1280 (O_1280,N_19942,N_19861);
and UO_1281 (O_1281,N_19495,N_19705);
and UO_1282 (O_1282,N_19985,N_19284);
nand UO_1283 (O_1283,N_19474,N_19448);
nand UO_1284 (O_1284,N_19282,N_19336);
nand UO_1285 (O_1285,N_19232,N_19630);
nor UO_1286 (O_1286,N_19375,N_19394);
and UO_1287 (O_1287,N_19820,N_19635);
nand UO_1288 (O_1288,N_19733,N_19740);
nor UO_1289 (O_1289,N_19252,N_19768);
nand UO_1290 (O_1290,N_19713,N_19693);
nor UO_1291 (O_1291,N_19480,N_19633);
nand UO_1292 (O_1292,N_19423,N_19943);
nand UO_1293 (O_1293,N_19267,N_19503);
nand UO_1294 (O_1294,N_19561,N_19286);
and UO_1295 (O_1295,N_19344,N_19615);
nor UO_1296 (O_1296,N_19292,N_19278);
or UO_1297 (O_1297,N_19517,N_19278);
and UO_1298 (O_1298,N_19742,N_19547);
and UO_1299 (O_1299,N_19950,N_19512);
and UO_1300 (O_1300,N_19684,N_19227);
nor UO_1301 (O_1301,N_19704,N_19994);
and UO_1302 (O_1302,N_19932,N_19875);
or UO_1303 (O_1303,N_19610,N_19855);
nor UO_1304 (O_1304,N_19726,N_19393);
and UO_1305 (O_1305,N_19256,N_19242);
and UO_1306 (O_1306,N_19841,N_19570);
nand UO_1307 (O_1307,N_19809,N_19353);
and UO_1308 (O_1308,N_19374,N_19932);
nor UO_1309 (O_1309,N_19401,N_19259);
and UO_1310 (O_1310,N_19303,N_19529);
and UO_1311 (O_1311,N_19726,N_19914);
and UO_1312 (O_1312,N_19376,N_19580);
or UO_1313 (O_1313,N_19253,N_19764);
nor UO_1314 (O_1314,N_19353,N_19431);
and UO_1315 (O_1315,N_19972,N_19419);
nor UO_1316 (O_1316,N_19304,N_19920);
or UO_1317 (O_1317,N_19570,N_19479);
nor UO_1318 (O_1318,N_19992,N_19485);
nor UO_1319 (O_1319,N_19923,N_19590);
xor UO_1320 (O_1320,N_19907,N_19500);
and UO_1321 (O_1321,N_19657,N_19276);
nor UO_1322 (O_1322,N_19929,N_19228);
and UO_1323 (O_1323,N_19665,N_19579);
and UO_1324 (O_1324,N_19350,N_19730);
or UO_1325 (O_1325,N_19509,N_19344);
and UO_1326 (O_1326,N_19228,N_19583);
or UO_1327 (O_1327,N_19927,N_19408);
nor UO_1328 (O_1328,N_19695,N_19790);
nand UO_1329 (O_1329,N_19447,N_19640);
nand UO_1330 (O_1330,N_19545,N_19390);
or UO_1331 (O_1331,N_19508,N_19662);
nand UO_1332 (O_1332,N_19802,N_19496);
or UO_1333 (O_1333,N_19332,N_19903);
or UO_1334 (O_1334,N_19649,N_19583);
or UO_1335 (O_1335,N_19768,N_19991);
and UO_1336 (O_1336,N_19439,N_19850);
nand UO_1337 (O_1337,N_19500,N_19552);
and UO_1338 (O_1338,N_19808,N_19841);
nand UO_1339 (O_1339,N_19528,N_19889);
or UO_1340 (O_1340,N_19375,N_19528);
and UO_1341 (O_1341,N_19459,N_19646);
and UO_1342 (O_1342,N_19511,N_19664);
or UO_1343 (O_1343,N_19353,N_19207);
or UO_1344 (O_1344,N_19356,N_19362);
or UO_1345 (O_1345,N_19581,N_19269);
nand UO_1346 (O_1346,N_19523,N_19370);
or UO_1347 (O_1347,N_19599,N_19871);
xor UO_1348 (O_1348,N_19937,N_19976);
nand UO_1349 (O_1349,N_19711,N_19242);
or UO_1350 (O_1350,N_19571,N_19250);
or UO_1351 (O_1351,N_19919,N_19990);
nor UO_1352 (O_1352,N_19733,N_19713);
nor UO_1353 (O_1353,N_19228,N_19562);
nor UO_1354 (O_1354,N_19730,N_19389);
nand UO_1355 (O_1355,N_19734,N_19813);
and UO_1356 (O_1356,N_19403,N_19835);
and UO_1357 (O_1357,N_19271,N_19241);
or UO_1358 (O_1358,N_19842,N_19672);
and UO_1359 (O_1359,N_19923,N_19627);
and UO_1360 (O_1360,N_19999,N_19537);
or UO_1361 (O_1361,N_19773,N_19998);
nor UO_1362 (O_1362,N_19323,N_19382);
and UO_1363 (O_1363,N_19782,N_19235);
nand UO_1364 (O_1364,N_19667,N_19467);
or UO_1365 (O_1365,N_19392,N_19650);
or UO_1366 (O_1366,N_19668,N_19932);
xor UO_1367 (O_1367,N_19737,N_19630);
and UO_1368 (O_1368,N_19575,N_19694);
or UO_1369 (O_1369,N_19787,N_19992);
nor UO_1370 (O_1370,N_19639,N_19715);
or UO_1371 (O_1371,N_19440,N_19233);
nand UO_1372 (O_1372,N_19260,N_19610);
nor UO_1373 (O_1373,N_19977,N_19211);
nand UO_1374 (O_1374,N_19396,N_19401);
nand UO_1375 (O_1375,N_19372,N_19812);
and UO_1376 (O_1376,N_19918,N_19806);
and UO_1377 (O_1377,N_19995,N_19583);
or UO_1378 (O_1378,N_19344,N_19666);
nor UO_1379 (O_1379,N_19529,N_19754);
nand UO_1380 (O_1380,N_19896,N_19927);
and UO_1381 (O_1381,N_19571,N_19626);
or UO_1382 (O_1382,N_19723,N_19466);
nand UO_1383 (O_1383,N_19725,N_19498);
or UO_1384 (O_1384,N_19445,N_19324);
nor UO_1385 (O_1385,N_19990,N_19366);
nand UO_1386 (O_1386,N_19597,N_19360);
and UO_1387 (O_1387,N_19593,N_19369);
and UO_1388 (O_1388,N_19938,N_19487);
nand UO_1389 (O_1389,N_19945,N_19834);
nor UO_1390 (O_1390,N_19880,N_19485);
or UO_1391 (O_1391,N_19977,N_19835);
or UO_1392 (O_1392,N_19221,N_19902);
nand UO_1393 (O_1393,N_19955,N_19569);
or UO_1394 (O_1394,N_19614,N_19950);
and UO_1395 (O_1395,N_19830,N_19711);
nor UO_1396 (O_1396,N_19606,N_19753);
or UO_1397 (O_1397,N_19586,N_19470);
nor UO_1398 (O_1398,N_19308,N_19947);
nor UO_1399 (O_1399,N_19726,N_19544);
nand UO_1400 (O_1400,N_19222,N_19714);
and UO_1401 (O_1401,N_19539,N_19466);
nand UO_1402 (O_1402,N_19202,N_19216);
or UO_1403 (O_1403,N_19516,N_19756);
and UO_1404 (O_1404,N_19932,N_19250);
and UO_1405 (O_1405,N_19936,N_19454);
or UO_1406 (O_1406,N_19263,N_19207);
nand UO_1407 (O_1407,N_19361,N_19911);
and UO_1408 (O_1408,N_19849,N_19371);
nand UO_1409 (O_1409,N_19260,N_19512);
and UO_1410 (O_1410,N_19505,N_19472);
or UO_1411 (O_1411,N_19230,N_19500);
and UO_1412 (O_1412,N_19672,N_19591);
nor UO_1413 (O_1413,N_19843,N_19961);
or UO_1414 (O_1414,N_19510,N_19645);
and UO_1415 (O_1415,N_19432,N_19640);
nand UO_1416 (O_1416,N_19898,N_19419);
and UO_1417 (O_1417,N_19706,N_19597);
xor UO_1418 (O_1418,N_19335,N_19951);
nor UO_1419 (O_1419,N_19811,N_19523);
or UO_1420 (O_1420,N_19695,N_19556);
or UO_1421 (O_1421,N_19790,N_19589);
nand UO_1422 (O_1422,N_19882,N_19652);
and UO_1423 (O_1423,N_19524,N_19497);
and UO_1424 (O_1424,N_19470,N_19388);
or UO_1425 (O_1425,N_19621,N_19887);
nand UO_1426 (O_1426,N_19963,N_19223);
nand UO_1427 (O_1427,N_19396,N_19329);
or UO_1428 (O_1428,N_19839,N_19632);
nand UO_1429 (O_1429,N_19290,N_19320);
and UO_1430 (O_1430,N_19234,N_19996);
and UO_1431 (O_1431,N_19865,N_19539);
or UO_1432 (O_1432,N_19537,N_19345);
and UO_1433 (O_1433,N_19701,N_19496);
and UO_1434 (O_1434,N_19842,N_19433);
and UO_1435 (O_1435,N_19270,N_19509);
and UO_1436 (O_1436,N_19757,N_19805);
and UO_1437 (O_1437,N_19977,N_19645);
nor UO_1438 (O_1438,N_19289,N_19523);
or UO_1439 (O_1439,N_19619,N_19919);
and UO_1440 (O_1440,N_19487,N_19273);
nor UO_1441 (O_1441,N_19727,N_19639);
nor UO_1442 (O_1442,N_19739,N_19488);
nor UO_1443 (O_1443,N_19784,N_19446);
nor UO_1444 (O_1444,N_19451,N_19940);
or UO_1445 (O_1445,N_19953,N_19856);
nor UO_1446 (O_1446,N_19729,N_19843);
nor UO_1447 (O_1447,N_19703,N_19511);
nand UO_1448 (O_1448,N_19477,N_19413);
nor UO_1449 (O_1449,N_19322,N_19658);
and UO_1450 (O_1450,N_19564,N_19229);
nor UO_1451 (O_1451,N_19570,N_19248);
nor UO_1452 (O_1452,N_19293,N_19676);
nor UO_1453 (O_1453,N_19274,N_19559);
or UO_1454 (O_1454,N_19341,N_19720);
and UO_1455 (O_1455,N_19829,N_19994);
nand UO_1456 (O_1456,N_19369,N_19271);
nor UO_1457 (O_1457,N_19743,N_19856);
nor UO_1458 (O_1458,N_19961,N_19225);
nor UO_1459 (O_1459,N_19491,N_19759);
nand UO_1460 (O_1460,N_19529,N_19500);
or UO_1461 (O_1461,N_19365,N_19450);
or UO_1462 (O_1462,N_19577,N_19618);
nor UO_1463 (O_1463,N_19786,N_19346);
nor UO_1464 (O_1464,N_19926,N_19689);
and UO_1465 (O_1465,N_19997,N_19763);
and UO_1466 (O_1466,N_19543,N_19471);
or UO_1467 (O_1467,N_19483,N_19721);
or UO_1468 (O_1468,N_19902,N_19350);
or UO_1469 (O_1469,N_19305,N_19680);
or UO_1470 (O_1470,N_19487,N_19608);
or UO_1471 (O_1471,N_19636,N_19551);
nand UO_1472 (O_1472,N_19326,N_19646);
nor UO_1473 (O_1473,N_19479,N_19539);
nor UO_1474 (O_1474,N_19805,N_19589);
nand UO_1475 (O_1475,N_19378,N_19888);
and UO_1476 (O_1476,N_19543,N_19862);
nand UO_1477 (O_1477,N_19242,N_19541);
and UO_1478 (O_1478,N_19974,N_19888);
nor UO_1479 (O_1479,N_19918,N_19490);
nand UO_1480 (O_1480,N_19527,N_19470);
nor UO_1481 (O_1481,N_19358,N_19536);
and UO_1482 (O_1482,N_19305,N_19335);
nand UO_1483 (O_1483,N_19746,N_19453);
nor UO_1484 (O_1484,N_19562,N_19333);
nand UO_1485 (O_1485,N_19764,N_19799);
and UO_1486 (O_1486,N_19317,N_19254);
and UO_1487 (O_1487,N_19704,N_19991);
or UO_1488 (O_1488,N_19706,N_19517);
nand UO_1489 (O_1489,N_19478,N_19651);
nand UO_1490 (O_1490,N_19607,N_19446);
or UO_1491 (O_1491,N_19938,N_19577);
nor UO_1492 (O_1492,N_19570,N_19866);
and UO_1493 (O_1493,N_19328,N_19348);
or UO_1494 (O_1494,N_19635,N_19809);
or UO_1495 (O_1495,N_19931,N_19497);
or UO_1496 (O_1496,N_19766,N_19390);
and UO_1497 (O_1497,N_19752,N_19726);
or UO_1498 (O_1498,N_19236,N_19814);
nand UO_1499 (O_1499,N_19744,N_19805);
and UO_1500 (O_1500,N_19839,N_19276);
and UO_1501 (O_1501,N_19824,N_19839);
and UO_1502 (O_1502,N_19372,N_19642);
and UO_1503 (O_1503,N_19323,N_19412);
nor UO_1504 (O_1504,N_19206,N_19262);
and UO_1505 (O_1505,N_19303,N_19930);
or UO_1506 (O_1506,N_19385,N_19440);
or UO_1507 (O_1507,N_19378,N_19209);
or UO_1508 (O_1508,N_19291,N_19958);
and UO_1509 (O_1509,N_19945,N_19647);
nor UO_1510 (O_1510,N_19235,N_19219);
and UO_1511 (O_1511,N_19549,N_19435);
or UO_1512 (O_1512,N_19778,N_19334);
or UO_1513 (O_1513,N_19381,N_19725);
or UO_1514 (O_1514,N_19947,N_19524);
and UO_1515 (O_1515,N_19502,N_19881);
nor UO_1516 (O_1516,N_19291,N_19302);
nand UO_1517 (O_1517,N_19774,N_19878);
and UO_1518 (O_1518,N_19387,N_19337);
nor UO_1519 (O_1519,N_19996,N_19545);
nand UO_1520 (O_1520,N_19591,N_19378);
nand UO_1521 (O_1521,N_19250,N_19712);
nand UO_1522 (O_1522,N_19857,N_19812);
and UO_1523 (O_1523,N_19401,N_19941);
nor UO_1524 (O_1524,N_19833,N_19496);
or UO_1525 (O_1525,N_19795,N_19576);
nor UO_1526 (O_1526,N_19858,N_19961);
and UO_1527 (O_1527,N_19489,N_19962);
and UO_1528 (O_1528,N_19894,N_19213);
nand UO_1529 (O_1529,N_19676,N_19413);
nor UO_1530 (O_1530,N_19818,N_19895);
nor UO_1531 (O_1531,N_19830,N_19854);
nand UO_1532 (O_1532,N_19911,N_19204);
or UO_1533 (O_1533,N_19586,N_19756);
nor UO_1534 (O_1534,N_19332,N_19920);
nor UO_1535 (O_1535,N_19574,N_19572);
nand UO_1536 (O_1536,N_19265,N_19262);
and UO_1537 (O_1537,N_19716,N_19971);
nand UO_1538 (O_1538,N_19230,N_19714);
nor UO_1539 (O_1539,N_19403,N_19642);
nand UO_1540 (O_1540,N_19781,N_19895);
nand UO_1541 (O_1541,N_19500,N_19603);
nand UO_1542 (O_1542,N_19749,N_19932);
nor UO_1543 (O_1543,N_19606,N_19771);
and UO_1544 (O_1544,N_19261,N_19386);
or UO_1545 (O_1545,N_19360,N_19247);
nor UO_1546 (O_1546,N_19503,N_19927);
nor UO_1547 (O_1547,N_19717,N_19811);
nand UO_1548 (O_1548,N_19677,N_19614);
nor UO_1549 (O_1549,N_19393,N_19642);
nand UO_1550 (O_1550,N_19752,N_19380);
nand UO_1551 (O_1551,N_19943,N_19309);
or UO_1552 (O_1552,N_19659,N_19472);
and UO_1553 (O_1553,N_19697,N_19404);
or UO_1554 (O_1554,N_19989,N_19230);
or UO_1555 (O_1555,N_19762,N_19258);
nor UO_1556 (O_1556,N_19534,N_19506);
or UO_1557 (O_1557,N_19837,N_19371);
nand UO_1558 (O_1558,N_19839,N_19206);
nor UO_1559 (O_1559,N_19522,N_19739);
or UO_1560 (O_1560,N_19336,N_19549);
nor UO_1561 (O_1561,N_19793,N_19659);
nor UO_1562 (O_1562,N_19931,N_19594);
or UO_1563 (O_1563,N_19421,N_19402);
and UO_1564 (O_1564,N_19591,N_19274);
or UO_1565 (O_1565,N_19676,N_19958);
nor UO_1566 (O_1566,N_19270,N_19502);
nand UO_1567 (O_1567,N_19877,N_19452);
nand UO_1568 (O_1568,N_19973,N_19533);
or UO_1569 (O_1569,N_19288,N_19961);
or UO_1570 (O_1570,N_19998,N_19905);
or UO_1571 (O_1571,N_19831,N_19501);
or UO_1572 (O_1572,N_19932,N_19576);
nor UO_1573 (O_1573,N_19764,N_19631);
and UO_1574 (O_1574,N_19972,N_19647);
nand UO_1575 (O_1575,N_19633,N_19966);
nand UO_1576 (O_1576,N_19355,N_19715);
and UO_1577 (O_1577,N_19212,N_19388);
nor UO_1578 (O_1578,N_19502,N_19643);
nand UO_1579 (O_1579,N_19719,N_19977);
or UO_1580 (O_1580,N_19560,N_19340);
and UO_1581 (O_1581,N_19753,N_19839);
or UO_1582 (O_1582,N_19557,N_19681);
nor UO_1583 (O_1583,N_19692,N_19480);
or UO_1584 (O_1584,N_19932,N_19457);
and UO_1585 (O_1585,N_19612,N_19291);
nor UO_1586 (O_1586,N_19976,N_19972);
xnor UO_1587 (O_1587,N_19446,N_19573);
nor UO_1588 (O_1588,N_19377,N_19354);
and UO_1589 (O_1589,N_19887,N_19345);
or UO_1590 (O_1590,N_19672,N_19987);
nand UO_1591 (O_1591,N_19736,N_19597);
nor UO_1592 (O_1592,N_19297,N_19843);
and UO_1593 (O_1593,N_19495,N_19801);
or UO_1594 (O_1594,N_19301,N_19893);
nand UO_1595 (O_1595,N_19820,N_19850);
or UO_1596 (O_1596,N_19601,N_19850);
nand UO_1597 (O_1597,N_19243,N_19621);
or UO_1598 (O_1598,N_19888,N_19295);
or UO_1599 (O_1599,N_19781,N_19391);
and UO_1600 (O_1600,N_19308,N_19303);
xor UO_1601 (O_1601,N_19778,N_19395);
or UO_1602 (O_1602,N_19797,N_19503);
or UO_1603 (O_1603,N_19943,N_19524);
or UO_1604 (O_1604,N_19842,N_19755);
and UO_1605 (O_1605,N_19205,N_19937);
nor UO_1606 (O_1606,N_19928,N_19982);
and UO_1607 (O_1607,N_19262,N_19700);
nand UO_1608 (O_1608,N_19498,N_19915);
nor UO_1609 (O_1609,N_19403,N_19892);
or UO_1610 (O_1610,N_19549,N_19651);
or UO_1611 (O_1611,N_19556,N_19287);
or UO_1612 (O_1612,N_19440,N_19333);
nor UO_1613 (O_1613,N_19923,N_19939);
nand UO_1614 (O_1614,N_19508,N_19877);
nand UO_1615 (O_1615,N_19217,N_19467);
nor UO_1616 (O_1616,N_19375,N_19409);
nor UO_1617 (O_1617,N_19501,N_19711);
nor UO_1618 (O_1618,N_19247,N_19547);
or UO_1619 (O_1619,N_19922,N_19630);
nand UO_1620 (O_1620,N_19384,N_19497);
nor UO_1621 (O_1621,N_19253,N_19593);
nand UO_1622 (O_1622,N_19760,N_19668);
or UO_1623 (O_1623,N_19290,N_19363);
nand UO_1624 (O_1624,N_19506,N_19641);
or UO_1625 (O_1625,N_19343,N_19911);
nor UO_1626 (O_1626,N_19629,N_19521);
or UO_1627 (O_1627,N_19668,N_19735);
nand UO_1628 (O_1628,N_19395,N_19435);
or UO_1629 (O_1629,N_19706,N_19485);
and UO_1630 (O_1630,N_19701,N_19545);
nand UO_1631 (O_1631,N_19353,N_19735);
or UO_1632 (O_1632,N_19967,N_19802);
nor UO_1633 (O_1633,N_19972,N_19918);
and UO_1634 (O_1634,N_19991,N_19349);
and UO_1635 (O_1635,N_19702,N_19765);
xor UO_1636 (O_1636,N_19433,N_19607);
nand UO_1637 (O_1637,N_19955,N_19503);
and UO_1638 (O_1638,N_19357,N_19624);
or UO_1639 (O_1639,N_19371,N_19780);
or UO_1640 (O_1640,N_19711,N_19686);
or UO_1641 (O_1641,N_19491,N_19405);
and UO_1642 (O_1642,N_19957,N_19483);
or UO_1643 (O_1643,N_19332,N_19626);
nor UO_1644 (O_1644,N_19260,N_19462);
nor UO_1645 (O_1645,N_19478,N_19552);
nand UO_1646 (O_1646,N_19823,N_19216);
or UO_1647 (O_1647,N_19755,N_19987);
nand UO_1648 (O_1648,N_19400,N_19209);
nand UO_1649 (O_1649,N_19663,N_19775);
and UO_1650 (O_1650,N_19752,N_19295);
or UO_1651 (O_1651,N_19549,N_19694);
or UO_1652 (O_1652,N_19924,N_19585);
nor UO_1653 (O_1653,N_19848,N_19652);
nor UO_1654 (O_1654,N_19674,N_19644);
or UO_1655 (O_1655,N_19894,N_19968);
nand UO_1656 (O_1656,N_19636,N_19936);
and UO_1657 (O_1657,N_19340,N_19493);
nor UO_1658 (O_1658,N_19895,N_19269);
nand UO_1659 (O_1659,N_19667,N_19681);
nand UO_1660 (O_1660,N_19969,N_19856);
nand UO_1661 (O_1661,N_19792,N_19587);
or UO_1662 (O_1662,N_19332,N_19263);
nor UO_1663 (O_1663,N_19654,N_19253);
nor UO_1664 (O_1664,N_19504,N_19667);
and UO_1665 (O_1665,N_19367,N_19286);
and UO_1666 (O_1666,N_19486,N_19781);
and UO_1667 (O_1667,N_19321,N_19714);
and UO_1668 (O_1668,N_19600,N_19819);
nor UO_1669 (O_1669,N_19307,N_19842);
and UO_1670 (O_1670,N_19542,N_19971);
nor UO_1671 (O_1671,N_19960,N_19307);
or UO_1672 (O_1672,N_19734,N_19808);
and UO_1673 (O_1673,N_19998,N_19921);
or UO_1674 (O_1674,N_19638,N_19306);
and UO_1675 (O_1675,N_19267,N_19739);
nand UO_1676 (O_1676,N_19459,N_19781);
or UO_1677 (O_1677,N_19980,N_19586);
or UO_1678 (O_1678,N_19581,N_19869);
nor UO_1679 (O_1679,N_19728,N_19296);
nor UO_1680 (O_1680,N_19917,N_19696);
or UO_1681 (O_1681,N_19894,N_19273);
or UO_1682 (O_1682,N_19881,N_19906);
or UO_1683 (O_1683,N_19404,N_19869);
nor UO_1684 (O_1684,N_19218,N_19979);
nand UO_1685 (O_1685,N_19502,N_19792);
and UO_1686 (O_1686,N_19490,N_19340);
and UO_1687 (O_1687,N_19264,N_19855);
or UO_1688 (O_1688,N_19677,N_19330);
and UO_1689 (O_1689,N_19658,N_19254);
nor UO_1690 (O_1690,N_19631,N_19882);
nand UO_1691 (O_1691,N_19580,N_19850);
xor UO_1692 (O_1692,N_19777,N_19544);
nand UO_1693 (O_1693,N_19958,N_19410);
nand UO_1694 (O_1694,N_19536,N_19387);
nor UO_1695 (O_1695,N_19292,N_19496);
nand UO_1696 (O_1696,N_19753,N_19977);
and UO_1697 (O_1697,N_19981,N_19270);
and UO_1698 (O_1698,N_19532,N_19851);
nand UO_1699 (O_1699,N_19624,N_19977);
or UO_1700 (O_1700,N_19932,N_19601);
nand UO_1701 (O_1701,N_19391,N_19643);
nor UO_1702 (O_1702,N_19822,N_19281);
nor UO_1703 (O_1703,N_19512,N_19996);
and UO_1704 (O_1704,N_19230,N_19685);
or UO_1705 (O_1705,N_19495,N_19697);
and UO_1706 (O_1706,N_19202,N_19709);
or UO_1707 (O_1707,N_19775,N_19414);
nor UO_1708 (O_1708,N_19275,N_19814);
or UO_1709 (O_1709,N_19890,N_19893);
and UO_1710 (O_1710,N_19530,N_19721);
and UO_1711 (O_1711,N_19218,N_19861);
or UO_1712 (O_1712,N_19277,N_19835);
nand UO_1713 (O_1713,N_19430,N_19332);
or UO_1714 (O_1714,N_19980,N_19816);
nor UO_1715 (O_1715,N_19486,N_19947);
nor UO_1716 (O_1716,N_19775,N_19474);
nand UO_1717 (O_1717,N_19611,N_19206);
nor UO_1718 (O_1718,N_19303,N_19821);
nand UO_1719 (O_1719,N_19718,N_19270);
nor UO_1720 (O_1720,N_19423,N_19880);
nor UO_1721 (O_1721,N_19383,N_19326);
nand UO_1722 (O_1722,N_19976,N_19382);
nor UO_1723 (O_1723,N_19890,N_19529);
and UO_1724 (O_1724,N_19500,N_19583);
nor UO_1725 (O_1725,N_19316,N_19569);
nand UO_1726 (O_1726,N_19276,N_19993);
nor UO_1727 (O_1727,N_19354,N_19342);
nand UO_1728 (O_1728,N_19512,N_19435);
nand UO_1729 (O_1729,N_19318,N_19640);
nand UO_1730 (O_1730,N_19239,N_19203);
and UO_1731 (O_1731,N_19266,N_19699);
nor UO_1732 (O_1732,N_19983,N_19713);
nand UO_1733 (O_1733,N_19928,N_19960);
or UO_1734 (O_1734,N_19826,N_19620);
nand UO_1735 (O_1735,N_19664,N_19725);
or UO_1736 (O_1736,N_19364,N_19982);
nand UO_1737 (O_1737,N_19840,N_19564);
nor UO_1738 (O_1738,N_19687,N_19365);
nor UO_1739 (O_1739,N_19667,N_19353);
or UO_1740 (O_1740,N_19470,N_19696);
and UO_1741 (O_1741,N_19653,N_19457);
or UO_1742 (O_1742,N_19445,N_19270);
and UO_1743 (O_1743,N_19406,N_19899);
nand UO_1744 (O_1744,N_19609,N_19954);
nand UO_1745 (O_1745,N_19988,N_19613);
nor UO_1746 (O_1746,N_19439,N_19573);
nand UO_1747 (O_1747,N_19430,N_19716);
and UO_1748 (O_1748,N_19248,N_19718);
nor UO_1749 (O_1749,N_19628,N_19678);
or UO_1750 (O_1750,N_19937,N_19523);
nor UO_1751 (O_1751,N_19624,N_19407);
or UO_1752 (O_1752,N_19221,N_19541);
nand UO_1753 (O_1753,N_19309,N_19358);
and UO_1754 (O_1754,N_19437,N_19398);
or UO_1755 (O_1755,N_19766,N_19842);
nor UO_1756 (O_1756,N_19471,N_19909);
nor UO_1757 (O_1757,N_19274,N_19348);
nand UO_1758 (O_1758,N_19676,N_19430);
and UO_1759 (O_1759,N_19506,N_19502);
nor UO_1760 (O_1760,N_19424,N_19966);
and UO_1761 (O_1761,N_19892,N_19621);
nand UO_1762 (O_1762,N_19669,N_19919);
and UO_1763 (O_1763,N_19408,N_19700);
or UO_1764 (O_1764,N_19573,N_19587);
nand UO_1765 (O_1765,N_19258,N_19667);
nand UO_1766 (O_1766,N_19424,N_19772);
nand UO_1767 (O_1767,N_19315,N_19831);
and UO_1768 (O_1768,N_19506,N_19877);
and UO_1769 (O_1769,N_19697,N_19409);
nor UO_1770 (O_1770,N_19442,N_19551);
or UO_1771 (O_1771,N_19995,N_19940);
or UO_1772 (O_1772,N_19242,N_19588);
nor UO_1773 (O_1773,N_19448,N_19285);
nand UO_1774 (O_1774,N_19633,N_19449);
and UO_1775 (O_1775,N_19357,N_19950);
or UO_1776 (O_1776,N_19704,N_19603);
nor UO_1777 (O_1777,N_19306,N_19791);
and UO_1778 (O_1778,N_19466,N_19357);
or UO_1779 (O_1779,N_19320,N_19982);
xor UO_1780 (O_1780,N_19798,N_19492);
nand UO_1781 (O_1781,N_19369,N_19245);
or UO_1782 (O_1782,N_19760,N_19627);
and UO_1783 (O_1783,N_19390,N_19838);
nand UO_1784 (O_1784,N_19563,N_19364);
or UO_1785 (O_1785,N_19506,N_19997);
or UO_1786 (O_1786,N_19972,N_19316);
nor UO_1787 (O_1787,N_19985,N_19979);
nor UO_1788 (O_1788,N_19748,N_19488);
or UO_1789 (O_1789,N_19717,N_19382);
nand UO_1790 (O_1790,N_19372,N_19559);
nor UO_1791 (O_1791,N_19842,N_19905);
nand UO_1792 (O_1792,N_19509,N_19497);
and UO_1793 (O_1793,N_19909,N_19211);
nand UO_1794 (O_1794,N_19507,N_19431);
and UO_1795 (O_1795,N_19234,N_19445);
and UO_1796 (O_1796,N_19499,N_19362);
and UO_1797 (O_1797,N_19514,N_19934);
nand UO_1798 (O_1798,N_19923,N_19833);
or UO_1799 (O_1799,N_19625,N_19287);
nor UO_1800 (O_1800,N_19975,N_19429);
or UO_1801 (O_1801,N_19746,N_19559);
nor UO_1802 (O_1802,N_19433,N_19367);
nand UO_1803 (O_1803,N_19682,N_19235);
nand UO_1804 (O_1804,N_19256,N_19246);
nand UO_1805 (O_1805,N_19453,N_19255);
or UO_1806 (O_1806,N_19244,N_19242);
and UO_1807 (O_1807,N_19466,N_19816);
nand UO_1808 (O_1808,N_19713,N_19398);
or UO_1809 (O_1809,N_19406,N_19751);
and UO_1810 (O_1810,N_19378,N_19841);
or UO_1811 (O_1811,N_19919,N_19849);
nor UO_1812 (O_1812,N_19967,N_19249);
nand UO_1813 (O_1813,N_19403,N_19970);
and UO_1814 (O_1814,N_19919,N_19428);
nand UO_1815 (O_1815,N_19554,N_19273);
nand UO_1816 (O_1816,N_19660,N_19206);
nand UO_1817 (O_1817,N_19915,N_19711);
nor UO_1818 (O_1818,N_19438,N_19317);
and UO_1819 (O_1819,N_19818,N_19808);
nand UO_1820 (O_1820,N_19353,N_19610);
and UO_1821 (O_1821,N_19478,N_19700);
or UO_1822 (O_1822,N_19260,N_19698);
nand UO_1823 (O_1823,N_19811,N_19361);
nor UO_1824 (O_1824,N_19960,N_19402);
and UO_1825 (O_1825,N_19355,N_19948);
nand UO_1826 (O_1826,N_19397,N_19561);
or UO_1827 (O_1827,N_19205,N_19485);
nor UO_1828 (O_1828,N_19441,N_19558);
or UO_1829 (O_1829,N_19594,N_19378);
and UO_1830 (O_1830,N_19917,N_19545);
nand UO_1831 (O_1831,N_19745,N_19478);
nor UO_1832 (O_1832,N_19721,N_19991);
or UO_1833 (O_1833,N_19702,N_19363);
nor UO_1834 (O_1834,N_19317,N_19623);
or UO_1835 (O_1835,N_19817,N_19341);
nand UO_1836 (O_1836,N_19399,N_19207);
xor UO_1837 (O_1837,N_19625,N_19285);
nand UO_1838 (O_1838,N_19755,N_19531);
or UO_1839 (O_1839,N_19882,N_19341);
nor UO_1840 (O_1840,N_19631,N_19475);
nand UO_1841 (O_1841,N_19637,N_19516);
nand UO_1842 (O_1842,N_19881,N_19392);
nor UO_1843 (O_1843,N_19509,N_19221);
and UO_1844 (O_1844,N_19899,N_19245);
and UO_1845 (O_1845,N_19472,N_19531);
or UO_1846 (O_1846,N_19965,N_19386);
or UO_1847 (O_1847,N_19472,N_19230);
and UO_1848 (O_1848,N_19478,N_19299);
and UO_1849 (O_1849,N_19804,N_19700);
nand UO_1850 (O_1850,N_19526,N_19943);
or UO_1851 (O_1851,N_19358,N_19885);
and UO_1852 (O_1852,N_19320,N_19654);
and UO_1853 (O_1853,N_19976,N_19497);
nand UO_1854 (O_1854,N_19708,N_19302);
or UO_1855 (O_1855,N_19816,N_19727);
nand UO_1856 (O_1856,N_19599,N_19695);
and UO_1857 (O_1857,N_19418,N_19497);
and UO_1858 (O_1858,N_19493,N_19265);
or UO_1859 (O_1859,N_19873,N_19552);
nor UO_1860 (O_1860,N_19564,N_19727);
and UO_1861 (O_1861,N_19548,N_19619);
nand UO_1862 (O_1862,N_19721,N_19288);
nor UO_1863 (O_1863,N_19327,N_19461);
nand UO_1864 (O_1864,N_19886,N_19538);
and UO_1865 (O_1865,N_19259,N_19977);
nor UO_1866 (O_1866,N_19336,N_19397);
and UO_1867 (O_1867,N_19234,N_19314);
nand UO_1868 (O_1868,N_19905,N_19505);
nor UO_1869 (O_1869,N_19874,N_19975);
nand UO_1870 (O_1870,N_19305,N_19586);
nor UO_1871 (O_1871,N_19994,N_19406);
nor UO_1872 (O_1872,N_19520,N_19580);
and UO_1873 (O_1873,N_19916,N_19553);
and UO_1874 (O_1874,N_19662,N_19972);
nand UO_1875 (O_1875,N_19298,N_19661);
nor UO_1876 (O_1876,N_19218,N_19995);
or UO_1877 (O_1877,N_19346,N_19302);
nand UO_1878 (O_1878,N_19392,N_19291);
nor UO_1879 (O_1879,N_19938,N_19229);
and UO_1880 (O_1880,N_19845,N_19512);
and UO_1881 (O_1881,N_19659,N_19706);
or UO_1882 (O_1882,N_19551,N_19657);
nand UO_1883 (O_1883,N_19429,N_19408);
nor UO_1884 (O_1884,N_19487,N_19832);
or UO_1885 (O_1885,N_19948,N_19256);
and UO_1886 (O_1886,N_19482,N_19255);
or UO_1887 (O_1887,N_19998,N_19203);
and UO_1888 (O_1888,N_19673,N_19494);
nor UO_1889 (O_1889,N_19701,N_19849);
nor UO_1890 (O_1890,N_19538,N_19609);
nor UO_1891 (O_1891,N_19323,N_19474);
and UO_1892 (O_1892,N_19256,N_19823);
or UO_1893 (O_1893,N_19215,N_19991);
nand UO_1894 (O_1894,N_19857,N_19269);
nand UO_1895 (O_1895,N_19540,N_19327);
and UO_1896 (O_1896,N_19339,N_19690);
nand UO_1897 (O_1897,N_19719,N_19994);
nand UO_1898 (O_1898,N_19472,N_19254);
nand UO_1899 (O_1899,N_19989,N_19779);
nand UO_1900 (O_1900,N_19723,N_19816);
nand UO_1901 (O_1901,N_19354,N_19965);
or UO_1902 (O_1902,N_19964,N_19577);
nand UO_1903 (O_1903,N_19983,N_19507);
and UO_1904 (O_1904,N_19769,N_19834);
nand UO_1905 (O_1905,N_19747,N_19263);
nand UO_1906 (O_1906,N_19709,N_19365);
or UO_1907 (O_1907,N_19348,N_19286);
and UO_1908 (O_1908,N_19402,N_19394);
or UO_1909 (O_1909,N_19427,N_19756);
nor UO_1910 (O_1910,N_19717,N_19742);
nor UO_1911 (O_1911,N_19920,N_19468);
or UO_1912 (O_1912,N_19820,N_19383);
and UO_1913 (O_1913,N_19297,N_19816);
nor UO_1914 (O_1914,N_19938,N_19367);
and UO_1915 (O_1915,N_19362,N_19841);
nand UO_1916 (O_1916,N_19505,N_19670);
or UO_1917 (O_1917,N_19932,N_19533);
nor UO_1918 (O_1918,N_19343,N_19556);
nor UO_1919 (O_1919,N_19856,N_19235);
nand UO_1920 (O_1920,N_19589,N_19324);
and UO_1921 (O_1921,N_19751,N_19272);
nor UO_1922 (O_1922,N_19411,N_19374);
or UO_1923 (O_1923,N_19350,N_19835);
and UO_1924 (O_1924,N_19264,N_19530);
nor UO_1925 (O_1925,N_19547,N_19205);
or UO_1926 (O_1926,N_19964,N_19366);
and UO_1927 (O_1927,N_19898,N_19593);
nor UO_1928 (O_1928,N_19642,N_19588);
nand UO_1929 (O_1929,N_19403,N_19383);
or UO_1930 (O_1930,N_19668,N_19279);
and UO_1931 (O_1931,N_19724,N_19907);
and UO_1932 (O_1932,N_19410,N_19684);
or UO_1933 (O_1933,N_19620,N_19236);
nor UO_1934 (O_1934,N_19367,N_19373);
nand UO_1935 (O_1935,N_19484,N_19267);
or UO_1936 (O_1936,N_19348,N_19624);
nor UO_1937 (O_1937,N_19328,N_19807);
nand UO_1938 (O_1938,N_19514,N_19721);
nor UO_1939 (O_1939,N_19365,N_19310);
nor UO_1940 (O_1940,N_19782,N_19742);
nand UO_1941 (O_1941,N_19279,N_19786);
xor UO_1942 (O_1942,N_19802,N_19509);
or UO_1943 (O_1943,N_19625,N_19806);
nand UO_1944 (O_1944,N_19780,N_19370);
nand UO_1945 (O_1945,N_19272,N_19894);
nand UO_1946 (O_1946,N_19312,N_19638);
or UO_1947 (O_1947,N_19792,N_19791);
or UO_1948 (O_1948,N_19858,N_19915);
nor UO_1949 (O_1949,N_19838,N_19873);
or UO_1950 (O_1950,N_19492,N_19869);
or UO_1951 (O_1951,N_19814,N_19752);
and UO_1952 (O_1952,N_19800,N_19768);
and UO_1953 (O_1953,N_19739,N_19529);
or UO_1954 (O_1954,N_19771,N_19356);
and UO_1955 (O_1955,N_19363,N_19223);
and UO_1956 (O_1956,N_19840,N_19753);
nor UO_1957 (O_1957,N_19616,N_19852);
nand UO_1958 (O_1958,N_19724,N_19799);
nor UO_1959 (O_1959,N_19227,N_19481);
or UO_1960 (O_1960,N_19404,N_19298);
or UO_1961 (O_1961,N_19726,N_19461);
nand UO_1962 (O_1962,N_19243,N_19293);
nand UO_1963 (O_1963,N_19373,N_19660);
nor UO_1964 (O_1964,N_19650,N_19688);
nand UO_1965 (O_1965,N_19937,N_19798);
nor UO_1966 (O_1966,N_19782,N_19242);
nand UO_1967 (O_1967,N_19803,N_19799);
nand UO_1968 (O_1968,N_19238,N_19757);
nor UO_1969 (O_1969,N_19873,N_19537);
or UO_1970 (O_1970,N_19836,N_19250);
nand UO_1971 (O_1971,N_19956,N_19468);
nand UO_1972 (O_1972,N_19424,N_19901);
and UO_1973 (O_1973,N_19569,N_19394);
and UO_1974 (O_1974,N_19266,N_19779);
nand UO_1975 (O_1975,N_19977,N_19218);
nand UO_1976 (O_1976,N_19871,N_19925);
or UO_1977 (O_1977,N_19892,N_19796);
or UO_1978 (O_1978,N_19581,N_19693);
nor UO_1979 (O_1979,N_19944,N_19257);
or UO_1980 (O_1980,N_19515,N_19252);
or UO_1981 (O_1981,N_19322,N_19350);
and UO_1982 (O_1982,N_19336,N_19843);
or UO_1983 (O_1983,N_19963,N_19705);
nor UO_1984 (O_1984,N_19639,N_19923);
nor UO_1985 (O_1985,N_19319,N_19677);
nor UO_1986 (O_1986,N_19431,N_19204);
or UO_1987 (O_1987,N_19469,N_19488);
nand UO_1988 (O_1988,N_19932,N_19361);
nand UO_1989 (O_1989,N_19774,N_19213);
nor UO_1990 (O_1990,N_19808,N_19232);
nand UO_1991 (O_1991,N_19468,N_19990);
nand UO_1992 (O_1992,N_19309,N_19737);
or UO_1993 (O_1993,N_19971,N_19522);
nor UO_1994 (O_1994,N_19218,N_19469);
nor UO_1995 (O_1995,N_19685,N_19207);
or UO_1996 (O_1996,N_19834,N_19962);
and UO_1997 (O_1997,N_19210,N_19590);
or UO_1998 (O_1998,N_19479,N_19422);
nand UO_1999 (O_1999,N_19696,N_19325);
nand UO_2000 (O_2000,N_19894,N_19297);
nor UO_2001 (O_2001,N_19654,N_19596);
nand UO_2002 (O_2002,N_19735,N_19549);
or UO_2003 (O_2003,N_19825,N_19576);
and UO_2004 (O_2004,N_19452,N_19692);
xnor UO_2005 (O_2005,N_19970,N_19237);
and UO_2006 (O_2006,N_19717,N_19507);
or UO_2007 (O_2007,N_19348,N_19784);
or UO_2008 (O_2008,N_19759,N_19603);
or UO_2009 (O_2009,N_19666,N_19852);
and UO_2010 (O_2010,N_19889,N_19735);
and UO_2011 (O_2011,N_19201,N_19589);
or UO_2012 (O_2012,N_19262,N_19930);
or UO_2013 (O_2013,N_19994,N_19350);
or UO_2014 (O_2014,N_19683,N_19917);
and UO_2015 (O_2015,N_19552,N_19784);
and UO_2016 (O_2016,N_19774,N_19890);
and UO_2017 (O_2017,N_19895,N_19245);
or UO_2018 (O_2018,N_19457,N_19472);
nor UO_2019 (O_2019,N_19790,N_19933);
or UO_2020 (O_2020,N_19506,N_19267);
or UO_2021 (O_2021,N_19297,N_19931);
nor UO_2022 (O_2022,N_19589,N_19926);
nand UO_2023 (O_2023,N_19724,N_19564);
and UO_2024 (O_2024,N_19389,N_19285);
and UO_2025 (O_2025,N_19400,N_19532);
nor UO_2026 (O_2026,N_19593,N_19772);
or UO_2027 (O_2027,N_19581,N_19552);
nor UO_2028 (O_2028,N_19825,N_19780);
or UO_2029 (O_2029,N_19451,N_19217);
or UO_2030 (O_2030,N_19923,N_19765);
and UO_2031 (O_2031,N_19722,N_19959);
and UO_2032 (O_2032,N_19623,N_19274);
nand UO_2033 (O_2033,N_19782,N_19847);
or UO_2034 (O_2034,N_19892,N_19597);
nand UO_2035 (O_2035,N_19244,N_19502);
or UO_2036 (O_2036,N_19898,N_19465);
xnor UO_2037 (O_2037,N_19815,N_19539);
nand UO_2038 (O_2038,N_19718,N_19813);
or UO_2039 (O_2039,N_19909,N_19369);
and UO_2040 (O_2040,N_19586,N_19657);
or UO_2041 (O_2041,N_19593,N_19385);
or UO_2042 (O_2042,N_19930,N_19217);
nor UO_2043 (O_2043,N_19480,N_19803);
or UO_2044 (O_2044,N_19537,N_19815);
nand UO_2045 (O_2045,N_19888,N_19703);
and UO_2046 (O_2046,N_19901,N_19262);
nor UO_2047 (O_2047,N_19359,N_19264);
or UO_2048 (O_2048,N_19289,N_19871);
nor UO_2049 (O_2049,N_19476,N_19543);
nor UO_2050 (O_2050,N_19730,N_19292);
nand UO_2051 (O_2051,N_19531,N_19752);
and UO_2052 (O_2052,N_19871,N_19923);
nor UO_2053 (O_2053,N_19925,N_19748);
nor UO_2054 (O_2054,N_19712,N_19692);
nor UO_2055 (O_2055,N_19329,N_19640);
or UO_2056 (O_2056,N_19410,N_19507);
nor UO_2057 (O_2057,N_19619,N_19433);
or UO_2058 (O_2058,N_19616,N_19637);
nor UO_2059 (O_2059,N_19479,N_19834);
nor UO_2060 (O_2060,N_19227,N_19578);
and UO_2061 (O_2061,N_19820,N_19629);
nand UO_2062 (O_2062,N_19350,N_19554);
and UO_2063 (O_2063,N_19435,N_19642);
and UO_2064 (O_2064,N_19506,N_19358);
or UO_2065 (O_2065,N_19246,N_19225);
or UO_2066 (O_2066,N_19807,N_19453);
xnor UO_2067 (O_2067,N_19571,N_19748);
and UO_2068 (O_2068,N_19690,N_19868);
nand UO_2069 (O_2069,N_19204,N_19569);
and UO_2070 (O_2070,N_19466,N_19669);
nand UO_2071 (O_2071,N_19791,N_19689);
and UO_2072 (O_2072,N_19927,N_19236);
or UO_2073 (O_2073,N_19689,N_19258);
nand UO_2074 (O_2074,N_19657,N_19699);
nor UO_2075 (O_2075,N_19901,N_19563);
nand UO_2076 (O_2076,N_19456,N_19922);
nand UO_2077 (O_2077,N_19828,N_19393);
and UO_2078 (O_2078,N_19849,N_19768);
or UO_2079 (O_2079,N_19565,N_19274);
or UO_2080 (O_2080,N_19218,N_19869);
or UO_2081 (O_2081,N_19508,N_19804);
nor UO_2082 (O_2082,N_19480,N_19937);
nand UO_2083 (O_2083,N_19827,N_19271);
nand UO_2084 (O_2084,N_19339,N_19471);
or UO_2085 (O_2085,N_19337,N_19795);
nand UO_2086 (O_2086,N_19660,N_19274);
and UO_2087 (O_2087,N_19902,N_19871);
or UO_2088 (O_2088,N_19523,N_19420);
or UO_2089 (O_2089,N_19294,N_19463);
and UO_2090 (O_2090,N_19571,N_19342);
or UO_2091 (O_2091,N_19786,N_19626);
and UO_2092 (O_2092,N_19365,N_19506);
or UO_2093 (O_2093,N_19410,N_19459);
nand UO_2094 (O_2094,N_19722,N_19622);
and UO_2095 (O_2095,N_19780,N_19451);
xor UO_2096 (O_2096,N_19655,N_19793);
nor UO_2097 (O_2097,N_19297,N_19542);
and UO_2098 (O_2098,N_19949,N_19367);
nor UO_2099 (O_2099,N_19905,N_19688);
and UO_2100 (O_2100,N_19889,N_19933);
nand UO_2101 (O_2101,N_19623,N_19782);
or UO_2102 (O_2102,N_19785,N_19348);
and UO_2103 (O_2103,N_19515,N_19539);
nor UO_2104 (O_2104,N_19433,N_19501);
and UO_2105 (O_2105,N_19567,N_19933);
or UO_2106 (O_2106,N_19985,N_19267);
and UO_2107 (O_2107,N_19899,N_19479);
and UO_2108 (O_2108,N_19877,N_19335);
and UO_2109 (O_2109,N_19835,N_19798);
and UO_2110 (O_2110,N_19707,N_19692);
nor UO_2111 (O_2111,N_19539,N_19350);
nor UO_2112 (O_2112,N_19845,N_19376);
or UO_2113 (O_2113,N_19845,N_19396);
nand UO_2114 (O_2114,N_19292,N_19378);
nor UO_2115 (O_2115,N_19914,N_19823);
and UO_2116 (O_2116,N_19623,N_19993);
nor UO_2117 (O_2117,N_19805,N_19897);
or UO_2118 (O_2118,N_19298,N_19998);
or UO_2119 (O_2119,N_19727,N_19349);
and UO_2120 (O_2120,N_19498,N_19291);
or UO_2121 (O_2121,N_19363,N_19390);
and UO_2122 (O_2122,N_19320,N_19322);
and UO_2123 (O_2123,N_19886,N_19841);
nand UO_2124 (O_2124,N_19738,N_19983);
nand UO_2125 (O_2125,N_19640,N_19508);
nand UO_2126 (O_2126,N_19786,N_19704);
or UO_2127 (O_2127,N_19334,N_19505);
and UO_2128 (O_2128,N_19272,N_19380);
nand UO_2129 (O_2129,N_19402,N_19870);
and UO_2130 (O_2130,N_19337,N_19391);
nor UO_2131 (O_2131,N_19445,N_19850);
or UO_2132 (O_2132,N_19838,N_19479);
nand UO_2133 (O_2133,N_19818,N_19666);
nor UO_2134 (O_2134,N_19201,N_19343);
or UO_2135 (O_2135,N_19814,N_19392);
nand UO_2136 (O_2136,N_19839,N_19651);
and UO_2137 (O_2137,N_19808,N_19282);
nor UO_2138 (O_2138,N_19586,N_19288);
and UO_2139 (O_2139,N_19360,N_19805);
nand UO_2140 (O_2140,N_19621,N_19749);
nand UO_2141 (O_2141,N_19284,N_19300);
nor UO_2142 (O_2142,N_19466,N_19290);
xnor UO_2143 (O_2143,N_19657,N_19929);
nand UO_2144 (O_2144,N_19594,N_19437);
nand UO_2145 (O_2145,N_19618,N_19222);
and UO_2146 (O_2146,N_19243,N_19668);
or UO_2147 (O_2147,N_19343,N_19639);
nor UO_2148 (O_2148,N_19302,N_19530);
xor UO_2149 (O_2149,N_19533,N_19208);
nand UO_2150 (O_2150,N_19729,N_19656);
nand UO_2151 (O_2151,N_19338,N_19654);
and UO_2152 (O_2152,N_19639,N_19387);
nor UO_2153 (O_2153,N_19997,N_19923);
and UO_2154 (O_2154,N_19394,N_19704);
nand UO_2155 (O_2155,N_19640,N_19424);
nand UO_2156 (O_2156,N_19891,N_19526);
nand UO_2157 (O_2157,N_19442,N_19652);
nand UO_2158 (O_2158,N_19336,N_19682);
or UO_2159 (O_2159,N_19301,N_19987);
and UO_2160 (O_2160,N_19417,N_19595);
nor UO_2161 (O_2161,N_19274,N_19594);
nor UO_2162 (O_2162,N_19229,N_19826);
and UO_2163 (O_2163,N_19304,N_19983);
or UO_2164 (O_2164,N_19784,N_19717);
nor UO_2165 (O_2165,N_19586,N_19954);
nor UO_2166 (O_2166,N_19391,N_19404);
and UO_2167 (O_2167,N_19540,N_19963);
and UO_2168 (O_2168,N_19657,N_19814);
and UO_2169 (O_2169,N_19290,N_19246);
and UO_2170 (O_2170,N_19293,N_19353);
or UO_2171 (O_2171,N_19350,N_19310);
or UO_2172 (O_2172,N_19541,N_19635);
nand UO_2173 (O_2173,N_19451,N_19776);
nor UO_2174 (O_2174,N_19683,N_19505);
or UO_2175 (O_2175,N_19750,N_19343);
or UO_2176 (O_2176,N_19372,N_19269);
and UO_2177 (O_2177,N_19801,N_19324);
nor UO_2178 (O_2178,N_19520,N_19377);
and UO_2179 (O_2179,N_19313,N_19382);
or UO_2180 (O_2180,N_19624,N_19354);
nand UO_2181 (O_2181,N_19501,N_19628);
or UO_2182 (O_2182,N_19787,N_19268);
and UO_2183 (O_2183,N_19551,N_19355);
and UO_2184 (O_2184,N_19237,N_19836);
or UO_2185 (O_2185,N_19815,N_19271);
nor UO_2186 (O_2186,N_19314,N_19953);
and UO_2187 (O_2187,N_19913,N_19809);
or UO_2188 (O_2188,N_19834,N_19905);
nand UO_2189 (O_2189,N_19711,N_19365);
and UO_2190 (O_2190,N_19776,N_19285);
nor UO_2191 (O_2191,N_19513,N_19520);
and UO_2192 (O_2192,N_19737,N_19667);
nand UO_2193 (O_2193,N_19584,N_19272);
xnor UO_2194 (O_2194,N_19789,N_19409);
nor UO_2195 (O_2195,N_19345,N_19886);
or UO_2196 (O_2196,N_19761,N_19375);
nor UO_2197 (O_2197,N_19711,N_19446);
nand UO_2198 (O_2198,N_19345,N_19678);
and UO_2199 (O_2199,N_19317,N_19455);
nor UO_2200 (O_2200,N_19230,N_19619);
and UO_2201 (O_2201,N_19859,N_19860);
nand UO_2202 (O_2202,N_19806,N_19593);
and UO_2203 (O_2203,N_19323,N_19645);
nor UO_2204 (O_2204,N_19334,N_19734);
or UO_2205 (O_2205,N_19249,N_19388);
or UO_2206 (O_2206,N_19514,N_19663);
and UO_2207 (O_2207,N_19292,N_19964);
nor UO_2208 (O_2208,N_19328,N_19827);
nor UO_2209 (O_2209,N_19307,N_19254);
xor UO_2210 (O_2210,N_19806,N_19357);
or UO_2211 (O_2211,N_19909,N_19859);
nand UO_2212 (O_2212,N_19898,N_19855);
nand UO_2213 (O_2213,N_19345,N_19550);
or UO_2214 (O_2214,N_19483,N_19760);
nor UO_2215 (O_2215,N_19477,N_19395);
nand UO_2216 (O_2216,N_19765,N_19340);
and UO_2217 (O_2217,N_19218,N_19457);
and UO_2218 (O_2218,N_19436,N_19900);
or UO_2219 (O_2219,N_19537,N_19433);
nor UO_2220 (O_2220,N_19370,N_19699);
nand UO_2221 (O_2221,N_19216,N_19321);
or UO_2222 (O_2222,N_19850,N_19524);
nand UO_2223 (O_2223,N_19935,N_19616);
nor UO_2224 (O_2224,N_19747,N_19684);
or UO_2225 (O_2225,N_19689,N_19741);
or UO_2226 (O_2226,N_19668,N_19345);
nor UO_2227 (O_2227,N_19945,N_19490);
and UO_2228 (O_2228,N_19804,N_19796);
nand UO_2229 (O_2229,N_19295,N_19286);
or UO_2230 (O_2230,N_19646,N_19756);
nand UO_2231 (O_2231,N_19670,N_19327);
or UO_2232 (O_2232,N_19951,N_19720);
and UO_2233 (O_2233,N_19304,N_19676);
nor UO_2234 (O_2234,N_19661,N_19886);
or UO_2235 (O_2235,N_19964,N_19946);
or UO_2236 (O_2236,N_19615,N_19387);
nand UO_2237 (O_2237,N_19588,N_19977);
or UO_2238 (O_2238,N_19353,N_19327);
and UO_2239 (O_2239,N_19624,N_19469);
nor UO_2240 (O_2240,N_19710,N_19771);
xor UO_2241 (O_2241,N_19687,N_19364);
or UO_2242 (O_2242,N_19618,N_19299);
nor UO_2243 (O_2243,N_19280,N_19339);
nor UO_2244 (O_2244,N_19618,N_19317);
nor UO_2245 (O_2245,N_19602,N_19321);
nor UO_2246 (O_2246,N_19279,N_19997);
or UO_2247 (O_2247,N_19784,N_19405);
or UO_2248 (O_2248,N_19932,N_19825);
nor UO_2249 (O_2249,N_19252,N_19899);
nor UO_2250 (O_2250,N_19818,N_19452);
and UO_2251 (O_2251,N_19345,N_19756);
nor UO_2252 (O_2252,N_19250,N_19669);
or UO_2253 (O_2253,N_19983,N_19562);
and UO_2254 (O_2254,N_19251,N_19573);
or UO_2255 (O_2255,N_19406,N_19662);
nor UO_2256 (O_2256,N_19957,N_19575);
nor UO_2257 (O_2257,N_19420,N_19505);
nand UO_2258 (O_2258,N_19659,N_19385);
nor UO_2259 (O_2259,N_19418,N_19404);
or UO_2260 (O_2260,N_19384,N_19330);
nor UO_2261 (O_2261,N_19894,N_19902);
nand UO_2262 (O_2262,N_19225,N_19687);
or UO_2263 (O_2263,N_19911,N_19883);
nor UO_2264 (O_2264,N_19783,N_19336);
nor UO_2265 (O_2265,N_19698,N_19640);
nand UO_2266 (O_2266,N_19879,N_19780);
nor UO_2267 (O_2267,N_19553,N_19677);
nor UO_2268 (O_2268,N_19274,N_19907);
and UO_2269 (O_2269,N_19649,N_19474);
and UO_2270 (O_2270,N_19212,N_19288);
nand UO_2271 (O_2271,N_19308,N_19492);
nor UO_2272 (O_2272,N_19575,N_19369);
nand UO_2273 (O_2273,N_19584,N_19225);
nand UO_2274 (O_2274,N_19228,N_19478);
nand UO_2275 (O_2275,N_19904,N_19976);
and UO_2276 (O_2276,N_19205,N_19312);
nand UO_2277 (O_2277,N_19223,N_19893);
and UO_2278 (O_2278,N_19497,N_19235);
nor UO_2279 (O_2279,N_19674,N_19755);
nand UO_2280 (O_2280,N_19302,N_19330);
or UO_2281 (O_2281,N_19205,N_19766);
or UO_2282 (O_2282,N_19370,N_19795);
or UO_2283 (O_2283,N_19764,N_19294);
and UO_2284 (O_2284,N_19558,N_19220);
or UO_2285 (O_2285,N_19694,N_19756);
nand UO_2286 (O_2286,N_19854,N_19222);
nand UO_2287 (O_2287,N_19525,N_19768);
or UO_2288 (O_2288,N_19729,N_19502);
nand UO_2289 (O_2289,N_19296,N_19823);
nor UO_2290 (O_2290,N_19917,N_19441);
or UO_2291 (O_2291,N_19880,N_19513);
and UO_2292 (O_2292,N_19691,N_19532);
nor UO_2293 (O_2293,N_19829,N_19305);
and UO_2294 (O_2294,N_19488,N_19602);
and UO_2295 (O_2295,N_19322,N_19706);
nor UO_2296 (O_2296,N_19351,N_19789);
or UO_2297 (O_2297,N_19770,N_19263);
or UO_2298 (O_2298,N_19753,N_19693);
nor UO_2299 (O_2299,N_19395,N_19369);
nand UO_2300 (O_2300,N_19541,N_19341);
and UO_2301 (O_2301,N_19841,N_19298);
nor UO_2302 (O_2302,N_19842,N_19368);
or UO_2303 (O_2303,N_19415,N_19646);
and UO_2304 (O_2304,N_19253,N_19270);
and UO_2305 (O_2305,N_19432,N_19769);
nand UO_2306 (O_2306,N_19637,N_19759);
nand UO_2307 (O_2307,N_19523,N_19962);
or UO_2308 (O_2308,N_19845,N_19445);
nor UO_2309 (O_2309,N_19729,N_19202);
and UO_2310 (O_2310,N_19379,N_19434);
nand UO_2311 (O_2311,N_19273,N_19514);
and UO_2312 (O_2312,N_19231,N_19326);
and UO_2313 (O_2313,N_19588,N_19439);
and UO_2314 (O_2314,N_19399,N_19406);
nand UO_2315 (O_2315,N_19770,N_19327);
and UO_2316 (O_2316,N_19474,N_19697);
and UO_2317 (O_2317,N_19261,N_19611);
or UO_2318 (O_2318,N_19931,N_19288);
nor UO_2319 (O_2319,N_19271,N_19456);
nand UO_2320 (O_2320,N_19362,N_19591);
nor UO_2321 (O_2321,N_19289,N_19476);
or UO_2322 (O_2322,N_19870,N_19465);
or UO_2323 (O_2323,N_19314,N_19366);
nor UO_2324 (O_2324,N_19565,N_19502);
nand UO_2325 (O_2325,N_19909,N_19792);
nand UO_2326 (O_2326,N_19368,N_19453);
and UO_2327 (O_2327,N_19285,N_19295);
or UO_2328 (O_2328,N_19612,N_19373);
nand UO_2329 (O_2329,N_19405,N_19249);
xnor UO_2330 (O_2330,N_19334,N_19206);
nand UO_2331 (O_2331,N_19679,N_19917);
nor UO_2332 (O_2332,N_19433,N_19892);
nor UO_2333 (O_2333,N_19535,N_19258);
and UO_2334 (O_2334,N_19483,N_19489);
nand UO_2335 (O_2335,N_19962,N_19612);
nand UO_2336 (O_2336,N_19994,N_19227);
or UO_2337 (O_2337,N_19516,N_19887);
and UO_2338 (O_2338,N_19749,N_19885);
and UO_2339 (O_2339,N_19744,N_19551);
or UO_2340 (O_2340,N_19462,N_19883);
nor UO_2341 (O_2341,N_19781,N_19590);
nor UO_2342 (O_2342,N_19289,N_19296);
nand UO_2343 (O_2343,N_19611,N_19804);
and UO_2344 (O_2344,N_19482,N_19558);
nand UO_2345 (O_2345,N_19592,N_19576);
nand UO_2346 (O_2346,N_19737,N_19957);
and UO_2347 (O_2347,N_19630,N_19867);
nand UO_2348 (O_2348,N_19800,N_19890);
or UO_2349 (O_2349,N_19573,N_19282);
nand UO_2350 (O_2350,N_19634,N_19950);
or UO_2351 (O_2351,N_19885,N_19823);
or UO_2352 (O_2352,N_19259,N_19429);
nor UO_2353 (O_2353,N_19404,N_19306);
nor UO_2354 (O_2354,N_19243,N_19926);
nor UO_2355 (O_2355,N_19653,N_19421);
nand UO_2356 (O_2356,N_19767,N_19268);
nor UO_2357 (O_2357,N_19867,N_19672);
and UO_2358 (O_2358,N_19288,N_19258);
nand UO_2359 (O_2359,N_19823,N_19577);
nand UO_2360 (O_2360,N_19314,N_19604);
or UO_2361 (O_2361,N_19723,N_19995);
or UO_2362 (O_2362,N_19423,N_19463);
nand UO_2363 (O_2363,N_19682,N_19681);
nand UO_2364 (O_2364,N_19419,N_19837);
nor UO_2365 (O_2365,N_19457,N_19370);
nand UO_2366 (O_2366,N_19232,N_19943);
nand UO_2367 (O_2367,N_19587,N_19527);
and UO_2368 (O_2368,N_19615,N_19804);
or UO_2369 (O_2369,N_19423,N_19302);
and UO_2370 (O_2370,N_19476,N_19347);
and UO_2371 (O_2371,N_19735,N_19754);
nand UO_2372 (O_2372,N_19345,N_19233);
nor UO_2373 (O_2373,N_19569,N_19686);
or UO_2374 (O_2374,N_19429,N_19361);
nand UO_2375 (O_2375,N_19807,N_19618);
nand UO_2376 (O_2376,N_19704,N_19472);
nor UO_2377 (O_2377,N_19859,N_19247);
and UO_2378 (O_2378,N_19994,N_19305);
nand UO_2379 (O_2379,N_19218,N_19868);
nand UO_2380 (O_2380,N_19866,N_19948);
nand UO_2381 (O_2381,N_19779,N_19532);
or UO_2382 (O_2382,N_19457,N_19590);
nor UO_2383 (O_2383,N_19467,N_19256);
or UO_2384 (O_2384,N_19747,N_19284);
nor UO_2385 (O_2385,N_19547,N_19932);
nand UO_2386 (O_2386,N_19714,N_19880);
nand UO_2387 (O_2387,N_19431,N_19618);
and UO_2388 (O_2388,N_19345,N_19805);
xnor UO_2389 (O_2389,N_19759,N_19849);
or UO_2390 (O_2390,N_19562,N_19202);
xor UO_2391 (O_2391,N_19604,N_19562);
and UO_2392 (O_2392,N_19775,N_19870);
and UO_2393 (O_2393,N_19984,N_19497);
nor UO_2394 (O_2394,N_19392,N_19661);
and UO_2395 (O_2395,N_19236,N_19861);
nand UO_2396 (O_2396,N_19756,N_19421);
nor UO_2397 (O_2397,N_19823,N_19990);
or UO_2398 (O_2398,N_19475,N_19343);
nor UO_2399 (O_2399,N_19866,N_19555);
and UO_2400 (O_2400,N_19443,N_19481);
nor UO_2401 (O_2401,N_19645,N_19294);
nor UO_2402 (O_2402,N_19450,N_19620);
or UO_2403 (O_2403,N_19991,N_19927);
or UO_2404 (O_2404,N_19640,N_19431);
nor UO_2405 (O_2405,N_19285,N_19698);
nor UO_2406 (O_2406,N_19753,N_19289);
nand UO_2407 (O_2407,N_19349,N_19725);
or UO_2408 (O_2408,N_19496,N_19820);
and UO_2409 (O_2409,N_19920,N_19752);
xor UO_2410 (O_2410,N_19914,N_19225);
and UO_2411 (O_2411,N_19428,N_19379);
or UO_2412 (O_2412,N_19457,N_19695);
and UO_2413 (O_2413,N_19244,N_19694);
and UO_2414 (O_2414,N_19316,N_19738);
nor UO_2415 (O_2415,N_19467,N_19407);
xor UO_2416 (O_2416,N_19787,N_19308);
nand UO_2417 (O_2417,N_19468,N_19418);
nor UO_2418 (O_2418,N_19838,N_19759);
or UO_2419 (O_2419,N_19481,N_19421);
nor UO_2420 (O_2420,N_19739,N_19939);
nor UO_2421 (O_2421,N_19852,N_19729);
nand UO_2422 (O_2422,N_19769,N_19414);
nor UO_2423 (O_2423,N_19200,N_19685);
nor UO_2424 (O_2424,N_19427,N_19998);
nand UO_2425 (O_2425,N_19970,N_19686);
nand UO_2426 (O_2426,N_19398,N_19702);
nor UO_2427 (O_2427,N_19529,N_19507);
nand UO_2428 (O_2428,N_19532,N_19387);
nor UO_2429 (O_2429,N_19340,N_19614);
or UO_2430 (O_2430,N_19288,N_19498);
and UO_2431 (O_2431,N_19260,N_19400);
nor UO_2432 (O_2432,N_19831,N_19700);
nor UO_2433 (O_2433,N_19680,N_19492);
and UO_2434 (O_2434,N_19447,N_19927);
nand UO_2435 (O_2435,N_19732,N_19560);
nand UO_2436 (O_2436,N_19525,N_19547);
or UO_2437 (O_2437,N_19997,N_19891);
nor UO_2438 (O_2438,N_19396,N_19654);
nor UO_2439 (O_2439,N_19685,N_19488);
nor UO_2440 (O_2440,N_19946,N_19986);
nor UO_2441 (O_2441,N_19438,N_19567);
nand UO_2442 (O_2442,N_19402,N_19941);
and UO_2443 (O_2443,N_19397,N_19635);
and UO_2444 (O_2444,N_19254,N_19493);
or UO_2445 (O_2445,N_19944,N_19278);
and UO_2446 (O_2446,N_19855,N_19885);
and UO_2447 (O_2447,N_19359,N_19613);
nand UO_2448 (O_2448,N_19572,N_19532);
nor UO_2449 (O_2449,N_19299,N_19980);
and UO_2450 (O_2450,N_19339,N_19818);
nand UO_2451 (O_2451,N_19981,N_19879);
nand UO_2452 (O_2452,N_19272,N_19329);
or UO_2453 (O_2453,N_19376,N_19958);
and UO_2454 (O_2454,N_19581,N_19248);
or UO_2455 (O_2455,N_19633,N_19732);
or UO_2456 (O_2456,N_19350,N_19945);
nand UO_2457 (O_2457,N_19725,N_19982);
nor UO_2458 (O_2458,N_19205,N_19578);
nand UO_2459 (O_2459,N_19607,N_19332);
or UO_2460 (O_2460,N_19987,N_19377);
or UO_2461 (O_2461,N_19381,N_19881);
or UO_2462 (O_2462,N_19218,N_19237);
nor UO_2463 (O_2463,N_19493,N_19960);
nand UO_2464 (O_2464,N_19225,N_19626);
nor UO_2465 (O_2465,N_19628,N_19909);
or UO_2466 (O_2466,N_19849,N_19554);
nand UO_2467 (O_2467,N_19763,N_19557);
nand UO_2468 (O_2468,N_19456,N_19932);
nor UO_2469 (O_2469,N_19538,N_19680);
or UO_2470 (O_2470,N_19677,N_19810);
and UO_2471 (O_2471,N_19456,N_19302);
nand UO_2472 (O_2472,N_19338,N_19423);
nor UO_2473 (O_2473,N_19239,N_19669);
nand UO_2474 (O_2474,N_19760,N_19606);
nor UO_2475 (O_2475,N_19405,N_19788);
and UO_2476 (O_2476,N_19898,N_19600);
nor UO_2477 (O_2477,N_19901,N_19895);
and UO_2478 (O_2478,N_19517,N_19599);
nor UO_2479 (O_2479,N_19330,N_19264);
or UO_2480 (O_2480,N_19624,N_19290);
and UO_2481 (O_2481,N_19288,N_19500);
and UO_2482 (O_2482,N_19551,N_19637);
and UO_2483 (O_2483,N_19613,N_19692);
nor UO_2484 (O_2484,N_19935,N_19810);
nand UO_2485 (O_2485,N_19396,N_19472);
nor UO_2486 (O_2486,N_19387,N_19280);
nor UO_2487 (O_2487,N_19996,N_19691);
or UO_2488 (O_2488,N_19453,N_19242);
xor UO_2489 (O_2489,N_19318,N_19945);
nor UO_2490 (O_2490,N_19908,N_19793);
nor UO_2491 (O_2491,N_19774,N_19775);
nand UO_2492 (O_2492,N_19208,N_19407);
or UO_2493 (O_2493,N_19712,N_19809);
or UO_2494 (O_2494,N_19398,N_19384);
nand UO_2495 (O_2495,N_19690,N_19483);
and UO_2496 (O_2496,N_19776,N_19338);
and UO_2497 (O_2497,N_19800,N_19266);
xnor UO_2498 (O_2498,N_19928,N_19845);
or UO_2499 (O_2499,N_19873,N_19213);
endmodule