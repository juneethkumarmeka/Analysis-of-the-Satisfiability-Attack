module basic_1000_10000_1500_100_levels_10xor_5(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999;
xnor U0 (N_0,In_837,In_752);
nor U1 (N_1,In_588,In_912);
nand U2 (N_2,In_304,In_476);
nor U3 (N_3,In_737,In_964);
or U4 (N_4,In_281,In_343);
or U5 (N_5,In_832,In_215);
xnor U6 (N_6,In_455,In_928);
nand U7 (N_7,In_448,In_956);
and U8 (N_8,In_214,In_623);
xnor U9 (N_9,In_272,In_469);
and U10 (N_10,In_236,In_449);
and U11 (N_11,In_187,In_653);
nand U12 (N_12,In_447,In_855);
xnor U13 (N_13,In_1,In_435);
nor U14 (N_14,In_944,In_471);
nand U15 (N_15,In_152,In_287);
and U16 (N_16,In_799,In_38);
or U17 (N_17,In_609,In_58);
xnor U18 (N_18,In_725,In_717);
nor U19 (N_19,In_391,In_104);
and U20 (N_20,In_267,In_950);
and U21 (N_21,In_11,In_536);
nor U22 (N_22,In_194,In_617);
xor U23 (N_23,In_744,In_923);
nor U24 (N_24,In_999,In_315);
xnor U25 (N_25,In_513,In_254);
and U26 (N_26,In_940,In_19);
xor U27 (N_27,In_136,In_683);
nand U28 (N_28,In_419,In_137);
nor U29 (N_29,In_125,In_258);
nand U30 (N_30,In_159,In_169);
and U31 (N_31,In_650,In_547);
xnor U32 (N_32,In_972,In_568);
nor U33 (N_33,In_577,In_593);
or U34 (N_34,In_569,In_616);
or U35 (N_35,In_199,In_161);
or U36 (N_36,In_173,In_835);
and U37 (N_37,In_308,In_635);
xnor U38 (N_38,In_76,In_882);
xnor U39 (N_39,In_396,In_771);
nand U40 (N_40,In_28,In_528);
nor U41 (N_41,In_442,In_997);
nand U42 (N_42,In_458,In_305);
and U43 (N_43,In_671,In_175);
nor U44 (N_44,In_823,In_792);
nor U45 (N_45,In_81,In_255);
or U46 (N_46,In_981,In_530);
nand U47 (N_47,In_693,In_193);
nor U48 (N_48,In_402,In_178);
and U49 (N_49,In_0,In_498);
nand U50 (N_50,In_390,In_25);
xor U51 (N_51,In_116,In_167);
nand U52 (N_52,In_910,In_660);
xor U53 (N_53,In_526,In_993);
and U54 (N_54,In_144,In_603);
or U55 (N_55,In_392,In_895);
or U56 (N_56,In_395,In_793);
or U57 (N_57,In_45,In_881);
nor U58 (N_58,In_439,In_283);
or U59 (N_59,In_428,In_244);
nand U60 (N_60,In_292,In_93);
nand U61 (N_61,In_774,In_559);
xnor U62 (N_62,In_711,In_704);
and U63 (N_63,In_658,In_755);
xnor U64 (N_64,In_840,In_994);
nand U65 (N_65,In_628,In_301);
nand U66 (N_66,In_566,In_669);
and U67 (N_67,In_812,In_631);
nor U68 (N_68,In_539,In_730);
and U69 (N_69,In_845,In_722);
nand U70 (N_70,In_432,In_443);
or U71 (N_71,In_885,In_649);
nor U72 (N_72,In_801,In_239);
xor U73 (N_73,In_815,In_60);
or U74 (N_74,In_374,In_461);
xnor U75 (N_75,In_268,In_376);
or U76 (N_76,In_777,In_366);
nand U77 (N_77,In_772,In_445);
nor U78 (N_78,In_869,In_791);
nand U79 (N_79,In_219,In_942);
xor U80 (N_80,In_618,In_949);
xor U81 (N_81,In_784,In_259);
nor U82 (N_82,In_652,In_94);
xor U83 (N_83,In_499,In_251);
and U84 (N_84,In_921,In_90);
and U85 (N_85,In_758,In_110);
or U86 (N_86,In_647,In_984);
nand U87 (N_87,In_800,In_998);
nor U88 (N_88,In_838,In_676);
nor U89 (N_89,In_555,In_30);
xnor U90 (N_90,In_198,In_665);
nand U91 (N_91,In_467,In_421);
or U92 (N_92,In_284,In_70);
or U93 (N_93,In_824,In_311);
or U94 (N_94,In_702,In_870);
xnor U95 (N_95,In_10,In_830);
nor U96 (N_96,In_289,In_403);
or U97 (N_97,In_645,In_68);
or U98 (N_98,In_222,In_889);
nor U99 (N_99,In_487,In_627);
nand U100 (N_100,In_86,In_378);
and U101 (N_101,In_692,In_629);
and U102 (N_102,In_92,In_689);
nor U103 (N_103,N_91,N_75);
nand U104 (N_104,In_15,N_74);
xor U105 (N_105,In_328,In_831);
or U106 (N_106,In_166,In_765);
nor U107 (N_107,In_242,In_454);
or U108 (N_108,N_50,In_365);
or U109 (N_109,In_651,In_899);
xor U110 (N_110,In_249,In_579);
xor U111 (N_111,In_333,In_231);
xor U112 (N_112,In_856,In_462);
xnor U113 (N_113,In_280,In_210);
and U114 (N_114,In_423,In_560);
nand U115 (N_115,N_72,In_522);
xnor U116 (N_116,In_174,In_779);
nand U117 (N_117,In_293,N_82);
xor U118 (N_118,In_191,In_973);
or U119 (N_119,In_868,In_633);
and U120 (N_120,N_31,In_786);
and U121 (N_121,In_608,In_361);
nor U122 (N_122,In_794,N_57);
nor U123 (N_123,In_319,N_19);
or U124 (N_124,In_426,In_269);
nand U125 (N_125,In_313,In_74);
and U126 (N_126,In_575,In_22);
xor U127 (N_127,In_8,In_596);
xnor U128 (N_128,In_873,In_584);
nand U129 (N_129,In_122,In_389);
nor U130 (N_130,In_783,In_14);
and U131 (N_131,N_42,In_678);
nand U132 (N_132,In_156,N_51);
and U133 (N_133,In_517,In_553);
and U134 (N_134,In_197,In_907);
and U135 (N_135,In_80,In_637);
nor U136 (N_136,In_282,In_5);
nand U137 (N_137,In_848,In_183);
and U138 (N_138,In_728,In_252);
nor U139 (N_139,In_422,In_814);
nand U140 (N_140,In_27,In_501);
xor U141 (N_141,In_71,In_370);
nand U142 (N_142,In_126,In_531);
xnor U143 (N_143,N_56,In_908);
or U144 (N_144,In_84,In_803);
nor U145 (N_145,In_24,In_929);
or U146 (N_146,In_226,In_682);
nor U147 (N_147,In_241,In_773);
nor U148 (N_148,In_906,In_766);
nand U149 (N_149,N_21,N_95);
nor U150 (N_150,In_349,In_288);
xnor U151 (N_151,In_695,In_638);
nor U152 (N_152,In_549,In_300);
nor U153 (N_153,In_79,N_20);
and U154 (N_154,In_317,In_232);
xnor U155 (N_155,N_69,N_58);
nand U156 (N_156,N_1,In_844);
or U157 (N_157,In_385,In_897);
and U158 (N_158,In_35,In_595);
nor U159 (N_159,In_586,In_83);
nand U160 (N_160,In_229,In_453);
xnor U161 (N_161,In_516,In_820);
nor U162 (N_162,In_271,In_223);
or U163 (N_163,N_61,In_257);
xnor U164 (N_164,In_53,In_731);
or U165 (N_165,In_337,In_431);
or U166 (N_166,In_277,In_141);
nand U167 (N_167,In_974,In_310);
and U168 (N_168,N_40,In_464);
and U169 (N_169,In_312,In_514);
or U170 (N_170,In_713,In_642);
or U171 (N_171,In_871,N_47);
xor U172 (N_172,In_238,In_452);
nand U173 (N_173,In_630,In_346);
xnor U174 (N_174,In_276,In_7);
nand U175 (N_175,In_880,In_32);
or U176 (N_176,In_55,In_170);
xnor U177 (N_177,In_316,In_357);
nand U178 (N_178,In_508,In_734);
nand U179 (N_179,In_967,In_935);
nor U180 (N_180,In_567,In_200);
nor U181 (N_181,In_675,In_988);
nor U182 (N_182,In_359,N_79);
xnor U183 (N_183,In_741,In_966);
nor U184 (N_184,In_331,In_933);
or U185 (N_185,In_205,In_996);
or U186 (N_186,In_163,In_479);
nand U187 (N_187,N_67,In_106);
nand U188 (N_188,In_770,In_474);
and U189 (N_189,In_490,In_158);
or U190 (N_190,In_580,In_892);
or U191 (N_191,In_925,In_781);
or U192 (N_192,In_959,In_457);
nor U193 (N_193,In_668,In_404);
or U194 (N_194,N_84,In_594);
or U195 (N_195,In_424,In_934);
and U196 (N_196,In_203,In_667);
nor U197 (N_197,In_468,In_118);
nand U198 (N_198,In_648,In_138);
nand U199 (N_199,In_919,In_738);
or U200 (N_200,In_411,In_550);
and U201 (N_201,N_59,N_76);
nand U202 (N_202,N_130,In_545);
or U203 (N_203,In_839,In_565);
xor U204 (N_204,N_142,In_583);
and U205 (N_205,In_177,In_684);
xnor U206 (N_206,In_813,In_336);
and U207 (N_207,In_548,In_506);
nand U208 (N_208,In_930,In_209);
xnor U209 (N_209,In_952,N_107);
or U210 (N_210,In_57,In_915);
xor U211 (N_211,In_822,In_495);
nand U212 (N_212,In_825,N_169);
or U213 (N_213,In_763,In_380);
xor U214 (N_214,In_903,N_196);
nand U215 (N_215,In_444,In_554);
and U216 (N_216,N_116,N_88);
and U217 (N_217,In_379,In_523);
xor U218 (N_218,In_4,In_393);
or U219 (N_219,In_485,N_103);
nor U220 (N_220,In_878,In_278);
nand U221 (N_221,N_12,In_805);
xnor U222 (N_222,In_342,In_954);
nand U223 (N_223,N_23,In_698);
and U224 (N_224,N_183,In_953);
or U225 (N_225,In_334,In_503);
and U226 (N_226,In_371,In_329);
and U227 (N_227,In_425,In_847);
nand U228 (N_228,In_165,N_45);
nor U229 (N_229,N_155,N_176);
or U230 (N_230,In_482,N_16);
nand U231 (N_231,N_70,In_400);
or U232 (N_232,In_821,In_888);
xnor U233 (N_233,In_348,In_240);
xor U234 (N_234,N_98,In_386);
nor U235 (N_235,In_49,In_286);
nor U236 (N_236,In_733,N_141);
xor U237 (N_237,In_440,In_742);
and U238 (N_238,In_557,In_480);
nand U239 (N_239,In_775,In_123);
xor U240 (N_240,In_512,In_26);
and U241 (N_241,In_417,In_463);
nand U242 (N_242,In_625,In_207);
nand U243 (N_243,In_989,In_597);
nor U244 (N_244,N_14,N_182);
xor U245 (N_245,In_275,In_97);
nand U246 (N_246,In_63,In_397);
and U247 (N_247,In_641,In_927);
nor U248 (N_248,In_690,In_708);
and U249 (N_249,In_811,In_938);
xnor U250 (N_250,In_230,In_573);
xor U251 (N_251,In_353,In_410);
and U252 (N_252,In_634,In_978);
and U253 (N_253,In_686,In_932);
or U254 (N_254,In_296,N_99);
or U255 (N_255,In_279,In_714);
nand U256 (N_256,N_78,In_322);
nand U257 (N_257,In_904,In_291);
nor U258 (N_258,In_795,N_53);
and U259 (N_259,In_192,In_561);
and U260 (N_260,In_502,In_963);
xor U261 (N_261,In_558,In_128);
xor U262 (N_262,In_412,In_891);
and U263 (N_263,In_767,In_681);
and U264 (N_264,In_436,In_802);
xor U265 (N_265,In_700,In_228);
nor U266 (N_266,In_664,In_88);
nor U267 (N_267,N_139,N_73);
xor U268 (N_268,In_434,In_105);
nand U269 (N_269,In_872,N_127);
nor U270 (N_270,In_544,In_829);
nand U271 (N_271,In_75,In_510);
xor U272 (N_272,In_776,N_97);
xor U273 (N_273,In_537,In_253);
nand U274 (N_274,In_739,In_82);
nand U275 (N_275,In_44,In_644);
and U276 (N_276,In_819,In_12);
nor U277 (N_277,N_46,In_245);
or U278 (N_278,N_151,N_64);
and U279 (N_279,In_540,In_612);
xor U280 (N_280,In_656,In_43);
nand U281 (N_281,N_124,N_118);
or U282 (N_282,In_902,In_626);
and U283 (N_283,In_754,In_712);
nand U284 (N_284,In_201,N_62);
and U285 (N_285,In_862,In_362);
nand U286 (N_286,In_188,N_122);
or U287 (N_287,N_184,In_373);
nand U288 (N_288,In_751,In_894);
nand U289 (N_289,In_901,N_152);
nor U290 (N_290,N_161,In_475);
nand U291 (N_291,In_108,In_808);
and U292 (N_292,In_451,In_607);
or U293 (N_293,In_429,In_858);
nor U294 (N_294,In_914,N_109);
xnor U295 (N_295,In_17,N_4);
and U296 (N_296,In_796,In_13);
nand U297 (N_297,N_160,In_971);
xnor U298 (N_298,In_157,In_538);
or U299 (N_299,In_500,In_399);
xor U300 (N_300,N_266,In_21);
nor U301 (N_301,In_217,N_270);
xnor U302 (N_302,In_661,In_91);
or U303 (N_303,N_128,N_110);
and U304 (N_304,N_112,In_89);
or U305 (N_305,In_854,In_941);
or U306 (N_306,In_33,In_34);
nand U307 (N_307,In_290,N_35);
or U308 (N_308,N_30,In_606);
nor U309 (N_309,In_325,In_127);
xnor U310 (N_310,In_833,In_976);
and U311 (N_311,In_666,In_350);
and U312 (N_312,In_320,N_167);
xor U313 (N_313,N_229,In_706);
or U314 (N_314,In_955,N_81);
and U315 (N_315,N_195,In_716);
nor U316 (N_316,N_34,In_204);
or U317 (N_317,In_114,N_290);
or U318 (N_318,N_234,In_248);
nand U319 (N_319,N_9,N_163);
nor U320 (N_320,In_578,In_154);
nor U321 (N_321,In_715,In_562);
and U322 (N_322,N_179,In_330);
and U323 (N_323,N_285,N_241);
or U324 (N_324,In_41,N_252);
nor U325 (N_325,In_149,N_37);
and U326 (N_326,In_979,N_221);
xnor U327 (N_327,In_190,In_103);
nand U328 (N_328,In_657,N_213);
nand U329 (N_329,N_232,In_563);
or U330 (N_330,In_29,In_383);
xnor U331 (N_331,In_401,In_576);
xnor U332 (N_332,In_757,In_619);
xor U333 (N_333,N_224,In_504);
and U334 (N_334,In_769,In_64);
nor U335 (N_335,N_39,In_340);
xnor U336 (N_336,In_418,In_990);
nand U337 (N_337,N_111,In_905);
or U338 (N_338,In_18,N_41);
and U339 (N_339,In_797,In_99);
nand U340 (N_340,In_977,In_851);
nand U341 (N_341,In_827,In_727);
nor U342 (N_342,In_818,In_785);
and U343 (N_343,N_233,N_96);
nand U344 (N_344,N_89,N_90);
or U345 (N_345,In_505,In_655);
and U346 (N_346,N_185,N_106);
and U347 (N_347,N_120,In_176);
nand U348 (N_348,N_7,In_816);
nor U349 (N_349,In_124,N_68);
xor U350 (N_350,In_195,In_931);
xnor U351 (N_351,In_151,In_867);
or U352 (N_352,In_314,N_220);
nor U353 (N_353,In_16,In_863);
nand U354 (N_354,N_131,N_134);
nor U355 (N_355,N_236,In_162);
nor U356 (N_356,In_624,N_216);
xnor U357 (N_357,N_256,In_51);
nor U358 (N_358,In_111,In_677);
nor U359 (N_359,N_71,N_284);
nor U360 (N_360,In_788,In_970);
nand U361 (N_361,In_360,In_859);
or U362 (N_362,In_581,In_384);
and U363 (N_363,In_218,N_114);
and U364 (N_364,N_294,In_220);
and U365 (N_365,In_48,In_817);
xnor U366 (N_366,In_438,In_145);
and U367 (N_367,N_173,In_102);
xor U368 (N_368,N_295,In_893);
xnor U369 (N_369,In_377,In_787);
xor U370 (N_370,N_104,N_210);
or U371 (N_371,In_171,In_213);
or U372 (N_372,In_918,In_968);
and U373 (N_373,N_247,N_86);
nand U374 (N_374,In_143,N_65);
nor U375 (N_375,N_276,N_254);
nand U376 (N_376,In_992,In_225);
nor U377 (N_377,In_488,In_496);
nor U378 (N_378,N_299,N_145);
nor U379 (N_379,N_94,In_142);
nor U380 (N_380,N_48,In_745);
xor U381 (N_381,In_810,N_255);
and U382 (N_382,In_726,In_909);
and U383 (N_383,In_759,In_420);
and U384 (N_384,N_49,N_293);
or U385 (N_385,In_985,N_192);
and U386 (N_386,N_244,In_615);
nor U387 (N_387,N_148,In_147);
or U388 (N_388,In_890,In_306);
xor U389 (N_389,N_87,In_153);
and U390 (N_390,In_266,In_599);
xor U391 (N_391,In_489,In_592);
nor U392 (N_392,N_105,N_267);
and U393 (N_393,In_69,In_355);
nand U394 (N_394,N_248,N_217);
nand U395 (N_395,N_194,In_509);
and U396 (N_396,N_162,In_408);
and U397 (N_397,In_78,In_674);
nand U398 (N_398,In_721,In_323);
xor U399 (N_399,In_246,In_427);
nand U400 (N_400,N_117,N_157);
xor U401 (N_401,In_570,N_239);
nor U402 (N_402,N_260,N_159);
nor U403 (N_403,In_224,In_247);
nor U404 (N_404,N_135,N_323);
or U405 (N_405,In_962,N_150);
nor U406 (N_406,N_358,N_357);
xor U407 (N_407,N_231,In_764);
nor U408 (N_408,In_875,In_261);
or U409 (N_409,In_98,In_129);
or U410 (N_410,In_636,In_62);
or U411 (N_411,In_564,N_380);
and U412 (N_412,N_273,N_168);
or U413 (N_413,N_129,In_294);
and U414 (N_414,In_916,N_360);
xnor U415 (N_415,N_33,In_729);
or U416 (N_416,In_233,In_743);
and U417 (N_417,N_100,In_332);
or U418 (N_418,In_663,N_296);
and U419 (N_419,In_23,In_756);
xnor U420 (N_420,In_208,In_874);
xor U421 (N_421,In_46,In_849);
xor U422 (N_422,N_342,In_478);
nor U423 (N_423,In_843,In_216);
and U424 (N_424,In_39,In_459);
nor U425 (N_425,In_552,In_96);
nand U426 (N_426,In_265,N_92);
xnor U427 (N_427,In_632,N_251);
nor U428 (N_428,In_600,In_836);
nor U429 (N_429,N_376,In_639);
or U430 (N_430,In_87,N_237);
nand U431 (N_431,In_446,In_234);
nor U432 (N_432,In_250,In_66);
and U433 (N_433,In_995,N_17);
and U434 (N_434,N_337,N_271);
or U435 (N_435,In_969,In_413);
xnor U436 (N_436,N_43,In_120);
xnor U437 (N_437,In_9,In_227);
and U438 (N_438,In_181,In_132);
and U439 (N_439,In_768,In_605);
nor U440 (N_440,N_303,In_318);
and U441 (N_441,In_943,In_922);
and U442 (N_442,In_338,N_102);
nand U443 (N_443,In_50,In_95);
nor U444 (N_444,In_256,In_351);
xnor U445 (N_445,N_26,In_611);
xnor U446 (N_446,In_524,N_138);
and U447 (N_447,N_370,In_375);
and U448 (N_448,In_551,In_507);
or U449 (N_449,N_378,N_190);
or U450 (N_450,In_946,N_166);
nand U451 (N_451,N_329,In_324);
or U452 (N_452,N_18,In_134);
xor U453 (N_453,In_986,In_659);
nor U454 (N_454,N_334,N_274);
nand U455 (N_455,In_465,N_8);
or U456 (N_456,In_735,N_340);
nand U457 (N_457,N_347,In_913);
or U458 (N_458,In_621,In_975);
xor U459 (N_459,N_60,N_202);
xor U460 (N_460,N_396,N_77);
and U461 (N_461,In_493,In_694);
or U462 (N_462,N_363,In_834);
or U463 (N_463,In_965,In_852);
or U464 (N_464,In_980,N_101);
nor U465 (N_465,N_140,In_521);
nand U466 (N_466,In_42,N_52);
nor U467 (N_467,N_275,In_347);
and U468 (N_468,N_388,N_258);
nand U469 (N_469,In_100,N_15);
xnor U470 (N_470,In_541,N_136);
nand U471 (N_471,In_520,N_355);
or U472 (N_472,N_149,In_515);
or U473 (N_473,In_67,N_392);
xor U474 (N_474,In_243,In_719);
xnor U475 (N_475,In_723,N_200);
or U476 (N_476,N_143,N_368);
and U477 (N_477,N_126,N_364);
nand U478 (N_478,N_191,N_304);
or U479 (N_479,In_470,N_158);
and U480 (N_480,N_399,N_343);
xnor U481 (N_481,In_101,In_168);
xnor U482 (N_482,N_319,In_481);
or U483 (N_483,N_390,N_333);
nand U484 (N_484,N_375,In_860);
and U485 (N_485,N_310,In_61);
and U486 (N_486,In_691,In_673);
or U487 (N_487,N_208,In_703);
nor U488 (N_488,N_356,In_662);
nor U489 (N_489,N_309,In_117);
xor U490 (N_490,In_363,In_887);
or U491 (N_491,In_133,In_842);
and U492 (N_492,N_345,N_223);
or U493 (N_493,N_315,N_242);
or U494 (N_494,In_680,In_525);
and U495 (N_495,In_148,In_947);
xor U496 (N_496,In_358,N_336);
nand U497 (N_497,In_688,In_937);
nand U498 (N_498,In_491,In_534);
xnor U499 (N_499,N_377,N_339);
and U500 (N_500,N_259,N_331);
nand U501 (N_501,In_598,N_414);
or U502 (N_502,N_431,N_415);
nor U503 (N_503,In_879,In_518);
or U504 (N_504,N_123,In_221);
nor U505 (N_505,In_483,In_303);
nand U506 (N_506,In_3,In_760);
and U507 (N_507,In_211,In_622);
or U508 (N_508,In_709,In_896);
nor U509 (N_509,N_230,In_533);
nand U510 (N_510,In_546,N_379);
xor U511 (N_511,In_920,N_235);
and U512 (N_512,N_286,In_160);
nor U513 (N_513,N_205,In_52);
nand U514 (N_514,In_382,In_782);
nor U515 (N_515,N_463,In_585);
or U516 (N_516,N_307,In_73);
or U517 (N_517,In_556,N_426);
nor U518 (N_518,N_466,In_273);
nand U519 (N_519,In_237,N_383);
xnor U520 (N_520,In_262,N_344);
nand U521 (N_521,In_535,N_288);
nor U522 (N_522,In_139,In_884);
nand U523 (N_523,N_429,N_38);
nor U524 (N_524,N_3,N_289);
nand U525 (N_525,N_312,N_197);
or U526 (N_526,N_215,In_460);
nand U527 (N_527,N_409,N_434);
and U528 (N_528,In_749,N_257);
nand U529 (N_529,In_807,In_936);
or U530 (N_530,N_449,In_65);
and U531 (N_531,N_13,N_448);
xor U532 (N_532,In_699,N_172);
xor U533 (N_533,In_924,N_402);
or U534 (N_534,In_672,In_394);
nor U535 (N_535,N_490,In_846);
nor U536 (N_536,N_228,In_841);
or U537 (N_537,N_214,In_352);
and U538 (N_538,N_367,N_486);
or U539 (N_539,N_253,In_433);
or U540 (N_540,In_687,N_207);
nand U541 (N_541,In_960,In_643);
nor U542 (N_542,In_235,N_411);
or U543 (N_543,N_218,N_459);
xnor U544 (N_544,In_987,In_718);
nor U545 (N_545,In_155,N_445);
or U546 (N_546,In_130,In_297);
and U547 (N_547,In_298,N_262);
nand U548 (N_548,N_461,N_25);
xor U549 (N_549,N_427,N_22);
or U550 (N_550,N_322,In_701);
xnor U551 (N_551,N_397,N_361);
nand U552 (N_552,N_327,In_184);
or U553 (N_553,N_417,N_308);
nand U554 (N_554,N_133,In_112);
nor U555 (N_555,In_762,In_886);
or U556 (N_556,In_59,N_470);
xnor U557 (N_557,In_206,In_415);
or U558 (N_558,In_260,N_226);
or U559 (N_559,In_604,In_414);
xor U560 (N_560,N_272,In_724);
nand U561 (N_561,N_297,In_646);
nor U562 (N_562,In_542,In_911);
and U563 (N_563,N_119,In_778);
and U564 (N_564,N_443,N_475);
nor U565 (N_565,In_640,N_264);
and U566 (N_566,N_291,In_339);
nor U567 (N_567,N_206,N_468);
nor U568 (N_568,In_409,In_179);
or U569 (N_569,In_532,N_212);
nor U570 (N_570,N_187,N_432);
nor U571 (N_571,N_0,In_335);
nor U572 (N_572,N_428,N_467);
nand U573 (N_573,N_211,In_602);
xor U574 (N_574,N_209,N_404);
or U575 (N_575,In_654,N_365);
nor U576 (N_576,N_325,In_20);
xnor U577 (N_577,In_790,In_345);
nand U578 (N_578,In_857,N_283);
and U579 (N_579,N_317,N_341);
or U580 (N_580,N_125,In_828);
nor U581 (N_581,N_451,In_850);
xor U582 (N_582,In_364,N_298);
xnor U583 (N_583,N_366,In_406);
nor U584 (N_584,In_798,In_77);
nor U585 (N_585,N_204,N_238);
or U586 (N_586,In_574,N_362);
or U587 (N_587,N_11,In_341);
or U588 (N_588,N_137,N_444);
or U589 (N_589,N_246,N_391);
nand U590 (N_590,N_240,In_740);
and U591 (N_591,N_372,N_483);
xnor U592 (N_592,N_386,N_313);
xnor U593 (N_593,N_416,In_270);
nand U594 (N_594,In_589,In_614);
nor U595 (N_595,N_66,In_864);
and U596 (N_596,N_287,In_748);
and U597 (N_597,In_140,In_900);
xor U598 (N_598,N_408,N_387);
and U599 (N_599,N_2,N_227);
nand U600 (N_600,In_450,N_507);
or U601 (N_601,In_948,In_877);
nand U602 (N_602,N_292,In_961);
xor U603 (N_603,N_527,In_182);
or U604 (N_604,N_165,N_198);
nor U605 (N_605,N_523,N_6);
xnor U606 (N_606,N_520,N_539);
or U607 (N_607,N_472,N_588);
xnor U608 (N_608,N_85,In_732);
nand U609 (N_609,N_306,N_575);
and U610 (N_610,In_761,N_460);
or U611 (N_611,In_295,N_497);
xnor U612 (N_612,N_484,In_610);
nand U613 (N_613,N_586,N_423);
or U614 (N_614,In_587,In_180);
xnor U615 (N_615,N_596,N_164);
xor U616 (N_616,N_381,N_433);
nor U617 (N_617,In_274,In_119);
nor U618 (N_618,N_54,In_437);
nor U619 (N_619,N_577,N_464);
or U620 (N_620,N_593,N_538);
and U621 (N_621,N_351,N_543);
or U622 (N_622,In_307,N_403);
or U623 (N_623,N_435,N_108);
nand U624 (N_624,N_422,N_598);
xnor U625 (N_625,In_2,N_203);
or U626 (N_626,N_324,N_245);
xor U627 (N_627,In_951,In_263);
or U628 (N_628,N_534,N_595);
nand U629 (N_629,N_265,N_513);
xor U630 (N_630,N_541,N_5);
xnor U631 (N_631,N_186,In_670);
and U632 (N_632,In_750,N_385);
nor U633 (N_633,In_543,N_263);
and U634 (N_634,In_477,N_302);
xor U635 (N_635,In_866,In_705);
xor U636 (N_636,In_113,N_556);
nor U637 (N_637,N_115,N_510);
and U638 (N_638,In_302,N_560);
and U639 (N_639,N_406,In_696);
and U640 (N_640,N_582,N_592);
xnor U641 (N_641,N_268,In_590);
or U642 (N_642,N_563,N_132);
and U643 (N_643,N_371,In_85);
xnor U644 (N_644,N_83,In_613);
xor U645 (N_645,In_441,In_387);
or U646 (N_646,N_454,N_328);
or U647 (N_647,N_441,N_436);
nor U648 (N_648,N_373,N_508);
or U649 (N_649,N_178,N_547);
nand U650 (N_650,N_544,In_146);
xnor U651 (N_651,N_80,N_153);
or U652 (N_652,N_500,N_576);
xnor U653 (N_653,In_405,N_559);
nand U654 (N_654,N_574,In_876);
nor U655 (N_655,N_174,In_983);
xor U656 (N_656,In_486,N_447);
nor U657 (N_657,N_453,In_135);
xnor U658 (N_658,N_479,N_219);
xnor U659 (N_659,N_584,N_532);
or U660 (N_660,N_516,N_32);
xor U661 (N_661,In_47,In_806);
nand U662 (N_662,In_529,In_591);
or U663 (N_663,N_476,In_31);
and U664 (N_664,N_502,N_424);
or U665 (N_665,N_320,N_551);
xor U666 (N_666,In_826,N_430);
nor U667 (N_667,N_525,N_481);
nand U668 (N_668,In_527,N_359);
xor U669 (N_669,N_55,In_809);
nand U670 (N_670,N_316,In_582);
or U671 (N_671,In_381,N_222);
nand U672 (N_672,N_121,N_369);
xor U673 (N_673,N_393,In_309);
and U674 (N_674,N_571,N_587);
nor U675 (N_675,N_154,In_571);
xor U676 (N_676,N_597,N_530);
nand U677 (N_677,N_318,N_407);
and U678 (N_678,In_354,In_720);
nand U679 (N_679,N_225,N_548);
nand U680 (N_680,N_280,In_861);
nor U681 (N_681,N_420,N_512);
nand U682 (N_682,N_583,In_494);
and U683 (N_683,N_589,N_578);
and U684 (N_684,In_753,N_144);
xor U685 (N_685,In_196,N_305);
or U686 (N_686,N_389,In_473);
xnor U687 (N_687,In_40,N_458);
nor U688 (N_688,In_746,N_554);
nor U689 (N_689,In_186,N_332);
nor U690 (N_690,N_495,In_326);
xor U691 (N_691,N_63,N_269);
nand U692 (N_692,N_522,N_199);
nor U693 (N_693,N_425,N_281);
nand U694 (N_694,In_697,N_491);
and U695 (N_695,N_489,N_405);
xor U696 (N_696,N_579,In_685);
and U697 (N_697,N_353,N_469);
nand U698 (N_698,N_395,N_537);
nor U699 (N_699,N_439,N_36);
or U700 (N_700,In_164,N_542);
nand U701 (N_701,N_637,N_24);
xor U702 (N_702,N_465,N_671);
and U703 (N_703,N_634,N_658);
xor U704 (N_704,N_485,N_664);
or U705 (N_705,In_185,In_56);
or U706 (N_706,In_572,N_648);
or U707 (N_707,N_677,N_509);
nor U708 (N_708,N_696,In_679);
or U709 (N_709,In_321,N_581);
nor U710 (N_710,N_349,N_580);
or U711 (N_711,N_501,In_601);
nor U712 (N_712,N_676,N_243);
xnor U713 (N_713,N_279,N_650);
xnor U714 (N_714,N_504,N_695);
xnor U715 (N_715,N_201,N_644);
or U716 (N_716,N_622,N_619);
nor U717 (N_717,N_660,N_565);
nor U718 (N_718,N_496,N_626);
nor U719 (N_719,N_564,N_147);
nor U720 (N_720,N_550,N_410);
nor U721 (N_721,In_883,In_430);
or U722 (N_722,N_528,N_511);
xnor U723 (N_723,N_646,N_697);
nor U724 (N_724,N_655,In_865);
xnor U725 (N_725,N_519,N_614);
nand U726 (N_726,N_682,In_747);
nor U727 (N_727,N_529,N_685);
or U728 (N_728,N_609,N_352);
nor U729 (N_729,N_535,N_606);
nand U730 (N_730,N_350,N_667);
xor U731 (N_731,N_610,N_301);
or U732 (N_732,In_109,N_630);
nand U733 (N_733,N_514,N_193);
xnor U734 (N_734,N_557,N_418);
xnor U735 (N_735,N_540,In_991);
or U736 (N_736,N_533,N_477);
xor U737 (N_737,N_638,N_536);
nor U738 (N_738,In_407,N_665);
nand U739 (N_739,In_416,N_633);
nor U740 (N_740,In_72,In_6);
xnor U741 (N_741,N_446,In_789);
and U742 (N_742,N_636,N_515);
or U743 (N_743,In_37,N_493);
and U744 (N_744,N_545,N_518);
and U745 (N_745,N_27,N_346);
or U746 (N_746,N_604,In_804);
and U747 (N_747,N_674,In_36);
and U748 (N_748,N_555,In_958);
xnor U749 (N_749,N_338,In_131);
nand U750 (N_750,N_613,N_440);
or U751 (N_751,N_615,N_384);
or U752 (N_752,N_678,In_299);
nand U753 (N_753,N_531,N_679);
nor U754 (N_754,In_497,N_663);
nor U755 (N_755,N_602,N_282);
nor U756 (N_756,N_691,N_627);
xnor U757 (N_757,In_939,N_642);
xor U758 (N_758,N_552,N_455);
and U759 (N_759,N_651,In_356);
nand U760 (N_760,N_698,N_321);
xor U761 (N_761,N_488,N_649);
xor U762 (N_762,N_478,In_780);
nand U763 (N_763,N_492,N_625);
nor U764 (N_764,N_93,In_372);
and U765 (N_765,N_694,N_681);
or U766 (N_766,N_311,N_689);
xnor U767 (N_767,N_526,N_573);
nor U768 (N_768,N_546,N_673);
xor U769 (N_769,N_659,N_639);
xor U770 (N_770,N_421,N_688);
nor U771 (N_771,N_473,In_620);
or U772 (N_772,N_498,N_146);
xor U773 (N_773,In_484,In_945);
nor U774 (N_774,N_641,In_264);
or U775 (N_775,N_635,N_629);
xor U776 (N_776,N_300,N_632);
xnor U777 (N_777,N_686,N_558);
nand U778 (N_778,In_456,N_620);
and U779 (N_779,N_623,N_585);
nand U780 (N_780,In_917,N_456);
xnor U781 (N_781,N_438,In_736);
or U782 (N_782,In_388,N_569);
xor U783 (N_783,N_631,N_669);
xor U784 (N_784,In_511,In_107);
xor U785 (N_785,N_562,N_643);
or U786 (N_786,N_640,N_189);
and U787 (N_787,N_398,N_692);
xor U788 (N_788,N_314,N_277);
xor U789 (N_789,N_616,N_394);
xnor U790 (N_790,In_285,N_590);
nand U791 (N_791,N_177,N_645);
nor U792 (N_792,In_189,N_450);
nand U793 (N_793,N_419,N_505);
and U794 (N_794,N_666,N_278);
nor U795 (N_795,N_653,N_611);
and U796 (N_796,N_471,N_374);
nand U797 (N_797,N_561,N_684);
xor U798 (N_798,N_600,N_28);
xor U799 (N_799,N_335,N_499);
and U800 (N_800,In_898,N_784);
or U801 (N_801,N_437,N_732);
or U802 (N_802,N_762,N_794);
nor U803 (N_803,In_982,N_728);
or U804 (N_804,N_782,N_722);
and U805 (N_805,N_594,N_180);
xor U806 (N_806,In_172,N_768);
and U807 (N_807,N_752,N_700);
or U808 (N_808,N_710,N_754);
and U809 (N_809,N_693,N_10);
or U810 (N_810,In_54,N_731);
nor U811 (N_811,N_781,N_755);
and U812 (N_812,N_793,N_707);
nand U813 (N_813,N_772,N_798);
nor U814 (N_814,In_150,N_687);
nand U815 (N_815,N_733,In_212);
nor U816 (N_816,N_442,N_702);
xor U817 (N_817,N_382,N_503);
nand U818 (N_818,In_710,N_743);
xor U819 (N_819,N_668,N_553);
and U820 (N_820,N_662,N_680);
nand U821 (N_821,N_757,N_717);
or U822 (N_822,N_788,N_474);
nor U823 (N_823,N_764,N_761);
or U824 (N_824,N_714,N_601);
nand U825 (N_825,N_29,N_618);
nand U826 (N_826,N_740,N_796);
or U827 (N_827,N_725,N_773);
or U828 (N_828,In_853,N_400);
nand U829 (N_829,N_480,N_736);
xnor U830 (N_830,N_739,N_672);
or U831 (N_831,N_624,N_494);
or U832 (N_832,N_724,N_566);
nor U833 (N_833,N_715,N_795);
or U834 (N_834,N_789,N_113);
nor U835 (N_835,N_683,N_799);
xnor U836 (N_836,N_767,N_621);
and U837 (N_837,N_774,N_628);
and U838 (N_838,N_744,N_171);
nand U839 (N_839,In_121,N_401);
nor U840 (N_840,In_344,N_250);
nor U841 (N_841,N_787,N_771);
xnor U842 (N_842,N_249,N_617);
nand U843 (N_843,N_699,N_711);
nand U844 (N_844,N_776,N_570);
and U845 (N_845,N_748,N_721);
xor U846 (N_846,N_261,N_413);
nand U847 (N_847,N_462,N_779);
nor U848 (N_848,N_723,N_741);
or U849 (N_849,N_517,N_482);
nand U850 (N_850,In_367,N_452);
or U851 (N_851,N_701,N_705);
nand U852 (N_852,N_652,N_612);
nor U853 (N_853,N_747,N_777);
nor U854 (N_854,N_647,N_170);
xor U855 (N_855,N_758,N_457);
and U856 (N_856,N_745,N_751);
nand U857 (N_857,N_703,N_603);
xnor U858 (N_858,In_472,N_790);
xnor U859 (N_859,N_709,N_607);
or U860 (N_860,N_770,N_354);
nor U861 (N_861,N_750,N_181);
nand U862 (N_862,In_957,N_742);
and U863 (N_863,N_749,N_737);
xor U864 (N_864,N_769,N_783);
xnor U865 (N_865,N_726,N_780);
nor U866 (N_866,In_368,N_654);
or U867 (N_867,N_756,N_706);
or U868 (N_868,N_608,In_398);
nor U869 (N_869,N_605,In_369);
or U870 (N_870,N_704,N_729);
nand U871 (N_871,N_730,N_572);
or U872 (N_872,N_44,N_657);
nor U873 (N_873,In_466,N_785);
and U874 (N_874,N_708,N_712);
and U875 (N_875,N_719,N_487);
or U876 (N_876,N_797,N_720);
nor U877 (N_877,N_713,N_330);
or U878 (N_878,N_326,N_656);
and U879 (N_879,N_734,N_412);
nand U880 (N_880,N_568,N_661);
nor U881 (N_881,N_188,N_524);
nor U882 (N_882,N_791,N_727);
xor U883 (N_883,N_591,N_746);
and U884 (N_884,N_786,N_690);
or U885 (N_885,In_327,N_670);
xnor U886 (N_886,In_519,In_926);
nand U887 (N_887,N_506,N_567);
nand U888 (N_888,N_675,N_778);
nor U889 (N_889,N_753,N_775);
xor U890 (N_890,In_202,N_735);
nand U891 (N_891,N_716,N_763);
and U892 (N_892,N_760,In_115);
or U893 (N_893,N_521,N_156);
and U894 (N_894,N_599,N_792);
and U895 (N_895,In_492,N_348);
nand U896 (N_896,N_766,In_707);
nor U897 (N_897,N_759,N_549);
and U898 (N_898,N_738,N_175);
and U899 (N_899,N_765,N_718);
or U900 (N_900,N_851,N_842);
xor U901 (N_901,N_843,N_817);
nand U902 (N_902,N_892,N_801);
nand U903 (N_903,N_897,N_857);
and U904 (N_904,N_832,N_846);
xnor U905 (N_905,N_803,N_877);
nand U906 (N_906,N_896,N_863);
and U907 (N_907,N_881,N_885);
xor U908 (N_908,N_879,N_860);
and U909 (N_909,N_878,N_893);
xor U910 (N_910,N_856,N_859);
xnor U911 (N_911,N_871,N_870);
nor U912 (N_912,N_862,N_895);
or U913 (N_913,N_814,N_808);
nand U914 (N_914,N_866,N_849);
or U915 (N_915,N_840,N_848);
and U916 (N_916,N_899,N_839);
nor U917 (N_917,N_815,N_804);
nand U918 (N_918,N_819,N_887);
and U919 (N_919,N_811,N_812);
xor U920 (N_920,N_854,N_824);
nand U921 (N_921,N_889,N_888);
nor U922 (N_922,N_872,N_821);
nor U923 (N_923,N_898,N_809);
nor U924 (N_924,N_837,N_886);
nand U925 (N_925,N_858,N_822);
nand U926 (N_926,N_813,N_835);
nand U927 (N_927,N_802,N_805);
and U928 (N_928,N_828,N_841);
nor U929 (N_929,N_867,N_836);
or U930 (N_930,N_826,N_847);
nor U931 (N_931,N_831,N_861);
and U932 (N_932,N_869,N_823);
and U933 (N_933,N_894,N_865);
and U934 (N_934,N_845,N_883);
xnor U935 (N_935,N_800,N_864);
and U936 (N_936,N_880,N_882);
or U937 (N_937,N_853,N_807);
xnor U938 (N_938,N_838,N_806);
xor U939 (N_939,N_825,N_818);
nor U940 (N_940,N_830,N_850);
xor U941 (N_941,N_820,N_868);
nor U942 (N_942,N_875,N_827);
xor U943 (N_943,N_829,N_834);
and U944 (N_944,N_873,N_874);
nor U945 (N_945,N_833,N_876);
nand U946 (N_946,N_844,N_816);
nor U947 (N_947,N_884,N_890);
or U948 (N_948,N_855,N_852);
nand U949 (N_949,N_891,N_810);
nor U950 (N_950,N_868,N_840);
and U951 (N_951,N_851,N_830);
nor U952 (N_952,N_828,N_867);
or U953 (N_953,N_848,N_853);
and U954 (N_954,N_870,N_848);
xor U955 (N_955,N_840,N_851);
nand U956 (N_956,N_897,N_852);
or U957 (N_957,N_822,N_802);
xnor U958 (N_958,N_809,N_897);
nor U959 (N_959,N_835,N_852);
nor U960 (N_960,N_887,N_812);
and U961 (N_961,N_859,N_874);
and U962 (N_962,N_854,N_858);
nor U963 (N_963,N_818,N_884);
or U964 (N_964,N_873,N_847);
and U965 (N_965,N_824,N_840);
and U966 (N_966,N_891,N_809);
xor U967 (N_967,N_819,N_849);
or U968 (N_968,N_808,N_854);
nand U969 (N_969,N_843,N_842);
nand U970 (N_970,N_852,N_867);
or U971 (N_971,N_808,N_841);
nand U972 (N_972,N_860,N_822);
xor U973 (N_973,N_867,N_830);
and U974 (N_974,N_897,N_827);
and U975 (N_975,N_826,N_855);
or U976 (N_976,N_848,N_847);
xor U977 (N_977,N_893,N_872);
or U978 (N_978,N_884,N_847);
and U979 (N_979,N_871,N_812);
nand U980 (N_980,N_808,N_820);
xnor U981 (N_981,N_857,N_891);
nor U982 (N_982,N_875,N_807);
and U983 (N_983,N_872,N_858);
and U984 (N_984,N_895,N_815);
and U985 (N_985,N_899,N_894);
xnor U986 (N_986,N_832,N_859);
and U987 (N_987,N_826,N_823);
nand U988 (N_988,N_885,N_820);
nand U989 (N_989,N_889,N_817);
or U990 (N_990,N_883,N_881);
xor U991 (N_991,N_875,N_825);
nor U992 (N_992,N_883,N_880);
and U993 (N_993,N_885,N_836);
or U994 (N_994,N_837,N_860);
or U995 (N_995,N_837,N_826);
or U996 (N_996,N_855,N_839);
or U997 (N_997,N_810,N_829);
xor U998 (N_998,N_807,N_899);
and U999 (N_999,N_815,N_820);
and U1000 (N_1000,N_949,N_904);
nor U1001 (N_1001,N_979,N_958);
and U1002 (N_1002,N_971,N_951);
and U1003 (N_1003,N_961,N_959);
nor U1004 (N_1004,N_974,N_999);
nand U1005 (N_1005,N_977,N_942);
nand U1006 (N_1006,N_947,N_980);
xnor U1007 (N_1007,N_931,N_950);
nand U1008 (N_1008,N_903,N_948);
nand U1009 (N_1009,N_927,N_969);
nand U1010 (N_1010,N_986,N_917);
nand U1011 (N_1011,N_905,N_989);
and U1012 (N_1012,N_993,N_988);
nor U1013 (N_1013,N_900,N_910);
or U1014 (N_1014,N_992,N_919);
nor U1015 (N_1015,N_929,N_975);
or U1016 (N_1016,N_956,N_946);
nand U1017 (N_1017,N_998,N_906);
nand U1018 (N_1018,N_916,N_907);
or U1019 (N_1019,N_920,N_963);
and U1020 (N_1020,N_918,N_960);
xor U1021 (N_1021,N_926,N_945);
nand U1022 (N_1022,N_972,N_911);
nor U1023 (N_1023,N_994,N_964);
or U1024 (N_1024,N_968,N_913);
nand U1025 (N_1025,N_982,N_928);
or U1026 (N_1026,N_921,N_965);
nor U1027 (N_1027,N_933,N_941);
xor U1028 (N_1028,N_944,N_955);
nor U1029 (N_1029,N_991,N_909);
nor U1030 (N_1030,N_970,N_962);
or U1031 (N_1031,N_935,N_936);
nor U1032 (N_1032,N_981,N_908);
or U1033 (N_1033,N_966,N_983);
nand U1034 (N_1034,N_990,N_924);
xnor U1035 (N_1035,N_987,N_967);
xor U1036 (N_1036,N_934,N_976);
xnor U1037 (N_1037,N_997,N_925);
nor U1038 (N_1038,N_938,N_978);
or U1039 (N_1039,N_902,N_923);
xor U1040 (N_1040,N_940,N_995);
or U1041 (N_1041,N_939,N_937);
and U1042 (N_1042,N_973,N_930);
and U1043 (N_1043,N_932,N_901);
or U1044 (N_1044,N_954,N_915);
and U1045 (N_1045,N_953,N_922);
nand U1046 (N_1046,N_957,N_943);
xor U1047 (N_1047,N_984,N_952);
nand U1048 (N_1048,N_912,N_996);
and U1049 (N_1049,N_914,N_985);
xor U1050 (N_1050,N_914,N_945);
xor U1051 (N_1051,N_937,N_938);
and U1052 (N_1052,N_970,N_930);
nand U1053 (N_1053,N_949,N_970);
nand U1054 (N_1054,N_951,N_902);
nor U1055 (N_1055,N_968,N_962);
and U1056 (N_1056,N_919,N_994);
and U1057 (N_1057,N_970,N_956);
or U1058 (N_1058,N_943,N_951);
nand U1059 (N_1059,N_943,N_928);
or U1060 (N_1060,N_977,N_901);
and U1061 (N_1061,N_961,N_983);
nor U1062 (N_1062,N_973,N_962);
and U1063 (N_1063,N_956,N_940);
and U1064 (N_1064,N_957,N_942);
and U1065 (N_1065,N_942,N_936);
nor U1066 (N_1066,N_909,N_982);
nor U1067 (N_1067,N_954,N_923);
nand U1068 (N_1068,N_939,N_907);
and U1069 (N_1069,N_923,N_979);
nor U1070 (N_1070,N_997,N_915);
xor U1071 (N_1071,N_962,N_948);
nand U1072 (N_1072,N_972,N_903);
and U1073 (N_1073,N_934,N_963);
xor U1074 (N_1074,N_971,N_913);
xnor U1075 (N_1075,N_926,N_954);
xnor U1076 (N_1076,N_953,N_955);
nor U1077 (N_1077,N_907,N_904);
nand U1078 (N_1078,N_926,N_942);
or U1079 (N_1079,N_935,N_906);
xnor U1080 (N_1080,N_951,N_928);
or U1081 (N_1081,N_910,N_950);
or U1082 (N_1082,N_969,N_977);
nor U1083 (N_1083,N_913,N_922);
nand U1084 (N_1084,N_921,N_908);
and U1085 (N_1085,N_953,N_931);
or U1086 (N_1086,N_913,N_955);
nor U1087 (N_1087,N_994,N_951);
and U1088 (N_1088,N_901,N_964);
xnor U1089 (N_1089,N_903,N_915);
or U1090 (N_1090,N_950,N_926);
or U1091 (N_1091,N_959,N_941);
nor U1092 (N_1092,N_958,N_915);
and U1093 (N_1093,N_947,N_995);
and U1094 (N_1094,N_905,N_935);
nor U1095 (N_1095,N_956,N_988);
xor U1096 (N_1096,N_944,N_961);
and U1097 (N_1097,N_979,N_924);
or U1098 (N_1098,N_984,N_974);
xor U1099 (N_1099,N_923,N_958);
nor U1100 (N_1100,N_1095,N_1031);
nor U1101 (N_1101,N_1010,N_1092);
nor U1102 (N_1102,N_1057,N_1078);
or U1103 (N_1103,N_1071,N_1087);
or U1104 (N_1104,N_1015,N_1068);
or U1105 (N_1105,N_1086,N_1016);
xnor U1106 (N_1106,N_1050,N_1021);
nor U1107 (N_1107,N_1012,N_1089);
nor U1108 (N_1108,N_1045,N_1077);
nor U1109 (N_1109,N_1048,N_1017);
nand U1110 (N_1110,N_1080,N_1065);
nor U1111 (N_1111,N_1076,N_1070);
nor U1112 (N_1112,N_1083,N_1096);
and U1113 (N_1113,N_1001,N_1082);
and U1114 (N_1114,N_1099,N_1066);
and U1115 (N_1115,N_1052,N_1014);
nor U1116 (N_1116,N_1011,N_1049);
nand U1117 (N_1117,N_1022,N_1008);
nor U1118 (N_1118,N_1039,N_1094);
xnor U1119 (N_1119,N_1032,N_1058);
and U1120 (N_1120,N_1030,N_1042);
or U1121 (N_1121,N_1046,N_1055);
nor U1122 (N_1122,N_1038,N_1003);
nor U1123 (N_1123,N_1067,N_1059);
nand U1124 (N_1124,N_1097,N_1025);
nand U1125 (N_1125,N_1007,N_1043);
xor U1126 (N_1126,N_1036,N_1023);
xnor U1127 (N_1127,N_1020,N_1081);
or U1128 (N_1128,N_1024,N_1053);
xor U1129 (N_1129,N_1013,N_1074);
nor U1130 (N_1130,N_1027,N_1028);
and U1131 (N_1131,N_1093,N_1075);
and U1132 (N_1132,N_1054,N_1079);
nand U1133 (N_1133,N_1051,N_1091);
nor U1134 (N_1134,N_1061,N_1063);
nor U1135 (N_1135,N_1073,N_1018);
xor U1136 (N_1136,N_1069,N_1035);
and U1137 (N_1137,N_1002,N_1009);
and U1138 (N_1138,N_1004,N_1019);
nor U1139 (N_1139,N_1072,N_1041);
or U1140 (N_1140,N_1084,N_1085);
and U1141 (N_1141,N_1064,N_1000);
xor U1142 (N_1142,N_1098,N_1029);
or U1143 (N_1143,N_1040,N_1026);
nand U1144 (N_1144,N_1056,N_1090);
or U1145 (N_1145,N_1033,N_1005);
or U1146 (N_1146,N_1037,N_1062);
and U1147 (N_1147,N_1047,N_1034);
and U1148 (N_1148,N_1088,N_1060);
nor U1149 (N_1149,N_1006,N_1044);
xnor U1150 (N_1150,N_1094,N_1031);
nand U1151 (N_1151,N_1078,N_1023);
and U1152 (N_1152,N_1099,N_1060);
or U1153 (N_1153,N_1008,N_1029);
xor U1154 (N_1154,N_1059,N_1077);
nand U1155 (N_1155,N_1052,N_1051);
nand U1156 (N_1156,N_1015,N_1076);
xor U1157 (N_1157,N_1033,N_1016);
nand U1158 (N_1158,N_1030,N_1097);
or U1159 (N_1159,N_1028,N_1039);
and U1160 (N_1160,N_1078,N_1058);
nand U1161 (N_1161,N_1019,N_1002);
nor U1162 (N_1162,N_1048,N_1001);
or U1163 (N_1163,N_1010,N_1043);
xnor U1164 (N_1164,N_1070,N_1039);
and U1165 (N_1165,N_1070,N_1042);
nand U1166 (N_1166,N_1026,N_1052);
and U1167 (N_1167,N_1028,N_1012);
or U1168 (N_1168,N_1019,N_1046);
xnor U1169 (N_1169,N_1040,N_1057);
nand U1170 (N_1170,N_1031,N_1044);
nor U1171 (N_1171,N_1012,N_1088);
nand U1172 (N_1172,N_1055,N_1031);
xnor U1173 (N_1173,N_1061,N_1007);
xor U1174 (N_1174,N_1073,N_1094);
and U1175 (N_1175,N_1023,N_1048);
xor U1176 (N_1176,N_1097,N_1033);
nor U1177 (N_1177,N_1089,N_1018);
xnor U1178 (N_1178,N_1026,N_1081);
xnor U1179 (N_1179,N_1071,N_1048);
and U1180 (N_1180,N_1065,N_1031);
nor U1181 (N_1181,N_1093,N_1028);
or U1182 (N_1182,N_1024,N_1095);
nor U1183 (N_1183,N_1085,N_1063);
nor U1184 (N_1184,N_1065,N_1014);
nand U1185 (N_1185,N_1022,N_1032);
xor U1186 (N_1186,N_1011,N_1024);
and U1187 (N_1187,N_1016,N_1010);
nor U1188 (N_1188,N_1074,N_1068);
nor U1189 (N_1189,N_1070,N_1086);
and U1190 (N_1190,N_1003,N_1068);
and U1191 (N_1191,N_1038,N_1052);
and U1192 (N_1192,N_1030,N_1017);
nor U1193 (N_1193,N_1039,N_1072);
nor U1194 (N_1194,N_1036,N_1062);
and U1195 (N_1195,N_1038,N_1049);
nor U1196 (N_1196,N_1057,N_1056);
nor U1197 (N_1197,N_1037,N_1014);
nor U1198 (N_1198,N_1092,N_1050);
nor U1199 (N_1199,N_1097,N_1003);
and U1200 (N_1200,N_1169,N_1111);
and U1201 (N_1201,N_1132,N_1130);
and U1202 (N_1202,N_1112,N_1160);
nand U1203 (N_1203,N_1171,N_1143);
or U1204 (N_1204,N_1176,N_1159);
and U1205 (N_1205,N_1128,N_1134);
and U1206 (N_1206,N_1166,N_1153);
xor U1207 (N_1207,N_1102,N_1149);
nor U1208 (N_1208,N_1126,N_1145);
and U1209 (N_1209,N_1100,N_1189);
or U1210 (N_1210,N_1154,N_1165);
nor U1211 (N_1211,N_1155,N_1148);
xnor U1212 (N_1212,N_1182,N_1170);
nor U1213 (N_1213,N_1192,N_1172);
nor U1214 (N_1214,N_1174,N_1163);
and U1215 (N_1215,N_1103,N_1115);
or U1216 (N_1216,N_1152,N_1181);
or U1217 (N_1217,N_1198,N_1119);
nor U1218 (N_1218,N_1183,N_1196);
or U1219 (N_1219,N_1121,N_1157);
or U1220 (N_1220,N_1187,N_1197);
and U1221 (N_1221,N_1193,N_1168);
or U1222 (N_1222,N_1151,N_1150);
xor U1223 (N_1223,N_1129,N_1188);
nor U1224 (N_1224,N_1120,N_1108);
xnor U1225 (N_1225,N_1156,N_1118);
xor U1226 (N_1226,N_1180,N_1135);
nand U1227 (N_1227,N_1141,N_1139);
or U1228 (N_1228,N_1127,N_1158);
and U1229 (N_1229,N_1113,N_1179);
nor U1230 (N_1230,N_1186,N_1125);
nand U1231 (N_1231,N_1164,N_1194);
nor U1232 (N_1232,N_1137,N_1124);
nor U1233 (N_1233,N_1147,N_1140);
nand U1234 (N_1234,N_1178,N_1195);
nor U1235 (N_1235,N_1131,N_1185);
or U1236 (N_1236,N_1101,N_1106);
and U1237 (N_1237,N_1142,N_1146);
nand U1238 (N_1238,N_1175,N_1136);
nor U1239 (N_1239,N_1123,N_1167);
nand U1240 (N_1240,N_1122,N_1133);
and U1241 (N_1241,N_1144,N_1114);
nand U1242 (N_1242,N_1107,N_1161);
nand U1243 (N_1243,N_1109,N_1191);
xnor U1244 (N_1244,N_1138,N_1116);
nand U1245 (N_1245,N_1199,N_1117);
nand U1246 (N_1246,N_1104,N_1105);
nor U1247 (N_1247,N_1173,N_1190);
nand U1248 (N_1248,N_1184,N_1110);
nor U1249 (N_1249,N_1177,N_1162);
nor U1250 (N_1250,N_1150,N_1146);
nor U1251 (N_1251,N_1188,N_1134);
nand U1252 (N_1252,N_1172,N_1193);
or U1253 (N_1253,N_1117,N_1113);
and U1254 (N_1254,N_1191,N_1190);
nand U1255 (N_1255,N_1160,N_1116);
xnor U1256 (N_1256,N_1173,N_1193);
xor U1257 (N_1257,N_1118,N_1123);
or U1258 (N_1258,N_1147,N_1110);
or U1259 (N_1259,N_1168,N_1155);
and U1260 (N_1260,N_1192,N_1104);
and U1261 (N_1261,N_1128,N_1153);
or U1262 (N_1262,N_1110,N_1173);
or U1263 (N_1263,N_1128,N_1152);
nand U1264 (N_1264,N_1111,N_1145);
xor U1265 (N_1265,N_1129,N_1106);
xnor U1266 (N_1266,N_1148,N_1178);
nand U1267 (N_1267,N_1183,N_1144);
nor U1268 (N_1268,N_1105,N_1122);
or U1269 (N_1269,N_1124,N_1167);
nand U1270 (N_1270,N_1171,N_1187);
nand U1271 (N_1271,N_1180,N_1111);
nor U1272 (N_1272,N_1127,N_1136);
or U1273 (N_1273,N_1145,N_1162);
or U1274 (N_1274,N_1133,N_1168);
and U1275 (N_1275,N_1175,N_1139);
xor U1276 (N_1276,N_1124,N_1190);
nand U1277 (N_1277,N_1198,N_1190);
nand U1278 (N_1278,N_1191,N_1170);
or U1279 (N_1279,N_1191,N_1188);
xor U1280 (N_1280,N_1131,N_1111);
nand U1281 (N_1281,N_1194,N_1156);
or U1282 (N_1282,N_1192,N_1135);
nor U1283 (N_1283,N_1159,N_1144);
and U1284 (N_1284,N_1161,N_1193);
or U1285 (N_1285,N_1132,N_1160);
nand U1286 (N_1286,N_1183,N_1133);
nand U1287 (N_1287,N_1100,N_1180);
or U1288 (N_1288,N_1178,N_1101);
and U1289 (N_1289,N_1152,N_1133);
xor U1290 (N_1290,N_1161,N_1134);
or U1291 (N_1291,N_1145,N_1120);
nand U1292 (N_1292,N_1132,N_1148);
nand U1293 (N_1293,N_1108,N_1199);
or U1294 (N_1294,N_1175,N_1119);
nand U1295 (N_1295,N_1125,N_1179);
xor U1296 (N_1296,N_1190,N_1123);
nand U1297 (N_1297,N_1171,N_1144);
or U1298 (N_1298,N_1187,N_1169);
nor U1299 (N_1299,N_1130,N_1131);
nor U1300 (N_1300,N_1246,N_1256);
and U1301 (N_1301,N_1299,N_1251);
xor U1302 (N_1302,N_1286,N_1247);
nand U1303 (N_1303,N_1273,N_1260);
or U1304 (N_1304,N_1232,N_1224);
nor U1305 (N_1305,N_1205,N_1230);
xor U1306 (N_1306,N_1211,N_1234);
nor U1307 (N_1307,N_1225,N_1278);
or U1308 (N_1308,N_1279,N_1239);
xnor U1309 (N_1309,N_1258,N_1214);
xor U1310 (N_1310,N_1261,N_1271);
or U1311 (N_1311,N_1235,N_1281);
nor U1312 (N_1312,N_1298,N_1257);
nor U1313 (N_1313,N_1226,N_1242);
and U1314 (N_1314,N_1275,N_1292);
nor U1315 (N_1315,N_1266,N_1289);
nor U1316 (N_1316,N_1253,N_1296);
xor U1317 (N_1317,N_1215,N_1243);
xor U1318 (N_1318,N_1297,N_1203);
xor U1319 (N_1319,N_1227,N_1216);
xor U1320 (N_1320,N_1213,N_1240);
or U1321 (N_1321,N_1245,N_1284);
and U1322 (N_1322,N_1268,N_1290);
nand U1323 (N_1323,N_1208,N_1221);
xor U1324 (N_1324,N_1233,N_1294);
nand U1325 (N_1325,N_1237,N_1200);
or U1326 (N_1326,N_1272,N_1217);
or U1327 (N_1327,N_1228,N_1291);
xor U1328 (N_1328,N_1274,N_1295);
nor U1329 (N_1329,N_1250,N_1259);
nand U1330 (N_1330,N_1201,N_1285);
nor U1331 (N_1331,N_1264,N_1223);
nor U1332 (N_1332,N_1276,N_1222);
nand U1333 (N_1333,N_1229,N_1207);
xnor U1334 (N_1334,N_1288,N_1219);
nand U1335 (N_1335,N_1293,N_1204);
nor U1336 (N_1336,N_1249,N_1282);
or U1337 (N_1337,N_1287,N_1248);
nor U1338 (N_1338,N_1267,N_1236);
xor U1339 (N_1339,N_1220,N_1209);
xnor U1340 (N_1340,N_1202,N_1277);
or U1341 (N_1341,N_1238,N_1269);
and U1342 (N_1342,N_1255,N_1270);
nor U1343 (N_1343,N_1263,N_1231);
or U1344 (N_1344,N_1210,N_1265);
or U1345 (N_1345,N_1241,N_1206);
nor U1346 (N_1346,N_1254,N_1218);
nand U1347 (N_1347,N_1280,N_1283);
nand U1348 (N_1348,N_1212,N_1262);
nor U1349 (N_1349,N_1244,N_1252);
and U1350 (N_1350,N_1239,N_1206);
xnor U1351 (N_1351,N_1265,N_1285);
xor U1352 (N_1352,N_1224,N_1297);
nand U1353 (N_1353,N_1221,N_1231);
nor U1354 (N_1354,N_1278,N_1237);
nor U1355 (N_1355,N_1295,N_1293);
xnor U1356 (N_1356,N_1202,N_1266);
and U1357 (N_1357,N_1274,N_1215);
nand U1358 (N_1358,N_1208,N_1295);
or U1359 (N_1359,N_1250,N_1211);
and U1360 (N_1360,N_1206,N_1282);
and U1361 (N_1361,N_1251,N_1279);
xnor U1362 (N_1362,N_1242,N_1267);
nand U1363 (N_1363,N_1244,N_1263);
nand U1364 (N_1364,N_1209,N_1244);
nand U1365 (N_1365,N_1263,N_1276);
and U1366 (N_1366,N_1232,N_1264);
nand U1367 (N_1367,N_1274,N_1269);
and U1368 (N_1368,N_1257,N_1210);
xor U1369 (N_1369,N_1238,N_1251);
nand U1370 (N_1370,N_1238,N_1208);
nand U1371 (N_1371,N_1252,N_1207);
nand U1372 (N_1372,N_1232,N_1286);
nand U1373 (N_1373,N_1218,N_1298);
xnor U1374 (N_1374,N_1235,N_1256);
and U1375 (N_1375,N_1239,N_1221);
nor U1376 (N_1376,N_1252,N_1276);
xnor U1377 (N_1377,N_1249,N_1295);
or U1378 (N_1378,N_1226,N_1200);
or U1379 (N_1379,N_1221,N_1218);
nor U1380 (N_1380,N_1253,N_1244);
and U1381 (N_1381,N_1299,N_1233);
nor U1382 (N_1382,N_1278,N_1245);
or U1383 (N_1383,N_1246,N_1290);
and U1384 (N_1384,N_1207,N_1239);
nor U1385 (N_1385,N_1202,N_1207);
nand U1386 (N_1386,N_1290,N_1261);
nand U1387 (N_1387,N_1285,N_1247);
or U1388 (N_1388,N_1236,N_1289);
or U1389 (N_1389,N_1262,N_1228);
xor U1390 (N_1390,N_1287,N_1256);
nor U1391 (N_1391,N_1284,N_1286);
or U1392 (N_1392,N_1282,N_1233);
xor U1393 (N_1393,N_1246,N_1241);
nor U1394 (N_1394,N_1282,N_1271);
and U1395 (N_1395,N_1236,N_1217);
and U1396 (N_1396,N_1275,N_1229);
or U1397 (N_1397,N_1253,N_1236);
nand U1398 (N_1398,N_1249,N_1220);
xnor U1399 (N_1399,N_1261,N_1232);
xnor U1400 (N_1400,N_1341,N_1369);
and U1401 (N_1401,N_1330,N_1360);
nand U1402 (N_1402,N_1326,N_1317);
or U1403 (N_1403,N_1352,N_1331);
nand U1404 (N_1404,N_1374,N_1332);
nand U1405 (N_1405,N_1398,N_1371);
nor U1406 (N_1406,N_1388,N_1380);
and U1407 (N_1407,N_1372,N_1324);
nor U1408 (N_1408,N_1322,N_1311);
or U1409 (N_1409,N_1384,N_1382);
and U1410 (N_1410,N_1399,N_1368);
nand U1411 (N_1411,N_1329,N_1370);
nor U1412 (N_1412,N_1357,N_1385);
and U1413 (N_1413,N_1347,N_1363);
and U1414 (N_1414,N_1361,N_1336);
nand U1415 (N_1415,N_1390,N_1378);
xnor U1416 (N_1416,N_1349,N_1320);
nand U1417 (N_1417,N_1309,N_1327);
and U1418 (N_1418,N_1387,N_1393);
nand U1419 (N_1419,N_1337,N_1379);
and U1420 (N_1420,N_1306,N_1328);
nor U1421 (N_1421,N_1315,N_1373);
and U1422 (N_1422,N_1386,N_1300);
or U1423 (N_1423,N_1367,N_1321);
nor U1424 (N_1424,N_1344,N_1362);
or U1425 (N_1425,N_1354,N_1343);
or U1426 (N_1426,N_1376,N_1308);
nor U1427 (N_1427,N_1377,N_1314);
and U1428 (N_1428,N_1391,N_1323);
nand U1429 (N_1429,N_1350,N_1364);
nand U1430 (N_1430,N_1395,N_1383);
and U1431 (N_1431,N_1304,N_1339);
and U1432 (N_1432,N_1358,N_1303);
nor U1433 (N_1433,N_1353,N_1365);
xnor U1434 (N_1434,N_1338,N_1397);
or U1435 (N_1435,N_1325,N_1316);
xor U1436 (N_1436,N_1381,N_1312);
and U1437 (N_1437,N_1318,N_1319);
nand U1438 (N_1438,N_1334,N_1356);
or U1439 (N_1439,N_1333,N_1340);
nand U1440 (N_1440,N_1375,N_1392);
nand U1441 (N_1441,N_1313,N_1342);
or U1442 (N_1442,N_1307,N_1351);
xor U1443 (N_1443,N_1301,N_1394);
or U1444 (N_1444,N_1305,N_1302);
nor U1445 (N_1445,N_1345,N_1355);
xnor U1446 (N_1446,N_1389,N_1359);
xnor U1447 (N_1447,N_1346,N_1310);
and U1448 (N_1448,N_1366,N_1396);
or U1449 (N_1449,N_1348,N_1335);
nor U1450 (N_1450,N_1352,N_1356);
xnor U1451 (N_1451,N_1319,N_1355);
xor U1452 (N_1452,N_1362,N_1374);
nand U1453 (N_1453,N_1389,N_1357);
and U1454 (N_1454,N_1332,N_1336);
nand U1455 (N_1455,N_1388,N_1362);
nor U1456 (N_1456,N_1395,N_1390);
or U1457 (N_1457,N_1310,N_1343);
xor U1458 (N_1458,N_1359,N_1385);
or U1459 (N_1459,N_1386,N_1362);
nor U1460 (N_1460,N_1322,N_1353);
and U1461 (N_1461,N_1353,N_1370);
and U1462 (N_1462,N_1309,N_1393);
and U1463 (N_1463,N_1378,N_1381);
nand U1464 (N_1464,N_1337,N_1383);
and U1465 (N_1465,N_1369,N_1385);
or U1466 (N_1466,N_1346,N_1354);
nand U1467 (N_1467,N_1385,N_1334);
xnor U1468 (N_1468,N_1366,N_1372);
and U1469 (N_1469,N_1399,N_1371);
nor U1470 (N_1470,N_1322,N_1375);
and U1471 (N_1471,N_1339,N_1307);
and U1472 (N_1472,N_1344,N_1349);
xnor U1473 (N_1473,N_1358,N_1388);
nand U1474 (N_1474,N_1336,N_1368);
nand U1475 (N_1475,N_1361,N_1376);
and U1476 (N_1476,N_1394,N_1326);
nand U1477 (N_1477,N_1383,N_1379);
nor U1478 (N_1478,N_1355,N_1399);
nor U1479 (N_1479,N_1392,N_1333);
xnor U1480 (N_1480,N_1308,N_1398);
nand U1481 (N_1481,N_1399,N_1377);
nor U1482 (N_1482,N_1330,N_1318);
nor U1483 (N_1483,N_1375,N_1311);
and U1484 (N_1484,N_1359,N_1325);
and U1485 (N_1485,N_1381,N_1333);
nand U1486 (N_1486,N_1387,N_1334);
nand U1487 (N_1487,N_1343,N_1345);
nand U1488 (N_1488,N_1371,N_1338);
or U1489 (N_1489,N_1346,N_1320);
or U1490 (N_1490,N_1354,N_1370);
and U1491 (N_1491,N_1315,N_1344);
or U1492 (N_1492,N_1328,N_1314);
or U1493 (N_1493,N_1350,N_1392);
or U1494 (N_1494,N_1395,N_1310);
or U1495 (N_1495,N_1395,N_1399);
and U1496 (N_1496,N_1398,N_1315);
or U1497 (N_1497,N_1310,N_1326);
or U1498 (N_1498,N_1320,N_1326);
and U1499 (N_1499,N_1325,N_1369);
and U1500 (N_1500,N_1454,N_1430);
nor U1501 (N_1501,N_1492,N_1402);
or U1502 (N_1502,N_1470,N_1477);
or U1503 (N_1503,N_1417,N_1429);
or U1504 (N_1504,N_1458,N_1446);
and U1505 (N_1505,N_1411,N_1447);
xor U1506 (N_1506,N_1467,N_1490);
nor U1507 (N_1507,N_1401,N_1440);
nor U1508 (N_1508,N_1413,N_1474);
nand U1509 (N_1509,N_1443,N_1442);
nand U1510 (N_1510,N_1487,N_1419);
and U1511 (N_1511,N_1416,N_1426);
and U1512 (N_1512,N_1455,N_1475);
xnor U1513 (N_1513,N_1476,N_1462);
or U1514 (N_1514,N_1421,N_1439);
xor U1515 (N_1515,N_1479,N_1434);
nand U1516 (N_1516,N_1445,N_1465);
and U1517 (N_1517,N_1423,N_1472);
nand U1518 (N_1518,N_1485,N_1456);
or U1519 (N_1519,N_1463,N_1457);
nor U1520 (N_1520,N_1420,N_1450);
and U1521 (N_1521,N_1433,N_1405);
and U1522 (N_1522,N_1441,N_1486);
nand U1523 (N_1523,N_1469,N_1495);
or U1524 (N_1524,N_1428,N_1412);
nor U1525 (N_1525,N_1491,N_1400);
and U1526 (N_1526,N_1482,N_1488);
and U1527 (N_1527,N_1466,N_1478);
nand U1528 (N_1528,N_1494,N_1493);
or U1529 (N_1529,N_1408,N_1415);
and U1530 (N_1530,N_1452,N_1448);
nor U1531 (N_1531,N_1407,N_1438);
and U1532 (N_1532,N_1459,N_1435);
nand U1533 (N_1533,N_1414,N_1461);
or U1534 (N_1534,N_1409,N_1444);
and U1535 (N_1535,N_1431,N_1483);
nand U1536 (N_1536,N_1424,N_1453);
xnor U1537 (N_1537,N_1451,N_1471);
and U1538 (N_1538,N_1427,N_1497);
or U1539 (N_1539,N_1425,N_1432);
xor U1540 (N_1540,N_1473,N_1404);
nand U1541 (N_1541,N_1481,N_1496);
nand U1542 (N_1542,N_1484,N_1480);
or U1543 (N_1543,N_1422,N_1464);
xnor U1544 (N_1544,N_1410,N_1460);
xor U1545 (N_1545,N_1437,N_1449);
nor U1546 (N_1546,N_1403,N_1418);
nand U1547 (N_1547,N_1489,N_1406);
nor U1548 (N_1548,N_1498,N_1436);
nand U1549 (N_1549,N_1499,N_1468);
or U1550 (N_1550,N_1473,N_1412);
nand U1551 (N_1551,N_1417,N_1494);
nor U1552 (N_1552,N_1434,N_1416);
nand U1553 (N_1553,N_1426,N_1417);
or U1554 (N_1554,N_1473,N_1441);
xnor U1555 (N_1555,N_1478,N_1406);
xor U1556 (N_1556,N_1422,N_1468);
or U1557 (N_1557,N_1403,N_1480);
and U1558 (N_1558,N_1452,N_1474);
nand U1559 (N_1559,N_1429,N_1423);
xor U1560 (N_1560,N_1405,N_1461);
xor U1561 (N_1561,N_1457,N_1472);
xor U1562 (N_1562,N_1444,N_1439);
nor U1563 (N_1563,N_1429,N_1483);
xnor U1564 (N_1564,N_1412,N_1457);
or U1565 (N_1565,N_1447,N_1438);
and U1566 (N_1566,N_1464,N_1491);
xor U1567 (N_1567,N_1490,N_1493);
nand U1568 (N_1568,N_1453,N_1451);
and U1569 (N_1569,N_1419,N_1481);
and U1570 (N_1570,N_1448,N_1412);
or U1571 (N_1571,N_1400,N_1412);
or U1572 (N_1572,N_1437,N_1446);
or U1573 (N_1573,N_1422,N_1411);
and U1574 (N_1574,N_1422,N_1465);
nor U1575 (N_1575,N_1425,N_1440);
xor U1576 (N_1576,N_1445,N_1409);
xnor U1577 (N_1577,N_1491,N_1441);
xnor U1578 (N_1578,N_1439,N_1456);
xnor U1579 (N_1579,N_1469,N_1476);
and U1580 (N_1580,N_1438,N_1414);
xnor U1581 (N_1581,N_1461,N_1403);
nor U1582 (N_1582,N_1427,N_1478);
nand U1583 (N_1583,N_1460,N_1417);
nor U1584 (N_1584,N_1490,N_1486);
or U1585 (N_1585,N_1447,N_1431);
or U1586 (N_1586,N_1413,N_1449);
nand U1587 (N_1587,N_1426,N_1439);
nand U1588 (N_1588,N_1489,N_1460);
nand U1589 (N_1589,N_1424,N_1470);
or U1590 (N_1590,N_1427,N_1460);
nand U1591 (N_1591,N_1463,N_1411);
xor U1592 (N_1592,N_1438,N_1412);
xnor U1593 (N_1593,N_1477,N_1493);
nor U1594 (N_1594,N_1484,N_1458);
or U1595 (N_1595,N_1475,N_1417);
nand U1596 (N_1596,N_1453,N_1403);
nand U1597 (N_1597,N_1460,N_1444);
or U1598 (N_1598,N_1403,N_1483);
nor U1599 (N_1599,N_1420,N_1438);
xnor U1600 (N_1600,N_1518,N_1515);
nand U1601 (N_1601,N_1564,N_1556);
nand U1602 (N_1602,N_1568,N_1533);
or U1603 (N_1603,N_1592,N_1598);
nand U1604 (N_1604,N_1576,N_1546);
or U1605 (N_1605,N_1561,N_1593);
nor U1606 (N_1606,N_1560,N_1509);
nor U1607 (N_1607,N_1532,N_1535);
xnor U1608 (N_1608,N_1545,N_1500);
nand U1609 (N_1609,N_1544,N_1536);
or U1610 (N_1610,N_1505,N_1577);
nand U1611 (N_1611,N_1552,N_1534);
xor U1612 (N_1612,N_1583,N_1559);
nand U1613 (N_1613,N_1585,N_1588);
xor U1614 (N_1614,N_1538,N_1589);
xor U1615 (N_1615,N_1525,N_1595);
nand U1616 (N_1616,N_1516,N_1597);
and U1617 (N_1617,N_1530,N_1562);
nand U1618 (N_1618,N_1529,N_1548);
or U1619 (N_1619,N_1501,N_1506);
and U1620 (N_1620,N_1537,N_1541);
and U1621 (N_1621,N_1521,N_1514);
nor U1622 (N_1622,N_1555,N_1539);
nor U1623 (N_1623,N_1566,N_1550);
nor U1624 (N_1624,N_1526,N_1519);
xnor U1625 (N_1625,N_1591,N_1586);
nand U1626 (N_1626,N_1596,N_1503);
or U1627 (N_1627,N_1573,N_1565);
xor U1628 (N_1628,N_1512,N_1553);
nor U1629 (N_1629,N_1524,N_1581);
nor U1630 (N_1630,N_1563,N_1574);
nand U1631 (N_1631,N_1557,N_1547);
xor U1632 (N_1632,N_1502,N_1549);
nor U1633 (N_1633,N_1504,N_1554);
xnor U1634 (N_1634,N_1531,N_1522);
xor U1635 (N_1635,N_1579,N_1508);
nand U1636 (N_1636,N_1594,N_1572);
or U1637 (N_1637,N_1567,N_1527);
and U1638 (N_1638,N_1575,N_1520);
nand U1639 (N_1639,N_1590,N_1551);
nand U1640 (N_1640,N_1569,N_1511);
nor U1641 (N_1641,N_1543,N_1542);
and U1642 (N_1642,N_1599,N_1571);
and U1643 (N_1643,N_1582,N_1513);
xor U1644 (N_1644,N_1540,N_1578);
nor U1645 (N_1645,N_1517,N_1580);
nand U1646 (N_1646,N_1570,N_1523);
and U1647 (N_1647,N_1584,N_1587);
xnor U1648 (N_1648,N_1510,N_1507);
nor U1649 (N_1649,N_1528,N_1558);
xnor U1650 (N_1650,N_1597,N_1581);
or U1651 (N_1651,N_1528,N_1500);
nor U1652 (N_1652,N_1509,N_1506);
nand U1653 (N_1653,N_1550,N_1535);
xor U1654 (N_1654,N_1535,N_1522);
nor U1655 (N_1655,N_1537,N_1558);
nor U1656 (N_1656,N_1513,N_1567);
nor U1657 (N_1657,N_1510,N_1572);
and U1658 (N_1658,N_1564,N_1565);
and U1659 (N_1659,N_1506,N_1587);
or U1660 (N_1660,N_1541,N_1529);
nor U1661 (N_1661,N_1577,N_1527);
xor U1662 (N_1662,N_1514,N_1575);
xnor U1663 (N_1663,N_1569,N_1503);
and U1664 (N_1664,N_1513,N_1598);
and U1665 (N_1665,N_1531,N_1588);
nand U1666 (N_1666,N_1523,N_1567);
xor U1667 (N_1667,N_1565,N_1587);
xor U1668 (N_1668,N_1533,N_1521);
xnor U1669 (N_1669,N_1544,N_1588);
nand U1670 (N_1670,N_1512,N_1501);
nor U1671 (N_1671,N_1506,N_1521);
nor U1672 (N_1672,N_1539,N_1586);
xor U1673 (N_1673,N_1576,N_1549);
xor U1674 (N_1674,N_1503,N_1591);
xnor U1675 (N_1675,N_1572,N_1582);
or U1676 (N_1676,N_1507,N_1535);
nand U1677 (N_1677,N_1558,N_1580);
and U1678 (N_1678,N_1590,N_1504);
nor U1679 (N_1679,N_1530,N_1584);
xor U1680 (N_1680,N_1559,N_1565);
nand U1681 (N_1681,N_1550,N_1506);
or U1682 (N_1682,N_1554,N_1561);
nor U1683 (N_1683,N_1575,N_1559);
nor U1684 (N_1684,N_1580,N_1551);
xor U1685 (N_1685,N_1578,N_1541);
nand U1686 (N_1686,N_1549,N_1571);
nor U1687 (N_1687,N_1597,N_1510);
and U1688 (N_1688,N_1542,N_1510);
or U1689 (N_1689,N_1587,N_1511);
nor U1690 (N_1690,N_1541,N_1572);
or U1691 (N_1691,N_1535,N_1502);
nand U1692 (N_1692,N_1569,N_1550);
nand U1693 (N_1693,N_1557,N_1561);
nand U1694 (N_1694,N_1510,N_1500);
xor U1695 (N_1695,N_1502,N_1596);
nand U1696 (N_1696,N_1571,N_1562);
or U1697 (N_1697,N_1573,N_1564);
nand U1698 (N_1698,N_1582,N_1588);
or U1699 (N_1699,N_1581,N_1507);
and U1700 (N_1700,N_1649,N_1678);
and U1701 (N_1701,N_1637,N_1650);
and U1702 (N_1702,N_1660,N_1616);
or U1703 (N_1703,N_1614,N_1673);
nor U1704 (N_1704,N_1626,N_1686);
or U1705 (N_1705,N_1674,N_1623);
nand U1706 (N_1706,N_1611,N_1665);
nor U1707 (N_1707,N_1646,N_1690);
xnor U1708 (N_1708,N_1671,N_1612);
and U1709 (N_1709,N_1651,N_1622);
nor U1710 (N_1710,N_1619,N_1648);
nand U1711 (N_1711,N_1602,N_1644);
nand U1712 (N_1712,N_1654,N_1663);
or U1713 (N_1713,N_1600,N_1694);
or U1714 (N_1714,N_1681,N_1653);
nand U1715 (N_1715,N_1672,N_1669);
or U1716 (N_1716,N_1693,N_1610);
and U1717 (N_1717,N_1680,N_1683);
or U1718 (N_1718,N_1642,N_1675);
and U1719 (N_1719,N_1630,N_1655);
nand U1720 (N_1720,N_1696,N_1647);
nor U1721 (N_1721,N_1620,N_1661);
or U1722 (N_1722,N_1617,N_1621);
nor U1723 (N_1723,N_1613,N_1641);
xnor U1724 (N_1724,N_1664,N_1636);
or U1725 (N_1725,N_1692,N_1605);
and U1726 (N_1726,N_1666,N_1657);
xor U1727 (N_1727,N_1601,N_1699);
nor U1728 (N_1728,N_1697,N_1645);
and U1729 (N_1729,N_1670,N_1625);
and U1730 (N_1730,N_1633,N_1691);
nand U1731 (N_1731,N_1632,N_1689);
xnor U1732 (N_1732,N_1668,N_1679);
xor U1733 (N_1733,N_1634,N_1606);
xnor U1734 (N_1734,N_1652,N_1624);
xor U1735 (N_1735,N_1659,N_1631);
nor U1736 (N_1736,N_1684,N_1604);
nand U1737 (N_1737,N_1640,N_1635);
and U1738 (N_1738,N_1629,N_1656);
nor U1739 (N_1739,N_1615,N_1608);
nand U1740 (N_1740,N_1688,N_1603);
xor U1741 (N_1741,N_1687,N_1658);
nor U1742 (N_1742,N_1698,N_1695);
nor U1743 (N_1743,N_1662,N_1643);
and U1744 (N_1744,N_1677,N_1682);
nand U1745 (N_1745,N_1685,N_1627);
and U1746 (N_1746,N_1607,N_1667);
and U1747 (N_1747,N_1618,N_1639);
nor U1748 (N_1748,N_1609,N_1628);
or U1749 (N_1749,N_1638,N_1676);
nand U1750 (N_1750,N_1618,N_1681);
or U1751 (N_1751,N_1679,N_1696);
and U1752 (N_1752,N_1637,N_1627);
xor U1753 (N_1753,N_1631,N_1693);
or U1754 (N_1754,N_1632,N_1680);
and U1755 (N_1755,N_1626,N_1675);
xor U1756 (N_1756,N_1689,N_1654);
xnor U1757 (N_1757,N_1612,N_1619);
nand U1758 (N_1758,N_1682,N_1655);
or U1759 (N_1759,N_1640,N_1606);
nor U1760 (N_1760,N_1665,N_1662);
xor U1761 (N_1761,N_1653,N_1643);
xor U1762 (N_1762,N_1696,N_1680);
and U1763 (N_1763,N_1618,N_1642);
or U1764 (N_1764,N_1640,N_1637);
nor U1765 (N_1765,N_1682,N_1666);
or U1766 (N_1766,N_1622,N_1664);
or U1767 (N_1767,N_1629,N_1675);
or U1768 (N_1768,N_1645,N_1623);
and U1769 (N_1769,N_1647,N_1680);
nand U1770 (N_1770,N_1675,N_1622);
and U1771 (N_1771,N_1642,N_1667);
xor U1772 (N_1772,N_1652,N_1665);
nand U1773 (N_1773,N_1618,N_1664);
and U1774 (N_1774,N_1626,N_1645);
nand U1775 (N_1775,N_1618,N_1603);
nand U1776 (N_1776,N_1686,N_1631);
or U1777 (N_1777,N_1696,N_1663);
xor U1778 (N_1778,N_1637,N_1664);
nor U1779 (N_1779,N_1638,N_1600);
xnor U1780 (N_1780,N_1629,N_1622);
nand U1781 (N_1781,N_1661,N_1682);
xor U1782 (N_1782,N_1626,N_1682);
or U1783 (N_1783,N_1652,N_1694);
and U1784 (N_1784,N_1613,N_1676);
and U1785 (N_1785,N_1681,N_1670);
and U1786 (N_1786,N_1642,N_1653);
nand U1787 (N_1787,N_1669,N_1626);
nor U1788 (N_1788,N_1692,N_1697);
nor U1789 (N_1789,N_1664,N_1696);
or U1790 (N_1790,N_1694,N_1630);
nor U1791 (N_1791,N_1692,N_1690);
xnor U1792 (N_1792,N_1647,N_1672);
nand U1793 (N_1793,N_1666,N_1627);
nand U1794 (N_1794,N_1683,N_1603);
or U1795 (N_1795,N_1648,N_1681);
and U1796 (N_1796,N_1688,N_1611);
xnor U1797 (N_1797,N_1669,N_1697);
and U1798 (N_1798,N_1698,N_1696);
or U1799 (N_1799,N_1686,N_1627);
nor U1800 (N_1800,N_1777,N_1792);
or U1801 (N_1801,N_1763,N_1720);
nand U1802 (N_1802,N_1758,N_1793);
or U1803 (N_1803,N_1790,N_1728);
nor U1804 (N_1804,N_1779,N_1746);
or U1805 (N_1805,N_1707,N_1731);
and U1806 (N_1806,N_1729,N_1776);
or U1807 (N_1807,N_1741,N_1782);
nor U1808 (N_1808,N_1752,N_1744);
or U1809 (N_1809,N_1775,N_1736);
or U1810 (N_1810,N_1724,N_1730);
and U1811 (N_1811,N_1787,N_1750);
nor U1812 (N_1812,N_1702,N_1713);
xnor U1813 (N_1813,N_1740,N_1797);
nor U1814 (N_1814,N_1761,N_1711);
or U1815 (N_1815,N_1700,N_1719);
xor U1816 (N_1816,N_1715,N_1789);
nor U1817 (N_1817,N_1703,N_1771);
nand U1818 (N_1818,N_1751,N_1721);
and U1819 (N_1819,N_1734,N_1739);
xnor U1820 (N_1820,N_1783,N_1705);
nand U1821 (N_1821,N_1706,N_1738);
xor U1822 (N_1822,N_1766,N_1768);
or U1823 (N_1823,N_1795,N_1749);
xnor U1824 (N_1824,N_1725,N_1743);
xnor U1825 (N_1825,N_1732,N_1722);
xor U1826 (N_1826,N_1774,N_1754);
and U1827 (N_1827,N_1769,N_1760);
nand U1828 (N_1828,N_1745,N_1767);
or U1829 (N_1829,N_1784,N_1717);
or U1830 (N_1830,N_1742,N_1798);
or U1831 (N_1831,N_1716,N_1748);
nor U1832 (N_1832,N_1791,N_1773);
or U1833 (N_1833,N_1727,N_1710);
and U1834 (N_1834,N_1714,N_1718);
xor U1835 (N_1835,N_1799,N_1709);
xnor U1836 (N_1836,N_1735,N_1708);
nor U1837 (N_1837,N_1755,N_1759);
and U1838 (N_1838,N_1772,N_1712);
xnor U1839 (N_1839,N_1762,N_1786);
and U1840 (N_1840,N_1781,N_1747);
and U1841 (N_1841,N_1794,N_1764);
nor U1842 (N_1842,N_1756,N_1788);
and U1843 (N_1843,N_1737,N_1778);
xor U1844 (N_1844,N_1785,N_1765);
and U1845 (N_1845,N_1733,N_1757);
nand U1846 (N_1846,N_1753,N_1701);
xor U1847 (N_1847,N_1796,N_1770);
nand U1848 (N_1848,N_1780,N_1726);
xor U1849 (N_1849,N_1704,N_1723);
or U1850 (N_1850,N_1735,N_1718);
or U1851 (N_1851,N_1705,N_1778);
nor U1852 (N_1852,N_1787,N_1761);
nand U1853 (N_1853,N_1784,N_1703);
nand U1854 (N_1854,N_1720,N_1767);
nand U1855 (N_1855,N_1753,N_1792);
nor U1856 (N_1856,N_1741,N_1723);
nor U1857 (N_1857,N_1796,N_1767);
or U1858 (N_1858,N_1741,N_1779);
or U1859 (N_1859,N_1719,N_1721);
xor U1860 (N_1860,N_1750,N_1705);
xnor U1861 (N_1861,N_1722,N_1788);
nand U1862 (N_1862,N_1788,N_1793);
or U1863 (N_1863,N_1778,N_1784);
nor U1864 (N_1864,N_1774,N_1728);
or U1865 (N_1865,N_1753,N_1761);
and U1866 (N_1866,N_1783,N_1762);
nand U1867 (N_1867,N_1755,N_1781);
nor U1868 (N_1868,N_1793,N_1756);
or U1869 (N_1869,N_1783,N_1722);
and U1870 (N_1870,N_1706,N_1702);
nor U1871 (N_1871,N_1778,N_1785);
and U1872 (N_1872,N_1770,N_1785);
nand U1873 (N_1873,N_1759,N_1787);
nor U1874 (N_1874,N_1795,N_1743);
and U1875 (N_1875,N_1792,N_1733);
nand U1876 (N_1876,N_1740,N_1755);
xnor U1877 (N_1877,N_1756,N_1703);
and U1878 (N_1878,N_1769,N_1775);
xnor U1879 (N_1879,N_1793,N_1708);
xor U1880 (N_1880,N_1793,N_1795);
xnor U1881 (N_1881,N_1738,N_1701);
and U1882 (N_1882,N_1719,N_1776);
or U1883 (N_1883,N_1713,N_1710);
and U1884 (N_1884,N_1766,N_1778);
nor U1885 (N_1885,N_1736,N_1755);
xor U1886 (N_1886,N_1703,N_1714);
nor U1887 (N_1887,N_1795,N_1762);
nor U1888 (N_1888,N_1745,N_1729);
nand U1889 (N_1889,N_1772,N_1740);
or U1890 (N_1890,N_1741,N_1762);
or U1891 (N_1891,N_1799,N_1775);
xor U1892 (N_1892,N_1757,N_1723);
xor U1893 (N_1893,N_1777,N_1799);
nor U1894 (N_1894,N_1719,N_1707);
and U1895 (N_1895,N_1774,N_1717);
xor U1896 (N_1896,N_1702,N_1701);
or U1897 (N_1897,N_1721,N_1715);
nor U1898 (N_1898,N_1775,N_1772);
xor U1899 (N_1899,N_1781,N_1729);
nand U1900 (N_1900,N_1833,N_1822);
or U1901 (N_1901,N_1855,N_1858);
xnor U1902 (N_1902,N_1883,N_1896);
nand U1903 (N_1903,N_1878,N_1888);
xnor U1904 (N_1904,N_1824,N_1847);
nand U1905 (N_1905,N_1856,N_1830);
xor U1906 (N_1906,N_1897,N_1826);
xnor U1907 (N_1907,N_1850,N_1835);
or U1908 (N_1908,N_1805,N_1898);
xnor U1909 (N_1909,N_1802,N_1862);
nand U1910 (N_1910,N_1872,N_1825);
nor U1911 (N_1911,N_1866,N_1861);
nand U1912 (N_1912,N_1844,N_1867);
xor U1913 (N_1913,N_1841,N_1879);
xor U1914 (N_1914,N_1853,N_1836);
nand U1915 (N_1915,N_1840,N_1891);
or U1916 (N_1916,N_1804,N_1877);
and U1917 (N_1917,N_1859,N_1848);
nand U1918 (N_1918,N_1865,N_1893);
and U1919 (N_1919,N_1827,N_1870);
nor U1920 (N_1920,N_1813,N_1814);
nand U1921 (N_1921,N_1876,N_1846);
nand U1922 (N_1922,N_1837,N_1812);
xor U1923 (N_1923,N_1887,N_1834);
xor U1924 (N_1924,N_1828,N_1863);
and U1925 (N_1925,N_1845,N_1818);
or U1926 (N_1926,N_1803,N_1852);
or U1927 (N_1927,N_1821,N_1808);
and U1928 (N_1928,N_1871,N_1801);
nor U1929 (N_1929,N_1882,N_1869);
xor U1930 (N_1930,N_1875,N_1899);
or U1931 (N_1931,N_1809,N_1864);
or U1932 (N_1932,N_1831,N_1815);
xor U1933 (N_1933,N_1857,N_1895);
nor U1934 (N_1934,N_1881,N_1823);
and U1935 (N_1935,N_1884,N_1874);
nor U1936 (N_1936,N_1811,N_1819);
or U1937 (N_1937,N_1894,N_1868);
and U1938 (N_1938,N_1832,N_1820);
nand U1939 (N_1939,N_1839,N_1890);
and U1940 (N_1940,N_1816,N_1807);
xnor U1941 (N_1941,N_1892,N_1829);
xnor U1942 (N_1942,N_1817,N_1810);
nor U1943 (N_1943,N_1885,N_1860);
xor U1944 (N_1944,N_1849,N_1842);
nor U1945 (N_1945,N_1843,N_1886);
nor U1946 (N_1946,N_1806,N_1800);
or U1947 (N_1947,N_1854,N_1880);
or U1948 (N_1948,N_1873,N_1889);
nand U1949 (N_1949,N_1838,N_1851);
and U1950 (N_1950,N_1873,N_1894);
nand U1951 (N_1951,N_1810,N_1831);
nor U1952 (N_1952,N_1866,N_1872);
xor U1953 (N_1953,N_1885,N_1839);
nor U1954 (N_1954,N_1894,N_1826);
and U1955 (N_1955,N_1880,N_1871);
nor U1956 (N_1956,N_1816,N_1885);
nor U1957 (N_1957,N_1815,N_1876);
nor U1958 (N_1958,N_1870,N_1872);
xnor U1959 (N_1959,N_1805,N_1822);
nand U1960 (N_1960,N_1836,N_1823);
nor U1961 (N_1961,N_1850,N_1861);
or U1962 (N_1962,N_1812,N_1896);
and U1963 (N_1963,N_1808,N_1843);
nand U1964 (N_1964,N_1813,N_1827);
and U1965 (N_1965,N_1821,N_1850);
xnor U1966 (N_1966,N_1810,N_1866);
nand U1967 (N_1967,N_1823,N_1894);
nor U1968 (N_1968,N_1884,N_1801);
xor U1969 (N_1969,N_1802,N_1883);
xor U1970 (N_1970,N_1809,N_1804);
xnor U1971 (N_1971,N_1847,N_1858);
xnor U1972 (N_1972,N_1891,N_1849);
or U1973 (N_1973,N_1812,N_1808);
or U1974 (N_1974,N_1803,N_1832);
and U1975 (N_1975,N_1800,N_1832);
nand U1976 (N_1976,N_1830,N_1861);
nand U1977 (N_1977,N_1892,N_1807);
nor U1978 (N_1978,N_1836,N_1890);
or U1979 (N_1979,N_1841,N_1830);
xor U1980 (N_1980,N_1820,N_1856);
xor U1981 (N_1981,N_1810,N_1881);
xor U1982 (N_1982,N_1815,N_1839);
nor U1983 (N_1983,N_1823,N_1891);
and U1984 (N_1984,N_1835,N_1886);
xor U1985 (N_1985,N_1886,N_1809);
or U1986 (N_1986,N_1899,N_1866);
nor U1987 (N_1987,N_1834,N_1850);
nor U1988 (N_1988,N_1820,N_1879);
or U1989 (N_1989,N_1849,N_1894);
or U1990 (N_1990,N_1818,N_1828);
nand U1991 (N_1991,N_1886,N_1896);
xor U1992 (N_1992,N_1893,N_1804);
and U1993 (N_1993,N_1895,N_1811);
and U1994 (N_1994,N_1875,N_1817);
and U1995 (N_1995,N_1801,N_1808);
and U1996 (N_1996,N_1888,N_1833);
and U1997 (N_1997,N_1887,N_1888);
xor U1998 (N_1998,N_1860,N_1846);
nand U1999 (N_1999,N_1882,N_1870);
or U2000 (N_2000,N_1932,N_1924);
xor U2001 (N_2001,N_1900,N_1955);
and U2002 (N_2002,N_1986,N_1912);
nand U2003 (N_2003,N_1998,N_1918);
nor U2004 (N_2004,N_1979,N_1907);
nand U2005 (N_2005,N_1981,N_1992);
or U2006 (N_2006,N_1977,N_1919);
xor U2007 (N_2007,N_1911,N_1965);
nor U2008 (N_2008,N_1936,N_1927);
or U2009 (N_2009,N_1967,N_1949);
nor U2010 (N_2010,N_1996,N_1970);
nor U2011 (N_2011,N_1956,N_1929);
xor U2012 (N_2012,N_1997,N_1994);
nor U2013 (N_2013,N_1957,N_1974);
nand U2014 (N_2014,N_1964,N_1990);
and U2015 (N_2015,N_1931,N_1940);
or U2016 (N_2016,N_1989,N_1922);
or U2017 (N_2017,N_1944,N_1937);
nand U2018 (N_2018,N_1953,N_1909);
xnor U2019 (N_2019,N_1901,N_1993);
or U2020 (N_2020,N_1969,N_1991);
nand U2021 (N_2021,N_1920,N_1948);
nor U2022 (N_2022,N_1903,N_1950);
xnor U2023 (N_2023,N_1954,N_1988);
or U2024 (N_2024,N_1943,N_1942);
and U2025 (N_2025,N_1985,N_1961);
and U2026 (N_2026,N_1925,N_1951);
or U2027 (N_2027,N_1984,N_1966);
and U2028 (N_2028,N_1938,N_1975);
nand U2029 (N_2029,N_1930,N_1982);
nor U2030 (N_2030,N_1959,N_1971);
nand U2031 (N_2031,N_1973,N_1960);
nand U2032 (N_2032,N_1978,N_1952);
nand U2033 (N_2033,N_1972,N_1934);
and U2034 (N_2034,N_1921,N_1935);
nor U2035 (N_2035,N_1999,N_1968);
and U2036 (N_2036,N_1963,N_1905);
xor U2037 (N_2037,N_1916,N_1995);
and U2038 (N_2038,N_1933,N_1980);
xnor U2039 (N_2039,N_1941,N_1946);
and U2040 (N_2040,N_1939,N_1947);
nor U2041 (N_2041,N_1917,N_1908);
nor U2042 (N_2042,N_1928,N_1913);
or U2043 (N_2043,N_1914,N_1910);
nor U2044 (N_2044,N_1915,N_1945);
or U2045 (N_2045,N_1976,N_1906);
nor U2046 (N_2046,N_1926,N_1904);
or U2047 (N_2047,N_1983,N_1962);
nand U2048 (N_2048,N_1958,N_1902);
or U2049 (N_2049,N_1987,N_1923);
nor U2050 (N_2050,N_1964,N_1934);
nor U2051 (N_2051,N_1970,N_1932);
and U2052 (N_2052,N_1911,N_1933);
nand U2053 (N_2053,N_1966,N_1965);
and U2054 (N_2054,N_1970,N_1989);
nor U2055 (N_2055,N_1968,N_1972);
and U2056 (N_2056,N_1981,N_1997);
xnor U2057 (N_2057,N_1989,N_1984);
and U2058 (N_2058,N_1932,N_1955);
and U2059 (N_2059,N_1962,N_1913);
or U2060 (N_2060,N_1984,N_1983);
xor U2061 (N_2061,N_1961,N_1992);
xor U2062 (N_2062,N_1946,N_1990);
or U2063 (N_2063,N_1979,N_1903);
nand U2064 (N_2064,N_1913,N_1955);
or U2065 (N_2065,N_1923,N_1956);
xnor U2066 (N_2066,N_1914,N_1958);
xor U2067 (N_2067,N_1985,N_1934);
or U2068 (N_2068,N_1926,N_1947);
nor U2069 (N_2069,N_1910,N_1998);
or U2070 (N_2070,N_1953,N_1947);
and U2071 (N_2071,N_1959,N_1935);
nor U2072 (N_2072,N_1994,N_1902);
nand U2073 (N_2073,N_1937,N_1966);
or U2074 (N_2074,N_1994,N_1904);
xnor U2075 (N_2075,N_1910,N_1941);
nor U2076 (N_2076,N_1959,N_1958);
or U2077 (N_2077,N_1963,N_1960);
and U2078 (N_2078,N_1955,N_1946);
nor U2079 (N_2079,N_1922,N_1980);
or U2080 (N_2080,N_1928,N_1914);
and U2081 (N_2081,N_1991,N_1984);
nor U2082 (N_2082,N_1909,N_1933);
nand U2083 (N_2083,N_1912,N_1957);
and U2084 (N_2084,N_1946,N_1983);
or U2085 (N_2085,N_1947,N_1912);
xor U2086 (N_2086,N_1997,N_1960);
or U2087 (N_2087,N_1919,N_1910);
and U2088 (N_2088,N_1919,N_1937);
and U2089 (N_2089,N_1927,N_1973);
and U2090 (N_2090,N_1970,N_1971);
and U2091 (N_2091,N_1975,N_1916);
or U2092 (N_2092,N_1945,N_1939);
xnor U2093 (N_2093,N_1983,N_1957);
nor U2094 (N_2094,N_1936,N_1910);
nor U2095 (N_2095,N_1913,N_1929);
nand U2096 (N_2096,N_1967,N_1927);
or U2097 (N_2097,N_1982,N_1962);
xnor U2098 (N_2098,N_1956,N_1937);
nor U2099 (N_2099,N_1991,N_1971);
xor U2100 (N_2100,N_2046,N_2048);
or U2101 (N_2101,N_2036,N_2038);
nand U2102 (N_2102,N_2085,N_2014);
or U2103 (N_2103,N_2027,N_2071);
xnor U2104 (N_2104,N_2096,N_2063);
nor U2105 (N_2105,N_2025,N_2033);
nand U2106 (N_2106,N_2062,N_2007);
and U2107 (N_2107,N_2020,N_2052);
nor U2108 (N_2108,N_2029,N_2082);
nand U2109 (N_2109,N_2001,N_2043);
nor U2110 (N_2110,N_2010,N_2009);
or U2111 (N_2111,N_2037,N_2054);
or U2112 (N_2112,N_2034,N_2053);
nand U2113 (N_2113,N_2057,N_2067);
and U2114 (N_2114,N_2090,N_2031);
and U2115 (N_2115,N_2069,N_2022);
nor U2116 (N_2116,N_2086,N_2042);
xor U2117 (N_2117,N_2081,N_2028);
or U2118 (N_2118,N_2066,N_2044);
nand U2119 (N_2119,N_2019,N_2015);
or U2120 (N_2120,N_2091,N_2041);
or U2121 (N_2121,N_2084,N_2060);
nor U2122 (N_2122,N_2018,N_2047);
nand U2123 (N_2123,N_2077,N_2040);
nor U2124 (N_2124,N_2032,N_2070);
nand U2125 (N_2125,N_2058,N_2087);
nand U2126 (N_2126,N_2049,N_2094);
nand U2127 (N_2127,N_2000,N_2012);
nand U2128 (N_2128,N_2075,N_2039);
and U2129 (N_2129,N_2098,N_2061);
and U2130 (N_2130,N_2003,N_2002);
nand U2131 (N_2131,N_2079,N_2076);
and U2132 (N_2132,N_2072,N_2021);
or U2133 (N_2133,N_2051,N_2006);
or U2134 (N_2134,N_2088,N_2083);
or U2135 (N_2135,N_2099,N_2097);
nand U2136 (N_2136,N_2093,N_2089);
xnor U2137 (N_2137,N_2026,N_2092);
nor U2138 (N_2138,N_2078,N_2030);
nor U2139 (N_2139,N_2080,N_2065);
and U2140 (N_2140,N_2073,N_2059);
xor U2141 (N_2141,N_2045,N_2050);
nand U2142 (N_2142,N_2023,N_2005);
nor U2143 (N_2143,N_2095,N_2017);
or U2144 (N_2144,N_2004,N_2055);
xor U2145 (N_2145,N_2013,N_2064);
or U2146 (N_2146,N_2008,N_2035);
or U2147 (N_2147,N_2011,N_2068);
or U2148 (N_2148,N_2074,N_2056);
or U2149 (N_2149,N_2024,N_2016);
nor U2150 (N_2150,N_2001,N_2051);
nor U2151 (N_2151,N_2067,N_2010);
or U2152 (N_2152,N_2029,N_2024);
xnor U2153 (N_2153,N_2088,N_2051);
or U2154 (N_2154,N_2016,N_2064);
or U2155 (N_2155,N_2002,N_2006);
nor U2156 (N_2156,N_2047,N_2008);
or U2157 (N_2157,N_2026,N_2024);
or U2158 (N_2158,N_2058,N_2011);
xor U2159 (N_2159,N_2011,N_2034);
xnor U2160 (N_2160,N_2058,N_2035);
nand U2161 (N_2161,N_2012,N_2066);
or U2162 (N_2162,N_2015,N_2058);
nand U2163 (N_2163,N_2023,N_2018);
nor U2164 (N_2164,N_2031,N_2002);
or U2165 (N_2165,N_2053,N_2077);
and U2166 (N_2166,N_2066,N_2075);
and U2167 (N_2167,N_2075,N_2083);
or U2168 (N_2168,N_2057,N_2096);
nand U2169 (N_2169,N_2045,N_2087);
nand U2170 (N_2170,N_2011,N_2017);
xnor U2171 (N_2171,N_2087,N_2078);
or U2172 (N_2172,N_2061,N_2046);
or U2173 (N_2173,N_2063,N_2047);
xor U2174 (N_2174,N_2092,N_2093);
xnor U2175 (N_2175,N_2093,N_2038);
nand U2176 (N_2176,N_2049,N_2059);
nor U2177 (N_2177,N_2034,N_2070);
and U2178 (N_2178,N_2049,N_2046);
nand U2179 (N_2179,N_2035,N_2030);
or U2180 (N_2180,N_2015,N_2020);
or U2181 (N_2181,N_2083,N_2004);
nor U2182 (N_2182,N_2032,N_2088);
xor U2183 (N_2183,N_2012,N_2090);
and U2184 (N_2184,N_2015,N_2081);
or U2185 (N_2185,N_2004,N_2046);
xnor U2186 (N_2186,N_2052,N_2027);
nor U2187 (N_2187,N_2067,N_2094);
nand U2188 (N_2188,N_2049,N_2058);
nand U2189 (N_2189,N_2045,N_2076);
xor U2190 (N_2190,N_2038,N_2033);
or U2191 (N_2191,N_2025,N_2042);
xor U2192 (N_2192,N_2001,N_2096);
xor U2193 (N_2193,N_2047,N_2029);
xnor U2194 (N_2194,N_2016,N_2036);
xnor U2195 (N_2195,N_2065,N_2047);
or U2196 (N_2196,N_2087,N_2099);
xor U2197 (N_2197,N_2059,N_2027);
or U2198 (N_2198,N_2065,N_2036);
xnor U2199 (N_2199,N_2065,N_2012);
nor U2200 (N_2200,N_2199,N_2149);
nor U2201 (N_2201,N_2134,N_2106);
and U2202 (N_2202,N_2125,N_2104);
or U2203 (N_2203,N_2141,N_2160);
and U2204 (N_2204,N_2120,N_2135);
nor U2205 (N_2205,N_2157,N_2158);
nand U2206 (N_2206,N_2165,N_2152);
or U2207 (N_2207,N_2118,N_2105);
nor U2208 (N_2208,N_2191,N_2183);
nor U2209 (N_2209,N_2185,N_2151);
xor U2210 (N_2210,N_2146,N_2132);
xor U2211 (N_2211,N_2192,N_2142);
nor U2212 (N_2212,N_2147,N_2176);
nand U2213 (N_2213,N_2189,N_2170);
nand U2214 (N_2214,N_2186,N_2187);
nand U2215 (N_2215,N_2167,N_2195);
xor U2216 (N_2216,N_2113,N_2115);
nor U2217 (N_2217,N_2168,N_2145);
nand U2218 (N_2218,N_2179,N_2100);
and U2219 (N_2219,N_2119,N_2178);
nand U2220 (N_2220,N_2153,N_2198);
or U2221 (N_2221,N_2171,N_2116);
or U2222 (N_2222,N_2144,N_2112);
and U2223 (N_2223,N_2193,N_2137);
nand U2224 (N_2224,N_2129,N_2127);
nor U2225 (N_2225,N_2182,N_2111);
and U2226 (N_2226,N_2156,N_2103);
nor U2227 (N_2227,N_2163,N_2130);
nor U2228 (N_2228,N_2107,N_2140);
or U2229 (N_2229,N_2122,N_2194);
nor U2230 (N_2230,N_2102,N_2175);
nand U2231 (N_2231,N_2184,N_2166);
and U2232 (N_2232,N_2150,N_2133);
or U2233 (N_2233,N_2143,N_2154);
or U2234 (N_2234,N_2139,N_2190);
nor U2235 (N_2235,N_2136,N_2108);
xor U2236 (N_2236,N_2197,N_2117);
and U2237 (N_2237,N_2109,N_2128);
nand U2238 (N_2238,N_2121,N_2101);
xnor U2239 (N_2239,N_2159,N_2123);
nor U2240 (N_2240,N_2174,N_2124);
xor U2241 (N_2241,N_2172,N_2181);
or U2242 (N_2242,N_2164,N_2180);
and U2243 (N_2243,N_2148,N_2196);
nor U2244 (N_2244,N_2162,N_2138);
or U2245 (N_2245,N_2173,N_2155);
xnor U2246 (N_2246,N_2177,N_2161);
or U2247 (N_2247,N_2131,N_2169);
and U2248 (N_2248,N_2188,N_2126);
or U2249 (N_2249,N_2114,N_2110);
xor U2250 (N_2250,N_2115,N_2121);
nand U2251 (N_2251,N_2142,N_2106);
xor U2252 (N_2252,N_2157,N_2159);
or U2253 (N_2253,N_2110,N_2113);
nand U2254 (N_2254,N_2101,N_2154);
or U2255 (N_2255,N_2123,N_2143);
nand U2256 (N_2256,N_2129,N_2105);
or U2257 (N_2257,N_2170,N_2125);
xnor U2258 (N_2258,N_2132,N_2154);
or U2259 (N_2259,N_2199,N_2185);
xnor U2260 (N_2260,N_2115,N_2187);
or U2261 (N_2261,N_2165,N_2183);
nor U2262 (N_2262,N_2187,N_2112);
and U2263 (N_2263,N_2194,N_2165);
nand U2264 (N_2264,N_2117,N_2175);
nand U2265 (N_2265,N_2179,N_2115);
nand U2266 (N_2266,N_2134,N_2148);
nor U2267 (N_2267,N_2129,N_2180);
and U2268 (N_2268,N_2115,N_2180);
or U2269 (N_2269,N_2197,N_2188);
and U2270 (N_2270,N_2196,N_2101);
and U2271 (N_2271,N_2110,N_2177);
nand U2272 (N_2272,N_2139,N_2114);
xnor U2273 (N_2273,N_2138,N_2107);
and U2274 (N_2274,N_2122,N_2133);
nand U2275 (N_2275,N_2109,N_2187);
nand U2276 (N_2276,N_2107,N_2196);
nor U2277 (N_2277,N_2126,N_2106);
xor U2278 (N_2278,N_2187,N_2108);
or U2279 (N_2279,N_2125,N_2119);
nand U2280 (N_2280,N_2153,N_2156);
or U2281 (N_2281,N_2190,N_2177);
or U2282 (N_2282,N_2191,N_2115);
nor U2283 (N_2283,N_2149,N_2171);
or U2284 (N_2284,N_2121,N_2182);
nand U2285 (N_2285,N_2189,N_2188);
nor U2286 (N_2286,N_2147,N_2188);
xnor U2287 (N_2287,N_2102,N_2131);
and U2288 (N_2288,N_2179,N_2188);
nor U2289 (N_2289,N_2175,N_2129);
or U2290 (N_2290,N_2109,N_2112);
and U2291 (N_2291,N_2126,N_2123);
or U2292 (N_2292,N_2115,N_2143);
and U2293 (N_2293,N_2179,N_2132);
nand U2294 (N_2294,N_2130,N_2110);
or U2295 (N_2295,N_2114,N_2184);
xor U2296 (N_2296,N_2157,N_2122);
or U2297 (N_2297,N_2125,N_2151);
or U2298 (N_2298,N_2116,N_2188);
xor U2299 (N_2299,N_2134,N_2120);
xor U2300 (N_2300,N_2278,N_2243);
and U2301 (N_2301,N_2239,N_2223);
nand U2302 (N_2302,N_2268,N_2226);
nor U2303 (N_2303,N_2242,N_2252);
xor U2304 (N_2304,N_2263,N_2274);
and U2305 (N_2305,N_2200,N_2281);
and U2306 (N_2306,N_2244,N_2230);
xnor U2307 (N_2307,N_2295,N_2249);
xnor U2308 (N_2308,N_2280,N_2257);
nand U2309 (N_2309,N_2270,N_2292);
nor U2310 (N_2310,N_2262,N_2228);
nand U2311 (N_2311,N_2279,N_2222);
or U2312 (N_2312,N_2221,N_2210);
nand U2313 (N_2313,N_2241,N_2253);
xor U2314 (N_2314,N_2238,N_2251);
nand U2315 (N_2315,N_2258,N_2291);
nand U2316 (N_2316,N_2259,N_2276);
xor U2317 (N_2317,N_2273,N_2256);
or U2318 (N_2318,N_2247,N_2240);
and U2319 (N_2319,N_2267,N_2203);
nor U2320 (N_2320,N_2261,N_2293);
nand U2321 (N_2321,N_2212,N_2275);
nor U2322 (N_2322,N_2250,N_2246);
or U2323 (N_2323,N_2287,N_2206);
xor U2324 (N_2324,N_2205,N_2211);
and U2325 (N_2325,N_2294,N_2285);
or U2326 (N_2326,N_2237,N_2214);
or U2327 (N_2327,N_2218,N_2269);
and U2328 (N_2328,N_2227,N_2233);
nor U2329 (N_2329,N_2208,N_2201);
nand U2330 (N_2330,N_2266,N_2289);
nand U2331 (N_2331,N_2283,N_2282);
nand U2332 (N_2332,N_2209,N_2216);
or U2333 (N_2333,N_2229,N_2297);
xnor U2334 (N_2334,N_2299,N_2213);
and U2335 (N_2335,N_2296,N_2245);
nor U2336 (N_2336,N_2255,N_2231);
xor U2337 (N_2337,N_2298,N_2284);
nand U2338 (N_2338,N_2224,N_2265);
xnor U2339 (N_2339,N_2264,N_2288);
and U2340 (N_2340,N_2277,N_2286);
and U2341 (N_2341,N_2215,N_2236);
xor U2342 (N_2342,N_2207,N_2232);
nor U2343 (N_2343,N_2204,N_2217);
xor U2344 (N_2344,N_2272,N_2234);
or U2345 (N_2345,N_2225,N_2202);
and U2346 (N_2346,N_2290,N_2248);
nand U2347 (N_2347,N_2235,N_2219);
or U2348 (N_2348,N_2220,N_2271);
nor U2349 (N_2349,N_2260,N_2254);
nand U2350 (N_2350,N_2242,N_2239);
or U2351 (N_2351,N_2227,N_2258);
and U2352 (N_2352,N_2250,N_2239);
or U2353 (N_2353,N_2255,N_2259);
or U2354 (N_2354,N_2288,N_2273);
nor U2355 (N_2355,N_2238,N_2223);
xnor U2356 (N_2356,N_2281,N_2203);
and U2357 (N_2357,N_2258,N_2208);
or U2358 (N_2358,N_2237,N_2299);
nor U2359 (N_2359,N_2291,N_2231);
nand U2360 (N_2360,N_2220,N_2289);
nor U2361 (N_2361,N_2229,N_2276);
xor U2362 (N_2362,N_2234,N_2278);
and U2363 (N_2363,N_2267,N_2236);
nand U2364 (N_2364,N_2259,N_2219);
xor U2365 (N_2365,N_2274,N_2256);
xnor U2366 (N_2366,N_2236,N_2201);
nand U2367 (N_2367,N_2290,N_2279);
nand U2368 (N_2368,N_2283,N_2226);
nor U2369 (N_2369,N_2253,N_2297);
and U2370 (N_2370,N_2290,N_2249);
nor U2371 (N_2371,N_2224,N_2248);
nor U2372 (N_2372,N_2280,N_2212);
nor U2373 (N_2373,N_2278,N_2281);
xor U2374 (N_2374,N_2275,N_2239);
xor U2375 (N_2375,N_2284,N_2288);
or U2376 (N_2376,N_2257,N_2228);
or U2377 (N_2377,N_2257,N_2226);
nand U2378 (N_2378,N_2267,N_2222);
or U2379 (N_2379,N_2246,N_2226);
and U2380 (N_2380,N_2211,N_2201);
xnor U2381 (N_2381,N_2241,N_2279);
nand U2382 (N_2382,N_2252,N_2283);
and U2383 (N_2383,N_2262,N_2234);
nand U2384 (N_2384,N_2266,N_2268);
and U2385 (N_2385,N_2210,N_2269);
or U2386 (N_2386,N_2264,N_2267);
nand U2387 (N_2387,N_2265,N_2258);
xnor U2388 (N_2388,N_2211,N_2297);
or U2389 (N_2389,N_2221,N_2248);
or U2390 (N_2390,N_2271,N_2291);
xor U2391 (N_2391,N_2201,N_2202);
nand U2392 (N_2392,N_2229,N_2245);
and U2393 (N_2393,N_2230,N_2223);
xnor U2394 (N_2394,N_2226,N_2218);
or U2395 (N_2395,N_2244,N_2226);
and U2396 (N_2396,N_2235,N_2289);
nand U2397 (N_2397,N_2206,N_2285);
and U2398 (N_2398,N_2207,N_2214);
xor U2399 (N_2399,N_2257,N_2275);
nand U2400 (N_2400,N_2386,N_2363);
or U2401 (N_2401,N_2322,N_2326);
nor U2402 (N_2402,N_2341,N_2397);
nor U2403 (N_2403,N_2387,N_2331);
or U2404 (N_2404,N_2372,N_2343);
xnor U2405 (N_2405,N_2394,N_2328);
nor U2406 (N_2406,N_2351,N_2303);
nand U2407 (N_2407,N_2356,N_2307);
xor U2408 (N_2408,N_2396,N_2318);
or U2409 (N_2409,N_2361,N_2384);
nor U2410 (N_2410,N_2395,N_2357);
and U2411 (N_2411,N_2316,N_2374);
and U2412 (N_2412,N_2347,N_2306);
xor U2413 (N_2413,N_2308,N_2360);
nand U2414 (N_2414,N_2364,N_2305);
or U2415 (N_2415,N_2353,N_2368);
or U2416 (N_2416,N_2332,N_2345);
and U2417 (N_2417,N_2339,N_2329);
or U2418 (N_2418,N_2348,N_2389);
xnor U2419 (N_2419,N_2390,N_2323);
or U2420 (N_2420,N_2362,N_2385);
nand U2421 (N_2421,N_2349,N_2315);
nor U2422 (N_2422,N_2317,N_2312);
nor U2423 (N_2423,N_2301,N_2314);
and U2424 (N_2424,N_2330,N_2393);
nand U2425 (N_2425,N_2373,N_2336);
nor U2426 (N_2426,N_2365,N_2380);
or U2427 (N_2427,N_2378,N_2346);
and U2428 (N_2428,N_2392,N_2311);
nand U2429 (N_2429,N_2302,N_2366);
nor U2430 (N_2430,N_2382,N_2335);
nor U2431 (N_2431,N_2370,N_2388);
and U2432 (N_2432,N_2321,N_2379);
and U2433 (N_2433,N_2355,N_2334);
nor U2434 (N_2434,N_2376,N_2383);
nand U2435 (N_2435,N_2337,N_2359);
nor U2436 (N_2436,N_2304,N_2352);
nand U2437 (N_2437,N_2371,N_2319);
or U2438 (N_2438,N_2320,N_2327);
nand U2439 (N_2439,N_2340,N_2300);
xor U2440 (N_2440,N_2309,N_2369);
or U2441 (N_2441,N_2367,N_2333);
or U2442 (N_2442,N_2358,N_2399);
nand U2443 (N_2443,N_2313,N_2350);
nand U2444 (N_2444,N_2338,N_2324);
and U2445 (N_2445,N_2381,N_2342);
or U2446 (N_2446,N_2375,N_2377);
or U2447 (N_2447,N_2310,N_2391);
and U2448 (N_2448,N_2398,N_2325);
or U2449 (N_2449,N_2354,N_2344);
nand U2450 (N_2450,N_2318,N_2343);
and U2451 (N_2451,N_2378,N_2334);
or U2452 (N_2452,N_2377,N_2340);
and U2453 (N_2453,N_2391,N_2390);
nand U2454 (N_2454,N_2327,N_2391);
and U2455 (N_2455,N_2317,N_2343);
nand U2456 (N_2456,N_2348,N_2338);
nor U2457 (N_2457,N_2349,N_2371);
and U2458 (N_2458,N_2331,N_2332);
nor U2459 (N_2459,N_2357,N_2301);
and U2460 (N_2460,N_2389,N_2321);
and U2461 (N_2461,N_2383,N_2337);
xor U2462 (N_2462,N_2357,N_2379);
nor U2463 (N_2463,N_2384,N_2360);
or U2464 (N_2464,N_2306,N_2315);
nand U2465 (N_2465,N_2322,N_2396);
xnor U2466 (N_2466,N_2377,N_2301);
and U2467 (N_2467,N_2385,N_2345);
nand U2468 (N_2468,N_2333,N_2384);
and U2469 (N_2469,N_2373,N_2327);
or U2470 (N_2470,N_2332,N_2371);
and U2471 (N_2471,N_2326,N_2347);
nand U2472 (N_2472,N_2370,N_2324);
or U2473 (N_2473,N_2374,N_2336);
and U2474 (N_2474,N_2375,N_2320);
xnor U2475 (N_2475,N_2365,N_2351);
or U2476 (N_2476,N_2344,N_2397);
or U2477 (N_2477,N_2376,N_2391);
or U2478 (N_2478,N_2355,N_2371);
nand U2479 (N_2479,N_2330,N_2370);
or U2480 (N_2480,N_2301,N_2383);
nor U2481 (N_2481,N_2312,N_2363);
and U2482 (N_2482,N_2330,N_2329);
and U2483 (N_2483,N_2383,N_2391);
nor U2484 (N_2484,N_2335,N_2339);
nand U2485 (N_2485,N_2387,N_2316);
nor U2486 (N_2486,N_2330,N_2320);
nor U2487 (N_2487,N_2355,N_2382);
nor U2488 (N_2488,N_2302,N_2348);
nand U2489 (N_2489,N_2394,N_2397);
nor U2490 (N_2490,N_2317,N_2361);
nand U2491 (N_2491,N_2372,N_2373);
xor U2492 (N_2492,N_2331,N_2329);
xor U2493 (N_2493,N_2312,N_2340);
nor U2494 (N_2494,N_2342,N_2399);
or U2495 (N_2495,N_2355,N_2313);
nand U2496 (N_2496,N_2327,N_2390);
or U2497 (N_2497,N_2391,N_2305);
and U2498 (N_2498,N_2393,N_2340);
and U2499 (N_2499,N_2335,N_2333);
xnor U2500 (N_2500,N_2465,N_2402);
nand U2501 (N_2501,N_2451,N_2426);
nand U2502 (N_2502,N_2441,N_2473);
nand U2503 (N_2503,N_2420,N_2437);
nor U2504 (N_2504,N_2416,N_2461);
and U2505 (N_2505,N_2459,N_2482);
nor U2506 (N_2506,N_2483,N_2462);
or U2507 (N_2507,N_2492,N_2455);
nor U2508 (N_2508,N_2425,N_2464);
nand U2509 (N_2509,N_2417,N_2466);
and U2510 (N_2510,N_2495,N_2481);
nand U2511 (N_2511,N_2443,N_2468);
nand U2512 (N_2512,N_2438,N_2419);
nor U2513 (N_2513,N_2496,N_2401);
xor U2514 (N_2514,N_2439,N_2424);
nand U2515 (N_2515,N_2427,N_2412);
xnor U2516 (N_2516,N_2403,N_2474);
nand U2517 (N_2517,N_2400,N_2484);
nand U2518 (N_2518,N_2435,N_2479);
nand U2519 (N_2519,N_2422,N_2405);
nor U2520 (N_2520,N_2454,N_2447);
nor U2521 (N_2521,N_2491,N_2470);
and U2522 (N_2522,N_2429,N_2449);
nand U2523 (N_2523,N_2406,N_2497);
and U2524 (N_2524,N_2411,N_2457);
nor U2525 (N_2525,N_2452,N_2456);
and U2526 (N_2526,N_2440,N_2488);
nor U2527 (N_2527,N_2409,N_2480);
nor U2528 (N_2528,N_2444,N_2493);
nand U2529 (N_2529,N_2442,N_2490);
nor U2530 (N_2530,N_2428,N_2487);
xnor U2531 (N_2531,N_2430,N_2436);
nor U2532 (N_2532,N_2494,N_2453);
nor U2533 (N_2533,N_2489,N_2460);
nand U2534 (N_2534,N_2458,N_2434);
or U2535 (N_2535,N_2463,N_2485);
xnor U2536 (N_2536,N_2450,N_2445);
nor U2537 (N_2537,N_2446,N_2448);
nand U2538 (N_2538,N_2499,N_2431);
nand U2539 (N_2539,N_2413,N_2432);
xnor U2540 (N_2540,N_2498,N_2478);
nand U2541 (N_2541,N_2433,N_2476);
nand U2542 (N_2542,N_2467,N_2477);
xor U2543 (N_2543,N_2423,N_2475);
xor U2544 (N_2544,N_2471,N_2418);
and U2545 (N_2545,N_2404,N_2414);
nand U2546 (N_2546,N_2415,N_2486);
xnor U2547 (N_2547,N_2410,N_2472);
nor U2548 (N_2548,N_2469,N_2408);
xnor U2549 (N_2549,N_2421,N_2407);
or U2550 (N_2550,N_2489,N_2479);
and U2551 (N_2551,N_2433,N_2485);
or U2552 (N_2552,N_2467,N_2472);
or U2553 (N_2553,N_2470,N_2487);
and U2554 (N_2554,N_2499,N_2488);
or U2555 (N_2555,N_2451,N_2497);
or U2556 (N_2556,N_2420,N_2424);
or U2557 (N_2557,N_2484,N_2449);
and U2558 (N_2558,N_2450,N_2482);
or U2559 (N_2559,N_2442,N_2415);
nand U2560 (N_2560,N_2473,N_2475);
nand U2561 (N_2561,N_2488,N_2487);
nor U2562 (N_2562,N_2449,N_2462);
or U2563 (N_2563,N_2445,N_2483);
or U2564 (N_2564,N_2446,N_2498);
nand U2565 (N_2565,N_2439,N_2417);
xnor U2566 (N_2566,N_2460,N_2421);
nor U2567 (N_2567,N_2452,N_2427);
nor U2568 (N_2568,N_2438,N_2481);
or U2569 (N_2569,N_2496,N_2428);
or U2570 (N_2570,N_2463,N_2460);
nor U2571 (N_2571,N_2401,N_2408);
nand U2572 (N_2572,N_2423,N_2460);
nor U2573 (N_2573,N_2474,N_2469);
xor U2574 (N_2574,N_2416,N_2455);
nor U2575 (N_2575,N_2442,N_2418);
or U2576 (N_2576,N_2409,N_2492);
xnor U2577 (N_2577,N_2400,N_2414);
or U2578 (N_2578,N_2422,N_2438);
xnor U2579 (N_2579,N_2473,N_2435);
and U2580 (N_2580,N_2467,N_2447);
xnor U2581 (N_2581,N_2483,N_2488);
nand U2582 (N_2582,N_2416,N_2442);
or U2583 (N_2583,N_2446,N_2490);
and U2584 (N_2584,N_2476,N_2478);
or U2585 (N_2585,N_2435,N_2485);
or U2586 (N_2586,N_2430,N_2406);
or U2587 (N_2587,N_2402,N_2478);
or U2588 (N_2588,N_2491,N_2493);
nor U2589 (N_2589,N_2457,N_2431);
nand U2590 (N_2590,N_2458,N_2405);
nor U2591 (N_2591,N_2413,N_2496);
nor U2592 (N_2592,N_2497,N_2445);
and U2593 (N_2593,N_2428,N_2481);
or U2594 (N_2594,N_2415,N_2420);
or U2595 (N_2595,N_2496,N_2452);
nand U2596 (N_2596,N_2451,N_2417);
xor U2597 (N_2597,N_2477,N_2485);
xnor U2598 (N_2598,N_2474,N_2462);
xnor U2599 (N_2599,N_2488,N_2462);
xnor U2600 (N_2600,N_2504,N_2562);
nor U2601 (N_2601,N_2535,N_2542);
nor U2602 (N_2602,N_2528,N_2516);
xor U2603 (N_2603,N_2508,N_2578);
or U2604 (N_2604,N_2559,N_2569);
nand U2605 (N_2605,N_2538,N_2551);
nor U2606 (N_2606,N_2541,N_2586);
nand U2607 (N_2607,N_2573,N_2530);
nor U2608 (N_2608,N_2544,N_2579);
nor U2609 (N_2609,N_2583,N_2552);
or U2610 (N_2610,N_2576,N_2506);
xnor U2611 (N_2611,N_2507,N_2532);
xnor U2612 (N_2612,N_2533,N_2522);
nand U2613 (N_2613,N_2539,N_2513);
xnor U2614 (N_2614,N_2519,N_2596);
nor U2615 (N_2615,N_2589,N_2582);
or U2616 (N_2616,N_2547,N_2570);
nor U2617 (N_2617,N_2501,N_2590);
nand U2618 (N_2618,N_2593,N_2564);
nand U2619 (N_2619,N_2568,N_2521);
nand U2620 (N_2620,N_2554,N_2580);
or U2621 (N_2621,N_2536,N_2550);
or U2622 (N_2622,N_2502,N_2581);
nor U2623 (N_2623,N_2598,N_2571);
xnor U2624 (N_2624,N_2561,N_2577);
nor U2625 (N_2625,N_2597,N_2540);
xnor U2626 (N_2626,N_2537,N_2531);
or U2627 (N_2627,N_2505,N_2574);
nor U2628 (N_2628,N_2553,N_2594);
nor U2629 (N_2629,N_2563,N_2557);
and U2630 (N_2630,N_2509,N_2592);
xor U2631 (N_2631,N_2575,N_2587);
xor U2632 (N_2632,N_2514,N_2503);
nor U2633 (N_2633,N_2525,N_2595);
and U2634 (N_2634,N_2591,N_2512);
nor U2635 (N_2635,N_2527,N_2588);
and U2636 (N_2636,N_2566,N_2560);
xnor U2637 (N_2637,N_2534,N_2558);
nor U2638 (N_2638,N_2584,N_2585);
and U2639 (N_2639,N_2526,N_2510);
or U2640 (N_2640,N_2549,N_2546);
nor U2641 (N_2641,N_2523,N_2500);
nor U2642 (N_2642,N_2599,N_2543);
or U2643 (N_2643,N_2515,N_2511);
or U2644 (N_2644,N_2524,N_2565);
nand U2645 (N_2645,N_2572,N_2529);
and U2646 (N_2646,N_2517,N_2545);
nand U2647 (N_2647,N_2520,N_2548);
xor U2648 (N_2648,N_2556,N_2555);
or U2649 (N_2649,N_2518,N_2567);
or U2650 (N_2650,N_2573,N_2590);
xor U2651 (N_2651,N_2532,N_2596);
and U2652 (N_2652,N_2509,N_2523);
or U2653 (N_2653,N_2541,N_2592);
nand U2654 (N_2654,N_2536,N_2598);
nand U2655 (N_2655,N_2581,N_2538);
or U2656 (N_2656,N_2585,N_2527);
and U2657 (N_2657,N_2512,N_2586);
nor U2658 (N_2658,N_2530,N_2586);
nor U2659 (N_2659,N_2567,N_2548);
and U2660 (N_2660,N_2573,N_2595);
and U2661 (N_2661,N_2534,N_2583);
and U2662 (N_2662,N_2540,N_2594);
nor U2663 (N_2663,N_2537,N_2577);
xor U2664 (N_2664,N_2573,N_2580);
nand U2665 (N_2665,N_2500,N_2501);
and U2666 (N_2666,N_2524,N_2584);
xor U2667 (N_2667,N_2567,N_2527);
nand U2668 (N_2668,N_2506,N_2502);
xnor U2669 (N_2669,N_2521,N_2561);
and U2670 (N_2670,N_2596,N_2504);
nor U2671 (N_2671,N_2579,N_2561);
nor U2672 (N_2672,N_2558,N_2567);
nand U2673 (N_2673,N_2564,N_2590);
xnor U2674 (N_2674,N_2533,N_2521);
xor U2675 (N_2675,N_2593,N_2538);
and U2676 (N_2676,N_2518,N_2515);
nand U2677 (N_2677,N_2527,N_2596);
and U2678 (N_2678,N_2544,N_2580);
and U2679 (N_2679,N_2500,N_2557);
and U2680 (N_2680,N_2534,N_2545);
or U2681 (N_2681,N_2531,N_2505);
or U2682 (N_2682,N_2543,N_2526);
and U2683 (N_2683,N_2546,N_2543);
nor U2684 (N_2684,N_2520,N_2578);
and U2685 (N_2685,N_2569,N_2524);
and U2686 (N_2686,N_2575,N_2539);
nand U2687 (N_2687,N_2522,N_2505);
nand U2688 (N_2688,N_2599,N_2577);
nand U2689 (N_2689,N_2544,N_2540);
nand U2690 (N_2690,N_2550,N_2500);
xor U2691 (N_2691,N_2578,N_2583);
xor U2692 (N_2692,N_2569,N_2577);
and U2693 (N_2693,N_2514,N_2557);
xor U2694 (N_2694,N_2568,N_2551);
nor U2695 (N_2695,N_2520,N_2509);
xor U2696 (N_2696,N_2564,N_2560);
nor U2697 (N_2697,N_2571,N_2537);
xor U2698 (N_2698,N_2584,N_2563);
nand U2699 (N_2699,N_2538,N_2522);
xnor U2700 (N_2700,N_2641,N_2613);
nor U2701 (N_2701,N_2648,N_2696);
nor U2702 (N_2702,N_2658,N_2630);
nand U2703 (N_2703,N_2697,N_2656);
nor U2704 (N_2704,N_2603,N_2633);
or U2705 (N_2705,N_2614,N_2672);
and U2706 (N_2706,N_2654,N_2622);
and U2707 (N_2707,N_2615,N_2694);
nor U2708 (N_2708,N_2651,N_2604);
nand U2709 (N_2709,N_2608,N_2660);
and U2710 (N_2710,N_2634,N_2682);
and U2711 (N_2711,N_2629,N_2670);
xnor U2712 (N_2712,N_2671,N_2624);
and U2713 (N_2713,N_2665,N_2681);
nor U2714 (N_2714,N_2606,N_2684);
nor U2715 (N_2715,N_2695,N_2659);
nor U2716 (N_2716,N_2657,N_2626);
and U2717 (N_2717,N_2668,N_2649);
xnor U2718 (N_2718,N_2647,N_2685);
nor U2719 (N_2719,N_2616,N_2643);
nand U2720 (N_2720,N_2644,N_2688);
or U2721 (N_2721,N_2652,N_2601);
or U2722 (N_2722,N_2687,N_2605);
nor U2723 (N_2723,N_2664,N_2617);
xor U2724 (N_2724,N_2683,N_2698);
xor U2725 (N_2725,N_2669,N_2632);
nand U2726 (N_2726,N_2693,N_2636);
nor U2727 (N_2727,N_2607,N_2686);
xnor U2728 (N_2728,N_2610,N_2642);
and U2729 (N_2729,N_2663,N_2655);
and U2730 (N_2730,N_2666,N_2677);
nor U2731 (N_2731,N_2646,N_2653);
xnor U2732 (N_2732,N_2675,N_2692);
xor U2733 (N_2733,N_2667,N_2627);
nor U2734 (N_2734,N_2635,N_2650);
nor U2735 (N_2735,N_2625,N_2619);
nand U2736 (N_2736,N_2640,N_2618);
xor U2737 (N_2737,N_2674,N_2637);
or U2738 (N_2738,N_2611,N_2621);
nand U2739 (N_2739,N_2691,N_2678);
xnor U2740 (N_2740,N_2623,N_2600);
nand U2741 (N_2741,N_2638,N_2602);
or U2742 (N_2742,N_2680,N_2662);
or U2743 (N_2743,N_2645,N_2690);
nor U2744 (N_2744,N_2661,N_2620);
nand U2745 (N_2745,N_2612,N_2679);
nand U2746 (N_2746,N_2628,N_2639);
nor U2747 (N_2747,N_2699,N_2673);
or U2748 (N_2748,N_2676,N_2689);
or U2749 (N_2749,N_2609,N_2631);
and U2750 (N_2750,N_2615,N_2647);
xnor U2751 (N_2751,N_2644,N_2695);
and U2752 (N_2752,N_2685,N_2626);
nand U2753 (N_2753,N_2623,N_2698);
or U2754 (N_2754,N_2639,N_2652);
xnor U2755 (N_2755,N_2622,N_2625);
nand U2756 (N_2756,N_2630,N_2666);
nor U2757 (N_2757,N_2692,N_2644);
nand U2758 (N_2758,N_2691,N_2681);
and U2759 (N_2759,N_2688,N_2659);
xor U2760 (N_2760,N_2632,N_2604);
and U2761 (N_2761,N_2679,N_2690);
nand U2762 (N_2762,N_2648,N_2609);
and U2763 (N_2763,N_2626,N_2617);
or U2764 (N_2764,N_2610,N_2608);
nor U2765 (N_2765,N_2618,N_2664);
nand U2766 (N_2766,N_2662,N_2623);
nand U2767 (N_2767,N_2601,N_2643);
nor U2768 (N_2768,N_2677,N_2620);
and U2769 (N_2769,N_2612,N_2675);
and U2770 (N_2770,N_2634,N_2613);
and U2771 (N_2771,N_2682,N_2608);
and U2772 (N_2772,N_2654,N_2690);
and U2773 (N_2773,N_2664,N_2637);
xnor U2774 (N_2774,N_2648,N_2670);
nor U2775 (N_2775,N_2610,N_2635);
nor U2776 (N_2776,N_2696,N_2685);
or U2777 (N_2777,N_2691,N_2612);
xor U2778 (N_2778,N_2616,N_2699);
nand U2779 (N_2779,N_2660,N_2646);
xor U2780 (N_2780,N_2621,N_2623);
and U2781 (N_2781,N_2661,N_2652);
xor U2782 (N_2782,N_2686,N_2630);
and U2783 (N_2783,N_2651,N_2643);
xor U2784 (N_2784,N_2693,N_2609);
or U2785 (N_2785,N_2617,N_2676);
nor U2786 (N_2786,N_2621,N_2615);
nand U2787 (N_2787,N_2694,N_2619);
or U2788 (N_2788,N_2604,N_2683);
nor U2789 (N_2789,N_2636,N_2652);
or U2790 (N_2790,N_2646,N_2601);
and U2791 (N_2791,N_2615,N_2657);
and U2792 (N_2792,N_2676,N_2660);
or U2793 (N_2793,N_2657,N_2662);
nor U2794 (N_2794,N_2687,N_2607);
nor U2795 (N_2795,N_2656,N_2616);
xor U2796 (N_2796,N_2618,N_2685);
nor U2797 (N_2797,N_2663,N_2657);
nand U2798 (N_2798,N_2679,N_2630);
nand U2799 (N_2799,N_2635,N_2638);
and U2800 (N_2800,N_2704,N_2791);
and U2801 (N_2801,N_2734,N_2721);
xor U2802 (N_2802,N_2788,N_2797);
and U2803 (N_2803,N_2723,N_2781);
nor U2804 (N_2804,N_2722,N_2768);
or U2805 (N_2805,N_2758,N_2727);
xnor U2806 (N_2806,N_2700,N_2799);
nand U2807 (N_2807,N_2772,N_2708);
nand U2808 (N_2808,N_2713,N_2787);
or U2809 (N_2809,N_2728,N_2779);
xor U2810 (N_2810,N_2756,N_2754);
xor U2811 (N_2811,N_2798,N_2729);
and U2812 (N_2812,N_2715,N_2706);
nand U2813 (N_2813,N_2751,N_2710);
or U2814 (N_2814,N_2794,N_2744);
xor U2815 (N_2815,N_2764,N_2720);
nand U2816 (N_2816,N_2741,N_2780);
nand U2817 (N_2817,N_2748,N_2725);
nand U2818 (N_2818,N_2765,N_2774);
and U2819 (N_2819,N_2757,N_2735);
or U2820 (N_2820,N_2709,N_2712);
nand U2821 (N_2821,N_2777,N_2739);
xnor U2822 (N_2822,N_2778,N_2753);
nand U2823 (N_2823,N_2747,N_2782);
and U2824 (N_2824,N_2743,N_2795);
nand U2825 (N_2825,N_2724,N_2752);
xnor U2826 (N_2826,N_2784,N_2783);
nor U2827 (N_2827,N_2755,N_2786);
xnor U2828 (N_2828,N_2759,N_2726);
or U2829 (N_2829,N_2796,N_2750);
xor U2830 (N_2830,N_2730,N_2738);
nor U2831 (N_2831,N_2760,N_2707);
and U2832 (N_2832,N_2731,N_2773);
nor U2833 (N_2833,N_2771,N_2711);
nand U2834 (N_2834,N_2716,N_2732);
or U2835 (N_2835,N_2746,N_2703);
xor U2836 (N_2836,N_2776,N_2717);
or U2837 (N_2837,N_2736,N_2719);
and U2838 (N_2838,N_2718,N_2766);
and U2839 (N_2839,N_2767,N_2762);
nor U2840 (N_2840,N_2733,N_2785);
nor U2841 (N_2841,N_2702,N_2749);
and U2842 (N_2842,N_2705,N_2742);
and U2843 (N_2843,N_2770,N_2789);
nand U2844 (N_2844,N_2790,N_2701);
nand U2845 (N_2845,N_2763,N_2769);
nand U2846 (N_2846,N_2714,N_2761);
and U2847 (N_2847,N_2775,N_2792);
nand U2848 (N_2848,N_2793,N_2745);
nand U2849 (N_2849,N_2740,N_2737);
or U2850 (N_2850,N_2710,N_2760);
xor U2851 (N_2851,N_2744,N_2743);
and U2852 (N_2852,N_2798,N_2797);
xor U2853 (N_2853,N_2731,N_2766);
or U2854 (N_2854,N_2781,N_2737);
nand U2855 (N_2855,N_2757,N_2766);
or U2856 (N_2856,N_2772,N_2741);
and U2857 (N_2857,N_2753,N_2772);
and U2858 (N_2858,N_2741,N_2795);
nor U2859 (N_2859,N_2718,N_2736);
nand U2860 (N_2860,N_2702,N_2757);
or U2861 (N_2861,N_2718,N_2710);
xor U2862 (N_2862,N_2755,N_2732);
and U2863 (N_2863,N_2751,N_2785);
nand U2864 (N_2864,N_2767,N_2737);
and U2865 (N_2865,N_2736,N_2712);
xnor U2866 (N_2866,N_2737,N_2725);
or U2867 (N_2867,N_2780,N_2716);
or U2868 (N_2868,N_2701,N_2785);
and U2869 (N_2869,N_2717,N_2790);
nor U2870 (N_2870,N_2744,N_2766);
nor U2871 (N_2871,N_2777,N_2748);
xnor U2872 (N_2872,N_2722,N_2708);
nand U2873 (N_2873,N_2726,N_2781);
nor U2874 (N_2874,N_2791,N_2759);
xnor U2875 (N_2875,N_2796,N_2797);
or U2876 (N_2876,N_2742,N_2708);
nor U2877 (N_2877,N_2709,N_2703);
nand U2878 (N_2878,N_2773,N_2786);
nand U2879 (N_2879,N_2753,N_2716);
xor U2880 (N_2880,N_2740,N_2704);
or U2881 (N_2881,N_2788,N_2721);
or U2882 (N_2882,N_2789,N_2772);
nor U2883 (N_2883,N_2772,N_2760);
nor U2884 (N_2884,N_2779,N_2787);
or U2885 (N_2885,N_2778,N_2700);
nand U2886 (N_2886,N_2770,N_2733);
xnor U2887 (N_2887,N_2740,N_2713);
xnor U2888 (N_2888,N_2776,N_2760);
xnor U2889 (N_2889,N_2702,N_2796);
or U2890 (N_2890,N_2760,N_2733);
nand U2891 (N_2891,N_2711,N_2730);
and U2892 (N_2892,N_2716,N_2777);
nor U2893 (N_2893,N_2778,N_2761);
nor U2894 (N_2894,N_2720,N_2778);
nor U2895 (N_2895,N_2725,N_2762);
xor U2896 (N_2896,N_2795,N_2739);
nand U2897 (N_2897,N_2745,N_2712);
nor U2898 (N_2898,N_2738,N_2791);
nand U2899 (N_2899,N_2747,N_2772);
or U2900 (N_2900,N_2819,N_2873);
or U2901 (N_2901,N_2892,N_2861);
xnor U2902 (N_2902,N_2804,N_2838);
xor U2903 (N_2903,N_2826,N_2832);
or U2904 (N_2904,N_2863,N_2836);
xor U2905 (N_2905,N_2834,N_2806);
nand U2906 (N_2906,N_2866,N_2825);
or U2907 (N_2907,N_2855,N_2850);
nor U2908 (N_2908,N_2817,N_2833);
xnor U2909 (N_2909,N_2829,N_2800);
nor U2910 (N_2910,N_2827,N_2824);
and U2911 (N_2911,N_2860,N_2883);
nor U2912 (N_2912,N_2835,N_2816);
and U2913 (N_2913,N_2812,N_2823);
xor U2914 (N_2914,N_2805,N_2875);
and U2915 (N_2915,N_2813,N_2888);
and U2916 (N_2916,N_2881,N_2877);
and U2917 (N_2917,N_2842,N_2871);
and U2918 (N_2918,N_2899,N_2845);
nand U2919 (N_2919,N_2814,N_2895);
nor U2920 (N_2920,N_2885,N_2803);
or U2921 (N_2921,N_2821,N_2893);
or U2922 (N_2922,N_2839,N_2851);
nor U2923 (N_2923,N_2856,N_2894);
xnor U2924 (N_2924,N_2882,N_2862);
nand U2925 (N_2925,N_2808,N_2849);
nand U2926 (N_2926,N_2859,N_2870);
nand U2927 (N_2927,N_2874,N_2865);
nor U2928 (N_2928,N_2879,N_2828);
and U2929 (N_2929,N_2841,N_2853);
or U2930 (N_2930,N_2844,N_2815);
and U2931 (N_2931,N_2872,N_2848);
and U2932 (N_2932,N_2846,N_2847);
nor U2933 (N_2933,N_2852,N_2810);
and U2934 (N_2934,N_2897,N_2887);
nor U2935 (N_2935,N_2898,N_2889);
nor U2936 (N_2936,N_2890,N_2822);
and U2937 (N_2937,N_2857,N_2811);
nand U2938 (N_2938,N_2867,N_2830);
and U2939 (N_2939,N_2818,N_2868);
xor U2940 (N_2940,N_2864,N_2831);
and U2941 (N_2941,N_2809,N_2807);
or U2942 (N_2942,N_2854,N_2858);
nor U2943 (N_2943,N_2878,N_2843);
or U2944 (N_2944,N_2876,N_2840);
nand U2945 (N_2945,N_2801,N_2802);
nor U2946 (N_2946,N_2884,N_2837);
xor U2947 (N_2947,N_2896,N_2869);
and U2948 (N_2948,N_2880,N_2820);
and U2949 (N_2949,N_2891,N_2886);
or U2950 (N_2950,N_2869,N_2846);
nor U2951 (N_2951,N_2846,N_2858);
nor U2952 (N_2952,N_2898,N_2821);
xor U2953 (N_2953,N_2827,N_2804);
nand U2954 (N_2954,N_2841,N_2875);
xor U2955 (N_2955,N_2892,N_2822);
nand U2956 (N_2956,N_2837,N_2858);
nor U2957 (N_2957,N_2874,N_2805);
and U2958 (N_2958,N_2840,N_2828);
or U2959 (N_2959,N_2827,N_2805);
xnor U2960 (N_2960,N_2871,N_2810);
nand U2961 (N_2961,N_2880,N_2870);
and U2962 (N_2962,N_2859,N_2874);
nor U2963 (N_2963,N_2820,N_2857);
nand U2964 (N_2964,N_2862,N_2836);
nor U2965 (N_2965,N_2824,N_2802);
nand U2966 (N_2966,N_2888,N_2829);
or U2967 (N_2967,N_2844,N_2871);
nor U2968 (N_2968,N_2863,N_2855);
and U2969 (N_2969,N_2845,N_2826);
xor U2970 (N_2970,N_2811,N_2876);
nand U2971 (N_2971,N_2845,N_2828);
and U2972 (N_2972,N_2813,N_2894);
and U2973 (N_2973,N_2876,N_2870);
nand U2974 (N_2974,N_2813,N_2805);
xnor U2975 (N_2975,N_2892,N_2881);
xnor U2976 (N_2976,N_2867,N_2891);
nand U2977 (N_2977,N_2898,N_2813);
or U2978 (N_2978,N_2813,N_2881);
and U2979 (N_2979,N_2897,N_2806);
nor U2980 (N_2980,N_2878,N_2816);
and U2981 (N_2981,N_2881,N_2885);
and U2982 (N_2982,N_2896,N_2871);
nand U2983 (N_2983,N_2850,N_2892);
and U2984 (N_2984,N_2893,N_2862);
nand U2985 (N_2985,N_2852,N_2842);
xor U2986 (N_2986,N_2844,N_2860);
nand U2987 (N_2987,N_2823,N_2836);
nand U2988 (N_2988,N_2820,N_2835);
xnor U2989 (N_2989,N_2870,N_2812);
xnor U2990 (N_2990,N_2827,N_2816);
nand U2991 (N_2991,N_2866,N_2897);
or U2992 (N_2992,N_2879,N_2813);
nand U2993 (N_2993,N_2829,N_2862);
nand U2994 (N_2994,N_2802,N_2841);
nand U2995 (N_2995,N_2843,N_2865);
nor U2996 (N_2996,N_2864,N_2840);
and U2997 (N_2997,N_2856,N_2845);
nand U2998 (N_2998,N_2823,N_2828);
or U2999 (N_2999,N_2816,N_2826);
and U3000 (N_3000,N_2993,N_2935);
or U3001 (N_3001,N_2937,N_2907);
xnor U3002 (N_3002,N_2920,N_2951);
and U3003 (N_3003,N_2917,N_2979);
or U3004 (N_3004,N_2909,N_2938);
xnor U3005 (N_3005,N_2973,N_2959);
xnor U3006 (N_3006,N_2901,N_2911);
or U3007 (N_3007,N_2903,N_2918);
xor U3008 (N_3008,N_2966,N_2980);
and U3009 (N_3009,N_2957,N_2974);
xnor U3010 (N_3010,N_2900,N_2978);
nand U3011 (N_3011,N_2945,N_2949);
nand U3012 (N_3012,N_2961,N_2924);
or U3013 (N_3013,N_2997,N_2971);
or U3014 (N_3014,N_2926,N_2929);
nor U3015 (N_3015,N_2915,N_2950);
and U3016 (N_3016,N_2994,N_2941);
xnor U3017 (N_3017,N_2912,N_2932);
xor U3018 (N_3018,N_2972,N_2928);
xnor U3019 (N_3019,N_2925,N_2962);
and U3020 (N_3020,N_2944,N_2977);
nand U3021 (N_3021,N_2967,N_2914);
and U3022 (N_3022,N_2958,N_2981);
nor U3023 (N_3023,N_2999,N_2975);
nand U3024 (N_3024,N_2948,N_2908);
nand U3025 (N_3025,N_2947,N_2998);
nand U3026 (N_3026,N_2939,N_2969);
or U3027 (N_3027,N_2990,N_2919);
or U3028 (N_3028,N_2982,N_2905);
nand U3029 (N_3029,N_2984,N_2988);
nor U3030 (N_3030,N_2934,N_2970);
nand U3031 (N_3031,N_2933,N_2946);
xor U3032 (N_3032,N_2976,N_2921);
xnor U3033 (N_3033,N_2960,N_2916);
or U3034 (N_3034,N_2952,N_2983);
and U3035 (N_3035,N_2904,N_2954);
xor U3036 (N_3036,N_2913,N_2953);
xor U3037 (N_3037,N_2930,N_2910);
xor U3038 (N_3038,N_2922,N_2931);
xor U3039 (N_3039,N_2989,N_2943);
nor U3040 (N_3040,N_2906,N_2956);
xnor U3041 (N_3041,N_2995,N_2902);
xnor U3042 (N_3042,N_2986,N_2965);
xnor U3043 (N_3043,N_2923,N_2992);
nor U3044 (N_3044,N_2955,N_2991);
xnor U3045 (N_3045,N_2996,N_2968);
and U3046 (N_3046,N_2927,N_2942);
or U3047 (N_3047,N_2936,N_2987);
nand U3048 (N_3048,N_2940,N_2963);
xor U3049 (N_3049,N_2964,N_2985);
nor U3050 (N_3050,N_2945,N_2985);
and U3051 (N_3051,N_2968,N_2953);
nor U3052 (N_3052,N_2905,N_2993);
and U3053 (N_3053,N_2932,N_2936);
nor U3054 (N_3054,N_2945,N_2926);
and U3055 (N_3055,N_2907,N_2933);
xor U3056 (N_3056,N_2908,N_2930);
xor U3057 (N_3057,N_2916,N_2947);
nor U3058 (N_3058,N_2936,N_2912);
xor U3059 (N_3059,N_2997,N_2915);
nor U3060 (N_3060,N_2903,N_2945);
or U3061 (N_3061,N_2946,N_2988);
xor U3062 (N_3062,N_2946,N_2919);
and U3063 (N_3063,N_2931,N_2945);
xor U3064 (N_3064,N_2902,N_2932);
and U3065 (N_3065,N_2943,N_2931);
or U3066 (N_3066,N_2921,N_2998);
nor U3067 (N_3067,N_2998,N_2927);
or U3068 (N_3068,N_2985,N_2918);
or U3069 (N_3069,N_2958,N_2961);
and U3070 (N_3070,N_2965,N_2942);
or U3071 (N_3071,N_2935,N_2919);
nor U3072 (N_3072,N_2909,N_2976);
nand U3073 (N_3073,N_2993,N_2901);
xnor U3074 (N_3074,N_2984,N_2900);
nand U3075 (N_3075,N_2917,N_2975);
xnor U3076 (N_3076,N_2987,N_2946);
or U3077 (N_3077,N_2920,N_2937);
nor U3078 (N_3078,N_2967,N_2995);
xnor U3079 (N_3079,N_2908,N_2958);
nor U3080 (N_3080,N_2988,N_2909);
xor U3081 (N_3081,N_2930,N_2953);
and U3082 (N_3082,N_2976,N_2999);
and U3083 (N_3083,N_2903,N_2935);
or U3084 (N_3084,N_2923,N_2998);
or U3085 (N_3085,N_2958,N_2925);
xnor U3086 (N_3086,N_2908,N_2993);
nor U3087 (N_3087,N_2992,N_2935);
and U3088 (N_3088,N_2968,N_2949);
or U3089 (N_3089,N_2913,N_2946);
nand U3090 (N_3090,N_2908,N_2934);
nand U3091 (N_3091,N_2953,N_2905);
nor U3092 (N_3092,N_2969,N_2979);
and U3093 (N_3093,N_2928,N_2996);
nand U3094 (N_3094,N_2931,N_2902);
nand U3095 (N_3095,N_2967,N_2989);
nor U3096 (N_3096,N_2931,N_2981);
xnor U3097 (N_3097,N_2915,N_2963);
nand U3098 (N_3098,N_2951,N_2981);
or U3099 (N_3099,N_2965,N_2932);
nand U3100 (N_3100,N_3033,N_3026);
xnor U3101 (N_3101,N_3061,N_3097);
nor U3102 (N_3102,N_3057,N_3081);
nand U3103 (N_3103,N_3018,N_3087);
xnor U3104 (N_3104,N_3086,N_3085);
xor U3105 (N_3105,N_3049,N_3054);
or U3106 (N_3106,N_3064,N_3059);
and U3107 (N_3107,N_3052,N_3005);
and U3108 (N_3108,N_3007,N_3040);
nand U3109 (N_3109,N_3088,N_3084);
xor U3110 (N_3110,N_3060,N_3068);
xnor U3111 (N_3111,N_3021,N_3048);
nand U3112 (N_3112,N_3069,N_3014);
xnor U3113 (N_3113,N_3053,N_3055);
nand U3114 (N_3114,N_3001,N_3082);
nand U3115 (N_3115,N_3029,N_3056);
and U3116 (N_3116,N_3028,N_3091);
nand U3117 (N_3117,N_3000,N_3076);
or U3118 (N_3118,N_3078,N_3070);
or U3119 (N_3119,N_3008,N_3047);
and U3120 (N_3120,N_3023,N_3094);
nor U3121 (N_3121,N_3031,N_3051);
xor U3122 (N_3122,N_3024,N_3046);
nand U3123 (N_3123,N_3090,N_3043);
or U3124 (N_3124,N_3067,N_3062);
or U3125 (N_3125,N_3095,N_3071);
or U3126 (N_3126,N_3025,N_3027);
or U3127 (N_3127,N_3022,N_3039);
and U3128 (N_3128,N_3017,N_3019);
xnor U3129 (N_3129,N_3063,N_3073);
xnor U3130 (N_3130,N_3016,N_3009);
nand U3131 (N_3131,N_3020,N_3050);
nor U3132 (N_3132,N_3012,N_3099);
or U3133 (N_3133,N_3036,N_3030);
nor U3134 (N_3134,N_3006,N_3011);
nand U3135 (N_3135,N_3002,N_3044);
or U3136 (N_3136,N_3066,N_3080);
nand U3137 (N_3137,N_3035,N_3092);
nor U3138 (N_3138,N_3010,N_3037);
and U3139 (N_3139,N_3032,N_3074);
or U3140 (N_3140,N_3072,N_3075);
xnor U3141 (N_3141,N_3083,N_3004);
nor U3142 (N_3142,N_3077,N_3003);
or U3143 (N_3143,N_3041,N_3058);
nor U3144 (N_3144,N_3098,N_3015);
and U3145 (N_3145,N_3045,N_3065);
nand U3146 (N_3146,N_3079,N_3038);
nand U3147 (N_3147,N_3034,N_3096);
xnor U3148 (N_3148,N_3089,N_3013);
nand U3149 (N_3149,N_3042,N_3093);
nand U3150 (N_3150,N_3007,N_3016);
or U3151 (N_3151,N_3021,N_3018);
and U3152 (N_3152,N_3053,N_3015);
xnor U3153 (N_3153,N_3062,N_3080);
nor U3154 (N_3154,N_3074,N_3093);
nor U3155 (N_3155,N_3025,N_3088);
and U3156 (N_3156,N_3091,N_3096);
nand U3157 (N_3157,N_3065,N_3057);
xor U3158 (N_3158,N_3094,N_3071);
nand U3159 (N_3159,N_3081,N_3074);
xnor U3160 (N_3160,N_3099,N_3091);
nand U3161 (N_3161,N_3079,N_3064);
and U3162 (N_3162,N_3057,N_3041);
nand U3163 (N_3163,N_3094,N_3051);
nor U3164 (N_3164,N_3087,N_3017);
or U3165 (N_3165,N_3027,N_3060);
and U3166 (N_3166,N_3026,N_3013);
and U3167 (N_3167,N_3087,N_3032);
xor U3168 (N_3168,N_3067,N_3037);
xnor U3169 (N_3169,N_3036,N_3046);
and U3170 (N_3170,N_3090,N_3080);
nor U3171 (N_3171,N_3021,N_3054);
nor U3172 (N_3172,N_3040,N_3054);
nand U3173 (N_3173,N_3062,N_3034);
nand U3174 (N_3174,N_3078,N_3033);
nor U3175 (N_3175,N_3050,N_3078);
nand U3176 (N_3176,N_3097,N_3091);
nor U3177 (N_3177,N_3052,N_3057);
xnor U3178 (N_3178,N_3074,N_3070);
nor U3179 (N_3179,N_3087,N_3091);
or U3180 (N_3180,N_3073,N_3086);
nor U3181 (N_3181,N_3014,N_3030);
and U3182 (N_3182,N_3082,N_3015);
nor U3183 (N_3183,N_3082,N_3004);
nand U3184 (N_3184,N_3099,N_3085);
or U3185 (N_3185,N_3090,N_3047);
nor U3186 (N_3186,N_3085,N_3027);
or U3187 (N_3187,N_3004,N_3065);
xnor U3188 (N_3188,N_3028,N_3030);
nand U3189 (N_3189,N_3034,N_3037);
nor U3190 (N_3190,N_3009,N_3062);
or U3191 (N_3191,N_3098,N_3086);
nand U3192 (N_3192,N_3069,N_3009);
nor U3193 (N_3193,N_3000,N_3063);
xor U3194 (N_3194,N_3031,N_3026);
and U3195 (N_3195,N_3038,N_3037);
nor U3196 (N_3196,N_3094,N_3016);
xnor U3197 (N_3197,N_3026,N_3054);
or U3198 (N_3198,N_3018,N_3016);
xor U3199 (N_3199,N_3079,N_3026);
or U3200 (N_3200,N_3124,N_3123);
and U3201 (N_3201,N_3175,N_3153);
nor U3202 (N_3202,N_3146,N_3167);
xor U3203 (N_3203,N_3177,N_3154);
nand U3204 (N_3204,N_3162,N_3188);
xor U3205 (N_3205,N_3144,N_3158);
nand U3206 (N_3206,N_3134,N_3117);
and U3207 (N_3207,N_3184,N_3130);
or U3208 (N_3208,N_3190,N_3108);
nand U3209 (N_3209,N_3139,N_3186);
or U3210 (N_3210,N_3121,N_3129);
or U3211 (N_3211,N_3128,N_3161);
nor U3212 (N_3212,N_3169,N_3142);
nor U3213 (N_3213,N_3170,N_3189);
nand U3214 (N_3214,N_3152,N_3166);
and U3215 (N_3215,N_3187,N_3103);
nand U3216 (N_3216,N_3197,N_3172);
nor U3217 (N_3217,N_3136,N_3131);
or U3218 (N_3218,N_3122,N_3173);
nor U3219 (N_3219,N_3183,N_3176);
or U3220 (N_3220,N_3126,N_3198);
xor U3221 (N_3221,N_3148,N_3137);
or U3222 (N_3222,N_3157,N_3192);
and U3223 (N_3223,N_3151,N_3109);
or U3224 (N_3224,N_3111,N_3182);
nand U3225 (N_3225,N_3181,N_3135);
nand U3226 (N_3226,N_3195,N_3138);
xnor U3227 (N_3227,N_3194,N_3106);
xnor U3228 (N_3228,N_3110,N_3143);
or U3229 (N_3229,N_3133,N_3163);
and U3230 (N_3230,N_3105,N_3141);
or U3231 (N_3231,N_3101,N_3116);
nor U3232 (N_3232,N_3191,N_3164);
and U3233 (N_3233,N_3193,N_3145);
nor U3234 (N_3234,N_3171,N_3119);
xor U3235 (N_3235,N_3125,N_3165);
or U3236 (N_3236,N_3160,N_3113);
and U3237 (N_3237,N_3132,N_3199);
and U3238 (N_3238,N_3156,N_3149);
xor U3239 (N_3239,N_3114,N_3150);
nand U3240 (N_3240,N_3155,N_3196);
xor U3241 (N_3241,N_3112,N_3127);
and U3242 (N_3242,N_3178,N_3120);
and U3243 (N_3243,N_3180,N_3118);
and U3244 (N_3244,N_3159,N_3115);
nor U3245 (N_3245,N_3104,N_3100);
nor U3246 (N_3246,N_3179,N_3174);
or U3247 (N_3247,N_3147,N_3102);
nand U3248 (N_3248,N_3107,N_3140);
and U3249 (N_3249,N_3185,N_3168);
and U3250 (N_3250,N_3170,N_3169);
nand U3251 (N_3251,N_3155,N_3172);
xnor U3252 (N_3252,N_3147,N_3131);
nand U3253 (N_3253,N_3159,N_3130);
or U3254 (N_3254,N_3143,N_3166);
nor U3255 (N_3255,N_3101,N_3121);
nand U3256 (N_3256,N_3144,N_3166);
and U3257 (N_3257,N_3195,N_3111);
nand U3258 (N_3258,N_3186,N_3128);
nand U3259 (N_3259,N_3147,N_3150);
nor U3260 (N_3260,N_3198,N_3114);
or U3261 (N_3261,N_3142,N_3127);
nor U3262 (N_3262,N_3163,N_3134);
nor U3263 (N_3263,N_3144,N_3197);
nand U3264 (N_3264,N_3188,N_3103);
and U3265 (N_3265,N_3189,N_3123);
xor U3266 (N_3266,N_3102,N_3107);
and U3267 (N_3267,N_3184,N_3191);
or U3268 (N_3268,N_3109,N_3164);
and U3269 (N_3269,N_3143,N_3161);
nor U3270 (N_3270,N_3140,N_3146);
nand U3271 (N_3271,N_3157,N_3111);
xnor U3272 (N_3272,N_3139,N_3101);
or U3273 (N_3273,N_3164,N_3126);
or U3274 (N_3274,N_3111,N_3135);
nand U3275 (N_3275,N_3133,N_3132);
and U3276 (N_3276,N_3105,N_3111);
xnor U3277 (N_3277,N_3178,N_3194);
or U3278 (N_3278,N_3139,N_3140);
or U3279 (N_3279,N_3189,N_3181);
or U3280 (N_3280,N_3198,N_3131);
and U3281 (N_3281,N_3150,N_3101);
nor U3282 (N_3282,N_3162,N_3167);
nand U3283 (N_3283,N_3188,N_3107);
and U3284 (N_3284,N_3174,N_3158);
or U3285 (N_3285,N_3154,N_3110);
nor U3286 (N_3286,N_3160,N_3112);
nor U3287 (N_3287,N_3149,N_3168);
nor U3288 (N_3288,N_3164,N_3122);
or U3289 (N_3289,N_3135,N_3110);
or U3290 (N_3290,N_3186,N_3175);
nor U3291 (N_3291,N_3153,N_3135);
or U3292 (N_3292,N_3186,N_3111);
xor U3293 (N_3293,N_3197,N_3195);
or U3294 (N_3294,N_3198,N_3121);
nor U3295 (N_3295,N_3185,N_3184);
nand U3296 (N_3296,N_3116,N_3107);
or U3297 (N_3297,N_3103,N_3135);
nand U3298 (N_3298,N_3105,N_3183);
nor U3299 (N_3299,N_3113,N_3157);
and U3300 (N_3300,N_3232,N_3211);
nor U3301 (N_3301,N_3231,N_3261);
or U3302 (N_3302,N_3205,N_3204);
and U3303 (N_3303,N_3296,N_3244);
nand U3304 (N_3304,N_3268,N_3215);
nor U3305 (N_3305,N_3285,N_3280);
nand U3306 (N_3306,N_3256,N_3259);
nand U3307 (N_3307,N_3288,N_3284);
nor U3308 (N_3308,N_3247,N_3218);
or U3309 (N_3309,N_3200,N_3295);
or U3310 (N_3310,N_3254,N_3278);
nand U3311 (N_3311,N_3283,N_3286);
nor U3312 (N_3312,N_3269,N_3212);
xor U3313 (N_3313,N_3248,N_3226);
and U3314 (N_3314,N_3209,N_3263);
nor U3315 (N_3315,N_3237,N_3234);
and U3316 (N_3316,N_3277,N_3238);
nand U3317 (N_3317,N_3281,N_3274);
or U3318 (N_3318,N_3233,N_3293);
or U3319 (N_3319,N_3279,N_3221);
nand U3320 (N_3320,N_3250,N_3219);
and U3321 (N_3321,N_3236,N_3207);
nor U3322 (N_3322,N_3216,N_3217);
nand U3323 (N_3323,N_3242,N_3294);
or U3324 (N_3324,N_3223,N_3297);
xnor U3325 (N_3325,N_3246,N_3228);
and U3326 (N_3326,N_3298,N_3257);
or U3327 (N_3327,N_3255,N_3210);
and U3328 (N_3328,N_3276,N_3271);
xnor U3329 (N_3329,N_3273,N_3222);
nor U3330 (N_3330,N_3202,N_3272);
or U3331 (N_3331,N_3225,N_3262);
nand U3332 (N_3332,N_3220,N_3230);
xor U3333 (N_3333,N_3206,N_3266);
nand U3334 (N_3334,N_3201,N_3260);
or U3335 (N_3335,N_3265,N_3214);
or U3336 (N_3336,N_3224,N_3249);
nor U3337 (N_3337,N_3245,N_3241);
nor U3338 (N_3338,N_3243,N_3289);
or U3339 (N_3339,N_3208,N_3213);
nand U3340 (N_3340,N_3275,N_3235);
nand U3341 (N_3341,N_3287,N_3240);
and U3342 (N_3342,N_3229,N_3203);
nor U3343 (N_3343,N_3267,N_3270);
nor U3344 (N_3344,N_3227,N_3290);
xnor U3345 (N_3345,N_3252,N_3239);
or U3346 (N_3346,N_3251,N_3291);
nor U3347 (N_3347,N_3282,N_3264);
or U3348 (N_3348,N_3253,N_3292);
or U3349 (N_3349,N_3299,N_3258);
xor U3350 (N_3350,N_3257,N_3207);
and U3351 (N_3351,N_3216,N_3255);
nand U3352 (N_3352,N_3286,N_3224);
or U3353 (N_3353,N_3260,N_3265);
nor U3354 (N_3354,N_3213,N_3258);
and U3355 (N_3355,N_3240,N_3233);
nor U3356 (N_3356,N_3276,N_3212);
and U3357 (N_3357,N_3235,N_3216);
xnor U3358 (N_3358,N_3268,N_3233);
and U3359 (N_3359,N_3237,N_3217);
nand U3360 (N_3360,N_3244,N_3258);
xnor U3361 (N_3361,N_3224,N_3235);
and U3362 (N_3362,N_3289,N_3221);
or U3363 (N_3363,N_3299,N_3249);
nand U3364 (N_3364,N_3270,N_3287);
xor U3365 (N_3365,N_3273,N_3201);
or U3366 (N_3366,N_3225,N_3212);
or U3367 (N_3367,N_3257,N_3280);
xor U3368 (N_3368,N_3262,N_3246);
nand U3369 (N_3369,N_3268,N_3228);
and U3370 (N_3370,N_3288,N_3215);
and U3371 (N_3371,N_3201,N_3242);
nor U3372 (N_3372,N_3247,N_3207);
nor U3373 (N_3373,N_3261,N_3266);
or U3374 (N_3374,N_3261,N_3272);
xor U3375 (N_3375,N_3285,N_3283);
or U3376 (N_3376,N_3295,N_3279);
or U3377 (N_3377,N_3211,N_3207);
or U3378 (N_3378,N_3221,N_3230);
nand U3379 (N_3379,N_3201,N_3281);
or U3380 (N_3380,N_3265,N_3211);
and U3381 (N_3381,N_3295,N_3209);
and U3382 (N_3382,N_3200,N_3220);
nand U3383 (N_3383,N_3249,N_3295);
nor U3384 (N_3384,N_3224,N_3226);
xor U3385 (N_3385,N_3276,N_3254);
and U3386 (N_3386,N_3228,N_3294);
nor U3387 (N_3387,N_3247,N_3298);
nor U3388 (N_3388,N_3273,N_3211);
nor U3389 (N_3389,N_3295,N_3290);
nand U3390 (N_3390,N_3229,N_3295);
nor U3391 (N_3391,N_3263,N_3214);
xnor U3392 (N_3392,N_3221,N_3203);
and U3393 (N_3393,N_3286,N_3267);
nand U3394 (N_3394,N_3258,N_3268);
nand U3395 (N_3395,N_3222,N_3260);
nor U3396 (N_3396,N_3210,N_3286);
or U3397 (N_3397,N_3261,N_3201);
nand U3398 (N_3398,N_3204,N_3276);
nand U3399 (N_3399,N_3276,N_3222);
nor U3400 (N_3400,N_3321,N_3311);
and U3401 (N_3401,N_3307,N_3343);
or U3402 (N_3402,N_3356,N_3323);
xor U3403 (N_3403,N_3391,N_3353);
and U3404 (N_3404,N_3339,N_3303);
or U3405 (N_3405,N_3351,N_3317);
and U3406 (N_3406,N_3397,N_3377);
or U3407 (N_3407,N_3330,N_3362);
nand U3408 (N_3408,N_3385,N_3398);
nor U3409 (N_3409,N_3386,N_3383);
and U3410 (N_3410,N_3369,N_3325);
nand U3411 (N_3411,N_3324,N_3352);
nand U3412 (N_3412,N_3335,N_3322);
nor U3413 (N_3413,N_3380,N_3389);
and U3414 (N_3414,N_3372,N_3300);
or U3415 (N_3415,N_3337,N_3308);
and U3416 (N_3416,N_3341,N_3350);
or U3417 (N_3417,N_3387,N_3364);
or U3418 (N_3418,N_3390,N_3310);
nor U3419 (N_3419,N_3381,N_3320);
nand U3420 (N_3420,N_3370,N_3306);
nor U3421 (N_3421,N_3319,N_3312);
xor U3422 (N_3422,N_3327,N_3318);
and U3423 (N_3423,N_3309,N_3365);
and U3424 (N_3424,N_3378,N_3355);
nand U3425 (N_3425,N_3315,N_3344);
nor U3426 (N_3426,N_3368,N_3328);
nand U3427 (N_3427,N_3302,N_3360);
or U3428 (N_3428,N_3396,N_3345);
and U3429 (N_3429,N_3338,N_3301);
and U3430 (N_3430,N_3392,N_3395);
nor U3431 (N_3431,N_3333,N_3342);
nand U3432 (N_3432,N_3366,N_3316);
and U3433 (N_3433,N_3314,N_3313);
nor U3434 (N_3434,N_3384,N_3393);
and U3435 (N_3435,N_3359,N_3399);
xnor U3436 (N_3436,N_3379,N_3357);
nand U3437 (N_3437,N_3371,N_3349);
or U3438 (N_3438,N_3340,N_3367);
nand U3439 (N_3439,N_3326,N_3334);
xor U3440 (N_3440,N_3332,N_3376);
nor U3441 (N_3441,N_3346,N_3347);
nand U3442 (N_3442,N_3305,N_3358);
nor U3443 (N_3443,N_3382,N_3354);
and U3444 (N_3444,N_3375,N_3394);
xor U3445 (N_3445,N_3361,N_3331);
or U3446 (N_3446,N_3348,N_3363);
nand U3447 (N_3447,N_3329,N_3388);
nor U3448 (N_3448,N_3373,N_3304);
or U3449 (N_3449,N_3374,N_3336);
nand U3450 (N_3450,N_3365,N_3353);
or U3451 (N_3451,N_3399,N_3363);
or U3452 (N_3452,N_3300,N_3318);
and U3453 (N_3453,N_3386,N_3371);
nor U3454 (N_3454,N_3345,N_3301);
or U3455 (N_3455,N_3336,N_3370);
nor U3456 (N_3456,N_3336,N_3371);
and U3457 (N_3457,N_3399,N_3368);
nand U3458 (N_3458,N_3328,N_3393);
nor U3459 (N_3459,N_3385,N_3316);
nand U3460 (N_3460,N_3382,N_3312);
and U3461 (N_3461,N_3362,N_3354);
or U3462 (N_3462,N_3350,N_3398);
xnor U3463 (N_3463,N_3390,N_3356);
or U3464 (N_3464,N_3311,N_3345);
xor U3465 (N_3465,N_3349,N_3303);
xor U3466 (N_3466,N_3304,N_3316);
xnor U3467 (N_3467,N_3305,N_3355);
nor U3468 (N_3468,N_3342,N_3340);
and U3469 (N_3469,N_3308,N_3371);
nand U3470 (N_3470,N_3309,N_3366);
nand U3471 (N_3471,N_3391,N_3342);
nor U3472 (N_3472,N_3398,N_3315);
nor U3473 (N_3473,N_3316,N_3319);
and U3474 (N_3474,N_3355,N_3333);
nand U3475 (N_3475,N_3365,N_3386);
and U3476 (N_3476,N_3344,N_3312);
nand U3477 (N_3477,N_3393,N_3351);
or U3478 (N_3478,N_3392,N_3364);
nor U3479 (N_3479,N_3382,N_3344);
nor U3480 (N_3480,N_3385,N_3363);
or U3481 (N_3481,N_3349,N_3358);
xnor U3482 (N_3482,N_3358,N_3362);
and U3483 (N_3483,N_3363,N_3355);
and U3484 (N_3484,N_3336,N_3332);
nand U3485 (N_3485,N_3381,N_3393);
or U3486 (N_3486,N_3394,N_3343);
or U3487 (N_3487,N_3333,N_3381);
xnor U3488 (N_3488,N_3339,N_3383);
nand U3489 (N_3489,N_3320,N_3350);
nor U3490 (N_3490,N_3317,N_3337);
nand U3491 (N_3491,N_3336,N_3373);
and U3492 (N_3492,N_3372,N_3358);
xnor U3493 (N_3493,N_3344,N_3306);
xor U3494 (N_3494,N_3323,N_3340);
xor U3495 (N_3495,N_3376,N_3319);
or U3496 (N_3496,N_3338,N_3334);
or U3497 (N_3497,N_3300,N_3373);
or U3498 (N_3498,N_3328,N_3361);
nor U3499 (N_3499,N_3398,N_3303);
nor U3500 (N_3500,N_3489,N_3470);
and U3501 (N_3501,N_3406,N_3416);
nand U3502 (N_3502,N_3497,N_3437);
nand U3503 (N_3503,N_3403,N_3432);
nand U3504 (N_3504,N_3421,N_3477);
nand U3505 (N_3505,N_3492,N_3499);
or U3506 (N_3506,N_3481,N_3436);
nor U3507 (N_3507,N_3417,N_3400);
xnor U3508 (N_3508,N_3482,N_3467);
or U3509 (N_3509,N_3486,N_3404);
and U3510 (N_3510,N_3483,N_3488);
nand U3511 (N_3511,N_3485,N_3453);
nand U3512 (N_3512,N_3475,N_3454);
or U3513 (N_3513,N_3465,N_3402);
and U3514 (N_3514,N_3476,N_3455);
xnor U3515 (N_3515,N_3443,N_3431);
nor U3516 (N_3516,N_3424,N_3474);
nand U3517 (N_3517,N_3444,N_3407);
xnor U3518 (N_3518,N_3445,N_3411);
xnor U3519 (N_3519,N_3464,N_3426);
or U3520 (N_3520,N_3423,N_3409);
xor U3521 (N_3521,N_3447,N_3408);
nor U3522 (N_3522,N_3468,N_3433);
nor U3523 (N_3523,N_3466,N_3401);
or U3524 (N_3524,N_3422,N_3452);
nand U3525 (N_3525,N_3461,N_3484);
xnor U3526 (N_3526,N_3439,N_3435);
nand U3527 (N_3527,N_3420,N_3456);
or U3528 (N_3528,N_3472,N_3412);
nand U3529 (N_3529,N_3418,N_3496);
nor U3530 (N_3530,N_3480,N_3425);
nand U3531 (N_3531,N_3441,N_3490);
and U3532 (N_3532,N_3491,N_3434);
and U3533 (N_3533,N_3448,N_3430);
and U3534 (N_3534,N_3462,N_3413);
nand U3535 (N_3535,N_3438,N_3429);
and U3536 (N_3536,N_3469,N_3419);
or U3537 (N_3537,N_3498,N_3427);
nor U3538 (N_3538,N_3446,N_3410);
nand U3539 (N_3539,N_3460,N_3463);
xor U3540 (N_3540,N_3495,N_3478);
xor U3541 (N_3541,N_3415,N_3471);
nand U3542 (N_3542,N_3442,N_3458);
nand U3543 (N_3543,N_3493,N_3405);
or U3544 (N_3544,N_3479,N_3457);
and U3545 (N_3545,N_3440,N_3494);
nor U3546 (N_3546,N_3449,N_3450);
or U3547 (N_3547,N_3428,N_3414);
nand U3548 (N_3548,N_3451,N_3459);
xnor U3549 (N_3549,N_3473,N_3487);
nor U3550 (N_3550,N_3498,N_3434);
xnor U3551 (N_3551,N_3401,N_3427);
xor U3552 (N_3552,N_3435,N_3466);
xnor U3553 (N_3553,N_3435,N_3497);
and U3554 (N_3554,N_3469,N_3467);
xor U3555 (N_3555,N_3425,N_3412);
or U3556 (N_3556,N_3407,N_3469);
xor U3557 (N_3557,N_3455,N_3447);
xor U3558 (N_3558,N_3497,N_3482);
nor U3559 (N_3559,N_3469,N_3457);
and U3560 (N_3560,N_3443,N_3491);
nor U3561 (N_3561,N_3431,N_3450);
and U3562 (N_3562,N_3498,N_3499);
nand U3563 (N_3563,N_3447,N_3430);
nor U3564 (N_3564,N_3458,N_3404);
and U3565 (N_3565,N_3457,N_3432);
or U3566 (N_3566,N_3451,N_3429);
nand U3567 (N_3567,N_3480,N_3490);
and U3568 (N_3568,N_3411,N_3467);
nor U3569 (N_3569,N_3409,N_3446);
and U3570 (N_3570,N_3413,N_3460);
or U3571 (N_3571,N_3401,N_3485);
and U3572 (N_3572,N_3421,N_3424);
nor U3573 (N_3573,N_3427,N_3479);
nand U3574 (N_3574,N_3480,N_3478);
and U3575 (N_3575,N_3465,N_3489);
nand U3576 (N_3576,N_3424,N_3468);
or U3577 (N_3577,N_3421,N_3429);
nand U3578 (N_3578,N_3451,N_3443);
nand U3579 (N_3579,N_3413,N_3482);
xnor U3580 (N_3580,N_3468,N_3403);
or U3581 (N_3581,N_3480,N_3402);
or U3582 (N_3582,N_3420,N_3475);
and U3583 (N_3583,N_3446,N_3418);
and U3584 (N_3584,N_3419,N_3425);
nand U3585 (N_3585,N_3467,N_3436);
xnor U3586 (N_3586,N_3497,N_3477);
nand U3587 (N_3587,N_3459,N_3449);
or U3588 (N_3588,N_3451,N_3445);
xor U3589 (N_3589,N_3462,N_3441);
or U3590 (N_3590,N_3411,N_3468);
xor U3591 (N_3591,N_3470,N_3420);
nand U3592 (N_3592,N_3496,N_3443);
nor U3593 (N_3593,N_3464,N_3400);
nand U3594 (N_3594,N_3472,N_3409);
and U3595 (N_3595,N_3411,N_3403);
xor U3596 (N_3596,N_3408,N_3485);
and U3597 (N_3597,N_3415,N_3403);
nand U3598 (N_3598,N_3406,N_3475);
and U3599 (N_3599,N_3486,N_3421);
or U3600 (N_3600,N_3503,N_3542);
xor U3601 (N_3601,N_3505,N_3533);
nor U3602 (N_3602,N_3572,N_3546);
and U3603 (N_3603,N_3501,N_3527);
xor U3604 (N_3604,N_3580,N_3579);
nor U3605 (N_3605,N_3512,N_3528);
xnor U3606 (N_3606,N_3565,N_3581);
nor U3607 (N_3607,N_3507,N_3545);
or U3608 (N_3608,N_3595,N_3568);
nand U3609 (N_3609,N_3564,N_3582);
nor U3610 (N_3610,N_3514,N_3555);
xnor U3611 (N_3611,N_3571,N_3547);
nor U3612 (N_3612,N_3518,N_3543);
and U3613 (N_3613,N_3583,N_3500);
and U3614 (N_3614,N_3526,N_3540);
or U3615 (N_3615,N_3589,N_3531);
nor U3616 (N_3616,N_3515,N_3576);
nor U3617 (N_3617,N_3521,N_3520);
nor U3618 (N_3618,N_3563,N_3567);
xnor U3619 (N_3619,N_3506,N_3508);
nor U3620 (N_3620,N_3502,N_3590);
nor U3621 (N_3621,N_3516,N_3551);
nand U3622 (N_3622,N_3525,N_3561);
or U3623 (N_3623,N_3592,N_3596);
xnor U3624 (N_3624,N_3534,N_3522);
xor U3625 (N_3625,N_3559,N_3544);
or U3626 (N_3626,N_3593,N_3578);
and U3627 (N_3627,N_3585,N_3536);
xnor U3628 (N_3628,N_3530,N_3511);
nor U3629 (N_3629,N_3558,N_3510);
nand U3630 (N_3630,N_3566,N_3541);
nand U3631 (N_3631,N_3560,N_3594);
or U3632 (N_3632,N_3519,N_3537);
nand U3633 (N_3633,N_3587,N_3548);
nand U3634 (N_3634,N_3554,N_3517);
and U3635 (N_3635,N_3538,N_3539);
nand U3636 (N_3636,N_3529,N_3588);
nand U3637 (N_3637,N_3552,N_3586);
nand U3638 (N_3638,N_3557,N_3597);
nand U3639 (N_3639,N_3524,N_3556);
nor U3640 (N_3640,N_3535,N_3599);
nand U3641 (N_3641,N_3562,N_3504);
or U3642 (N_3642,N_3513,N_3553);
xor U3643 (N_3643,N_3549,N_3577);
xor U3644 (N_3644,N_3574,N_3575);
nor U3645 (N_3645,N_3591,N_3550);
or U3646 (N_3646,N_3598,N_3509);
or U3647 (N_3647,N_3569,N_3573);
and U3648 (N_3648,N_3570,N_3584);
nor U3649 (N_3649,N_3523,N_3532);
xor U3650 (N_3650,N_3525,N_3539);
xnor U3651 (N_3651,N_3550,N_3554);
and U3652 (N_3652,N_3586,N_3563);
nor U3653 (N_3653,N_3570,N_3503);
nor U3654 (N_3654,N_3511,N_3594);
xnor U3655 (N_3655,N_3578,N_3557);
or U3656 (N_3656,N_3580,N_3545);
nor U3657 (N_3657,N_3509,N_3522);
or U3658 (N_3658,N_3529,N_3533);
nand U3659 (N_3659,N_3537,N_3544);
nand U3660 (N_3660,N_3500,N_3596);
or U3661 (N_3661,N_3520,N_3572);
and U3662 (N_3662,N_3560,N_3508);
or U3663 (N_3663,N_3540,N_3549);
or U3664 (N_3664,N_3567,N_3536);
xor U3665 (N_3665,N_3579,N_3528);
nand U3666 (N_3666,N_3529,N_3587);
and U3667 (N_3667,N_3551,N_3570);
or U3668 (N_3668,N_3555,N_3585);
or U3669 (N_3669,N_3590,N_3577);
or U3670 (N_3670,N_3513,N_3541);
and U3671 (N_3671,N_3501,N_3578);
nor U3672 (N_3672,N_3598,N_3552);
nand U3673 (N_3673,N_3555,N_3515);
xnor U3674 (N_3674,N_3500,N_3580);
and U3675 (N_3675,N_3573,N_3599);
nor U3676 (N_3676,N_3525,N_3517);
or U3677 (N_3677,N_3518,N_3550);
and U3678 (N_3678,N_3563,N_3548);
or U3679 (N_3679,N_3507,N_3566);
xnor U3680 (N_3680,N_3559,N_3502);
nand U3681 (N_3681,N_3504,N_3520);
nor U3682 (N_3682,N_3590,N_3597);
and U3683 (N_3683,N_3538,N_3506);
nand U3684 (N_3684,N_3590,N_3596);
or U3685 (N_3685,N_3567,N_3588);
nand U3686 (N_3686,N_3589,N_3528);
nand U3687 (N_3687,N_3508,N_3590);
or U3688 (N_3688,N_3530,N_3577);
nand U3689 (N_3689,N_3542,N_3508);
and U3690 (N_3690,N_3566,N_3592);
nand U3691 (N_3691,N_3562,N_3518);
nand U3692 (N_3692,N_3520,N_3574);
nor U3693 (N_3693,N_3539,N_3528);
xnor U3694 (N_3694,N_3556,N_3539);
or U3695 (N_3695,N_3581,N_3589);
or U3696 (N_3696,N_3595,N_3532);
and U3697 (N_3697,N_3540,N_3521);
xnor U3698 (N_3698,N_3512,N_3583);
and U3699 (N_3699,N_3515,N_3556);
nor U3700 (N_3700,N_3617,N_3600);
and U3701 (N_3701,N_3653,N_3632);
or U3702 (N_3702,N_3657,N_3626);
nand U3703 (N_3703,N_3665,N_3672);
nand U3704 (N_3704,N_3631,N_3640);
and U3705 (N_3705,N_3614,N_3642);
nor U3706 (N_3706,N_3644,N_3694);
nor U3707 (N_3707,N_3636,N_3683);
and U3708 (N_3708,N_3684,N_3629);
or U3709 (N_3709,N_3655,N_3690);
xor U3710 (N_3710,N_3661,N_3609);
or U3711 (N_3711,N_3627,N_3681);
and U3712 (N_3712,N_3678,N_3602);
and U3713 (N_3713,N_3620,N_3658);
nand U3714 (N_3714,N_3676,N_3688);
xor U3715 (N_3715,N_3605,N_3686);
or U3716 (N_3716,N_3603,N_3639);
nand U3717 (N_3717,N_3666,N_3618);
and U3718 (N_3718,N_3662,N_3638);
nand U3719 (N_3719,N_3669,N_3622);
nand U3720 (N_3720,N_3668,N_3673);
nand U3721 (N_3721,N_3635,N_3660);
xor U3722 (N_3722,N_3651,N_3659);
nand U3723 (N_3723,N_3611,N_3606);
xnor U3724 (N_3724,N_3652,N_3610);
nand U3725 (N_3725,N_3647,N_3675);
and U3726 (N_3726,N_3654,N_3619);
or U3727 (N_3727,N_3692,N_3615);
and U3728 (N_3728,N_3634,N_3641);
nand U3729 (N_3729,N_3685,N_3637);
nor U3730 (N_3730,N_3696,N_3648);
and U3731 (N_3731,N_3643,N_3671);
and U3732 (N_3732,N_3616,N_3656);
nand U3733 (N_3733,N_3645,N_3679);
xor U3734 (N_3734,N_3667,N_3698);
nor U3735 (N_3735,N_3682,N_3630);
nand U3736 (N_3736,N_3691,N_3612);
and U3737 (N_3737,N_3699,N_3650);
nand U3738 (N_3738,N_3625,N_3664);
xor U3739 (N_3739,N_3677,N_3693);
xnor U3740 (N_3740,N_3646,N_3624);
or U3741 (N_3741,N_3689,N_3680);
or U3742 (N_3742,N_3628,N_3695);
and U3743 (N_3743,N_3674,N_3613);
nand U3744 (N_3744,N_3621,N_3687);
nand U3745 (N_3745,N_3663,N_3670);
and U3746 (N_3746,N_3604,N_3649);
and U3747 (N_3747,N_3601,N_3623);
xnor U3748 (N_3748,N_3607,N_3697);
xor U3749 (N_3749,N_3608,N_3633);
xor U3750 (N_3750,N_3689,N_3684);
nor U3751 (N_3751,N_3615,N_3602);
nand U3752 (N_3752,N_3646,N_3670);
nand U3753 (N_3753,N_3620,N_3678);
and U3754 (N_3754,N_3619,N_3633);
nand U3755 (N_3755,N_3634,N_3669);
or U3756 (N_3756,N_3644,N_3646);
or U3757 (N_3757,N_3650,N_3680);
or U3758 (N_3758,N_3606,N_3687);
and U3759 (N_3759,N_3688,N_3675);
nand U3760 (N_3760,N_3609,N_3622);
or U3761 (N_3761,N_3652,N_3616);
xor U3762 (N_3762,N_3623,N_3621);
nand U3763 (N_3763,N_3613,N_3600);
and U3764 (N_3764,N_3606,N_3683);
or U3765 (N_3765,N_3631,N_3645);
xnor U3766 (N_3766,N_3618,N_3660);
nor U3767 (N_3767,N_3626,N_3691);
xor U3768 (N_3768,N_3609,N_3637);
xnor U3769 (N_3769,N_3690,N_3637);
xor U3770 (N_3770,N_3643,N_3645);
and U3771 (N_3771,N_3600,N_3697);
or U3772 (N_3772,N_3696,N_3659);
nand U3773 (N_3773,N_3605,N_3626);
or U3774 (N_3774,N_3650,N_3687);
nand U3775 (N_3775,N_3602,N_3626);
nor U3776 (N_3776,N_3601,N_3685);
nand U3777 (N_3777,N_3684,N_3620);
or U3778 (N_3778,N_3687,N_3636);
or U3779 (N_3779,N_3656,N_3675);
and U3780 (N_3780,N_3657,N_3670);
and U3781 (N_3781,N_3656,N_3613);
or U3782 (N_3782,N_3636,N_3663);
xnor U3783 (N_3783,N_3688,N_3628);
and U3784 (N_3784,N_3654,N_3635);
or U3785 (N_3785,N_3655,N_3685);
and U3786 (N_3786,N_3670,N_3625);
xor U3787 (N_3787,N_3650,N_3636);
nor U3788 (N_3788,N_3622,N_3678);
nor U3789 (N_3789,N_3698,N_3605);
nor U3790 (N_3790,N_3624,N_3633);
or U3791 (N_3791,N_3610,N_3615);
nand U3792 (N_3792,N_3665,N_3615);
or U3793 (N_3793,N_3675,N_3614);
nand U3794 (N_3794,N_3674,N_3626);
or U3795 (N_3795,N_3686,N_3687);
nand U3796 (N_3796,N_3679,N_3671);
or U3797 (N_3797,N_3649,N_3660);
nor U3798 (N_3798,N_3620,N_3672);
nor U3799 (N_3799,N_3699,N_3635);
nand U3800 (N_3800,N_3706,N_3760);
or U3801 (N_3801,N_3785,N_3787);
xnor U3802 (N_3802,N_3708,N_3759);
and U3803 (N_3803,N_3773,N_3744);
nor U3804 (N_3804,N_3761,N_3743);
nand U3805 (N_3805,N_3788,N_3745);
xnor U3806 (N_3806,N_3752,N_3724);
or U3807 (N_3807,N_3741,N_3723);
xor U3808 (N_3808,N_3707,N_3795);
or U3809 (N_3809,N_3799,N_3784);
and U3810 (N_3810,N_3746,N_3711);
nor U3811 (N_3811,N_3767,N_3715);
xor U3812 (N_3812,N_3792,N_3753);
nand U3813 (N_3813,N_3726,N_3778);
and U3814 (N_3814,N_3733,N_3734);
and U3815 (N_3815,N_3716,N_3789);
nor U3816 (N_3816,N_3727,N_3779);
xnor U3817 (N_3817,N_3751,N_3776);
and U3818 (N_3818,N_3754,N_3771);
and U3819 (N_3819,N_3703,N_3702);
nor U3820 (N_3820,N_3762,N_3765);
or U3821 (N_3821,N_3731,N_3705);
xnor U3822 (N_3822,N_3719,N_3797);
xnor U3823 (N_3823,N_3732,N_3735);
or U3824 (N_3824,N_3783,N_3710);
nor U3825 (N_3825,N_3747,N_3701);
nor U3826 (N_3826,N_3748,N_3737);
xor U3827 (N_3827,N_3739,N_3780);
xnor U3828 (N_3828,N_3791,N_3736);
and U3829 (N_3829,N_3722,N_3730);
nand U3830 (N_3830,N_3777,N_3728);
nand U3831 (N_3831,N_3755,N_3709);
and U3832 (N_3832,N_3794,N_3781);
and U3833 (N_3833,N_3796,N_3772);
and U3834 (N_3834,N_3793,N_3718);
and U3835 (N_3835,N_3782,N_3774);
and U3836 (N_3836,N_3770,N_3757);
nor U3837 (N_3837,N_3704,N_3700);
xor U3838 (N_3838,N_3764,N_3714);
nand U3839 (N_3839,N_3798,N_3756);
xnor U3840 (N_3840,N_3763,N_3720);
xnor U3841 (N_3841,N_3740,N_3775);
and U3842 (N_3842,N_3749,N_3717);
nor U3843 (N_3843,N_3729,N_3712);
nor U3844 (N_3844,N_3721,N_3766);
nand U3845 (N_3845,N_3786,N_3738);
or U3846 (N_3846,N_3758,N_3768);
or U3847 (N_3847,N_3790,N_3742);
nand U3848 (N_3848,N_3713,N_3769);
or U3849 (N_3849,N_3750,N_3725);
nor U3850 (N_3850,N_3764,N_3728);
nand U3851 (N_3851,N_3720,N_3732);
and U3852 (N_3852,N_3774,N_3780);
or U3853 (N_3853,N_3778,N_3793);
nor U3854 (N_3854,N_3745,N_3770);
nand U3855 (N_3855,N_3786,N_3744);
and U3856 (N_3856,N_3751,N_3713);
xnor U3857 (N_3857,N_3755,N_3729);
and U3858 (N_3858,N_3799,N_3709);
nor U3859 (N_3859,N_3759,N_3739);
and U3860 (N_3860,N_3729,N_3783);
xor U3861 (N_3861,N_3753,N_3703);
nor U3862 (N_3862,N_3772,N_3706);
nand U3863 (N_3863,N_3735,N_3795);
and U3864 (N_3864,N_3773,N_3791);
nand U3865 (N_3865,N_3778,N_3786);
or U3866 (N_3866,N_3754,N_3762);
nor U3867 (N_3867,N_3736,N_3757);
nand U3868 (N_3868,N_3753,N_3763);
nand U3869 (N_3869,N_3740,N_3745);
xor U3870 (N_3870,N_3715,N_3745);
and U3871 (N_3871,N_3757,N_3795);
xor U3872 (N_3872,N_3727,N_3740);
nand U3873 (N_3873,N_3739,N_3773);
or U3874 (N_3874,N_3753,N_3729);
nand U3875 (N_3875,N_3721,N_3759);
nand U3876 (N_3876,N_3706,N_3757);
or U3877 (N_3877,N_3711,N_3725);
nor U3878 (N_3878,N_3757,N_3785);
or U3879 (N_3879,N_3706,N_3779);
nand U3880 (N_3880,N_3784,N_3744);
nor U3881 (N_3881,N_3748,N_3786);
or U3882 (N_3882,N_3771,N_3744);
nor U3883 (N_3883,N_3703,N_3717);
nand U3884 (N_3884,N_3761,N_3702);
and U3885 (N_3885,N_3731,N_3778);
xor U3886 (N_3886,N_3721,N_3714);
nand U3887 (N_3887,N_3730,N_3716);
or U3888 (N_3888,N_3702,N_3738);
nor U3889 (N_3889,N_3763,N_3769);
xnor U3890 (N_3890,N_3795,N_3765);
xor U3891 (N_3891,N_3712,N_3750);
and U3892 (N_3892,N_3735,N_3744);
nor U3893 (N_3893,N_3709,N_3741);
nor U3894 (N_3894,N_3748,N_3799);
nand U3895 (N_3895,N_3719,N_3703);
and U3896 (N_3896,N_3767,N_3732);
xor U3897 (N_3897,N_3796,N_3742);
nand U3898 (N_3898,N_3752,N_3764);
nand U3899 (N_3899,N_3746,N_3720);
xor U3900 (N_3900,N_3819,N_3864);
nor U3901 (N_3901,N_3886,N_3821);
nand U3902 (N_3902,N_3883,N_3820);
and U3903 (N_3903,N_3870,N_3854);
xor U3904 (N_3904,N_3803,N_3810);
and U3905 (N_3905,N_3892,N_3859);
nand U3906 (N_3906,N_3836,N_3815);
nand U3907 (N_3907,N_3863,N_3869);
nand U3908 (N_3908,N_3804,N_3835);
or U3909 (N_3909,N_3889,N_3805);
or U3910 (N_3910,N_3827,N_3816);
xor U3911 (N_3911,N_3817,N_3801);
or U3912 (N_3912,N_3822,N_3885);
and U3913 (N_3913,N_3865,N_3808);
nor U3914 (N_3914,N_3813,N_3880);
nand U3915 (N_3915,N_3826,N_3847);
or U3916 (N_3916,N_3830,N_3856);
nor U3917 (N_3917,N_3882,N_3894);
or U3918 (N_3918,N_3838,N_3843);
or U3919 (N_3919,N_3895,N_3832);
nand U3920 (N_3920,N_3867,N_3834);
nand U3921 (N_3921,N_3839,N_3876);
xor U3922 (N_3922,N_3855,N_3861);
nand U3923 (N_3923,N_3858,N_3850);
and U3924 (N_3924,N_3831,N_3860);
xor U3925 (N_3925,N_3833,N_3828);
and U3926 (N_3926,N_3898,N_3806);
or U3927 (N_3927,N_3812,N_3891);
nor U3928 (N_3928,N_3872,N_3851);
nand U3929 (N_3929,N_3809,N_3897);
nor U3930 (N_3930,N_3884,N_3823);
xnor U3931 (N_3931,N_3893,N_3840);
or U3932 (N_3932,N_3879,N_3814);
nand U3933 (N_3933,N_3888,N_3874);
nor U3934 (N_3934,N_3852,N_3849);
nor U3935 (N_3935,N_3866,N_3887);
or U3936 (N_3936,N_3873,N_3846);
nor U3937 (N_3937,N_3845,N_3824);
and U3938 (N_3938,N_3811,N_3841);
or U3939 (N_3939,N_3890,N_3853);
nand U3940 (N_3940,N_3871,N_3899);
xor U3941 (N_3941,N_3829,N_3857);
nand U3942 (N_3942,N_3875,N_3868);
nor U3943 (N_3943,N_3825,N_3862);
and U3944 (N_3944,N_3800,N_3877);
or U3945 (N_3945,N_3848,N_3842);
xnor U3946 (N_3946,N_3896,N_3807);
and U3947 (N_3947,N_3881,N_3818);
and U3948 (N_3948,N_3802,N_3844);
nand U3949 (N_3949,N_3837,N_3878);
xor U3950 (N_3950,N_3808,N_3872);
xor U3951 (N_3951,N_3897,N_3880);
nand U3952 (N_3952,N_3855,N_3892);
xor U3953 (N_3953,N_3805,N_3884);
and U3954 (N_3954,N_3836,N_3807);
nand U3955 (N_3955,N_3848,N_3859);
or U3956 (N_3956,N_3872,N_3844);
xnor U3957 (N_3957,N_3821,N_3893);
xor U3958 (N_3958,N_3878,N_3832);
nor U3959 (N_3959,N_3852,N_3831);
or U3960 (N_3960,N_3812,N_3885);
nor U3961 (N_3961,N_3801,N_3896);
xor U3962 (N_3962,N_3863,N_3895);
and U3963 (N_3963,N_3894,N_3838);
xor U3964 (N_3964,N_3857,N_3818);
xnor U3965 (N_3965,N_3856,N_3848);
nand U3966 (N_3966,N_3826,N_3803);
or U3967 (N_3967,N_3861,N_3841);
and U3968 (N_3968,N_3888,N_3890);
xnor U3969 (N_3969,N_3875,N_3897);
and U3970 (N_3970,N_3812,N_3841);
or U3971 (N_3971,N_3871,N_3885);
or U3972 (N_3972,N_3877,N_3884);
or U3973 (N_3973,N_3827,N_3847);
or U3974 (N_3974,N_3866,N_3880);
nand U3975 (N_3975,N_3840,N_3835);
nor U3976 (N_3976,N_3826,N_3822);
nor U3977 (N_3977,N_3875,N_3888);
nand U3978 (N_3978,N_3857,N_3817);
or U3979 (N_3979,N_3864,N_3842);
nand U3980 (N_3980,N_3884,N_3857);
and U3981 (N_3981,N_3849,N_3820);
xnor U3982 (N_3982,N_3845,N_3813);
or U3983 (N_3983,N_3854,N_3801);
and U3984 (N_3984,N_3857,N_3840);
xor U3985 (N_3985,N_3878,N_3825);
xor U3986 (N_3986,N_3827,N_3868);
nand U3987 (N_3987,N_3870,N_3837);
and U3988 (N_3988,N_3894,N_3811);
or U3989 (N_3989,N_3866,N_3804);
xor U3990 (N_3990,N_3861,N_3888);
or U3991 (N_3991,N_3833,N_3865);
xnor U3992 (N_3992,N_3861,N_3807);
or U3993 (N_3993,N_3829,N_3849);
xor U3994 (N_3994,N_3869,N_3833);
nand U3995 (N_3995,N_3853,N_3840);
and U3996 (N_3996,N_3844,N_3875);
nand U3997 (N_3997,N_3882,N_3868);
nor U3998 (N_3998,N_3838,N_3866);
nand U3999 (N_3999,N_3887,N_3833);
or U4000 (N_4000,N_3990,N_3969);
or U4001 (N_4001,N_3904,N_3961);
and U4002 (N_4002,N_3992,N_3993);
and U4003 (N_4003,N_3922,N_3979);
nor U4004 (N_4004,N_3938,N_3900);
or U4005 (N_4005,N_3920,N_3980);
and U4006 (N_4006,N_3937,N_3978);
nor U4007 (N_4007,N_3928,N_3952);
nand U4008 (N_4008,N_3913,N_3956);
or U4009 (N_4009,N_3929,N_3935);
and U4010 (N_4010,N_3974,N_3940);
and U4011 (N_4011,N_3989,N_3964);
xnor U4012 (N_4012,N_3965,N_3986);
nor U4013 (N_4013,N_3977,N_3941);
and U4014 (N_4014,N_3946,N_3912);
nand U4015 (N_4015,N_3909,N_3983);
or U4016 (N_4016,N_3963,N_3925);
nor U4017 (N_4017,N_3995,N_3936);
xnor U4018 (N_4018,N_3973,N_3906);
xnor U4019 (N_4019,N_3947,N_3923);
nand U4020 (N_4020,N_3960,N_3931);
nand U4021 (N_4021,N_3958,N_3939);
nand U4022 (N_4022,N_3998,N_3996);
nand U4023 (N_4023,N_3988,N_3950);
and U4024 (N_4024,N_3901,N_3970);
and U4025 (N_4025,N_3934,N_3966);
and U4026 (N_4026,N_3902,N_3933);
nand U4027 (N_4027,N_3943,N_3953);
and U4028 (N_4028,N_3907,N_3945);
or U4029 (N_4029,N_3984,N_3914);
and U4030 (N_4030,N_3955,N_3930);
or U4031 (N_4031,N_3962,N_3949);
nor U4032 (N_4032,N_3903,N_3919);
nor U4033 (N_4033,N_3976,N_3917);
nor U4034 (N_4034,N_3916,N_3926);
nand U4035 (N_4035,N_3971,N_3982);
and U4036 (N_4036,N_3987,N_3944);
and U4037 (N_4037,N_3959,N_3927);
nand U4038 (N_4038,N_3951,N_3968);
and U4039 (N_4039,N_3911,N_3997);
nand U4040 (N_4040,N_3985,N_3918);
or U4041 (N_4041,N_3957,N_3991);
or U4042 (N_4042,N_3954,N_3932);
and U4043 (N_4043,N_3972,N_3994);
and U4044 (N_4044,N_3910,N_3905);
nor U4045 (N_4045,N_3948,N_3908);
nor U4046 (N_4046,N_3942,N_3967);
nand U4047 (N_4047,N_3975,N_3924);
xor U4048 (N_4048,N_3915,N_3981);
and U4049 (N_4049,N_3999,N_3921);
or U4050 (N_4050,N_3934,N_3967);
nand U4051 (N_4051,N_3925,N_3998);
nand U4052 (N_4052,N_3953,N_3962);
and U4053 (N_4053,N_3954,N_3984);
xor U4054 (N_4054,N_3908,N_3905);
nor U4055 (N_4055,N_3961,N_3912);
or U4056 (N_4056,N_3952,N_3938);
nand U4057 (N_4057,N_3998,N_3928);
nor U4058 (N_4058,N_3906,N_3920);
nor U4059 (N_4059,N_3921,N_3904);
or U4060 (N_4060,N_3998,N_3933);
or U4061 (N_4061,N_3903,N_3993);
and U4062 (N_4062,N_3925,N_3959);
xnor U4063 (N_4063,N_3967,N_3922);
nor U4064 (N_4064,N_3972,N_3909);
nor U4065 (N_4065,N_3939,N_3999);
nor U4066 (N_4066,N_3964,N_3977);
nand U4067 (N_4067,N_3966,N_3982);
nor U4068 (N_4068,N_3977,N_3956);
or U4069 (N_4069,N_3996,N_3966);
nand U4070 (N_4070,N_3963,N_3919);
xnor U4071 (N_4071,N_3991,N_3920);
nand U4072 (N_4072,N_3957,N_3982);
and U4073 (N_4073,N_3967,N_3914);
nor U4074 (N_4074,N_3903,N_3989);
and U4075 (N_4075,N_3916,N_3940);
or U4076 (N_4076,N_3990,N_3961);
nand U4077 (N_4077,N_3982,N_3952);
nor U4078 (N_4078,N_3924,N_3921);
nand U4079 (N_4079,N_3983,N_3931);
nand U4080 (N_4080,N_3956,N_3992);
nor U4081 (N_4081,N_3925,N_3906);
xnor U4082 (N_4082,N_3975,N_3927);
xnor U4083 (N_4083,N_3991,N_3945);
nor U4084 (N_4084,N_3951,N_3957);
nand U4085 (N_4085,N_3941,N_3975);
xor U4086 (N_4086,N_3949,N_3906);
xor U4087 (N_4087,N_3979,N_3999);
nand U4088 (N_4088,N_3976,N_3929);
nor U4089 (N_4089,N_3944,N_3911);
xnor U4090 (N_4090,N_3907,N_3990);
xor U4091 (N_4091,N_3988,N_3936);
nor U4092 (N_4092,N_3984,N_3964);
nor U4093 (N_4093,N_3990,N_3981);
nand U4094 (N_4094,N_3910,N_3993);
nand U4095 (N_4095,N_3984,N_3988);
and U4096 (N_4096,N_3958,N_3967);
nor U4097 (N_4097,N_3903,N_3943);
or U4098 (N_4098,N_3960,N_3924);
or U4099 (N_4099,N_3970,N_3962);
xor U4100 (N_4100,N_4056,N_4085);
and U4101 (N_4101,N_4026,N_4042);
nand U4102 (N_4102,N_4006,N_4064);
nand U4103 (N_4103,N_4054,N_4076);
and U4104 (N_4104,N_4019,N_4034);
or U4105 (N_4105,N_4015,N_4000);
nor U4106 (N_4106,N_4066,N_4024);
nor U4107 (N_4107,N_4005,N_4004);
xor U4108 (N_4108,N_4047,N_4014);
and U4109 (N_4109,N_4091,N_4067);
and U4110 (N_4110,N_4025,N_4074);
nor U4111 (N_4111,N_4037,N_4075);
or U4112 (N_4112,N_4045,N_4063);
nand U4113 (N_4113,N_4093,N_4071);
and U4114 (N_4114,N_4028,N_4048);
or U4115 (N_4115,N_4090,N_4013);
nor U4116 (N_4116,N_4009,N_4084);
nor U4117 (N_4117,N_4046,N_4082);
xnor U4118 (N_4118,N_4031,N_4052);
nor U4119 (N_4119,N_4007,N_4057);
and U4120 (N_4120,N_4043,N_4092);
xor U4121 (N_4121,N_4053,N_4080);
nor U4122 (N_4122,N_4001,N_4039);
nor U4123 (N_4123,N_4088,N_4073);
and U4124 (N_4124,N_4017,N_4069);
xor U4125 (N_4125,N_4035,N_4072);
nand U4126 (N_4126,N_4018,N_4065);
or U4127 (N_4127,N_4038,N_4041);
nor U4128 (N_4128,N_4081,N_4083);
and U4129 (N_4129,N_4099,N_4036);
or U4130 (N_4130,N_4087,N_4050);
nor U4131 (N_4131,N_4094,N_4098);
nor U4132 (N_4132,N_4020,N_4002);
nor U4133 (N_4133,N_4077,N_4062);
nor U4134 (N_4134,N_4027,N_4061);
nor U4135 (N_4135,N_4079,N_4070);
and U4136 (N_4136,N_4023,N_4089);
or U4137 (N_4137,N_4016,N_4044);
or U4138 (N_4138,N_4049,N_4032);
nor U4139 (N_4139,N_4095,N_4086);
nand U4140 (N_4140,N_4033,N_4059);
nand U4141 (N_4141,N_4097,N_4029);
nand U4142 (N_4142,N_4022,N_4011);
or U4143 (N_4143,N_4051,N_4030);
nand U4144 (N_4144,N_4008,N_4055);
nor U4145 (N_4145,N_4010,N_4012);
nor U4146 (N_4146,N_4068,N_4021);
xnor U4147 (N_4147,N_4040,N_4096);
or U4148 (N_4148,N_4060,N_4003);
xor U4149 (N_4149,N_4078,N_4058);
nor U4150 (N_4150,N_4048,N_4049);
nor U4151 (N_4151,N_4057,N_4010);
xor U4152 (N_4152,N_4031,N_4058);
or U4153 (N_4153,N_4054,N_4015);
nor U4154 (N_4154,N_4073,N_4089);
or U4155 (N_4155,N_4006,N_4038);
or U4156 (N_4156,N_4059,N_4029);
nand U4157 (N_4157,N_4088,N_4056);
and U4158 (N_4158,N_4051,N_4045);
and U4159 (N_4159,N_4097,N_4066);
xnor U4160 (N_4160,N_4075,N_4021);
nor U4161 (N_4161,N_4013,N_4029);
and U4162 (N_4162,N_4082,N_4022);
nand U4163 (N_4163,N_4032,N_4020);
nor U4164 (N_4164,N_4009,N_4000);
or U4165 (N_4165,N_4039,N_4052);
nand U4166 (N_4166,N_4038,N_4095);
and U4167 (N_4167,N_4072,N_4081);
and U4168 (N_4168,N_4086,N_4096);
xnor U4169 (N_4169,N_4061,N_4011);
xnor U4170 (N_4170,N_4050,N_4035);
xor U4171 (N_4171,N_4065,N_4061);
nor U4172 (N_4172,N_4030,N_4087);
nand U4173 (N_4173,N_4093,N_4021);
nor U4174 (N_4174,N_4036,N_4021);
and U4175 (N_4175,N_4037,N_4098);
or U4176 (N_4176,N_4072,N_4059);
xor U4177 (N_4177,N_4083,N_4089);
or U4178 (N_4178,N_4061,N_4022);
xnor U4179 (N_4179,N_4010,N_4039);
and U4180 (N_4180,N_4052,N_4063);
and U4181 (N_4181,N_4011,N_4040);
nor U4182 (N_4182,N_4086,N_4044);
xor U4183 (N_4183,N_4034,N_4082);
or U4184 (N_4184,N_4072,N_4033);
or U4185 (N_4185,N_4087,N_4022);
nor U4186 (N_4186,N_4083,N_4009);
or U4187 (N_4187,N_4028,N_4082);
or U4188 (N_4188,N_4031,N_4088);
and U4189 (N_4189,N_4086,N_4010);
nor U4190 (N_4190,N_4020,N_4061);
xnor U4191 (N_4191,N_4017,N_4026);
or U4192 (N_4192,N_4020,N_4087);
xnor U4193 (N_4193,N_4007,N_4084);
xor U4194 (N_4194,N_4063,N_4005);
nor U4195 (N_4195,N_4029,N_4031);
xor U4196 (N_4196,N_4043,N_4087);
nor U4197 (N_4197,N_4052,N_4081);
and U4198 (N_4198,N_4005,N_4079);
nand U4199 (N_4199,N_4041,N_4003);
or U4200 (N_4200,N_4124,N_4175);
nor U4201 (N_4201,N_4122,N_4168);
xnor U4202 (N_4202,N_4162,N_4189);
nand U4203 (N_4203,N_4135,N_4178);
nand U4204 (N_4204,N_4113,N_4126);
or U4205 (N_4205,N_4153,N_4125);
and U4206 (N_4206,N_4185,N_4106);
nor U4207 (N_4207,N_4105,N_4161);
and U4208 (N_4208,N_4128,N_4154);
xnor U4209 (N_4209,N_4192,N_4197);
and U4210 (N_4210,N_4134,N_4163);
xnor U4211 (N_4211,N_4127,N_4101);
or U4212 (N_4212,N_4144,N_4182);
nor U4213 (N_4213,N_4167,N_4119);
nor U4214 (N_4214,N_4160,N_4100);
nor U4215 (N_4215,N_4142,N_4186);
and U4216 (N_4216,N_4117,N_4133);
nand U4217 (N_4217,N_4151,N_4136);
nand U4218 (N_4218,N_4174,N_4116);
or U4219 (N_4219,N_4103,N_4183);
or U4220 (N_4220,N_4169,N_4152);
nor U4221 (N_4221,N_4145,N_4199);
or U4222 (N_4222,N_4176,N_4165);
xnor U4223 (N_4223,N_4157,N_4111);
or U4224 (N_4224,N_4188,N_4121);
xor U4225 (N_4225,N_4141,N_4147);
nor U4226 (N_4226,N_4173,N_4109);
or U4227 (N_4227,N_4158,N_4179);
or U4228 (N_4228,N_4143,N_4139);
nand U4229 (N_4229,N_4150,N_4120);
nand U4230 (N_4230,N_4123,N_4164);
and U4231 (N_4231,N_4132,N_4156);
xor U4232 (N_4232,N_4115,N_4102);
nor U4233 (N_4233,N_4130,N_4131);
xor U4234 (N_4234,N_4180,N_4170);
nor U4235 (N_4235,N_4110,N_4198);
xnor U4236 (N_4236,N_4172,N_4193);
xnor U4237 (N_4237,N_4155,N_4146);
xnor U4238 (N_4238,N_4171,N_4114);
or U4239 (N_4239,N_4194,N_4177);
xor U4240 (N_4240,N_4112,N_4159);
nand U4241 (N_4241,N_4137,N_4129);
or U4242 (N_4242,N_4140,N_4104);
xnor U4243 (N_4243,N_4190,N_4138);
or U4244 (N_4244,N_4187,N_4108);
nand U4245 (N_4245,N_4166,N_4107);
and U4246 (N_4246,N_4195,N_4149);
nor U4247 (N_4247,N_4196,N_4118);
nor U4248 (N_4248,N_4148,N_4184);
xor U4249 (N_4249,N_4181,N_4191);
and U4250 (N_4250,N_4109,N_4137);
nand U4251 (N_4251,N_4164,N_4140);
and U4252 (N_4252,N_4164,N_4167);
nor U4253 (N_4253,N_4131,N_4103);
xor U4254 (N_4254,N_4128,N_4184);
nor U4255 (N_4255,N_4172,N_4188);
nor U4256 (N_4256,N_4139,N_4190);
xnor U4257 (N_4257,N_4126,N_4172);
xor U4258 (N_4258,N_4124,N_4151);
nand U4259 (N_4259,N_4107,N_4112);
and U4260 (N_4260,N_4131,N_4176);
or U4261 (N_4261,N_4177,N_4179);
xor U4262 (N_4262,N_4153,N_4194);
nor U4263 (N_4263,N_4117,N_4118);
or U4264 (N_4264,N_4130,N_4172);
xnor U4265 (N_4265,N_4144,N_4123);
or U4266 (N_4266,N_4183,N_4195);
nand U4267 (N_4267,N_4102,N_4178);
nor U4268 (N_4268,N_4113,N_4119);
and U4269 (N_4269,N_4168,N_4157);
nor U4270 (N_4270,N_4138,N_4108);
or U4271 (N_4271,N_4185,N_4137);
nor U4272 (N_4272,N_4124,N_4188);
nor U4273 (N_4273,N_4104,N_4186);
and U4274 (N_4274,N_4148,N_4175);
or U4275 (N_4275,N_4117,N_4163);
or U4276 (N_4276,N_4185,N_4103);
nand U4277 (N_4277,N_4153,N_4120);
xnor U4278 (N_4278,N_4180,N_4188);
and U4279 (N_4279,N_4110,N_4199);
nor U4280 (N_4280,N_4186,N_4128);
or U4281 (N_4281,N_4170,N_4182);
nand U4282 (N_4282,N_4135,N_4164);
and U4283 (N_4283,N_4191,N_4106);
nor U4284 (N_4284,N_4114,N_4192);
xnor U4285 (N_4285,N_4144,N_4164);
and U4286 (N_4286,N_4168,N_4117);
and U4287 (N_4287,N_4184,N_4121);
or U4288 (N_4288,N_4122,N_4151);
and U4289 (N_4289,N_4151,N_4144);
nand U4290 (N_4290,N_4165,N_4121);
xnor U4291 (N_4291,N_4185,N_4128);
or U4292 (N_4292,N_4158,N_4153);
xor U4293 (N_4293,N_4197,N_4115);
and U4294 (N_4294,N_4151,N_4198);
or U4295 (N_4295,N_4180,N_4166);
or U4296 (N_4296,N_4151,N_4111);
nor U4297 (N_4297,N_4124,N_4101);
or U4298 (N_4298,N_4105,N_4193);
and U4299 (N_4299,N_4103,N_4191);
xor U4300 (N_4300,N_4220,N_4257);
and U4301 (N_4301,N_4236,N_4278);
or U4302 (N_4302,N_4281,N_4201);
and U4303 (N_4303,N_4210,N_4294);
and U4304 (N_4304,N_4237,N_4226);
and U4305 (N_4305,N_4268,N_4297);
xor U4306 (N_4306,N_4252,N_4285);
or U4307 (N_4307,N_4258,N_4263);
and U4308 (N_4308,N_4235,N_4261);
nand U4309 (N_4309,N_4292,N_4229);
nand U4310 (N_4310,N_4290,N_4291);
nand U4311 (N_4311,N_4203,N_4205);
and U4312 (N_4312,N_4223,N_4260);
nand U4313 (N_4313,N_4286,N_4299);
and U4314 (N_4314,N_4295,N_4274);
nand U4315 (N_4315,N_4250,N_4200);
xor U4316 (N_4316,N_4206,N_4249);
and U4317 (N_4317,N_4224,N_4244);
nand U4318 (N_4318,N_4221,N_4230);
and U4319 (N_4319,N_4298,N_4233);
nand U4320 (N_4320,N_4219,N_4264);
nand U4321 (N_4321,N_4265,N_4251);
or U4322 (N_4322,N_4241,N_4288);
xor U4323 (N_4323,N_4208,N_4202);
or U4324 (N_4324,N_4246,N_4267);
or U4325 (N_4325,N_4283,N_4204);
nand U4326 (N_4326,N_4289,N_4216);
nand U4327 (N_4327,N_4214,N_4217);
nand U4328 (N_4328,N_4245,N_4287);
nor U4329 (N_4329,N_4272,N_4227);
or U4330 (N_4330,N_4222,N_4215);
nand U4331 (N_4331,N_4228,N_4273);
nor U4332 (N_4332,N_4266,N_4243);
xor U4333 (N_4333,N_4212,N_4240);
or U4334 (N_4334,N_4262,N_4270);
or U4335 (N_4335,N_4209,N_4234);
and U4336 (N_4336,N_4253,N_4231);
or U4337 (N_4337,N_4275,N_4279);
nor U4338 (N_4338,N_4211,N_4277);
and U4339 (N_4339,N_4242,N_4269);
nor U4340 (N_4340,N_4282,N_4256);
xor U4341 (N_4341,N_4296,N_4213);
xor U4342 (N_4342,N_4218,N_4284);
xor U4343 (N_4343,N_4248,N_4280);
nand U4344 (N_4344,N_4225,N_4293);
and U4345 (N_4345,N_4254,N_4207);
nor U4346 (N_4346,N_4232,N_4238);
and U4347 (N_4347,N_4259,N_4247);
and U4348 (N_4348,N_4255,N_4276);
xnor U4349 (N_4349,N_4239,N_4271);
or U4350 (N_4350,N_4247,N_4296);
nand U4351 (N_4351,N_4285,N_4261);
nor U4352 (N_4352,N_4280,N_4263);
xnor U4353 (N_4353,N_4296,N_4255);
and U4354 (N_4354,N_4272,N_4203);
and U4355 (N_4355,N_4229,N_4271);
nand U4356 (N_4356,N_4267,N_4239);
or U4357 (N_4357,N_4253,N_4212);
nand U4358 (N_4358,N_4282,N_4285);
xnor U4359 (N_4359,N_4246,N_4231);
nand U4360 (N_4360,N_4204,N_4293);
and U4361 (N_4361,N_4216,N_4263);
nand U4362 (N_4362,N_4243,N_4280);
nor U4363 (N_4363,N_4206,N_4290);
or U4364 (N_4364,N_4212,N_4223);
and U4365 (N_4365,N_4223,N_4279);
or U4366 (N_4366,N_4258,N_4252);
xnor U4367 (N_4367,N_4251,N_4218);
or U4368 (N_4368,N_4209,N_4278);
nor U4369 (N_4369,N_4213,N_4227);
and U4370 (N_4370,N_4239,N_4255);
or U4371 (N_4371,N_4208,N_4225);
or U4372 (N_4372,N_4297,N_4205);
nand U4373 (N_4373,N_4234,N_4203);
or U4374 (N_4374,N_4298,N_4241);
and U4375 (N_4375,N_4220,N_4245);
xnor U4376 (N_4376,N_4233,N_4260);
nor U4377 (N_4377,N_4278,N_4231);
and U4378 (N_4378,N_4211,N_4289);
nand U4379 (N_4379,N_4236,N_4258);
or U4380 (N_4380,N_4298,N_4212);
and U4381 (N_4381,N_4296,N_4222);
nor U4382 (N_4382,N_4290,N_4232);
nor U4383 (N_4383,N_4200,N_4263);
nor U4384 (N_4384,N_4293,N_4256);
nand U4385 (N_4385,N_4283,N_4274);
xnor U4386 (N_4386,N_4254,N_4222);
and U4387 (N_4387,N_4266,N_4205);
xor U4388 (N_4388,N_4236,N_4282);
xnor U4389 (N_4389,N_4235,N_4296);
nor U4390 (N_4390,N_4218,N_4230);
xnor U4391 (N_4391,N_4231,N_4243);
nand U4392 (N_4392,N_4227,N_4223);
and U4393 (N_4393,N_4221,N_4265);
and U4394 (N_4394,N_4280,N_4235);
or U4395 (N_4395,N_4264,N_4272);
nor U4396 (N_4396,N_4287,N_4212);
nand U4397 (N_4397,N_4229,N_4233);
nand U4398 (N_4398,N_4223,N_4271);
or U4399 (N_4399,N_4257,N_4214);
nand U4400 (N_4400,N_4340,N_4360);
and U4401 (N_4401,N_4377,N_4324);
xnor U4402 (N_4402,N_4396,N_4373);
nand U4403 (N_4403,N_4332,N_4342);
nand U4404 (N_4404,N_4326,N_4375);
nand U4405 (N_4405,N_4321,N_4305);
or U4406 (N_4406,N_4381,N_4329);
nand U4407 (N_4407,N_4341,N_4389);
and U4408 (N_4408,N_4334,N_4315);
nor U4409 (N_4409,N_4346,N_4313);
and U4410 (N_4410,N_4322,N_4367);
and U4411 (N_4411,N_4333,N_4309);
nor U4412 (N_4412,N_4314,N_4331);
nor U4413 (N_4413,N_4385,N_4301);
nor U4414 (N_4414,N_4368,N_4393);
or U4415 (N_4415,N_4383,N_4353);
nand U4416 (N_4416,N_4372,N_4366);
and U4417 (N_4417,N_4387,N_4356);
xor U4418 (N_4418,N_4330,N_4394);
nor U4419 (N_4419,N_4398,N_4318);
nand U4420 (N_4420,N_4312,N_4308);
and U4421 (N_4421,N_4364,N_4316);
nand U4422 (N_4422,N_4325,N_4350);
xnor U4423 (N_4423,N_4397,N_4344);
nand U4424 (N_4424,N_4358,N_4378);
nand U4425 (N_4425,N_4300,N_4328);
or U4426 (N_4426,N_4370,N_4369);
nor U4427 (N_4427,N_4319,N_4382);
and U4428 (N_4428,N_4302,N_4371);
or U4429 (N_4429,N_4336,N_4338);
xor U4430 (N_4430,N_4395,N_4359);
nand U4431 (N_4431,N_4380,N_4354);
xnor U4432 (N_4432,N_4392,N_4391);
nand U4433 (N_4433,N_4365,N_4339);
nor U4434 (N_4434,N_4399,N_4390);
and U4435 (N_4435,N_4310,N_4327);
xnor U4436 (N_4436,N_4352,N_4347);
or U4437 (N_4437,N_4307,N_4343);
or U4438 (N_4438,N_4337,N_4317);
and U4439 (N_4439,N_4374,N_4355);
or U4440 (N_4440,N_4388,N_4363);
and U4441 (N_4441,N_4304,N_4349);
nand U4442 (N_4442,N_4386,N_4303);
nor U4443 (N_4443,N_4379,N_4335);
nand U4444 (N_4444,N_4323,N_4376);
nand U4445 (N_4445,N_4320,N_4351);
nor U4446 (N_4446,N_4361,N_4311);
nor U4447 (N_4447,N_4362,N_4348);
nand U4448 (N_4448,N_4306,N_4384);
nor U4449 (N_4449,N_4345,N_4357);
nand U4450 (N_4450,N_4336,N_4366);
xor U4451 (N_4451,N_4324,N_4367);
and U4452 (N_4452,N_4306,N_4378);
nor U4453 (N_4453,N_4374,N_4347);
or U4454 (N_4454,N_4389,N_4394);
nand U4455 (N_4455,N_4322,N_4313);
nor U4456 (N_4456,N_4343,N_4321);
nand U4457 (N_4457,N_4312,N_4371);
and U4458 (N_4458,N_4398,N_4356);
nand U4459 (N_4459,N_4337,N_4391);
xnor U4460 (N_4460,N_4379,N_4350);
and U4461 (N_4461,N_4397,N_4332);
or U4462 (N_4462,N_4327,N_4321);
xor U4463 (N_4463,N_4324,N_4360);
and U4464 (N_4464,N_4355,N_4319);
nor U4465 (N_4465,N_4376,N_4328);
or U4466 (N_4466,N_4328,N_4388);
or U4467 (N_4467,N_4376,N_4370);
xor U4468 (N_4468,N_4374,N_4376);
and U4469 (N_4469,N_4387,N_4336);
nor U4470 (N_4470,N_4365,N_4342);
or U4471 (N_4471,N_4346,N_4304);
nand U4472 (N_4472,N_4338,N_4378);
nor U4473 (N_4473,N_4371,N_4374);
or U4474 (N_4474,N_4398,N_4330);
or U4475 (N_4475,N_4362,N_4340);
nor U4476 (N_4476,N_4321,N_4399);
nor U4477 (N_4477,N_4386,N_4375);
nand U4478 (N_4478,N_4360,N_4389);
or U4479 (N_4479,N_4384,N_4341);
xnor U4480 (N_4480,N_4313,N_4369);
nand U4481 (N_4481,N_4313,N_4304);
nand U4482 (N_4482,N_4304,N_4316);
and U4483 (N_4483,N_4376,N_4324);
nand U4484 (N_4484,N_4358,N_4341);
and U4485 (N_4485,N_4313,N_4363);
nor U4486 (N_4486,N_4384,N_4327);
and U4487 (N_4487,N_4395,N_4310);
nand U4488 (N_4488,N_4353,N_4384);
nor U4489 (N_4489,N_4340,N_4335);
nor U4490 (N_4490,N_4312,N_4350);
and U4491 (N_4491,N_4394,N_4318);
nand U4492 (N_4492,N_4319,N_4373);
nor U4493 (N_4493,N_4331,N_4302);
or U4494 (N_4494,N_4392,N_4316);
or U4495 (N_4495,N_4376,N_4357);
and U4496 (N_4496,N_4332,N_4336);
nand U4497 (N_4497,N_4320,N_4333);
nor U4498 (N_4498,N_4378,N_4339);
xnor U4499 (N_4499,N_4323,N_4345);
or U4500 (N_4500,N_4407,N_4423);
nor U4501 (N_4501,N_4485,N_4484);
nor U4502 (N_4502,N_4413,N_4489);
nand U4503 (N_4503,N_4471,N_4480);
and U4504 (N_4504,N_4454,N_4482);
nor U4505 (N_4505,N_4488,N_4462);
nor U4506 (N_4506,N_4494,N_4401);
nand U4507 (N_4507,N_4479,N_4490);
nand U4508 (N_4508,N_4461,N_4436);
nand U4509 (N_4509,N_4404,N_4425);
xnor U4510 (N_4510,N_4476,N_4492);
nand U4511 (N_4511,N_4409,N_4410);
nor U4512 (N_4512,N_4431,N_4403);
and U4513 (N_4513,N_4496,N_4438);
or U4514 (N_4514,N_4405,N_4415);
xnor U4515 (N_4515,N_4495,N_4458);
or U4516 (N_4516,N_4427,N_4439);
and U4517 (N_4517,N_4422,N_4419);
and U4518 (N_4518,N_4420,N_4466);
nor U4519 (N_4519,N_4448,N_4414);
nand U4520 (N_4520,N_4478,N_4464);
nor U4521 (N_4521,N_4441,N_4468);
nand U4522 (N_4522,N_4408,N_4450);
and U4523 (N_4523,N_4412,N_4421);
and U4524 (N_4524,N_4446,N_4470);
nand U4525 (N_4525,N_4474,N_4444);
nor U4526 (N_4526,N_4497,N_4445);
or U4527 (N_4527,N_4437,N_4428);
or U4528 (N_4528,N_4467,N_4440);
and U4529 (N_4529,N_4416,N_4477);
or U4530 (N_4530,N_4481,N_4430);
and U4531 (N_4531,N_4447,N_4465);
nor U4532 (N_4532,N_4463,N_4498);
nand U4533 (N_4533,N_4426,N_4491);
or U4534 (N_4534,N_4487,N_4455);
xor U4535 (N_4535,N_4493,N_4456);
nand U4536 (N_4536,N_4434,N_4499);
nand U4537 (N_4537,N_4418,N_4453);
xnor U4538 (N_4538,N_4459,N_4435);
and U4539 (N_4539,N_4472,N_4433);
xnor U4540 (N_4540,N_4473,N_4411);
or U4541 (N_4541,N_4457,N_4475);
and U4542 (N_4542,N_4443,N_4469);
and U4543 (N_4543,N_4417,N_4486);
xnor U4544 (N_4544,N_4400,N_4429);
and U4545 (N_4545,N_4406,N_4452);
nor U4546 (N_4546,N_4451,N_4432);
or U4547 (N_4547,N_4483,N_4442);
nand U4548 (N_4548,N_4460,N_4424);
nor U4549 (N_4549,N_4402,N_4449);
nor U4550 (N_4550,N_4452,N_4404);
nand U4551 (N_4551,N_4491,N_4463);
or U4552 (N_4552,N_4454,N_4446);
nor U4553 (N_4553,N_4465,N_4467);
nor U4554 (N_4554,N_4458,N_4438);
nor U4555 (N_4555,N_4438,N_4430);
and U4556 (N_4556,N_4415,N_4489);
or U4557 (N_4557,N_4447,N_4424);
or U4558 (N_4558,N_4463,N_4479);
or U4559 (N_4559,N_4469,N_4476);
or U4560 (N_4560,N_4441,N_4401);
xor U4561 (N_4561,N_4426,N_4466);
or U4562 (N_4562,N_4486,N_4419);
nor U4563 (N_4563,N_4464,N_4445);
and U4564 (N_4564,N_4403,N_4442);
xor U4565 (N_4565,N_4411,N_4446);
nand U4566 (N_4566,N_4429,N_4418);
and U4567 (N_4567,N_4493,N_4402);
or U4568 (N_4568,N_4440,N_4402);
xor U4569 (N_4569,N_4479,N_4409);
and U4570 (N_4570,N_4458,N_4421);
and U4571 (N_4571,N_4490,N_4455);
xnor U4572 (N_4572,N_4417,N_4490);
xor U4573 (N_4573,N_4499,N_4424);
or U4574 (N_4574,N_4429,N_4473);
nand U4575 (N_4575,N_4486,N_4446);
nand U4576 (N_4576,N_4477,N_4495);
or U4577 (N_4577,N_4411,N_4429);
and U4578 (N_4578,N_4406,N_4401);
xor U4579 (N_4579,N_4474,N_4469);
and U4580 (N_4580,N_4468,N_4480);
nor U4581 (N_4581,N_4483,N_4405);
xnor U4582 (N_4582,N_4479,N_4476);
nand U4583 (N_4583,N_4447,N_4421);
nor U4584 (N_4584,N_4458,N_4449);
or U4585 (N_4585,N_4420,N_4495);
and U4586 (N_4586,N_4499,N_4444);
nor U4587 (N_4587,N_4403,N_4416);
xnor U4588 (N_4588,N_4486,N_4412);
nand U4589 (N_4589,N_4457,N_4437);
nor U4590 (N_4590,N_4477,N_4451);
nor U4591 (N_4591,N_4442,N_4462);
nand U4592 (N_4592,N_4432,N_4438);
xor U4593 (N_4593,N_4458,N_4451);
and U4594 (N_4594,N_4451,N_4444);
xor U4595 (N_4595,N_4461,N_4422);
or U4596 (N_4596,N_4493,N_4499);
or U4597 (N_4597,N_4491,N_4452);
xnor U4598 (N_4598,N_4471,N_4429);
nand U4599 (N_4599,N_4498,N_4405);
and U4600 (N_4600,N_4506,N_4525);
and U4601 (N_4601,N_4557,N_4591);
nor U4602 (N_4602,N_4544,N_4594);
nand U4603 (N_4603,N_4555,N_4562);
or U4604 (N_4604,N_4598,N_4567);
nor U4605 (N_4605,N_4595,N_4512);
xnor U4606 (N_4606,N_4530,N_4560);
nand U4607 (N_4607,N_4569,N_4574);
xor U4608 (N_4608,N_4552,N_4582);
and U4609 (N_4609,N_4540,N_4536);
nor U4610 (N_4610,N_4563,N_4593);
and U4611 (N_4611,N_4527,N_4502);
xor U4612 (N_4612,N_4577,N_4568);
or U4613 (N_4613,N_4592,N_4546);
xor U4614 (N_4614,N_4551,N_4597);
xor U4615 (N_4615,N_4514,N_4545);
xor U4616 (N_4616,N_4583,N_4505);
xnor U4617 (N_4617,N_4541,N_4570);
and U4618 (N_4618,N_4504,N_4585);
nor U4619 (N_4619,N_4571,N_4538);
xor U4620 (N_4620,N_4501,N_4559);
nor U4621 (N_4621,N_4547,N_4579);
nor U4622 (N_4622,N_4510,N_4507);
nand U4623 (N_4623,N_4556,N_4573);
nand U4624 (N_4624,N_4586,N_4508);
nand U4625 (N_4625,N_4529,N_4519);
xnor U4626 (N_4626,N_4500,N_4539);
or U4627 (N_4627,N_4587,N_4542);
nor U4628 (N_4628,N_4564,N_4599);
nor U4629 (N_4629,N_4581,N_4589);
nor U4630 (N_4630,N_4575,N_4553);
or U4631 (N_4631,N_4503,N_4523);
and U4632 (N_4632,N_4543,N_4532);
xnor U4633 (N_4633,N_4537,N_4550);
nor U4634 (N_4634,N_4549,N_4566);
xnor U4635 (N_4635,N_4520,N_4535);
nor U4636 (N_4636,N_4572,N_4511);
or U4637 (N_4637,N_4565,N_4518);
and U4638 (N_4638,N_4524,N_4534);
or U4639 (N_4639,N_4516,N_4513);
and U4640 (N_4640,N_4517,N_4548);
nor U4641 (N_4641,N_4580,N_4588);
nor U4642 (N_4642,N_4533,N_4521);
nand U4643 (N_4643,N_4561,N_4578);
or U4644 (N_4644,N_4526,N_4584);
xor U4645 (N_4645,N_4596,N_4576);
or U4646 (N_4646,N_4531,N_4554);
and U4647 (N_4647,N_4528,N_4558);
and U4648 (N_4648,N_4509,N_4590);
nor U4649 (N_4649,N_4515,N_4522);
and U4650 (N_4650,N_4522,N_4588);
nor U4651 (N_4651,N_4599,N_4586);
and U4652 (N_4652,N_4518,N_4566);
or U4653 (N_4653,N_4596,N_4571);
and U4654 (N_4654,N_4595,N_4502);
nor U4655 (N_4655,N_4532,N_4508);
or U4656 (N_4656,N_4526,N_4533);
or U4657 (N_4657,N_4501,N_4574);
nor U4658 (N_4658,N_4539,N_4583);
and U4659 (N_4659,N_4514,N_4594);
xnor U4660 (N_4660,N_4507,N_4548);
xnor U4661 (N_4661,N_4537,N_4572);
nand U4662 (N_4662,N_4534,N_4543);
nor U4663 (N_4663,N_4565,N_4543);
nor U4664 (N_4664,N_4510,N_4534);
and U4665 (N_4665,N_4583,N_4585);
or U4666 (N_4666,N_4597,N_4508);
and U4667 (N_4667,N_4505,N_4517);
or U4668 (N_4668,N_4522,N_4579);
xnor U4669 (N_4669,N_4592,N_4523);
and U4670 (N_4670,N_4596,N_4562);
or U4671 (N_4671,N_4576,N_4599);
xnor U4672 (N_4672,N_4572,N_4574);
xor U4673 (N_4673,N_4553,N_4501);
xnor U4674 (N_4674,N_4598,N_4540);
xor U4675 (N_4675,N_4531,N_4549);
nand U4676 (N_4676,N_4524,N_4538);
or U4677 (N_4677,N_4575,N_4586);
nand U4678 (N_4678,N_4522,N_4536);
xor U4679 (N_4679,N_4516,N_4565);
or U4680 (N_4680,N_4553,N_4538);
xnor U4681 (N_4681,N_4551,N_4559);
xor U4682 (N_4682,N_4521,N_4565);
or U4683 (N_4683,N_4551,N_4546);
nor U4684 (N_4684,N_4560,N_4548);
and U4685 (N_4685,N_4526,N_4552);
and U4686 (N_4686,N_4525,N_4509);
nor U4687 (N_4687,N_4543,N_4511);
xnor U4688 (N_4688,N_4522,N_4541);
and U4689 (N_4689,N_4509,N_4536);
and U4690 (N_4690,N_4553,N_4543);
and U4691 (N_4691,N_4504,N_4597);
nor U4692 (N_4692,N_4548,N_4528);
and U4693 (N_4693,N_4588,N_4516);
or U4694 (N_4694,N_4505,N_4522);
nand U4695 (N_4695,N_4514,N_4528);
or U4696 (N_4696,N_4599,N_4587);
or U4697 (N_4697,N_4589,N_4540);
xnor U4698 (N_4698,N_4598,N_4559);
and U4699 (N_4699,N_4532,N_4542);
xnor U4700 (N_4700,N_4681,N_4662);
nand U4701 (N_4701,N_4693,N_4645);
or U4702 (N_4702,N_4635,N_4651);
nor U4703 (N_4703,N_4600,N_4605);
or U4704 (N_4704,N_4695,N_4668);
xor U4705 (N_4705,N_4607,N_4684);
nor U4706 (N_4706,N_4633,N_4614);
nand U4707 (N_4707,N_4661,N_4694);
nor U4708 (N_4708,N_4674,N_4613);
or U4709 (N_4709,N_4689,N_4634);
or U4710 (N_4710,N_4655,N_4618);
and U4711 (N_4711,N_4646,N_4626);
or U4712 (N_4712,N_4636,N_4680);
nor U4713 (N_4713,N_4615,N_4606);
nand U4714 (N_4714,N_4686,N_4643);
and U4715 (N_4715,N_4664,N_4624);
nand U4716 (N_4716,N_4676,N_4660);
nand U4717 (N_4717,N_4699,N_4698);
or U4718 (N_4718,N_4628,N_4673);
xnor U4719 (N_4719,N_4621,N_4677);
and U4720 (N_4720,N_4669,N_4644);
nand U4721 (N_4721,N_4640,N_4620);
nand U4722 (N_4722,N_4627,N_4666);
and U4723 (N_4723,N_4604,N_4649);
nand U4724 (N_4724,N_4617,N_4632);
or U4725 (N_4725,N_4631,N_4685);
and U4726 (N_4726,N_4637,N_4663);
nor U4727 (N_4727,N_4625,N_4641);
and U4728 (N_4728,N_4638,N_4648);
nand U4729 (N_4729,N_4678,N_4687);
or U4730 (N_4730,N_4601,N_4642);
nand U4731 (N_4731,N_4667,N_4630);
nor U4732 (N_4732,N_4658,N_4623);
nand U4733 (N_4733,N_4692,N_4653);
nand U4734 (N_4734,N_4690,N_4616);
xor U4735 (N_4735,N_4608,N_4683);
nor U4736 (N_4736,N_4682,N_4611);
nand U4737 (N_4737,N_4659,N_4612);
xor U4738 (N_4738,N_4609,N_4650);
or U4739 (N_4739,N_4691,N_4629);
nor U4740 (N_4740,N_4675,N_4652);
nor U4741 (N_4741,N_4665,N_4657);
nand U4742 (N_4742,N_4656,N_4697);
nand U4743 (N_4743,N_4679,N_4672);
nand U4744 (N_4744,N_4671,N_4610);
and U4745 (N_4745,N_4602,N_4603);
nand U4746 (N_4746,N_4670,N_4639);
and U4747 (N_4747,N_4619,N_4654);
and U4748 (N_4748,N_4688,N_4622);
and U4749 (N_4749,N_4647,N_4696);
and U4750 (N_4750,N_4637,N_4692);
and U4751 (N_4751,N_4651,N_4632);
and U4752 (N_4752,N_4600,N_4611);
nand U4753 (N_4753,N_4680,N_4624);
nand U4754 (N_4754,N_4676,N_4671);
xnor U4755 (N_4755,N_4692,N_4696);
or U4756 (N_4756,N_4630,N_4673);
or U4757 (N_4757,N_4697,N_4605);
nand U4758 (N_4758,N_4671,N_4618);
nor U4759 (N_4759,N_4681,N_4650);
nor U4760 (N_4760,N_4697,N_4613);
nand U4761 (N_4761,N_4664,N_4615);
xnor U4762 (N_4762,N_4643,N_4673);
nand U4763 (N_4763,N_4655,N_4699);
nor U4764 (N_4764,N_4631,N_4605);
and U4765 (N_4765,N_4696,N_4611);
xnor U4766 (N_4766,N_4664,N_4662);
xor U4767 (N_4767,N_4628,N_4618);
nand U4768 (N_4768,N_4623,N_4693);
nor U4769 (N_4769,N_4633,N_4668);
or U4770 (N_4770,N_4620,N_4634);
and U4771 (N_4771,N_4663,N_4692);
nand U4772 (N_4772,N_4676,N_4648);
nand U4773 (N_4773,N_4639,N_4695);
nor U4774 (N_4774,N_4600,N_4652);
xor U4775 (N_4775,N_4689,N_4616);
or U4776 (N_4776,N_4601,N_4605);
nor U4777 (N_4777,N_4611,N_4688);
and U4778 (N_4778,N_4663,N_4604);
nand U4779 (N_4779,N_4685,N_4683);
xnor U4780 (N_4780,N_4689,N_4687);
xor U4781 (N_4781,N_4654,N_4613);
nand U4782 (N_4782,N_4657,N_4696);
xnor U4783 (N_4783,N_4602,N_4676);
nor U4784 (N_4784,N_4662,N_4645);
nand U4785 (N_4785,N_4667,N_4665);
and U4786 (N_4786,N_4629,N_4662);
xor U4787 (N_4787,N_4669,N_4681);
and U4788 (N_4788,N_4679,N_4689);
nor U4789 (N_4789,N_4631,N_4681);
nor U4790 (N_4790,N_4663,N_4648);
nand U4791 (N_4791,N_4611,N_4624);
nor U4792 (N_4792,N_4648,N_4667);
xor U4793 (N_4793,N_4692,N_4620);
nor U4794 (N_4794,N_4685,N_4678);
or U4795 (N_4795,N_4631,N_4660);
or U4796 (N_4796,N_4668,N_4652);
nand U4797 (N_4797,N_4655,N_4698);
xor U4798 (N_4798,N_4660,N_4678);
nor U4799 (N_4799,N_4678,N_4663);
nand U4800 (N_4800,N_4782,N_4743);
nand U4801 (N_4801,N_4774,N_4752);
xor U4802 (N_4802,N_4799,N_4716);
and U4803 (N_4803,N_4745,N_4706);
and U4804 (N_4804,N_4797,N_4733);
xor U4805 (N_4805,N_4718,N_4777);
or U4806 (N_4806,N_4735,N_4754);
xnor U4807 (N_4807,N_4707,N_4702);
xnor U4808 (N_4808,N_4728,N_4779);
and U4809 (N_4809,N_4786,N_4776);
and U4810 (N_4810,N_4784,N_4717);
or U4811 (N_4811,N_4744,N_4762);
nor U4812 (N_4812,N_4773,N_4710);
and U4813 (N_4813,N_4704,N_4725);
and U4814 (N_4814,N_4768,N_4739);
xor U4815 (N_4815,N_4737,N_4723);
nand U4816 (N_4816,N_4787,N_4775);
nor U4817 (N_4817,N_4724,N_4793);
nand U4818 (N_4818,N_4714,N_4751);
nand U4819 (N_4819,N_4700,N_4761);
nand U4820 (N_4820,N_4713,N_4709);
or U4821 (N_4821,N_4778,N_4755);
xnor U4822 (N_4822,N_4742,N_4765);
nor U4823 (N_4823,N_4763,N_4701);
and U4824 (N_4824,N_4746,N_4727);
and U4825 (N_4825,N_4705,N_4764);
nand U4826 (N_4826,N_4790,N_4720);
nand U4827 (N_4827,N_4788,N_4740);
nor U4828 (N_4828,N_4721,N_4741);
and U4829 (N_4829,N_4760,N_4753);
and U4830 (N_4830,N_4791,N_4781);
or U4831 (N_4831,N_4708,N_4757);
and U4832 (N_4832,N_4792,N_4703);
xor U4833 (N_4833,N_4747,N_4722);
or U4834 (N_4834,N_4738,N_4772);
xnor U4835 (N_4835,N_4715,N_4748);
xor U4836 (N_4836,N_4789,N_4756);
or U4837 (N_4837,N_4759,N_4736);
nand U4838 (N_4838,N_4771,N_4785);
nor U4839 (N_4839,N_4758,N_4719);
and U4840 (N_4840,N_4734,N_4726);
nand U4841 (N_4841,N_4766,N_4712);
and U4842 (N_4842,N_4769,N_4731);
or U4843 (N_4843,N_4711,N_4795);
nand U4844 (N_4844,N_4794,N_4749);
and U4845 (N_4845,N_4729,N_4796);
nand U4846 (N_4846,N_4767,N_4780);
nand U4847 (N_4847,N_4783,N_4770);
xnor U4848 (N_4848,N_4750,N_4732);
nand U4849 (N_4849,N_4798,N_4730);
xnor U4850 (N_4850,N_4714,N_4731);
or U4851 (N_4851,N_4725,N_4767);
and U4852 (N_4852,N_4792,N_4748);
or U4853 (N_4853,N_4753,N_4733);
nand U4854 (N_4854,N_4733,N_4744);
xor U4855 (N_4855,N_4753,N_4763);
xor U4856 (N_4856,N_4709,N_4747);
nor U4857 (N_4857,N_4718,N_4771);
xnor U4858 (N_4858,N_4721,N_4719);
and U4859 (N_4859,N_4764,N_4715);
and U4860 (N_4860,N_4712,N_4774);
xnor U4861 (N_4861,N_4718,N_4745);
or U4862 (N_4862,N_4784,N_4733);
nor U4863 (N_4863,N_4735,N_4752);
and U4864 (N_4864,N_4774,N_4715);
xnor U4865 (N_4865,N_4780,N_4722);
or U4866 (N_4866,N_4715,N_4770);
and U4867 (N_4867,N_4761,N_4798);
and U4868 (N_4868,N_4744,N_4718);
xnor U4869 (N_4869,N_4754,N_4706);
nor U4870 (N_4870,N_4725,N_4765);
nor U4871 (N_4871,N_4760,N_4715);
and U4872 (N_4872,N_4747,N_4780);
nor U4873 (N_4873,N_4740,N_4771);
nor U4874 (N_4874,N_4748,N_4779);
or U4875 (N_4875,N_4730,N_4702);
nand U4876 (N_4876,N_4761,N_4724);
nor U4877 (N_4877,N_4776,N_4790);
and U4878 (N_4878,N_4701,N_4770);
nand U4879 (N_4879,N_4716,N_4705);
and U4880 (N_4880,N_4736,N_4754);
xnor U4881 (N_4881,N_4745,N_4701);
nand U4882 (N_4882,N_4734,N_4793);
nand U4883 (N_4883,N_4734,N_4747);
or U4884 (N_4884,N_4761,N_4795);
and U4885 (N_4885,N_4752,N_4715);
or U4886 (N_4886,N_4752,N_4737);
nand U4887 (N_4887,N_4750,N_4757);
and U4888 (N_4888,N_4745,N_4746);
xor U4889 (N_4889,N_4791,N_4718);
or U4890 (N_4890,N_4760,N_4723);
nand U4891 (N_4891,N_4767,N_4784);
nor U4892 (N_4892,N_4755,N_4743);
or U4893 (N_4893,N_4745,N_4738);
nand U4894 (N_4894,N_4723,N_4751);
and U4895 (N_4895,N_4766,N_4768);
xor U4896 (N_4896,N_4767,N_4751);
nor U4897 (N_4897,N_4715,N_4734);
nor U4898 (N_4898,N_4721,N_4766);
and U4899 (N_4899,N_4772,N_4791);
nor U4900 (N_4900,N_4838,N_4811);
nor U4901 (N_4901,N_4852,N_4844);
nand U4902 (N_4902,N_4881,N_4822);
xnor U4903 (N_4903,N_4856,N_4813);
or U4904 (N_4904,N_4876,N_4850);
and U4905 (N_4905,N_4834,N_4840);
xnor U4906 (N_4906,N_4863,N_4864);
and U4907 (N_4907,N_4898,N_4827);
nor U4908 (N_4908,N_4891,N_4873);
xnor U4909 (N_4909,N_4804,N_4867);
nor U4910 (N_4910,N_4824,N_4897);
xnor U4911 (N_4911,N_4814,N_4800);
or U4912 (N_4912,N_4835,N_4877);
nand U4913 (N_4913,N_4847,N_4869);
nand U4914 (N_4914,N_4888,N_4825);
and U4915 (N_4915,N_4892,N_4816);
and U4916 (N_4916,N_4870,N_4865);
xor U4917 (N_4917,N_4842,N_4801);
xor U4918 (N_4918,N_4836,N_4830);
xor U4919 (N_4919,N_4846,N_4875);
or U4920 (N_4920,N_4832,N_4872);
nor U4921 (N_4921,N_4848,N_4862);
nor U4922 (N_4922,N_4899,N_4895);
nand U4923 (N_4923,N_4805,N_4874);
or U4924 (N_4924,N_4896,N_4878);
and U4925 (N_4925,N_4860,N_4831);
xor U4926 (N_4926,N_4879,N_4871);
and U4927 (N_4927,N_4829,N_4817);
nand U4928 (N_4928,N_4808,N_4883);
and U4929 (N_4929,N_4857,N_4802);
and U4930 (N_4930,N_4884,N_4815);
nand U4931 (N_4931,N_4861,N_4843);
and U4932 (N_4932,N_4826,N_4858);
nor U4933 (N_4933,N_4807,N_4886);
nand U4934 (N_4934,N_4812,N_4820);
nand U4935 (N_4935,N_4851,N_4885);
nand U4936 (N_4936,N_4845,N_4880);
xor U4937 (N_4937,N_4806,N_4890);
nand U4938 (N_4938,N_4853,N_4849);
nand U4939 (N_4939,N_4868,N_4833);
nor U4940 (N_4940,N_4866,N_4889);
xor U4941 (N_4941,N_4841,N_4894);
or U4942 (N_4942,N_4821,N_4823);
or U4943 (N_4943,N_4828,N_4859);
xnor U4944 (N_4944,N_4818,N_4803);
and U4945 (N_4945,N_4893,N_4839);
or U4946 (N_4946,N_4855,N_4819);
and U4947 (N_4947,N_4837,N_4887);
nor U4948 (N_4948,N_4809,N_4810);
or U4949 (N_4949,N_4854,N_4882);
and U4950 (N_4950,N_4841,N_4883);
xor U4951 (N_4951,N_4840,N_4870);
and U4952 (N_4952,N_4809,N_4835);
xor U4953 (N_4953,N_4891,N_4841);
or U4954 (N_4954,N_4816,N_4884);
nand U4955 (N_4955,N_4807,N_4885);
or U4956 (N_4956,N_4816,N_4819);
or U4957 (N_4957,N_4821,N_4882);
and U4958 (N_4958,N_4887,N_4846);
and U4959 (N_4959,N_4821,N_4853);
and U4960 (N_4960,N_4832,N_4876);
or U4961 (N_4961,N_4803,N_4864);
nor U4962 (N_4962,N_4836,N_4891);
and U4963 (N_4963,N_4899,N_4844);
or U4964 (N_4964,N_4819,N_4820);
xor U4965 (N_4965,N_4807,N_4892);
nand U4966 (N_4966,N_4808,N_4835);
xnor U4967 (N_4967,N_4887,N_4824);
nor U4968 (N_4968,N_4809,N_4868);
or U4969 (N_4969,N_4867,N_4854);
or U4970 (N_4970,N_4892,N_4850);
or U4971 (N_4971,N_4842,N_4827);
or U4972 (N_4972,N_4898,N_4817);
xnor U4973 (N_4973,N_4830,N_4870);
and U4974 (N_4974,N_4883,N_4840);
xor U4975 (N_4975,N_4811,N_4831);
or U4976 (N_4976,N_4829,N_4880);
and U4977 (N_4977,N_4816,N_4893);
nand U4978 (N_4978,N_4893,N_4837);
and U4979 (N_4979,N_4821,N_4819);
or U4980 (N_4980,N_4893,N_4874);
nor U4981 (N_4981,N_4866,N_4816);
and U4982 (N_4982,N_4831,N_4814);
xnor U4983 (N_4983,N_4824,N_4878);
nor U4984 (N_4984,N_4810,N_4811);
xnor U4985 (N_4985,N_4893,N_4824);
and U4986 (N_4986,N_4832,N_4818);
nor U4987 (N_4987,N_4822,N_4837);
xnor U4988 (N_4988,N_4838,N_4832);
nand U4989 (N_4989,N_4808,N_4878);
nand U4990 (N_4990,N_4813,N_4833);
nand U4991 (N_4991,N_4832,N_4899);
xnor U4992 (N_4992,N_4811,N_4852);
xnor U4993 (N_4993,N_4845,N_4883);
nand U4994 (N_4994,N_4896,N_4867);
nand U4995 (N_4995,N_4869,N_4842);
xnor U4996 (N_4996,N_4872,N_4830);
nand U4997 (N_4997,N_4874,N_4850);
and U4998 (N_4998,N_4867,N_4838);
xnor U4999 (N_4999,N_4884,N_4890);
nand U5000 (N_5000,N_4933,N_4960);
and U5001 (N_5001,N_4977,N_4934);
or U5002 (N_5002,N_4940,N_4908);
or U5003 (N_5003,N_4913,N_4956);
xor U5004 (N_5004,N_4937,N_4950);
xnor U5005 (N_5005,N_4967,N_4927);
nand U5006 (N_5006,N_4915,N_4961);
nand U5007 (N_5007,N_4947,N_4918);
and U5008 (N_5008,N_4952,N_4968);
nor U5009 (N_5009,N_4974,N_4938);
xor U5010 (N_5010,N_4944,N_4939);
or U5011 (N_5011,N_4982,N_4926);
xor U5012 (N_5012,N_4986,N_4964);
nand U5013 (N_5013,N_4997,N_4910);
nand U5014 (N_5014,N_4949,N_4920);
xnor U5015 (N_5015,N_4941,N_4923);
xnor U5016 (N_5016,N_4989,N_4995);
nor U5017 (N_5017,N_4979,N_4988);
nor U5018 (N_5018,N_4987,N_4980);
nor U5019 (N_5019,N_4901,N_4951);
xnor U5020 (N_5020,N_4978,N_4966);
and U5021 (N_5021,N_4991,N_4984);
or U5022 (N_5022,N_4921,N_4929);
nor U5023 (N_5023,N_4914,N_4962);
xnor U5024 (N_5024,N_4999,N_4975);
nor U5025 (N_5025,N_4993,N_4943);
nand U5026 (N_5026,N_4985,N_4998);
or U5027 (N_5027,N_4930,N_4983);
nor U5028 (N_5028,N_4942,N_4994);
xor U5029 (N_5029,N_4972,N_4928);
and U5030 (N_5030,N_4946,N_4903);
and U5031 (N_5031,N_4925,N_4973);
or U5032 (N_5032,N_4976,N_4924);
or U5033 (N_5033,N_4945,N_4909);
nor U5034 (N_5034,N_4996,N_4912);
nor U5035 (N_5035,N_4970,N_4907);
and U5036 (N_5036,N_4965,N_4969);
or U5037 (N_5037,N_4957,N_4922);
nand U5038 (N_5038,N_4953,N_4948);
nand U5039 (N_5039,N_4963,N_4906);
xor U5040 (N_5040,N_4905,N_4936);
nor U5041 (N_5041,N_4902,N_4990);
or U5042 (N_5042,N_4911,N_4992);
nor U5043 (N_5043,N_4900,N_4958);
xnor U5044 (N_5044,N_4955,N_4917);
nor U5045 (N_5045,N_4932,N_4904);
xnor U5046 (N_5046,N_4954,N_4981);
xnor U5047 (N_5047,N_4931,N_4959);
nor U5048 (N_5048,N_4919,N_4935);
or U5049 (N_5049,N_4971,N_4916);
nor U5050 (N_5050,N_4938,N_4947);
nand U5051 (N_5051,N_4920,N_4950);
nand U5052 (N_5052,N_4913,N_4960);
and U5053 (N_5053,N_4923,N_4983);
xnor U5054 (N_5054,N_4957,N_4966);
or U5055 (N_5055,N_4971,N_4941);
nor U5056 (N_5056,N_4924,N_4986);
xor U5057 (N_5057,N_4930,N_4910);
nand U5058 (N_5058,N_4931,N_4982);
xnor U5059 (N_5059,N_4904,N_4971);
and U5060 (N_5060,N_4906,N_4930);
xor U5061 (N_5061,N_4910,N_4994);
and U5062 (N_5062,N_4949,N_4985);
nor U5063 (N_5063,N_4981,N_4979);
nand U5064 (N_5064,N_4998,N_4920);
and U5065 (N_5065,N_4925,N_4983);
nor U5066 (N_5066,N_4950,N_4982);
and U5067 (N_5067,N_4933,N_4965);
nor U5068 (N_5068,N_4980,N_4913);
nand U5069 (N_5069,N_4976,N_4973);
and U5070 (N_5070,N_4971,N_4902);
xor U5071 (N_5071,N_4999,N_4984);
or U5072 (N_5072,N_4947,N_4902);
xor U5073 (N_5073,N_4975,N_4970);
or U5074 (N_5074,N_4912,N_4935);
xor U5075 (N_5075,N_4935,N_4932);
and U5076 (N_5076,N_4951,N_4966);
nand U5077 (N_5077,N_4969,N_4934);
and U5078 (N_5078,N_4917,N_4995);
and U5079 (N_5079,N_4936,N_4988);
nand U5080 (N_5080,N_4996,N_4966);
nand U5081 (N_5081,N_4949,N_4934);
nor U5082 (N_5082,N_4901,N_4993);
nor U5083 (N_5083,N_4978,N_4900);
and U5084 (N_5084,N_4952,N_4954);
xor U5085 (N_5085,N_4914,N_4950);
or U5086 (N_5086,N_4963,N_4954);
or U5087 (N_5087,N_4942,N_4971);
nor U5088 (N_5088,N_4926,N_4953);
nand U5089 (N_5089,N_4918,N_4933);
or U5090 (N_5090,N_4916,N_4995);
or U5091 (N_5091,N_4967,N_4966);
nand U5092 (N_5092,N_4973,N_4946);
nor U5093 (N_5093,N_4936,N_4929);
nand U5094 (N_5094,N_4947,N_4960);
nand U5095 (N_5095,N_4982,N_4981);
and U5096 (N_5096,N_4963,N_4902);
nor U5097 (N_5097,N_4959,N_4924);
xnor U5098 (N_5098,N_4935,N_4966);
xnor U5099 (N_5099,N_4926,N_4954);
or U5100 (N_5100,N_5082,N_5004);
nand U5101 (N_5101,N_5052,N_5036);
or U5102 (N_5102,N_5064,N_5041);
xnor U5103 (N_5103,N_5077,N_5057);
xor U5104 (N_5104,N_5032,N_5094);
nand U5105 (N_5105,N_5070,N_5062);
or U5106 (N_5106,N_5030,N_5002);
nor U5107 (N_5107,N_5010,N_5055);
nor U5108 (N_5108,N_5067,N_5044);
and U5109 (N_5109,N_5048,N_5013);
and U5110 (N_5110,N_5021,N_5091);
xnor U5111 (N_5111,N_5079,N_5034);
and U5112 (N_5112,N_5012,N_5072);
and U5113 (N_5113,N_5088,N_5029);
nor U5114 (N_5114,N_5066,N_5085);
or U5115 (N_5115,N_5003,N_5065);
nand U5116 (N_5116,N_5018,N_5045);
and U5117 (N_5117,N_5089,N_5001);
nand U5118 (N_5118,N_5078,N_5071);
nand U5119 (N_5119,N_5084,N_5073);
and U5120 (N_5120,N_5087,N_5043);
and U5121 (N_5121,N_5017,N_5099);
xnor U5122 (N_5122,N_5027,N_5031);
or U5123 (N_5123,N_5011,N_5015);
nand U5124 (N_5124,N_5046,N_5028);
xor U5125 (N_5125,N_5007,N_5075);
nand U5126 (N_5126,N_5093,N_5086);
or U5127 (N_5127,N_5020,N_5000);
or U5128 (N_5128,N_5054,N_5056);
nand U5129 (N_5129,N_5035,N_5005);
and U5130 (N_5130,N_5033,N_5083);
xor U5131 (N_5131,N_5042,N_5080);
nand U5132 (N_5132,N_5039,N_5060);
nand U5133 (N_5133,N_5040,N_5051);
nor U5134 (N_5134,N_5053,N_5024);
xnor U5135 (N_5135,N_5061,N_5059);
xnor U5136 (N_5136,N_5016,N_5076);
and U5137 (N_5137,N_5092,N_5074);
nand U5138 (N_5138,N_5037,N_5008);
xor U5139 (N_5139,N_5019,N_5023);
nand U5140 (N_5140,N_5025,N_5006);
nand U5141 (N_5141,N_5097,N_5022);
nand U5142 (N_5142,N_5050,N_5049);
nand U5143 (N_5143,N_5095,N_5069);
xor U5144 (N_5144,N_5063,N_5026);
nor U5145 (N_5145,N_5090,N_5096);
and U5146 (N_5146,N_5081,N_5014);
nand U5147 (N_5147,N_5038,N_5047);
nor U5148 (N_5148,N_5068,N_5009);
xor U5149 (N_5149,N_5058,N_5098);
xnor U5150 (N_5150,N_5041,N_5082);
or U5151 (N_5151,N_5048,N_5049);
nand U5152 (N_5152,N_5004,N_5073);
nand U5153 (N_5153,N_5016,N_5008);
and U5154 (N_5154,N_5011,N_5097);
and U5155 (N_5155,N_5072,N_5076);
or U5156 (N_5156,N_5007,N_5093);
nor U5157 (N_5157,N_5057,N_5025);
nor U5158 (N_5158,N_5010,N_5021);
nor U5159 (N_5159,N_5070,N_5046);
nand U5160 (N_5160,N_5068,N_5019);
nand U5161 (N_5161,N_5053,N_5046);
or U5162 (N_5162,N_5071,N_5036);
nand U5163 (N_5163,N_5064,N_5005);
nand U5164 (N_5164,N_5077,N_5052);
nor U5165 (N_5165,N_5095,N_5067);
and U5166 (N_5166,N_5063,N_5058);
nand U5167 (N_5167,N_5088,N_5052);
xor U5168 (N_5168,N_5094,N_5077);
nor U5169 (N_5169,N_5058,N_5027);
xnor U5170 (N_5170,N_5022,N_5047);
and U5171 (N_5171,N_5071,N_5067);
nor U5172 (N_5172,N_5064,N_5015);
nor U5173 (N_5173,N_5030,N_5017);
nor U5174 (N_5174,N_5058,N_5017);
nor U5175 (N_5175,N_5051,N_5037);
or U5176 (N_5176,N_5056,N_5046);
nand U5177 (N_5177,N_5048,N_5019);
and U5178 (N_5178,N_5001,N_5034);
xnor U5179 (N_5179,N_5084,N_5012);
and U5180 (N_5180,N_5092,N_5041);
or U5181 (N_5181,N_5043,N_5008);
or U5182 (N_5182,N_5035,N_5024);
or U5183 (N_5183,N_5063,N_5089);
xnor U5184 (N_5184,N_5099,N_5062);
or U5185 (N_5185,N_5029,N_5039);
xor U5186 (N_5186,N_5061,N_5078);
and U5187 (N_5187,N_5050,N_5099);
and U5188 (N_5188,N_5069,N_5021);
nor U5189 (N_5189,N_5032,N_5088);
and U5190 (N_5190,N_5045,N_5081);
or U5191 (N_5191,N_5010,N_5017);
xor U5192 (N_5192,N_5029,N_5038);
nand U5193 (N_5193,N_5040,N_5059);
xor U5194 (N_5194,N_5072,N_5047);
nor U5195 (N_5195,N_5003,N_5015);
and U5196 (N_5196,N_5064,N_5044);
or U5197 (N_5197,N_5099,N_5069);
or U5198 (N_5198,N_5030,N_5034);
or U5199 (N_5199,N_5037,N_5046);
xor U5200 (N_5200,N_5182,N_5154);
and U5201 (N_5201,N_5100,N_5128);
nor U5202 (N_5202,N_5189,N_5101);
and U5203 (N_5203,N_5193,N_5157);
or U5204 (N_5204,N_5191,N_5121);
and U5205 (N_5205,N_5141,N_5125);
nand U5206 (N_5206,N_5156,N_5116);
and U5207 (N_5207,N_5178,N_5143);
nand U5208 (N_5208,N_5151,N_5163);
xnor U5209 (N_5209,N_5166,N_5170);
xor U5210 (N_5210,N_5167,N_5175);
xnor U5211 (N_5211,N_5146,N_5152);
and U5212 (N_5212,N_5195,N_5180);
nand U5213 (N_5213,N_5155,N_5105);
nor U5214 (N_5214,N_5111,N_5169);
xnor U5215 (N_5215,N_5153,N_5177);
and U5216 (N_5216,N_5199,N_5122);
nor U5217 (N_5217,N_5132,N_5174);
xnor U5218 (N_5218,N_5119,N_5168);
and U5219 (N_5219,N_5188,N_5103);
nand U5220 (N_5220,N_5123,N_5127);
and U5221 (N_5221,N_5149,N_5131);
and U5222 (N_5222,N_5135,N_5139);
or U5223 (N_5223,N_5138,N_5120);
nand U5224 (N_5224,N_5117,N_5184);
or U5225 (N_5225,N_5161,N_5126);
or U5226 (N_5226,N_5145,N_5124);
nor U5227 (N_5227,N_5136,N_5183);
xor U5228 (N_5228,N_5194,N_5172);
nor U5229 (N_5229,N_5165,N_5187);
nor U5230 (N_5230,N_5129,N_5134);
nor U5231 (N_5231,N_5160,N_5144);
nor U5232 (N_5232,N_5162,N_5114);
nand U5233 (N_5233,N_5137,N_5107);
nor U5234 (N_5234,N_5173,N_5106);
and U5235 (N_5235,N_5102,N_5115);
nor U5236 (N_5236,N_5181,N_5185);
nor U5237 (N_5237,N_5192,N_5179);
nand U5238 (N_5238,N_5109,N_5112);
or U5239 (N_5239,N_5190,N_5140);
xor U5240 (N_5240,N_5104,N_5110);
or U5241 (N_5241,N_5186,N_5176);
xnor U5242 (N_5242,N_5133,N_5147);
nor U5243 (N_5243,N_5164,N_5130);
or U5244 (N_5244,N_5159,N_5171);
nand U5245 (N_5245,N_5108,N_5196);
nand U5246 (N_5246,N_5150,N_5148);
nor U5247 (N_5247,N_5113,N_5197);
and U5248 (N_5248,N_5158,N_5142);
or U5249 (N_5249,N_5118,N_5198);
or U5250 (N_5250,N_5199,N_5127);
and U5251 (N_5251,N_5143,N_5119);
or U5252 (N_5252,N_5136,N_5110);
and U5253 (N_5253,N_5172,N_5158);
or U5254 (N_5254,N_5162,N_5167);
nand U5255 (N_5255,N_5100,N_5184);
nand U5256 (N_5256,N_5106,N_5170);
or U5257 (N_5257,N_5137,N_5108);
nand U5258 (N_5258,N_5175,N_5100);
xor U5259 (N_5259,N_5185,N_5102);
xnor U5260 (N_5260,N_5191,N_5116);
nand U5261 (N_5261,N_5108,N_5118);
and U5262 (N_5262,N_5108,N_5105);
nor U5263 (N_5263,N_5159,N_5111);
xnor U5264 (N_5264,N_5161,N_5174);
or U5265 (N_5265,N_5125,N_5152);
xor U5266 (N_5266,N_5126,N_5107);
and U5267 (N_5267,N_5115,N_5145);
nand U5268 (N_5268,N_5162,N_5102);
nand U5269 (N_5269,N_5146,N_5131);
xor U5270 (N_5270,N_5146,N_5101);
or U5271 (N_5271,N_5110,N_5138);
xnor U5272 (N_5272,N_5137,N_5135);
and U5273 (N_5273,N_5111,N_5122);
nor U5274 (N_5274,N_5104,N_5144);
nand U5275 (N_5275,N_5196,N_5194);
and U5276 (N_5276,N_5166,N_5163);
and U5277 (N_5277,N_5130,N_5186);
and U5278 (N_5278,N_5197,N_5118);
or U5279 (N_5279,N_5151,N_5136);
or U5280 (N_5280,N_5115,N_5117);
and U5281 (N_5281,N_5110,N_5188);
or U5282 (N_5282,N_5105,N_5158);
xnor U5283 (N_5283,N_5125,N_5108);
and U5284 (N_5284,N_5124,N_5158);
or U5285 (N_5285,N_5170,N_5160);
or U5286 (N_5286,N_5155,N_5111);
or U5287 (N_5287,N_5131,N_5180);
and U5288 (N_5288,N_5171,N_5179);
nor U5289 (N_5289,N_5146,N_5148);
and U5290 (N_5290,N_5150,N_5184);
nand U5291 (N_5291,N_5194,N_5124);
nand U5292 (N_5292,N_5159,N_5160);
nor U5293 (N_5293,N_5191,N_5130);
xnor U5294 (N_5294,N_5109,N_5190);
and U5295 (N_5295,N_5106,N_5132);
or U5296 (N_5296,N_5194,N_5109);
nor U5297 (N_5297,N_5165,N_5120);
nor U5298 (N_5298,N_5172,N_5125);
and U5299 (N_5299,N_5110,N_5164);
nand U5300 (N_5300,N_5220,N_5268);
nor U5301 (N_5301,N_5246,N_5205);
nand U5302 (N_5302,N_5261,N_5248);
xnor U5303 (N_5303,N_5203,N_5207);
or U5304 (N_5304,N_5292,N_5237);
nand U5305 (N_5305,N_5286,N_5296);
xnor U5306 (N_5306,N_5210,N_5263);
xor U5307 (N_5307,N_5253,N_5249);
and U5308 (N_5308,N_5265,N_5211);
and U5309 (N_5309,N_5290,N_5272);
and U5310 (N_5310,N_5280,N_5289);
xor U5311 (N_5311,N_5262,N_5215);
nor U5312 (N_5312,N_5226,N_5206);
and U5313 (N_5313,N_5235,N_5209);
nand U5314 (N_5314,N_5297,N_5266);
and U5315 (N_5315,N_5256,N_5257);
nor U5316 (N_5316,N_5240,N_5299);
and U5317 (N_5317,N_5267,N_5239);
and U5318 (N_5318,N_5287,N_5202);
and U5319 (N_5319,N_5217,N_5204);
xnor U5320 (N_5320,N_5284,N_5278);
nor U5321 (N_5321,N_5252,N_5244);
xnor U5322 (N_5322,N_5282,N_5295);
or U5323 (N_5323,N_5255,N_5293);
xnor U5324 (N_5324,N_5258,N_5264);
nand U5325 (N_5325,N_5288,N_5283);
xor U5326 (N_5326,N_5231,N_5281);
or U5327 (N_5327,N_5270,N_5219);
nand U5328 (N_5328,N_5247,N_5277);
or U5329 (N_5329,N_5233,N_5200);
or U5330 (N_5330,N_5276,N_5298);
nor U5331 (N_5331,N_5271,N_5201);
and U5332 (N_5332,N_5228,N_5285);
or U5333 (N_5333,N_5294,N_5245);
and U5334 (N_5334,N_5251,N_5218);
xor U5335 (N_5335,N_5242,N_5250);
xnor U5336 (N_5336,N_5230,N_5269);
and U5337 (N_5337,N_5213,N_5234);
nand U5338 (N_5338,N_5274,N_5243);
or U5339 (N_5339,N_5212,N_5227);
or U5340 (N_5340,N_5229,N_5222);
and U5341 (N_5341,N_5236,N_5223);
nand U5342 (N_5342,N_5275,N_5225);
nor U5343 (N_5343,N_5232,N_5291);
and U5344 (N_5344,N_5238,N_5224);
or U5345 (N_5345,N_5214,N_5279);
and U5346 (N_5346,N_5260,N_5273);
nor U5347 (N_5347,N_5241,N_5259);
nand U5348 (N_5348,N_5216,N_5221);
nand U5349 (N_5349,N_5254,N_5208);
xor U5350 (N_5350,N_5269,N_5232);
nand U5351 (N_5351,N_5248,N_5290);
nand U5352 (N_5352,N_5226,N_5237);
nor U5353 (N_5353,N_5253,N_5230);
nand U5354 (N_5354,N_5268,N_5243);
nor U5355 (N_5355,N_5257,N_5251);
or U5356 (N_5356,N_5274,N_5264);
or U5357 (N_5357,N_5200,N_5202);
and U5358 (N_5358,N_5218,N_5223);
and U5359 (N_5359,N_5225,N_5203);
xor U5360 (N_5360,N_5253,N_5261);
xor U5361 (N_5361,N_5229,N_5209);
nand U5362 (N_5362,N_5212,N_5295);
and U5363 (N_5363,N_5235,N_5280);
nor U5364 (N_5364,N_5265,N_5230);
and U5365 (N_5365,N_5223,N_5283);
nand U5366 (N_5366,N_5299,N_5269);
nand U5367 (N_5367,N_5285,N_5247);
or U5368 (N_5368,N_5211,N_5212);
and U5369 (N_5369,N_5232,N_5295);
nand U5370 (N_5370,N_5254,N_5297);
and U5371 (N_5371,N_5284,N_5276);
nand U5372 (N_5372,N_5250,N_5257);
and U5373 (N_5373,N_5294,N_5250);
and U5374 (N_5374,N_5205,N_5268);
xnor U5375 (N_5375,N_5231,N_5267);
xor U5376 (N_5376,N_5200,N_5249);
nand U5377 (N_5377,N_5296,N_5233);
or U5378 (N_5378,N_5209,N_5291);
nor U5379 (N_5379,N_5267,N_5200);
xor U5380 (N_5380,N_5201,N_5267);
and U5381 (N_5381,N_5219,N_5231);
and U5382 (N_5382,N_5278,N_5256);
or U5383 (N_5383,N_5260,N_5220);
nand U5384 (N_5384,N_5240,N_5248);
or U5385 (N_5385,N_5213,N_5230);
nand U5386 (N_5386,N_5244,N_5212);
xor U5387 (N_5387,N_5251,N_5222);
xor U5388 (N_5388,N_5276,N_5222);
and U5389 (N_5389,N_5277,N_5242);
xor U5390 (N_5390,N_5296,N_5282);
nor U5391 (N_5391,N_5285,N_5219);
nor U5392 (N_5392,N_5249,N_5260);
nand U5393 (N_5393,N_5235,N_5269);
xnor U5394 (N_5394,N_5286,N_5249);
nor U5395 (N_5395,N_5243,N_5218);
xor U5396 (N_5396,N_5251,N_5236);
nor U5397 (N_5397,N_5215,N_5263);
xnor U5398 (N_5398,N_5266,N_5209);
xor U5399 (N_5399,N_5281,N_5283);
nor U5400 (N_5400,N_5376,N_5394);
or U5401 (N_5401,N_5320,N_5391);
xor U5402 (N_5402,N_5360,N_5301);
nor U5403 (N_5403,N_5367,N_5378);
xor U5404 (N_5404,N_5363,N_5395);
or U5405 (N_5405,N_5342,N_5302);
xnor U5406 (N_5406,N_5377,N_5331);
and U5407 (N_5407,N_5328,N_5371);
nand U5408 (N_5408,N_5312,N_5350);
xor U5409 (N_5409,N_5336,N_5348);
nor U5410 (N_5410,N_5368,N_5315);
nand U5411 (N_5411,N_5384,N_5339);
or U5412 (N_5412,N_5345,N_5399);
and U5413 (N_5413,N_5372,N_5310);
xor U5414 (N_5414,N_5313,N_5326);
xnor U5415 (N_5415,N_5323,N_5398);
and U5416 (N_5416,N_5358,N_5316);
nand U5417 (N_5417,N_5383,N_5352);
and U5418 (N_5418,N_5362,N_5396);
and U5419 (N_5419,N_5340,N_5357);
nand U5420 (N_5420,N_5341,N_5355);
xor U5421 (N_5421,N_5303,N_5351);
xor U5422 (N_5422,N_5389,N_5385);
or U5423 (N_5423,N_5318,N_5374);
or U5424 (N_5424,N_5397,N_5337);
nand U5425 (N_5425,N_5305,N_5319);
nor U5426 (N_5426,N_5364,N_5366);
and U5427 (N_5427,N_5325,N_5324);
nand U5428 (N_5428,N_5304,N_5365);
nor U5429 (N_5429,N_5300,N_5307);
xor U5430 (N_5430,N_5346,N_5322);
and U5431 (N_5431,N_5361,N_5390);
nor U5432 (N_5432,N_5317,N_5354);
and U5433 (N_5433,N_5386,N_5321);
nand U5434 (N_5434,N_5369,N_5379);
xnor U5435 (N_5435,N_5388,N_5343);
and U5436 (N_5436,N_5392,N_5334);
nor U5437 (N_5437,N_5306,N_5308);
xnor U5438 (N_5438,N_5332,N_5327);
nand U5439 (N_5439,N_5338,N_5329);
xnor U5440 (N_5440,N_5344,N_5373);
nor U5441 (N_5441,N_5393,N_5333);
xnor U5442 (N_5442,N_5353,N_5330);
or U5443 (N_5443,N_5314,N_5370);
nand U5444 (N_5444,N_5387,N_5375);
or U5445 (N_5445,N_5382,N_5380);
nor U5446 (N_5446,N_5311,N_5335);
nor U5447 (N_5447,N_5309,N_5359);
or U5448 (N_5448,N_5347,N_5349);
and U5449 (N_5449,N_5381,N_5356);
nand U5450 (N_5450,N_5385,N_5372);
nand U5451 (N_5451,N_5366,N_5319);
nand U5452 (N_5452,N_5303,N_5316);
nand U5453 (N_5453,N_5377,N_5376);
or U5454 (N_5454,N_5368,N_5369);
and U5455 (N_5455,N_5347,N_5326);
nand U5456 (N_5456,N_5349,N_5318);
nor U5457 (N_5457,N_5329,N_5303);
nor U5458 (N_5458,N_5300,N_5356);
nand U5459 (N_5459,N_5336,N_5323);
nand U5460 (N_5460,N_5390,N_5394);
and U5461 (N_5461,N_5303,N_5356);
xor U5462 (N_5462,N_5354,N_5384);
nor U5463 (N_5463,N_5305,N_5310);
nor U5464 (N_5464,N_5355,N_5368);
and U5465 (N_5465,N_5363,N_5372);
nand U5466 (N_5466,N_5399,N_5379);
xor U5467 (N_5467,N_5357,N_5341);
or U5468 (N_5468,N_5307,N_5351);
and U5469 (N_5469,N_5348,N_5355);
xnor U5470 (N_5470,N_5340,N_5367);
nand U5471 (N_5471,N_5357,N_5344);
or U5472 (N_5472,N_5380,N_5336);
and U5473 (N_5473,N_5396,N_5342);
nor U5474 (N_5474,N_5300,N_5385);
xnor U5475 (N_5475,N_5343,N_5383);
or U5476 (N_5476,N_5302,N_5330);
nand U5477 (N_5477,N_5388,N_5316);
or U5478 (N_5478,N_5331,N_5333);
and U5479 (N_5479,N_5345,N_5321);
nor U5480 (N_5480,N_5364,N_5301);
and U5481 (N_5481,N_5351,N_5387);
nand U5482 (N_5482,N_5300,N_5306);
nor U5483 (N_5483,N_5396,N_5334);
xnor U5484 (N_5484,N_5317,N_5326);
xor U5485 (N_5485,N_5302,N_5345);
nand U5486 (N_5486,N_5383,N_5363);
or U5487 (N_5487,N_5394,N_5377);
nand U5488 (N_5488,N_5333,N_5349);
or U5489 (N_5489,N_5358,N_5337);
nand U5490 (N_5490,N_5331,N_5350);
and U5491 (N_5491,N_5383,N_5350);
xnor U5492 (N_5492,N_5397,N_5353);
xnor U5493 (N_5493,N_5345,N_5314);
and U5494 (N_5494,N_5335,N_5346);
and U5495 (N_5495,N_5363,N_5379);
xor U5496 (N_5496,N_5385,N_5338);
xnor U5497 (N_5497,N_5361,N_5371);
and U5498 (N_5498,N_5314,N_5394);
nor U5499 (N_5499,N_5374,N_5357);
or U5500 (N_5500,N_5450,N_5444);
xnor U5501 (N_5501,N_5422,N_5489);
and U5502 (N_5502,N_5423,N_5467);
nand U5503 (N_5503,N_5436,N_5468);
or U5504 (N_5504,N_5420,N_5427);
or U5505 (N_5505,N_5481,N_5484);
xor U5506 (N_5506,N_5456,N_5466);
nand U5507 (N_5507,N_5400,N_5414);
and U5508 (N_5508,N_5446,N_5453);
and U5509 (N_5509,N_5485,N_5417);
or U5510 (N_5510,N_5435,N_5447);
and U5511 (N_5511,N_5425,N_5432);
and U5512 (N_5512,N_5461,N_5402);
nand U5513 (N_5513,N_5454,N_5452);
nor U5514 (N_5514,N_5424,N_5410);
and U5515 (N_5515,N_5415,N_5445);
nor U5516 (N_5516,N_5463,N_5443);
nand U5517 (N_5517,N_5421,N_5449);
and U5518 (N_5518,N_5477,N_5403);
or U5519 (N_5519,N_5473,N_5470);
xnor U5520 (N_5520,N_5472,N_5458);
or U5521 (N_5521,N_5406,N_5442);
xor U5522 (N_5522,N_5469,N_5482);
nor U5523 (N_5523,N_5478,N_5437);
or U5524 (N_5524,N_5412,N_5475);
xnor U5525 (N_5525,N_5408,N_5440);
nand U5526 (N_5526,N_5495,N_5413);
and U5527 (N_5527,N_5457,N_5430);
xnor U5528 (N_5528,N_5494,N_5497);
and U5529 (N_5529,N_5431,N_5419);
xor U5530 (N_5530,N_5492,N_5439);
xnor U5531 (N_5531,N_5459,N_5438);
or U5532 (N_5532,N_5476,N_5483);
nor U5533 (N_5533,N_5471,N_5462);
nor U5534 (N_5534,N_5409,N_5499);
and U5535 (N_5535,N_5401,N_5460);
nand U5536 (N_5536,N_5487,N_5465);
or U5537 (N_5537,N_5486,N_5411);
nor U5538 (N_5538,N_5405,N_5429);
or U5539 (N_5539,N_5490,N_5479);
or U5540 (N_5540,N_5416,N_5493);
xnor U5541 (N_5541,N_5464,N_5488);
nand U5542 (N_5542,N_5451,N_5404);
nor U5543 (N_5543,N_5428,N_5480);
nor U5544 (N_5544,N_5441,N_5426);
or U5545 (N_5545,N_5474,N_5498);
xor U5546 (N_5546,N_5496,N_5448);
and U5547 (N_5547,N_5491,N_5455);
and U5548 (N_5548,N_5434,N_5407);
and U5549 (N_5549,N_5418,N_5433);
nor U5550 (N_5550,N_5420,N_5442);
xor U5551 (N_5551,N_5454,N_5479);
or U5552 (N_5552,N_5444,N_5457);
xnor U5553 (N_5553,N_5431,N_5496);
nor U5554 (N_5554,N_5498,N_5448);
xnor U5555 (N_5555,N_5436,N_5419);
and U5556 (N_5556,N_5486,N_5463);
and U5557 (N_5557,N_5450,N_5460);
xnor U5558 (N_5558,N_5411,N_5467);
nand U5559 (N_5559,N_5442,N_5405);
and U5560 (N_5560,N_5466,N_5492);
nor U5561 (N_5561,N_5491,N_5495);
and U5562 (N_5562,N_5417,N_5447);
xor U5563 (N_5563,N_5468,N_5425);
nor U5564 (N_5564,N_5470,N_5410);
xnor U5565 (N_5565,N_5475,N_5442);
xor U5566 (N_5566,N_5401,N_5471);
and U5567 (N_5567,N_5466,N_5477);
and U5568 (N_5568,N_5485,N_5461);
xor U5569 (N_5569,N_5496,N_5427);
xnor U5570 (N_5570,N_5447,N_5440);
nand U5571 (N_5571,N_5407,N_5453);
nor U5572 (N_5572,N_5467,N_5442);
and U5573 (N_5573,N_5435,N_5461);
and U5574 (N_5574,N_5487,N_5421);
or U5575 (N_5575,N_5494,N_5436);
nand U5576 (N_5576,N_5479,N_5463);
nand U5577 (N_5577,N_5408,N_5476);
nand U5578 (N_5578,N_5466,N_5404);
and U5579 (N_5579,N_5499,N_5427);
nor U5580 (N_5580,N_5478,N_5414);
or U5581 (N_5581,N_5490,N_5461);
or U5582 (N_5582,N_5408,N_5432);
nor U5583 (N_5583,N_5464,N_5424);
nor U5584 (N_5584,N_5489,N_5466);
and U5585 (N_5585,N_5488,N_5403);
or U5586 (N_5586,N_5403,N_5421);
nand U5587 (N_5587,N_5480,N_5474);
nand U5588 (N_5588,N_5486,N_5427);
or U5589 (N_5589,N_5480,N_5430);
nor U5590 (N_5590,N_5444,N_5435);
and U5591 (N_5591,N_5456,N_5440);
or U5592 (N_5592,N_5471,N_5433);
or U5593 (N_5593,N_5430,N_5489);
and U5594 (N_5594,N_5471,N_5436);
and U5595 (N_5595,N_5440,N_5419);
and U5596 (N_5596,N_5476,N_5445);
xnor U5597 (N_5597,N_5476,N_5423);
nor U5598 (N_5598,N_5457,N_5476);
nand U5599 (N_5599,N_5493,N_5442);
or U5600 (N_5600,N_5585,N_5574);
nand U5601 (N_5601,N_5568,N_5515);
or U5602 (N_5602,N_5598,N_5590);
xor U5603 (N_5603,N_5527,N_5524);
nor U5604 (N_5604,N_5554,N_5559);
nand U5605 (N_5605,N_5544,N_5528);
nor U5606 (N_5606,N_5511,N_5556);
xor U5607 (N_5607,N_5517,N_5580);
xor U5608 (N_5608,N_5567,N_5504);
and U5609 (N_5609,N_5513,N_5583);
and U5610 (N_5610,N_5566,N_5584);
nor U5611 (N_5611,N_5582,N_5549);
and U5612 (N_5612,N_5561,N_5514);
and U5613 (N_5613,N_5550,N_5599);
nand U5614 (N_5614,N_5505,N_5593);
nor U5615 (N_5615,N_5553,N_5597);
xor U5616 (N_5616,N_5538,N_5577);
nand U5617 (N_5617,N_5516,N_5520);
nor U5618 (N_5618,N_5589,N_5571);
xnor U5619 (N_5619,N_5572,N_5581);
nor U5620 (N_5620,N_5510,N_5573);
nor U5621 (N_5621,N_5588,N_5587);
and U5622 (N_5622,N_5547,N_5551);
or U5623 (N_5623,N_5569,N_5503);
nand U5624 (N_5624,N_5578,N_5500);
and U5625 (N_5625,N_5531,N_5579);
and U5626 (N_5626,N_5595,N_5521);
xor U5627 (N_5627,N_5540,N_5563);
and U5628 (N_5628,N_5560,N_5506);
nand U5629 (N_5629,N_5548,N_5507);
nor U5630 (N_5630,N_5552,N_5529);
or U5631 (N_5631,N_5539,N_5512);
and U5632 (N_5632,N_5523,N_5525);
nor U5633 (N_5633,N_5534,N_5558);
and U5634 (N_5634,N_5519,N_5502);
and U5635 (N_5635,N_5501,N_5576);
xor U5636 (N_5636,N_5526,N_5592);
nand U5637 (N_5637,N_5508,N_5537);
xnor U5638 (N_5638,N_5542,N_5545);
nand U5639 (N_5639,N_5541,N_5594);
nor U5640 (N_5640,N_5555,N_5536);
xor U5641 (N_5641,N_5596,N_5530);
and U5642 (N_5642,N_5575,N_5509);
or U5643 (N_5643,N_5586,N_5564);
or U5644 (N_5644,N_5562,N_5565);
xor U5645 (N_5645,N_5591,N_5543);
nor U5646 (N_5646,N_5570,N_5557);
nor U5647 (N_5647,N_5532,N_5546);
or U5648 (N_5648,N_5533,N_5522);
nand U5649 (N_5649,N_5535,N_5518);
nand U5650 (N_5650,N_5519,N_5500);
nor U5651 (N_5651,N_5508,N_5573);
and U5652 (N_5652,N_5563,N_5560);
or U5653 (N_5653,N_5541,N_5527);
xnor U5654 (N_5654,N_5545,N_5569);
or U5655 (N_5655,N_5538,N_5568);
xnor U5656 (N_5656,N_5534,N_5571);
nand U5657 (N_5657,N_5526,N_5528);
xor U5658 (N_5658,N_5597,N_5539);
xnor U5659 (N_5659,N_5598,N_5527);
or U5660 (N_5660,N_5540,N_5549);
and U5661 (N_5661,N_5554,N_5506);
nand U5662 (N_5662,N_5511,N_5536);
or U5663 (N_5663,N_5575,N_5546);
xor U5664 (N_5664,N_5567,N_5587);
xnor U5665 (N_5665,N_5559,N_5509);
xnor U5666 (N_5666,N_5557,N_5569);
nor U5667 (N_5667,N_5527,N_5510);
nor U5668 (N_5668,N_5502,N_5538);
or U5669 (N_5669,N_5598,N_5550);
xor U5670 (N_5670,N_5567,N_5565);
nand U5671 (N_5671,N_5555,N_5561);
nor U5672 (N_5672,N_5539,N_5581);
nor U5673 (N_5673,N_5598,N_5542);
xor U5674 (N_5674,N_5516,N_5566);
or U5675 (N_5675,N_5555,N_5562);
and U5676 (N_5676,N_5520,N_5568);
nor U5677 (N_5677,N_5595,N_5587);
nand U5678 (N_5678,N_5586,N_5546);
or U5679 (N_5679,N_5583,N_5580);
xor U5680 (N_5680,N_5587,N_5598);
nand U5681 (N_5681,N_5544,N_5565);
nor U5682 (N_5682,N_5587,N_5536);
nand U5683 (N_5683,N_5505,N_5501);
nor U5684 (N_5684,N_5560,N_5511);
nand U5685 (N_5685,N_5546,N_5509);
nor U5686 (N_5686,N_5536,N_5551);
and U5687 (N_5687,N_5565,N_5510);
xor U5688 (N_5688,N_5555,N_5589);
nor U5689 (N_5689,N_5500,N_5506);
nand U5690 (N_5690,N_5516,N_5559);
or U5691 (N_5691,N_5538,N_5517);
and U5692 (N_5692,N_5568,N_5523);
or U5693 (N_5693,N_5535,N_5591);
nor U5694 (N_5694,N_5563,N_5504);
xor U5695 (N_5695,N_5581,N_5523);
nand U5696 (N_5696,N_5592,N_5567);
xor U5697 (N_5697,N_5585,N_5513);
and U5698 (N_5698,N_5502,N_5589);
or U5699 (N_5699,N_5514,N_5546);
and U5700 (N_5700,N_5683,N_5691);
xor U5701 (N_5701,N_5639,N_5600);
and U5702 (N_5702,N_5671,N_5633);
nand U5703 (N_5703,N_5653,N_5609);
or U5704 (N_5704,N_5643,N_5635);
and U5705 (N_5705,N_5605,N_5672);
nand U5706 (N_5706,N_5625,N_5640);
xnor U5707 (N_5707,N_5622,N_5692);
and U5708 (N_5708,N_5620,N_5649);
nor U5709 (N_5709,N_5624,N_5694);
and U5710 (N_5710,N_5681,N_5665);
or U5711 (N_5711,N_5675,N_5606);
or U5712 (N_5712,N_5618,N_5646);
xor U5713 (N_5713,N_5603,N_5604);
or U5714 (N_5714,N_5697,N_5647);
nand U5715 (N_5715,N_5661,N_5686);
nor U5716 (N_5716,N_5641,N_5687);
nor U5717 (N_5717,N_5616,N_5684);
nand U5718 (N_5718,N_5601,N_5663);
and U5719 (N_5719,N_5614,N_5630);
xor U5720 (N_5720,N_5638,N_5612);
or U5721 (N_5721,N_5607,N_5696);
nand U5722 (N_5722,N_5657,N_5682);
nor U5723 (N_5723,N_5652,N_5654);
xor U5724 (N_5724,N_5636,N_5623);
or U5725 (N_5725,N_5674,N_5617);
nor U5726 (N_5726,N_5698,N_5673);
and U5727 (N_5727,N_5664,N_5676);
xor U5728 (N_5728,N_5666,N_5695);
xor U5729 (N_5729,N_5689,N_5637);
nand U5730 (N_5730,N_5608,N_5677);
nand U5731 (N_5731,N_5644,N_5650);
nor U5732 (N_5732,N_5628,N_5659);
and U5733 (N_5733,N_5667,N_5621);
xnor U5734 (N_5734,N_5627,N_5626);
nor U5735 (N_5735,N_5648,N_5662);
nand U5736 (N_5736,N_5655,N_5693);
nor U5737 (N_5737,N_5615,N_5619);
nand U5738 (N_5738,N_5632,N_5634);
nand U5739 (N_5739,N_5631,N_5688);
and U5740 (N_5740,N_5610,N_5651);
or U5741 (N_5741,N_5660,N_5668);
xnor U5742 (N_5742,N_5645,N_5611);
nor U5743 (N_5743,N_5629,N_5658);
and U5744 (N_5744,N_5613,N_5679);
or U5745 (N_5745,N_5678,N_5690);
xor U5746 (N_5746,N_5670,N_5602);
or U5747 (N_5747,N_5669,N_5685);
and U5748 (N_5748,N_5656,N_5642);
nor U5749 (N_5749,N_5699,N_5680);
xnor U5750 (N_5750,N_5673,N_5661);
nand U5751 (N_5751,N_5661,N_5611);
or U5752 (N_5752,N_5629,N_5644);
or U5753 (N_5753,N_5605,N_5607);
and U5754 (N_5754,N_5642,N_5685);
nand U5755 (N_5755,N_5677,N_5665);
or U5756 (N_5756,N_5651,N_5611);
nor U5757 (N_5757,N_5682,N_5600);
and U5758 (N_5758,N_5686,N_5660);
nand U5759 (N_5759,N_5636,N_5681);
or U5760 (N_5760,N_5675,N_5658);
or U5761 (N_5761,N_5662,N_5604);
xnor U5762 (N_5762,N_5619,N_5616);
or U5763 (N_5763,N_5614,N_5664);
nor U5764 (N_5764,N_5603,N_5613);
and U5765 (N_5765,N_5626,N_5606);
and U5766 (N_5766,N_5625,N_5611);
nor U5767 (N_5767,N_5620,N_5664);
nor U5768 (N_5768,N_5662,N_5675);
and U5769 (N_5769,N_5639,N_5693);
and U5770 (N_5770,N_5633,N_5694);
or U5771 (N_5771,N_5602,N_5617);
nor U5772 (N_5772,N_5673,N_5644);
xor U5773 (N_5773,N_5693,N_5619);
nand U5774 (N_5774,N_5647,N_5673);
xnor U5775 (N_5775,N_5673,N_5643);
and U5776 (N_5776,N_5669,N_5620);
or U5777 (N_5777,N_5641,N_5610);
and U5778 (N_5778,N_5687,N_5696);
and U5779 (N_5779,N_5653,N_5680);
xor U5780 (N_5780,N_5622,N_5650);
or U5781 (N_5781,N_5670,N_5618);
nand U5782 (N_5782,N_5669,N_5652);
or U5783 (N_5783,N_5634,N_5625);
or U5784 (N_5784,N_5640,N_5670);
and U5785 (N_5785,N_5641,N_5670);
and U5786 (N_5786,N_5695,N_5603);
nand U5787 (N_5787,N_5677,N_5615);
xnor U5788 (N_5788,N_5660,N_5626);
nor U5789 (N_5789,N_5694,N_5644);
xor U5790 (N_5790,N_5607,N_5677);
nor U5791 (N_5791,N_5651,N_5675);
xnor U5792 (N_5792,N_5690,N_5626);
nand U5793 (N_5793,N_5646,N_5622);
or U5794 (N_5794,N_5655,N_5663);
or U5795 (N_5795,N_5634,N_5608);
or U5796 (N_5796,N_5697,N_5671);
nor U5797 (N_5797,N_5660,N_5655);
or U5798 (N_5798,N_5698,N_5685);
nand U5799 (N_5799,N_5618,N_5611);
and U5800 (N_5800,N_5750,N_5745);
and U5801 (N_5801,N_5719,N_5781);
nand U5802 (N_5802,N_5712,N_5732);
nor U5803 (N_5803,N_5763,N_5785);
and U5804 (N_5804,N_5722,N_5746);
xnor U5805 (N_5805,N_5773,N_5713);
nor U5806 (N_5806,N_5771,N_5721);
nor U5807 (N_5807,N_5736,N_5783);
and U5808 (N_5808,N_5729,N_5747);
xnor U5809 (N_5809,N_5707,N_5727);
and U5810 (N_5810,N_5751,N_5743);
xor U5811 (N_5811,N_5738,N_5795);
or U5812 (N_5812,N_5733,N_5759);
nor U5813 (N_5813,N_5708,N_5702);
xor U5814 (N_5814,N_5737,N_5764);
xnor U5815 (N_5815,N_5770,N_5797);
nand U5816 (N_5816,N_5789,N_5793);
or U5817 (N_5817,N_5752,N_5776);
or U5818 (N_5818,N_5774,N_5724);
nor U5819 (N_5819,N_5756,N_5742);
nand U5820 (N_5820,N_5777,N_5768);
nand U5821 (N_5821,N_5786,N_5758);
nand U5822 (N_5822,N_5717,N_5739);
and U5823 (N_5823,N_5705,N_5772);
and U5824 (N_5824,N_5779,N_5778);
and U5825 (N_5825,N_5725,N_5715);
xnor U5826 (N_5826,N_5798,N_5788);
and U5827 (N_5827,N_5731,N_5767);
and U5828 (N_5828,N_5766,N_5741);
nand U5829 (N_5829,N_5792,N_5799);
or U5830 (N_5830,N_5734,N_5706);
nor U5831 (N_5831,N_5749,N_5761);
xor U5832 (N_5832,N_5726,N_5791);
or U5833 (N_5833,N_5790,N_5765);
xor U5834 (N_5834,N_5744,N_5775);
xnor U5835 (N_5835,N_5704,N_5730);
nor U5836 (N_5836,N_5760,N_5794);
or U5837 (N_5837,N_5740,N_5769);
or U5838 (N_5838,N_5710,N_5784);
xnor U5839 (N_5839,N_5757,N_5753);
xnor U5840 (N_5840,N_5782,N_5716);
nor U5841 (N_5841,N_5700,N_5735);
nor U5842 (N_5842,N_5755,N_5701);
or U5843 (N_5843,N_5720,N_5703);
nor U5844 (N_5844,N_5787,N_5718);
and U5845 (N_5845,N_5796,N_5762);
and U5846 (N_5846,N_5780,N_5754);
and U5847 (N_5847,N_5714,N_5748);
and U5848 (N_5848,N_5728,N_5709);
nor U5849 (N_5849,N_5711,N_5723);
or U5850 (N_5850,N_5741,N_5775);
and U5851 (N_5851,N_5740,N_5756);
and U5852 (N_5852,N_5738,N_5781);
and U5853 (N_5853,N_5712,N_5747);
xor U5854 (N_5854,N_5750,N_5785);
or U5855 (N_5855,N_5726,N_5772);
and U5856 (N_5856,N_5752,N_5757);
and U5857 (N_5857,N_5750,N_5777);
nand U5858 (N_5858,N_5788,N_5780);
xnor U5859 (N_5859,N_5759,N_5742);
or U5860 (N_5860,N_5767,N_5710);
nor U5861 (N_5861,N_5757,N_5778);
xor U5862 (N_5862,N_5738,N_5784);
xnor U5863 (N_5863,N_5786,N_5793);
nor U5864 (N_5864,N_5711,N_5767);
xor U5865 (N_5865,N_5734,N_5710);
and U5866 (N_5866,N_5765,N_5774);
nor U5867 (N_5867,N_5738,N_5791);
nor U5868 (N_5868,N_5764,N_5755);
nor U5869 (N_5869,N_5710,N_5757);
nand U5870 (N_5870,N_5744,N_5726);
xor U5871 (N_5871,N_5749,N_5797);
xnor U5872 (N_5872,N_5770,N_5761);
and U5873 (N_5873,N_5734,N_5720);
and U5874 (N_5874,N_5707,N_5703);
and U5875 (N_5875,N_5791,N_5713);
and U5876 (N_5876,N_5736,N_5768);
and U5877 (N_5877,N_5789,N_5764);
or U5878 (N_5878,N_5785,N_5719);
xor U5879 (N_5879,N_5722,N_5719);
nor U5880 (N_5880,N_5773,N_5756);
or U5881 (N_5881,N_5775,N_5719);
and U5882 (N_5882,N_5748,N_5722);
or U5883 (N_5883,N_5726,N_5788);
nand U5884 (N_5884,N_5767,N_5706);
and U5885 (N_5885,N_5725,N_5783);
xnor U5886 (N_5886,N_5700,N_5738);
xor U5887 (N_5887,N_5716,N_5787);
nor U5888 (N_5888,N_5795,N_5759);
xnor U5889 (N_5889,N_5726,N_5719);
or U5890 (N_5890,N_5701,N_5763);
nand U5891 (N_5891,N_5757,N_5727);
xor U5892 (N_5892,N_5714,N_5736);
nor U5893 (N_5893,N_5762,N_5770);
or U5894 (N_5894,N_5793,N_5799);
and U5895 (N_5895,N_5714,N_5738);
and U5896 (N_5896,N_5791,N_5717);
nand U5897 (N_5897,N_5774,N_5763);
and U5898 (N_5898,N_5783,N_5740);
xor U5899 (N_5899,N_5742,N_5703);
xor U5900 (N_5900,N_5882,N_5894);
and U5901 (N_5901,N_5871,N_5869);
xor U5902 (N_5902,N_5830,N_5877);
and U5903 (N_5903,N_5856,N_5893);
or U5904 (N_5904,N_5885,N_5810);
xor U5905 (N_5905,N_5870,N_5861);
or U5906 (N_5906,N_5897,N_5864);
nand U5907 (N_5907,N_5868,N_5878);
or U5908 (N_5908,N_5883,N_5895);
or U5909 (N_5909,N_5823,N_5816);
nor U5910 (N_5910,N_5881,N_5844);
or U5911 (N_5911,N_5814,N_5845);
nor U5912 (N_5912,N_5804,N_5889);
or U5913 (N_5913,N_5824,N_5859);
xor U5914 (N_5914,N_5840,N_5827);
nand U5915 (N_5915,N_5819,N_5835);
xnor U5916 (N_5916,N_5862,N_5821);
xnor U5917 (N_5917,N_5801,N_5880);
xor U5918 (N_5918,N_5837,N_5863);
and U5919 (N_5919,N_5805,N_5826);
or U5920 (N_5920,N_5806,N_5839);
nor U5921 (N_5921,N_5833,N_5803);
and U5922 (N_5922,N_5831,N_5812);
nand U5923 (N_5923,N_5853,N_5884);
or U5924 (N_5924,N_5836,N_5843);
xnor U5925 (N_5925,N_5825,N_5820);
nand U5926 (N_5926,N_5842,N_5874);
and U5927 (N_5927,N_5809,N_5832);
nand U5928 (N_5928,N_5811,N_5815);
nor U5929 (N_5929,N_5800,N_5898);
and U5930 (N_5930,N_5860,N_5857);
nor U5931 (N_5931,N_5852,N_5802);
and U5932 (N_5932,N_5866,N_5838);
xnor U5933 (N_5933,N_5886,N_5847);
nand U5934 (N_5934,N_5890,N_5873);
or U5935 (N_5935,N_5896,N_5879);
xnor U5936 (N_5936,N_5846,N_5841);
xnor U5937 (N_5937,N_5848,N_5822);
or U5938 (N_5938,N_5899,N_5865);
nand U5939 (N_5939,N_5818,N_5813);
and U5940 (N_5940,N_5858,N_5829);
and U5941 (N_5941,N_5872,N_5888);
nor U5942 (N_5942,N_5855,N_5850);
nand U5943 (N_5943,N_5834,N_5851);
or U5944 (N_5944,N_5828,N_5807);
nand U5945 (N_5945,N_5892,N_5817);
and U5946 (N_5946,N_5876,N_5891);
nor U5947 (N_5947,N_5849,N_5854);
or U5948 (N_5948,N_5875,N_5867);
xor U5949 (N_5949,N_5887,N_5808);
nor U5950 (N_5950,N_5857,N_5879);
or U5951 (N_5951,N_5832,N_5876);
nand U5952 (N_5952,N_5853,N_5894);
and U5953 (N_5953,N_5833,N_5809);
and U5954 (N_5954,N_5873,N_5834);
and U5955 (N_5955,N_5807,N_5855);
xor U5956 (N_5956,N_5870,N_5884);
nor U5957 (N_5957,N_5879,N_5861);
nand U5958 (N_5958,N_5890,N_5877);
nand U5959 (N_5959,N_5838,N_5884);
xor U5960 (N_5960,N_5832,N_5824);
nand U5961 (N_5961,N_5892,N_5853);
nor U5962 (N_5962,N_5891,N_5872);
nor U5963 (N_5963,N_5851,N_5852);
and U5964 (N_5964,N_5881,N_5821);
nand U5965 (N_5965,N_5841,N_5818);
nand U5966 (N_5966,N_5881,N_5891);
xor U5967 (N_5967,N_5802,N_5890);
nand U5968 (N_5968,N_5854,N_5839);
and U5969 (N_5969,N_5868,N_5844);
nand U5970 (N_5970,N_5816,N_5869);
nand U5971 (N_5971,N_5859,N_5844);
and U5972 (N_5972,N_5825,N_5886);
and U5973 (N_5973,N_5871,N_5874);
nand U5974 (N_5974,N_5881,N_5875);
xnor U5975 (N_5975,N_5847,N_5816);
and U5976 (N_5976,N_5849,N_5846);
nand U5977 (N_5977,N_5826,N_5827);
nand U5978 (N_5978,N_5860,N_5816);
or U5979 (N_5979,N_5828,N_5818);
and U5980 (N_5980,N_5843,N_5859);
and U5981 (N_5981,N_5817,N_5802);
xor U5982 (N_5982,N_5894,N_5829);
nor U5983 (N_5983,N_5883,N_5868);
nand U5984 (N_5984,N_5872,N_5803);
and U5985 (N_5985,N_5863,N_5871);
xor U5986 (N_5986,N_5873,N_5823);
xor U5987 (N_5987,N_5889,N_5857);
nor U5988 (N_5988,N_5825,N_5800);
and U5989 (N_5989,N_5818,N_5805);
nor U5990 (N_5990,N_5866,N_5822);
nand U5991 (N_5991,N_5882,N_5864);
and U5992 (N_5992,N_5856,N_5811);
nor U5993 (N_5993,N_5834,N_5835);
xnor U5994 (N_5994,N_5891,N_5805);
xnor U5995 (N_5995,N_5821,N_5825);
or U5996 (N_5996,N_5834,N_5896);
and U5997 (N_5997,N_5819,N_5870);
and U5998 (N_5998,N_5827,N_5866);
or U5999 (N_5999,N_5884,N_5827);
nor U6000 (N_6000,N_5979,N_5910);
and U6001 (N_6001,N_5926,N_5901);
xnor U6002 (N_6002,N_5900,N_5902);
or U6003 (N_6003,N_5909,N_5952);
nor U6004 (N_6004,N_5996,N_5954);
nand U6005 (N_6005,N_5949,N_5940);
nand U6006 (N_6006,N_5946,N_5989);
or U6007 (N_6007,N_5939,N_5933);
and U6008 (N_6008,N_5918,N_5987);
nor U6009 (N_6009,N_5923,N_5994);
nand U6010 (N_6010,N_5990,N_5958);
nor U6011 (N_6011,N_5930,N_5924);
xor U6012 (N_6012,N_5961,N_5932);
nand U6013 (N_6013,N_5984,N_5972);
xnor U6014 (N_6014,N_5938,N_5986);
nand U6015 (N_6015,N_5964,N_5966);
or U6016 (N_6016,N_5908,N_5929);
or U6017 (N_6017,N_5965,N_5967);
or U6018 (N_6018,N_5983,N_5981);
nor U6019 (N_6019,N_5985,N_5944);
nor U6020 (N_6020,N_5971,N_5945);
nand U6021 (N_6021,N_5947,N_5974);
nand U6022 (N_6022,N_5980,N_5913);
and U6023 (N_6023,N_5912,N_5917);
and U6024 (N_6024,N_5935,N_5920);
xnor U6025 (N_6025,N_5937,N_5904);
nor U6026 (N_6026,N_5905,N_5992);
xor U6027 (N_6027,N_5915,N_5960);
and U6028 (N_6028,N_5953,N_5993);
or U6029 (N_6029,N_5903,N_5936);
and U6030 (N_6030,N_5982,N_5907);
and U6031 (N_6031,N_5977,N_5957);
or U6032 (N_6032,N_5956,N_5997);
and U6033 (N_6033,N_5928,N_5925);
xor U6034 (N_6034,N_5931,N_5973);
xnor U6035 (N_6035,N_5919,N_5955);
nand U6036 (N_6036,N_5969,N_5941);
nand U6037 (N_6037,N_5975,N_5978);
or U6038 (N_6038,N_5976,N_5991);
xnor U6039 (N_6039,N_5943,N_5914);
or U6040 (N_6040,N_5962,N_5959);
xnor U6041 (N_6041,N_5922,N_5942);
nand U6042 (N_6042,N_5999,N_5998);
and U6043 (N_6043,N_5927,N_5934);
nor U6044 (N_6044,N_5963,N_5906);
nand U6045 (N_6045,N_5921,N_5995);
and U6046 (N_6046,N_5911,N_5968);
or U6047 (N_6047,N_5916,N_5988);
nor U6048 (N_6048,N_5970,N_5948);
xnor U6049 (N_6049,N_5951,N_5950);
nor U6050 (N_6050,N_5938,N_5974);
nor U6051 (N_6051,N_5979,N_5930);
nor U6052 (N_6052,N_5908,N_5950);
or U6053 (N_6053,N_5937,N_5981);
or U6054 (N_6054,N_5986,N_5989);
nand U6055 (N_6055,N_5978,N_5907);
nor U6056 (N_6056,N_5935,N_5945);
or U6057 (N_6057,N_5962,N_5921);
xor U6058 (N_6058,N_5906,N_5900);
and U6059 (N_6059,N_5949,N_5984);
xor U6060 (N_6060,N_5961,N_5995);
xor U6061 (N_6061,N_5986,N_5950);
nand U6062 (N_6062,N_5989,N_5903);
xor U6063 (N_6063,N_5903,N_5985);
nor U6064 (N_6064,N_5973,N_5938);
nand U6065 (N_6065,N_5933,N_5944);
or U6066 (N_6066,N_5985,N_5922);
nor U6067 (N_6067,N_5912,N_5945);
and U6068 (N_6068,N_5960,N_5926);
or U6069 (N_6069,N_5938,N_5979);
xor U6070 (N_6070,N_5988,N_5953);
nor U6071 (N_6071,N_5976,N_5908);
xor U6072 (N_6072,N_5949,N_5928);
nand U6073 (N_6073,N_5977,N_5930);
nor U6074 (N_6074,N_5935,N_5984);
and U6075 (N_6075,N_5954,N_5952);
or U6076 (N_6076,N_5984,N_5977);
xor U6077 (N_6077,N_5963,N_5958);
nor U6078 (N_6078,N_5905,N_5925);
nor U6079 (N_6079,N_5931,N_5996);
or U6080 (N_6080,N_5940,N_5996);
or U6081 (N_6081,N_5958,N_5933);
nand U6082 (N_6082,N_5959,N_5968);
nor U6083 (N_6083,N_5971,N_5921);
xnor U6084 (N_6084,N_5929,N_5904);
and U6085 (N_6085,N_5903,N_5928);
nand U6086 (N_6086,N_5986,N_5908);
and U6087 (N_6087,N_5986,N_5970);
xnor U6088 (N_6088,N_5943,N_5951);
nor U6089 (N_6089,N_5955,N_5938);
xor U6090 (N_6090,N_5966,N_5982);
xor U6091 (N_6091,N_5950,N_5970);
and U6092 (N_6092,N_5918,N_5928);
or U6093 (N_6093,N_5944,N_5963);
or U6094 (N_6094,N_5925,N_5989);
and U6095 (N_6095,N_5942,N_5930);
nand U6096 (N_6096,N_5995,N_5981);
xor U6097 (N_6097,N_5916,N_5917);
and U6098 (N_6098,N_5935,N_5934);
xnor U6099 (N_6099,N_5911,N_5967);
xnor U6100 (N_6100,N_6043,N_6082);
or U6101 (N_6101,N_6031,N_6090);
nand U6102 (N_6102,N_6051,N_6064);
and U6103 (N_6103,N_6045,N_6055);
or U6104 (N_6104,N_6089,N_6060);
xor U6105 (N_6105,N_6014,N_6079);
xor U6106 (N_6106,N_6024,N_6067);
or U6107 (N_6107,N_6026,N_6019);
xor U6108 (N_6108,N_6007,N_6080);
and U6109 (N_6109,N_6041,N_6081);
nand U6110 (N_6110,N_6094,N_6027);
or U6111 (N_6111,N_6099,N_6063);
or U6112 (N_6112,N_6002,N_6049);
xnor U6113 (N_6113,N_6038,N_6058);
nand U6114 (N_6114,N_6071,N_6098);
and U6115 (N_6115,N_6036,N_6062);
or U6116 (N_6116,N_6065,N_6010);
and U6117 (N_6117,N_6069,N_6011);
or U6118 (N_6118,N_6075,N_6048);
or U6119 (N_6119,N_6066,N_6013);
or U6120 (N_6120,N_6018,N_6050);
and U6121 (N_6121,N_6088,N_6005);
nor U6122 (N_6122,N_6040,N_6070);
nor U6123 (N_6123,N_6061,N_6093);
nand U6124 (N_6124,N_6003,N_6012);
and U6125 (N_6125,N_6087,N_6015);
and U6126 (N_6126,N_6095,N_6053);
nand U6127 (N_6127,N_6035,N_6085);
nor U6128 (N_6128,N_6008,N_6059);
xnor U6129 (N_6129,N_6020,N_6009);
nor U6130 (N_6130,N_6023,N_6032);
and U6131 (N_6131,N_6073,N_6047);
xnor U6132 (N_6132,N_6037,N_6016);
or U6133 (N_6133,N_6004,N_6052);
and U6134 (N_6134,N_6046,N_6030);
or U6135 (N_6135,N_6039,N_6074);
or U6136 (N_6136,N_6097,N_6056);
nor U6137 (N_6137,N_6017,N_6084);
and U6138 (N_6138,N_6091,N_6042);
nand U6139 (N_6139,N_6000,N_6033);
nor U6140 (N_6140,N_6078,N_6001);
xor U6141 (N_6141,N_6068,N_6083);
nand U6142 (N_6142,N_6034,N_6086);
xnor U6143 (N_6143,N_6057,N_6077);
xor U6144 (N_6144,N_6072,N_6029);
xor U6145 (N_6145,N_6021,N_6025);
and U6146 (N_6146,N_6006,N_6092);
nand U6147 (N_6147,N_6096,N_6022);
nand U6148 (N_6148,N_6076,N_6044);
nor U6149 (N_6149,N_6054,N_6028);
nor U6150 (N_6150,N_6072,N_6061);
nor U6151 (N_6151,N_6007,N_6078);
or U6152 (N_6152,N_6027,N_6032);
and U6153 (N_6153,N_6092,N_6029);
or U6154 (N_6154,N_6094,N_6007);
xor U6155 (N_6155,N_6044,N_6053);
nand U6156 (N_6156,N_6035,N_6022);
and U6157 (N_6157,N_6083,N_6007);
or U6158 (N_6158,N_6011,N_6035);
or U6159 (N_6159,N_6098,N_6041);
or U6160 (N_6160,N_6064,N_6095);
xor U6161 (N_6161,N_6031,N_6054);
nand U6162 (N_6162,N_6027,N_6054);
xor U6163 (N_6163,N_6000,N_6091);
and U6164 (N_6164,N_6073,N_6084);
or U6165 (N_6165,N_6032,N_6052);
or U6166 (N_6166,N_6069,N_6084);
nor U6167 (N_6167,N_6023,N_6020);
and U6168 (N_6168,N_6019,N_6052);
xor U6169 (N_6169,N_6041,N_6066);
xnor U6170 (N_6170,N_6059,N_6019);
xnor U6171 (N_6171,N_6014,N_6023);
nand U6172 (N_6172,N_6046,N_6053);
nor U6173 (N_6173,N_6037,N_6095);
or U6174 (N_6174,N_6055,N_6058);
xor U6175 (N_6175,N_6047,N_6045);
and U6176 (N_6176,N_6039,N_6048);
nor U6177 (N_6177,N_6019,N_6079);
and U6178 (N_6178,N_6073,N_6040);
xor U6179 (N_6179,N_6036,N_6068);
and U6180 (N_6180,N_6001,N_6058);
and U6181 (N_6181,N_6011,N_6034);
or U6182 (N_6182,N_6079,N_6020);
nor U6183 (N_6183,N_6034,N_6009);
or U6184 (N_6184,N_6091,N_6053);
and U6185 (N_6185,N_6008,N_6067);
and U6186 (N_6186,N_6039,N_6032);
nand U6187 (N_6187,N_6072,N_6046);
nor U6188 (N_6188,N_6022,N_6005);
nor U6189 (N_6189,N_6089,N_6059);
nor U6190 (N_6190,N_6001,N_6003);
and U6191 (N_6191,N_6071,N_6003);
and U6192 (N_6192,N_6016,N_6091);
nor U6193 (N_6193,N_6094,N_6083);
nand U6194 (N_6194,N_6001,N_6013);
or U6195 (N_6195,N_6067,N_6055);
xor U6196 (N_6196,N_6040,N_6057);
nand U6197 (N_6197,N_6024,N_6026);
nand U6198 (N_6198,N_6047,N_6054);
or U6199 (N_6199,N_6051,N_6091);
or U6200 (N_6200,N_6142,N_6111);
nand U6201 (N_6201,N_6101,N_6176);
nand U6202 (N_6202,N_6149,N_6190);
nor U6203 (N_6203,N_6148,N_6146);
xnor U6204 (N_6204,N_6186,N_6113);
nand U6205 (N_6205,N_6127,N_6136);
nand U6206 (N_6206,N_6118,N_6126);
and U6207 (N_6207,N_6189,N_6117);
nand U6208 (N_6208,N_6191,N_6160);
nand U6209 (N_6209,N_6165,N_6158);
xor U6210 (N_6210,N_6133,N_6131);
and U6211 (N_6211,N_6192,N_6153);
and U6212 (N_6212,N_6132,N_6102);
xor U6213 (N_6213,N_6152,N_6174);
nor U6214 (N_6214,N_6139,N_6169);
nand U6215 (N_6215,N_6163,N_6172);
nor U6216 (N_6216,N_6107,N_6156);
nor U6217 (N_6217,N_6123,N_6137);
nand U6218 (N_6218,N_6144,N_6100);
nand U6219 (N_6219,N_6180,N_6150);
and U6220 (N_6220,N_6129,N_6183);
xnor U6221 (N_6221,N_6106,N_6162);
or U6222 (N_6222,N_6110,N_6143);
nand U6223 (N_6223,N_6159,N_6104);
or U6224 (N_6224,N_6121,N_6194);
or U6225 (N_6225,N_6181,N_6140);
xnor U6226 (N_6226,N_6125,N_6161);
or U6227 (N_6227,N_6119,N_6134);
nor U6228 (N_6228,N_6173,N_6167);
and U6229 (N_6229,N_6195,N_6154);
nor U6230 (N_6230,N_6155,N_6177);
and U6231 (N_6231,N_6108,N_6138);
and U6232 (N_6232,N_6145,N_6151);
nand U6233 (N_6233,N_6179,N_6157);
nor U6234 (N_6234,N_6112,N_6135);
or U6235 (N_6235,N_6128,N_6182);
nand U6236 (N_6236,N_6187,N_6197);
xor U6237 (N_6237,N_6166,N_6116);
nand U6238 (N_6238,N_6170,N_6105);
and U6239 (N_6239,N_6115,N_6175);
nand U6240 (N_6240,N_6196,N_6168);
xnor U6241 (N_6241,N_6130,N_6185);
xor U6242 (N_6242,N_6171,N_6193);
or U6243 (N_6243,N_6199,N_6164);
nand U6244 (N_6244,N_6114,N_6120);
xor U6245 (N_6245,N_6109,N_6178);
xor U6246 (N_6246,N_6141,N_6124);
nand U6247 (N_6247,N_6147,N_6103);
nor U6248 (N_6248,N_6122,N_6198);
nand U6249 (N_6249,N_6188,N_6184);
xor U6250 (N_6250,N_6119,N_6171);
nand U6251 (N_6251,N_6103,N_6161);
xnor U6252 (N_6252,N_6130,N_6100);
nand U6253 (N_6253,N_6135,N_6136);
xnor U6254 (N_6254,N_6107,N_6180);
nor U6255 (N_6255,N_6169,N_6162);
nand U6256 (N_6256,N_6167,N_6157);
or U6257 (N_6257,N_6118,N_6135);
and U6258 (N_6258,N_6120,N_6142);
nor U6259 (N_6259,N_6131,N_6146);
nand U6260 (N_6260,N_6166,N_6126);
or U6261 (N_6261,N_6163,N_6187);
and U6262 (N_6262,N_6162,N_6195);
and U6263 (N_6263,N_6182,N_6116);
or U6264 (N_6264,N_6133,N_6100);
xor U6265 (N_6265,N_6188,N_6116);
nand U6266 (N_6266,N_6123,N_6101);
and U6267 (N_6267,N_6128,N_6111);
and U6268 (N_6268,N_6140,N_6180);
and U6269 (N_6269,N_6102,N_6173);
xnor U6270 (N_6270,N_6177,N_6148);
nor U6271 (N_6271,N_6129,N_6109);
nor U6272 (N_6272,N_6113,N_6106);
nand U6273 (N_6273,N_6179,N_6194);
or U6274 (N_6274,N_6107,N_6144);
or U6275 (N_6275,N_6197,N_6166);
xnor U6276 (N_6276,N_6154,N_6100);
nand U6277 (N_6277,N_6164,N_6156);
and U6278 (N_6278,N_6165,N_6140);
or U6279 (N_6279,N_6119,N_6172);
and U6280 (N_6280,N_6132,N_6136);
and U6281 (N_6281,N_6169,N_6195);
and U6282 (N_6282,N_6158,N_6109);
or U6283 (N_6283,N_6148,N_6120);
nor U6284 (N_6284,N_6196,N_6140);
nand U6285 (N_6285,N_6121,N_6186);
xor U6286 (N_6286,N_6176,N_6190);
xnor U6287 (N_6287,N_6102,N_6183);
or U6288 (N_6288,N_6107,N_6193);
nor U6289 (N_6289,N_6142,N_6106);
and U6290 (N_6290,N_6114,N_6124);
nand U6291 (N_6291,N_6194,N_6141);
nand U6292 (N_6292,N_6100,N_6157);
nor U6293 (N_6293,N_6165,N_6123);
and U6294 (N_6294,N_6125,N_6152);
nand U6295 (N_6295,N_6116,N_6142);
xnor U6296 (N_6296,N_6118,N_6146);
nand U6297 (N_6297,N_6146,N_6143);
or U6298 (N_6298,N_6108,N_6188);
and U6299 (N_6299,N_6180,N_6176);
or U6300 (N_6300,N_6235,N_6206);
xnor U6301 (N_6301,N_6213,N_6296);
nor U6302 (N_6302,N_6286,N_6249);
and U6303 (N_6303,N_6278,N_6259);
nand U6304 (N_6304,N_6240,N_6284);
nor U6305 (N_6305,N_6254,N_6255);
nand U6306 (N_6306,N_6241,N_6247);
nand U6307 (N_6307,N_6211,N_6214);
xor U6308 (N_6308,N_6280,N_6230);
nor U6309 (N_6309,N_6208,N_6225);
nor U6310 (N_6310,N_6231,N_6262);
xor U6311 (N_6311,N_6258,N_6229);
nor U6312 (N_6312,N_6282,N_6222);
nor U6313 (N_6313,N_6243,N_6217);
or U6314 (N_6314,N_6242,N_6268);
or U6315 (N_6315,N_6277,N_6244);
nand U6316 (N_6316,N_6294,N_6276);
nor U6317 (N_6317,N_6234,N_6273);
nor U6318 (N_6318,N_6203,N_6266);
nor U6319 (N_6319,N_6232,N_6238);
or U6320 (N_6320,N_6201,N_6223);
xor U6321 (N_6321,N_6256,N_6248);
and U6322 (N_6322,N_6272,N_6263);
nor U6323 (N_6323,N_6252,N_6290);
or U6324 (N_6324,N_6253,N_6228);
xor U6325 (N_6325,N_6200,N_6215);
nor U6326 (N_6326,N_6226,N_6298);
nor U6327 (N_6327,N_6218,N_6246);
xor U6328 (N_6328,N_6251,N_6270);
and U6329 (N_6329,N_6289,N_6267);
and U6330 (N_6330,N_6239,N_6293);
nor U6331 (N_6331,N_6269,N_6221);
and U6332 (N_6332,N_6204,N_6292);
nor U6333 (N_6333,N_6224,N_6260);
nor U6334 (N_6334,N_6219,N_6245);
xor U6335 (N_6335,N_6210,N_6205);
nor U6336 (N_6336,N_6236,N_6275);
xor U6337 (N_6337,N_6207,N_6237);
nor U6338 (N_6338,N_6216,N_6265);
and U6339 (N_6339,N_6250,N_6288);
nand U6340 (N_6340,N_6297,N_6257);
nand U6341 (N_6341,N_6212,N_6287);
nand U6342 (N_6342,N_6281,N_6227);
nor U6343 (N_6343,N_6283,N_6271);
xnor U6344 (N_6344,N_6295,N_6291);
nand U6345 (N_6345,N_6274,N_6233);
or U6346 (N_6346,N_6220,N_6202);
xor U6347 (N_6347,N_6299,N_6261);
xnor U6348 (N_6348,N_6279,N_6209);
xnor U6349 (N_6349,N_6285,N_6264);
nand U6350 (N_6350,N_6239,N_6257);
nor U6351 (N_6351,N_6242,N_6287);
xnor U6352 (N_6352,N_6241,N_6259);
nor U6353 (N_6353,N_6247,N_6204);
or U6354 (N_6354,N_6222,N_6276);
nor U6355 (N_6355,N_6281,N_6205);
nand U6356 (N_6356,N_6206,N_6273);
xnor U6357 (N_6357,N_6270,N_6211);
nor U6358 (N_6358,N_6290,N_6231);
nand U6359 (N_6359,N_6219,N_6218);
nor U6360 (N_6360,N_6265,N_6213);
xnor U6361 (N_6361,N_6297,N_6242);
or U6362 (N_6362,N_6201,N_6275);
nor U6363 (N_6363,N_6207,N_6254);
nand U6364 (N_6364,N_6238,N_6247);
or U6365 (N_6365,N_6257,N_6270);
nand U6366 (N_6366,N_6202,N_6283);
xnor U6367 (N_6367,N_6202,N_6249);
and U6368 (N_6368,N_6273,N_6210);
and U6369 (N_6369,N_6217,N_6230);
nand U6370 (N_6370,N_6230,N_6226);
nor U6371 (N_6371,N_6235,N_6220);
nand U6372 (N_6372,N_6288,N_6280);
xnor U6373 (N_6373,N_6292,N_6252);
and U6374 (N_6374,N_6297,N_6246);
and U6375 (N_6375,N_6257,N_6219);
nor U6376 (N_6376,N_6281,N_6222);
nor U6377 (N_6377,N_6241,N_6200);
nand U6378 (N_6378,N_6256,N_6228);
nand U6379 (N_6379,N_6275,N_6262);
nor U6380 (N_6380,N_6227,N_6201);
xor U6381 (N_6381,N_6205,N_6213);
xor U6382 (N_6382,N_6254,N_6217);
nand U6383 (N_6383,N_6221,N_6276);
nand U6384 (N_6384,N_6289,N_6237);
xor U6385 (N_6385,N_6234,N_6291);
nor U6386 (N_6386,N_6241,N_6248);
or U6387 (N_6387,N_6282,N_6205);
nor U6388 (N_6388,N_6251,N_6224);
nor U6389 (N_6389,N_6279,N_6296);
xor U6390 (N_6390,N_6225,N_6226);
or U6391 (N_6391,N_6214,N_6241);
and U6392 (N_6392,N_6269,N_6203);
xor U6393 (N_6393,N_6214,N_6277);
or U6394 (N_6394,N_6256,N_6235);
and U6395 (N_6395,N_6229,N_6272);
or U6396 (N_6396,N_6200,N_6291);
nand U6397 (N_6397,N_6272,N_6234);
nor U6398 (N_6398,N_6234,N_6285);
nand U6399 (N_6399,N_6214,N_6227);
xor U6400 (N_6400,N_6302,N_6310);
xnor U6401 (N_6401,N_6397,N_6352);
and U6402 (N_6402,N_6304,N_6359);
or U6403 (N_6403,N_6327,N_6356);
nand U6404 (N_6404,N_6312,N_6399);
or U6405 (N_6405,N_6364,N_6348);
or U6406 (N_6406,N_6370,N_6301);
or U6407 (N_6407,N_6335,N_6340);
xnor U6408 (N_6408,N_6372,N_6366);
xnor U6409 (N_6409,N_6319,N_6326);
and U6410 (N_6410,N_6334,N_6383);
nand U6411 (N_6411,N_6368,N_6306);
nand U6412 (N_6412,N_6393,N_6392);
xor U6413 (N_6413,N_6365,N_6363);
or U6414 (N_6414,N_6336,N_6394);
nand U6415 (N_6415,N_6307,N_6344);
or U6416 (N_6416,N_6305,N_6330);
and U6417 (N_6417,N_6398,N_6373);
xnor U6418 (N_6418,N_6314,N_6390);
xnor U6419 (N_6419,N_6379,N_6369);
nor U6420 (N_6420,N_6382,N_6384);
or U6421 (N_6421,N_6362,N_6331);
nand U6422 (N_6422,N_6388,N_6343);
nor U6423 (N_6423,N_6376,N_6317);
nor U6424 (N_6424,N_6349,N_6357);
nor U6425 (N_6425,N_6371,N_6367);
and U6426 (N_6426,N_6309,N_6389);
xnor U6427 (N_6427,N_6391,N_6300);
xor U6428 (N_6428,N_6361,N_6323);
xor U6429 (N_6429,N_6375,N_6328);
or U6430 (N_6430,N_6347,N_6345);
xnor U6431 (N_6431,N_6346,N_6377);
or U6432 (N_6432,N_6318,N_6316);
nor U6433 (N_6433,N_6341,N_6338);
xnor U6434 (N_6434,N_6321,N_6396);
and U6435 (N_6435,N_6381,N_6303);
xor U6436 (N_6436,N_6322,N_6308);
or U6437 (N_6437,N_6353,N_6315);
xnor U6438 (N_6438,N_6378,N_6351);
nor U6439 (N_6439,N_6320,N_6354);
xnor U6440 (N_6440,N_6395,N_6325);
nand U6441 (N_6441,N_6329,N_6360);
or U6442 (N_6442,N_6333,N_6313);
nor U6443 (N_6443,N_6385,N_6350);
or U6444 (N_6444,N_6380,N_6324);
nor U6445 (N_6445,N_6339,N_6374);
or U6446 (N_6446,N_6342,N_6386);
and U6447 (N_6447,N_6337,N_6355);
nand U6448 (N_6448,N_6311,N_6387);
and U6449 (N_6449,N_6358,N_6332);
and U6450 (N_6450,N_6355,N_6333);
nand U6451 (N_6451,N_6373,N_6305);
xnor U6452 (N_6452,N_6331,N_6340);
nand U6453 (N_6453,N_6339,N_6376);
or U6454 (N_6454,N_6389,N_6399);
nand U6455 (N_6455,N_6301,N_6337);
xor U6456 (N_6456,N_6330,N_6370);
or U6457 (N_6457,N_6306,N_6334);
nor U6458 (N_6458,N_6350,N_6306);
nor U6459 (N_6459,N_6363,N_6393);
nand U6460 (N_6460,N_6377,N_6386);
or U6461 (N_6461,N_6375,N_6387);
xnor U6462 (N_6462,N_6368,N_6399);
and U6463 (N_6463,N_6315,N_6351);
xnor U6464 (N_6464,N_6334,N_6386);
and U6465 (N_6465,N_6359,N_6344);
and U6466 (N_6466,N_6381,N_6364);
and U6467 (N_6467,N_6362,N_6352);
or U6468 (N_6468,N_6392,N_6398);
nand U6469 (N_6469,N_6306,N_6351);
nor U6470 (N_6470,N_6349,N_6394);
and U6471 (N_6471,N_6315,N_6396);
nand U6472 (N_6472,N_6345,N_6367);
and U6473 (N_6473,N_6335,N_6308);
and U6474 (N_6474,N_6378,N_6309);
nand U6475 (N_6475,N_6338,N_6310);
nand U6476 (N_6476,N_6394,N_6319);
xor U6477 (N_6477,N_6381,N_6329);
or U6478 (N_6478,N_6366,N_6380);
xnor U6479 (N_6479,N_6318,N_6378);
and U6480 (N_6480,N_6388,N_6378);
xor U6481 (N_6481,N_6397,N_6355);
nor U6482 (N_6482,N_6340,N_6355);
nand U6483 (N_6483,N_6366,N_6393);
nor U6484 (N_6484,N_6334,N_6378);
nor U6485 (N_6485,N_6369,N_6361);
or U6486 (N_6486,N_6360,N_6375);
nand U6487 (N_6487,N_6374,N_6324);
nand U6488 (N_6488,N_6334,N_6329);
and U6489 (N_6489,N_6353,N_6347);
and U6490 (N_6490,N_6321,N_6356);
nand U6491 (N_6491,N_6308,N_6381);
xor U6492 (N_6492,N_6387,N_6391);
xor U6493 (N_6493,N_6317,N_6303);
nand U6494 (N_6494,N_6315,N_6394);
nand U6495 (N_6495,N_6354,N_6334);
nand U6496 (N_6496,N_6377,N_6315);
nor U6497 (N_6497,N_6391,N_6384);
nor U6498 (N_6498,N_6301,N_6395);
or U6499 (N_6499,N_6352,N_6358);
or U6500 (N_6500,N_6481,N_6491);
nor U6501 (N_6501,N_6425,N_6448);
nor U6502 (N_6502,N_6476,N_6403);
nand U6503 (N_6503,N_6456,N_6486);
xnor U6504 (N_6504,N_6424,N_6437);
nand U6505 (N_6505,N_6413,N_6487);
and U6506 (N_6506,N_6400,N_6494);
and U6507 (N_6507,N_6428,N_6469);
nand U6508 (N_6508,N_6479,N_6452);
or U6509 (N_6509,N_6466,N_6451);
xnor U6510 (N_6510,N_6474,N_6453);
xnor U6511 (N_6511,N_6478,N_6426);
and U6512 (N_6512,N_6421,N_6444);
and U6513 (N_6513,N_6431,N_6475);
nand U6514 (N_6514,N_6446,N_6498);
nand U6515 (N_6515,N_6454,N_6410);
and U6516 (N_6516,N_6439,N_6449);
nor U6517 (N_6517,N_6422,N_6485);
xor U6518 (N_6518,N_6427,N_6461);
xor U6519 (N_6519,N_6489,N_6460);
nor U6520 (N_6520,N_6408,N_6401);
xor U6521 (N_6521,N_6416,N_6418);
nor U6522 (N_6522,N_6441,N_6471);
and U6523 (N_6523,N_6407,N_6457);
nand U6524 (N_6524,N_6462,N_6455);
xnor U6525 (N_6525,N_6402,N_6482);
nand U6526 (N_6526,N_6432,N_6490);
and U6527 (N_6527,N_6405,N_6488);
or U6528 (N_6528,N_6409,N_6419);
nand U6529 (N_6529,N_6499,N_6470);
nand U6530 (N_6530,N_6468,N_6434);
or U6531 (N_6531,N_6406,N_6483);
and U6532 (N_6532,N_6411,N_6433);
or U6533 (N_6533,N_6430,N_6442);
xor U6534 (N_6534,N_6473,N_6484);
nand U6535 (N_6535,N_6492,N_6463);
and U6536 (N_6536,N_6493,N_6495);
or U6537 (N_6537,N_6429,N_6414);
xor U6538 (N_6538,N_6465,N_6459);
nor U6539 (N_6539,N_6497,N_6417);
or U6540 (N_6540,N_6443,N_6436);
nand U6541 (N_6541,N_6464,N_6480);
xor U6542 (N_6542,N_6472,N_6435);
nand U6543 (N_6543,N_6440,N_6412);
and U6544 (N_6544,N_6458,N_6447);
or U6545 (N_6545,N_6415,N_6423);
and U6546 (N_6546,N_6445,N_6477);
or U6547 (N_6547,N_6438,N_6496);
nor U6548 (N_6548,N_6404,N_6467);
or U6549 (N_6549,N_6420,N_6450);
nand U6550 (N_6550,N_6495,N_6435);
xor U6551 (N_6551,N_6479,N_6425);
nor U6552 (N_6552,N_6495,N_6483);
and U6553 (N_6553,N_6441,N_6492);
nand U6554 (N_6554,N_6498,N_6455);
and U6555 (N_6555,N_6431,N_6483);
nand U6556 (N_6556,N_6428,N_6435);
and U6557 (N_6557,N_6461,N_6404);
xnor U6558 (N_6558,N_6416,N_6407);
and U6559 (N_6559,N_6430,N_6405);
or U6560 (N_6560,N_6449,N_6457);
nand U6561 (N_6561,N_6403,N_6444);
and U6562 (N_6562,N_6499,N_6425);
nor U6563 (N_6563,N_6493,N_6462);
xnor U6564 (N_6564,N_6413,N_6473);
or U6565 (N_6565,N_6462,N_6428);
nor U6566 (N_6566,N_6496,N_6452);
and U6567 (N_6567,N_6406,N_6401);
and U6568 (N_6568,N_6474,N_6469);
or U6569 (N_6569,N_6413,N_6498);
xor U6570 (N_6570,N_6460,N_6439);
and U6571 (N_6571,N_6413,N_6472);
nor U6572 (N_6572,N_6463,N_6473);
nor U6573 (N_6573,N_6431,N_6412);
nand U6574 (N_6574,N_6420,N_6432);
nand U6575 (N_6575,N_6489,N_6457);
xnor U6576 (N_6576,N_6424,N_6491);
or U6577 (N_6577,N_6447,N_6424);
nand U6578 (N_6578,N_6432,N_6413);
nor U6579 (N_6579,N_6466,N_6465);
nand U6580 (N_6580,N_6415,N_6400);
nand U6581 (N_6581,N_6449,N_6415);
nor U6582 (N_6582,N_6450,N_6497);
or U6583 (N_6583,N_6450,N_6459);
and U6584 (N_6584,N_6418,N_6493);
xnor U6585 (N_6585,N_6425,N_6465);
xor U6586 (N_6586,N_6480,N_6474);
nor U6587 (N_6587,N_6460,N_6468);
nor U6588 (N_6588,N_6484,N_6498);
or U6589 (N_6589,N_6448,N_6434);
xor U6590 (N_6590,N_6471,N_6411);
nor U6591 (N_6591,N_6441,N_6424);
nand U6592 (N_6592,N_6484,N_6476);
nor U6593 (N_6593,N_6426,N_6441);
nand U6594 (N_6594,N_6404,N_6471);
or U6595 (N_6595,N_6496,N_6484);
nor U6596 (N_6596,N_6430,N_6441);
xor U6597 (N_6597,N_6467,N_6472);
nand U6598 (N_6598,N_6434,N_6415);
nor U6599 (N_6599,N_6496,N_6445);
and U6600 (N_6600,N_6540,N_6573);
and U6601 (N_6601,N_6523,N_6539);
nand U6602 (N_6602,N_6521,N_6530);
nand U6603 (N_6603,N_6544,N_6520);
nor U6604 (N_6604,N_6555,N_6579);
nor U6605 (N_6605,N_6576,N_6558);
or U6606 (N_6606,N_6567,N_6587);
nand U6607 (N_6607,N_6598,N_6514);
or U6608 (N_6608,N_6593,N_6525);
xnor U6609 (N_6609,N_6568,N_6528);
and U6610 (N_6610,N_6585,N_6550);
and U6611 (N_6611,N_6564,N_6578);
nand U6612 (N_6612,N_6575,N_6554);
xnor U6613 (N_6613,N_6592,N_6590);
xnor U6614 (N_6614,N_6556,N_6542);
nor U6615 (N_6615,N_6547,N_6599);
nor U6616 (N_6616,N_6561,N_6529);
nand U6617 (N_6617,N_6511,N_6526);
and U6618 (N_6618,N_6553,N_6566);
or U6619 (N_6619,N_6524,N_6580);
xnor U6620 (N_6620,N_6594,N_6583);
nor U6621 (N_6621,N_6535,N_6551);
nand U6622 (N_6622,N_6517,N_6506);
or U6623 (N_6623,N_6513,N_6571);
and U6624 (N_6624,N_6502,N_6577);
or U6625 (N_6625,N_6512,N_6559);
or U6626 (N_6626,N_6565,N_6563);
xnor U6627 (N_6627,N_6508,N_6536);
and U6628 (N_6628,N_6569,N_6515);
nor U6629 (N_6629,N_6538,N_6545);
nor U6630 (N_6630,N_6533,N_6503);
xnor U6631 (N_6631,N_6591,N_6522);
nand U6632 (N_6632,N_6501,N_6516);
nor U6633 (N_6633,N_6531,N_6509);
and U6634 (N_6634,N_6543,N_6510);
or U6635 (N_6635,N_6562,N_6596);
nand U6636 (N_6636,N_6589,N_6552);
or U6637 (N_6637,N_6504,N_6532);
and U6638 (N_6638,N_6519,N_6582);
nor U6639 (N_6639,N_6574,N_6549);
nand U6640 (N_6640,N_6570,N_6541);
xor U6641 (N_6641,N_6527,N_6548);
xor U6642 (N_6642,N_6588,N_6518);
nand U6643 (N_6643,N_6572,N_6534);
nand U6644 (N_6644,N_6597,N_6507);
and U6645 (N_6645,N_6581,N_6595);
and U6646 (N_6646,N_6500,N_6586);
or U6647 (N_6647,N_6546,N_6560);
or U6648 (N_6648,N_6537,N_6584);
xnor U6649 (N_6649,N_6505,N_6557);
and U6650 (N_6650,N_6528,N_6502);
xnor U6651 (N_6651,N_6580,N_6597);
xor U6652 (N_6652,N_6573,N_6590);
or U6653 (N_6653,N_6514,N_6587);
and U6654 (N_6654,N_6594,N_6540);
nand U6655 (N_6655,N_6515,N_6575);
nand U6656 (N_6656,N_6501,N_6555);
and U6657 (N_6657,N_6544,N_6545);
or U6658 (N_6658,N_6554,N_6541);
and U6659 (N_6659,N_6583,N_6517);
and U6660 (N_6660,N_6567,N_6508);
xor U6661 (N_6661,N_6574,N_6536);
or U6662 (N_6662,N_6597,N_6518);
xor U6663 (N_6663,N_6515,N_6580);
and U6664 (N_6664,N_6513,N_6501);
and U6665 (N_6665,N_6511,N_6589);
or U6666 (N_6666,N_6576,N_6569);
nor U6667 (N_6667,N_6522,N_6594);
xor U6668 (N_6668,N_6577,N_6584);
nor U6669 (N_6669,N_6587,N_6516);
and U6670 (N_6670,N_6515,N_6534);
nor U6671 (N_6671,N_6598,N_6541);
nor U6672 (N_6672,N_6571,N_6558);
nand U6673 (N_6673,N_6549,N_6504);
and U6674 (N_6674,N_6589,N_6505);
nand U6675 (N_6675,N_6544,N_6566);
nand U6676 (N_6676,N_6519,N_6549);
nand U6677 (N_6677,N_6523,N_6597);
xor U6678 (N_6678,N_6510,N_6598);
nand U6679 (N_6679,N_6519,N_6515);
nor U6680 (N_6680,N_6563,N_6556);
and U6681 (N_6681,N_6518,N_6504);
nor U6682 (N_6682,N_6562,N_6513);
nor U6683 (N_6683,N_6529,N_6585);
and U6684 (N_6684,N_6518,N_6572);
nand U6685 (N_6685,N_6514,N_6512);
nor U6686 (N_6686,N_6579,N_6509);
xor U6687 (N_6687,N_6501,N_6588);
or U6688 (N_6688,N_6534,N_6599);
nor U6689 (N_6689,N_6598,N_6559);
or U6690 (N_6690,N_6581,N_6527);
and U6691 (N_6691,N_6546,N_6541);
nand U6692 (N_6692,N_6530,N_6508);
xnor U6693 (N_6693,N_6570,N_6542);
nor U6694 (N_6694,N_6546,N_6595);
and U6695 (N_6695,N_6548,N_6572);
xor U6696 (N_6696,N_6522,N_6589);
nand U6697 (N_6697,N_6543,N_6558);
nor U6698 (N_6698,N_6596,N_6547);
and U6699 (N_6699,N_6541,N_6594);
xor U6700 (N_6700,N_6674,N_6683);
nor U6701 (N_6701,N_6623,N_6648);
or U6702 (N_6702,N_6620,N_6660);
nand U6703 (N_6703,N_6645,N_6621);
and U6704 (N_6704,N_6639,N_6666);
or U6705 (N_6705,N_6644,N_6695);
nand U6706 (N_6706,N_6676,N_6687);
and U6707 (N_6707,N_6668,N_6651);
or U6708 (N_6708,N_6664,N_6632);
nor U6709 (N_6709,N_6698,N_6633);
nor U6710 (N_6710,N_6663,N_6671);
nand U6711 (N_6711,N_6619,N_6694);
and U6712 (N_6712,N_6605,N_6679);
xor U6713 (N_6713,N_6691,N_6685);
and U6714 (N_6714,N_6653,N_6613);
or U6715 (N_6715,N_6675,N_6690);
nor U6716 (N_6716,N_6641,N_6678);
xor U6717 (N_6717,N_6681,N_6670);
and U6718 (N_6718,N_6657,N_6684);
nand U6719 (N_6719,N_6600,N_6680);
or U6720 (N_6720,N_6649,N_6667);
nor U6721 (N_6721,N_6661,N_6672);
or U6722 (N_6722,N_6601,N_6636);
and U6723 (N_6723,N_6617,N_6658);
or U6724 (N_6724,N_6665,N_6616);
nand U6725 (N_6725,N_6618,N_6608);
or U6726 (N_6726,N_6693,N_6630);
xor U6727 (N_6727,N_6642,N_6686);
nor U6728 (N_6728,N_6647,N_6629);
and U6729 (N_6729,N_6602,N_6606);
xor U6730 (N_6730,N_6699,N_6638);
xor U6731 (N_6731,N_6628,N_6614);
nand U6732 (N_6732,N_6626,N_6688);
and U6733 (N_6733,N_6662,N_6615);
nor U6734 (N_6734,N_6677,N_6656);
xor U6735 (N_6735,N_6655,N_6610);
nand U6736 (N_6736,N_6682,N_6609);
or U6737 (N_6737,N_6692,N_6697);
nor U6738 (N_6738,N_6673,N_6627);
and U6739 (N_6739,N_6631,N_6603);
or U6740 (N_6740,N_6640,N_6652);
nand U6741 (N_6741,N_6624,N_6637);
nand U6742 (N_6742,N_6689,N_6607);
or U6743 (N_6743,N_6604,N_6696);
and U6744 (N_6744,N_6646,N_6612);
and U6745 (N_6745,N_6659,N_6634);
nor U6746 (N_6746,N_6635,N_6669);
nor U6747 (N_6747,N_6625,N_6643);
nand U6748 (N_6748,N_6611,N_6650);
nand U6749 (N_6749,N_6654,N_6622);
and U6750 (N_6750,N_6657,N_6665);
xor U6751 (N_6751,N_6634,N_6635);
xor U6752 (N_6752,N_6644,N_6615);
and U6753 (N_6753,N_6641,N_6698);
and U6754 (N_6754,N_6677,N_6636);
nor U6755 (N_6755,N_6619,N_6668);
nand U6756 (N_6756,N_6697,N_6677);
and U6757 (N_6757,N_6688,N_6641);
xor U6758 (N_6758,N_6637,N_6686);
or U6759 (N_6759,N_6645,N_6675);
nand U6760 (N_6760,N_6652,N_6649);
nor U6761 (N_6761,N_6648,N_6681);
or U6762 (N_6762,N_6668,N_6638);
or U6763 (N_6763,N_6652,N_6675);
or U6764 (N_6764,N_6674,N_6646);
nor U6765 (N_6765,N_6625,N_6618);
or U6766 (N_6766,N_6661,N_6665);
xor U6767 (N_6767,N_6639,N_6600);
xor U6768 (N_6768,N_6639,N_6648);
nand U6769 (N_6769,N_6689,N_6690);
nor U6770 (N_6770,N_6642,N_6690);
and U6771 (N_6771,N_6638,N_6675);
nand U6772 (N_6772,N_6613,N_6684);
xor U6773 (N_6773,N_6670,N_6693);
and U6774 (N_6774,N_6659,N_6658);
nand U6775 (N_6775,N_6663,N_6625);
xnor U6776 (N_6776,N_6616,N_6645);
nand U6777 (N_6777,N_6612,N_6698);
nor U6778 (N_6778,N_6648,N_6689);
and U6779 (N_6779,N_6671,N_6612);
or U6780 (N_6780,N_6603,N_6677);
or U6781 (N_6781,N_6683,N_6671);
xor U6782 (N_6782,N_6621,N_6656);
and U6783 (N_6783,N_6684,N_6602);
nor U6784 (N_6784,N_6636,N_6625);
and U6785 (N_6785,N_6681,N_6636);
xnor U6786 (N_6786,N_6691,N_6661);
nand U6787 (N_6787,N_6644,N_6658);
or U6788 (N_6788,N_6695,N_6696);
and U6789 (N_6789,N_6643,N_6627);
nand U6790 (N_6790,N_6680,N_6605);
nand U6791 (N_6791,N_6650,N_6685);
xnor U6792 (N_6792,N_6690,N_6614);
xnor U6793 (N_6793,N_6672,N_6602);
or U6794 (N_6794,N_6630,N_6622);
xor U6795 (N_6795,N_6638,N_6647);
nand U6796 (N_6796,N_6628,N_6698);
or U6797 (N_6797,N_6637,N_6673);
xor U6798 (N_6798,N_6652,N_6646);
or U6799 (N_6799,N_6651,N_6694);
and U6800 (N_6800,N_6702,N_6796);
nand U6801 (N_6801,N_6715,N_6778);
and U6802 (N_6802,N_6795,N_6794);
nand U6803 (N_6803,N_6741,N_6714);
and U6804 (N_6804,N_6746,N_6770);
and U6805 (N_6805,N_6747,N_6776);
nor U6806 (N_6806,N_6701,N_6716);
and U6807 (N_6807,N_6768,N_6775);
xor U6808 (N_6808,N_6729,N_6744);
nand U6809 (N_6809,N_6756,N_6750);
xor U6810 (N_6810,N_6751,N_6738);
nor U6811 (N_6811,N_6748,N_6730);
xor U6812 (N_6812,N_6766,N_6703);
xnor U6813 (N_6813,N_6718,N_6725);
and U6814 (N_6814,N_6710,N_6798);
xor U6815 (N_6815,N_6784,N_6742);
nand U6816 (N_6816,N_6743,N_6781);
nand U6817 (N_6817,N_6779,N_6731);
or U6818 (N_6818,N_6787,N_6704);
or U6819 (N_6819,N_6723,N_6722);
or U6820 (N_6820,N_6732,N_6760);
xor U6821 (N_6821,N_6792,N_6758);
xor U6822 (N_6822,N_6774,N_6736);
or U6823 (N_6823,N_6745,N_6724);
xor U6824 (N_6824,N_6783,N_6734);
nor U6825 (N_6825,N_6720,N_6777);
xnor U6826 (N_6826,N_6754,N_6739);
and U6827 (N_6827,N_6790,N_6762);
or U6828 (N_6828,N_6717,N_6761);
nand U6829 (N_6829,N_6728,N_6763);
and U6830 (N_6830,N_6772,N_6764);
nor U6831 (N_6831,N_6767,N_6769);
nand U6832 (N_6832,N_6719,N_6785);
nor U6833 (N_6833,N_6780,N_6727);
nand U6834 (N_6834,N_6735,N_6757);
and U6835 (N_6835,N_6786,N_6713);
nor U6836 (N_6836,N_6733,N_6711);
nand U6837 (N_6837,N_6782,N_6706);
and U6838 (N_6838,N_6705,N_6712);
nand U6839 (N_6839,N_6753,N_6740);
nand U6840 (N_6840,N_6737,N_6708);
or U6841 (N_6841,N_6771,N_6726);
nor U6842 (N_6842,N_6759,N_6755);
nor U6843 (N_6843,N_6721,N_6765);
xnor U6844 (N_6844,N_6700,N_6749);
nand U6845 (N_6845,N_6788,N_6707);
nor U6846 (N_6846,N_6793,N_6789);
and U6847 (N_6847,N_6709,N_6752);
xnor U6848 (N_6848,N_6799,N_6797);
xnor U6849 (N_6849,N_6791,N_6773);
nor U6850 (N_6850,N_6749,N_6725);
or U6851 (N_6851,N_6792,N_6721);
nand U6852 (N_6852,N_6795,N_6721);
nand U6853 (N_6853,N_6715,N_6714);
xor U6854 (N_6854,N_6712,N_6787);
nand U6855 (N_6855,N_6771,N_6792);
nor U6856 (N_6856,N_6749,N_6751);
or U6857 (N_6857,N_6742,N_6733);
and U6858 (N_6858,N_6712,N_6745);
or U6859 (N_6859,N_6777,N_6738);
nand U6860 (N_6860,N_6773,N_6799);
and U6861 (N_6861,N_6773,N_6760);
or U6862 (N_6862,N_6763,N_6723);
xnor U6863 (N_6863,N_6782,N_6769);
and U6864 (N_6864,N_6772,N_6769);
or U6865 (N_6865,N_6731,N_6755);
nor U6866 (N_6866,N_6707,N_6722);
and U6867 (N_6867,N_6722,N_6700);
or U6868 (N_6868,N_6712,N_6795);
nand U6869 (N_6869,N_6798,N_6768);
and U6870 (N_6870,N_6767,N_6729);
xnor U6871 (N_6871,N_6700,N_6736);
and U6872 (N_6872,N_6767,N_6725);
and U6873 (N_6873,N_6711,N_6764);
or U6874 (N_6874,N_6765,N_6738);
or U6875 (N_6875,N_6741,N_6754);
or U6876 (N_6876,N_6712,N_6761);
nor U6877 (N_6877,N_6743,N_6744);
and U6878 (N_6878,N_6775,N_6742);
xor U6879 (N_6879,N_6731,N_6703);
nand U6880 (N_6880,N_6739,N_6779);
nor U6881 (N_6881,N_6791,N_6703);
and U6882 (N_6882,N_6790,N_6764);
or U6883 (N_6883,N_6759,N_6770);
xnor U6884 (N_6884,N_6727,N_6752);
nor U6885 (N_6885,N_6781,N_6706);
nand U6886 (N_6886,N_6744,N_6724);
nand U6887 (N_6887,N_6718,N_6777);
and U6888 (N_6888,N_6731,N_6727);
xor U6889 (N_6889,N_6760,N_6762);
nor U6890 (N_6890,N_6758,N_6762);
nand U6891 (N_6891,N_6747,N_6710);
and U6892 (N_6892,N_6709,N_6726);
xnor U6893 (N_6893,N_6750,N_6724);
and U6894 (N_6894,N_6749,N_6762);
nor U6895 (N_6895,N_6793,N_6780);
or U6896 (N_6896,N_6760,N_6796);
and U6897 (N_6897,N_6731,N_6788);
xor U6898 (N_6898,N_6737,N_6749);
nand U6899 (N_6899,N_6715,N_6745);
xor U6900 (N_6900,N_6896,N_6865);
nand U6901 (N_6901,N_6873,N_6877);
xnor U6902 (N_6902,N_6843,N_6881);
nand U6903 (N_6903,N_6889,N_6888);
xnor U6904 (N_6904,N_6810,N_6812);
or U6905 (N_6905,N_6808,N_6869);
xor U6906 (N_6906,N_6803,N_6833);
nor U6907 (N_6907,N_6838,N_6826);
and U6908 (N_6908,N_6832,N_6847);
and U6909 (N_6909,N_6876,N_6858);
nor U6910 (N_6910,N_6872,N_6837);
and U6911 (N_6911,N_6874,N_6816);
nand U6912 (N_6912,N_6886,N_6897);
and U6913 (N_6913,N_6829,N_6887);
nand U6914 (N_6914,N_6892,N_6890);
and U6915 (N_6915,N_6862,N_6813);
and U6916 (N_6916,N_6854,N_6822);
nor U6917 (N_6917,N_6853,N_6864);
nor U6918 (N_6918,N_6861,N_6821);
nand U6919 (N_6919,N_6806,N_6866);
xor U6920 (N_6920,N_6805,N_6856);
nor U6921 (N_6921,N_6840,N_6824);
or U6922 (N_6922,N_6834,N_6857);
or U6923 (N_6923,N_6885,N_6894);
nand U6924 (N_6924,N_6804,N_6819);
and U6925 (N_6925,N_6802,N_6817);
or U6926 (N_6926,N_6844,N_6851);
and U6927 (N_6927,N_6898,N_6875);
nor U6928 (N_6928,N_6823,N_6883);
nor U6929 (N_6929,N_6839,N_6882);
and U6930 (N_6930,N_6818,N_6871);
or U6931 (N_6931,N_6878,N_6842);
or U6932 (N_6932,N_6893,N_6841);
nand U6933 (N_6933,N_6846,N_6863);
nor U6934 (N_6934,N_6868,N_6849);
nand U6935 (N_6935,N_6855,N_6830);
xor U6936 (N_6936,N_6801,N_6811);
nor U6937 (N_6937,N_6850,N_6867);
and U6938 (N_6938,N_6827,N_6880);
and U6939 (N_6939,N_6828,N_6859);
or U6940 (N_6940,N_6879,N_6835);
xnor U6941 (N_6941,N_6891,N_6860);
or U6942 (N_6942,N_6845,N_6825);
xnor U6943 (N_6943,N_6815,N_6831);
nand U6944 (N_6944,N_6809,N_6848);
or U6945 (N_6945,N_6820,N_6895);
and U6946 (N_6946,N_6870,N_6884);
xnor U6947 (N_6947,N_6836,N_6852);
and U6948 (N_6948,N_6899,N_6814);
or U6949 (N_6949,N_6807,N_6800);
nor U6950 (N_6950,N_6828,N_6812);
xor U6951 (N_6951,N_6875,N_6831);
or U6952 (N_6952,N_6849,N_6801);
xor U6953 (N_6953,N_6827,N_6856);
or U6954 (N_6954,N_6871,N_6809);
or U6955 (N_6955,N_6899,N_6862);
nand U6956 (N_6956,N_6858,N_6837);
or U6957 (N_6957,N_6882,N_6800);
nor U6958 (N_6958,N_6895,N_6801);
and U6959 (N_6959,N_6841,N_6830);
xnor U6960 (N_6960,N_6890,N_6806);
nand U6961 (N_6961,N_6850,N_6815);
xnor U6962 (N_6962,N_6827,N_6862);
nand U6963 (N_6963,N_6895,N_6880);
or U6964 (N_6964,N_6837,N_6852);
nor U6965 (N_6965,N_6800,N_6841);
or U6966 (N_6966,N_6827,N_6819);
nand U6967 (N_6967,N_6894,N_6800);
nand U6968 (N_6968,N_6886,N_6830);
or U6969 (N_6969,N_6876,N_6809);
nand U6970 (N_6970,N_6849,N_6880);
nor U6971 (N_6971,N_6824,N_6867);
and U6972 (N_6972,N_6880,N_6815);
xor U6973 (N_6973,N_6885,N_6829);
and U6974 (N_6974,N_6852,N_6891);
xnor U6975 (N_6975,N_6816,N_6831);
and U6976 (N_6976,N_6866,N_6864);
xor U6977 (N_6977,N_6844,N_6892);
nand U6978 (N_6978,N_6845,N_6807);
xor U6979 (N_6979,N_6810,N_6872);
nand U6980 (N_6980,N_6869,N_6839);
and U6981 (N_6981,N_6832,N_6817);
xnor U6982 (N_6982,N_6805,N_6825);
nor U6983 (N_6983,N_6868,N_6881);
or U6984 (N_6984,N_6870,N_6815);
or U6985 (N_6985,N_6800,N_6837);
nand U6986 (N_6986,N_6882,N_6812);
nor U6987 (N_6987,N_6830,N_6836);
xor U6988 (N_6988,N_6872,N_6877);
nor U6989 (N_6989,N_6827,N_6871);
xnor U6990 (N_6990,N_6824,N_6893);
xnor U6991 (N_6991,N_6822,N_6808);
or U6992 (N_6992,N_6825,N_6868);
nor U6993 (N_6993,N_6870,N_6883);
nand U6994 (N_6994,N_6812,N_6893);
nor U6995 (N_6995,N_6845,N_6867);
or U6996 (N_6996,N_6805,N_6867);
nand U6997 (N_6997,N_6833,N_6812);
or U6998 (N_6998,N_6849,N_6881);
xnor U6999 (N_6999,N_6801,N_6826);
nor U7000 (N_7000,N_6990,N_6932);
and U7001 (N_7001,N_6948,N_6911);
nand U7002 (N_7002,N_6902,N_6951);
and U7003 (N_7003,N_6942,N_6927);
nor U7004 (N_7004,N_6936,N_6999);
nor U7005 (N_7005,N_6979,N_6986);
and U7006 (N_7006,N_6925,N_6916);
nor U7007 (N_7007,N_6947,N_6995);
nor U7008 (N_7008,N_6973,N_6929);
and U7009 (N_7009,N_6949,N_6970);
and U7010 (N_7010,N_6953,N_6921);
nand U7011 (N_7011,N_6993,N_6908);
and U7012 (N_7012,N_6981,N_6969);
or U7013 (N_7013,N_6987,N_6914);
nor U7014 (N_7014,N_6904,N_6923);
and U7015 (N_7015,N_6919,N_6937);
xor U7016 (N_7016,N_6913,N_6955);
nor U7017 (N_7017,N_6985,N_6954);
nand U7018 (N_7018,N_6906,N_6940);
xnor U7019 (N_7019,N_6938,N_6967);
and U7020 (N_7020,N_6971,N_6997);
nor U7021 (N_7021,N_6945,N_6968);
nor U7022 (N_7022,N_6909,N_6966);
xor U7023 (N_7023,N_6978,N_6934);
xor U7024 (N_7024,N_6939,N_6918);
or U7025 (N_7025,N_6996,N_6984);
nor U7026 (N_7026,N_6964,N_6912);
and U7027 (N_7027,N_6907,N_6980);
or U7028 (N_7028,N_6983,N_6952);
nor U7029 (N_7029,N_6900,N_6910);
or U7030 (N_7030,N_6957,N_6962);
or U7031 (N_7031,N_6950,N_6961);
or U7032 (N_7032,N_6920,N_6931);
xor U7033 (N_7033,N_6956,N_6989);
and U7034 (N_7034,N_6905,N_6901);
and U7035 (N_7035,N_6958,N_6965);
and U7036 (N_7036,N_6998,N_6992);
and U7037 (N_7037,N_6928,N_6994);
xnor U7038 (N_7038,N_6935,N_6922);
xnor U7039 (N_7039,N_6988,N_6975);
xnor U7040 (N_7040,N_6915,N_6959);
nand U7041 (N_7041,N_6972,N_6924);
or U7042 (N_7042,N_6944,N_6963);
nor U7043 (N_7043,N_6943,N_6976);
or U7044 (N_7044,N_6926,N_6933);
xor U7045 (N_7045,N_6946,N_6903);
or U7046 (N_7046,N_6982,N_6941);
and U7047 (N_7047,N_6917,N_6977);
nor U7048 (N_7048,N_6991,N_6930);
or U7049 (N_7049,N_6960,N_6974);
or U7050 (N_7050,N_6953,N_6975);
or U7051 (N_7051,N_6966,N_6986);
or U7052 (N_7052,N_6945,N_6961);
xor U7053 (N_7053,N_6983,N_6997);
or U7054 (N_7054,N_6937,N_6954);
or U7055 (N_7055,N_6916,N_6994);
or U7056 (N_7056,N_6937,N_6952);
and U7057 (N_7057,N_6960,N_6933);
and U7058 (N_7058,N_6980,N_6994);
and U7059 (N_7059,N_6922,N_6939);
and U7060 (N_7060,N_6967,N_6911);
xnor U7061 (N_7061,N_6991,N_6999);
nor U7062 (N_7062,N_6926,N_6979);
and U7063 (N_7063,N_6939,N_6949);
or U7064 (N_7064,N_6980,N_6937);
and U7065 (N_7065,N_6941,N_6954);
or U7066 (N_7066,N_6997,N_6994);
nand U7067 (N_7067,N_6908,N_6977);
or U7068 (N_7068,N_6965,N_6988);
or U7069 (N_7069,N_6940,N_6900);
and U7070 (N_7070,N_6915,N_6985);
nor U7071 (N_7071,N_6998,N_6959);
nor U7072 (N_7072,N_6918,N_6952);
or U7073 (N_7073,N_6902,N_6914);
and U7074 (N_7074,N_6901,N_6951);
and U7075 (N_7075,N_6958,N_6911);
and U7076 (N_7076,N_6904,N_6976);
nand U7077 (N_7077,N_6978,N_6963);
xnor U7078 (N_7078,N_6908,N_6912);
nor U7079 (N_7079,N_6994,N_6990);
and U7080 (N_7080,N_6906,N_6949);
xor U7081 (N_7081,N_6917,N_6953);
nand U7082 (N_7082,N_6967,N_6939);
xor U7083 (N_7083,N_6971,N_6932);
or U7084 (N_7084,N_6956,N_6904);
or U7085 (N_7085,N_6967,N_6916);
nand U7086 (N_7086,N_6932,N_6931);
or U7087 (N_7087,N_6971,N_6937);
nand U7088 (N_7088,N_6950,N_6980);
nand U7089 (N_7089,N_6980,N_6959);
nor U7090 (N_7090,N_6975,N_6940);
xnor U7091 (N_7091,N_6967,N_6958);
nand U7092 (N_7092,N_6951,N_6989);
nor U7093 (N_7093,N_6979,N_6911);
nor U7094 (N_7094,N_6922,N_6987);
or U7095 (N_7095,N_6957,N_6943);
nor U7096 (N_7096,N_6936,N_6993);
or U7097 (N_7097,N_6915,N_6968);
nor U7098 (N_7098,N_6939,N_6974);
xor U7099 (N_7099,N_6938,N_6901);
or U7100 (N_7100,N_7071,N_7083);
nor U7101 (N_7101,N_7064,N_7041);
nand U7102 (N_7102,N_7079,N_7056);
nand U7103 (N_7103,N_7075,N_7039);
and U7104 (N_7104,N_7050,N_7043);
nand U7105 (N_7105,N_7065,N_7017);
and U7106 (N_7106,N_7091,N_7057);
nand U7107 (N_7107,N_7018,N_7035);
nand U7108 (N_7108,N_7037,N_7098);
and U7109 (N_7109,N_7070,N_7021);
or U7110 (N_7110,N_7047,N_7006);
xor U7111 (N_7111,N_7090,N_7030);
xnor U7112 (N_7112,N_7012,N_7024);
xnor U7113 (N_7113,N_7088,N_7069);
or U7114 (N_7114,N_7027,N_7080);
or U7115 (N_7115,N_7093,N_7082);
xor U7116 (N_7116,N_7084,N_7058);
and U7117 (N_7117,N_7061,N_7092);
nand U7118 (N_7118,N_7087,N_7042);
nand U7119 (N_7119,N_7044,N_7010);
or U7120 (N_7120,N_7081,N_7066);
xnor U7121 (N_7121,N_7029,N_7094);
or U7122 (N_7122,N_7063,N_7004);
nand U7123 (N_7123,N_7074,N_7099);
xnor U7124 (N_7124,N_7073,N_7055);
and U7125 (N_7125,N_7023,N_7059);
xnor U7126 (N_7126,N_7005,N_7048);
nor U7127 (N_7127,N_7009,N_7095);
xor U7128 (N_7128,N_7013,N_7001);
nand U7129 (N_7129,N_7068,N_7078);
nand U7130 (N_7130,N_7089,N_7034);
nand U7131 (N_7131,N_7000,N_7077);
or U7132 (N_7132,N_7049,N_7085);
xor U7133 (N_7133,N_7015,N_7019);
or U7134 (N_7134,N_7003,N_7002);
or U7135 (N_7135,N_7067,N_7026);
or U7136 (N_7136,N_7045,N_7038);
nand U7137 (N_7137,N_7086,N_7040);
or U7138 (N_7138,N_7060,N_7076);
or U7139 (N_7139,N_7072,N_7062);
or U7140 (N_7140,N_7007,N_7097);
nor U7141 (N_7141,N_7016,N_7096);
nor U7142 (N_7142,N_7022,N_7025);
xor U7143 (N_7143,N_7032,N_7033);
and U7144 (N_7144,N_7031,N_7054);
and U7145 (N_7145,N_7053,N_7028);
and U7146 (N_7146,N_7046,N_7014);
nand U7147 (N_7147,N_7020,N_7052);
nor U7148 (N_7148,N_7036,N_7011);
nand U7149 (N_7149,N_7051,N_7008);
and U7150 (N_7150,N_7037,N_7070);
nor U7151 (N_7151,N_7073,N_7005);
nor U7152 (N_7152,N_7054,N_7099);
nor U7153 (N_7153,N_7016,N_7020);
and U7154 (N_7154,N_7055,N_7029);
nor U7155 (N_7155,N_7070,N_7066);
nor U7156 (N_7156,N_7033,N_7036);
or U7157 (N_7157,N_7052,N_7019);
nor U7158 (N_7158,N_7033,N_7010);
nor U7159 (N_7159,N_7091,N_7090);
and U7160 (N_7160,N_7096,N_7014);
xor U7161 (N_7161,N_7084,N_7047);
nand U7162 (N_7162,N_7080,N_7049);
or U7163 (N_7163,N_7034,N_7076);
nor U7164 (N_7164,N_7060,N_7036);
xnor U7165 (N_7165,N_7016,N_7064);
nand U7166 (N_7166,N_7041,N_7069);
nand U7167 (N_7167,N_7041,N_7003);
and U7168 (N_7168,N_7048,N_7084);
nor U7169 (N_7169,N_7037,N_7042);
xnor U7170 (N_7170,N_7004,N_7013);
nor U7171 (N_7171,N_7016,N_7089);
xor U7172 (N_7172,N_7021,N_7071);
nand U7173 (N_7173,N_7000,N_7082);
nand U7174 (N_7174,N_7001,N_7023);
nand U7175 (N_7175,N_7010,N_7003);
nor U7176 (N_7176,N_7014,N_7048);
xnor U7177 (N_7177,N_7016,N_7042);
nand U7178 (N_7178,N_7005,N_7034);
nand U7179 (N_7179,N_7001,N_7091);
nand U7180 (N_7180,N_7058,N_7032);
nor U7181 (N_7181,N_7002,N_7013);
nand U7182 (N_7182,N_7015,N_7086);
and U7183 (N_7183,N_7042,N_7094);
nor U7184 (N_7184,N_7082,N_7008);
nand U7185 (N_7185,N_7026,N_7078);
xnor U7186 (N_7186,N_7092,N_7088);
nand U7187 (N_7187,N_7030,N_7008);
and U7188 (N_7188,N_7044,N_7091);
or U7189 (N_7189,N_7084,N_7083);
or U7190 (N_7190,N_7010,N_7041);
nor U7191 (N_7191,N_7068,N_7037);
or U7192 (N_7192,N_7066,N_7054);
nor U7193 (N_7193,N_7017,N_7069);
nor U7194 (N_7194,N_7057,N_7065);
xnor U7195 (N_7195,N_7019,N_7083);
and U7196 (N_7196,N_7024,N_7022);
nand U7197 (N_7197,N_7043,N_7021);
nor U7198 (N_7198,N_7090,N_7003);
nor U7199 (N_7199,N_7050,N_7033);
xor U7200 (N_7200,N_7196,N_7169);
xnor U7201 (N_7201,N_7178,N_7154);
or U7202 (N_7202,N_7129,N_7122);
and U7203 (N_7203,N_7137,N_7174);
and U7204 (N_7204,N_7111,N_7160);
and U7205 (N_7205,N_7181,N_7172);
and U7206 (N_7206,N_7188,N_7130);
xor U7207 (N_7207,N_7110,N_7125);
xor U7208 (N_7208,N_7153,N_7197);
or U7209 (N_7209,N_7113,N_7162);
and U7210 (N_7210,N_7107,N_7164);
or U7211 (N_7211,N_7141,N_7190);
nand U7212 (N_7212,N_7185,N_7195);
or U7213 (N_7213,N_7100,N_7134);
nor U7214 (N_7214,N_7124,N_7186);
nand U7215 (N_7215,N_7118,N_7131);
xor U7216 (N_7216,N_7191,N_7170);
xor U7217 (N_7217,N_7147,N_7187);
nand U7218 (N_7218,N_7114,N_7192);
or U7219 (N_7219,N_7126,N_7123);
nand U7220 (N_7220,N_7158,N_7199);
or U7221 (N_7221,N_7183,N_7151);
xor U7222 (N_7222,N_7136,N_7109);
nor U7223 (N_7223,N_7142,N_7152);
nor U7224 (N_7224,N_7193,N_7106);
or U7225 (N_7225,N_7104,N_7117);
and U7226 (N_7226,N_7182,N_7133);
xnor U7227 (N_7227,N_7144,N_7140);
nand U7228 (N_7228,N_7177,N_7116);
xor U7229 (N_7229,N_7179,N_7156);
nor U7230 (N_7230,N_7120,N_7128);
nor U7231 (N_7231,N_7161,N_7119);
or U7232 (N_7232,N_7139,N_7115);
or U7233 (N_7233,N_7102,N_7103);
xnor U7234 (N_7234,N_7155,N_7108);
and U7235 (N_7235,N_7132,N_7145);
nor U7236 (N_7236,N_7105,N_7135);
nand U7237 (N_7237,N_7173,N_7112);
nor U7238 (N_7238,N_7167,N_7143);
and U7239 (N_7239,N_7138,N_7149);
nor U7240 (N_7240,N_7175,N_7157);
nor U7241 (N_7241,N_7146,N_7184);
xnor U7242 (N_7242,N_7127,N_7163);
xnor U7243 (N_7243,N_7176,N_7101);
nor U7244 (N_7244,N_7180,N_7171);
nand U7245 (N_7245,N_7189,N_7198);
xnor U7246 (N_7246,N_7159,N_7148);
xnor U7247 (N_7247,N_7168,N_7121);
nand U7248 (N_7248,N_7194,N_7166);
xor U7249 (N_7249,N_7150,N_7165);
nand U7250 (N_7250,N_7135,N_7136);
nand U7251 (N_7251,N_7173,N_7178);
and U7252 (N_7252,N_7181,N_7158);
or U7253 (N_7253,N_7169,N_7189);
nand U7254 (N_7254,N_7132,N_7144);
or U7255 (N_7255,N_7197,N_7110);
and U7256 (N_7256,N_7175,N_7156);
and U7257 (N_7257,N_7164,N_7115);
and U7258 (N_7258,N_7173,N_7117);
or U7259 (N_7259,N_7172,N_7113);
and U7260 (N_7260,N_7130,N_7143);
or U7261 (N_7261,N_7108,N_7193);
or U7262 (N_7262,N_7190,N_7170);
nand U7263 (N_7263,N_7128,N_7110);
nor U7264 (N_7264,N_7120,N_7198);
or U7265 (N_7265,N_7124,N_7183);
nand U7266 (N_7266,N_7172,N_7176);
nor U7267 (N_7267,N_7109,N_7187);
or U7268 (N_7268,N_7108,N_7158);
or U7269 (N_7269,N_7189,N_7171);
and U7270 (N_7270,N_7129,N_7137);
xnor U7271 (N_7271,N_7119,N_7125);
xnor U7272 (N_7272,N_7116,N_7169);
or U7273 (N_7273,N_7103,N_7195);
nand U7274 (N_7274,N_7107,N_7150);
and U7275 (N_7275,N_7124,N_7108);
xnor U7276 (N_7276,N_7177,N_7162);
or U7277 (N_7277,N_7159,N_7115);
and U7278 (N_7278,N_7172,N_7125);
xor U7279 (N_7279,N_7104,N_7142);
nand U7280 (N_7280,N_7172,N_7153);
or U7281 (N_7281,N_7195,N_7176);
nor U7282 (N_7282,N_7192,N_7167);
xnor U7283 (N_7283,N_7154,N_7132);
nor U7284 (N_7284,N_7120,N_7174);
nand U7285 (N_7285,N_7144,N_7124);
nor U7286 (N_7286,N_7158,N_7176);
or U7287 (N_7287,N_7166,N_7171);
or U7288 (N_7288,N_7134,N_7141);
and U7289 (N_7289,N_7130,N_7115);
xor U7290 (N_7290,N_7121,N_7135);
nand U7291 (N_7291,N_7121,N_7107);
xor U7292 (N_7292,N_7166,N_7193);
xor U7293 (N_7293,N_7161,N_7110);
xor U7294 (N_7294,N_7120,N_7148);
xor U7295 (N_7295,N_7110,N_7136);
nor U7296 (N_7296,N_7169,N_7184);
or U7297 (N_7297,N_7151,N_7144);
xnor U7298 (N_7298,N_7125,N_7147);
nand U7299 (N_7299,N_7127,N_7162);
and U7300 (N_7300,N_7213,N_7212);
nand U7301 (N_7301,N_7205,N_7224);
or U7302 (N_7302,N_7215,N_7277);
nand U7303 (N_7303,N_7241,N_7225);
nor U7304 (N_7304,N_7229,N_7282);
nand U7305 (N_7305,N_7231,N_7246);
xor U7306 (N_7306,N_7264,N_7216);
or U7307 (N_7307,N_7263,N_7297);
nand U7308 (N_7308,N_7296,N_7257);
and U7309 (N_7309,N_7242,N_7208);
or U7310 (N_7310,N_7261,N_7283);
xnor U7311 (N_7311,N_7221,N_7291);
and U7312 (N_7312,N_7244,N_7211);
nand U7313 (N_7313,N_7201,N_7295);
nor U7314 (N_7314,N_7299,N_7259);
nand U7315 (N_7315,N_7218,N_7293);
nand U7316 (N_7316,N_7265,N_7228);
nor U7317 (N_7317,N_7274,N_7279);
nand U7318 (N_7318,N_7234,N_7220);
and U7319 (N_7319,N_7253,N_7239);
nand U7320 (N_7320,N_7247,N_7210);
nand U7321 (N_7321,N_7203,N_7271);
or U7322 (N_7322,N_7272,N_7290);
nor U7323 (N_7323,N_7285,N_7280);
and U7324 (N_7324,N_7245,N_7238);
nand U7325 (N_7325,N_7266,N_7204);
and U7326 (N_7326,N_7226,N_7292);
xor U7327 (N_7327,N_7209,N_7260);
or U7328 (N_7328,N_7281,N_7276);
and U7329 (N_7329,N_7219,N_7236);
nand U7330 (N_7330,N_7217,N_7250);
xnor U7331 (N_7331,N_7235,N_7227);
and U7332 (N_7332,N_7243,N_7268);
nor U7333 (N_7333,N_7255,N_7294);
nand U7334 (N_7334,N_7237,N_7230);
xor U7335 (N_7335,N_7262,N_7233);
nand U7336 (N_7336,N_7275,N_7286);
xor U7337 (N_7337,N_7287,N_7240);
xnor U7338 (N_7338,N_7258,N_7232);
nor U7339 (N_7339,N_7270,N_7222);
and U7340 (N_7340,N_7249,N_7288);
xor U7341 (N_7341,N_7206,N_7289);
nor U7342 (N_7342,N_7251,N_7256);
or U7343 (N_7343,N_7267,N_7298);
or U7344 (N_7344,N_7214,N_7200);
nor U7345 (N_7345,N_7254,N_7207);
or U7346 (N_7346,N_7223,N_7269);
nand U7347 (N_7347,N_7284,N_7278);
and U7348 (N_7348,N_7248,N_7273);
nor U7349 (N_7349,N_7252,N_7202);
nand U7350 (N_7350,N_7204,N_7241);
xnor U7351 (N_7351,N_7269,N_7202);
nand U7352 (N_7352,N_7233,N_7268);
xor U7353 (N_7353,N_7211,N_7221);
nand U7354 (N_7354,N_7254,N_7274);
xnor U7355 (N_7355,N_7239,N_7256);
nor U7356 (N_7356,N_7233,N_7251);
xnor U7357 (N_7357,N_7282,N_7240);
xnor U7358 (N_7358,N_7234,N_7283);
and U7359 (N_7359,N_7258,N_7245);
xor U7360 (N_7360,N_7291,N_7238);
xor U7361 (N_7361,N_7259,N_7220);
or U7362 (N_7362,N_7259,N_7241);
nor U7363 (N_7363,N_7230,N_7238);
nor U7364 (N_7364,N_7268,N_7262);
nand U7365 (N_7365,N_7259,N_7240);
xor U7366 (N_7366,N_7299,N_7242);
or U7367 (N_7367,N_7250,N_7287);
and U7368 (N_7368,N_7245,N_7296);
or U7369 (N_7369,N_7225,N_7251);
xor U7370 (N_7370,N_7285,N_7256);
nand U7371 (N_7371,N_7243,N_7204);
nand U7372 (N_7372,N_7226,N_7275);
nor U7373 (N_7373,N_7229,N_7208);
or U7374 (N_7374,N_7231,N_7243);
nand U7375 (N_7375,N_7242,N_7247);
nor U7376 (N_7376,N_7248,N_7200);
nor U7377 (N_7377,N_7229,N_7262);
and U7378 (N_7378,N_7262,N_7289);
and U7379 (N_7379,N_7246,N_7260);
nand U7380 (N_7380,N_7242,N_7269);
or U7381 (N_7381,N_7277,N_7228);
xor U7382 (N_7382,N_7264,N_7203);
nor U7383 (N_7383,N_7253,N_7201);
nor U7384 (N_7384,N_7213,N_7246);
nand U7385 (N_7385,N_7251,N_7203);
or U7386 (N_7386,N_7266,N_7296);
xnor U7387 (N_7387,N_7267,N_7250);
or U7388 (N_7388,N_7264,N_7261);
and U7389 (N_7389,N_7269,N_7296);
and U7390 (N_7390,N_7298,N_7278);
and U7391 (N_7391,N_7236,N_7229);
and U7392 (N_7392,N_7282,N_7222);
nand U7393 (N_7393,N_7230,N_7222);
xor U7394 (N_7394,N_7228,N_7291);
or U7395 (N_7395,N_7224,N_7276);
or U7396 (N_7396,N_7223,N_7273);
nor U7397 (N_7397,N_7280,N_7223);
nor U7398 (N_7398,N_7224,N_7265);
nand U7399 (N_7399,N_7230,N_7245);
nor U7400 (N_7400,N_7331,N_7386);
nor U7401 (N_7401,N_7380,N_7322);
xnor U7402 (N_7402,N_7327,N_7345);
or U7403 (N_7403,N_7328,N_7318);
or U7404 (N_7404,N_7377,N_7316);
and U7405 (N_7405,N_7398,N_7301);
xor U7406 (N_7406,N_7361,N_7336);
nand U7407 (N_7407,N_7310,N_7329);
or U7408 (N_7408,N_7325,N_7399);
nand U7409 (N_7409,N_7306,N_7384);
or U7410 (N_7410,N_7346,N_7334);
nor U7411 (N_7411,N_7348,N_7326);
xor U7412 (N_7412,N_7372,N_7341);
and U7413 (N_7413,N_7309,N_7375);
xor U7414 (N_7414,N_7302,N_7353);
xor U7415 (N_7415,N_7330,N_7347);
or U7416 (N_7416,N_7305,N_7396);
and U7417 (N_7417,N_7338,N_7317);
nand U7418 (N_7418,N_7323,N_7314);
nor U7419 (N_7419,N_7324,N_7351);
or U7420 (N_7420,N_7383,N_7382);
nand U7421 (N_7421,N_7392,N_7315);
nor U7422 (N_7422,N_7359,N_7354);
and U7423 (N_7423,N_7387,N_7366);
nor U7424 (N_7424,N_7389,N_7393);
or U7425 (N_7425,N_7394,N_7319);
xnor U7426 (N_7426,N_7357,N_7332);
and U7427 (N_7427,N_7376,N_7312);
and U7428 (N_7428,N_7313,N_7321);
xor U7429 (N_7429,N_7342,N_7349);
nor U7430 (N_7430,N_7369,N_7368);
or U7431 (N_7431,N_7340,N_7355);
and U7432 (N_7432,N_7373,N_7311);
and U7433 (N_7433,N_7320,N_7390);
nor U7434 (N_7434,N_7300,N_7363);
and U7435 (N_7435,N_7362,N_7339);
nor U7436 (N_7436,N_7344,N_7379);
nor U7437 (N_7437,N_7303,N_7395);
xnor U7438 (N_7438,N_7370,N_7352);
and U7439 (N_7439,N_7364,N_7335);
or U7440 (N_7440,N_7356,N_7365);
nor U7441 (N_7441,N_7374,N_7343);
or U7442 (N_7442,N_7333,N_7397);
nand U7443 (N_7443,N_7360,N_7378);
nand U7444 (N_7444,N_7358,N_7350);
nor U7445 (N_7445,N_7388,N_7367);
nor U7446 (N_7446,N_7304,N_7308);
or U7447 (N_7447,N_7391,N_7381);
nand U7448 (N_7448,N_7385,N_7371);
nand U7449 (N_7449,N_7337,N_7307);
nor U7450 (N_7450,N_7338,N_7302);
and U7451 (N_7451,N_7322,N_7381);
nor U7452 (N_7452,N_7315,N_7395);
nor U7453 (N_7453,N_7318,N_7372);
nor U7454 (N_7454,N_7380,N_7330);
nand U7455 (N_7455,N_7373,N_7333);
xor U7456 (N_7456,N_7301,N_7399);
or U7457 (N_7457,N_7322,N_7324);
nand U7458 (N_7458,N_7321,N_7304);
nor U7459 (N_7459,N_7312,N_7365);
xnor U7460 (N_7460,N_7384,N_7304);
nor U7461 (N_7461,N_7367,N_7332);
and U7462 (N_7462,N_7332,N_7335);
xnor U7463 (N_7463,N_7356,N_7320);
or U7464 (N_7464,N_7309,N_7380);
nor U7465 (N_7465,N_7312,N_7394);
xor U7466 (N_7466,N_7337,N_7395);
or U7467 (N_7467,N_7311,N_7352);
nand U7468 (N_7468,N_7324,N_7334);
and U7469 (N_7469,N_7379,N_7332);
or U7470 (N_7470,N_7304,N_7350);
nand U7471 (N_7471,N_7351,N_7388);
or U7472 (N_7472,N_7399,N_7347);
nand U7473 (N_7473,N_7342,N_7321);
and U7474 (N_7474,N_7391,N_7318);
xnor U7475 (N_7475,N_7337,N_7351);
nand U7476 (N_7476,N_7354,N_7399);
or U7477 (N_7477,N_7305,N_7323);
nor U7478 (N_7478,N_7391,N_7369);
or U7479 (N_7479,N_7394,N_7307);
and U7480 (N_7480,N_7344,N_7391);
or U7481 (N_7481,N_7362,N_7369);
xnor U7482 (N_7482,N_7389,N_7352);
and U7483 (N_7483,N_7378,N_7365);
nand U7484 (N_7484,N_7318,N_7377);
nor U7485 (N_7485,N_7392,N_7355);
and U7486 (N_7486,N_7397,N_7357);
xnor U7487 (N_7487,N_7353,N_7334);
nor U7488 (N_7488,N_7348,N_7306);
nand U7489 (N_7489,N_7358,N_7310);
xor U7490 (N_7490,N_7326,N_7322);
xnor U7491 (N_7491,N_7357,N_7346);
and U7492 (N_7492,N_7395,N_7379);
nand U7493 (N_7493,N_7355,N_7308);
xnor U7494 (N_7494,N_7327,N_7310);
and U7495 (N_7495,N_7304,N_7317);
and U7496 (N_7496,N_7363,N_7315);
nor U7497 (N_7497,N_7351,N_7390);
or U7498 (N_7498,N_7385,N_7325);
or U7499 (N_7499,N_7393,N_7303);
and U7500 (N_7500,N_7466,N_7411);
nor U7501 (N_7501,N_7495,N_7476);
or U7502 (N_7502,N_7467,N_7434);
or U7503 (N_7503,N_7456,N_7428);
xor U7504 (N_7504,N_7446,N_7482);
nor U7505 (N_7505,N_7496,N_7481);
nand U7506 (N_7506,N_7477,N_7404);
or U7507 (N_7507,N_7448,N_7405);
nor U7508 (N_7508,N_7490,N_7400);
nand U7509 (N_7509,N_7410,N_7450);
nor U7510 (N_7510,N_7408,N_7461);
and U7511 (N_7511,N_7435,N_7460);
xor U7512 (N_7512,N_7437,N_7449);
nor U7513 (N_7513,N_7420,N_7478);
or U7514 (N_7514,N_7489,N_7484);
and U7515 (N_7515,N_7415,N_7479);
nor U7516 (N_7516,N_7459,N_7473);
nor U7517 (N_7517,N_7421,N_7457);
and U7518 (N_7518,N_7438,N_7417);
and U7519 (N_7519,N_7402,N_7418);
nand U7520 (N_7520,N_7406,N_7469);
nor U7521 (N_7521,N_7431,N_7494);
nand U7522 (N_7522,N_7444,N_7475);
nor U7523 (N_7523,N_7403,N_7430);
nand U7524 (N_7524,N_7474,N_7414);
nor U7525 (N_7525,N_7483,N_7465);
and U7526 (N_7526,N_7470,N_7499);
nor U7527 (N_7527,N_7487,N_7452);
xor U7528 (N_7528,N_7462,N_7425);
or U7529 (N_7529,N_7458,N_7442);
xnor U7530 (N_7530,N_7439,N_7454);
and U7531 (N_7531,N_7485,N_7409);
nor U7532 (N_7532,N_7464,N_7455);
nor U7533 (N_7533,N_7445,N_7429);
nand U7534 (N_7534,N_7413,N_7451);
nand U7535 (N_7535,N_7424,N_7419);
or U7536 (N_7536,N_7471,N_7407);
nand U7537 (N_7537,N_7447,N_7493);
and U7538 (N_7538,N_7443,N_7463);
nand U7539 (N_7539,N_7426,N_7433);
or U7540 (N_7540,N_7472,N_7432);
nor U7541 (N_7541,N_7401,N_7427);
and U7542 (N_7542,N_7491,N_7440);
xnor U7543 (N_7543,N_7436,N_7492);
xnor U7544 (N_7544,N_7468,N_7412);
nand U7545 (N_7545,N_7441,N_7422);
xor U7546 (N_7546,N_7416,N_7486);
or U7547 (N_7547,N_7497,N_7498);
and U7548 (N_7548,N_7480,N_7453);
or U7549 (N_7549,N_7423,N_7488);
or U7550 (N_7550,N_7499,N_7495);
and U7551 (N_7551,N_7485,N_7460);
and U7552 (N_7552,N_7480,N_7432);
xnor U7553 (N_7553,N_7476,N_7418);
nor U7554 (N_7554,N_7458,N_7482);
nor U7555 (N_7555,N_7478,N_7498);
or U7556 (N_7556,N_7482,N_7412);
xnor U7557 (N_7557,N_7431,N_7456);
or U7558 (N_7558,N_7486,N_7457);
or U7559 (N_7559,N_7493,N_7422);
nand U7560 (N_7560,N_7437,N_7422);
nor U7561 (N_7561,N_7457,N_7478);
or U7562 (N_7562,N_7442,N_7468);
or U7563 (N_7563,N_7461,N_7411);
nand U7564 (N_7564,N_7465,N_7436);
xnor U7565 (N_7565,N_7490,N_7482);
or U7566 (N_7566,N_7412,N_7453);
nor U7567 (N_7567,N_7449,N_7460);
or U7568 (N_7568,N_7409,N_7438);
nand U7569 (N_7569,N_7404,N_7444);
nand U7570 (N_7570,N_7463,N_7484);
nor U7571 (N_7571,N_7418,N_7414);
and U7572 (N_7572,N_7464,N_7470);
or U7573 (N_7573,N_7488,N_7461);
nor U7574 (N_7574,N_7494,N_7412);
nor U7575 (N_7575,N_7435,N_7431);
nor U7576 (N_7576,N_7464,N_7400);
nand U7577 (N_7577,N_7467,N_7460);
or U7578 (N_7578,N_7439,N_7417);
nand U7579 (N_7579,N_7471,N_7423);
nor U7580 (N_7580,N_7422,N_7489);
and U7581 (N_7581,N_7458,N_7464);
or U7582 (N_7582,N_7430,N_7422);
nand U7583 (N_7583,N_7455,N_7400);
and U7584 (N_7584,N_7493,N_7441);
or U7585 (N_7585,N_7459,N_7485);
nand U7586 (N_7586,N_7488,N_7464);
and U7587 (N_7587,N_7440,N_7426);
and U7588 (N_7588,N_7479,N_7451);
nand U7589 (N_7589,N_7496,N_7455);
xnor U7590 (N_7590,N_7423,N_7438);
and U7591 (N_7591,N_7474,N_7401);
or U7592 (N_7592,N_7439,N_7402);
nand U7593 (N_7593,N_7494,N_7429);
xor U7594 (N_7594,N_7475,N_7498);
xor U7595 (N_7595,N_7444,N_7493);
nor U7596 (N_7596,N_7451,N_7417);
or U7597 (N_7597,N_7409,N_7420);
xnor U7598 (N_7598,N_7416,N_7494);
nor U7599 (N_7599,N_7427,N_7453);
or U7600 (N_7600,N_7542,N_7580);
and U7601 (N_7601,N_7559,N_7560);
and U7602 (N_7602,N_7592,N_7596);
or U7603 (N_7603,N_7576,N_7584);
xnor U7604 (N_7604,N_7507,N_7543);
xor U7605 (N_7605,N_7572,N_7546);
xor U7606 (N_7606,N_7531,N_7519);
and U7607 (N_7607,N_7553,N_7574);
nand U7608 (N_7608,N_7561,N_7594);
xor U7609 (N_7609,N_7586,N_7565);
or U7610 (N_7610,N_7551,N_7547);
xor U7611 (N_7611,N_7571,N_7532);
and U7612 (N_7612,N_7583,N_7522);
or U7613 (N_7613,N_7511,N_7529);
nor U7614 (N_7614,N_7539,N_7570);
xnor U7615 (N_7615,N_7587,N_7503);
and U7616 (N_7616,N_7521,N_7536);
xor U7617 (N_7617,N_7534,N_7556);
nor U7618 (N_7618,N_7506,N_7504);
or U7619 (N_7619,N_7567,N_7528);
nor U7620 (N_7620,N_7520,N_7598);
nand U7621 (N_7621,N_7518,N_7558);
and U7622 (N_7622,N_7515,N_7509);
nand U7623 (N_7623,N_7595,N_7544);
or U7624 (N_7624,N_7505,N_7590);
nor U7625 (N_7625,N_7554,N_7523);
nand U7626 (N_7626,N_7568,N_7538);
or U7627 (N_7627,N_7575,N_7501);
xor U7628 (N_7628,N_7564,N_7526);
nor U7629 (N_7629,N_7530,N_7540);
nand U7630 (N_7630,N_7566,N_7527);
nand U7631 (N_7631,N_7557,N_7585);
nor U7632 (N_7632,N_7512,N_7502);
nand U7633 (N_7633,N_7545,N_7577);
nand U7634 (N_7634,N_7513,N_7569);
xnor U7635 (N_7635,N_7578,N_7550);
nor U7636 (N_7636,N_7581,N_7537);
nand U7637 (N_7637,N_7533,N_7517);
nand U7638 (N_7638,N_7562,N_7510);
and U7639 (N_7639,N_7588,N_7591);
and U7640 (N_7640,N_7541,N_7589);
nor U7641 (N_7641,N_7555,N_7597);
nand U7642 (N_7642,N_7593,N_7535);
or U7643 (N_7643,N_7524,N_7500);
nand U7644 (N_7644,N_7525,N_7514);
nor U7645 (N_7645,N_7549,N_7573);
and U7646 (N_7646,N_7548,N_7579);
nand U7647 (N_7647,N_7516,N_7563);
or U7648 (N_7648,N_7582,N_7508);
or U7649 (N_7649,N_7599,N_7552);
and U7650 (N_7650,N_7522,N_7504);
xor U7651 (N_7651,N_7597,N_7537);
xnor U7652 (N_7652,N_7519,N_7592);
nand U7653 (N_7653,N_7513,N_7532);
xor U7654 (N_7654,N_7536,N_7511);
or U7655 (N_7655,N_7502,N_7555);
or U7656 (N_7656,N_7535,N_7511);
or U7657 (N_7657,N_7587,N_7596);
nor U7658 (N_7658,N_7531,N_7533);
nand U7659 (N_7659,N_7534,N_7539);
and U7660 (N_7660,N_7590,N_7521);
nor U7661 (N_7661,N_7570,N_7587);
nor U7662 (N_7662,N_7577,N_7592);
and U7663 (N_7663,N_7535,N_7540);
xor U7664 (N_7664,N_7519,N_7507);
or U7665 (N_7665,N_7568,N_7527);
and U7666 (N_7666,N_7537,N_7550);
nand U7667 (N_7667,N_7547,N_7546);
nor U7668 (N_7668,N_7509,N_7594);
nand U7669 (N_7669,N_7500,N_7589);
nor U7670 (N_7670,N_7592,N_7564);
nor U7671 (N_7671,N_7542,N_7511);
and U7672 (N_7672,N_7589,N_7560);
or U7673 (N_7673,N_7583,N_7532);
or U7674 (N_7674,N_7537,N_7562);
nand U7675 (N_7675,N_7531,N_7565);
and U7676 (N_7676,N_7561,N_7520);
nor U7677 (N_7677,N_7554,N_7537);
and U7678 (N_7678,N_7592,N_7526);
or U7679 (N_7679,N_7546,N_7515);
nand U7680 (N_7680,N_7579,N_7595);
and U7681 (N_7681,N_7541,N_7553);
nand U7682 (N_7682,N_7522,N_7523);
and U7683 (N_7683,N_7583,N_7536);
and U7684 (N_7684,N_7510,N_7545);
and U7685 (N_7685,N_7521,N_7517);
or U7686 (N_7686,N_7500,N_7501);
and U7687 (N_7687,N_7590,N_7589);
or U7688 (N_7688,N_7558,N_7544);
or U7689 (N_7689,N_7559,N_7517);
nor U7690 (N_7690,N_7526,N_7519);
and U7691 (N_7691,N_7547,N_7530);
and U7692 (N_7692,N_7503,N_7586);
xor U7693 (N_7693,N_7538,N_7512);
or U7694 (N_7694,N_7515,N_7591);
xnor U7695 (N_7695,N_7524,N_7508);
or U7696 (N_7696,N_7542,N_7561);
nor U7697 (N_7697,N_7538,N_7574);
nor U7698 (N_7698,N_7530,N_7533);
nor U7699 (N_7699,N_7561,N_7574);
or U7700 (N_7700,N_7673,N_7638);
nand U7701 (N_7701,N_7618,N_7625);
nand U7702 (N_7702,N_7664,N_7657);
nand U7703 (N_7703,N_7674,N_7659);
and U7704 (N_7704,N_7602,N_7608);
nor U7705 (N_7705,N_7653,N_7620);
and U7706 (N_7706,N_7611,N_7637);
and U7707 (N_7707,N_7670,N_7656);
nand U7708 (N_7708,N_7683,N_7684);
nor U7709 (N_7709,N_7612,N_7619);
nor U7710 (N_7710,N_7676,N_7689);
and U7711 (N_7711,N_7627,N_7650);
and U7712 (N_7712,N_7606,N_7698);
nor U7713 (N_7713,N_7636,N_7681);
nand U7714 (N_7714,N_7661,N_7632);
nor U7715 (N_7715,N_7623,N_7658);
and U7716 (N_7716,N_7668,N_7691);
xnor U7717 (N_7717,N_7624,N_7639);
xor U7718 (N_7718,N_7693,N_7617);
xnor U7719 (N_7719,N_7640,N_7692);
nand U7720 (N_7720,N_7616,N_7685);
xnor U7721 (N_7721,N_7682,N_7671);
nor U7722 (N_7722,N_7631,N_7669);
nand U7723 (N_7723,N_7672,N_7687);
and U7724 (N_7724,N_7678,N_7699);
or U7725 (N_7725,N_7622,N_7614);
nand U7726 (N_7726,N_7635,N_7628);
or U7727 (N_7727,N_7626,N_7690);
xor U7728 (N_7728,N_7679,N_7696);
and U7729 (N_7729,N_7642,N_7694);
nand U7730 (N_7730,N_7607,N_7662);
nor U7731 (N_7731,N_7645,N_7605);
and U7732 (N_7732,N_7641,N_7649);
and U7733 (N_7733,N_7677,N_7630);
nor U7734 (N_7734,N_7610,N_7655);
or U7735 (N_7735,N_7697,N_7643);
or U7736 (N_7736,N_7654,N_7647);
and U7737 (N_7737,N_7660,N_7646);
nand U7738 (N_7738,N_7621,N_7666);
or U7739 (N_7739,N_7613,N_7601);
or U7740 (N_7740,N_7686,N_7680);
or U7741 (N_7741,N_7663,N_7634);
nor U7742 (N_7742,N_7644,N_7665);
nand U7743 (N_7743,N_7603,N_7648);
nor U7744 (N_7744,N_7695,N_7688);
nand U7745 (N_7745,N_7600,N_7652);
nand U7746 (N_7746,N_7633,N_7629);
nor U7747 (N_7747,N_7651,N_7667);
nor U7748 (N_7748,N_7604,N_7615);
nor U7749 (N_7749,N_7675,N_7609);
or U7750 (N_7750,N_7617,N_7681);
nand U7751 (N_7751,N_7619,N_7694);
nor U7752 (N_7752,N_7677,N_7668);
or U7753 (N_7753,N_7697,N_7611);
xor U7754 (N_7754,N_7649,N_7650);
nand U7755 (N_7755,N_7692,N_7602);
xor U7756 (N_7756,N_7665,N_7606);
and U7757 (N_7757,N_7690,N_7699);
nand U7758 (N_7758,N_7663,N_7697);
xor U7759 (N_7759,N_7677,N_7687);
or U7760 (N_7760,N_7659,N_7670);
and U7761 (N_7761,N_7694,N_7621);
xnor U7762 (N_7762,N_7656,N_7678);
or U7763 (N_7763,N_7654,N_7651);
and U7764 (N_7764,N_7640,N_7614);
xnor U7765 (N_7765,N_7689,N_7614);
or U7766 (N_7766,N_7633,N_7602);
xor U7767 (N_7767,N_7604,N_7641);
and U7768 (N_7768,N_7696,N_7690);
or U7769 (N_7769,N_7664,N_7641);
xnor U7770 (N_7770,N_7655,N_7692);
or U7771 (N_7771,N_7613,N_7699);
nand U7772 (N_7772,N_7618,N_7640);
and U7773 (N_7773,N_7603,N_7694);
nor U7774 (N_7774,N_7602,N_7622);
nor U7775 (N_7775,N_7673,N_7687);
xor U7776 (N_7776,N_7640,N_7657);
xor U7777 (N_7777,N_7640,N_7619);
and U7778 (N_7778,N_7600,N_7648);
and U7779 (N_7779,N_7688,N_7604);
nor U7780 (N_7780,N_7657,N_7611);
nor U7781 (N_7781,N_7648,N_7608);
xnor U7782 (N_7782,N_7615,N_7661);
and U7783 (N_7783,N_7640,N_7602);
nand U7784 (N_7784,N_7665,N_7696);
nand U7785 (N_7785,N_7683,N_7638);
or U7786 (N_7786,N_7645,N_7639);
nor U7787 (N_7787,N_7691,N_7638);
xor U7788 (N_7788,N_7677,N_7617);
and U7789 (N_7789,N_7651,N_7604);
or U7790 (N_7790,N_7699,N_7676);
nor U7791 (N_7791,N_7617,N_7674);
xnor U7792 (N_7792,N_7675,N_7673);
nand U7793 (N_7793,N_7613,N_7623);
nor U7794 (N_7794,N_7619,N_7699);
nand U7795 (N_7795,N_7618,N_7650);
nand U7796 (N_7796,N_7667,N_7600);
xor U7797 (N_7797,N_7644,N_7686);
and U7798 (N_7798,N_7624,N_7609);
and U7799 (N_7799,N_7611,N_7642);
or U7800 (N_7800,N_7746,N_7785);
or U7801 (N_7801,N_7736,N_7710);
nor U7802 (N_7802,N_7707,N_7730);
nand U7803 (N_7803,N_7720,N_7793);
nand U7804 (N_7804,N_7709,N_7773);
and U7805 (N_7805,N_7788,N_7741);
xor U7806 (N_7806,N_7711,N_7783);
and U7807 (N_7807,N_7787,N_7708);
xnor U7808 (N_7808,N_7705,N_7747);
xor U7809 (N_7809,N_7791,N_7799);
and U7810 (N_7810,N_7718,N_7731);
xnor U7811 (N_7811,N_7740,N_7797);
nor U7812 (N_7812,N_7766,N_7722);
and U7813 (N_7813,N_7701,N_7742);
nor U7814 (N_7814,N_7752,N_7702);
nand U7815 (N_7815,N_7756,N_7732);
nand U7816 (N_7816,N_7703,N_7751);
nor U7817 (N_7817,N_7765,N_7761);
nor U7818 (N_7818,N_7776,N_7760);
or U7819 (N_7819,N_7735,N_7743);
nand U7820 (N_7820,N_7777,N_7771);
xor U7821 (N_7821,N_7734,N_7774);
nand U7822 (N_7822,N_7769,N_7784);
xor U7823 (N_7823,N_7755,N_7749);
or U7824 (N_7824,N_7719,N_7700);
nand U7825 (N_7825,N_7779,N_7759);
nor U7826 (N_7826,N_7714,N_7750);
or U7827 (N_7827,N_7717,N_7762);
and U7828 (N_7828,N_7728,N_7782);
nor U7829 (N_7829,N_7794,N_7754);
nor U7830 (N_7830,N_7712,N_7772);
nand U7831 (N_7831,N_7796,N_7723);
nor U7832 (N_7832,N_7738,N_7715);
nand U7833 (N_7833,N_7745,N_7770);
xor U7834 (N_7834,N_7781,N_7763);
nand U7835 (N_7835,N_7706,N_7780);
nand U7836 (N_7836,N_7753,N_7768);
nand U7837 (N_7837,N_7739,N_7786);
and U7838 (N_7838,N_7727,N_7733);
and U7839 (N_7839,N_7790,N_7758);
or U7840 (N_7840,N_7789,N_7798);
and U7841 (N_7841,N_7725,N_7767);
or U7842 (N_7842,N_7721,N_7792);
nor U7843 (N_7843,N_7764,N_7729);
nor U7844 (N_7844,N_7778,N_7775);
xor U7845 (N_7845,N_7716,N_7704);
xor U7846 (N_7846,N_7724,N_7795);
nor U7847 (N_7847,N_7757,N_7737);
and U7848 (N_7848,N_7748,N_7713);
xor U7849 (N_7849,N_7744,N_7726);
nor U7850 (N_7850,N_7794,N_7750);
xor U7851 (N_7851,N_7722,N_7764);
nand U7852 (N_7852,N_7765,N_7724);
xor U7853 (N_7853,N_7769,N_7741);
nand U7854 (N_7854,N_7712,N_7786);
nand U7855 (N_7855,N_7792,N_7716);
xor U7856 (N_7856,N_7760,N_7772);
nor U7857 (N_7857,N_7714,N_7788);
xor U7858 (N_7858,N_7749,N_7774);
or U7859 (N_7859,N_7719,N_7768);
and U7860 (N_7860,N_7724,N_7740);
and U7861 (N_7861,N_7778,N_7707);
nor U7862 (N_7862,N_7744,N_7754);
nor U7863 (N_7863,N_7748,N_7792);
xor U7864 (N_7864,N_7721,N_7790);
xnor U7865 (N_7865,N_7725,N_7713);
nand U7866 (N_7866,N_7710,N_7745);
nor U7867 (N_7867,N_7763,N_7707);
nor U7868 (N_7868,N_7729,N_7777);
nor U7869 (N_7869,N_7757,N_7718);
nor U7870 (N_7870,N_7717,N_7708);
or U7871 (N_7871,N_7744,N_7771);
xnor U7872 (N_7872,N_7796,N_7765);
xor U7873 (N_7873,N_7740,N_7711);
and U7874 (N_7874,N_7736,N_7712);
xnor U7875 (N_7875,N_7700,N_7799);
nand U7876 (N_7876,N_7793,N_7708);
xnor U7877 (N_7877,N_7771,N_7769);
or U7878 (N_7878,N_7750,N_7748);
nand U7879 (N_7879,N_7783,N_7738);
xor U7880 (N_7880,N_7704,N_7756);
nand U7881 (N_7881,N_7719,N_7743);
xnor U7882 (N_7882,N_7750,N_7732);
and U7883 (N_7883,N_7768,N_7714);
or U7884 (N_7884,N_7751,N_7773);
xor U7885 (N_7885,N_7774,N_7733);
nand U7886 (N_7886,N_7796,N_7734);
nor U7887 (N_7887,N_7767,N_7726);
xnor U7888 (N_7888,N_7749,N_7747);
nand U7889 (N_7889,N_7734,N_7745);
nand U7890 (N_7890,N_7774,N_7761);
nor U7891 (N_7891,N_7741,N_7765);
and U7892 (N_7892,N_7714,N_7739);
nand U7893 (N_7893,N_7740,N_7735);
xor U7894 (N_7894,N_7739,N_7754);
xnor U7895 (N_7895,N_7717,N_7707);
nor U7896 (N_7896,N_7737,N_7773);
nand U7897 (N_7897,N_7766,N_7745);
nand U7898 (N_7898,N_7755,N_7715);
nand U7899 (N_7899,N_7784,N_7773);
xnor U7900 (N_7900,N_7810,N_7857);
or U7901 (N_7901,N_7813,N_7853);
nor U7902 (N_7902,N_7849,N_7879);
nand U7903 (N_7903,N_7873,N_7837);
xor U7904 (N_7904,N_7891,N_7854);
xnor U7905 (N_7905,N_7882,N_7884);
nand U7906 (N_7906,N_7818,N_7869);
and U7907 (N_7907,N_7819,N_7823);
nand U7908 (N_7908,N_7824,N_7880);
xnor U7909 (N_7909,N_7840,N_7886);
or U7910 (N_7910,N_7826,N_7856);
or U7911 (N_7911,N_7883,N_7808);
nand U7912 (N_7912,N_7841,N_7865);
nand U7913 (N_7913,N_7862,N_7843);
or U7914 (N_7914,N_7838,N_7852);
xnor U7915 (N_7915,N_7892,N_7821);
xnor U7916 (N_7916,N_7888,N_7814);
or U7917 (N_7917,N_7801,N_7805);
and U7918 (N_7918,N_7887,N_7851);
nand U7919 (N_7919,N_7815,N_7831);
xor U7920 (N_7920,N_7816,N_7890);
xor U7921 (N_7921,N_7812,N_7800);
nor U7922 (N_7922,N_7842,N_7874);
or U7923 (N_7923,N_7859,N_7829);
or U7924 (N_7924,N_7822,N_7825);
nor U7925 (N_7925,N_7834,N_7802);
xnor U7926 (N_7926,N_7827,N_7809);
or U7927 (N_7927,N_7863,N_7885);
and U7928 (N_7928,N_7868,N_7861);
xnor U7929 (N_7929,N_7846,N_7807);
and U7930 (N_7930,N_7847,N_7878);
nand U7931 (N_7931,N_7835,N_7806);
nor U7932 (N_7932,N_7844,N_7817);
nand U7933 (N_7933,N_7867,N_7875);
or U7934 (N_7934,N_7830,N_7897);
nand U7935 (N_7935,N_7832,N_7804);
or U7936 (N_7936,N_7855,N_7820);
nand U7937 (N_7937,N_7866,N_7877);
nand U7938 (N_7938,N_7871,N_7828);
xor U7939 (N_7939,N_7848,N_7858);
xor U7940 (N_7940,N_7850,N_7860);
or U7941 (N_7941,N_7811,N_7803);
nand U7942 (N_7942,N_7845,N_7896);
and U7943 (N_7943,N_7836,N_7889);
or U7944 (N_7944,N_7864,N_7899);
nand U7945 (N_7945,N_7870,N_7839);
or U7946 (N_7946,N_7876,N_7872);
or U7947 (N_7947,N_7893,N_7895);
xor U7948 (N_7948,N_7881,N_7898);
xnor U7949 (N_7949,N_7833,N_7894);
nor U7950 (N_7950,N_7839,N_7882);
or U7951 (N_7951,N_7897,N_7838);
or U7952 (N_7952,N_7824,N_7895);
and U7953 (N_7953,N_7879,N_7883);
xnor U7954 (N_7954,N_7805,N_7854);
and U7955 (N_7955,N_7847,N_7881);
and U7956 (N_7956,N_7860,N_7818);
nand U7957 (N_7957,N_7882,N_7815);
and U7958 (N_7958,N_7860,N_7838);
and U7959 (N_7959,N_7871,N_7806);
or U7960 (N_7960,N_7872,N_7819);
xor U7961 (N_7961,N_7860,N_7869);
nor U7962 (N_7962,N_7854,N_7819);
or U7963 (N_7963,N_7876,N_7864);
nor U7964 (N_7964,N_7892,N_7801);
nor U7965 (N_7965,N_7809,N_7845);
or U7966 (N_7966,N_7826,N_7834);
nand U7967 (N_7967,N_7846,N_7840);
nor U7968 (N_7968,N_7883,N_7822);
and U7969 (N_7969,N_7897,N_7870);
nand U7970 (N_7970,N_7833,N_7868);
nand U7971 (N_7971,N_7858,N_7893);
nor U7972 (N_7972,N_7890,N_7874);
or U7973 (N_7973,N_7899,N_7821);
or U7974 (N_7974,N_7862,N_7832);
and U7975 (N_7975,N_7821,N_7835);
nor U7976 (N_7976,N_7851,N_7863);
and U7977 (N_7977,N_7878,N_7835);
xor U7978 (N_7978,N_7894,N_7873);
xor U7979 (N_7979,N_7839,N_7858);
xnor U7980 (N_7980,N_7842,N_7876);
nor U7981 (N_7981,N_7854,N_7865);
or U7982 (N_7982,N_7804,N_7852);
nand U7983 (N_7983,N_7839,N_7807);
xor U7984 (N_7984,N_7870,N_7824);
nand U7985 (N_7985,N_7884,N_7890);
or U7986 (N_7986,N_7862,N_7892);
xor U7987 (N_7987,N_7893,N_7847);
xor U7988 (N_7988,N_7877,N_7858);
nor U7989 (N_7989,N_7878,N_7825);
and U7990 (N_7990,N_7813,N_7849);
nand U7991 (N_7991,N_7895,N_7829);
or U7992 (N_7992,N_7878,N_7823);
nand U7993 (N_7993,N_7812,N_7803);
or U7994 (N_7994,N_7813,N_7810);
or U7995 (N_7995,N_7848,N_7831);
xnor U7996 (N_7996,N_7812,N_7850);
xor U7997 (N_7997,N_7881,N_7808);
nor U7998 (N_7998,N_7813,N_7811);
nor U7999 (N_7999,N_7895,N_7888);
and U8000 (N_8000,N_7951,N_7902);
or U8001 (N_8001,N_7905,N_7988);
xnor U8002 (N_8002,N_7939,N_7904);
nor U8003 (N_8003,N_7914,N_7907);
nor U8004 (N_8004,N_7969,N_7986);
or U8005 (N_8005,N_7930,N_7979);
nor U8006 (N_8006,N_7948,N_7924);
nor U8007 (N_8007,N_7961,N_7974);
or U8008 (N_8008,N_7959,N_7998);
nor U8009 (N_8009,N_7926,N_7993);
or U8010 (N_8010,N_7970,N_7923);
nor U8011 (N_8011,N_7965,N_7921);
and U8012 (N_8012,N_7908,N_7967);
nand U8013 (N_8013,N_7981,N_7937);
nor U8014 (N_8014,N_7972,N_7940);
nor U8015 (N_8015,N_7991,N_7945);
nor U8016 (N_8016,N_7934,N_7996);
nor U8017 (N_8017,N_7973,N_7913);
xor U8018 (N_8018,N_7947,N_7915);
xor U8019 (N_8019,N_7960,N_7971);
nor U8020 (N_8020,N_7955,N_7916);
xor U8021 (N_8021,N_7964,N_7912);
xnor U8022 (N_8022,N_7976,N_7978);
and U8023 (N_8023,N_7929,N_7950);
xnor U8024 (N_8024,N_7963,N_7935);
nor U8025 (N_8025,N_7906,N_7966);
xor U8026 (N_8026,N_7931,N_7990);
nor U8027 (N_8027,N_7941,N_7992);
or U8028 (N_8028,N_7933,N_7909);
and U8029 (N_8029,N_7900,N_7954);
xor U8030 (N_8030,N_7980,N_7910);
and U8031 (N_8031,N_7958,N_7953);
or U8032 (N_8032,N_7995,N_7922);
nand U8033 (N_8033,N_7927,N_7928);
nor U8034 (N_8034,N_7985,N_7903);
nor U8035 (N_8035,N_7943,N_7962);
or U8036 (N_8036,N_7982,N_7944);
nand U8037 (N_8037,N_7949,N_7956);
xor U8038 (N_8038,N_7987,N_7968);
xor U8039 (N_8039,N_7920,N_7957);
and U8040 (N_8040,N_7917,N_7919);
nor U8041 (N_8041,N_7983,N_7925);
and U8042 (N_8042,N_7938,N_7911);
xor U8043 (N_8043,N_7997,N_7936);
nand U8044 (N_8044,N_7932,N_7942);
nand U8045 (N_8045,N_7994,N_7977);
or U8046 (N_8046,N_7946,N_7999);
and U8047 (N_8047,N_7989,N_7952);
or U8048 (N_8048,N_7984,N_7901);
and U8049 (N_8049,N_7975,N_7918);
xnor U8050 (N_8050,N_7953,N_7970);
nor U8051 (N_8051,N_7946,N_7961);
and U8052 (N_8052,N_7948,N_7919);
nand U8053 (N_8053,N_7942,N_7934);
and U8054 (N_8054,N_7941,N_7922);
nand U8055 (N_8055,N_7907,N_7937);
nand U8056 (N_8056,N_7965,N_7928);
and U8057 (N_8057,N_7936,N_7970);
nor U8058 (N_8058,N_7984,N_7956);
or U8059 (N_8059,N_7999,N_7924);
or U8060 (N_8060,N_7921,N_7938);
and U8061 (N_8061,N_7951,N_7940);
xor U8062 (N_8062,N_7900,N_7950);
nand U8063 (N_8063,N_7962,N_7904);
and U8064 (N_8064,N_7935,N_7919);
xnor U8065 (N_8065,N_7953,N_7966);
xnor U8066 (N_8066,N_7946,N_7975);
nand U8067 (N_8067,N_7946,N_7907);
xnor U8068 (N_8068,N_7997,N_7910);
or U8069 (N_8069,N_7988,N_7969);
nand U8070 (N_8070,N_7918,N_7977);
nor U8071 (N_8071,N_7909,N_7944);
and U8072 (N_8072,N_7994,N_7931);
or U8073 (N_8073,N_7903,N_7904);
and U8074 (N_8074,N_7956,N_7996);
or U8075 (N_8075,N_7966,N_7920);
nand U8076 (N_8076,N_7994,N_7998);
or U8077 (N_8077,N_7993,N_7997);
or U8078 (N_8078,N_7964,N_7988);
nor U8079 (N_8079,N_7973,N_7991);
nor U8080 (N_8080,N_7973,N_7951);
nand U8081 (N_8081,N_7968,N_7941);
and U8082 (N_8082,N_7976,N_7974);
nor U8083 (N_8083,N_7954,N_7972);
nor U8084 (N_8084,N_7988,N_7957);
xnor U8085 (N_8085,N_7943,N_7984);
xor U8086 (N_8086,N_7929,N_7982);
or U8087 (N_8087,N_7911,N_7982);
xnor U8088 (N_8088,N_7924,N_7961);
and U8089 (N_8089,N_7954,N_7955);
or U8090 (N_8090,N_7929,N_7934);
nand U8091 (N_8091,N_7913,N_7914);
xor U8092 (N_8092,N_7940,N_7937);
xor U8093 (N_8093,N_7994,N_7922);
nand U8094 (N_8094,N_7909,N_7931);
or U8095 (N_8095,N_7935,N_7966);
and U8096 (N_8096,N_7906,N_7901);
nand U8097 (N_8097,N_7972,N_7932);
nand U8098 (N_8098,N_7906,N_7997);
nand U8099 (N_8099,N_7986,N_7998);
nand U8100 (N_8100,N_8057,N_8013);
nand U8101 (N_8101,N_8045,N_8083);
xnor U8102 (N_8102,N_8073,N_8078);
nor U8103 (N_8103,N_8038,N_8006);
or U8104 (N_8104,N_8070,N_8026);
nand U8105 (N_8105,N_8061,N_8022);
nor U8106 (N_8106,N_8003,N_8032);
xor U8107 (N_8107,N_8037,N_8067);
or U8108 (N_8108,N_8036,N_8018);
nand U8109 (N_8109,N_8058,N_8048);
xnor U8110 (N_8110,N_8056,N_8097);
or U8111 (N_8111,N_8088,N_8033);
xnor U8112 (N_8112,N_8077,N_8091);
and U8113 (N_8113,N_8095,N_8046);
nor U8114 (N_8114,N_8093,N_8023);
xnor U8115 (N_8115,N_8051,N_8011);
nor U8116 (N_8116,N_8065,N_8099);
nor U8117 (N_8117,N_8063,N_8008);
nor U8118 (N_8118,N_8081,N_8020);
xor U8119 (N_8119,N_8047,N_8071);
or U8120 (N_8120,N_8085,N_8090);
xnor U8121 (N_8121,N_8025,N_8080);
xnor U8122 (N_8122,N_8005,N_8086);
nor U8123 (N_8123,N_8010,N_8007);
nor U8124 (N_8124,N_8042,N_8012);
nand U8125 (N_8125,N_8060,N_8072);
nor U8126 (N_8126,N_8092,N_8054);
nand U8127 (N_8127,N_8049,N_8094);
or U8128 (N_8128,N_8015,N_8076);
nand U8129 (N_8129,N_8084,N_8004);
or U8130 (N_8130,N_8028,N_8027);
and U8131 (N_8131,N_8064,N_8021);
nand U8132 (N_8132,N_8089,N_8096);
or U8133 (N_8133,N_8016,N_8030);
nand U8134 (N_8134,N_8002,N_8087);
or U8135 (N_8135,N_8040,N_8014);
xor U8136 (N_8136,N_8052,N_8000);
xnor U8137 (N_8137,N_8039,N_8009);
xnor U8138 (N_8138,N_8069,N_8034);
xnor U8139 (N_8139,N_8082,N_8019);
xor U8140 (N_8140,N_8059,N_8043);
and U8141 (N_8141,N_8079,N_8031);
or U8142 (N_8142,N_8066,N_8041);
nand U8143 (N_8143,N_8055,N_8098);
nand U8144 (N_8144,N_8001,N_8062);
nand U8145 (N_8145,N_8068,N_8053);
nor U8146 (N_8146,N_8050,N_8017);
or U8147 (N_8147,N_8044,N_8075);
nand U8148 (N_8148,N_8074,N_8035);
xor U8149 (N_8149,N_8024,N_8029);
nor U8150 (N_8150,N_8096,N_8021);
nor U8151 (N_8151,N_8062,N_8038);
xor U8152 (N_8152,N_8028,N_8047);
or U8153 (N_8153,N_8045,N_8098);
nor U8154 (N_8154,N_8059,N_8091);
and U8155 (N_8155,N_8019,N_8003);
xnor U8156 (N_8156,N_8015,N_8086);
xor U8157 (N_8157,N_8012,N_8061);
xnor U8158 (N_8158,N_8099,N_8002);
nor U8159 (N_8159,N_8063,N_8010);
and U8160 (N_8160,N_8073,N_8017);
or U8161 (N_8161,N_8082,N_8012);
and U8162 (N_8162,N_8004,N_8039);
nor U8163 (N_8163,N_8008,N_8097);
nand U8164 (N_8164,N_8049,N_8034);
xor U8165 (N_8165,N_8094,N_8077);
nor U8166 (N_8166,N_8055,N_8043);
nand U8167 (N_8167,N_8070,N_8087);
nor U8168 (N_8168,N_8088,N_8051);
and U8169 (N_8169,N_8010,N_8001);
nand U8170 (N_8170,N_8019,N_8055);
nand U8171 (N_8171,N_8000,N_8010);
nand U8172 (N_8172,N_8046,N_8096);
nand U8173 (N_8173,N_8077,N_8097);
xnor U8174 (N_8174,N_8053,N_8013);
xor U8175 (N_8175,N_8055,N_8075);
and U8176 (N_8176,N_8047,N_8025);
xnor U8177 (N_8177,N_8002,N_8059);
and U8178 (N_8178,N_8083,N_8035);
nand U8179 (N_8179,N_8023,N_8098);
xnor U8180 (N_8180,N_8074,N_8050);
and U8181 (N_8181,N_8003,N_8051);
nand U8182 (N_8182,N_8076,N_8012);
nand U8183 (N_8183,N_8006,N_8080);
nor U8184 (N_8184,N_8064,N_8090);
and U8185 (N_8185,N_8072,N_8034);
nor U8186 (N_8186,N_8089,N_8006);
xnor U8187 (N_8187,N_8034,N_8050);
xor U8188 (N_8188,N_8038,N_8066);
or U8189 (N_8189,N_8088,N_8023);
and U8190 (N_8190,N_8016,N_8082);
and U8191 (N_8191,N_8061,N_8025);
or U8192 (N_8192,N_8018,N_8043);
nand U8193 (N_8193,N_8049,N_8086);
nor U8194 (N_8194,N_8054,N_8026);
nor U8195 (N_8195,N_8041,N_8048);
and U8196 (N_8196,N_8029,N_8051);
nand U8197 (N_8197,N_8014,N_8027);
or U8198 (N_8198,N_8083,N_8056);
nand U8199 (N_8199,N_8046,N_8007);
nand U8200 (N_8200,N_8100,N_8156);
nor U8201 (N_8201,N_8130,N_8119);
or U8202 (N_8202,N_8122,N_8171);
nor U8203 (N_8203,N_8142,N_8188);
or U8204 (N_8204,N_8179,N_8150);
xnor U8205 (N_8205,N_8104,N_8165);
and U8206 (N_8206,N_8185,N_8106);
and U8207 (N_8207,N_8153,N_8129);
and U8208 (N_8208,N_8161,N_8180);
or U8209 (N_8209,N_8102,N_8196);
and U8210 (N_8210,N_8191,N_8136);
xnor U8211 (N_8211,N_8169,N_8174);
or U8212 (N_8212,N_8110,N_8157);
xnor U8213 (N_8213,N_8141,N_8139);
nor U8214 (N_8214,N_8175,N_8197);
or U8215 (N_8215,N_8137,N_8101);
or U8216 (N_8216,N_8164,N_8109);
and U8217 (N_8217,N_8172,N_8155);
nand U8218 (N_8218,N_8194,N_8115);
xor U8219 (N_8219,N_8107,N_8151);
nor U8220 (N_8220,N_8138,N_8168);
and U8221 (N_8221,N_8114,N_8121);
and U8222 (N_8222,N_8118,N_8144);
xnor U8223 (N_8223,N_8170,N_8167);
and U8224 (N_8224,N_8123,N_8183);
or U8225 (N_8225,N_8103,N_8108);
nand U8226 (N_8226,N_8124,N_8113);
and U8227 (N_8227,N_8173,N_8135);
and U8228 (N_8228,N_8145,N_8178);
and U8229 (N_8229,N_8176,N_8186);
nand U8230 (N_8230,N_8190,N_8187);
and U8231 (N_8231,N_8112,N_8148);
nor U8232 (N_8232,N_8177,N_8162);
nand U8233 (N_8233,N_8143,N_8126);
xnor U8234 (N_8234,N_8128,N_8111);
xor U8235 (N_8235,N_8152,N_8163);
nor U8236 (N_8236,N_8182,N_8193);
nand U8237 (N_8237,N_8134,N_8158);
xor U8238 (N_8238,N_8189,N_8146);
or U8239 (N_8239,N_8149,N_8105);
xnor U8240 (N_8240,N_8154,N_8160);
nor U8241 (N_8241,N_8127,N_8131);
xnor U8242 (N_8242,N_8132,N_8166);
nand U8243 (N_8243,N_8184,N_8147);
or U8244 (N_8244,N_8140,N_8199);
nand U8245 (N_8245,N_8116,N_8120);
or U8246 (N_8246,N_8159,N_8198);
or U8247 (N_8247,N_8133,N_8192);
nand U8248 (N_8248,N_8181,N_8195);
or U8249 (N_8249,N_8125,N_8117);
nor U8250 (N_8250,N_8176,N_8141);
nand U8251 (N_8251,N_8150,N_8153);
nor U8252 (N_8252,N_8175,N_8195);
and U8253 (N_8253,N_8148,N_8159);
nor U8254 (N_8254,N_8120,N_8199);
and U8255 (N_8255,N_8184,N_8120);
xor U8256 (N_8256,N_8111,N_8120);
xor U8257 (N_8257,N_8157,N_8152);
xnor U8258 (N_8258,N_8102,N_8105);
nor U8259 (N_8259,N_8138,N_8195);
xnor U8260 (N_8260,N_8130,N_8106);
xor U8261 (N_8261,N_8139,N_8132);
xor U8262 (N_8262,N_8124,N_8153);
xnor U8263 (N_8263,N_8147,N_8151);
nand U8264 (N_8264,N_8180,N_8143);
and U8265 (N_8265,N_8157,N_8124);
nand U8266 (N_8266,N_8146,N_8125);
xor U8267 (N_8267,N_8182,N_8197);
nand U8268 (N_8268,N_8103,N_8156);
nand U8269 (N_8269,N_8175,N_8122);
xor U8270 (N_8270,N_8144,N_8161);
and U8271 (N_8271,N_8154,N_8134);
nor U8272 (N_8272,N_8108,N_8117);
or U8273 (N_8273,N_8174,N_8181);
xor U8274 (N_8274,N_8156,N_8182);
and U8275 (N_8275,N_8186,N_8198);
or U8276 (N_8276,N_8196,N_8136);
and U8277 (N_8277,N_8147,N_8121);
nand U8278 (N_8278,N_8155,N_8182);
nor U8279 (N_8279,N_8186,N_8111);
or U8280 (N_8280,N_8131,N_8140);
xnor U8281 (N_8281,N_8109,N_8187);
nor U8282 (N_8282,N_8112,N_8102);
nor U8283 (N_8283,N_8190,N_8111);
and U8284 (N_8284,N_8169,N_8118);
or U8285 (N_8285,N_8130,N_8118);
nor U8286 (N_8286,N_8154,N_8156);
nor U8287 (N_8287,N_8137,N_8184);
nand U8288 (N_8288,N_8159,N_8131);
xor U8289 (N_8289,N_8157,N_8174);
xor U8290 (N_8290,N_8175,N_8170);
or U8291 (N_8291,N_8121,N_8168);
xor U8292 (N_8292,N_8134,N_8115);
xor U8293 (N_8293,N_8145,N_8132);
nor U8294 (N_8294,N_8163,N_8137);
nand U8295 (N_8295,N_8159,N_8172);
nor U8296 (N_8296,N_8145,N_8144);
nor U8297 (N_8297,N_8133,N_8114);
nand U8298 (N_8298,N_8114,N_8141);
or U8299 (N_8299,N_8184,N_8125);
nor U8300 (N_8300,N_8215,N_8243);
nand U8301 (N_8301,N_8283,N_8225);
nand U8302 (N_8302,N_8237,N_8291);
xor U8303 (N_8303,N_8251,N_8207);
xnor U8304 (N_8304,N_8297,N_8254);
or U8305 (N_8305,N_8270,N_8234);
and U8306 (N_8306,N_8290,N_8273);
nand U8307 (N_8307,N_8238,N_8249);
nand U8308 (N_8308,N_8267,N_8213);
nand U8309 (N_8309,N_8221,N_8248);
or U8310 (N_8310,N_8271,N_8240);
xnor U8311 (N_8311,N_8292,N_8287);
nor U8312 (N_8312,N_8289,N_8284);
or U8313 (N_8313,N_8212,N_8241);
or U8314 (N_8314,N_8272,N_8210);
nand U8315 (N_8315,N_8204,N_8223);
nor U8316 (N_8316,N_8224,N_8252);
or U8317 (N_8317,N_8285,N_8260);
nor U8318 (N_8318,N_8259,N_8263);
nand U8319 (N_8319,N_8274,N_8230);
xnor U8320 (N_8320,N_8246,N_8266);
and U8321 (N_8321,N_8253,N_8233);
or U8322 (N_8322,N_8288,N_8218);
or U8323 (N_8323,N_8247,N_8217);
xor U8324 (N_8324,N_8277,N_8286);
nand U8325 (N_8325,N_8236,N_8276);
nand U8326 (N_8326,N_8235,N_8299);
or U8327 (N_8327,N_8232,N_8282);
or U8328 (N_8328,N_8205,N_8214);
nand U8329 (N_8329,N_8257,N_8226);
xnor U8330 (N_8330,N_8262,N_8268);
xnor U8331 (N_8331,N_8203,N_8245);
nor U8332 (N_8332,N_8269,N_8264);
and U8333 (N_8333,N_8298,N_8201);
xor U8334 (N_8334,N_8229,N_8220);
nand U8335 (N_8335,N_8293,N_8275);
nand U8336 (N_8336,N_8200,N_8278);
or U8337 (N_8337,N_8256,N_8239);
or U8338 (N_8338,N_8242,N_8279);
xor U8339 (N_8339,N_8211,N_8261);
and U8340 (N_8340,N_8228,N_8219);
or U8341 (N_8341,N_8280,N_8255);
xnor U8342 (N_8342,N_8209,N_8258);
xor U8343 (N_8343,N_8206,N_8296);
nand U8344 (N_8344,N_8244,N_8250);
xor U8345 (N_8345,N_8281,N_8216);
and U8346 (N_8346,N_8202,N_8227);
and U8347 (N_8347,N_8294,N_8231);
nor U8348 (N_8348,N_8265,N_8222);
xor U8349 (N_8349,N_8295,N_8208);
nor U8350 (N_8350,N_8220,N_8231);
nor U8351 (N_8351,N_8268,N_8282);
nand U8352 (N_8352,N_8267,N_8223);
or U8353 (N_8353,N_8260,N_8219);
and U8354 (N_8354,N_8233,N_8257);
nor U8355 (N_8355,N_8230,N_8233);
nor U8356 (N_8356,N_8228,N_8280);
or U8357 (N_8357,N_8252,N_8204);
nor U8358 (N_8358,N_8204,N_8228);
and U8359 (N_8359,N_8218,N_8240);
or U8360 (N_8360,N_8204,N_8240);
and U8361 (N_8361,N_8202,N_8217);
and U8362 (N_8362,N_8203,N_8227);
xor U8363 (N_8363,N_8256,N_8297);
or U8364 (N_8364,N_8206,N_8277);
or U8365 (N_8365,N_8209,N_8257);
xor U8366 (N_8366,N_8227,N_8213);
and U8367 (N_8367,N_8239,N_8282);
and U8368 (N_8368,N_8252,N_8212);
nand U8369 (N_8369,N_8218,N_8265);
and U8370 (N_8370,N_8298,N_8284);
nand U8371 (N_8371,N_8237,N_8290);
or U8372 (N_8372,N_8281,N_8284);
xor U8373 (N_8373,N_8217,N_8219);
xor U8374 (N_8374,N_8298,N_8281);
nor U8375 (N_8375,N_8271,N_8232);
nand U8376 (N_8376,N_8293,N_8247);
nor U8377 (N_8377,N_8266,N_8236);
and U8378 (N_8378,N_8222,N_8209);
nor U8379 (N_8379,N_8274,N_8218);
and U8380 (N_8380,N_8229,N_8264);
and U8381 (N_8381,N_8247,N_8202);
or U8382 (N_8382,N_8229,N_8273);
xnor U8383 (N_8383,N_8225,N_8220);
and U8384 (N_8384,N_8260,N_8242);
nand U8385 (N_8385,N_8270,N_8230);
xnor U8386 (N_8386,N_8282,N_8259);
nor U8387 (N_8387,N_8218,N_8257);
or U8388 (N_8388,N_8229,N_8266);
xor U8389 (N_8389,N_8263,N_8222);
nor U8390 (N_8390,N_8209,N_8292);
or U8391 (N_8391,N_8250,N_8204);
nor U8392 (N_8392,N_8235,N_8238);
nand U8393 (N_8393,N_8290,N_8263);
nand U8394 (N_8394,N_8263,N_8228);
or U8395 (N_8395,N_8241,N_8255);
nand U8396 (N_8396,N_8210,N_8228);
or U8397 (N_8397,N_8210,N_8235);
xnor U8398 (N_8398,N_8207,N_8288);
xnor U8399 (N_8399,N_8249,N_8288);
or U8400 (N_8400,N_8342,N_8345);
or U8401 (N_8401,N_8320,N_8388);
or U8402 (N_8402,N_8334,N_8385);
or U8403 (N_8403,N_8378,N_8379);
nand U8404 (N_8404,N_8351,N_8374);
nor U8405 (N_8405,N_8398,N_8317);
nor U8406 (N_8406,N_8354,N_8343);
xnor U8407 (N_8407,N_8375,N_8336);
and U8408 (N_8408,N_8363,N_8358);
or U8409 (N_8409,N_8356,N_8327);
or U8410 (N_8410,N_8310,N_8316);
xnor U8411 (N_8411,N_8326,N_8332);
xnor U8412 (N_8412,N_8384,N_8312);
or U8413 (N_8413,N_8355,N_8353);
and U8414 (N_8414,N_8302,N_8307);
xor U8415 (N_8415,N_8365,N_8382);
nor U8416 (N_8416,N_8367,N_8390);
and U8417 (N_8417,N_8318,N_8369);
nand U8418 (N_8418,N_8322,N_8377);
nor U8419 (N_8419,N_8364,N_8340);
nand U8420 (N_8420,N_8319,N_8399);
or U8421 (N_8421,N_8325,N_8339);
nor U8422 (N_8422,N_8372,N_8394);
and U8423 (N_8423,N_8357,N_8370);
xnor U8424 (N_8424,N_8389,N_8306);
or U8425 (N_8425,N_8338,N_8328);
nand U8426 (N_8426,N_8313,N_8348);
nand U8427 (N_8427,N_8315,N_8383);
or U8428 (N_8428,N_8335,N_8330);
xnor U8429 (N_8429,N_8300,N_8323);
or U8430 (N_8430,N_8349,N_8329);
or U8431 (N_8431,N_8333,N_8362);
nor U8432 (N_8432,N_8341,N_8350);
or U8433 (N_8433,N_8371,N_8380);
and U8434 (N_8434,N_8397,N_8314);
xor U8435 (N_8435,N_8393,N_8308);
or U8436 (N_8436,N_8321,N_8361);
and U8437 (N_8437,N_8301,N_8386);
or U8438 (N_8438,N_8309,N_8381);
nand U8439 (N_8439,N_8359,N_8396);
nor U8440 (N_8440,N_8395,N_8368);
nor U8441 (N_8441,N_8304,N_8324);
nor U8442 (N_8442,N_8376,N_8360);
and U8443 (N_8443,N_8346,N_8387);
and U8444 (N_8444,N_8352,N_8344);
and U8445 (N_8445,N_8303,N_8373);
or U8446 (N_8446,N_8337,N_8331);
and U8447 (N_8447,N_8392,N_8347);
nand U8448 (N_8448,N_8391,N_8311);
xor U8449 (N_8449,N_8366,N_8305);
xnor U8450 (N_8450,N_8381,N_8314);
nor U8451 (N_8451,N_8353,N_8318);
nor U8452 (N_8452,N_8375,N_8383);
and U8453 (N_8453,N_8393,N_8377);
and U8454 (N_8454,N_8360,N_8369);
nor U8455 (N_8455,N_8343,N_8391);
xor U8456 (N_8456,N_8314,N_8347);
nand U8457 (N_8457,N_8362,N_8340);
xnor U8458 (N_8458,N_8396,N_8379);
nor U8459 (N_8459,N_8389,N_8341);
nand U8460 (N_8460,N_8355,N_8371);
or U8461 (N_8461,N_8303,N_8307);
nand U8462 (N_8462,N_8369,N_8380);
nand U8463 (N_8463,N_8328,N_8330);
nor U8464 (N_8464,N_8354,N_8391);
nand U8465 (N_8465,N_8325,N_8379);
nor U8466 (N_8466,N_8323,N_8313);
nand U8467 (N_8467,N_8398,N_8314);
xor U8468 (N_8468,N_8377,N_8350);
or U8469 (N_8469,N_8301,N_8383);
xor U8470 (N_8470,N_8387,N_8343);
nand U8471 (N_8471,N_8337,N_8361);
nand U8472 (N_8472,N_8388,N_8360);
nor U8473 (N_8473,N_8360,N_8368);
and U8474 (N_8474,N_8303,N_8310);
or U8475 (N_8475,N_8307,N_8314);
and U8476 (N_8476,N_8361,N_8357);
nand U8477 (N_8477,N_8367,N_8315);
or U8478 (N_8478,N_8384,N_8338);
or U8479 (N_8479,N_8375,N_8365);
nor U8480 (N_8480,N_8399,N_8357);
xnor U8481 (N_8481,N_8312,N_8329);
xor U8482 (N_8482,N_8307,N_8318);
and U8483 (N_8483,N_8357,N_8346);
or U8484 (N_8484,N_8393,N_8326);
xnor U8485 (N_8485,N_8375,N_8364);
nand U8486 (N_8486,N_8354,N_8339);
or U8487 (N_8487,N_8366,N_8300);
xor U8488 (N_8488,N_8367,N_8364);
xnor U8489 (N_8489,N_8304,N_8354);
or U8490 (N_8490,N_8309,N_8393);
and U8491 (N_8491,N_8358,N_8365);
xor U8492 (N_8492,N_8327,N_8393);
or U8493 (N_8493,N_8353,N_8340);
nor U8494 (N_8494,N_8388,N_8367);
and U8495 (N_8495,N_8328,N_8394);
xor U8496 (N_8496,N_8389,N_8399);
and U8497 (N_8497,N_8300,N_8397);
and U8498 (N_8498,N_8336,N_8378);
xnor U8499 (N_8499,N_8373,N_8321);
nand U8500 (N_8500,N_8434,N_8476);
and U8501 (N_8501,N_8405,N_8478);
nand U8502 (N_8502,N_8407,N_8492);
and U8503 (N_8503,N_8458,N_8424);
xnor U8504 (N_8504,N_8401,N_8429);
and U8505 (N_8505,N_8426,N_8490);
nand U8506 (N_8506,N_8451,N_8443);
and U8507 (N_8507,N_8467,N_8499);
and U8508 (N_8508,N_8488,N_8436);
nand U8509 (N_8509,N_8420,N_8417);
and U8510 (N_8510,N_8452,N_8450);
nor U8511 (N_8511,N_8447,N_8442);
nand U8512 (N_8512,N_8462,N_8433);
xor U8513 (N_8513,N_8441,N_8494);
nor U8514 (N_8514,N_8482,N_8414);
nand U8515 (N_8515,N_8483,N_8409);
nor U8516 (N_8516,N_8425,N_8491);
nand U8517 (N_8517,N_8493,N_8431);
or U8518 (N_8518,N_8446,N_8470);
xor U8519 (N_8519,N_8416,N_8485);
nand U8520 (N_8520,N_8464,N_8468);
nand U8521 (N_8521,N_8496,N_8438);
nand U8522 (N_8522,N_8472,N_8456);
and U8523 (N_8523,N_8459,N_8466);
nand U8524 (N_8524,N_8413,N_8439);
and U8525 (N_8525,N_8453,N_8463);
xnor U8526 (N_8526,N_8444,N_8455);
or U8527 (N_8527,N_8477,N_8418);
or U8528 (N_8528,N_8486,N_8460);
and U8529 (N_8529,N_8435,N_8475);
or U8530 (N_8530,N_8403,N_8495);
nor U8531 (N_8531,N_8400,N_8497);
nor U8532 (N_8532,N_8481,N_8415);
or U8533 (N_8533,N_8484,N_8422);
and U8534 (N_8534,N_8408,N_8428);
nand U8535 (N_8535,N_8487,N_8474);
and U8536 (N_8536,N_8412,N_8498);
and U8537 (N_8537,N_8473,N_8430);
nor U8538 (N_8538,N_8419,N_8449);
nor U8539 (N_8539,N_8406,N_8421);
nand U8540 (N_8540,N_8404,N_8448);
nand U8541 (N_8541,N_8423,N_8461);
nor U8542 (N_8542,N_8471,N_8480);
nand U8543 (N_8543,N_8465,N_8411);
and U8544 (N_8544,N_8457,N_8402);
nor U8545 (N_8545,N_8454,N_8445);
or U8546 (N_8546,N_8469,N_8489);
nor U8547 (N_8547,N_8410,N_8427);
or U8548 (N_8548,N_8437,N_8432);
or U8549 (N_8549,N_8440,N_8479);
or U8550 (N_8550,N_8453,N_8480);
or U8551 (N_8551,N_8489,N_8480);
xor U8552 (N_8552,N_8461,N_8406);
and U8553 (N_8553,N_8498,N_8430);
and U8554 (N_8554,N_8444,N_8475);
or U8555 (N_8555,N_8448,N_8416);
and U8556 (N_8556,N_8487,N_8473);
and U8557 (N_8557,N_8476,N_8489);
or U8558 (N_8558,N_8452,N_8462);
nor U8559 (N_8559,N_8461,N_8441);
nor U8560 (N_8560,N_8402,N_8418);
nor U8561 (N_8561,N_8486,N_8412);
nor U8562 (N_8562,N_8490,N_8427);
or U8563 (N_8563,N_8415,N_8430);
nand U8564 (N_8564,N_8442,N_8413);
and U8565 (N_8565,N_8423,N_8402);
nand U8566 (N_8566,N_8433,N_8476);
and U8567 (N_8567,N_8404,N_8460);
xnor U8568 (N_8568,N_8480,N_8440);
nand U8569 (N_8569,N_8400,N_8464);
xnor U8570 (N_8570,N_8442,N_8438);
xor U8571 (N_8571,N_8410,N_8400);
and U8572 (N_8572,N_8473,N_8402);
and U8573 (N_8573,N_8470,N_8406);
nand U8574 (N_8574,N_8468,N_8451);
or U8575 (N_8575,N_8427,N_8406);
and U8576 (N_8576,N_8450,N_8404);
nor U8577 (N_8577,N_8423,N_8408);
xor U8578 (N_8578,N_8454,N_8453);
and U8579 (N_8579,N_8464,N_8431);
xor U8580 (N_8580,N_8430,N_8468);
or U8581 (N_8581,N_8424,N_8456);
xnor U8582 (N_8582,N_8439,N_8487);
xor U8583 (N_8583,N_8405,N_8473);
nand U8584 (N_8584,N_8412,N_8476);
and U8585 (N_8585,N_8416,N_8409);
nor U8586 (N_8586,N_8445,N_8434);
xnor U8587 (N_8587,N_8408,N_8430);
nor U8588 (N_8588,N_8484,N_8457);
nand U8589 (N_8589,N_8431,N_8415);
or U8590 (N_8590,N_8482,N_8459);
or U8591 (N_8591,N_8479,N_8400);
nand U8592 (N_8592,N_8417,N_8488);
and U8593 (N_8593,N_8448,N_8433);
nor U8594 (N_8594,N_8456,N_8447);
nor U8595 (N_8595,N_8420,N_8463);
xor U8596 (N_8596,N_8444,N_8496);
xnor U8597 (N_8597,N_8445,N_8487);
nand U8598 (N_8598,N_8475,N_8409);
nor U8599 (N_8599,N_8413,N_8489);
and U8600 (N_8600,N_8577,N_8585);
nand U8601 (N_8601,N_8516,N_8503);
nor U8602 (N_8602,N_8519,N_8551);
xnor U8603 (N_8603,N_8504,N_8562);
nor U8604 (N_8604,N_8525,N_8576);
or U8605 (N_8605,N_8534,N_8568);
nand U8606 (N_8606,N_8500,N_8587);
nand U8607 (N_8607,N_8540,N_8547);
nor U8608 (N_8608,N_8589,N_8512);
or U8609 (N_8609,N_8535,N_8506);
nand U8610 (N_8610,N_8537,N_8567);
or U8611 (N_8611,N_8505,N_8598);
xnor U8612 (N_8612,N_8565,N_8559);
or U8613 (N_8613,N_8550,N_8556);
or U8614 (N_8614,N_8592,N_8526);
xnor U8615 (N_8615,N_8513,N_8510);
nor U8616 (N_8616,N_8594,N_8569);
or U8617 (N_8617,N_8541,N_8524);
nor U8618 (N_8618,N_8578,N_8511);
and U8619 (N_8619,N_8501,N_8544);
or U8620 (N_8620,N_8579,N_8523);
nand U8621 (N_8621,N_8588,N_8560);
xor U8622 (N_8622,N_8502,N_8542);
nor U8623 (N_8623,N_8557,N_8521);
nor U8624 (N_8624,N_8546,N_8517);
and U8625 (N_8625,N_8520,N_8536);
and U8626 (N_8626,N_8518,N_8584);
nor U8627 (N_8627,N_8583,N_8533);
nand U8628 (N_8628,N_8528,N_8561);
and U8629 (N_8629,N_8596,N_8571);
nand U8630 (N_8630,N_8564,N_8509);
nor U8631 (N_8631,N_8580,N_8590);
xnor U8632 (N_8632,N_8573,N_8595);
or U8633 (N_8633,N_8597,N_8545);
nand U8634 (N_8634,N_8558,N_8543);
or U8635 (N_8635,N_8574,N_8527);
xnor U8636 (N_8636,N_8530,N_8514);
xnor U8637 (N_8637,N_8599,N_8563);
nor U8638 (N_8638,N_8591,N_8553);
or U8639 (N_8639,N_8531,N_8522);
or U8640 (N_8640,N_8566,N_8575);
or U8641 (N_8641,N_8548,N_8572);
xnor U8642 (N_8642,N_8570,N_8515);
and U8643 (N_8643,N_8552,N_8507);
and U8644 (N_8644,N_8539,N_8555);
nor U8645 (N_8645,N_8582,N_8554);
nand U8646 (N_8646,N_8508,N_8586);
or U8647 (N_8647,N_8529,N_8538);
and U8648 (N_8648,N_8581,N_8549);
or U8649 (N_8649,N_8593,N_8532);
nand U8650 (N_8650,N_8588,N_8519);
xnor U8651 (N_8651,N_8558,N_8539);
nand U8652 (N_8652,N_8534,N_8553);
xor U8653 (N_8653,N_8561,N_8543);
and U8654 (N_8654,N_8567,N_8538);
xor U8655 (N_8655,N_8566,N_8513);
nor U8656 (N_8656,N_8510,N_8534);
xor U8657 (N_8657,N_8573,N_8568);
xnor U8658 (N_8658,N_8506,N_8507);
and U8659 (N_8659,N_8505,N_8585);
nand U8660 (N_8660,N_8528,N_8508);
or U8661 (N_8661,N_8523,N_8558);
or U8662 (N_8662,N_8527,N_8598);
nor U8663 (N_8663,N_8515,N_8518);
and U8664 (N_8664,N_8530,N_8598);
or U8665 (N_8665,N_8511,N_8560);
nor U8666 (N_8666,N_8579,N_8526);
xor U8667 (N_8667,N_8539,N_8533);
nor U8668 (N_8668,N_8510,N_8512);
or U8669 (N_8669,N_8580,N_8593);
nor U8670 (N_8670,N_8576,N_8581);
nand U8671 (N_8671,N_8573,N_8534);
and U8672 (N_8672,N_8524,N_8562);
nand U8673 (N_8673,N_8563,N_8511);
nor U8674 (N_8674,N_8520,N_8559);
and U8675 (N_8675,N_8540,N_8516);
and U8676 (N_8676,N_8586,N_8537);
nand U8677 (N_8677,N_8588,N_8584);
nor U8678 (N_8678,N_8583,N_8555);
xor U8679 (N_8679,N_8502,N_8546);
nand U8680 (N_8680,N_8564,N_8591);
or U8681 (N_8681,N_8560,N_8529);
nor U8682 (N_8682,N_8597,N_8589);
or U8683 (N_8683,N_8516,N_8568);
nor U8684 (N_8684,N_8577,N_8598);
or U8685 (N_8685,N_8582,N_8558);
or U8686 (N_8686,N_8580,N_8551);
nor U8687 (N_8687,N_8562,N_8515);
nor U8688 (N_8688,N_8576,N_8598);
and U8689 (N_8689,N_8530,N_8599);
or U8690 (N_8690,N_8559,N_8556);
nand U8691 (N_8691,N_8535,N_8595);
nor U8692 (N_8692,N_8590,N_8583);
and U8693 (N_8693,N_8558,N_8552);
or U8694 (N_8694,N_8552,N_8599);
or U8695 (N_8695,N_8527,N_8541);
and U8696 (N_8696,N_8558,N_8560);
xor U8697 (N_8697,N_8503,N_8549);
or U8698 (N_8698,N_8517,N_8506);
nand U8699 (N_8699,N_8556,N_8529);
or U8700 (N_8700,N_8646,N_8640);
xnor U8701 (N_8701,N_8633,N_8624);
or U8702 (N_8702,N_8622,N_8605);
xor U8703 (N_8703,N_8601,N_8698);
nor U8704 (N_8704,N_8682,N_8650);
nor U8705 (N_8705,N_8612,N_8685);
or U8706 (N_8706,N_8630,N_8666);
and U8707 (N_8707,N_8672,N_8618);
or U8708 (N_8708,N_8679,N_8675);
xnor U8709 (N_8709,N_8694,N_8692);
nand U8710 (N_8710,N_8649,N_8623);
or U8711 (N_8711,N_8652,N_8603);
or U8712 (N_8712,N_8687,N_8637);
xor U8713 (N_8713,N_8639,N_8688);
xor U8714 (N_8714,N_8654,N_8689);
and U8715 (N_8715,N_8631,N_8684);
and U8716 (N_8716,N_8610,N_8670);
and U8717 (N_8717,N_8608,N_8647);
and U8718 (N_8718,N_8667,N_8665);
and U8719 (N_8719,N_8609,N_8607);
xnor U8720 (N_8720,N_8645,N_8660);
xor U8721 (N_8721,N_8634,N_8641);
nor U8722 (N_8722,N_8628,N_8600);
nand U8723 (N_8723,N_8655,N_8695);
nor U8724 (N_8724,N_8677,N_8669);
nand U8725 (N_8725,N_8602,N_8656);
xnor U8726 (N_8726,N_8611,N_8657);
nand U8727 (N_8727,N_8668,N_8659);
xor U8728 (N_8728,N_8614,N_8636);
nand U8729 (N_8729,N_8606,N_8680);
nor U8730 (N_8730,N_8693,N_8625);
xor U8731 (N_8731,N_8683,N_8619);
nand U8732 (N_8732,N_8615,N_8676);
and U8733 (N_8733,N_8697,N_8644);
xnor U8734 (N_8734,N_8696,N_8661);
or U8735 (N_8735,N_8658,N_8620);
or U8736 (N_8736,N_8627,N_8616);
or U8737 (N_8737,N_8663,N_8662);
xor U8738 (N_8738,N_8626,N_8629);
xnor U8739 (N_8739,N_8651,N_8690);
and U8740 (N_8740,N_8681,N_8642);
or U8741 (N_8741,N_8648,N_8632);
nor U8742 (N_8742,N_8686,N_8674);
and U8743 (N_8743,N_8673,N_8638);
xor U8744 (N_8744,N_8643,N_8691);
nor U8745 (N_8745,N_8653,N_8664);
nand U8746 (N_8746,N_8604,N_8678);
xor U8747 (N_8747,N_8635,N_8671);
or U8748 (N_8748,N_8699,N_8621);
or U8749 (N_8749,N_8617,N_8613);
or U8750 (N_8750,N_8680,N_8659);
or U8751 (N_8751,N_8618,N_8676);
or U8752 (N_8752,N_8628,N_8647);
xor U8753 (N_8753,N_8693,N_8673);
xnor U8754 (N_8754,N_8642,N_8611);
xor U8755 (N_8755,N_8696,N_8603);
or U8756 (N_8756,N_8663,N_8669);
xor U8757 (N_8757,N_8683,N_8632);
xnor U8758 (N_8758,N_8600,N_8686);
xor U8759 (N_8759,N_8670,N_8622);
or U8760 (N_8760,N_8643,N_8676);
or U8761 (N_8761,N_8616,N_8666);
and U8762 (N_8762,N_8646,N_8621);
and U8763 (N_8763,N_8622,N_8625);
nand U8764 (N_8764,N_8680,N_8611);
or U8765 (N_8765,N_8659,N_8644);
nand U8766 (N_8766,N_8683,N_8644);
or U8767 (N_8767,N_8647,N_8610);
nor U8768 (N_8768,N_8690,N_8637);
nand U8769 (N_8769,N_8685,N_8649);
xor U8770 (N_8770,N_8653,N_8665);
nor U8771 (N_8771,N_8616,N_8694);
nand U8772 (N_8772,N_8654,N_8619);
and U8773 (N_8773,N_8648,N_8638);
or U8774 (N_8774,N_8661,N_8692);
or U8775 (N_8775,N_8626,N_8645);
and U8776 (N_8776,N_8626,N_8684);
nand U8777 (N_8777,N_8672,N_8621);
nor U8778 (N_8778,N_8632,N_8659);
nand U8779 (N_8779,N_8615,N_8678);
xnor U8780 (N_8780,N_8658,N_8683);
or U8781 (N_8781,N_8634,N_8680);
and U8782 (N_8782,N_8692,N_8689);
nand U8783 (N_8783,N_8699,N_8667);
or U8784 (N_8784,N_8675,N_8608);
nand U8785 (N_8785,N_8699,N_8619);
nand U8786 (N_8786,N_8608,N_8602);
or U8787 (N_8787,N_8694,N_8619);
nor U8788 (N_8788,N_8667,N_8687);
xor U8789 (N_8789,N_8620,N_8675);
nand U8790 (N_8790,N_8688,N_8601);
nor U8791 (N_8791,N_8620,N_8611);
nand U8792 (N_8792,N_8698,N_8602);
xor U8793 (N_8793,N_8638,N_8633);
xor U8794 (N_8794,N_8628,N_8680);
or U8795 (N_8795,N_8605,N_8647);
or U8796 (N_8796,N_8636,N_8672);
or U8797 (N_8797,N_8674,N_8684);
and U8798 (N_8798,N_8683,N_8691);
and U8799 (N_8799,N_8649,N_8671);
and U8800 (N_8800,N_8768,N_8706);
nor U8801 (N_8801,N_8785,N_8742);
and U8802 (N_8802,N_8756,N_8751);
xor U8803 (N_8803,N_8708,N_8704);
nor U8804 (N_8804,N_8799,N_8783);
nand U8805 (N_8805,N_8792,N_8718);
or U8806 (N_8806,N_8720,N_8789);
nor U8807 (N_8807,N_8744,N_8724);
or U8808 (N_8808,N_8710,N_8726);
xnor U8809 (N_8809,N_8702,N_8764);
or U8810 (N_8810,N_8763,N_8762);
nor U8811 (N_8811,N_8771,N_8741);
and U8812 (N_8812,N_8758,N_8767);
and U8813 (N_8813,N_8759,N_8788);
xnor U8814 (N_8814,N_8773,N_8716);
nand U8815 (N_8815,N_8735,N_8750);
xor U8816 (N_8816,N_8700,N_8795);
nand U8817 (N_8817,N_8715,N_8757);
xor U8818 (N_8818,N_8780,N_8761);
nand U8819 (N_8819,N_8729,N_8745);
nor U8820 (N_8820,N_8717,N_8787);
nor U8821 (N_8821,N_8727,N_8711);
nor U8822 (N_8822,N_8743,N_8733);
nor U8823 (N_8823,N_8797,N_8793);
or U8824 (N_8824,N_8714,N_8734);
or U8825 (N_8825,N_8738,N_8746);
xor U8826 (N_8826,N_8769,N_8730);
nand U8827 (N_8827,N_8760,N_8798);
nand U8828 (N_8828,N_8731,N_8736);
xor U8829 (N_8829,N_8755,N_8747);
and U8830 (N_8830,N_8790,N_8732);
xor U8831 (N_8831,N_8739,N_8709);
or U8832 (N_8832,N_8740,N_8753);
nand U8833 (N_8833,N_8703,N_8701);
nor U8834 (N_8834,N_8772,N_8775);
and U8835 (N_8835,N_8737,N_8728);
or U8836 (N_8836,N_8782,N_8705);
nor U8837 (N_8837,N_8781,N_8719);
or U8838 (N_8838,N_8779,N_8784);
xnor U8839 (N_8839,N_8786,N_8777);
or U8840 (N_8840,N_8794,N_8748);
xnor U8841 (N_8841,N_8713,N_8712);
nor U8842 (N_8842,N_8752,N_8796);
and U8843 (N_8843,N_8754,N_8774);
and U8844 (N_8844,N_8749,N_8723);
nor U8845 (N_8845,N_8776,N_8770);
and U8846 (N_8846,N_8725,N_8722);
and U8847 (N_8847,N_8778,N_8707);
nor U8848 (N_8848,N_8721,N_8765);
xnor U8849 (N_8849,N_8791,N_8766);
xor U8850 (N_8850,N_8738,N_8761);
and U8851 (N_8851,N_8753,N_8717);
and U8852 (N_8852,N_8706,N_8781);
and U8853 (N_8853,N_8777,N_8709);
nor U8854 (N_8854,N_8774,N_8792);
or U8855 (N_8855,N_8725,N_8731);
xnor U8856 (N_8856,N_8785,N_8765);
xnor U8857 (N_8857,N_8779,N_8740);
or U8858 (N_8858,N_8798,N_8764);
xnor U8859 (N_8859,N_8777,N_8747);
nand U8860 (N_8860,N_8714,N_8747);
or U8861 (N_8861,N_8784,N_8701);
or U8862 (N_8862,N_8758,N_8745);
nor U8863 (N_8863,N_8721,N_8716);
or U8864 (N_8864,N_8700,N_8770);
or U8865 (N_8865,N_8717,N_8754);
or U8866 (N_8866,N_8708,N_8759);
nor U8867 (N_8867,N_8765,N_8715);
nor U8868 (N_8868,N_8780,N_8775);
or U8869 (N_8869,N_8729,N_8752);
nand U8870 (N_8870,N_8733,N_8750);
xor U8871 (N_8871,N_8756,N_8739);
xnor U8872 (N_8872,N_8757,N_8790);
nor U8873 (N_8873,N_8714,N_8720);
xnor U8874 (N_8874,N_8749,N_8790);
nor U8875 (N_8875,N_8744,N_8719);
nand U8876 (N_8876,N_8790,N_8796);
nand U8877 (N_8877,N_8777,N_8705);
and U8878 (N_8878,N_8756,N_8765);
or U8879 (N_8879,N_8727,N_8701);
xnor U8880 (N_8880,N_8751,N_8708);
xnor U8881 (N_8881,N_8735,N_8731);
xnor U8882 (N_8882,N_8729,N_8708);
xnor U8883 (N_8883,N_8746,N_8798);
nand U8884 (N_8884,N_8796,N_8723);
or U8885 (N_8885,N_8738,N_8718);
xor U8886 (N_8886,N_8787,N_8747);
xnor U8887 (N_8887,N_8703,N_8720);
nand U8888 (N_8888,N_8737,N_8796);
xor U8889 (N_8889,N_8797,N_8710);
xnor U8890 (N_8890,N_8750,N_8798);
or U8891 (N_8891,N_8779,N_8756);
or U8892 (N_8892,N_8735,N_8777);
nand U8893 (N_8893,N_8775,N_8729);
xnor U8894 (N_8894,N_8791,N_8748);
xor U8895 (N_8895,N_8770,N_8775);
and U8896 (N_8896,N_8779,N_8777);
xor U8897 (N_8897,N_8738,N_8767);
xnor U8898 (N_8898,N_8738,N_8712);
and U8899 (N_8899,N_8778,N_8773);
nor U8900 (N_8900,N_8836,N_8886);
or U8901 (N_8901,N_8894,N_8800);
and U8902 (N_8902,N_8827,N_8814);
and U8903 (N_8903,N_8875,N_8857);
xor U8904 (N_8904,N_8851,N_8834);
xnor U8905 (N_8905,N_8853,N_8861);
nand U8906 (N_8906,N_8896,N_8842);
or U8907 (N_8907,N_8813,N_8816);
xnor U8908 (N_8908,N_8845,N_8870);
or U8909 (N_8909,N_8890,N_8844);
nand U8910 (N_8910,N_8899,N_8806);
or U8911 (N_8911,N_8855,N_8868);
or U8912 (N_8912,N_8880,N_8881);
or U8913 (N_8913,N_8898,N_8849);
nand U8914 (N_8914,N_8815,N_8893);
nand U8915 (N_8915,N_8862,N_8883);
nor U8916 (N_8916,N_8877,N_8821);
and U8917 (N_8917,N_8804,N_8846);
and U8918 (N_8918,N_8879,N_8887);
nor U8919 (N_8919,N_8802,N_8865);
nor U8920 (N_8920,N_8869,N_8878);
or U8921 (N_8921,N_8805,N_8889);
xor U8922 (N_8922,N_8810,N_8830);
nor U8923 (N_8923,N_8837,N_8874);
xnor U8924 (N_8924,N_8848,N_8864);
nor U8925 (N_8925,N_8859,N_8854);
or U8926 (N_8926,N_8843,N_8825);
or U8927 (N_8927,N_8897,N_8803);
nor U8928 (N_8928,N_8847,N_8873);
nand U8929 (N_8929,N_8835,N_8867);
xnor U8930 (N_8930,N_8833,N_8812);
xnor U8931 (N_8931,N_8807,N_8820);
xor U8932 (N_8932,N_8871,N_8822);
and U8933 (N_8933,N_8882,N_8891);
and U8934 (N_8934,N_8892,N_8838);
or U8935 (N_8935,N_8824,N_8811);
or U8936 (N_8936,N_8829,N_8817);
and U8937 (N_8937,N_8819,N_8852);
or U8938 (N_8938,N_8885,N_8841);
nor U8939 (N_8939,N_8832,N_8828);
nand U8940 (N_8940,N_8866,N_8809);
or U8941 (N_8941,N_8801,N_8826);
or U8942 (N_8942,N_8895,N_8888);
nor U8943 (N_8943,N_8856,N_8831);
nand U8944 (N_8944,N_8872,N_8876);
or U8945 (N_8945,N_8823,N_8863);
xor U8946 (N_8946,N_8839,N_8818);
nand U8947 (N_8947,N_8884,N_8850);
xor U8948 (N_8948,N_8858,N_8860);
nor U8949 (N_8949,N_8808,N_8840);
or U8950 (N_8950,N_8832,N_8843);
xor U8951 (N_8951,N_8839,N_8866);
or U8952 (N_8952,N_8854,N_8824);
nand U8953 (N_8953,N_8875,N_8860);
xor U8954 (N_8954,N_8849,N_8865);
nor U8955 (N_8955,N_8878,N_8820);
nand U8956 (N_8956,N_8892,N_8821);
or U8957 (N_8957,N_8801,N_8897);
and U8958 (N_8958,N_8830,N_8868);
nand U8959 (N_8959,N_8814,N_8882);
and U8960 (N_8960,N_8811,N_8858);
and U8961 (N_8961,N_8885,N_8838);
nand U8962 (N_8962,N_8878,N_8844);
nand U8963 (N_8963,N_8847,N_8829);
xor U8964 (N_8964,N_8801,N_8838);
nor U8965 (N_8965,N_8889,N_8838);
nand U8966 (N_8966,N_8829,N_8819);
nand U8967 (N_8967,N_8881,N_8861);
xnor U8968 (N_8968,N_8804,N_8870);
and U8969 (N_8969,N_8801,N_8852);
nor U8970 (N_8970,N_8872,N_8816);
nand U8971 (N_8971,N_8837,N_8828);
and U8972 (N_8972,N_8859,N_8891);
or U8973 (N_8973,N_8809,N_8806);
nand U8974 (N_8974,N_8848,N_8877);
or U8975 (N_8975,N_8833,N_8885);
xnor U8976 (N_8976,N_8832,N_8858);
nor U8977 (N_8977,N_8897,N_8812);
and U8978 (N_8978,N_8808,N_8827);
nor U8979 (N_8979,N_8898,N_8857);
nand U8980 (N_8980,N_8827,N_8890);
nand U8981 (N_8981,N_8802,N_8892);
nand U8982 (N_8982,N_8879,N_8860);
nand U8983 (N_8983,N_8823,N_8860);
xnor U8984 (N_8984,N_8835,N_8825);
nand U8985 (N_8985,N_8801,N_8894);
and U8986 (N_8986,N_8811,N_8825);
nand U8987 (N_8987,N_8812,N_8803);
nor U8988 (N_8988,N_8842,N_8871);
nand U8989 (N_8989,N_8891,N_8895);
nor U8990 (N_8990,N_8826,N_8822);
xnor U8991 (N_8991,N_8842,N_8817);
nor U8992 (N_8992,N_8807,N_8861);
xnor U8993 (N_8993,N_8812,N_8843);
nor U8994 (N_8994,N_8805,N_8863);
or U8995 (N_8995,N_8870,N_8839);
xnor U8996 (N_8996,N_8820,N_8867);
or U8997 (N_8997,N_8848,N_8851);
and U8998 (N_8998,N_8851,N_8844);
or U8999 (N_8999,N_8878,N_8880);
and U9000 (N_9000,N_8972,N_8975);
nor U9001 (N_9001,N_8962,N_8993);
and U9002 (N_9002,N_8920,N_8958);
nand U9003 (N_9003,N_8997,N_8957);
or U9004 (N_9004,N_8982,N_8934);
xor U9005 (N_9005,N_8933,N_8990);
nor U9006 (N_9006,N_8900,N_8925);
nor U9007 (N_9007,N_8950,N_8952);
and U9008 (N_9008,N_8956,N_8977);
and U9009 (N_9009,N_8930,N_8943);
xnor U9010 (N_9010,N_8955,N_8953);
or U9011 (N_9011,N_8967,N_8968);
nand U9012 (N_9012,N_8991,N_8923);
or U9013 (N_9013,N_8909,N_8940);
nor U9014 (N_9014,N_8941,N_8939);
xnor U9015 (N_9015,N_8946,N_8919);
or U9016 (N_9016,N_8927,N_8981);
nor U9017 (N_9017,N_8903,N_8983);
or U9018 (N_9018,N_8986,N_8912);
nand U9019 (N_9019,N_8937,N_8987);
xor U9020 (N_9020,N_8947,N_8905);
nor U9021 (N_9021,N_8928,N_8918);
nor U9022 (N_9022,N_8942,N_8932);
and U9023 (N_9023,N_8964,N_8908);
or U9024 (N_9024,N_8963,N_8911);
and U9025 (N_9025,N_8954,N_8980);
and U9026 (N_9026,N_8974,N_8969);
and U9027 (N_9027,N_8935,N_8949);
nor U9028 (N_9028,N_8917,N_8966);
and U9029 (N_9029,N_8945,N_8936);
and U9030 (N_9030,N_8915,N_8929);
or U9031 (N_9031,N_8913,N_8902);
xnor U9032 (N_9032,N_8959,N_8914);
nand U9033 (N_9033,N_8984,N_8989);
xnor U9034 (N_9034,N_8960,N_8988);
or U9035 (N_9035,N_8995,N_8999);
nor U9036 (N_9036,N_8976,N_8921);
xnor U9037 (N_9037,N_8965,N_8985);
nor U9038 (N_9038,N_8996,N_8971);
nor U9039 (N_9039,N_8924,N_8961);
and U9040 (N_9040,N_8973,N_8994);
and U9041 (N_9041,N_8998,N_8926);
xor U9042 (N_9042,N_8931,N_8992);
and U9043 (N_9043,N_8938,N_8916);
nor U9044 (N_9044,N_8901,N_8979);
or U9045 (N_9045,N_8910,N_8951);
and U9046 (N_9046,N_8944,N_8948);
xnor U9047 (N_9047,N_8904,N_8906);
xnor U9048 (N_9048,N_8922,N_8907);
and U9049 (N_9049,N_8978,N_8970);
or U9050 (N_9050,N_8985,N_8995);
and U9051 (N_9051,N_8995,N_8925);
xnor U9052 (N_9052,N_8902,N_8933);
nand U9053 (N_9053,N_8942,N_8914);
or U9054 (N_9054,N_8965,N_8976);
nand U9055 (N_9055,N_8928,N_8934);
or U9056 (N_9056,N_8987,N_8983);
or U9057 (N_9057,N_8942,N_8967);
and U9058 (N_9058,N_8917,N_8941);
nor U9059 (N_9059,N_8991,N_8993);
or U9060 (N_9060,N_8946,N_8926);
nand U9061 (N_9061,N_8957,N_8947);
or U9062 (N_9062,N_8933,N_8951);
nand U9063 (N_9063,N_8972,N_8951);
nor U9064 (N_9064,N_8967,N_8955);
or U9065 (N_9065,N_8948,N_8956);
nor U9066 (N_9066,N_8938,N_8953);
or U9067 (N_9067,N_8951,N_8920);
nor U9068 (N_9068,N_8979,N_8968);
xor U9069 (N_9069,N_8985,N_8954);
nand U9070 (N_9070,N_8984,N_8924);
nand U9071 (N_9071,N_8966,N_8901);
xnor U9072 (N_9072,N_8987,N_8952);
xnor U9073 (N_9073,N_8976,N_8947);
nor U9074 (N_9074,N_8958,N_8969);
nand U9075 (N_9075,N_8948,N_8961);
nor U9076 (N_9076,N_8976,N_8920);
or U9077 (N_9077,N_8915,N_8943);
nand U9078 (N_9078,N_8934,N_8950);
and U9079 (N_9079,N_8984,N_8901);
nor U9080 (N_9080,N_8979,N_8912);
or U9081 (N_9081,N_8904,N_8910);
nor U9082 (N_9082,N_8906,N_8969);
and U9083 (N_9083,N_8914,N_8969);
nand U9084 (N_9084,N_8933,N_8976);
nand U9085 (N_9085,N_8984,N_8963);
nand U9086 (N_9086,N_8964,N_8951);
nor U9087 (N_9087,N_8924,N_8939);
nor U9088 (N_9088,N_8902,N_8909);
or U9089 (N_9089,N_8975,N_8934);
nor U9090 (N_9090,N_8932,N_8940);
and U9091 (N_9091,N_8974,N_8984);
nor U9092 (N_9092,N_8985,N_8988);
and U9093 (N_9093,N_8910,N_8925);
or U9094 (N_9094,N_8991,N_8920);
xnor U9095 (N_9095,N_8951,N_8919);
and U9096 (N_9096,N_8995,N_8906);
xor U9097 (N_9097,N_8908,N_8971);
and U9098 (N_9098,N_8926,N_8947);
or U9099 (N_9099,N_8992,N_8990);
or U9100 (N_9100,N_9017,N_9048);
or U9101 (N_9101,N_9085,N_9069);
nor U9102 (N_9102,N_9091,N_9074);
xor U9103 (N_9103,N_9066,N_9067);
nor U9104 (N_9104,N_9063,N_9098);
and U9105 (N_9105,N_9095,N_9092);
xor U9106 (N_9106,N_9007,N_9022);
and U9107 (N_9107,N_9009,N_9006);
nor U9108 (N_9108,N_9065,N_9028);
nand U9109 (N_9109,N_9050,N_9031);
xor U9110 (N_9110,N_9034,N_9082);
or U9111 (N_9111,N_9004,N_9099);
nand U9112 (N_9112,N_9057,N_9019);
nor U9113 (N_9113,N_9025,N_9011);
xor U9114 (N_9114,N_9027,N_9024);
nand U9115 (N_9115,N_9023,N_9077);
or U9116 (N_9116,N_9089,N_9052);
or U9117 (N_9117,N_9094,N_9042);
nand U9118 (N_9118,N_9093,N_9026);
nor U9119 (N_9119,N_9090,N_9029);
xor U9120 (N_9120,N_9043,N_9049);
nor U9121 (N_9121,N_9047,N_9015);
and U9122 (N_9122,N_9040,N_9014);
nand U9123 (N_9123,N_9075,N_9073);
and U9124 (N_9124,N_9058,N_9087);
nor U9125 (N_9125,N_9020,N_9037);
xnor U9126 (N_9126,N_9003,N_9084);
nand U9127 (N_9127,N_9096,N_9071);
nor U9128 (N_9128,N_9088,N_9080);
xor U9129 (N_9129,N_9072,N_9045);
or U9130 (N_9130,N_9081,N_9002);
or U9131 (N_9131,N_9044,N_9078);
xor U9132 (N_9132,N_9018,N_9000);
nor U9133 (N_9133,N_9001,N_9060);
nor U9134 (N_9134,N_9061,N_9041);
nand U9135 (N_9135,N_9046,N_9064);
xor U9136 (N_9136,N_9076,N_9053);
nand U9137 (N_9137,N_9038,N_9070);
or U9138 (N_9138,N_9021,N_9055);
nand U9139 (N_9139,N_9005,N_9079);
and U9140 (N_9140,N_9086,N_9032);
nand U9141 (N_9141,N_9039,N_9054);
nand U9142 (N_9142,N_9051,N_9013);
xnor U9143 (N_9143,N_9012,N_9035);
and U9144 (N_9144,N_9056,N_9008);
or U9145 (N_9145,N_9097,N_9068);
xor U9146 (N_9146,N_9033,N_9030);
nand U9147 (N_9147,N_9016,N_9083);
nor U9148 (N_9148,N_9010,N_9059);
or U9149 (N_9149,N_9062,N_9036);
or U9150 (N_9150,N_9093,N_9037);
or U9151 (N_9151,N_9086,N_9093);
xnor U9152 (N_9152,N_9077,N_9022);
nand U9153 (N_9153,N_9021,N_9010);
and U9154 (N_9154,N_9052,N_9098);
nand U9155 (N_9155,N_9039,N_9062);
nor U9156 (N_9156,N_9087,N_9065);
nor U9157 (N_9157,N_9081,N_9022);
nand U9158 (N_9158,N_9033,N_9075);
and U9159 (N_9159,N_9021,N_9098);
and U9160 (N_9160,N_9068,N_9044);
or U9161 (N_9161,N_9066,N_9051);
nor U9162 (N_9162,N_9043,N_9097);
or U9163 (N_9163,N_9046,N_9010);
nor U9164 (N_9164,N_9034,N_9092);
and U9165 (N_9165,N_9038,N_9008);
xor U9166 (N_9166,N_9088,N_9018);
or U9167 (N_9167,N_9048,N_9047);
or U9168 (N_9168,N_9045,N_9080);
nor U9169 (N_9169,N_9046,N_9091);
or U9170 (N_9170,N_9076,N_9041);
nand U9171 (N_9171,N_9029,N_9030);
or U9172 (N_9172,N_9022,N_9065);
or U9173 (N_9173,N_9025,N_9007);
xnor U9174 (N_9174,N_9005,N_9028);
nor U9175 (N_9175,N_9065,N_9017);
nand U9176 (N_9176,N_9020,N_9035);
or U9177 (N_9177,N_9030,N_9028);
nand U9178 (N_9178,N_9069,N_9062);
or U9179 (N_9179,N_9041,N_9088);
xor U9180 (N_9180,N_9055,N_9076);
xor U9181 (N_9181,N_9026,N_9018);
nor U9182 (N_9182,N_9075,N_9047);
nor U9183 (N_9183,N_9047,N_9090);
or U9184 (N_9184,N_9018,N_9037);
nand U9185 (N_9185,N_9070,N_9030);
xnor U9186 (N_9186,N_9059,N_9072);
xnor U9187 (N_9187,N_9056,N_9021);
or U9188 (N_9188,N_9043,N_9047);
or U9189 (N_9189,N_9010,N_9054);
nor U9190 (N_9190,N_9046,N_9017);
xor U9191 (N_9191,N_9067,N_9077);
or U9192 (N_9192,N_9044,N_9022);
nor U9193 (N_9193,N_9084,N_9047);
and U9194 (N_9194,N_9000,N_9004);
nor U9195 (N_9195,N_9075,N_9035);
nand U9196 (N_9196,N_9044,N_9075);
xnor U9197 (N_9197,N_9070,N_9076);
nor U9198 (N_9198,N_9015,N_9087);
or U9199 (N_9199,N_9073,N_9009);
and U9200 (N_9200,N_9132,N_9181);
nor U9201 (N_9201,N_9178,N_9164);
nand U9202 (N_9202,N_9190,N_9130);
and U9203 (N_9203,N_9148,N_9172);
and U9204 (N_9204,N_9146,N_9161);
or U9205 (N_9205,N_9145,N_9105);
nor U9206 (N_9206,N_9117,N_9183);
and U9207 (N_9207,N_9127,N_9100);
and U9208 (N_9208,N_9138,N_9174);
or U9209 (N_9209,N_9124,N_9166);
or U9210 (N_9210,N_9159,N_9133);
xor U9211 (N_9211,N_9151,N_9142);
nand U9212 (N_9212,N_9162,N_9179);
and U9213 (N_9213,N_9186,N_9171);
or U9214 (N_9214,N_9184,N_9197);
nand U9215 (N_9215,N_9180,N_9147);
nand U9216 (N_9216,N_9199,N_9177);
nor U9217 (N_9217,N_9118,N_9152);
nand U9218 (N_9218,N_9192,N_9125);
or U9219 (N_9219,N_9135,N_9113);
and U9220 (N_9220,N_9128,N_9139);
nor U9221 (N_9221,N_9110,N_9168);
nand U9222 (N_9222,N_9182,N_9119);
and U9223 (N_9223,N_9191,N_9116);
nor U9224 (N_9224,N_9144,N_9150);
and U9225 (N_9225,N_9131,N_9167);
and U9226 (N_9226,N_9189,N_9104);
nand U9227 (N_9227,N_9187,N_9103);
xor U9228 (N_9228,N_9165,N_9156);
and U9229 (N_9229,N_9195,N_9112);
nand U9230 (N_9230,N_9196,N_9153);
nand U9231 (N_9231,N_9137,N_9170);
nand U9232 (N_9232,N_9173,N_9102);
nand U9233 (N_9233,N_9107,N_9108);
and U9234 (N_9234,N_9134,N_9169);
or U9235 (N_9235,N_9193,N_9111);
xnor U9236 (N_9236,N_9176,N_9157);
or U9237 (N_9237,N_9120,N_9185);
xor U9238 (N_9238,N_9198,N_9194);
or U9239 (N_9239,N_9114,N_9154);
xnor U9240 (N_9240,N_9122,N_9160);
nor U9241 (N_9241,N_9188,N_9123);
xor U9242 (N_9242,N_9175,N_9141);
nor U9243 (N_9243,N_9155,N_9140);
or U9244 (N_9244,N_9126,N_9101);
and U9245 (N_9245,N_9136,N_9115);
xor U9246 (N_9246,N_9158,N_9106);
nand U9247 (N_9247,N_9143,N_9149);
nand U9248 (N_9248,N_9163,N_9129);
nand U9249 (N_9249,N_9109,N_9121);
nor U9250 (N_9250,N_9184,N_9189);
or U9251 (N_9251,N_9144,N_9182);
and U9252 (N_9252,N_9154,N_9129);
and U9253 (N_9253,N_9147,N_9198);
xor U9254 (N_9254,N_9140,N_9136);
nand U9255 (N_9255,N_9183,N_9148);
nand U9256 (N_9256,N_9139,N_9194);
and U9257 (N_9257,N_9198,N_9133);
xnor U9258 (N_9258,N_9109,N_9142);
xor U9259 (N_9259,N_9133,N_9111);
or U9260 (N_9260,N_9155,N_9176);
nand U9261 (N_9261,N_9190,N_9150);
nor U9262 (N_9262,N_9113,N_9156);
xor U9263 (N_9263,N_9131,N_9182);
or U9264 (N_9264,N_9178,N_9101);
and U9265 (N_9265,N_9185,N_9143);
nor U9266 (N_9266,N_9105,N_9102);
and U9267 (N_9267,N_9198,N_9112);
and U9268 (N_9268,N_9170,N_9190);
or U9269 (N_9269,N_9179,N_9153);
and U9270 (N_9270,N_9125,N_9129);
nand U9271 (N_9271,N_9152,N_9127);
nor U9272 (N_9272,N_9146,N_9172);
nand U9273 (N_9273,N_9192,N_9156);
or U9274 (N_9274,N_9167,N_9149);
or U9275 (N_9275,N_9114,N_9186);
nand U9276 (N_9276,N_9136,N_9116);
nand U9277 (N_9277,N_9119,N_9108);
xnor U9278 (N_9278,N_9187,N_9108);
and U9279 (N_9279,N_9105,N_9131);
xnor U9280 (N_9280,N_9113,N_9131);
nor U9281 (N_9281,N_9130,N_9148);
nor U9282 (N_9282,N_9120,N_9105);
and U9283 (N_9283,N_9143,N_9162);
and U9284 (N_9284,N_9107,N_9126);
and U9285 (N_9285,N_9127,N_9104);
xnor U9286 (N_9286,N_9145,N_9196);
or U9287 (N_9287,N_9149,N_9124);
and U9288 (N_9288,N_9151,N_9138);
nand U9289 (N_9289,N_9171,N_9199);
or U9290 (N_9290,N_9150,N_9118);
nand U9291 (N_9291,N_9116,N_9167);
or U9292 (N_9292,N_9146,N_9166);
and U9293 (N_9293,N_9129,N_9171);
nor U9294 (N_9294,N_9111,N_9187);
xnor U9295 (N_9295,N_9110,N_9166);
or U9296 (N_9296,N_9117,N_9171);
xor U9297 (N_9297,N_9109,N_9175);
xor U9298 (N_9298,N_9194,N_9179);
nand U9299 (N_9299,N_9101,N_9139);
nor U9300 (N_9300,N_9283,N_9236);
or U9301 (N_9301,N_9284,N_9253);
nand U9302 (N_9302,N_9299,N_9252);
nor U9303 (N_9303,N_9200,N_9229);
xor U9304 (N_9304,N_9263,N_9235);
and U9305 (N_9305,N_9297,N_9246);
or U9306 (N_9306,N_9226,N_9222);
nand U9307 (N_9307,N_9260,N_9230);
nor U9308 (N_9308,N_9291,N_9245);
and U9309 (N_9309,N_9287,N_9276);
and U9310 (N_9310,N_9261,N_9247);
nand U9311 (N_9311,N_9286,N_9242);
xor U9312 (N_9312,N_9214,N_9201);
nor U9313 (N_9313,N_9266,N_9249);
nand U9314 (N_9314,N_9233,N_9218);
nand U9315 (N_9315,N_9219,N_9264);
nand U9316 (N_9316,N_9231,N_9204);
xnor U9317 (N_9317,N_9290,N_9248);
xor U9318 (N_9318,N_9280,N_9238);
xnor U9319 (N_9319,N_9279,N_9209);
xor U9320 (N_9320,N_9221,N_9271);
and U9321 (N_9321,N_9289,N_9203);
nand U9322 (N_9322,N_9267,N_9211);
nor U9323 (N_9323,N_9216,N_9295);
nor U9324 (N_9324,N_9225,N_9293);
nor U9325 (N_9325,N_9240,N_9262);
nor U9326 (N_9326,N_9215,N_9288);
nor U9327 (N_9327,N_9298,N_9296);
nor U9328 (N_9328,N_9208,N_9255);
nor U9329 (N_9329,N_9207,N_9241);
or U9330 (N_9330,N_9244,N_9237);
nand U9331 (N_9331,N_9213,N_9275);
nand U9332 (N_9332,N_9270,N_9282);
nor U9333 (N_9333,N_9281,N_9227);
and U9334 (N_9334,N_9212,N_9251);
and U9335 (N_9335,N_9217,N_9265);
and U9336 (N_9336,N_9232,N_9223);
or U9337 (N_9337,N_9224,N_9272);
or U9338 (N_9338,N_9254,N_9258);
nand U9339 (N_9339,N_9228,N_9202);
xor U9340 (N_9340,N_9239,N_9220);
and U9341 (N_9341,N_9285,N_9294);
nand U9342 (N_9342,N_9250,N_9257);
nor U9343 (N_9343,N_9259,N_9206);
or U9344 (N_9344,N_9277,N_9273);
nand U9345 (N_9345,N_9256,N_9278);
or U9346 (N_9346,N_9274,N_9234);
nor U9347 (N_9347,N_9210,N_9292);
nand U9348 (N_9348,N_9269,N_9205);
or U9349 (N_9349,N_9268,N_9243);
nand U9350 (N_9350,N_9255,N_9247);
or U9351 (N_9351,N_9258,N_9299);
nor U9352 (N_9352,N_9204,N_9214);
or U9353 (N_9353,N_9259,N_9277);
or U9354 (N_9354,N_9237,N_9207);
xnor U9355 (N_9355,N_9270,N_9230);
or U9356 (N_9356,N_9290,N_9282);
and U9357 (N_9357,N_9246,N_9288);
nor U9358 (N_9358,N_9265,N_9216);
nand U9359 (N_9359,N_9215,N_9217);
nor U9360 (N_9360,N_9249,N_9289);
and U9361 (N_9361,N_9256,N_9210);
nand U9362 (N_9362,N_9222,N_9216);
or U9363 (N_9363,N_9284,N_9249);
nand U9364 (N_9364,N_9260,N_9226);
xnor U9365 (N_9365,N_9242,N_9234);
xor U9366 (N_9366,N_9286,N_9224);
or U9367 (N_9367,N_9232,N_9269);
and U9368 (N_9368,N_9285,N_9226);
and U9369 (N_9369,N_9218,N_9282);
nor U9370 (N_9370,N_9205,N_9276);
nor U9371 (N_9371,N_9218,N_9281);
xnor U9372 (N_9372,N_9243,N_9263);
nor U9373 (N_9373,N_9222,N_9225);
xor U9374 (N_9374,N_9220,N_9223);
and U9375 (N_9375,N_9267,N_9230);
nand U9376 (N_9376,N_9281,N_9216);
nand U9377 (N_9377,N_9204,N_9227);
or U9378 (N_9378,N_9215,N_9247);
nor U9379 (N_9379,N_9276,N_9216);
and U9380 (N_9380,N_9221,N_9297);
and U9381 (N_9381,N_9222,N_9292);
or U9382 (N_9382,N_9214,N_9266);
or U9383 (N_9383,N_9223,N_9227);
or U9384 (N_9384,N_9272,N_9237);
nand U9385 (N_9385,N_9237,N_9248);
xor U9386 (N_9386,N_9238,N_9233);
nand U9387 (N_9387,N_9200,N_9231);
nor U9388 (N_9388,N_9275,N_9240);
and U9389 (N_9389,N_9283,N_9222);
or U9390 (N_9390,N_9270,N_9249);
nand U9391 (N_9391,N_9285,N_9242);
and U9392 (N_9392,N_9262,N_9271);
and U9393 (N_9393,N_9202,N_9236);
xnor U9394 (N_9394,N_9288,N_9285);
nand U9395 (N_9395,N_9276,N_9269);
xor U9396 (N_9396,N_9227,N_9275);
nor U9397 (N_9397,N_9219,N_9254);
nand U9398 (N_9398,N_9266,N_9208);
xnor U9399 (N_9399,N_9206,N_9236);
xor U9400 (N_9400,N_9334,N_9398);
nor U9401 (N_9401,N_9387,N_9377);
or U9402 (N_9402,N_9325,N_9340);
xnor U9403 (N_9403,N_9358,N_9346);
or U9404 (N_9404,N_9338,N_9356);
and U9405 (N_9405,N_9335,N_9360);
xnor U9406 (N_9406,N_9316,N_9369);
nand U9407 (N_9407,N_9310,N_9308);
nor U9408 (N_9408,N_9317,N_9333);
nor U9409 (N_9409,N_9396,N_9330);
or U9410 (N_9410,N_9304,N_9327);
xor U9411 (N_9411,N_9319,N_9375);
and U9412 (N_9412,N_9314,N_9395);
and U9413 (N_9413,N_9382,N_9305);
xnor U9414 (N_9414,N_9370,N_9371);
nand U9415 (N_9415,N_9363,N_9303);
nand U9416 (N_9416,N_9384,N_9353);
and U9417 (N_9417,N_9348,N_9309);
and U9418 (N_9418,N_9328,N_9365);
xnor U9419 (N_9419,N_9343,N_9312);
nand U9420 (N_9420,N_9399,N_9366);
or U9421 (N_9421,N_9393,N_9329);
xor U9422 (N_9422,N_9339,N_9344);
nor U9423 (N_9423,N_9337,N_9379);
nor U9424 (N_9424,N_9342,N_9373);
or U9425 (N_9425,N_9389,N_9347);
or U9426 (N_9426,N_9364,N_9361);
nand U9427 (N_9427,N_9324,N_9311);
nor U9428 (N_9428,N_9367,N_9349);
and U9429 (N_9429,N_9378,N_9397);
and U9430 (N_9430,N_9352,N_9392);
or U9431 (N_9431,N_9318,N_9320);
xor U9432 (N_9432,N_9332,N_9383);
nand U9433 (N_9433,N_9350,N_9381);
nand U9434 (N_9434,N_9321,N_9302);
and U9435 (N_9435,N_9307,N_9390);
nor U9436 (N_9436,N_9362,N_9388);
and U9437 (N_9437,N_9376,N_9301);
nor U9438 (N_9438,N_9300,N_9331);
and U9439 (N_9439,N_9323,N_9394);
and U9440 (N_9440,N_9313,N_9374);
xnor U9441 (N_9441,N_9386,N_9359);
or U9442 (N_9442,N_9357,N_9385);
nand U9443 (N_9443,N_9368,N_9341);
nor U9444 (N_9444,N_9322,N_9372);
nor U9445 (N_9445,N_9355,N_9380);
nor U9446 (N_9446,N_9345,N_9354);
xnor U9447 (N_9447,N_9306,N_9351);
or U9448 (N_9448,N_9391,N_9315);
xor U9449 (N_9449,N_9336,N_9326);
nand U9450 (N_9450,N_9315,N_9308);
xnor U9451 (N_9451,N_9331,N_9347);
and U9452 (N_9452,N_9342,N_9362);
or U9453 (N_9453,N_9355,N_9359);
nor U9454 (N_9454,N_9348,N_9354);
nand U9455 (N_9455,N_9304,N_9381);
and U9456 (N_9456,N_9340,N_9367);
nor U9457 (N_9457,N_9386,N_9348);
nand U9458 (N_9458,N_9341,N_9396);
nand U9459 (N_9459,N_9366,N_9360);
or U9460 (N_9460,N_9392,N_9315);
nor U9461 (N_9461,N_9300,N_9354);
or U9462 (N_9462,N_9342,N_9392);
xnor U9463 (N_9463,N_9389,N_9340);
and U9464 (N_9464,N_9343,N_9356);
or U9465 (N_9465,N_9322,N_9341);
nand U9466 (N_9466,N_9317,N_9373);
and U9467 (N_9467,N_9392,N_9363);
xor U9468 (N_9468,N_9307,N_9326);
nor U9469 (N_9469,N_9326,N_9390);
xor U9470 (N_9470,N_9372,N_9356);
nand U9471 (N_9471,N_9384,N_9327);
xor U9472 (N_9472,N_9378,N_9382);
nand U9473 (N_9473,N_9392,N_9395);
and U9474 (N_9474,N_9351,N_9348);
nor U9475 (N_9475,N_9316,N_9301);
nand U9476 (N_9476,N_9345,N_9395);
and U9477 (N_9477,N_9375,N_9301);
nor U9478 (N_9478,N_9354,N_9395);
xor U9479 (N_9479,N_9330,N_9383);
nand U9480 (N_9480,N_9342,N_9321);
nand U9481 (N_9481,N_9350,N_9369);
and U9482 (N_9482,N_9309,N_9336);
xor U9483 (N_9483,N_9399,N_9348);
xor U9484 (N_9484,N_9396,N_9328);
xnor U9485 (N_9485,N_9327,N_9347);
and U9486 (N_9486,N_9369,N_9348);
nand U9487 (N_9487,N_9370,N_9340);
nor U9488 (N_9488,N_9344,N_9386);
xor U9489 (N_9489,N_9363,N_9366);
nor U9490 (N_9490,N_9365,N_9300);
and U9491 (N_9491,N_9321,N_9365);
nor U9492 (N_9492,N_9362,N_9338);
xor U9493 (N_9493,N_9388,N_9315);
or U9494 (N_9494,N_9325,N_9355);
xor U9495 (N_9495,N_9369,N_9330);
or U9496 (N_9496,N_9398,N_9354);
and U9497 (N_9497,N_9331,N_9369);
nor U9498 (N_9498,N_9387,N_9312);
xnor U9499 (N_9499,N_9306,N_9393);
xor U9500 (N_9500,N_9411,N_9429);
and U9501 (N_9501,N_9497,N_9453);
and U9502 (N_9502,N_9465,N_9489);
nor U9503 (N_9503,N_9435,N_9441);
xnor U9504 (N_9504,N_9461,N_9443);
nand U9505 (N_9505,N_9424,N_9417);
xor U9506 (N_9506,N_9472,N_9456);
or U9507 (N_9507,N_9496,N_9408);
or U9508 (N_9508,N_9467,N_9415);
and U9509 (N_9509,N_9402,N_9422);
and U9510 (N_9510,N_9482,N_9430);
or U9511 (N_9511,N_9477,N_9499);
nor U9512 (N_9512,N_9451,N_9440);
nor U9513 (N_9513,N_9475,N_9471);
nand U9514 (N_9514,N_9474,N_9442);
nand U9515 (N_9515,N_9473,N_9436);
xor U9516 (N_9516,N_9407,N_9405);
or U9517 (N_9517,N_9487,N_9438);
xnor U9518 (N_9518,N_9437,N_9463);
xnor U9519 (N_9519,N_9455,N_9427);
xnor U9520 (N_9520,N_9412,N_9485);
nor U9521 (N_9521,N_9469,N_9431);
nand U9522 (N_9522,N_9428,N_9498);
xnor U9523 (N_9523,N_9462,N_9448);
xnor U9524 (N_9524,N_9464,N_9468);
and U9525 (N_9525,N_9452,N_9490);
and U9526 (N_9526,N_9434,N_9400);
or U9527 (N_9527,N_9491,N_9479);
nand U9528 (N_9528,N_9493,N_9419);
nor U9529 (N_9529,N_9421,N_9433);
or U9530 (N_9530,N_9406,N_9480);
or U9531 (N_9531,N_9416,N_9439);
or U9532 (N_9532,N_9483,N_9481);
or U9533 (N_9533,N_9418,N_9450);
and U9534 (N_9534,N_9495,N_9447);
nand U9535 (N_9535,N_9449,N_9488);
nand U9536 (N_9536,N_9454,N_9457);
nor U9537 (N_9537,N_9410,N_9444);
nand U9538 (N_9538,N_9403,N_9486);
and U9539 (N_9539,N_9420,N_9492);
or U9540 (N_9540,N_9466,N_9476);
nor U9541 (N_9541,N_9425,N_9426);
xnor U9542 (N_9542,N_9458,N_9414);
nand U9543 (N_9543,N_9409,N_9459);
nand U9544 (N_9544,N_9445,N_9484);
or U9545 (N_9545,N_9446,N_9423);
xor U9546 (N_9546,N_9460,N_9413);
and U9547 (N_9547,N_9432,N_9404);
or U9548 (N_9548,N_9494,N_9401);
nand U9549 (N_9549,N_9478,N_9470);
xnor U9550 (N_9550,N_9474,N_9478);
or U9551 (N_9551,N_9405,N_9483);
xor U9552 (N_9552,N_9442,N_9400);
and U9553 (N_9553,N_9447,N_9476);
and U9554 (N_9554,N_9429,N_9422);
and U9555 (N_9555,N_9455,N_9437);
xnor U9556 (N_9556,N_9497,N_9479);
xnor U9557 (N_9557,N_9451,N_9411);
nand U9558 (N_9558,N_9416,N_9438);
and U9559 (N_9559,N_9401,N_9418);
and U9560 (N_9560,N_9411,N_9420);
and U9561 (N_9561,N_9468,N_9412);
xnor U9562 (N_9562,N_9453,N_9476);
or U9563 (N_9563,N_9472,N_9498);
or U9564 (N_9564,N_9458,N_9472);
nand U9565 (N_9565,N_9497,N_9443);
and U9566 (N_9566,N_9467,N_9458);
nand U9567 (N_9567,N_9440,N_9412);
nor U9568 (N_9568,N_9434,N_9418);
nand U9569 (N_9569,N_9464,N_9471);
xnor U9570 (N_9570,N_9419,N_9468);
xor U9571 (N_9571,N_9481,N_9405);
nor U9572 (N_9572,N_9439,N_9404);
and U9573 (N_9573,N_9454,N_9424);
xor U9574 (N_9574,N_9496,N_9430);
nor U9575 (N_9575,N_9435,N_9404);
or U9576 (N_9576,N_9413,N_9463);
xor U9577 (N_9577,N_9419,N_9430);
xor U9578 (N_9578,N_9471,N_9496);
and U9579 (N_9579,N_9432,N_9450);
nand U9580 (N_9580,N_9443,N_9495);
or U9581 (N_9581,N_9440,N_9483);
xnor U9582 (N_9582,N_9471,N_9434);
or U9583 (N_9583,N_9409,N_9451);
nor U9584 (N_9584,N_9426,N_9400);
nor U9585 (N_9585,N_9425,N_9435);
xnor U9586 (N_9586,N_9481,N_9458);
xor U9587 (N_9587,N_9444,N_9420);
nand U9588 (N_9588,N_9457,N_9428);
and U9589 (N_9589,N_9497,N_9417);
and U9590 (N_9590,N_9498,N_9406);
nor U9591 (N_9591,N_9481,N_9482);
nor U9592 (N_9592,N_9434,N_9402);
or U9593 (N_9593,N_9498,N_9416);
nand U9594 (N_9594,N_9420,N_9407);
nor U9595 (N_9595,N_9450,N_9442);
and U9596 (N_9596,N_9492,N_9464);
or U9597 (N_9597,N_9473,N_9491);
or U9598 (N_9598,N_9475,N_9435);
or U9599 (N_9599,N_9469,N_9483);
xnor U9600 (N_9600,N_9515,N_9560);
and U9601 (N_9601,N_9591,N_9597);
or U9602 (N_9602,N_9594,N_9502);
nor U9603 (N_9603,N_9583,N_9525);
nor U9604 (N_9604,N_9599,N_9568);
nand U9605 (N_9605,N_9545,N_9500);
xor U9606 (N_9606,N_9553,N_9596);
or U9607 (N_9607,N_9576,N_9524);
and U9608 (N_9608,N_9547,N_9561);
nand U9609 (N_9609,N_9587,N_9536);
and U9610 (N_9610,N_9510,N_9556);
xor U9611 (N_9611,N_9578,N_9552);
or U9612 (N_9612,N_9546,N_9528);
xnor U9613 (N_9613,N_9532,N_9521);
xor U9614 (N_9614,N_9529,N_9539);
and U9615 (N_9615,N_9555,N_9505);
and U9616 (N_9616,N_9562,N_9574);
nor U9617 (N_9617,N_9540,N_9589);
nand U9618 (N_9618,N_9571,N_9542);
or U9619 (N_9619,N_9509,N_9581);
or U9620 (N_9620,N_9541,N_9549);
and U9621 (N_9621,N_9586,N_9523);
nor U9622 (N_9622,N_9550,N_9557);
nor U9623 (N_9623,N_9580,N_9531);
and U9624 (N_9624,N_9534,N_9585);
xor U9625 (N_9625,N_9584,N_9554);
nor U9626 (N_9626,N_9513,N_9519);
or U9627 (N_9627,N_9564,N_9592);
nand U9628 (N_9628,N_9511,N_9503);
nor U9629 (N_9629,N_9544,N_9501);
nand U9630 (N_9630,N_9563,N_9543);
and U9631 (N_9631,N_9535,N_9506);
nand U9632 (N_9632,N_9514,N_9572);
and U9633 (N_9633,N_9567,N_9512);
nand U9634 (N_9634,N_9504,N_9559);
xor U9635 (N_9635,N_9533,N_9538);
or U9636 (N_9636,N_9537,N_9566);
and U9637 (N_9637,N_9573,N_9595);
nand U9638 (N_9638,N_9579,N_9558);
and U9639 (N_9639,N_9530,N_9520);
xor U9640 (N_9640,N_9507,N_9526);
or U9641 (N_9641,N_9516,N_9548);
nor U9642 (N_9642,N_9527,N_9522);
xor U9643 (N_9643,N_9598,N_9551);
xnor U9644 (N_9644,N_9517,N_9575);
xor U9645 (N_9645,N_9590,N_9582);
and U9646 (N_9646,N_9577,N_9588);
nand U9647 (N_9647,N_9565,N_9570);
and U9648 (N_9648,N_9593,N_9569);
xnor U9649 (N_9649,N_9518,N_9508);
and U9650 (N_9650,N_9532,N_9592);
nand U9651 (N_9651,N_9523,N_9507);
or U9652 (N_9652,N_9573,N_9596);
or U9653 (N_9653,N_9589,N_9560);
and U9654 (N_9654,N_9557,N_9544);
nand U9655 (N_9655,N_9530,N_9535);
or U9656 (N_9656,N_9548,N_9576);
and U9657 (N_9657,N_9523,N_9551);
nor U9658 (N_9658,N_9508,N_9516);
or U9659 (N_9659,N_9553,N_9556);
nand U9660 (N_9660,N_9566,N_9519);
and U9661 (N_9661,N_9500,N_9594);
nor U9662 (N_9662,N_9546,N_9575);
or U9663 (N_9663,N_9571,N_9556);
xnor U9664 (N_9664,N_9585,N_9527);
and U9665 (N_9665,N_9596,N_9502);
nand U9666 (N_9666,N_9509,N_9578);
xnor U9667 (N_9667,N_9590,N_9595);
and U9668 (N_9668,N_9588,N_9595);
nand U9669 (N_9669,N_9538,N_9532);
and U9670 (N_9670,N_9549,N_9584);
nand U9671 (N_9671,N_9504,N_9508);
nand U9672 (N_9672,N_9554,N_9536);
xnor U9673 (N_9673,N_9586,N_9504);
and U9674 (N_9674,N_9576,N_9536);
nand U9675 (N_9675,N_9591,N_9561);
nand U9676 (N_9676,N_9514,N_9509);
xnor U9677 (N_9677,N_9539,N_9566);
or U9678 (N_9678,N_9581,N_9548);
or U9679 (N_9679,N_9519,N_9535);
and U9680 (N_9680,N_9575,N_9567);
and U9681 (N_9681,N_9557,N_9541);
nor U9682 (N_9682,N_9515,N_9545);
or U9683 (N_9683,N_9596,N_9589);
and U9684 (N_9684,N_9524,N_9574);
and U9685 (N_9685,N_9512,N_9568);
xor U9686 (N_9686,N_9512,N_9587);
nand U9687 (N_9687,N_9550,N_9508);
nand U9688 (N_9688,N_9525,N_9577);
nor U9689 (N_9689,N_9525,N_9559);
and U9690 (N_9690,N_9587,N_9509);
or U9691 (N_9691,N_9536,N_9572);
and U9692 (N_9692,N_9592,N_9575);
nor U9693 (N_9693,N_9518,N_9589);
or U9694 (N_9694,N_9564,N_9517);
nor U9695 (N_9695,N_9567,N_9559);
or U9696 (N_9696,N_9532,N_9566);
and U9697 (N_9697,N_9530,N_9594);
or U9698 (N_9698,N_9564,N_9540);
or U9699 (N_9699,N_9542,N_9556);
nand U9700 (N_9700,N_9681,N_9625);
nor U9701 (N_9701,N_9617,N_9606);
nor U9702 (N_9702,N_9640,N_9602);
or U9703 (N_9703,N_9646,N_9654);
or U9704 (N_9704,N_9665,N_9688);
nand U9705 (N_9705,N_9686,N_9635);
nor U9706 (N_9706,N_9611,N_9669);
xnor U9707 (N_9707,N_9614,N_9643);
nand U9708 (N_9708,N_9687,N_9607);
or U9709 (N_9709,N_9622,N_9631);
and U9710 (N_9710,N_9673,N_9629);
nor U9711 (N_9711,N_9676,N_9632);
nand U9712 (N_9712,N_9671,N_9601);
or U9713 (N_9713,N_9609,N_9684);
nor U9714 (N_9714,N_9698,N_9668);
xnor U9715 (N_9715,N_9634,N_9695);
and U9716 (N_9716,N_9645,N_9618);
nor U9717 (N_9717,N_9610,N_9628);
and U9718 (N_9718,N_9664,N_9678);
nand U9719 (N_9719,N_9600,N_9692);
xnor U9720 (N_9720,N_9689,N_9694);
nor U9721 (N_9721,N_9624,N_9620);
xor U9722 (N_9722,N_9660,N_9697);
nand U9723 (N_9723,N_9612,N_9693);
xor U9724 (N_9724,N_9648,N_9642);
nand U9725 (N_9725,N_9655,N_9649);
xnor U9726 (N_9726,N_9650,N_9653);
nor U9727 (N_9727,N_9623,N_9644);
nand U9728 (N_9728,N_9696,N_9621);
and U9729 (N_9729,N_9675,N_9604);
xor U9730 (N_9730,N_9652,N_9605);
nor U9731 (N_9731,N_9674,N_9633);
nor U9732 (N_9732,N_9690,N_9627);
nor U9733 (N_9733,N_9657,N_9685);
xnor U9734 (N_9734,N_9616,N_9682);
or U9735 (N_9735,N_9658,N_9680);
or U9736 (N_9736,N_9647,N_9699);
nand U9737 (N_9737,N_9670,N_9608);
or U9738 (N_9738,N_9691,N_9613);
or U9739 (N_9739,N_9603,N_9637);
nor U9740 (N_9740,N_9638,N_9667);
or U9741 (N_9741,N_9677,N_9661);
nand U9742 (N_9742,N_9626,N_9641);
and U9743 (N_9743,N_9639,N_9615);
and U9744 (N_9744,N_9672,N_9662);
nand U9745 (N_9745,N_9663,N_9636);
nor U9746 (N_9746,N_9679,N_9619);
nor U9747 (N_9747,N_9683,N_9659);
nor U9748 (N_9748,N_9651,N_9656);
nand U9749 (N_9749,N_9630,N_9666);
nand U9750 (N_9750,N_9647,N_9605);
and U9751 (N_9751,N_9601,N_9646);
xnor U9752 (N_9752,N_9644,N_9637);
nor U9753 (N_9753,N_9601,N_9657);
nor U9754 (N_9754,N_9694,N_9605);
or U9755 (N_9755,N_9680,N_9608);
or U9756 (N_9756,N_9612,N_9603);
and U9757 (N_9757,N_9695,N_9611);
nand U9758 (N_9758,N_9679,N_9608);
and U9759 (N_9759,N_9655,N_9691);
or U9760 (N_9760,N_9642,N_9680);
and U9761 (N_9761,N_9665,N_9652);
nor U9762 (N_9762,N_9671,N_9632);
or U9763 (N_9763,N_9621,N_9666);
or U9764 (N_9764,N_9629,N_9616);
nand U9765 (N_9765,N_9659,N_9613);
xnor U9766 (N_9766,N_9665,N_9691);
xnor U9767 (N_9767,N_9674,N_9653);
nand U9768 (N_9768,N_9659,N_9697);
nor U9769 (N_9769,N_9605,N_9625);
or U9770 (N_9770,N_9664,N_9625);
or U9771 (N_9771,N_9647,N_9640);
or U9772 (N_9772,N_9619,N_9638);
and U9773 (N_9773,N_9689,N_9624);
and U9774 (N_9774,N_9668,N_9691);
or U9775 (N_9775,N_9681,N_9657);
nand U9776 (N_9776,N_9607,N_9643);
and U9777 (N_9777,N_9667,N_9609);
or U9778 (N_9778,N_9605,N_9688);
nor U9779 (N_9779,N_9613,N_9615);
or U9780 (N_9780,N_9692,N_9663);
xnor U9781 (N_9781,N_9604,N_9636);
nor U9782 (N_9782,N_9602,N_9660);
xnor U9783 (N_9783,N_9686,N_9650);
or U9784 (N_9784,N_9607,N_9637);
nor U9785 (N_9785,N_9608,N_9601);
or U9786 (N_9786,N_9604,N_9619);
nor U9787 (N_9787,N_9654,N_9695);
nor U9788 (N_9788,N_9603,N_9656);
and U9789 (N_9789,N_9675,N_9688);
xnor U9790 (N_9790,N_9618,N_9668);
or U9791 (N_9791,N_9699,N_9657);
or U9792 (N_9792,N_9605,N_9613);
xnor U9793 (N_9793,N_9612,N_9658);
nor U9794 (N_9794,N_9671,N_9695);
and U9795 (N_9795,N_9613,N_9646);
or U9796 (N_9796,N_9613,N_9642);
nand U9797 (N_9797,N_9646,N_9665);
or U9798 (N_9798,N_9665,N_9677);
nor U9799 (N_9799,N_9699,N_9606);
xnor U9800 (N_9800,N_9772,N_9708);
nand U9801 (N_9801,N_9742,N_9705);
or U9802 (N_9802,N_9728,N_9718);
nand U9803 (N_9803,N_9716,N_9725);
nand U9804 (N_9804,N_9738,N_9791);
and U9805 (N_9805,N_9789,N_9750);
or U9806 (N_9806,N_9798,N_9799);
nand U9807 (N_9807,N_9731,N_9763);
and U9808 (N_9808,N_9745,N_9777);
nand U9809 (N_9809,N_9704,N_9736);
xnor U9810 (N_9810,N_9709,N_9711);
or U9811 (N_9811,N_9747,N_9755);
or U9812 (N_9812,N_9788,N_9743);
nand U9813 (N_9813,N_9758,N_9715);
and U9814 (N_9814,N_9761,N_9720);
nor U9815 (N_9815,N_9723,N_9767);
or U9816 (N_9816,N_9754,N_9768);
nand U9817 (N_9817,N_9714,N_9737);
and U9818 (N_9818,N_9762,N_9775);
or U9819 (N_9819,N_9757,N_9719);
and U9820 (N_9820,N_9700,N_9751);
xor U9821 (N_9821,N_9796,N_9786);
nand U9822 (N_9822,N_9780,N_9733);
nand U9823 (N_9823,N_9722,N_9741);
and U9824 (N_9824,N_9753,N_9769);
nand U9825 (N_9825,N_9774,N_9779);
or U9826 (N_9826,N_9721,N_9794);
or U9827 (N_9827,N_9703,N_9782);
nand U9828 (N_9828,N_9702,N_9776);
nand U9829 (N_9829,N_9710,N_9744);
and U9830 (N_9830,N_9793,N_9783);
xor U9831 (N_9831,N_9740,N_9727);
or U9832 (N_9832,N_9781,N_9766);
and U9833 (N_9833,N_9726,N_9792);
nand U9834 (N_9834,N_9729,N_9701);
and U9835 (N_9835,N_9752,N_9734);
and U9836 (N_9836,N_9773,N_9797);
xor U9837 (N_9837,N_9756,N_9778);
nor U9838 (N_9838,N_9712,N_9785);
xor U9839 (N_9839,N_9784,N_9748);
nor U9840 (N_9840,N_9707,N_9717);
nand U9841 (N_9841,N_9746,N_9760);
xnor U9842 (N_9842,N_9759,N_9770);
nor U9843 (N_9843,N_9724,N_9730);
xor U9844 (N_9844,N_9706,N_9787);
nor U9845 (N_9845,N_9732,N_9713);
and U9846 (N_9846,N_9771,N_9795);
nor U9847 (N_9847,N_9790,N_9764);
xnor U9848 (N_9848,N_9735,N_9765);
nand U9849 (N_9849,N_9739,N_9749);
nor U9850 (N_9850,N_9711,N_9790);
nand U9851 (N_9851,N_9731,N_9761);
nor U9852 (N_9852,N_9778,N_9753);
or U9853 (N_9853,N_9765,N_9781);
or U9854 (N_9854,N_9786,N_9739);
nor U9855 (N_9855,N_9766,N_9783);
and U9856 (N_9856,N_9781,N_9779);
nand U9857 (N_9857,N_9714,N_9708);
or U9858 (N_9858,N_9721,N_9725);
or U9859 (N_9859,N_9716,N_9724);
nand U9860 (N_9860,N_9740,N_9737);
or U9861 (N_9861,N_9770,N_9712);
or U9862 (N_9862,N_9730,N_9764);
nor U9863 (N_9863,N_9794,N_9762);
nor U9864 (N_9864,N_9798,N_9730);
and U9865 (N_9865,N_9742,N_9771);
nand U9866 (N_9866,N_9777,N_9778);
or U9867 (N_9867,N_9795,N_9736);
nor U9868 (N_9868,N_9742,N_9766);
nand U9869 (N_9869,N_9792,N_9796);
nand U9870 (N_9870,N_9730,N_9729);
or U9871 (N_9871,N_9767,N_9781);
or U9872 (N_9872,N_9733,N_9755);
xnor U9873 (N_9873,N_9720,N_9786);
nand U9874 (N_9874,N_9751,N_9790);
and U9875 (N_9875,N_9759,N_9760);
or U9876 (N_9876,N_9765,N_9711);
nand U9877 (N_9877,N_9744,N_9767);
and U9878 (N_9878,N_9793,N_9709);
nand U9879 (N_9879,N_9795,N_9722);
nand U9880 (N_9880,N_9724,N_9784);
and U9881 (N_9881,N_9729,N_9734);
and U9882 (N_9882,N_9724,N_9729);
nand U9883 (N_9883,N_9741,N_9763);
xor U9884 (N_9884,N_9753,N_9771);
nor U9885 (N_9885,N_9712,N_9739);
nand U9886 (N_9886,N_9782,N_9722);
and U9887 (N_9887,N_9743,N_9732);
nand U9888 (N_9888,N_9737,N_9780);
or U9889 (N_9889,N_9735,N_9726);
and U9890 (N_9890,N_9701,N_9798);
or U9891 (N_9891,N_9709,N_9733);
nor U9892 (N_9892,N_9706,N_9762);
xnor U9893 (N_9893,N_9705,N_9757);
xnor U9894 (N_9894,N_9760,N_9755);
xnor U9895 (N_9895,N_9742,N_9738);
or U9896 (N_9896,N_9739,N_9732);
nor U9897 (N_9897,N_9705,N_9709);
or U9898 (N_9898,N_9785,N_9780);
and U9899 (N_9899,N_9794,N_9755);
nor U9900 (N_9900,N_9874,N_9834);
or U9901 (N_9901,N_9886,N_9807);
nand U9902 (N_9902,N_9820,N_9833);
nand U9903 (N_9903,N_9832,N_9880);
nor U9904 (N_9904,N_9811,N_9873);
xor U9905 (N_9905,N_9803,N_9854);
and U9906 (N_9906,N_9868,N_9867);
xor U9907 (N_9907,N_9809,N_9890);
or U9908 (N_9908,N_9876,N_9887);
nor U9909 (N_9909,N_9877,N_9851);
nor U9910 (N_9910,N_9821,N_9826);
or U9911 (N_9911,N_9825,N_9899);
and U9912 (N_9912,N_9848,N_9841);
xor U9913 (N_9913,N_9802,N_9853);
xor U9914 (N_9914,N_9801,N_9804);
or U9915 (N_9915,N_9823,N_9837);
or U9916 (N_9916,N_9893,N_9842);
nor U9917 (N_9917,N_9816,N_9845);
or U9918 (N_9918,N_9828,N_9818);
and U9919 (N_9919,N_9835,N_9831);
nor U9920 (N_9920,N_9819,N_9849);
xor U9921 (N_9921,N_9856,N_9895);
or U9922 (N_9922,N_9838,N_9896);
or U9923 (N_9923,N_9817,N_9883);
nand U9924 (N_9924,N_9829,N_9822);
nand U9925 (N_9925,N_9824,N_9894);
nand U9926 (N_9926,N_9875,N_9800);
nand U9927 (N_9927,N_9806,N_9839);
nand U9928 (N_9928,N_9861,N_9898);
and U9929 (N_9929,N_9855,N_9870);
xor U9930 (N_9930,N_9885,N_9852);
xnor U9931 (N_9931,N_9827,N_9888);
or U9932 (N_9932,N_9863,N_9815);
and U9933 (N_9933,N_9850,N_9860);
xnor U9934 (N_9934,N_9812,N_9872);
nor U9935 (N_9935,N_9881,N_9884);
and U9936 (N_9936,N_9889,N_9805);
or U9937 (N_9937,N_9840,N_9871);
nor U9938 (N_9938,N_9866,N_9892);
and U9939 (N_9939,N_9836,N_9865);
and U9940 (N_9940,N_9882,N_9847);
nor U9941 (N_9941,N_9864,N_9897);
xnor U9942 (N_9942,N_9813,N_9858);
or U9943 (N_9943,N_9862,N_9843);
nand U9944 (N_9944,N_9830,N_9844);
and U9945 (N_9945,N_9808,N_9859);
nor U9946 (N_9946,N_9878,N_9869);
or U9947 (N_9947,N_9814,N_9857);
nand U9948 (N_9948,N_9891,N_9879);
nor U9949 (N_9949,N_9810,N_9846);
or U9950 (N_9950,N_9834,N_9859);
nand U9951 (N_9951,N_9880,N_9895);
nor U9952 (N_9952,N_9866,N_9821);
and U9953 (N_9953,N_9888,N_9834);
nor U9954 (N_9954,N_9858,N_9817);
or U9955 (N_9955,N_9863,N_9860);
and U9956 (N_9956,N_9868,N_9878);
nor U9957 (N_9957,N_9856,N_9809);
or U9958 (N_9958,N_9828,N_9849);
xnor U9959 (N_9959,N_9805,N_9820);
nor U9960 (N_9960,N_9861,N_9852);
xor U9961 (N_9961,N_9881,N_9825);
nor U9962 (N_9962,N_9852,N_9838);
xor U9963 (N_9963,N_9862,N_9874);
nand U9964 (N_9964,N_9852,N_9867);
nor U9965 (N_9965,N_9808,N_9893);
xnor U9966 (N_9966,N_9814,N_9848);
nand U9967 (N_9967,N_9858,N_9845);
xnor U9968 (N_9968,N_9845,N_9879);
nand U9969 (N_9969,N_9862,N_9838);
and U9970 (N_9970,N_9805,N_9852);
and U9971 (N_9971,N_9841,N_9886);
nand U9972 (N_9972,N_9850,N_9874);
nand U9973 (N_9973,N_9860,N_9883);
nand U9974 (N_9974,N_9830,N_9810);
and U9975 (N_9975,N_9878,N_9886);
xnor U9976 (N_9976,N_9839,N_9867);
nor U9977 (N_9977,N_9839,N_9817);
nor U9978 (N_9978,N_9841,N_9891);
xor U9979 (N_9979,N_9879,N_9892);
xnor U9980 (N_9980,N_9805,N_9878);
nand U9981 (N_9981,N_9829,N_9882);
and U9982 (N_9982,N_9848,N_9800);
xnor U9983 (N_9983,N_9832,N_9820);
nor U9984 (N_9984,N_9892,N_9813);
nand U9985 (N_9985,N_9861,N_9886);
xnor U9986 (N_9986,N_9838,N_9836);
nand U9987 (N_9987,N_9889,N_9820);
and U9988 (N_9988,N_9819,N_9882);
nand U9989 (N_9989,N_9838,N_9827);
nand U9990 (N_9990,N_9861,N_9883);
nand U9991 (N_9991,N_9887,N_9840);
nand U9992 (N_9992,N_9839,N_9842);
nor U9993 (N_9993,N_9805,N_9834);
and U9994 (N_9994,N_9863,N_9856);
and U9995 (N_9995,N_9884,N_9844);
xor U9996 (N_9996,N_9859,N_9883);
and U9997 (N_9997,N_9812,N_9868);
xnor U9998 (N_9998,N_9822,N_9891);
or U9999 (N_9999,N_9854,N_9816);
nor UO_0 (O_0,N_9958,N_9938);
nand UO_1 (O_1,N_9956,N_9922);
or UO_2 (O_2,N_9909,N_9972);
nor UO_3 (O_3,N_9919,N_9921);
or UO_4 (O_4,N_9910,N_9994);
nor UO_5 (O_5,N_9961,N_9997);
xor UO_6 (O_6,N_9964,N_9966);
xor UO_7 (O_7,N_9944,N_9977);
or UO_8 (O_8,N_9960,N_9904);
nand UO_9 (O_9,N_9980,N_9978);
and UO_10 (O_10,N_9992,N_9962);
nand UO_11 (O_11,N_9989,N_9941);
or UO_12 (O_12,N_9914,N_9987);
nor UO_13 (O_13,N_9949,N_9990);
xnor UO_14 (O_14,N_9940,N_9999);
nand UO_15 (O_15,N_9985,N_9952);
or UO_16 (O_16,N_9953,N_9973);
nand UO_17 (O_17,N_9975,N_9937);
or UO_18 (O_18,N_9974,N_9923);
or UO_19 (O_19,N_9955,N_9943);
or UO_20 (O_20,N_9933,N_9959);
or UO_21 (O_21,N_9942,N_9979);
xnor UO_22 (O_22,N_9911,N_9947);
nand UO_23 (O_23,N_9946,N_9932);
and UO_24 (O_24,N_9954,N_9945);
nand UO_25 (O_25,N_9948,N_9920);
xor UO_26 (O_26,N_9928,N_9902);
and UO_27 (O_27,N_9982,N_9931);
nand UO_28 (O_28,N_9924,N_9930);
nand UO_29 (O_29,N_9901,N_9917);
nand UO_30 (O_30,N_9950,N_9984);
nand UO_31 (O_31,N_9935,N_9936);
xor UO_32 (O_32,N_9963,N_9995);
xor UO_33 (O_33,N_9900,N_9988);
nor UO_34 (O_34,N_9971,N_9957);
and UO_35 (O_35,N_9993,N_9912);
or UO_36 (O_36,N_9996,N_9986);
nand UO_37 (O_37,N_9929,N_9991);
or UO_38 (O_38,N_9906,N_9998);
xor UO_39 (O_39,N_9967,N_9907);
and UO_40 (O_40,N_9927,N_9926);
or UO_41 (O_41,N_9918,N_9915);
nand UO_42 (O_42,N_9939,N_9965);
and UO_43 (O_43,N_9981,N_9913);
nand UO_44 (O_44,N_9970,N_9925);
and UO_45 (O_45,N_9905,N_9968);
or UO_46 (O_46,N_9983,N_9976);
and UO_47 (O_47,N_9969,N_9951);
nand UO_48 (O_48,N_9903,N_9916);
nand UO_49 (O_49,N_9934,N_9908);
xnor UO_50 (O_50,N_9921,N_9941);
or UO_51 (O_51,N_9900,N_9974);
xnor UO_52 (O_52,N_9975,N_9993);
xnor UO_53 (O_53,N_9930,N_9945);
nor UO_54 (O_54,N_9973,N_9923);
nand UO_55 (O_55,N_9982,N_9949);
xor UO_56 (O_56,N_9920,N_9940);
nor UO_57 (O_57,N_9927,N_9956);
xnor UO_58 (O_58,N_9988,N_9998);
nand UO_59 (O_59,N_9928,N_9948);
xor UO_60 (O_60,N_9976,N_9937);
or UO_61 (O_61,N_9901,N_9908);
or UO_62 (O_62,N_9994,N_9996);
or UO_63 (O_63,N_9962,N_9923);
xor UO_64 (O_64,N_9936,N_9937);
nand UO_65 (O_65,N_9922,N_9993);
nor UO_66 (O_66,N_9974,N_9958);
and UO_67 (O_67,N_9961,N_9901);
xor UO_68 (O_68,N_9938,N_9925);
nand UO_69 (O_69,N_9941,N_9931);
nor UO_70 (O_70,N_9908,N_9935);
nand UO_71 (O_71,N_9990,N_9905);
nor UO_72 (O_72,N_9949,N_9993);
xor UO_73 (O_73,N_9981,N_9967);
xnor UO_74 (O_74,N_9952,N_9938);
or UO_75 (O_75,N_9935,N_9953);
and UO_76 (O_76,N_9946,N_9919);
nand UO_77 (O_77,N_9984,N_9936);
nand UO_78 (O_78,N_9968,N_9923);
nand UO_79 (O_79,N_9937,N_9902);
or UO_80 (O_80,N_9998,N_9971);
and UO_81 (O_81,N_9979,N_9971);
xor UO_82 (O_82,N_9960,N_9993);
and UO_83 (O_83,N_9904,N_9905);
nor UO_84 (O_84,N_9953,N_9958);
nand UO_85 (O_85,N_9923,N_9926);
nand UO_86 (O_86,N_9929,N_9908);
nor UO_87 (O_87,N_9961,N_9928);
or UO_88 (O_88,N_9948,N_9993);
or UO_89 (O_89,N_9923,N_9959);
xnor UO_90 (O_90,N_9996,N_9918);
nand UO_91 (O_91,N_9949,N_9945);
and UO_92 (O_92,N_9997,N_9991);
xnor UO_93 (O_93,N_9924,N_9942);
nor UO_94 (O_94,N_9943,N_9947);
and UO_95 (O_95,N_9944,N_9953);
nor UO_96 (O_96,N_9924,N_9907);
nand UO_97 (O_97,N_9962,N_9928);
or UO_98 (O_98,N_9914,N_9932);
nor UO_99 (O_99,N_9985,N_9931);
nand UO_100 (O_100,N_9915,N_9920);
nor UO_101 (O_101,N_9933,N_9975);
nor UO_102 (O_102,N_9927,N_9914);
xor UO_103 (O_103,N_9960,N_9980);
xor UO_104 (O_104,N_9953,N_9906);
nand UO_105 (O_105,N_9969,N_9968);
xnor UO_106 (O_106,N_9980,N_9985);
nor UO_107 (O_107,N_9916,N_9940);
nand UO_108 (O_108,N_9981,N_9950);
or UO_109 (O_109,N_9979,N_9937);
nand UO_110 (O_110,N_9940,N_9984);
or UO_111 (O_111,N_9945,N_9986);
xor UO_112 (O_112,N_9959,N_9948);
nand UO_113 (O_113,N_9938,N_9989);
or UO_114 (O_114,N_9986,N_9902);
or UO_115 (O_115,N_9992,N_9931);
or UO_116 (O_116,N_9920,N_9979);
or UO_117 (O_117,N_9921,N_9994);
or UO_118 (O_118,N_9935,N_9909);
nor UO_119 (O_119,N_9957,N_9913);
xnor UO_120 (O_120,N_9986,N_9943);
or UO_121 (O_121,N_9970,N_9905);
or UO_122 (O_122,N_9945,N_9955);
nor UO_123 (O_123,N_9988,N_9986);
nand UO_124 (O_124,N_9976,N_9997);
and UO_125 (O_125,N_9983,N_9921);
or UO_126 (O_126,N_9911,N_9960);
or UO_127 (O_127,N_9981,N_9998);
nor UO_128 (O_128,N_9985,N_9911);
or UO_129 (O_129,N_9977,N_9988);
xnor UO_130 (O_130,N_9960,N_9954);
and UO_131 (O_131,N_9998,N_9964);
xnor UO_132 (O_132,N_9945,N_9935);
nand UO_133 (O_133,N_9924,N_9936);
nor UO_134 (O_134,N_9939,N_9990);
nand UO_135 (O_135,N_9992,N_9957);
nor UO_136 (O_136,N_9974,N_9919);
nor UO_137 (O_137,N_9977,N_9930);
nand UO_138 (O_138,N_9952,N_9901);
nand UO_139 (O_139,N_9974,N_9924);
nand UO_140 (O_140,N_9964,N_9925);
nor UO_141 (O_141,N_9903,N_9905);
and UO_142 (O_142,N_9935,N_9991);
nand UO_143 (O_143,N_9965,N_9930);
and UO_144 (O_144,N_9958,N_9903);
or UO_145 (O_145,N_9933,N_9979);
xor UO_146 (O_146,N_9998,N_9955);
nor UO_147 (O_147,N_9937,N_9956);
or UO_148 (O_148,N_9934,N_9958);
nand UO_149 (O_149,N_9950,N_9995);
nor UO_150 (O_150,N_9964,N_9968);
nor UO_151 (O_151,N_9981,N_9978);
nand UO_152 (O_152,N_9928,N_9915);
nor UO_153 (O_153,N_9912,N_9932);
or UO_154 (O_154,N_9912,N_9982);
and UO_155 (O_155,N_9945,N_9988);
nor UO_156 (O_156,N_9984,N_9917);
xnor UO_157 (O_157,N_9984,N_9951);
and UO_158 (O_158,N_9990,N_9981);
nand UO_159 (O_159,N_9930,N_9946);
and UO_160 (O_160,N_9967,N_9915);
and UO_161 (O_161,N_9928,N_9971);
nor UO_162 (O_162,N_9911,N_9954);
or UO_163 (O_163,N_9930,N_9914);
nor UO_164 (O_164,N_9987,N_9926);
nor UO_165 (O_165,N_9906,N_9911);
nand UO_166 (O_166,N_9909,N_9986);
xor UO_167 (O_167,N_9981,N_9919);
or UO_168 (O_168,N_9953,N_9927);
and UO_169 (O_169,N_9988,N_9961);
nand UO_170 (O_170,N_9904,N_9983);
nor UO_171 (O_171,N_9901,N_9904);
and UO_172 (O_172,N_9976,N_9929);
nor UO_173 (O_173,N_9943,N_9905);
xor UO_174 (O_174,N_9955,N_9916);
nand UO_175 (O_175,N_9923,N_9984);
nor UO_176 (O_176,N_9901,N_9987);
nor UO_177 (O_177,N_9910,N_9978);
nand UO_178 (O_178,N_9964,N_9973);
nand UO_179 (O_179,N_9991,N_9968);
or UO_180 (O_180,N_9928,N_9963);
and UO_181 (O_181,N_9946,N_9979);
and UO_182 (O_182,N_9934,N_9918);
nor UO_183 (O_183,N_9948,N_9978);
nor UO_184 (O_184,N_9949,N_9980);
xnor UO_185 (O_185,N_9924,N_9965);
nand UO_186 (O_186,N_9971,N_9949);
and UO_187 (O_187,N_9987,N_9956);
nand UO_188 (O_188,N_9993,N_9910);
nor UO_189 (O_189,N_9989,N_9967);
nand UO_190 (O_190,N_9990,N_9934);
and UO_191 (O_191,N_9982,N_9925);
and UO_192 (O_192,N_9905,N_9967);
nand UO_193 (O_193,N_9983,N_9908);
nand UO_194 (O_194,N_9904,N_9957);
and UO_195 (O_195,N_9938,N_9960);
nand UO_196 (O_196,N_9962,N_9929);
or UO_197 (O_197,N_9909,N_9908);
nor UO_198 (O_198,N_9927,N_9912);
or UO_199 (O_199,N_9982,N_9926);
nand UO_200 (O_200,N_9937,N_9957);
nand UO_201 (O_201,N_9952,N_9935);
and UO_202 (O_202,N_9923,N_9907);
nand UO_203 (O_203,N_9987,N_9932);
or UO_204 (O_204,N_9917,N_9927);
and UO_205 (O_205,N_9943,N_9929);
or UO_206 (O_206,N_9945,N_9901);
and UO_207 (O_207,N_9946,N_9988);
nor UO_208 (O_208,N_9992,N_9952);
nor UO_209 (O_209,N_9939,N_9955);
xnor UO_210 (O_210,N_9966,N_9996);
nand UO_211 (O_211,N_9966,N_9959);
or UO_212 (O_212,N_9943,N_9989);
xor UO_213 (O_213,N_9921,N_9974);
nor UO_214 (O_214,N_9929,N_9928);
or UO_215 (O_215,N_9994,N_9919);
or UO_216 (O_216,N_9976,N_9980);
nor UO_217 (O_217,N_9957,N_9954);
xnor UO_218 (O_218,N_9985,N_9913);
nor UO_219 (O_219,N_9975,N_9935);
and UO_220 (O_220,N_9923,N_9966);
and UO_221 (O_221,N_9955,N_9947);
xnor UO_222 (O_222,N_9976,N_9918);
nand UO_223 (O_223,N_9989,N_9958);
xnor UO_224 (O_224,N_9980,N_9937);
or UO_225 (O_225,N_9993,N_9995);
xnor UO_226 (O_226,N_9992,N_9902);
or UO_227 (O_227,N_9915,N_9960);
nand UO_228 (O_228,N_9900,N_9964);
nor UO_229 (O_229,N_9904,N_9924);
nand UO_230 (O_230,N_9957,N_9960);
nand UO_231 (O_231,N_9933,N_9944);
nor UO_232 (O_232,N_9974,N_9942);
and UO_233 (O_233,N_9917,N_9918);
or UO_234 (O_234,N_9950,N_9919);
nor UO_235 (O_235,N_9926,N_9973);
nor UO_236 (O_236,N_9996,N_9910);
nor UO_237 (O_237,N_9968,N_9917);
nand UO_238 (O_238,N_9989,N_9937);
xnor UO_239 (O_239,N_9964,N_9989);
or UO_240 (O_240,N_9912,N_9980);
or UO_241 (O_241,N_9989,N_9981);
nor UO_242 (O_242,N_9914,N_9965);
nand UO_243 (O_243,N_9970,N_9921);
or UO_244 (O_244,N_9989,N_9992);
and UO_245 (O_245,N_9914,N_9976);
xor UO_246 (O_246,N_9998,N_9905);
xor UO_247 (O_247,N_9944,N_9986);
nor UO_248 (O_248,N_9905,N_9972);
nand UO_249 (O_249,N_9916,N_9911);
nand UO_250 (O_250,N_9989,N_9935);
or UO_251 (O_251,N_9904,N_9913);
and UO_252 (O_252,N_9903,N_9918);
and UO_253 (O_253,N_9924,N_9975);
or UO_254 (O_254,N_9930,N_9979);
nor UO_255 (O_255,N_9928,N_9957);
xor UO_256 (O_256,N_9955,N_9972);
xor UO_257 (O_257,N_9937,N_9977);
or UO_258 (O_258,N_9938,N_9976);
and UO_259 (O_259,N_9952,N_9931);
or UO_260 (O_260,N_9929,N_9914);
or UO_261 (O_261,N_9953,N_9997);
or UO_262 (O_262,N_9900,N_9922);
nand UO_263 (O_263,N_9976,N_9954);
or UO_264 (O_264,N_9965,N_9913);
and UO_265 (O_265,N_9956,N_9992);
and UO_266 (O_266,N_9912,N_9931);
xnor UO_267 (O_267,N_9940,N_9943);
and UO_268 (O_268,N_9969,N_9996);
and UO_269 (O_269,N_9962,N_9969);
nor UO_270 (O_270,N_9927,N_9936);
and UO_271 (O_271,N_9946,N_9992);
nand UO_272 (O_272,N_9919,N_9942);
nand UO_273 (O_273,N_9934,N_9970);
nand UO_274 (O_274,N_9914,N_9921);
or UO_275 (O_275,N_9993,N_9931);
nor UO_276 (O_276,N_9992,N_9993);
or UO_277 (O_277,N_9972,N_9900);
or UO_278 (O_278,N_9957,N_9910);
nor UO_279 (O_279,N_9909,N_9904);
nand UO_280 (O_280,N_9978,N_9983);
xor UO_281 (O_281,N_9918,N_9912);
nand UO_282 (O_282,N_9912,N_9967);
and UO_283 (O_283,N_9922,N_9980);
nand UO_284 (O_284,N_9990,N_9969);
xnor UO_285 (O_285,N_9952,N_9941);
nand UO_286 (O_286,N_9910,N_9975);
or UO_287 (O_287,N_9920,N_9974);
and UO_288 (O_288,N_9959,N_9978);
nor UO_289 (O_289,N_9940,N_9949);
or UO_290 (O_290,N_9910,N_9953);
and UO_291 (O_291,N_9948,N_9941);
and UO_292 (O_292,N_9997,N_9913);
or UO_293 (O_293,N_9994,N_9955);
and UO_294 (O_294,N_9955,N_9922);
nand UO_295 (O_295,N_9930,N_9919);
xor UO_296 (O_296,N_9977,N_9975);
nor UO_297 (O_297,N_9942,N_9918);
nor UO_298 (O_298,N_9953,N_9952);
nor UO_299 (O_299,N_9968,N_9944);
and UO_300 (O_300,N_9996,N_9982);
and UO_301 (O_301,N_9988,N_9962);
nor UO_302 (O_302,N_9977,N_9954);
or UO_303 (O_303,N_9943,N_9907);
and UO_304 (O_304,N_9910,N_9959);
nand UO_305 (O_305,N_9981,N_9961);
or UO_306 (O_306,N_9986,N_9920);
nor UO_307 (O_307,N_9953,N_9922);
nand UO_308 (O_308,N_9909,N_9954);
nand UO_309 (O_309,N_9958,N_9956);
or UO_310 (O_310,N_9976,N_9993);
or UO_311 (O_311,N_9912,N_9942);
xnor UO_312 (O_312,N_9955,N_9912);
or UO_313 (O_313,N_9926,N_9934);
and UO_314 (O_314,N_9957,N_9959);
xnor UO_315 (O_315,N_9921,N_9999);
nand UO_316 (O_316,N_9961,N_9979);
nand UO_317 (O_317,N_9986,N_9917);
or UO_318 (O_318,N_9966,N_9962);
nand UO_319 (O_319,N_9987,N_9905);
and UO_320 (O_320,N_9998,N_9951);
and UO_321 (O_321,N_9955,N_9960);
nor UO_322 (O_322,N_9944,N_9950);
nor UO_323 (O_323,N_9925,N_9921);
xor UO_324 (O_324,N_9963,N_9965);
or UO_325 (O_325,N_9912,N_9994);
nand UO_326 (O_326,N_9955,N_9999);
or UO_327 (O_327,N_9972,N_9929);
or UO_328 (O_328,N_9931,N_9942);
nand UO_329 (O_329,N_9980,N_9963);
nor UO_330 (O_330,N_9992,N_9912);
xor UO_331 (O_331,N_9935,N_9901);
and UO_332 (O_332,N_9937,N_9965);
and UO_333 (O_333,N_9998,N_9900);
nor UO_334 (O_334,N_9930,N_9909);
xnor UO_335 (O_335,N_9944,N_9985);
and UO_336 (O_336,N_9904,N_9907);
xnor UO_337 (O_337,N_9905,N_9928);
and UO_338 (O_338,N_9941,N_9903);
xnor UO_339 (O_339,N_9967,N_9926);
and UO_340 (O_340,N_9914,N_9955);
or UO_341 (O_341,N_9912,N_9904);
nand UO_342 (O_342,N_9936,N_9921);
and UO_343 (O_343,N_9975,N_9932);
or UO_344 (O_344,N_9907,N_9964);
xnor UO_345 (O_345,N_9910,N_9937);
nor UO_346 (O_346,N_9923,N_9902);
xnor UO_347 (O_347,N_9914,N_9992);
nand UO_348 (O_348,N_9924,N_9948);
or UO_349 (O_349,N_9926,N_9918);
nand UO_350 (O_350,N_9902,N_9910);
nand UO_351 (O_351,N_9930,N_9989);
nand UO_352 (O_352,N_9965,N_9952);
xnor UO_353 (O_353,N_9975,N_9954);
nor UO_354 (O_354,N_9982,N_9971);
nor UO_355 (O_355,N_9963,N_9903);
or UO_356 (O_356,N_9937,N_9966);
nand UO_357 (O_357,N_9910,N_9917);
nor UO_358 (O_358,N_9923,N_9919);
or UO_359 (O_359,N_9947,N_9935);
and UO_360 (O_360,N_9976,N_9999);
and UO_361 (O_361,N_9986,N_9911);
or UO_362 (O_362,N_9937,N_9932);
nand UO_363 (O_363,N_9951,N_9968);
or UO_364 (O_364,N_9999,N_9905);
xor UO_365 (O_365,N_9940,N_9955);
nor UO_366 (O_366,N_9999,N_9992);
xor UO_367 (O_367,N_9945,N_9906);
or UO_368 (O_368,N_9929,N_9935);
nor UO_369 (O_369,N_9928,N_9993);
and UO_370 (O_370,N_9923,N_9957);
xor UO_371 (O_371,N_9952,N_9951);
and UO_372 (O_372,N_9998,N_9974);
or UO_373 (O_373,N_9921,N_9951);
nor UO_374 (O_374,N_9928,N_9974);
and UO_375 (O_375,N_9920,N_9926);
nor UO_376 (O_376,N_9925,N_9992);
xnor UO_377 (O_377,N_9946,N_9940);
or UO_378 (O_378,N_9941,N_9913);
nand UO_379 (O_379,N_9946,N_9948);
or UO_380 (O_380,N_9950,N_9903);
xor UO_381 (O_381,N_9991,N_9999);
and UO_382 (O_382,N_9991,N_9986);
nand UO_383 (O_383,N_9910,N_9921);
or UO_384 (O_384,N_9949,N_9953);
nand UO_385 (O_385,N_9935,N_9910);
or UO_386 (O_386,N_9929,N_9905);
and UO_387 (O_387,N_9955,N_9975);
xnor UO_388 (O_388,N_9991,N_9921);
xor UO_389 (O_389,N_9997,N_9921);
nor UO_390 (O_390,N_9951,N_9973);
nand UO_391 (O_391,N_9948,N_9970);
nand UO_392 (O_392,N_9987,N_9924);
or UO_393 (O_393,N_9992,N_9977);
or UO_394 (O_394,N_9954,N_9993);
nor UO_395 (O_395,N_9992,N_9927);
nand UO_396 (O_396,N_9976,N_9989);
or UO_397 (O_397,N_9902,N_9987);
nand UO_398 (O_398,N_9991,N_9983);
xor UO_399 (O_399,N_9972,N_9937);
xnor UO_400 (O_400,N_9960,N_9931);
xnor UO_401 (O_401,N_9941,N_9957);
xnor UO_402 (O_402,N_9993,N_9914);
and UO_403 (O_403,N_9992,N_9995);
and UO_404 (O_404,N_9952,N_9939);
nor UO_405 (O_405,N_9968,N_9943);
xnor UO_406 (O_406,N_9951,N_9918);
or UO_407 (O_407,N_9904,N_9959);
or UO_408 (O_408,N_9925,N_9933);
nor UO_409 (O_409,N_9946,N_9928);
nand UO_410 (O_410,N_9990,N_9968);
nand UO_411 (O_411,N_9920,N_9959);
and UO_412 (O_412,N_9905,N_9906);
nand UO_413 (O_413,N_9930,N_9956);
or UO_414 (O_414,N_9986,N_9929);
or UO_415 (O_415,N_9923,N_9975);
nor UO_416 (O_416,N_9913,N_9938);
or UO_417 (O_417,N_9941,N_9995);
nand UO_418 (O_418,N_9962,N_9931);
nor UO_419 (O_419,N_9961,N_9995);
and UO_420 (O_420,N_9993,N_9998);
nor UO_421 (O_421,N_9963,N_9947);
nor UO_422 (O_422,N_9915,N_9965);
or UO_423 (O_423,N_9968,N_9976);
and UO_424 (O_424,N_9923,N_9988);
nand UO_425 (O_425,N_9946,N_9993);
nor UO_426 (O_426,N_9946,N_9968);
nor UO_427 (O_427,N_9976,N_9904);
and UO_428 (O_428,N_9954,N_9928);
xnor UO_429 (O_429,N_9961,N_9987);
and UO_430 (O_430,N_9966,N_9978);
nor UO_431 (O_431,N_9902,N_9921);
nand UO_432 (O_432,N_9971,N_9910);
xnor UO_433 (O_433,N_9924,N_9940);
or UO_434 (O_434,N_9995,N_9982);
or UO_435 (O_435,N_9963,N_9940);
nand UO_436 (O_436,N_9996,N_9903);
nand UO_437 (O_437,N_9913,N_9900);
nand UO_438 (O_438,N_9944,N_9943);
nand UO_439 (O_439,N_9990,N_9920);
and UO_440 (O_440,N_9933,N_9962);
nand UO_441 (O_441,N_9962,N_9968);
nor UO_442 (O_442,N_9952,N_9976);
xnor UO_443 (O_443,N_9905,N_9952);
nand UO_444 (O_444,N_9958,N_9900);
and UO_445 (O_445,N_9985,N_9949);
nand UO_446 (O_446,N_9938,N_9980);
nor UO_447 (O_447,N_9917,N_9938);
or UO_448 (O_448,N_9983,N_9975);
nand UO_449 (O_449,N_9940,N_9952);
nand UO_450 (O_450,N_9992,N_9909);
nand UO_451 (O_451,N_9944,N_9964);
xnor UO_452 (O_452,N_9974,N_9938);
xnor UO_453 (O_453,N_9970,N_9936);
nor UO_454 (O_454,N_9935,N_9993);
nor UO_455 (O_455,N_9958,N_9921);
nand UO_456 (O_456,N_9953,N_9971);
nor UO_457 (O_457,N_9935,N_9964);
and UO_458 (O_458,N_9978,N_9956);
nor UO_459 (O_459,N_9956,N_9983);
and UO_460 (O_460,N_9924,N_9921);
xnor UO_461 (O_461,N_9991,N_9907);
nor UO_462 (O_462,N_9961,N_9906);
and UO_463 (O_463,N_9962,N_9965);
nand UO_464 (O_464,N_9929,N_9900);
xor UO_465 (O_465,N_9941,N_9925);
xor UO_466 (O_466,N_9970,N_9965);
and UO_467 (O_467,N_9921,N_9926);
xor UO_468 (O_468,N_9922,N_9931);
and UO_469 (O_469,N_9933,N_9913);
nand UO_470 (O_470,N_9966,N_9912);
xor UO_471 (O_471,N_9964,N_9965);
xor UO_472 (O_472,N_9966,N_9908);
nor UO_473 (O_473,N_9925,N_9908);
nand UO_474 (O_474,N_9919,N_9983);
or UO_475 (O_475,N_9960,N_9912);
or UO_476 (O_476,N_9942,N_9908);
or UO_477 (O_477,N_9932,N_9972);
nand UO_478 (O_478,N_9961,N_9927);
nor UO_479 (O_479,N_9914,N_9952);
and UO_480 (O_480,N_9919,N_9987);
and UO_481 (O_481,N_9939,N_9932);
and UO_482 (O_482,N_9915,N_9964);
xor UO_483 (O_483,N_9948,N_9935);
nor UO_484 (O_484,N_9916,N_9923);
and UO_485 (O_485,N_9958,N_9968);
xnor UO_486 (O_486,N_9955,N_9954);
or UO_487 (O_487,N_9947,N_9903);
xnor UO_488 (O_488,N_9948,N_9963);
nand UO_489 (O_489,N_9921,N_9938);
and UO_490 (O_490,N_9969,N_9973);
nor UO_491 (O_491,N_9976,N_9936);
nand UO_492 (O_492,N_9903,N_9966);
or UO_493 (O_493,N_9966,N_9990);
or UO_494 (O_494,N_9931,N_9943);
and UO_495 (O_495,N_9981,N_9900);
xnor UO_496 (O_496,N_9925,N_9943);
xor UO_497 (O_497,N_9947,N_9931);
xor UO_498 (O_498,N_9998,N_9917);
or UO_499 (O_499,N_9985,N_9973);
or UO_500 (O_500,N_9997,N_9972);
and UO_501 (O_501,N_9991,N_9994);
xor UO_502 (O_502,N_9933,N_9936);
xnor UO_503 (O_503,N_9947,N_9989);
nand UO_504 (O_504,N_9910,N_9970);
and UO_505 (O_505,N_9972,N_9926);
xnor UO_506 (O_506,N_9972,N_9991);
xnor UO_507 (O_507,N_9911,N_9921);
xnor UO_508 (O_508,N_9977,N_9980);
nand UO_509 (O_509,N_9954,N_9901);
nor UO_510 (O_510,N_9945,N_9942);
or UO_511 (O_511,N_9914,N_9960);
nand UO_512 (O_512,N_9918,N_9923);
nor UO_513 (O_513,N_9994,N_9943);
nor UO_514 (O_514,N_9986,N_9922);
xor UO_515 (O_515,N_9978,N_9907);
and UO_516 (O_516,N_9996,N_9952);
nor UO_517 (O_517,N_9939,N_9973);
nor UO_518 (O_518,N_9948,N_9958);
nor UO_519 (O_519,N_9914,N_9988);
xnor UO_520 (O_520,N_9971,N_9951);
nand UO_521 (O_521,N_9966,N_9957);
or UO_522 (O_522,N_9924,N_9934);
nor UO_523 (O_523,N_9956,N_9969);
or UO_524 (O_524,N_9941,N_9922);
or UO_525 (O_525,N_9943,N_9950);
nand UO_526 (O_526,N_9990,N_9928);
xnor UO_527 (O_527,N_9991,N_9917);
or UO_528 (O_528,N_9931,N_9964);
and UO_529 (O_529,N_9975,N_9906);
and UO_530 (O_530,N_9996,N_9953);
and UO_531 (O_531,N_9942,N_9986);
nand UO_532 (O_532,N_9933,N_9932);
nand UO_533 (O_533,N_9922,N_9969);
nand UO_534 (O_534,N_9922,N_9913);
nor UO_535 (O_535,N_9997,N_9912);
or UO_536 (O_536,N_9941,N_9901);
or UO_537 (O_537,N_9966,N_9979);
and UO_538 (O_538,N_9900,N_9950);
or UO_539 (O_539,N_9946,N_9900);
or UO_540 (O_540,N_9979,N_9931);
or UO_541 (O_541,N_9927,N_9976);
and UO_542 (O_542,N_9963,N_9930);
nand UO_543 (O_543,N_9967,N_9909);
xnor UO_544 (O_544,N_9904,N_9953);
nor UO_545 (O_545,N_9909,N_9987);
nand UO_546 (O_546,N_9975,N_9980);
nand UO_547 (O_547,N_9946,N_9995);
nand UO_548 (O_548,N_9977,N_9948);
nor UO_549 (O_549,N_9949,N_9901);
nor UO_550 (O_550,N_9953,N_9916);
nand UO_551 (O_551,N_9942,N_9960);
nand UO_552 (O_552,N_9963,N_9993);
and UO_553 (O_553,N_9937,N_9940);
xor UO_554 (O_554,N_9909,N_9917);
nor UO_555 (O_555,N_9948,N_9974);
xnor UO_556 (O_556,N_9973,N_9932);
or UO_557 (O_557,N_9927,N_9921);
nor UO_558 (O_558,N_9962,N_9922);
or UO_559 (O_559,N_9913,N_9992);
or UO_560 (O_560,N_9991,N_9950);
nand UO_561 (O_561,N_9938,N_9911);
xnor UO_562 (O_562,N_9984,N_9904);
nand UO_563 (O_563,N_9906,N_9974);
or UO_564 (O_564,N_9992,N_9986);
or UO_565 (O_565,N_9935,N_9998);
nor UO_566 (O_566,N_9943,N_9938);
and UO_567 (O_567,N_9947,N_9940);
nand UO_568 (O_568,N_9978,N_9994);
or UO_569 (O_569,N_9957,N_9975);
nand UO_570 (O_570,N_9966,N_9945);
and UO_571 (O_571,N_9983,N_9920);
or UO_572 (O_572,N_9980,N_9969);
xor UO_573 (O_573,N_9987,N_9930);
or UO_574 (O_574,N_9981,N_9975);
nand UO_575 (O_575,N_9986,N_9963);
or UO_576 (O_576,N_9914,N_9973);
and UO_577 (O_577,N_9951,N_9963);
and UO_578 (O_578,N_9983,N_9951);
nor UO_579 (O_579,N_9997,N_9998);
and UO_580 (O_580,N_9918,N_9943);
nand UO_581 (O_581,N_9900,N_9956);
or UO_582 (O_582,N_9918,N_9983);
nand UO_583 (O_583,N_9908,N_9954);
xnor UO_584 (O_584,N_9906,N_9944);
and UO_585 (O_585,N_9916,N_9996);
nand UO_586 (O_586,N_9928,N_9926);
or UO_587 (O_587,N_9905,N_9955);
xnor UO_588 (O_588,N_9914,N_9915);
and UO_589 (O_589,N_9979,N_9949);
xor UO_590 (O_590,N_9999,N_9907);
and UO_591 (O_591,N_9918,N_9905);
or UO_592 (O_592,N_9967,N_9925);
nor UO_593 (O_593,N_9930,N_9991);
or UO_594 (O_594,N_9947,N_9978);
xnor UO_595 (O_595,N_9904,N_9945);
xor UO_596 (O_596,N_9982,N_9965);
or UO_597 (O_597,N_9906,N_9990);
nand UO_598 (O_598,N_9981,N_9916);
xnor UO_599 (O_599,N_9944,N_9916);
xnor UO_600 (O_600,N_9987,N_9988);
and UO_601 (O_601,N_9963,N_9970);
nor UO_602 (O_602,N_9931,N_9920);
and UO_603 (O_603,N_9947,N_9973);
and UO_604 (O_604,N_9947,N_9915);
or UO_605 (O_605,N_9935,N_9932);
xnor UO_606 (O_606,N_9985,N_9936);
and UO_607 (O_607,N_9960,N_9951);
or UO_608 (O_608,N_9983,N_9923);
xor UO_609 (O_609,N_9906,N_9957);
and UO_610 (O_610,N_9991,N_9915);
or UO_611 (O_611,N_9935,N_9927);
and UO_612 (O_612,N_9963,N_9997);
or UO_613 (O_613,N_9974,N_9912);
or UO_614 (O_614,N_9991,N_9952);
nand UO_615 (O_615,N_9933,N_9981);
xor UO_616 (O_616,N_9940,N_9977);
and UO_617 (O_617,N_9993,N_9918);
nor UO_618 (O_618,N_9952,N_9979);
nand UO_619 (O_619,N_9918,N_9970);
nor UO_620 (O_620,N_9927,N_9997);
and UO_621 (O_621,N_9983,N_9966);
and UO_622 (O_622,N_9960,N_9986);
xor UO_623 (O_623,N_9994,N_9949);
nor UO_624 (O_624,N_9944,N_9934);
xor UO_625 (O_625,N_9924,N_9978);
xnor UO_626 (O_626,N_9914,N_9963);
xnor UO_627 (O_627,N_9967,N_9956);
and UO_628 (O_628,N_9919,N_9967);
nor UO_629 (O_629,N_9974,N_9986);
or UO_630 (O_630,N_9921,N_9939);
xor UO_631 (O_631,N_9906,N_9979);
xnor UO_632 (O_632,N_9990,N_9979);
or UO_633 (O_633,N_9905,N_9900);
nor UO_634 (O_634,N_9965,N_9955);
xnor UO_635 (O_635,N_9902,N_9993);
nand UO_636 (O_636,N_9956,N_9945);
nor UO_637 (O_637,N_9904,N_9914);
and UO_638 (O_638,N_9979,N_9993);
nor UO_639 (O_639,N_9908,N_9956);
and UO_640 (O_640,N_9950,N_9930);
xnor UO_641 (O_641,N_9916,N_9932);
nor UO_642 (O_642,N_9916,N_9936);
and UO_643 (O_643,N_9981,N_9936);
xor UO_644 (O_644,N_9959,N_9952);
or UO_645 (O_645,N_9920,N_9966);
and UO_646 (O_646,N_9947,N_9902);
or UO_647 (O_647,N_9955,N_9988);
and UO_648 (O_648,N_9901,N_9938);
and UO_649 (O_649,N_9928,N_9909);
or UO_650 (O_650,N_9919,N_9949);
and UO_651 (O_651,N_9985,N_9946);
or UO_652 (O_652,N_9924,N_9979);
xnor UO_653 (O_653,N_9900,N_9939);
xnor UO_654 (O_654,N_9978,N_9934);
xnor UO_655 (O_655,N_9978,N_9963);
xnor UO_656 (O_656,N_9914,N_9924);
nor UO_657 (O_657,N_9907,N_9973);
xor UO_658 (O_658,N_9992,N_9990);
xor UO_659 (O_659,N_9944,N_9939);
xnor UO_660 (O_660,N_9941,N_9940);
nor UO_661 (O_661,N_9952,N_9932);
or UO_662 (O_662,N_9929,N_9995);
and UO_663 (O_663,N_9939,N_9924);
nor UO_664 (O_664,N_9959,N_9981);
and UO_665 (O_665,N_9974,N_9963);
nand UO_666 (O_666,N_9944,N_9957);
nor UO_667 (O_667,N_9903,N_9972);
xnor UO_668 (O_668,N_9973,N_9934);
nand UO_669 (O_669,N_9976,N_9958);
xnor UO_670 (O_670,N_9937,N_9986);
and UO_671 (O_671,N_9900,N_9987);
xor UO_672 (O_672,N_9979,N_9989);
nand UO_673 (O_673,N_9903,N_9952);
nand UO_674 (O_674,N_9940,N_9996);
or UO_675 (O_675,N_9951,N_9906);
and UO_676 (O_676,N_9918,N_9936);
nand UO_677 (O_677,N_9999,N_9994);
xnor UO_678 (O_678,N_9987,N_9946);
and UO_679 (O_679,N_9935,N_9949);
nand UO_680 (O_680,N_9980,N_9900);
or UO_681 (O_681,N_9984,N_9994);
nor UO_682 (O_682,N_9936,N_9934);
xor UO_683 (O_683,N_9919,N_9962);
nand UO_684 (O_684,N_9994,N_9915);
or UO_685 (O_685,N_9966,N_9938);
nor UO_686 (O_686,N_9998,N_9930);
nand UO_687 (O_687,N_9995,N_9977);
and UO_688 (O_688,N_9995,N_9933);
nor UO_689 (O_689,N_9995,N_9956);
nand UO_690 (O_690,N_9953,N_9993);
or UO_691 (O_691,N_9920,N_9928);
nor UO_692 (O_692,N_9936,N_9986);
nor UO_693 (O_693,N_9912,N_9950);
and UO_694 (O_694,N_9979,N_9955);
and UO_695 (O_695,N_9961,N_9989);
and UO_696 (O_696,N_9905,N_9958);
xnor UO_697 (O_697,N_9927,N_9990);
nand UO_698 (O_698,N_9970,N_9986);
or UO_699 (O_699,N_9932,N_9991);
xor UO_700 (O_700,N_9964,N_9951);
nor UO_701 (O_701,N_9996,N_9913);
nor UO_702 (O_702,N_9910,N_9999);
and UO_703 (O_703,N_9980,N_9911);
or UO_704 (O_704,N_9990,N_9907);
xor UO_705 (O_705,N_9950,N_9904);
or UO_706 (O_706,N_9920,N_9942);
nor UO_707 (O_707,N_9911,N_9924);
nand UO_708 (O_708,N_9923,N_9939);
xor UO_709 (O_709,N_9946,N_9942);
and UO_710 (O_710,N_9979,N_9900);
xor UO_711 (O_711,N_9983,N_9926);
nand UO_712 (O_712,N_9927,N_9905);
nand UO_713 (O_713,N_9912,N_9921);
nor UO_714 (O_714,N_9988,N_9903);
xor UO_715 (O_715,N_9995,N_9907);
or UO_716 (O_716,N_9920,N_9944);
nor UO_717 (O_717,N_9907,N_9996);
xnor UO_718 (O_718,N_9970,N_9946);
xnor UO_719 (O_719,N_9964,N_9916);
and UO_720 (O_720,N_9984,N_9969);
and UO_721 (O_721,N_9955,N_9996);
nand UO_722 (O_722,N_9993,N_9999);
and UO_723 (O_723,N_9957,N_9947);
xor UO_724 (O_724,N_9902,N_9965);
nor UO_725 (O_725,N_9922,N_9907);
and UO_726 (O_726,N_9980,N_9918);
nand UO_727 (O_727,N_9960,N_9962);
xnor UO_728 (O_728,N_9973,N_9952);
or UO_729 (O_729,N_9995,N_9918);
nor UO_730 (O_730,N_9945,N_9921);
nor UO_731 (O_731,N_9912,N_9946);
and UO_732 (O_732,N_9901,N_9998);
nor UO_733 (O_733,N_9941,N_9911);
nand UO_734 (O_734,N_9927,N_9909);
xor UO_735 (O_735,N_9903,N_9946);
or UO_736 (O_736,N_9902,N_9948);
nor UO_737 (O_737,N_9991,N_9901);
nor UO_738 (O_738,N_9976,N_9941);
and UO_739 (O_739,N_9994,N_9972);
and UO_740 (O_740,N_9966,N_9947);
nor UO_741 (O_741,N_9916,N_9947);
xor UO_742 (O_742,N_9967,N_9988);
xnor UO_743 (O_743,N_9959,N_9903);
xnor UO_744 (O_744,N_9915,N_9982);
xnor UO_745 (O_745,N_9927,N_9985);
xnor UO_746 (O_746,N_9935,N_9931);
or UO_747 (O_747,N_9917,N_9954);
nand UO_748 (O_748,N_9923,N_9950);
xnor UO_749 (O_749,N_9952,N_9981);
nor UO_750 (O_750,N_9986,N_9956);
and UO_751 (O_751,N_9923,N_9900);
or UO_752 (O_752,N_9955,N_9987);
nand UO_753 (O_753,N_9915,N_9951);
or UO_754 (O_754,N_9924,N_9969);
nor UO_755 (O_755,N_9985,N_9988);
xor UO_756 (O_756,N_9978,N_9908);
nand UO_757 (O_757,N_9958,N_9952);
nor UO_758 (O_758,N_9907,N_9972);
nand UO_759 (O_759,N_9956,N_9949);
nor UO_760 (O_760,N_9917,N_9999);
and UO_761 (O_761,N_9997,N_9905);
and UO_762 (O_762,N_9968,N_9947);
and UO_763 (O_763,N_9996,N_9959);
and UO_764 (O_764,N_9935,N_9971);
and UO_765 (O_765,N_9984,N_9915);
nand UO_766 (O_766,N_9969,N_9927);
and UO_767 (O_767,N_9943,N_9914);
nand UO_768 (O_768,N_9919,N_9920);
and UO_769 (O_769,N_9946,N_9933);
or UO_770 (O_770,N_9927,N_9907);
nand UO_771 (O_771,N_9925,N_9965);
and UO_772 (O_772,N_9984,N_9902);
or UO_773 (O_773,N_9985,N_9966);
or UO_774 (O_774,N_9921,N_9949);
nand UO_775 (O_775,N_9964,N_9924);
or UO_776 (O_776,N_9925,N_9949);
nand UO_777 (O_777,N_9971,N_9926);
and UO_778 (O_778,N_9910,N_9930);
or UO_779 (O_779,N_9957,N_9998);
and UO_780 (O_780,N_9941,N_9997);
nand UO_781 (O_781,N_9941,N_9994);
nor UO_782 (O_782,N_9930,N_9917);
xor UO_783 (O_783,N_9927,N_9928);
nand UO_784 (O_784,N_9985,N_9926);
and UO_785 (O_785,N_9949,N_9992);
and UO_786 (O_786,N_9909,N_9926);
and UO_787 (O_787,N_9917,N_9943);
and UO_788 (O_788,N_9957,N_9915);
xnor UO_789 (O_789,N_9977,N_9962);
nand UO_790 (O_790,N_9978,N_9952);
or UO_791 (O_791,N_9970,N_9952);
xor UO_792 (O_792,N_9911,N_9946);
nand UO_793 (O_793,N_9944,N_9992);
xnor UO_794 (O_794,N_9926,N_9933);
xor UO_795 (O_795,N_9956,N_9980);
and UO_796 (O_796,N_9959,N_9949);
nor UO_797 (O_797,N_9998,N_9995);
xnor UO_798 (O_798,N_9917,N_9977);
or UO_799 (O_799,N_9945,N_9964);
nand UO_800 (O_800,N_9930,N_9916);
and UO_801 (O_801,N_9943,N_9923);
and UO_802 (O_802,N_9919,N_9903);
xor UO_803 (O_803,N_9944,N_9963);
xor UO_804 (O_804,N_9949,N_9905);
nor UO_805 (O_805,N_9917,N_9994);
or UO_806 (O_806,N_9997,N_9928);
or UO_807 (O_807,N_9954,N_9931);
or UO_808 (O_808,N_9953,N_9985);
and UO_809 (O_809,N_9905,N_9971);
and UO_810 (O_810,N_9997,N_9904);
nand UO_811 (O_811,N_9927,N_9962);
nor UO_812 (O_812,N_9974,N_9917);
or UO_813 (O_813,N_9963,N_9915);
or UO_814 (O_814,N_9902,N_9994);
and UO_815 (O_815,N_9981,N_9905);
xor UO_816 (O_816,N_9969,N_9921);
nand UO_817 (O_817,N_9977,N_9945);
and UO_818 (O_818,N_9966,N_9998);
nor UO_819 (O_819,N_9916,N_9919);
nor UO_820 (O_820,N_9916,N_9974);
xor UO_821 (O_821,N_9970,N_9929);
xor UO_822 (O_822,N_9931,N_9913);
or UO_823 (O_823,N_9927,N_9998);
xor UO_824 (O_824,N_9906,N_9942);
nand UO_825 (O_825,N_9991,N_9940);
or UO_826 (O_826,N_9957,N_9986);
or UO_827 (O_827,N_9910,N_9907);
or UO_828 (O_828,N_9984,N_9912);
and UO_829 (O_829,N_9919,N_9992);
or UO_830 (O_830,N_9989,N_9969);
and UO_831 (O_831,N_9940,N_9965);
nor UO_832 (O_832,N_9992,N_9979);
and UO_833 (O_833,N_9913,N_9915);
xor UO_834 (O_834,N_9985,N_9977);
nor UO_835 (O_835,N_9908,N_9982);
nand UO_836 (O_836,N_9936,N_9962);
nor UO_837 (O_837,N_9921,N_9908);
nor UO_838 (O_838,N_9975,N_9938);
nand UO_839 (O_839,N_9941,N_9935);
and UO_840 (O_840,N_9957,N_9968);
xor UO_841 (O_841,N_9958,N_9942);
xnor UO_842 (O_842,N_9931,N_9932);
and UO_843 (O_843,N_9949,N_9941);
nand UO_844 (O_844,N_9911,N_9943);
or UO_845 (O_845,N_9935,N_9959);
or UO_846 (O_846,N_9977,N_9949);
nand UO_847 (O_847,N_9975,N_9988);
nor UO_848 (O_848,N_9970,N_9908);
and UO_849 (O_849,N_9973,N_9922);
nor UO_850 (O_850,N_9992,N_9953);
or UO_851 (O_851,N_9986,N_9907);
nor UO_852 (O_852,N_9987,N_9904);
and UO_853 (O_853,N_9943,N_9978);
xor UO_854 (O_854,N_9933,N_9939);
nand UO_855 (O_855,N_9981,N_9963);
and UO_856 (O_856,N_9911,N_9931);
or UO_857 (O_857,N_9912,N_9908);
nand UO_858 (O_858,N_9950,N_9934);
xnor UO_859 (O_859,N_9938,N_9985);
and UO_860 (O_860,N_9942,N_9965);
nand UO_861 (O_861,N_9918,N_9992);
nor UO_862 (O_862,N_9988,N_9968);
nand UO_863 (O_863,N_9971,N_9965);
xor UO_864 (O_864,N_9963,N_9962);
or UO_865 (O_865,N_9908,N_9932);
and UO_866 (O_866,N_9969,N_9906);
and UO_867 (O_867,N_9936,N_9901);
nand UO_868 (O_868,N_9949,N_9948);
nand UO_869 (O_869,N_9933,N_9902);
nand UO_870 (O_870,N_9903,N_9985);
nand UO_871 (O_871,N_9990,N_9967);
nand UO_872 (O_872,N_9913,N_9991);
or UO_873 (O_873,N_9936,N_9944);
xnor UO_874 (O_874,N_9942,N_9962);
and UO_875 (O_875,N_9927,N_9932);
xor UO_876 (O_876,N_9961,N_9982);
nor UO_877 (O_877,N_9920,N_9910);
nor UO_878 (O_878,N_9917,N_9972);
nand UO_879 (O_879,N_9979,N_9980);
nor UO_880 (O_880,N_9999,N_9918);
or UO_881 (O_881,N_9922,N_9904);
nor UO_882 (O_882,N_9920,N_9947);
nor UO_883 (O_883,N_9956,N_9904);
nor UO_884 (O_884,N_9943,N_9903);
xor UO_885 (O_885,N_9911,N_9904);
xnor UO_886 (O_886,N_9966,N_9951);
xnor UO_887 (O_887,N_9941,N_9944);
or UO_888 (O_888,N_9933,N_9927);
or UO_889 (O_889,N_9973,N_9977);
and UO_890 (O_890,N_9964,N_9903);
or UO_891 (O_891,N_9988,N_9940);
and UO_892 (O_892,N_9984,N_9956);
or UO_893 (O_893,N_9978,N_9913);
or UO_894 (O_894,N_9906,N_9989);
or UO_895 (O_895,N_9927,N_9906);
nand UO_896 (O_896,N_9921,N_9993);
nor UO_897 (O_897,N_9936,N_9926);
nand UO_898 (O_898,N_9906,N_9909);
and UO_899 (O_899,N_9946,N_9909);
nor UO_900 (O_900,N_9996,N_9980);
and UO_901 (O_901,N_9988,N_9937);
and UO_902 (O_902,N_9933,N_9969);
or UO_903 (O_903,N_9910,N_9911);
or UO_904 (O_904,N_9972,N_9925);
and UO_905 (O_905,N_9946,N_9997);
and UO_906 (O_906,N_9928,N_9965);
nand UO_907 (O_907,N_9962,N_9921);
nand UO_908 (O_908,N_9965,N_9979);
and UO_909 (O_909,N_9944,N_9909);
nor UO_910 (O_910,N_9946,N_9904);
xnor UO_911 (O_911,N_9929,N_9950);
nor UO_912 (O_912,N_9973,N_9991);
nor UO_913 (O_913,N_9999,N_9951);
nor UO_914 (O_914,N_9954,N_9964);
nand UO_915 (O_915,N_9991,N_9966);
xor UO_916 (O_916,N_9960,N_9988);
or UO_917 (O_917,N_9925,N_9919);
and UO_918 (O_918,N_9930,N_9992);
and UO_919 (O_919,N_9983,N_9947);
nor UO_920 (O_920,N_9908,N_9964);
xnor UO_921 (O_921,N_9971,N_9993);
and UO_922 (O_922,N_9960,N_9994);
xor UO_923 (O_923,N_9902,N_9905);
nand UO_924 (O_924,N_9903,N_9920);
xnor UO_925 (O_925,N_9950,N_9999);
and UO_926 (O_926,N_9983,N_9998);
or UO_927 (O_927,N_9998,N_9950);
or UO_928 (O_928,N_9933,N_9970);
nand UO_929 (O_929,N_9964,N_9923);
nor UO_930 (O_930,N_9940,N_9905);
and UO_931 (O_931,N_9901,N_9923);
xnor UO_932 (O_932,N_9943,N_9951);
nand UO_933 (O_933,N_9921,N_9904);
and UO_934 (O_934,N_9920,N_9962);
or UO_935 (O_935,N_9962,N_9926);
nor UO_936 (O_936,N_9988,N_9954);
xor UO_937 (O_937,N_9968,N_9906);
nand UO_938 (O_938,N_9974,N_9970);
or UO_939 (O_939,N_9920,N_9904);
and UO_940 (O_940,N_9903,N_9987);
and UO_941 (O_941,N_9999,N_9961);
and UO_942 (O_942,N_9938,N_9918);
or UO_943 (O_943,N_9920,N_9965);
nor UO_944 (O_944,N_9961,N_9950);
and UO_945 (O_945,N_9945,N_9993);
or UO_946 (O_946,N_9937,N_9951);
or UO_947 (O_947,N_9957,N_9996);
xnor UO_948 (O_948,N_9904,N_9926);
or UO_949 (O_949,N_9936,N_9911);
or UO_950 (O_950,N_9930,N_9937);
or UO_951 (O_951,N_9977,N_9958);
nand UO_952 (O_952,N_9954,N_9936);
and UO_953 (O_953,N_9927,N_9958);
and UO_954 (O_954,N_9961,N_9929);
or UO_955 (O_955,N_9959,N_9993);
nand UO_956 (O_956,N_9902,N_9958);
nand UO_957 (O_957,N_9916,N_9968);
and UO_958 (O_958,N_9987,N_9998);
xor UO_959 (O_959,N_9925,N_9903);
nor UO_960 (O_960,N_9915,N_9908);
and UO_961 (O_961,N_9944,N_9932);
xor UO_962 (O_962,N_9980,N_9973);
xnor UO_963 (O_963,N_9942,N_9909);
xor UO_964 (O_964,N_9937,N_9947);
and UO_965 (O_965,N_9924,N_9966);
nand UO_966 (O_966,N_9987,N_9947);
or UO_967 (O_967,N_9996,N_9924);
nor UO_968 (O_968,N_9994,N_9952);
xnor UO_969 (O_969,N_9945,N_9975);
xnor UO_970 (O_970,N_9935,N_9900);
xnor UO_971 (O_971,N_9928,N_9950);
xnor UO_972 (O_972,N_9937,N_9906);
nor UO_973 (O_973,N_9949,N_9976);
nand UO_974 (O_974,N_9939,N_9995);
nand UO_975 (O_975,N_9980,N_9942);
and UO_976 (O_976,N_9914,N_9990);
xnor UO_977 (O_977,N_9958,N_9964);
nand UO_978 (O_978,N_9907,N_9985);
nor UO_979 (O_979,N_9914,N_9922);
and UO_980 (O_980,N_9918,N_9932);
and UO_981 (O_981,N_9931,N_9956);
or UO_982 (O_982,N_9958,N_9922);
nand UO_983 (O_983,N_9925,N_9950);
and UO_984 (O_984,N_9935,N_9923);
nand UO_985 (O_985,N_9929,N_9959);
xor UO_986 (O_986,N_9924,N_9937);
or UO_987 (O_987,N_9947,N_9909);
xnor UO_988 (O_988,N_9970,N_9917);
nand UO_989 (O_989,N_9961,N_9910);
xor UO_990 (O_990,N_9955,N_9936);
nor UO_991 (O_991,N_9951,N_9912);
nand UO_992 (O_992,N_9971,N_9955);
xnor UO_993 (O_993,N_9981,N_9917);
or UO_994 (O_994,N_9963,N_9988);
and UO_995 (O_995,N_9936,N_9999);
and UO_996 (O_996,N_9992,N_9963);
nor UO_997 (O_997,N_9990,N_9959);
xor UO_998 (O_998,N_9962,N_9916);
xnor UO_999 (O_999,N_9964,N_9978);
and UO_1000 (O_1000,N_9995,N_9910);
nand UO_1001 (O_1001,N_9941,N_9982);
xnor UO_1002 (O_1002,N_9940,N_9961);
nor UO_1003 (O_1003,N_9947,N_9976);
xnor UO_1004 (O_1004,N_9940,N_9929);
or UO_1005 (O_1005,N_9994,N_9906);
and UO_1006 (O_1006,N_9950,N_9937);
and UO_1007 (O_1007,N_9953,N_9938);
or UO_1008 (O_1008,N_9964,N_9932);
and UO_1009 (O_1009,N_9933,N_9917);
nor UO_1010 (O_1010,N_9986,N_9967);
and UO_1011 (O_1011,N_9937,N_9929);
or UO_1012 (O_1012,N_9965,N_9948);
xnor UO_1013 (O_1013,N_9902,N_9912);
and UO_1014 (O_1014,N_9987,N_9971);
and UO_1015 (O_1015,N_9936,N_9951);
or UO_1016 (O_1016,N_9924,N_9989);
and UO_1017 (O_1017,N_9917,N_9971);
nor UO_1018 (O_1018,N_9928,N_9947);
nor UO_1019 (O_1019,N_9980,N_9910);
xnor UO_1020 (O_1020,N_9904,N_9965);
nor UO_1021 (O_1021,N_9980,N_9986);
nor UO_1022 (O_1022,N_9972,N_9915);
and UO_1023 (O_1023,N_9970,N_9945);
nor UO_1024 (O_1024,N_9988,N_9934);
nand UO_1025 (O_1025,N_9910,N_9944);
nor UO_1026 (O_1026,N_9962,N_9911);
or UO_1027 (O_1027,N_9959,N_9997);
nor UO_1028 (O_1028,N_9971,N_9975);
and UO_1029 (O_1029,N_9988,N_9950);
and UO_1030 (O_1030,N_9936,N_9957);
or UO_1031 (O_1031,N_9932,N_9953);
or UO_1032 (O_1032,N_9978,N_9970);
xnor UO_1033 (O_1033,N_9928,N_9904);
xor UO_1034 (O_1034,N_9941,N_9966);
nand UO_1035 (O_1035,N_9953,N_9919);
nand UO_1036 (O_1036,N_9958,N_9984);
and UO_1037 (O_1037,N_9940,N_9910);
or UO_1038 (O_1038,N_9927,N_9941);
nor UO_1039 (O_1039,N_9970,N_9958);
nand UO_1040 (O_1040,N_9964,N_9936);
nor UO_1041 (O_1041,N_9910,N_9974);
xnor UO_1042 (O_1042,N_9954,N_9904);
nor UO_1043 (O_1043,N_9993,N_9926);
nor UO_1044 (O_1044,N_9912,N_9903);
nor UO_1045 (O_1045,N_9981,N_9937);
xor UO_1046 (O_1046,N_9976,N_9924);
nor UO_1047 (O_1047,N_9963,N_9929);
and UO_1048 (O_1048,N_9964,N_9957);
or UO_1049 (O_1049,N_9919,N_9954);
nand UO_1050 (O_1050,N_9959,N_9991);
nand UO_1051 (O_1051,N_9927,N_9904);
xor UO_1052 (O_1052,N_9995,N_9960);
xnor UO_1053 (O_1053,N_9932,N_9917);
nor UO_1054 (O_1054,N_9971,N_9902);
nor UO_1055 (O_1055,N_9935,N_9940);
xnor UO_1056 (O_1056,N_9906,N_9972);
and UO_1057 (O_1057,N_9994,N_9927);
nor UO_1058 (O_1058,N_9927,N_9920);
nand UO_1059 (O_1059,N_9919,N_9984);
and UO_1060 (O_1060,N_9991,N_9928);
nand UO_1061 (O_1061,N_9930,N_9940);
and UO_1062 (O_1062,N_9901,N_9969);
and UO_1063 (O_1063,N_9952,N_9928);
nand UO_1064 (O_1064,N_9990,N_9994);
or UO_1065 (O_1065,N_9967,N_9998);
nand UO_1066 (O_1066,N_9985,N_9970);
or UO_1067 (O_1067,N_9997,N_9978);
nand UO_1068 (O_1068,N_9913,N_9928);
nand UO_1069 (O_1069,N_9920,N_9960);
xnor UO_1070 (O_1070,N_9919,N_9913);
xor UO_1071 (O_1071,N_9964,N_9991);
and UO_1072 (O_1072,N_9931,N_9957);
and UO_1073 (O_1073,N_9952,N_9945);
xor UO_1074 (O_1074,N_9997,N_9936);
and UO_1075 (O_1075,N_9910,N_9923);
nor UO_1076 (O_1076,N_9909,N_9936);
xor UO_1077 (O_1077,N_9908,N_9953);
and UO_1078 (O_1078,N_9939,N_9946);
xor UO_1079 (O_1079,N_9934,N_9982);
nand UO_1080 (O_1080,N_9943,N_9939);
and UO_1081 (O_1081,N_9959,N_9986);
nand UO_1082 (O_1082,N_9967,N_9995);
and UO_1083 (O_1083,N_9933,N_9912);
nand UO_1084 (O_1084,N_9991,N_9979);
nor UO_1085 (O_1085,N_9935,N_9926);
and UO_1086 (O_1086,N_9969,N_9982);
and UO_1087 (O_1087,N_9996,N_9908);
xnor UO_1088 (O_1088,N_9965,N_9976);
xor UO_1089 (O_1089,N_9915,N_9996);
or UO_1090 (O_1090,N_9941,N_9975);
or UO_1091 (O_1091,N_9994,N_9957);
xor UO_1092 (O_1092,N_9943,N_9906);
and UO_1093 (O_1093,N_9903,N_9989);
nor UO_1094 (O_1094,N_9999,N_9967);
and UO_1095 (O_1095,N_9958,N_9910);
xor UO_1096 (O_1096,N_9958,N_9909);
and UO_1097 (O_1097,N_9990,N_9929);
and UO_1098 (O_1098,N_9959,N_9950);
and UO_1099 (O_1099,N_9980,N_9992);
xor UO_1100 (O_1100,N_9976,N_9913);
or UO_1101 (O_1101,N_9970,N_9966);
nor UO_1102 (O_1102,N_9971,N_9929);
nor UO_1103 (O_1103,N_9998,N_9952);
nand UO_1104 (O_1104,N_9923,N_9912);
nor UO_1105 (O_1105,N_9958,N_9988);
nand UO_1106 (O_1106,N_9977,N_9925);
nand UO_1107 (O_1107,N_9942,N_9989);
or UO_1108 (O_1108,N_9993,N_9927);
or UO_1109 (O_1109,N_9965,N_9975);
xnor UO_1110 (O_1110,N_9977,N_9982);
nor UO_1111 (O_1111,N_9946,N_9996);
and UO_1112 (O_1112,N_9926,N_9901);
nand UO_1113 (O_1113,N_9932,N_9954);
xor UO_1114 (O_1114,N_9922,N_9991);
nand UO_1115 (O_1115,N_9997,N_9909);
or UO_1116 (O_1116,N_9936,N_9906);
and UO_1117 (O_1117,N_9938,N_9906);
or UO_1118 (O_1118,N_9977,N_9972);
nor UO_1119 (O_1119,N_9911,N_9940);
or UO_1120 (O_1120,N_9947,N_9942);
xnor UO_1121 (O_1121,N_9918,N_9914);
or UO_1122 (O_1122,N_9955,N_9951);
nand UO_1123 (O_1123,N_9981,N_9908);
or UO_1124 (O_1124,N_9997,N_9995);
xor UO_1125 (O_1125,N_9927,N_9999);
xnor UO_1126 (O_1126,N_9974,N_9931);
and UO_1127 (O_1127,N_9982,N_9919);
nor UO_1128 (O_1128,N_9958,N_9930);
nor UO_1129 (O_1129,N_9945,N_9907);
nand UO_1130 (O_1130,N_9980,N_9927);
and UO_1131 (O_1131,N_9954,N_9967);
nor UO_1132 (O_1132,N_9928,N_9983);
xnor UO_1133 (O_1133,N_9934,N_9948);
or UO_1134 (O_1134,N_9975,N_9992);
or UO_1135 (O_1135,N_9975,N_9967);
and UO_1136 (O_1136,N_9930,N_9926);
xnor UO_1137 (O_1137,N_9956,N_9964);
nand UO_1138 (O_1138,N_9956,N_9998);
or UO_1139 (O_1139,N_9970,N_9975);
and UO_1140 (O_1140,N_9969,N_9967);
or UO_1141 (O_1141,N_9997,N_9942);
or UO_1142 (O_1142,N_9924,N_9994);
and UO_1143 (O_1143,N_9996,N_9912);
or UO_1144 (O_1144,N_9936,N_9968);
nand UO_1145 (O_1145,N_9986,N_9958);
or UO_1146 (O_1146,N_9936,N_9952);
nand UO_1147 (O_1147,N_9924,N_9990);
nor UO_1148 (O_1148,N_9915,N_9988);
nand UO_1149 (O_1149,N_9943,N_9971);
xor UO_1150 (O_1150,N_9965,N_9981);
or UO_1151 (O_1151,N_9928,N_9959);
xor UO_1152 (O_1152,N_9934,N_9904);
or UO_1153 (O_1153,N_9976,N_9931);
or UO_1154 (O_1154,N_9945,N_9973);
nand UO_1155 (O_1155,N_9954,N_9958);
xnor UO_1156 (O_1156,N_9991,N_9981);
xor UO_1157 (O_1157,N_9955,N_9969);
and UO_1158 (O_1158,N_9977,N_9916);
or UO_1159 (O_1159,N_9920,N_9952);
nor UO_1160 (O_1160,N_9970,N_9950);
nand UO_1161 (O_1161,N_9938,N_9964);
or UO_1162 (O_1162,N_9912,N_9920);
xnor UO_1163 (O_1163,N_9988,N_9973);
xor UO_1164 (O_1164,N_9944,N_9994);
and UO_1165 (O_1165,N_9966,N_9993);
nor UO_1166 (O_1166,N_9987,N_9980);
and UO_1167 (O_1167,N_9929,N_9982);
xnor UO_1168 (O_1168,N_9948,N_9906);
nor UO_1169 (O_1169,N_9986,N_9941);
and UO_1170 (O_1170,N_9933,N_9972);
nand UO_1171 (O_1171,N_9948,N_9944);
nand UO_1172 (O_1172,N_9913,N_9952);
nand UO_1173 (O_1173,N_9935,N_9934);
xnor UO_1174 (O_1174,N_9959,N_9934);
and UO_1175 (O_1175,N_9972,N_9902);
nand UO_1176 (O_1176,N_9997,N_9993);
nand UO_1177 (O_1177,N_9957,N_9958);
nor UO_1178 (O_1178,N_9996,N_9933);
or UO_1179 (O_1179,N_9999,N_9923);
nor UO_1180 (O_1180,N_9914,N_9947);
or UO_1181 (O_1181,N_9999,N_9954);
or UO_1182 (O_1182,N_9995,N_9940);
nor UO_1183 (O_1183,N_9964,N_9985);
nor UO_1184 (O_1184,N_9952,N_9909);
xor UO_1185 (O_1185,N_9943,N_9983);
and UO_1186 (O_1186,N_9981,N_9979);
nor UO_1187 (O_1187,N_9911,N_9995);
and UO_1188 (O_1188,N_9913,N_9949);
and UO_1189 (O_1189,N_9943,N_9980);
or UO_1190 (O_1190,N_9943,N_9941);
nor UO_1191 (O_1191,N_9978,N_9938);
and UO_1192 (O_1192,N_9964,N_9910);
xnor UO_1193 (O_1193,N_9918,N_9913);
nand UO_1194 (O_1194,N_9955,N_9909);
or UO_1195 (O_1195,N_9952,N_9925);
and UO_1196 (O_1196,N_9930,N_9973);
and UO_1197 (O_1197,N_9982,N_9994);
xnor UO_1198 (O_1198,N_9937,N_9997);
xnor UO_1199 (O_1199,N_9990,N_9915);
nor UO_1200 (O_1200,N_9917,N_9907);
xnor UO_1201 (O_1201,N_9938,N_9950);
xor UO_1202 (O_1202,N_9980,N_9950);
and UO_1203 (O_1203,N_9969,N_9948);
or UO_1204 (O_1204,N_9912,N_9939);
nand UO_1205 (O_1205,N_9938,N_9907);
and UO_1206 (O_1206,N_9975,N_9922);
nor UO_1207 (O_1207,N_9981,N_9918);
nand UO_1208 (O_1208,N_9921,N_9990);
and UO_1209 (O_1209,N_9907,N_9914);
and UO_1210 (O_1210,N_9916,N_9963);
or UO_1211 (O_1211,N_9972,N_9999);
xnor UO_1212 (O_1212,N_9978,N_9914);
xnor UO_1213 (O_1213,N_9916,N_9958);
xor UO_1214 (O_1214,N_9996,N_9954);
xnor UO_1215 (O_1215,N_9910,N_9908);
xor UO_1216 (O_1216,N_9919,N_9951);
nand UO_1217 (O_1217,N_9971,N_9945);
and UO_1218 (O_1218,N_9920,N_9967);
or UO_1219 (O_1219,N_9913,N_9956);
and UO_1220 (O_1220,N_9900,N_9904);
and UO_1221 (O_1221,N_9986,N_9905);
xnor UO_1222 (O_1222,N_9941,N_9977);
nand UO_1223 (O_1223,N_9982,N_9923);
xor UO_1224 (O_1224,N_9975,N_9909);
nor UO_1225 (O_1225,N_9905,N_9992);
and UO_1226 (O_1226,N_9901,N_9909);
nor UO_1227 (O_1227,N_9986,N_9923);
nor UO_1228 (O_1228,N_9938,N_9930);
and UO_1229 (O_1229,N_9929,N_9960);
xnor UO_1230 (O_1230,N_9922,N_9987);
and UO_1231 (O_1231,N_9997,N_9979);
and UO_1232 (O_1232,N_9933,N_9997);
nor UO_1233 (O_1233,N_9994,N_9901);
xor UO_1234 (O_1234,N_9955,N_9983);
xnor UO_1235 (O_1235,N_9933,N_9954);
or UO_1236 (O_1236,N_9978,N_9904);
or UO_1237 (O_1237,N_9928,N_9942);
nor UO_1238 (O_1238,N_9913,N_9995);
or UO_1239 (O_1239,N_9919,N_9964);
and UO_1240 (O_1240,N_9966,N_9988);
or UO_1241 (O_1241,N_9933,N_9906);
nand UO_1242 (O_1242,N_9993,N_9980);
xnor UO_1243 (O_1243,N_9975,N_9969);
nand UO_1244 (O_1244,N_9981,N_9974);
and UO_1245 (O_1245,N_9915,N_9942);
nand UO_1246 (O_1246,N_9939,N_9901);
xor UO_1247 (O_1247,N_9918,N_9965);
or UO_1248 (O_1248,N_9984,N_9993);
xnor UO_1249 (O_1249,N_9907,N_9920);
and UO_1250 (O_1250,N_9974,N_9909);
nor UO_1251 (O_1251,N_9947,N_9986);
or UO_1252 (O_1252,N_9901,N_9986);
and UO_1253 (O_1253,N_9919,N_9999);
nand UO_1254 (O_1254,N_9997,N_9934);
nor UO_1255 (O_1255,N_9922,N_9948);
nand UO_1256 (O_1256,N_9937,N_9944);
nor UO_1257 (O_1257,N_9961,N_9970);
or UO_1258 (O_1258,N_9915,N_9956);
nor UO_1259 (O_1259,N_9943,N_9982);
and UO_1260 (O_1260,N_9960,N_9996);
nor UO_1261 (O_1261,N_9902,N_9951);
nand UO_1262 (O_1262,N_9990,N_9971);
or UO_1263 (O_1263,N_9933,N_9920);
nor UO_1264 (O_1264,N_9964,N_9929);
nand UO_1265 (O_1265,N_9958,N_9955);
and UO_1266 (O_1266,N_9956,N_9999);
xor UO_1267 (O_1267,N_9937,N_9942);
or UO_1268 (O_1268,N_9941,N_9984);
nand UO_1269 (O_1269,N_9931,N_9909);
and UO_1270 (O_1270,N_9970,N_9914);
xor UO_1271 (O_1271,N_9920,N_9946);
nand UO_1272 (O_1272,N_9958,N_9906);
nand UO_1273 (O_1273,N_9992,N_9984);
nand UO_1274 (O_1274,N_9940,N_9975);
or UO_1275 (O_1275,N_9916,N_9972);
nand UO_1276 (O_1276,N_9901,N_9937);
nor UO_1277 (O_1277,N_9939,N_9988);
or UO_1278 (O_1278,N_9991,N_9960);
nand UO_1279 (O_1279,N_9959,N_9947);
nand UO_1280 (O_1280,N_9960,N_9910);
xnor UO_1281 (O_1281,N_9953,N_9984);
and UO_1282 (O_1282,N_9912,N_9983);
or UO_1283 (O_1283,N_9946,N_9978);
and UO_1284 (O_1284,N_9958,N_9931);
xnor UO_1285 (O_1285,N_9914,N_9919);
xnor UO_1286 (O_1286,N_9978,N_9935);
and UO_1287 (O_1287,N_9934,N_9962);
nor UO_1288 (O_1288,N_9985,N_9914);
xor UO_1289 (O_1289,N_9970,N_9939);
xor UO_1290 (O_1290,N_9972,N_9936);
nor UO_1291 (O_1291,N_9907,N_9900);
xnor UO_1292 (O_1292,N_9901,N_9918);
or UO_1293 (O_1293,N_9921,N_9932);
xnor UO_1294 (O_1294,N_9991,N_9949);
xor UO_1295 (O_1295,N_9924,N_9906);
xnor UO_1296 (O_1296,N_9955,N_9977);
and UO_1297 (O_1297,N_9939,N_9962);
and UO_1298 (O_1298,N_9934,N_9917);
or UO_1299 (O_1299,N_9900,N_9994);
or UO_1300 (O_1300,N_9960,N_9963);
nor UO_1301 (O_1301,N_9915,N_9933);
nor UO_1302 (O_1302,N_9954,N_9971);
or UO_1303 (O_1303,N_9909,N_9933);
nand UO_1304 (O_1304,N_9975,N_9911);
xor UO_1305 (O_1305,N_9953,N_9965);
xnor UO_1306 (O_1306,N_9912,N_9930);
or UO_1307 (O_1307,N_9968,N_9948);
nor UO_1308 (O_1308,N_9954,N_9990);
and UO_1309 (O_1309,N_9997,N_9925);
xor UO_1310 (O_1310,N_9970,N_9919);
nor UO_1311 (O_1311,N_9937,N_9909);
nor UO_1312 (O_1312,N_9982,N_9954);
nand UO_1313 (O_1313,N_9919,N_9902);
xnor UO_1314 (O_1314,N_9953,N_9942);
or UO_1315 (O_1315,N_9992,N_9960);
and UO_1316 (O_1316,N_9983,N_9957);
xor UO_1317 (O_1317,N_9982,N_9944);
nand UO_1318 (O_1318,N_9917,N_9966);
or UO_1319 (O_1319,N_9930,N_9962);
nor UO_1320 (O_1320,N_9949,N_9915);
nor UO_1321 (O_1321,N_9903,N_9944);
and UO_1322 (O_1322,N_9929,N_9918);
xor UO_1323 (O_1323,N_9908,N_9917);
and UO_1324 (O_1324,N_9918,N_9921);
or UO_1325 (O_1325,N_9982,N_9902);
or UO_1326 (O_1326,N_9952,N_9915);
nand UO_1327 (O_1327,N_9953,N_9966);
and UO_1328 (O_1328,N_9981,N_9915);
and UO_1329 (O_1329,N_9979,N_9913);
xor UO_1330 (O_1330,N_9973,N_9942);
or UO_1331 (O_1331,N_9996,N_9970);
nand UO_1332 (O_1332,N_9996,N_9934);
or UO_1333 (O_1333,N_9909,N_9905);
nor UO_1334 (O_1334,N_9974,N_9951);
xnor UO_1335 (O_1335,N_9956,N_9920);
and UO_1336 (O_1336,N_9903,N_9981);
or UO_1337 (O_1337,N_9998,N_9943);
and UO_1338 (O_1338,N_9915,N_9986);
xnor UO_1339 (O_1339,N_9932,N_9960);
nor UO_1340 (O_1340,N_9940,N_9974);
and UO_1341 (O_1341,N_9973,N_9994);
xnor UO_1342 (O_1342,N_9911,N_9933);
nor UO_1343 (O_1343,N_9948,N_9979);
xor UO_1344 (O_1344,N_9923,N_9970);
nand UO_1345 (O_1345,N_9979,N_9944);
nor UO_1346 (O_1346,N_9996,N_9921);
and UO_1347 (O_1347,N_9974,N_9952);
and UO_1348 (O_1348,N_9954,N_9923);
xnor UO_1349 (O_1349,N_9924,N_9946);
nor UO_1350 (O_1350,N_9985,N_9940);
xor UO_1351 (O_1351,N_9976,N_9907);
nand UO_1352 (O_1352,N_9928,N_9921);
and UO_1353 (O_1353,N_9930,N_9966);
nor UO_1354 (O_1354,N_9965,N_9933);
xnor UO_1355 (O_1355,N_9933,N_9980);
xnor UO_1356 (O_1356,N_9967,N_9941);
nor UO_1357 (O_1357,N_9960,N_9936);
nand UO_1358 (O_1358,N_9908,N_9945);
nor UO_1359 (O_1359,N_9925,N_9904);
nand UO_1360 (O_1360,N_9967,N_9917);
nor UO_1361 (O_1361,N_9909,N_9923);
nand UO_1362 (O_1362,N_9988,N_9949);
and UO_1363 (O_1363,N_9959,N_9958);
or UO_1364 (O_1364,N_9947,N_9960);
or UO_1365 (O_1365,N_9950,N_9969);
or UO_1366 (O_1366,N_9965,N_9991);
xnor UO_1367 (O_1367,N_9933,N_9976);
or UO_1368 (O_1368,N_9939,N_9949);
or UO_1369 (O_1369,N_9990,N_9913);
and UO_1370 (O_1370,N_9981,N_9947);
nor UO_1371 (O_1371,N_9978,N_9975);
and UO_1372 (O_1372,N_9927,N_9924);
xor UO_1373 (O_1373,N_9993,N_9952);
xor UO_1374 (O_1374,N_9971,N_9930);
xnor UO_1375 (O_1375,N_9939,N_9959);
xor UO_1376 (O_1376,N_9995,N_9903);
nand UO_1377 (O_1377,N_9927,N_9937);
nand UO_1378 (O_1378,N_9907,N_9949);
or UO_1379 (O_1379,N_9975,N_9914);
and UO_1380 (O_1380,N_9909,N_9918);
or UO_1381 (O_1381,N_9922,N_9964);
or UO_1382 (O_1382,N_9936,N_9942);
nor UO_1383 (O_1383,N_9949,N_9998);
and UO_1384 (O_1384,N_9997,N_9968);
and UO_1385 (O_1385,N_9933,N_9931);
nor UO_1386 (O_1386,N_9973,N_9928);
xnor UO_1387 (O_1387,N_9953,N_9901);
nand UO_1388 (O_1388,N_9994,N_9983);
xnor UO_1389 (O_1389,N_9993,N_9907);
nor UO_1390 (O_1390,N_9981,N_9938);
xor UO_1391 (O_1391,N_9961,N_9923);
or UO_1392 (O_1392,N_9920,N_9971);
xor UO_1393 (O_1393,N_9931,N_9902);
xor UO_1394 (O_1394,N_9916,N_9922);
nand UO_1395 (O_1395,N_9978,N_9939);
or UO_1396 (O_1396,N_9949,N_9916);
xor UO_1397 (O_1397,N_9945,N_9934);
or UO_1398 (O_1398,N_9965,N_9911);
nand UO_1399 (O_1399,N_9961,N_9900);
nand UO_1400 (O_1400,N_9917,N_9955);
nor UO_1401 (O_1401,N_9933,N_9901);
and UO_1402 (O_1402,N_9984,N_9924);
nor UO_1403 (O_1403,N_9968,N_9961);
xnor UO_1404 (O_1404,N_9948,N_9903);
nor UO_1405 (O_1405,N_9960,N_9953);
and UO_1406 (O_1406,N_9922,N_9982);
xor UO_1407 (O_1407,N_9922,N_9925);
nor UO_1408 (O_1408,N_9901,N_9988);
or UO_1409 (O_1409,N_9918,N_9927);
nand UO_1410 (O_1410,N_9955,N_9981);
xor UO_1411 (O_1411,N_9905,N_9910);
xnor UO_1412 (O_1412,N_9910,N_9928);
and UO_1413 (O_1413,N_9944,N_9925);
and UO_1414 (O_1414,N_9922,N_9936);
or UO_1415 (O_1415,N_9908,N_9900);
or UO_1416 (O_1416,N_9997,N_9926);
nor UO_1417 (O_1417,N_9940,N_9912);
nor UO_1418 (O_1418,N_9917,N_9923);
or UO_1419 (O_1419,N_9960,N_9972);
xor UO_1420 (O_1420,N_9980,N_9925);
xnor UO_1421 (O_1421,N_9948,N_9989);
xnor UO_1422 (O_1422,N_9913,N_9998);
xor UO_1423 (O_1423,N_9995,N_9914);
xnor UO_1424 (O_1424,N_9979,N_9975);
nor UO_1425 (O_1425,N_9964,N_9930);
or UO_1426 (O_1426,N_9914,N_9954);
xor UO_1427 (O_1427,N_9989,N_9949);
nor UO_1428 (O_1428,N_9967,N_9901);
nand UO_1429 (O_1429,N_9932,N_9909);
and UO_1430 (O_1430,N_9943,N_9910);
and UO_1431 (O_1431,N_9979,N_9941);
xnor UO_1432 (O_1432,N_9933,N_9966);
nand UO_1433 (O_1433,N_9990,N_9911);
nor UO_1434 (O_1434,N_9908,N_9940);
and UO_1435 (O_1435,N_9937,N_9987);
and UO_1436 (O_1436,N_9995,N_9970);
and UO_1437 (O_1437,N_9908,N_9961);
and UO_1438 (O_1438,N_9903,N_9960);
nand UO_1439 (O_1439,N_9926,N_9955);
and UO_1440 (O_1440,N_9950,N_9983);
xnor UO_1441 (O_1441,N_9963,N_9990);
nand UO_1442 (O_1442,N_9967,N_9968);
or UO_1443 (O_1443,N_9958,N_9943);
nand UO_1444 (O_1444,N_9970,N_9969);
nor UO_1445 (O_1445,N_9990,N_9998);
nor UO_1446 (O_1446,N_9991,N_9933);
nand UO_1447 (O_1447,N_9995,N_9991);
xor UO_1448 (O_1448,N_9996,N_9900);
xnor UO_1449 (O_1449,N_9945,N_9932);
nor UO_1450 (O_1450,N_9965,N_9934);
nand UO_1451 (O_1451,N_9980,N_9902);
and UO_1452 (O_1452,N_9925,N_9983);
or UO_1453 (O_1453,N_9942,N_9970);
nor UO_1454 (O_1454,N_9917,N_9906);
or UO_1455 (O_1455,N_9950,N_9947);
nand UO_1456 (O_1456,N_9997,N_9917);
nor UO_1457 (O_1457,N_9938,N_9990);
or UO_1458 (O_1458,N_9998,N_9979);
xnor UO_1459 (O_1459,N_9928,N_9933);
xnor UO_1460 (O_1460,N_9990,N_9936);
xor UO_1461 (O_1461,N_9916,N_9950);
or UO_1462 (O_1462,N_9998,N_9938);
or UO_1463 (O_1463,N_9992,N_9988);
xnor UO_1464 (O_1464,N_9971,N_9973);
nand UO_1465 (O_1465,N_9962,N_9996);
xnor UO_1466 (O_1466,N_9944,N_9902);
or UO_1467 (O_1467,N_9948,N_9942);
xnor UO_1468 (O_1468,N_9987,N_9923);
xnor UO_1469 (O_1469,N_9945,N_9994);
xnor UO_1470 (O_1470,N_9903,N_9913);
and UO_1471 (O_1471,N_9985,N_9941);
or UO_1472 (O_1472,N_9929,N_9932);
nor UO_1473 (O_1473,N_9989,N_9991);
nor UO_1474 (O_1474,N_9982,N_9950);
nand UO_1475 (O_1475,N_9962,N_9973);
nand UO_1476 (O_1476,N_9950,N_9951);
nor UO_1477 (O_1477,N_9945,N_9983);
nor UO_1478 (O_1478,N_9936,N_9915);
nand UO_1479 (O_1479,N_9944,N_9959);
or UO_1480 (O_1480,N_9950,N_9945);
xnor UO_1481 (O_1481,N_9920,N_9918);
and UO_1482 (O_1482,N_9952,N_9906);
and UO_1483 (O_1483,N_9943,N_9948);
nor UO_1484 (O_1484,N_9905,N_9965);
or UO_1485 (O_1485,N_9955,N_9929);
or UO_1486 (O_1486,N_9967,N_9991);
or UO_1487 (O_1487,N_9988,N_9991);
and UO_1488 (O_1488,N_9952,N_9984);
or UO_1489 (O_1489,N_9931,N_9927);
and UO_1490 (O_1490,N_9908,N_9950);
xnor UO_1491 (O_1491,N_9989,N_9988);
or UO_1492 (O_1492,N_9933,N_9938);
nor UO_1493 (O_1493,N_9959,N_9973);
nand UO_1494 (O_1494,N_9918,N_9984);
nor UO_1495 (O_1495,N_9941,N_9928);
and UO_1496 (O_1496,N_9928,N_9967);
or UO_1497 (O_1497,N_9931,N_9949);
or UO_1498 (O_1498,N_9983,N_9969);
nor UO_1499 (O_1499,N_9932,N_9943);
endmodule